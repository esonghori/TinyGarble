
module MUX_N1024_0 ( A, B, S, O );
  input [1023:0] A;
  input [1023:0] B;
  output [1023:0] O;
  input S;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048;

  XOR U1 ( .A(A[9]), .B(n1), .Z(O[9]) );
  AND U2 ( .A(S), .B(n2), .Z(n1) );
  XOR U3 ( .A(B[9]), .B(A[9]), .Z(n2) );
  XOR U4 ( .A(A[99]), .B(n3), .Z(O[99]) );
  AND U5 ( .A(S), .B(n4), .Z(n3) );
  XOR U6 ( .A(B[99]), .B(A[99]), .Z(n4) );
  XOR U7 ( .A(A[999]), .B(n5), .Z(O[999]) );
  AND U8 ( .A(S), .B(n6), .Z(n5) );
  XOR U9 ( .A(B[999]), .B(A[999]), .Z(n6) );
  XOR U10 ( .A(A[998]), .B(n7), .Z(O[998]) );
  AND U11 ( .A(S), .B(n8), .Z(n7) );
  XOR U12 ( .A(B[998]), .B(A[998]), .Z(n8) );
  XOR U13 ( .A(A[997]), .B(n9), .Z(O[997]) );
  AND U14 ( .A(S), .B(n10), .Z(n9) );
  XOR U15 ( .A(B[997]), .B(A[997]), .Z(n10) );
  XOR U16 ( .A(A[996]), .B(n11), .Z(O[996]) );
  AND U17 ( .A(S), .B(n12), .Z(n11) );
  XOR U18 ( .A(B[996]), .B(A[996]), .Z(n12) );
  XOR U19 ( .A(A[995]), .B(n13), .Z(O[995]) );
  AND U20 ( .A(S), .B(n14), .Z(n13) );
  XOR U21 ( .A(B[995]), .B(A[995]), .Z(n14) );
  XOR U22 ( .A(A[994]), .B(n15), .Z(O[994]) );
  AND U23 ( .A(S), .B(n16), .Z(n15) );
  XOR U24 ( .A(B[994]), .B(A[994]), .Z(n16) );
  XOR U25 ( .A(A[993]), .B(n17), .Z(O[993]) );
  AND U26 ( .A(S), .B(n18), .Z(n17) );
  XOR U27 ( .A(B[993]), .B(A[993]), .Z(n18) );
  XOR U28 ( .A(A[992]), .B(n19), .Z(O[992]) );
  AND U29 ( .A(S), .B(n20), .Z(n19) );
  XOR U30 ( .A(B[992]), .B(A[992]), .Z(n20) );
  XOR U31 ( .A(A[991]), .B(n21), .Z(O[991]) );
  AND U32 ( .A(S), .B(n22), .Z(n21) );
  XOR U33 ( .A(B[991]), .B(A[991]), .Z(n22) );
  XOR U34 ( .A(A[990]), .B(n23), .Z(O[990]) );
  AND U35 ( .A(S), .B(n24), .Z(n23) );
  XOR U36 ( .A(B[990]), .B(A[990]), .Z(n24) );
  XOR U37 ( .A(A[98]), .B(n25), .Z(O[98]) );
  AND U38 ( .A(S), .B(n26), .Z(n25) );
  XOR U39 ( .A(B[98]), .B(A[98]), .Z(n26) );
  XOR U40 ( .A(A[989]), .B(n27), .Z(O[989]) );
  AND U41 ( .A(S), .B(n28), .Z(n27) );
  XOR U42 ( .A(B[989]), .B(A[989]), .Z(n28) );
  XOR U43 ( .A(A[988]), .B(n29), .Z(O[988]) );
  AND U44 ( .A(S), .B(n30), .Z(n29) );
  XOR U45 ( .A(B[988]), .B(A[988]), .Z(n30) );
  XOR U46 ( .A(A[987]), .B(n31), .Z(O[987]) );
  AND U47 ( .A(S), .B(n32), .Z(n31) );
  XOR U48 ( .A(B[987]), .B(A[987]), .Z(n32) );
  XOR U49 ( .A(A[986]), .B(n33), .Z(O[986]) );
  AND U50 ( .A(S), .B(n34), .Z(n33) );
  XOR U51 ( .A(B[986]), .B(A[986]), .Z(n34) );
  XOR U52 ( .A(A[985]), .B(n35), .Z(O[985]) );
  AND U53 ( .A(S), .B(n36), .Z(n35) );
  XOR U54 ( .A(B[985]), .B(A[985]), .Z(n36) );
  XOR U55 ( .A(A[984]), .B(n37), .Z(O[984]) );
  AND U56 ( .A(S), .B(n38), .Z(n37) );
  XOR U57 ( .A(B[984]), .B(A[984]), .Z(n38) );
  XOR U58 ( .A(A[983]), .B(n39), .Z(O[983]) );
  AND U59 ( .A(S), .B(n40), .Z(n39) );
  XOR U60 ( .A(B[983]), .B(A[983]), .Z(n40) );
  XOR U61 ( .A(A[982]), .B(n41), .Z(O[982]) );
  AND U62 ( .A(S), .B(n42), .Z(n41) );
  XOR U63 ( .A(B[982]), .B(A[982]), .Z(n42) );
  XOR U64 ( .A(A[981]), .B(n43), .Z(O[981]) );
  AND U65 ( .A(S), .B(n44), .Z(n43) );
  XOR U66 ( .A(B[981]), .B(A[981]), .Z(n44) );
  XOR U67 ( .A(A[980]), .B(n45), .Z(O[980]) );
  AND U68 ( .A(S), .B(n46), .Z(n45) );
  XOR U69 ( .A(B[980]), .B(A[980]), .Z(n46) );
  XOR U70 ( .A(A[97]), .B(n47), .Z(O[97]) );
  AND U71 ( .A(S), .B(n48), .Z(n47) );
  XOR U72 ( .A(B[97]), .B(A[97]), .Z(n48) );
  XOR U73 ( .A(A[979]), .B(n49), .Z(O[979]) );
  AND U74 ( .A(S), .B(n50), .Z(n49) );
  XOR U75 ( .A(B[979]), .B(A[979]), .Z(n50) );
  XOR U76 ( .A(A[978]), .B(n51), .Z(O[978]) );
  AND U77 ( .A(S), .B(n52), .Z(n51) );
  XOR U78 ( .A(B[978]), .B(A[978]), .Z(n52) );
  XOR U79 ( .A(A[977]), .B(n53), .Z(O[977]) );
  AND U80 ( .A(S), .B(n54), .Z(n53) );
  XOR U81 ( .A(B[977]), .B(A[977]), .Z(n54) );
  XOR U82 ( .A(A[976]), .B(n55), .Z(O[976]) );
  AND U83 ( .A(S), .B(n56), .Z(n55) );
  XOR U84 ( .A(B[976]), .B(A[976]), .Z(n56) );
  XOR U85 ( .A(A[975]), .B(n57), .Z(O[975]) );
  AND U86 ( .A(S), .B(n58), .Z(n57) );
  XOR U87 ( .A(B[975]), .B(A[975]), .Z(n58) );
  XOR U88 ( .A(A[974]), .B(n59), .Z(O[974]) );
  AND U89 ( .A(S), .B(n60), .Z(n59) );
  XOR U90 ( .A(B[974]), .B(A[974]), .Z(n60) );
  XOR U91 ( .A(A[973]), .B(n61), .Z(O[973]) );
  AND U92 ( .A(S), .B(n62), .Z(n61) );
  XOR U93 ( .A(B[973]), .B(A[973]), .Z(n62) );
  XOR U94 ( .A(A[972]), .B(n63), .Z(O[972]) );
  AND U95 ( .A(S), .B(n64), .Z(n63) );
  XOR U96 ( .A(B[972]), .B(A[972]), .Z(n64) );
  XOR U97 ( .A(A[971]), .B(n65), .Z(O[971]) );
  AND U98 ( .A(S), .B(n66), .Z(n65) );
  XOR U99 ( .A(B[971]), .B(A[971]), .Z(n66) );
  XOR U100 ( .A(A[970]), .B(n67), .Z(O[970]) );
  AND U101 ( .A(S), .B(n68), .Z(n67) );
  XOR U102 ( .A(B[970]), .B(A[970]), .Z(n68) );
  XOR U103 ( .A(A[96]), .B(n69), .Z(O[96]) );
  AND U104 ( .A(S), .B(n70), .Z(n69) );
  XOR U105 ( .A(B[96]), .B(A[96]), .Z(n70) );
  XOR U106 ( .A(A[969]), .B(n71), .Z(O[969]) );
  AND U107 ( .A(S), .B(n72), .Z(n71) );
  XOR U108 ( .A(B[969]), .B(A[969]), .Z(n72) );
  XOR U109 ( .A(A[968]), .B(n73), .Z(O[968]) );
  AND U110 ( .A(S), .B(n74), .Z(n73) );
  XOR U111 ( .A(B[968]), .B(A[968]), .Z(n74) );
  XOR U112 ( .A(A[967]), .B(n75), .Z(O[967]) );
  AND U113 ( .A(S), .B(n76), .Z(n75) );
  XOR U114 ( .A(B[967]), .B(A[967]), .Z(n76) );
  XOR U115 ( .A(A[966]), .B(n77), .Z(O[966]) );
  AND U116 ( .A(S), .B(n78), .Z(n77) );
  XOR U117 ( .A(B[966]), .B(A[966]), .Z(n78) );
  XOR U118 ( .A(A[965]), .B(n79), .Z(O[965]) );
  AND U119 ( .A(S), .B(n80), .Z(n79) );
  XOR U120 ( .A(B[965]), .B(A[965]), .Z(n80) );
  XOR U121 ( .A(A[964]), .B(n81), .Z(O[964]) );
  AND U122 ( .A(S), .B(n82), .Z(n81) );
  XOR U123 ( .A(B[964]), .B(A[964]), .Z(n82) );
  XOR U124 ( .A(A[963]), .B(n83), .Z(O[963]) );
  AND U125 ( .A(S), .B(n84), .Z(n83) );
  XOR U126 ( .A(B[963]), .B(A[963]), .Z(n84) );
  XOR U127 ( .A(A[962]), .B(n85), .Z(O[962]) );
  AND U128 ( .A(S), .B(n86), .Z(n85) );
  XOR U129 ( .A(B[962]), .B(A[962]), .Z(n86) );
  XOR U130 ( .A(A[961]), .B(n87), .Z(O[961]) );
  AND U131 ( .A(S), .B(n88), .Z(n87) );
  XOR U132 ( .A(B[961]), .B(A[961]), .Z(n88) );
  XOR U133 ( .A(A[960]), .B(n89), .Z(O[960]) );
  AND U134 ( .A(S), .B(n90), .Z(n89) );
  XOR U135 ( .A(B[960]), .B(A[960]), .Z(n90) );
  XOR U136 ( .A(A[95]), .B(n91), .Z(O[95]) );
  AND U137 ( .A(S), .B(n92), .Z(n91) );
  XOR U138 ( .A(B[95]), .B(A[95]), .Z(n92) );
  XOR U139 ( .A(A[959]), .B(n93), .Z(O[959]) );
  AND U140 ( .A(S), .B(n94), .Z(n93) );
  XOR U141 ( .A(B[959]), .B(A[959]), .Z(n94) );
  XOR U142 ( .A(A[958]), .B(n95), .Z(O[958]) );
  AND U143 ( .A(S), .B(n96), .Z(n95) );
  XOR U144 ( .A(B[958]), .B(A[958]), .Z(n96) );
  XOR U145 ( .A(A[957]), .B(n97), .Z(O[957]) );
  AND U146 ( .A(S), .B(n98), .Z(n97) );
  XOR U147 ( .A(B[957]), .B(A[957]), .Z(n98) );
  XOR U148 ( .A(A[956]), .B(n99), .Z(O[956]) );
  AND U149 ( .A(S), .B(n100), .Z(n99) );
  XOR U150 ( .A(B[956]), .B(A[956]), .Z(n100) );
  XOR U151 ( .A(A[955]), .B(n101), .Z(O[955]) );
  AND U152 ( .A(S), .B(n102), .Z(n101) );
  XOR U153 ( .A(B[955]), .B(A[955]), .Z(n102) );
  XOR U154 ( .A(A[954]), .B(n103), .Z(O[954]) );
  AND U155 ( .A(S), .B(n104), .Z(n103) );
  XOR U156 ( .A(B[954]), .B(A[954]), .Z(n104) );
  XOR U157 ( .A(A[953]), .B(n105), .Z(O[953]) );
  AND U158 ( .A(S), .B(n106), .Z(n105) );
  XOR U159 ( .A(B[953]), .B(A[953]), .Z(n106) );
  XOR U160 ( .A(A[952]), .B(n107), .Z(O[952]) );
  AND U161 ( .A(S), .B(n108), .Z(n107) );
  XOR U162 ( .A(B[952]), .B(A[952]), .Z(n108) );
  XOR U163 ( .A(A[951]), .B(n109), .Z(O[951]) );
  AND U164 ( .A(S), .B(n110), .Z(n109) );
  XOR U165 ( .A(B[951]), .B(A[951]), .Z(n110) );
  XOR U166 ( .A(A[950]), .B(n111), .Z(O[950]) );
  AND U167 ( .A(S), .B(n112), .Z(n111) );
  XOR U168 ( .A(B[950]), .B(A[950]), .Z(n112) );
  XOR U169 ( .A(A[94]), .B(n113), .Z(O[94]) );
  AND U170 ( .A(S), .B(n114), .Z(n113) );
  XOR U171 ( .A(B[94]), .B(A[94]), .Z(n114) );
  XOR U172 ( .A(A[949]), .B(n115), .Z(O[949]) );
  AND U173 ( .A(S), .B(n116), .Z(n115) );
  XOR U174 ( .A(B[949]), .B(A[949]), .Z(n116) );
  XOR U175 ( .A(A[948]), .B(n117), .Z(O[948]) );
  AND U176 ( .A(S), .B(n118), .Z(n117) );
  XOR U177 ( .A(B[948]), .B(A[948]), .Z(n118) );
  XOR U178 ( .A(A[947]), .B(n119), .Z(O[947]) );
  AND U179 ( .A(S), .B(n120), .Z(n119) );
  XOR U180 ( .A(B[947]), .B(A[947]), .Z(n120) );
  XOR U181 ( .A(A[946]), .B(n121), .Z(O[946]) );
  AND U182 ( .A(S), .B(n122), .Z(n121) );
  XOR U183 ( .A(B[946]), .B(A[946]), .Z(n122) );
  XOR U184 ( .A(A[945]), .B(n123), .Z(O[945]) );
  AND U185 ( .A(S), .B(n124), .Z(n123) );
  XOR U186 ( .A(B[945]), .B(A[945]), .Z(n124) );
  XOR U187 ( .A(A[944]), .B(n125), .Z(O[944]) );
  AND U188 ( .A(S), .B(n126), .Z(n125) );
  XOR U189 ( .A(B[944]), .B(A[944]), .Z(n126) );
  XOR U190 ( .A(A[943]), .B(n127), .Z(O[943]) );
  AND U191 ( .A(S), .B(n128), .Z(n127) );
  XOR U192 ( .A(B[943]), .B(A[943]), .Z(n128) );
  XOR U193 ( .A(A[942]), .B(n129), .Z(O[942]) );
  AND U194 ( .A(S), .B(n130), .Z(n129) );
  XOR U195 ( .A(B[942]), .B(A[942]), .Z(n130) );
  XOR U196 ( .A(A[941]), .B(n131), .Z(O[941]) );
  AND U197 ( .A(S), .B(n132), .Z(n131) );
  XOR U198 ( .A(B[941]), .B(A[941]), .Z(n132) );
  XOR U199 ( .A(A[940]), .B(n133), .Z(O[940]) );
  AND U200 ( .A(S), .B(n134), .Z(n133) );
  XOR U201 ( .A(B[940]), .B(A[940]), .Z(n134) );
  XOR U202 ( .A(A[93]), .B(n135), .Z(O[93]) );
  AND U203 ( .A(S), .B(n136), .Z(n135) );
  XOR U204 ( .A(B[93]), .B(A[93]), .Z(n136) );
  XOR U205 ( .A(A[939]), .B(n137), .Z(O[939]) );
  AND U206 ( .A(S), .B(n138), .Z(n137) );
  XOR U207 ( .A(B[939]), .B(A[939]), .Z(n138) );
  XOR U208 ( .A(A[938]), .B(n139), .Z(O[938]) );
  AND U209 ( .A(S), .B(n140), .Z(n139) );
  XOR U210 ( .A(B[938]), .B(A[938]), .Z(n140) );
  XOR U211 ( .A(A[937]), .B(n141), .Z(O[937]) );
  AND U212 ( .A(S), .B(n142), .Z(n141) );
  XOR U213 ( .A(B[937]), .B(A[937]), .Z(n142) );
  XOR U214 ( .A(A[936]), .B(n143), .Z(O[936]) );
  AND U215 ( .A(S), .B(n144), .Z(n143) );
  XOR U216 ( .A(B[936]), .B(A[936]), .Z(n144) );
  XOR U217 ( .A(A[935]), .B(n145), .Z(O[935]) );
  AND U218 ( .A(S), .B(n146), .Z(n145) );
  XOR U219 ( .A(B[935]), .B(A[935]), .Z(n146) );
  XOR U220 ( .A(A[934]), .B(n147), .Z(O[934]) );
  AND U221 ( .A(S), .B(n148), .Z(n147) );
  XOR U222 ( .A(B[934]), .B(A[934]), .Z(n148) );
  XOR U223 ( .A(A[933]), .B(n149), .Z(O[933]) );
  AND U224 ( .A(S), .B(n150), .Z(n149) );
  XOR U225 ( .A(B[933]), .B(A[933]), .Z(n150) );
  XOR U226 ( .A(A[932]), .B(n151), .Z(O[932]) );
  AND U227 ( .A(S), .B(n152), .Z(n151) );
  XOR U228 ( .A(B[932]), .B(A[932]), .Z(n152) );
  XOR U229 ( .A(A[931]), .B(n153), .Z(O[931]) );
  AND U230 ( .A(S), .B(n154), .Z(n153) );
  XOR U231 ( .A(B[931]), .B(A[931]), .Z(n154) );
  XOR U232 ( .A(A[930]), .B(n155), .Z(O[930]) );
  AND U233 ( .A(S), .B(n156), .Z(n155) );
  XOR U234 ( .A(B[930]), .B(A[930]), .Z(n156) );
  XOR U235 ( .A(A[92]), .B(n157), .Z(O[92]) );
  AND U236 ( .A(S), .B(n158), .Z(n157) );
  XOR U237 ( .A(B[92]), .B(A[92]), .Z(n158) );
  XOR U238 ( .A(A[929]), .B(n159), .Z(O[929]) );
  AND U239 ( .A(S), .B(n160), .Z(n159) );
  XOR U240 ( .A(B[929]), .B(A[929]), .Z(n160) );
  XOR U241 ( .A(A[928]), .B(n161), .Z(O[928]) );
  AND U242 ( .A(S), .B(n162), .Z(n161) );
  XOR U243 ( .A(B[928]), .B(A[928]), .Z(n162) );
  XOR U244 ( .A(A[927]), .B(n163), .Z(O[927]) );
  AND U245 ( .A(S), .B(n164), .Z(n163) );
  XOR U246 ( .A(B[927]), .B(A[927]), .Z(n164) );
  XOR U247 ( .A(A[926]), .B(n165), .Z(O[926]) );
  AND U248 ( .A(S), .B(n166), .Z(n165) );
  XOR U249 ( .A(B[926]), .B(A[926]), .Z(n166) );
  XOR U250 ( .A(A[925]), .B(n167), .Z(O[925]) );
  AND U251 ( .A(S), .B(n168), .Z(n167) );
  XOR U252 ( .A(B[925]), .B(A[925]), .Z(n168) );
  XOR U253 ( .A(A[924]), .B(n169), .Z(O[924]) );
  AND U254 ( .A(S), .B(n170), .Z(n169) );
  XOR U255 ( .A(B[924]), .B(A[924]), .Z(n170) );
  XOR U256 ( .A(A[923]), .B(n171), .Z(O[923]) );
  AND U257 ( .A(S), .B(n172), .Z(n171) );
  XOR U258 ( .A(B[923]), .B(A[923]), .Z(n172) );
  XOR U259 ( .A(A[922]), .B(n173), .Z(O[922]) );
  AND U260 ( .A(S), .B(n174), .Z(n173) );
  XOR U261 ( .A(B[922]), .B(A[922]), .Z(n174) );
  XOR U262 ( .A(A[921]), .B(n175), .Z(O[921]) );
  AND U263 ( .A(S), .B(n176), .Z(n175) );
  XOR U264 ( .A(B[921]), .B(A[921]), .Z(n176) );
  XOR U265 ( .A(A[920]), .B(n177), .Z(O[920]) );
  AND U266 ( .A(S), .B(n178), .Z(n177) );
  XOR U267 ( .A(B[920]), .B(A[920]), .Z(n178) );
  XOR U268 ( .A(A[91]), .B(n179), .Z(O[91]) );
  AND U269 ( .A(S), .B(n180), .Z(n179) );
  XOR U270 ( .A(B[91]), .B(A[91]), .Z(n180) );
  XOR U271 ( .A(A[919]), .B(n181), .Z(O[919]) );
  AND U272 ( .A(S), .B(n182), .Z(n181) );
  XOR U273 ( .A(B[919]), .B(A[919]), .Z(n182) );
  XOR U274 ( .A(A[918]), .B(n183), .Z(O[918]) );
  AND U275 ( .A(S), .B(n184), .Z(n183) );
  XOR U276 ( .A(B[918]), .B(A[918]), .Z(n184) );
  XOR U277 ( .A(A[917]), .B(n185), .Z(O[917]) );
  AND U278 ( .A(S), .B(n186), .Z(n185) );
  XOR U279 ( .A(B[917]), .B(A[917]), .Z(n186) );
  XOR U280 ( .A(A[916]), .B(n187), .Z(O[916]) );
  AND U281 ( .A(S), .B(n188), .Z(n187) );
  XOR U282 ( .A(B[916]), .B(A[916]), .Z(n188) );
  XOR U283 ( .A(A[915]), .B(n189), .Z(O[915]) );
  AND U284 ( .A(S), .B(n190), .Z(n189) );
  XOR U285 ( .A(B[915]), .B(A[915]), .Z(n190) );
  XOR U286 ( .A(A[914]), .B(n191), .Z(O[914]) );
  AND U287 ( .A(S), .B(n192), .Z(n191) );
  XOR U288 ( .A(B[914]), .B(A[914]), .Z(n192) );
  XOR U289 ( .A(A[913]), .B(n193), .Z(O[913]) );
  AND U290 ( .A(S), .B(n194), .Z(n193) );
  XOR U291 ( .A(B[913]), .B(A[913]), .Z(n194) );
  XOR U292 ( .A(A[912]), .B(n195), .Z(O[912]) );
  AND U293 ( .A(S), .B(n196), .Z(n195) );
  XOR U294 ( .A(B[912]), .B(A[912]), .Z(n196) );
  XOR U295 ( .A(A[911]), .B(n197), .Z(O[911]) );
  AND U296 ( .A(S), .B(n198), .Z(n197) );
  XOR U297 ( .A(B[911]), .B(A[911]), .Z(n198) );
  XOR U298 ( .A(A[910]), .B(n199), .Z(O[910]) );
  AND U299 ( .A(S), .B(n200), .Z(n199) );
  XOR U300 ( .A(B[910]), .B(A[910]), .Z(n200) );
  XOR U301 ( .A(A[90]), .B(n201), .Z(O[90]) );
  AND U302 ( .A(S), .B(n202), .Z(n201) );
  XOR U303 ( .A(B[90]), .B(A[90]), .Z(n202) );
  XOR U304 ( .A(A[909]), .B(n203), .Z(O[909]) );
  AND U305 ( .A(S), .B(n204), .Z(n203) );
  XOR U306 ( .A(B[909]), .B(A[909]), .Z(n204) );
  XOR U307 ( .A(A[908]), .B(n205), .Z(O[908]) );
  AND U308 ( .A(S), .B(n206), .Z(n205) );
  XOR U309 ( .A(B[908]), .B(A[908]), .Z(n206) );
  XOR U310 ( .A(A[907]), .B(n207), .Z(O[907]) );
  AND U311 ( .A(S), .B(n208), .Z(n207) );
  XOR U312 ( .A(B[907]), .B(A[907]), .Z(n208) );
  XOR U313 ( .A(A[906]), .B(n209), .Z(O[906]) );
  AND U314 ( .A(S), .B(n210), .Z(n209) );
  XOR U315 ( .A(B[906]), .B(A[906]), .Z(n210) );
  XOR U316 ( .A(A[905]), .B(n211), .Z(O[905]) );
  AND U317 ( .A(S), .B(n212), .Z(n211) );
  XOR U318 ( .A(B[905]), .B(A[905]), .Z(n212) );
  XOR U319 ( .A(A[904]), .B(n213), .Z(O[904]) );
  AND U320 ( .A(S), .B(n214), .Z(n213) );
  XOR U321 ( .A(B[904]), .B(A[904]), .Z(n214) );
  XOR U322 ( .A(A[903]), .B(n215), .Z(O[903]) );
  AND U323 ( .A(S), .B(n216), .Z(n215) );
  XOR U324 ( .A(B[903]), .B(A[903]), .Z(n216) );
  XOR U325 ( .A(A[902]), .B(n217), .Z(O[902]) );
  AND U326 ( .A(S), .B(n218), .Z(n217) );
  XOR U327 ( .A(B[902]), .B(A[902]), .Z(n218) );
  XOR U328 ( .A(A[901]), .B(n219), .Z(O[901]) );
  AND U329 ( .A(S), .B(n220), .Z(n219) );
  XOR U330 ( .A(B[901]), .B(A[901]), .Z(n220) );
  XOR U331 ( .A(A[900]), .B(n221), .Z(O[900]) );
  AND U332 ( .A(S), .B(n222), .Z(n221) );
  XOR U333 ( .A(B[900]), .B(A[900]), .Z(n222) );
  XOR U334 ( .A(A[8]), .B(n223), .Z(O[8]) );
  AND U335 ( .A(S), .B(n224), .Z(n223) );
  XOR U336 ( .A(B[8]), .B(A[8]), .Z(n224) );
  XOR U337 ( .A(A[89]), .B(n225), .Z(O[89]) );
  AND U338 ( .A(S), .B(n226), .Z(n225) );
  XOR U339 ( .A(B[89]), .B(A[89]), .Z(n226) );
  XOR U340 ( .A(A[899]), .B(n227), .Z(O[899]) );
  AND U341 ( .A(S), .B(n228), .Z(n227) );
  XOR U342 ( .A(B[899]), .B(A[899]), .Z(n228) );
  XOR U343 ( .A(A[898]), .B(n229), .Z(O[898]) );
  AND U344 ( .A(S), .B(n230), .Z(n229) );
  XOR U345 ( .A(B[898]), .B(A[898]), .Z(n230) );
  XOR U346 ( .A(A[897]), .B(n231), .Z(O[897]) );
  AND U347 ( .A(S), .B(n232), .Z(n231) );
  XOR U348 ( .A(B[897]), .B(A[897]), .Z(n232) );
  XOR U349 ( .A(A[896]), .B(n233), .Z(O[896]) );
  AND U350 ( .A(S), .B(n234), .Z(n233) );
  XOR U351 ( .A(B[896]), .B(A[896]), .Z(n234) );
  XOR U352 ( .A(A[895]), .B(n235), .Z(O[895]) );
  AND U353 ( .A(S), .B(n236), .Z(n235) );
  XOR U354 ( .A(B[895]), .B(A[895]), .Z(n236) );
  XOR U355 ( .A(A[894]), .B(n237), .Z(O[894]) );
  AND U356 ( .A(S), .B(n238), .Z(n237) );
  XOR U357 ( .A(B[894]), .B(A[894]), .Z(n238) );
  XOR U358 ( .A(A[893]), .B(n239), .Z(O[893]) );
  AND U359 ( .A(S), .B(n240), .Z(n239) );
  XOR U360 ( .A(B[893]), .B(A[893]), .Z(n240) );
  XOR U361 ( .A(A[892]), .B(n241), .Z(O[892]) );
  AND U362 ( .A(S), .B(n242), .Z(n241) );
  XOR U363 ( .A(B[892]), .B(A[892]), .Z(n242) );
  XOR U364 ( .A(A[891]), .B(n243), .Z(O[891]) );
  AND U365 ( .A(S), .B(n244), .Z(n243) );
  XOR U366 ( .A(B[891]), .B(A[891]), .Z(n244) );
  XOR U367 ( .A(A[890]), .B(n245), .Z(O[890]) );
  AND U368 ( .A(S), .B(n246), .Z(n245) );
  XOR U369 ( .A(B[890]), .B(A[890]), .Z(n246) );
  XOR U370 ( .A(A[88]), .B(n247), .Z(O[88]) );
  AND U371 ( .A(S), .B(n248), .Z(n247) );
  XOR U372 ( .A(B[88]), .B(A[88]), .Z(n248) );
  XOR U373 ( .A(A[889]), .B(n249), .Z(O[889]) );
  AND U374 ( .A(S), .B(n250), .Z(n249) );
  XOR U375 ( .A(B[889]), .B(A[889]), .Z(n250) );
  XOR U376 ( .A(A[888]), .B(n251), .Z(O[888]) );
  AND U377 ( .A(S), .B(n252), .Z(n251) );
  XOR U378 ( .A(B[888]), .B(A[888]), .Z(n252) );
  XOR U379 ( .A(A[887]), .B(n253), .Z(O[887]) );
  AND U380 ( .A(S), .B(n254), .Z(n253) );
  XOR U381 ( .A(B[887]), .B(A[887]), .Z(n254) );
  XOR U382 ( .A(A[886]), .B(n255), .Z(O[886]) );
  AND U383 ( .A(S), .B(n256), .Z(n255) );
  XOR U384 ( .A(B[886]), .B(A[886]), .Z(n256) );
  XOR U385 ( .A(A[885]), .B(n257), .Z(O[885]) );
  AND U386 ( .A(S), .B(n258), .Z(n257) );
  XOR U387 ( .A(B[885]), .B(A[885]), .Z(n258) );
  XOR U388 ( .A(A[884]), .B(n259), .Z(O[884]) );
  AND U389 ( .A(S), .B(n260), .Z(n259) );
  XOR U390 ( .A(B[884]), .B(A[884]), .Z(n260) );
  XOR U391 ( .A(A[883]), .B(n261), .Z(O[883]) );
  AND U392 ( .A(S), .B(n262), .Z(n261) );
  XOR U393 ( .A(B[883]), .B(A[883]), .Z(n262) );
  XOR U394 ( .A(A[882]), .B(n263), .Z(O[882]) );
  AND U395 ( .A(S), .B(n264), .Z(n263) );
  XOR U396 ( .A(B[882]), .B(A[882]), .Z(n264) );
  XOR U397 ( .A(A[881]), .B(n265), .Z(O[881]) );
  AND U398 ( .A(S), .B(n266), .Z(n265) );
  XOR U399 ( .A(B[881]), .B(A[881]), .Z(n266) );
  XOR U400 ( .A(A[880]), .B(n267), .Z(O[880]) );
  AND U401 ( .A(S), .B(n268), .Z(n267) );
  XOR U402 ( .A(B[880]), .B(A[880]), .Z(n268) );
  XOR U403 ( .A(A[87]), .B(n269), .Z(O[87]) );
  AND U404 ( .A(S), .B(n270), .Z(n269) );
  XOR U405 ( .A(B[87]), .B(A[87]), .Z(n270) );
  XOR U406 ( .A(A[879]), .B(n271), .Z(O[879]) );
  AND U407 ( .A(S), .B(n272), .Z(n271) );
  XOR U408 ( .A(B[879]), .B(A[879]), .Z(n272) );
  XOR U409 ( .A(A[878]), .B(n273), .Z(O[878]) );
  AND U410 ( .A(S), .B(n274), .Z(n273) );
  XOR U411 ( .A(B[878]), .B(A[878]), .Z(n274) );
  XOR U412 ( .A(A[877]), .B(n275), .Z(O[877]) );
  AND U413 ( .A(S), .B(n276), .Z(n275) );
  XOR U414 ( .A(B[877]), .B(A[877]), .Z(n276) );
  XOR U415 ( .A(A[876]), .B(n277), .Z(O[876]) );
  AND U416 ( .A(S), .B(n278), .Z(n277) );
  XOR U417 ( .A(B[876]), .B(A[876]), .Z(n278) );
  XOR U418 ( .A(A[875]), .B(n279), .Z(O[875]) );
  AND U419 ( .A(S), .B(n280), .Z(n279) );
  XOR U420 ( .A(B[875]), .B(A[875]), .Z(n280) );
  XOR U421 ( .A(A[874]), .B(n281), .Z(O[874]) );
  AND U422 ( .A(S), .B(n282), .Z(n281) );
  XOR U423 ( .A(B[874]), .B(A[874]), .Z(n282) );
  XOR U424 ( .A(A[873]), .B(n283), .Z(O[873]) );
  AND U425 ( .A(S), .B(n284), .Z(n283) );
  XOR U426 ( .A(B[873]), .B(A[873]), .Z(n284) );
  XOR U427 ( .A(A[872]), .B(n285), .Z(O[872]) );
  AND U428 ( .A(S), .B(n286), .Z(n285) );
  XOR U429 ( .A(B[872]), .B(A[872]), .Z(n286) );
  XOR U430 ( .A(A[871]), .B(n287), .Z(O[871]) );
  AND U431 ( .A(S), .B(n288), .Z(n287) );
  XOR U432 ( .A(B[871]), .B(A[871]), .Z(n288) );
  XOR U433 ( .A(A[870]), .B(n289), .Z(O[870]) );
  AND U434 ( .A(S), .B(n290), .Z(n289) );
  XOR U435 ( .A(B[870]), .B(A[870]), .Z(n290) );
  XOR U436 ( .A(A[86]), .B(n291), .Z(O[86]) );
  AND U437 ( .A(S), .B(n292), .Z(n291) );
  XOR U438 ( .A(B[86]), .B(A[86]), .Z(n292) );
  XOR U439 ( .A(A[869]), .B(n293), .Z(O[869]) );
  AND U440 ( .A(S), .B(n294), .Z(n293) );
  XOR U441 ( .A(B[869]), .B(A[869]), .Z(n294) );
  XOR U442 ( .A(A[868]), .B(n295), .Z(O[868]) );
  AND U443 ( .A(S), .B(n296), .Z(n295) );
  XOR U444 ( .A(B[868]), .B(A[868]), .Z(n296) );
  XOR U445 ( .A(A[867]), .B(n297), .Z(O[867]) );
  AND U446 ( .A(S), .B(n298), .Z(n297) );
  XOR U447 ( .A(B[867]), .B(A[867]), .Z(n298) );
  XOR U448 ( .A(A[866]), .B(n299), .Z(O[866]) );
  AND U449 ( .A(S), .B(n300), .Z(n299) );
  XOR U450 ( .A(B[866]), .B(A[866]), .Z(n300) );
  XOR U451 ( .A(A[865]), .B(n301), .Z(O[865]) );
  AND U452 ( .A(S), .B(n302), .Z(n301) );
  XOR U453 ( .A(B[865]), .B(A[865]), .Z(n302) );
  XOR U454 ( .A(A[864]), .B(n303), .Z(O[864]) );
  AND U455 ( .A(S), .B(n304), .Z(n303) );
  XOR U456 ( .A(B[864]), .B(A[864]), .Z(n304) );
  XOR U457 ( .A(A[863]), .B(n305), .Z(O[863]) );
  AND U458 ( .A(S), .B(n306), .Z(n305) );
  XOR U459 ( .A(B[863]), .B(A[863]), .Z(n306) );
  XOR U460 ( .A(A[862]), .B(n307), .Z(O[862]) );
  AND U461 ( .A(S), .B(n308), .Z(n307) );
  XOR U462 ( .A(B[862]), .B(A[862]), .Z(n308) );
  XOR U463 ( .A(A[861]), .B(n309), .Z(O[861]) );
  AND U464 ( .A(S), .B(n310), .Z(n309) );
  XOR U465 ( .A(B[861]), .B(A[861]), .Z(n310) );
  XOR U466 ( .A(A[860]), .B(n311), .Z(O[860]) );
  AND U467 ( .A(S), .B(n312), .Z(n311) );
  XOR U468 ( .A(B[860]), .B(A[860]), .Z(n312) );
  XOR U469 ( .A(A[85]), .B(n313), .Z(O[85]) );
  AND U470 ( .A(S), .B(n314), .Z(n313) );
  XOR U471 ( .A(B[85]), .B(A[85]), .Z(n314) );
  XOR U472 ( .A(A[859]), .B(n315), .Z(O[859]) );
  AND U473 ( .A(S), .B(n316), .Z(n315) );
  XOR U474 ( .A(B[859]), .B(A[859]), .Z(n316) );
  XOR U475 ( .A(A[858]), .B(n317), .Z(O[858]) );
  AND U476 ( .A(S), .B(n318), .Z(n317) );
  XOR U477 ( .A(B[858]), .B(A[858]), .Z(n318) );
  XOR U478 ( .A(A[857]), .B(n319), .Z(O[857]) );
  AND U479 ( .A(S), .B(n320), .Z(n319) );
  XOR U480 ( .A(B[857]), .B(A[857]), .Z(n320) );
  XOR U481 ( .A(A[856]), .B(n321), .Z(O[856]) );
  AND U482 ( .A(S), .B(n322), .Z(n321) );
  XOR U483 ( .A(B[856]), .B(A[856]), .Z(n322) );
  XOR U484 ( .A(A[855]), .B(n323), .Z(O[855]) );
  AND U485 ( .A(S), .B(n324), .Z(n323) );
  XOR U486 ( .A(B[855]), .B(A[855]), .Z(n324) );
  XOR U487 ( .A(A[854]), .B(n325), .Z(O[854]) );
  AND U488 ( .A(S), .B(n326), .Z(n325) );
  XOR U489 ( .A(B[854]), .B(A[854]), .Z(n326) );
  XOR U490 ( .A(A[853]), .B(n327), .Z(O[853]) );
  AND U491 ( .A(S), .B(n328), .Z(n327) );
  XOR U492 ( .A(B[853]), .B(A[853]), .Z(n328) );
  XOR U493 ( .A(A[852]), .B(n329), .Z(O[852]) );
  AND U494 ( .A(S), .B(n330), .Z(n329) );
  XOR U495 ( .A(B[852]), .B(A[852]), .Z(n330) );
  XOR U496 ( .A(A[851]), .B(n331), .Z(O[851]) );
  AND U497 ( .A(S), .B(n332), .Z(n331) );
  XOR U498 ( .A(B[851]), .B(A[851]), .Z(n332) );
  XOR U499 ( .A(A[850]), .B(n333), .Z(O[850]) );
  AND U500 ( .A(S), .B(n334), .Z(n333) );
  XOR U501 ( .A(B[850]), .B(A[850]), .Z(n334) );
  XOR U502 ( .A(A[84]), .B(n335), .Z(O[84]) );
  AND U503 ( .A(S), .B(n336), .Z(n335) );
  XOR U504 ( .A(B[84]), .B(A[84]), .Z(n336) );
  XOR U505 ( .A(A[849]), .B(n337), .Z(O[849]) );
  AND U506 ( .A(S), .B(n338), .Z(n337) );
  XOR U507 ( .A(B[849]), .B(A[849]), .Z(n338) );
  XOR U508 ( .A(A[848]), .B(n339), .Z(O[848]) );
  AND U509 ( .A(S), .B(n340), .Z(n339) );
  XOR U510 ( .A(B[848]), .B(A[848]), .Z(n340) );
  XOR U511 ( .A(A[847]), .B(n341), .Z(O[847]) );
  AND U512 ( .A(S), .B(n342), .Z(n341) );
  XOR U513 ( .A(B[847]), .B(A[847]), .Z(n342) );
  XOR U514 ( .A(A[846]), .B(n343), .Z(O[846]) );
  AND U515 ( .A(S), .B(n344), .Z(n343) );
  XOR U516 ( .A(B[846]), .B(A[846]), .Z(n344) );
  XOR U517 ( .A(A[845]), .B(n345), .Z(O[845]) );
  AND U518 ( .A(S), .B(n346), .Z(n345) );
  XOR U519 ( .A(B[845]), .B(A[845]), .Z(n346) );
  XOR U520 ( .A(A[844]), .B(n347), .Z(O[844]) );
  AND U521 ( .A(S), .B(n348), .Z(n347) );
  XOR U522 ( .A(B[844]), .B(A[844]), .Z(n348) );
  XOR U523 ( .A(A[843]), .B(n349), .Z(O[843]) );
  AND U524 ( .A(S), .B(n350), .Z(n349) );
  XOR U525 ( .A(B[843]), .B(A[843]), .Z(n350) );
  XOR U526 ( .A(A[842]), .B(n351), .Z(O[842]) );
  AND U527 ( .A(S), .B(n352), .Z(n351) );
  XOR U528 ( .A(B[842]), .B(A[842]), .Z(n352) );
  XOR U529 ( .A(A[841]), .B(n353), .Z(O[841]) );
  AND U530 ( .A(S), .B(n354), .Z(n353) );
  XOR U531 ( .A(B[841]), .B(A[841]), .Z(n354) );
  XOR U532 ( .A(A[840]), .B(n355), .Z(O[840]) );
  AND U533 ( .A(S), .B(n356), .Z(n355) );
  XOR U534 ( .A(B[840]), .B(A[840]), .Z(n356) );
  XOR U535 ( .A(A[83]), .B(n357), .Z(O[83]) );
  AND U536 ( .A(S), .B(n358), .Z(n357) );
  XOR U537 ( .A(B[83]), .B(A[83]), .Z(n358) );
  XOR U538 ( .A(A[839]), .B(n359), .Z(O[839]) );
  AND U539 ( .A(S), .B(n360), .Z(n359) );
  XOR U540 ( .A(B[839]), .B(A[839]), .Z(n360) );
  XOR U541 ( .A(A[838]), .B(n361), .Z(O[838]) );
  AND U542 ( .A(S), .B(n362), .Z(n361) );
  XOR U543 ( .A(B[838]), .B(A[838]), .Z(n362) );
  XOR U544 ( .A(A[837]), .B(n363), .Z(O[837]) );
  AND U545 ( .A(S), .B(n364), .Z(n363) );
  XOR U546 ( .A(B[837]), .B(A[837]), .Z(n364) );
  XOR U547 ( .A(A[836]), .B(n365), .Z(O[836]) );
  AND U548 ( .A(S), .B(n366), .Z(n365) );
  XOR U549 ( .A(B[836]), .B(A[836]), .Z(n366) );
  XOR U550 ( .A(A[835]), .B(n367), .Z(O[835]) );
  AND U551 ( .A(S), .B(n368), .Z(n367) );
  XOR U552 ( .A(B[835]), .B(A[835]), .Z(n368) );
  XOR U553 ( .A(A[834]), .B(n369), .Z(O[834]) );
  AND U554 ( .A(S), .B(n370), .Z(n369) );
  XOR U555 ( .A(B[834]), .B(A[834]), .Z(n370) );
  XOR U556 ( .A(A[833]), .B(n371), .Z(O[833]) );
  AND U557 ( .A(S), .B(n372), .Z(n371) );
  XOR U558 ( .A(B[833]), .B(A[833]), .Z(n372) );
  XOR U559 ( .A(A[832]), .B(n373), .Z(O[832]) );
  AND U560 ( .A(S), .B(n374), .Z(n373) );
  XOR U561 ( .A(B[832]), .B(A[832]), .Z(n374) );
  XOR U562 ( .A(A[831]), .B(n375), .Z(O[831]) );
  AND U563 ( .A(S), .B(n376), .Z(n375) );
  XOR U564 ( .A(B[831]), .B(A[831]), .Z(n376) );
  XOR U565 ( .A(A[830]), .B(n377), .Z(O[830]) );
  AND U566 ( .A(S), .B(n378), .Z(n377) );
  XOR U567 ( .A(B[830]), .B(A[830]), .Z(n378) );
  XOR U568 ( .A(A[82]), .B(n379), .Z(O[82]) );
  AND U569 ( .A(S), .B(n380), .Z(n379) );
  XOR U570 ( .A(B[82]), .B(A[82]), .Z(n380) );
  XOR U571 ( .A(A[829]), .B(n381), .Z(O[829]) );
  AND U572 ( .A(S), .B(n382), .Z(n381) );
  XOR U573 ( .A(B[829]), .B(A[829]), .Z(n382) );
  XOR U574 ( .A(A[828]), .B(n383), .Z(O[828]) );
  AND U575 ( .A(S), .B(n384), .Z(n383) );
  XOR U576 ( .A(B[828]), .B(A[828]), .Z(n384) );
  XOR U577 ( .A(A[827]), .B(n385), .Z(O[827]) );
  AND U578 ( .A(S), .B(n386), .Z(n385) );
  XOR U579 ( .A(B[827]), .B(A[827]), .Z(n386) );
  XOR U580 ( .A(A[826]), .B(n387), .Z(O[826]) );
  AND U581 ( .A(S), .B(n388), .Z(n387) );
  XOR U582 ( .A(B[826]), .B(A[826]), .Z(n388) );
  XOR U583 ( .A(A[825]), .B(n389), .Z(O[825]) );
  AND U584 ( .A(S), .B(n390), .Z(n389) );
  XOR U585 ( .A(B[825]), .B(A[825]), .Z(n390) );
  XOR U586 ( .A(A[824]), .B(n391), .Z(O[824]) );
  AND U587 ( .A(S), .B(n392), .Z(n391) );
  XOR U588 ( .A(B[824]), .B(A[824]), .Z(n392) );
  XOR U589 ( .A(A[823]), .B(n393), .Z(O[823]) );
  AND U590 ( .A(S), .B(n394), .Z(n393) );
  XOR U591 ( .A(B[823]), .B(A[823]), .Z(n394) );
  XOR U592 ( .A(A[822]), .B(n395), .Z(O[822]) );
  AND U593 ( .A(S), .B(n396), .Z(n395) );
  XOR U594 ( .A(B[822]), .B(A[822]), .Z(n396) );
  XOR U595 ( .A(A[821]), .B(n397), .Z(O[821]) );
  AND U596 ( .A(S), .B(n398), .Z(n397) );
  XOR U597 ( .A(B[821]), .B(A[821]), .Z(n398) );
  XOR U598 ( .A(A[820]), .B(n399), .Z(O[820]) );
  AND U599 ( .A(S), .B(n400), .Z(n399) );
  XOR U600 ( .A(B[820]), .B(A[820]), .Z(n400) );
  XOR U601 ( .A(A[81]), .B(n401), .Z(O[81]) );
  AND U602 ( .A(S), .B(n402), .Z(n401) );
  XOR U603 ( .A(B[81]), .B(A[81]), .Z(n402) );
  XOR U604 ( .A(A[819]), .B(n403), .Z(O[819]) );
  AND U605 ( .A(S), .B(n404), .Z(n403) );
  XOR U606 ( .A(B[819]), .B(A[819]), .Z(n404) );
  XOR U607 ( .A(A[818]), .B(n405), .Z(O[818]) );
  AND U608 ( .A(S), .B(n406), .Z(n405) );
  XOR U609 ( .A(B[818]), .B(A[818]), .Z(n406) );
  XOR U610 ( .A(A[817]), .B(n407), .Z(O[817]) );
  AND U611 ( .A(S), .B(n408), .Z(n407) );
  XOR U612 ( .A(B[817]), .B(A[817]), .Z(n408) );
  XOR U613 ( .A(A[816]), .B(n409), .Z(O[816]) );
  AND U614 ( .A(S), .B(n410), .Z(n409) );
  XOR U615 ( .A(B[816]), .B(A[816]), .Z(n410) );
  XOR U616 ( .A(A[815]), .B(n411), .Z(O[815]) );
  AND U617 ( .A(S), .B(n412), .Z(n411) );
  XOR U618 ( .A(B[815]), .B(A[815]), .Z(n412) );
  XOR U619 ( .A(A[814]), .B(n413), .Z(O[814]) );
  AND U620 ( .A(S), .B(n414), .Z(n413) );
  XOR U621 ( .A(B[814]), .B(A[814]), .Z(n414) );
  XOR U622 ( .A(A[813]), .B(n415), .Z(O[813]) );
  AND U623 ( .A(S), .B(n416), .Z(n415) );
  XOR U624 ( .A(B[813]), .B(A[813]), .Z(n416) );
  XOR U625 ( .A(A[812]), .B(n417), .Z(O[812]) );
  AND U626 ( .A(S), .B(n418), .Z(n417) );
  XOR U627 ( .A(B[812]), .B(A[812]), .Z(n418) );
  XOR U628 ( .A(A[811]), .B(n419), .Z(O[811]) );
  AND U629 ( .A(S), .B(n420), .Z(n419) );
  XOR U630 ( .A(B[811]), .B(A[811]), .Z(n420) );
  XOR U631 ( .A(A[810]), .B(n421), .Z(O[810]) );
  AND U632 ( .A(S), .B(n422), .Z(n421) );
  XOR U633 ( .A(B[810]), .B(A[810]), .Z(n422) );
  XOR U634 ( .A(A[80]), .B(n423), .Z(O[80]) );
  AND U635 ( .A(S), .B(n424), .Z(n423) );
  XOR U636 ( .A(B[80]), .B(A[80]), .Z(n424) );
  XOR U637 ( .A(A[809]), .B(n425), .Z(O[809]) );
  AND U638 ( .A(S), .B(n426), .Z(n425) );
  XOR U639 ( .A(B[809]), .B(A[809]), .Z(n426) );
  XOR U640 ( .A(A[808]), .B(n427), .Z(O[808]) );
  AND U641 ( .A(S), .B(n428), .Z(n427) );
  XOR U642 ( .A(B[808]), .B(A[808]), .Z(n428) );
  XOR U643 ( .A(A[807]), .B(n429), .Z(O[807]) );
  AND U644 ( .A(S), .B(n430), .Z(n429) );
  XOR U645 ( .A(B[807]), .B(A[807]), .Z(n430) );
  XOR U646 ( .A(A[806]), .B(n431), .Z(O[806]) );
  AND U647 ( .A(S), .B(n432), .Z(n431) );
  XOR U648 ( .A(B[806]), .B(A[806]), .Z(n432) );
  XOR U649 ( .A(A[805]), .B(n433), .Z(O[805]) );
  AND U650 ( .A(S), .B(n434), .Z(n433) );
  XOR U651 ( .A(B[805]), .B(A[805]), .Z(n434) );
  XOR U652 ( .A(A[804]), .B(n435), .Z(O[804]) );
  AND U653 ( .A(S), .B(n436), .Z(n435) );
  XOR U654 ( .A(B[804]), .B(A[804]), .Z(n436) );
  XOR U655 ( .A(A[803]), .B(n437), .Z(O[803]) );
  AND U656 ( .A(S), .B(n438), .Z(n437) );
  XOR U657 ( .A(B[803]), .B(A[803]), .Z(n438) );
  XOR U658 ( .A(A[802]), .B(n439), .Z(O[802]) );
  AND U659 ( .A(S), .B(n440), .Z(n439) );
  XOR U660 ( .A(B[802]), .B(A[802]), .Z(n440) );
  XOR U661 ( .A(A[801]), .B(n441), .Z(O[801]) );
  AND U662 ( .A(S), .B(n442), .Z(n441) );
  XOR U663 ( .A(B[801]), .B(A[801]), .Z(n442) );
  XOR U664 ( .A(A[800]), .B(n443), .Z(O[800]) );
  AND U665 ( .A(S), .B(n444), .Z(n443) );
  XOR U666 ( .A(B[800]), .B(A[800]), .Z(n444) );
  XOR U667 ( .A(A[7]), .B(n445), .Z(O[7]) );
  AND U668 ( .A(S), .B(n446), .Z(n445) );
  XOR U669 ( .A(B[7]), .B(A[7]), .Z(n446) );
  XOR U670 ( .A(A[79]), .B(n447), .Z(O[79]) );
  AND U671 ( .A(S), .B(n448), .Z(n447) );
  XOR U672 ( .A(B[79]), .B(A[79]), .Z(n448) );
  XOR U673 ( .A(A[799]), .B(n449), .Z(O[799]) );
  AND U674 ( .A(S), .B(n450), .Z(n449) );
  XOR U675 ( .A(B[799]), .B(A[799]), .Z(n450) );
  XOR U676 ( .A(A[798]), .B(n451), .Z(O[798]) );
  AND U677 ( .A(S), .B(n452), .Z(n451) );
  XOR U678 ( .A(B[798]), .B(A[798]), .Z(n452) );
  XOR U679 ( .A(A[797]), .B(n453), .Z(O[797]) );
  AND U680 ( .A(S), .B(n454), .Z(n453) );
  XOR U681 ( .A(B[797]), .B(A[797]), .Z(n454) );
  XOR U682 ( .A(A[796]), .B(n455), .Z(O[796]) );
  AND U683 ( .A(S), .B(n456), .Z(n455) );
  XOR U684 ( .A(B[796]), .B(A[796]), .Z(n456) );
  XOR U685 ( .A(A[795]), .B(n457), .Z(O[795]) );
  AND U686 ( .A(S), .B(n458), .Z(n457) );
  XOR U687 ( .A(B[795]), .B(A[795]), .Z(n458) );
  XOR U688 ( .A(A[794]), .B(n459), .Z(O[794]) );
  AND U689 ( .A(S), .B(n460), .Z(n459) );
  XOR U690 ( .A(B[794]), .B(A[794]), .Z(n460) );
  XOR U691 ( .A(A[793]), .B(n461), .Z(O[793]) );
  AND U692 ( .A(S), .B(n462), .Z(n461) );
  XOR U693 ( .A(B[793]), .B(A[793]), .Z(n462) );
  XOR U694 ( .A(A[792]), .B(n463), .Z(O[792]) );
  AND U695 ( .A(S), .B(n464), .Z(n463) );
  XOR U696 ( .A(B[792]), .B(A[792]), .Z(n464) );
  XOR U697 ( .A(A[791]), .B(n465), .Z(O[791]) );
  AND U698 ( .A(S), .B(n466), .Z(n465) );
  XOR U699 ( .A(B[791]), .B(A[791]), .Z(n466) );
  XOR U700 ( .A(A[790]), .B(n467), .Z(O[790]) );
  AND U701 ( .A(S), .B(n468), .Z(n467) );
  XOR U702 ( .A(B[790]), .B(A[790]), .Z(n468) );
  XOR U703 ( .A(A[78]), .B(n469), .Z(O[78]) );
  AND U704 ( .A(S), .B(n470), .Z(n469) );
  XOR U705 ( .A(B[78]), .B(A[78]), .Z(n470) );
  XOR U706 ( .A(A[789]), .B(n471), .Z(O[789]) );
  AND U707 ( .A(S), .B(n472), .Z(n471) );
  XOR U708 ( .A(B[789]), .B(A[789]), .Z(n472) );
  XOR U709 ( .A(A[788]), .B(n473), .Z(O[788]) );
  AND U710 ( .A(S), .B(n474), .Z(n473) );
  XOR U711 ( .A(B[788]), .B(A[788]), .Z(n474) );
  XOR U712 ( .A(A[787]), .B(n475), .Z(O[787]) );
  AND U713 ( .A(S), .B(n476), .Z(n475) );
  XOR U714 ( .A(B[787]), .B(A[787]), .Z(n476) );
  XOR U715 ( .A(A[786]), .B(n477), .Z(O[786]) );
  AND U716 ( .A(S), .B(n478), .Z(n477) );
  XOR U717 ( .A(B[786]), .B(A[786]), .Z(n478) );
  XOR U718 ( .A(A[785]), .B(n479), .Z(O[785]) );
  AND U719 ( .A(S), .B(n480), .Z(n479) );
  XOR U720 ( .A(B[785]), .B(A[785]), .Z(n480) );
  XOR U721 ( .A(A[784]), .B(n481), .Z(O[784]) );
  AND U722 ( .A(S), .B(n482), .Z(n481) );
  XOR U723 ( .A(B[784]), .B(A[784]), .Z(n482) );
  XOR U724 ( .A(A[783]), .B(n483), .Z(O[783]) );
  AND U725 ( .A(S), .B(n484), .Z(n483) );
  XOR U726 ( .A(B[783]), .B(A[783]), .Z(n484) );
  XOR U727 ( .A(A[782]), .B(n485), .Z(O[782]) );
  AND U728 ( .A(S), .B(n486), .Z(n485) );
  XOR U729 ( .A(B[782]), .B(A[782]), .Z(n486) );
  XOR U730 ( .A(A[781]), .B(n487), .Z(O[781]) );
  AND U731 ( .A(S), .B(n488), .Z(n487) );
  XOR U732 ( .A(B[781]), .B(A[781]), .Z(n488) );
  XOR U733 ( .A(A[780]), .B(n489), .Z(O[780]) );
  AND U734 ( .A(S), .B(n490), .Z(n489) );
  XOR U735 ( .A(B[780]), .B(A[780]), .Z(n490) );
  XOR U736 ( .A(A[77]), .B(n491), .Z(O[77]) );
  AND U737 ( .A(S), .B(n492), .Z(n491) );
  XOR U738 ( .A(B[77]), .B(A[77]), .Z(n492) );
  XOR U739 ( .A(A[779]), .B(n493), .Z(O[779]) );
  AND U740 ( .A(S), .B(n494), .Z(n493) );
  XOR U741 ( .A(B[779]), .B(A[779]), .Z(n494) );
  XOR U742 ( .A(A[778]), .B(n495), .Z(O[778]) );
  AND U743 ( .A(S), .B(n496), .Z(n495) );
  XOR U744 ( .A(B[778]), .B(A[778]), .Z(n496) );
  XOR U745 ( .A(A[777]), .B(n497), .Z(O[777]) );
  AND U746 ( .A(S), .B(n498), .Z(n497) );
  XOR U747 ( .A(B[777]), .B(A[777]), .Z(n498) );
  XOR U748 ( .A(A[776]), .B(n499), .Z(O[776]) );
  AND U749 ( .A(S), .B(n500), .Z(n499) );
  XOR U750 ( .A(B[776]), .B(A[776]), .Z(n500) );
  XOR U751 ( .A(A[775]), .B(n501), .Z(O[775]) );
  AND U752 ( .A(S), .B(n502), .Z(n501) );
  XOR U753 ( .A(B[775]), .B(A[775]), .Z(n502) );
  XOR U754 ( .A(A[774]), .B(n503), .Z(O[774]) );
  AND U755 ( .A(S), .B(n504), .Z(n503) );
  XOR U756 ( .A(B[774]), .B(A[774]), .Z(n504) );
  XOR U757 ( .A(A[773]), .B(n505), .Z(O[773]) );
  AND U758 ( .A(S), .B(n506), .Z(n505) );
  XOR U759 ( .A(B[773]), .B(A[773]), .Z(n506) );
  XOR U760 ( .A(A[772]), .B(n507), .Z(O[772]) );
  AND U761 ( .A(S), .B(n508), .Z(n507) );
  XOR U762 ( .A(B[772]), .B(A[772]), .Z(n508) );
  XOR U763 ( .A(A[771]), .B(n509), .Z(O[771]) );
  AND U764 ( .A(S), .B(n510), .Z(n509) );
  XOR U765 ( .A(B[771]), .B(A[771]), .Z(n510) );
  XOR U766 ( .A(A[770]), .B(n511), .Z(O[770]) );
  AND U767 ( .A(S), .B(n512), .Z(n511) );
  XOR U768 ( .A(B[770]), .B(A[770]), .Z(n512) );
  XOR U769 ( .A(A[76]), .B(n513), .Z(O[76]) );
  AND U770 ( .A(S), .B(n514), .Z(n513) );
  XOR U771 ( .A(B[76]), .B(A[76]), .Z(n514) );
  XOR U772 ( .A(A[769]), .B(n515), .Z(O[769]) );
  AND U773 ( .A(S), .B(n516), .Z(n515) );
  XOR U774 ( .A(B[769]), .B(A[769]), .Z(n516) );
  XOR U775 ( .A(A[768]), .B(n517), .Z(O[768]) );
  AND U776 ( .A(S), .B(n518), .Z(n517) );
  XOR U777 ( .A(B[768]), .B(A[768]), .Z(n518) );
  XOR U778 ( .A(A[767]), .B(n519), .Z(O[767]) );
  AND U779 ( .A(S), .B(n520), .Z(n519) );
  XOR U780 ( .A(B[767]), .B(A[767]), .Z(n520) );
  XOR U781 ( .A(A[766]), .B(n521), .Z(O[766]) );
  AND U782 ( .A(S), .B(n522), .Z(n521) );
  XOR U783 ( .A(B[766]), .B(A[766]), .Z(n522) );
  XOR U784 ( .A(A[765]), .B(n523), .Z(O[765]) );
  AND U785 ( .A(S), .B(n524), .Z(n523) );
  XOR U786 ( .A(B[765]), .B(A[765]), .Z(n524) );
  XOR U787 ( .A(A[764]), .B(n525), .Z(O[764]) );
  AND U788 ( .A(S), .B(n526), .Z(n525) );
  XOR U789 ( .A(B[764]), .B(A[764]), .Z(n526) );
  XOR U790 ( .A(A[763]), .B(n527), .Z(O[763]) );
  AND U791 ( .A(S), .B(n528), .Z(n527) );
  XOR U792 ( .A(B[763]), .B(A[763]), .Z(n528) );
  XOR U793 ( .A(A[762]), .B(n529), .Z(O[762]) );
  AND U794 ( .A(S), .B(n530), .Z(n529) );
  XOR U795 ( .A(B[762]), .B(A[762]), .Z(n530) );
  XOR U796 ( .A(A[761]), .B(n531), .Z(O[761]) );
  AND U797 ( .A(S), .B(n532), .Z(n531) );
  XOR U798 ( .A(B[761]), .B(A[761]), .Z(n532) );
  XOR U799 ( .A(A[760]), .B(n533), .Z(O[760]) );
  AND U800 ( .A(S), .B(n534), .Z(n533) );
  XOR U801 ( .A(B[760]), .B(A[760]), .Z(n534) );
  XOR U802 ( .A(A[75]), .B(n535), .Z(O[75]) );
  AND U803 ( .A(S), .B(n536), .Z(n535) );
  XOR U804 ( .A(B[75]), .B(A[75]), .Z(n536) );
  XOR U805 ( .A(A[759]), .B(n537), .Z(O[759]) );
  AND U806 ( .A(S), .B(n538), .Z(n537) );
  XOR U807 ( .A(B[759]), .B(A[759]), .Z(n538) );
  XOR U808 ( .A(A[758]), .B(n539), .Z(O[758]) );
  AND U809 ( .A(S), .B(n540), .Z(n539) );
  XOR U810 ( .A(B[758]), .B(A[758]), .Z(n540) );
  XOR U811 ( .A(A[757]), .B(n541), .Z(O[757]) );
  AND U812 ( .A(S), .B(n542), .Z(n541) );
  XOR U813 ( .A(B[757]), .B(A[757]), .Z(n542) );
  XOR U814 ( .A(A[756]), .B(n543), .Z(O[756]) );
  AND U815 ( .A(S), .B(n544), .Z(n543) );
  XOR U816 ( .A(B[756]), .B(A[756]), .Z(n544) );
  XOR U817 ( .A(A[755]), .B(n545), .Z(O[755]) );
  AND U818 ( .A(S), .B(n546), .Z(n545) );
  XOR U819 ( .A(B[755]), .B(A[755]), .Z(n546) );
  XOR U820 ( .A(A[754]), .B(n547), .Z(O[754]) );
  AND U821 ( .A(S), .B(n548), .Z(n547) );
  XOR U822 ( .A(B[754]), .B(A[754]), .Z(n548) );
  XOR U823 ( .A(A[753]), .B(n549), .Z(O[753]) );
  AND U824 ( .A(S), .B(n550), .Z(n549) );
  XOR U825 ( .A(B[753]), .B(A[753]), .Z(n550) );
  XOR U826 ( .A(A[752]), .B(n551), .Z(O[752]) );
  AND U827 ( .A(S), .B(n552), .Z(n551) );
  XOR U828 ( .A(B[752]), .B(A[752]), .Z(n552) );
  XOR U829 ( .A(A[751]), .B(n553), .Z(O[751]) );
  AND U830 ( .A(S), .B(n554), .Z(n553) );
  XOR U831 ( .A(B[751]), .B(A[751]), .Z(n554) );
  XOR U832 ( .A(A[750]), .B(n555), .Z(O[750]) );
  AND U833 ( .A(S), .B(n556), .Z(n555) );
  XOR U834 ( .A(B[750]), .B(A[750]), .Z(n556) );
  XOR U835 ( .A(A[74]), .B(n557), .Z(O[74]) );
  AND U836 ( .A(S), .B(n558), .Z(n557) );
  XOR U837 ( .A(B[74]), .B(A[74]), .Z(n558) );
  XOR U838 ( .A(A[749]), .B(n559), .Z(O[749]) );
  AND U839 ( .A(S), .B(n560), .Z(n559) );
  XOR U840 ( .A(B[749]), .B(A[749]), .Z(n560) );
  XOR U841 ( .A(A[748]), .B(n561), .Z(O[748]) );
  AND U842 ( .A(S), .B(n562), .Z(n561) );
  XOR U843 ( .A(B[748]), .B(A[748]), .Z(n562) );
  XOR U844 ( .A(A[747]), .B(n563), .Z(O[747]) );
  AND U845 ( .A(S), .B(n564), .Z(n563) );
  XOR U846 ( .A(B[747]), .B(A[747]), .Z(n564) );
  XOR U847 ( .A(A[746]), .B(n565), .Z(O[746]) );
  AND U848 ( .A(S), .B(n566), .Z(n565) );
  XOR U849 ( .A(B[746]), .B(A[746]), .Z(n566) );
  XOR U850 ( .A(A[745]), .B(n567), .Z(O[745]) );
  AND U851 ( .A(S), .B(n568), .Z(n567) );
  XOR U852 ( .A(B[745]), .B(A[745]), .Z(n568) );
  XOR U853 ( .A(A[744]), .B(n569), .Z(O[744]) );
  AND U854 ( .A(S), .B(n570), .Z(n569) );
  XOR U855 ( .A(B[744]), .B(A[744]), .Z(n570) );
  XOR U856 ( .A(A[743]), .B(n571), .Z(O[743]) );
  AND U857 ( .A(S), .B(n572), .Z(n571) );
  XOR U858 ( .A(B[743]), .B(A[743]), .Z(n572) );
  XOR U859 ( .A(A[742]), .B(n573), .Z(O[742]) );
  AND U860 ( .A(S), .B(n574), .Z(n573) );
  XOR U861 ( .A(B[742]), .B(A[742]), .Z(n574) );
  XOR U862 ( .A(A[741]), .B(n575), .Z(O[741]) );
  AND U863 ( .A(S), .B(n576), .Z(n575) );
  XOR U864 ( .A(B[741]), .B(A[741]), .Z(n576) );
  XOR U865 ( .A(A[740]), .B(n577), .Z(O[740]) );
  AND U866 ( .A(S), .B(n578), .Z(n577) );
  XOR U867 ( .A(B[740]), .B(A[740]), .Z(n578) );
  XOR U868 ( .A(A[73]), .B(n579), .Z(O[73]) );
  AND U869 ( .A(S), .B(n580), .Z(n579) );
  XOR U870 ( .A(B[73]), .B(A[73]), .Z(n580) );
  XOR U871 ( .A(A[739]), .B(n581), .Z(O[739]) );
  AND U872 ( .A(S), .B(n582), .Z(n581) );
  XOR U873 ( .A(B[739]), .B(A[739]), .Z(n582) );
  XOR U874 ( .A(A[738]), .B(n583), .Z(O[738]) );
  AND U875 ( .A(S), .B(n584), .Z(n583) );
  XOR U876 ( .A(B[738]), .B(A[738]), .Z(n584) );
  XOR U877 ( .A(A[737]), .B(n585), .Z(O[737]) );
  AND U878 ( .A(S), .B(n586), .Z(n585) );
  XOR U879 ( .A(B[737]), .B(A[737]), .Z(n586) );
  XOR U880 ( .A(A[736]), .B(n587), .Z(O[736]) );
  AND U881 ( .A(S), .B(n588), .Z(n587) );
  XOR U882 ( .A(B[736]), .B(A[736]), .Z(n588) );
  XOR U883 ( .A(A[735]), .B(n589), .Z(O[735]) );
  AND U884 ( .A(S), .B(n590), .Z(n589) );
  XOR U885 ( .A(B[735]), .B(A[735]), .Z(n590) );
  XOR U886 ( .A(A[734]), .B(n591), .Z(O[734]) );
  AND U887 ( .A(S), .B(n592), .Z(n591) );
  XOR U888 ( .A(B[734]), .B(A[734]), .Z(n592) );
  XOR U889 ( .A(A[733]), .B(n593), .Z(O[733]) );
  AND U890 ( .A(S), .B(n594), .Z(n593) );
  XOR U891 ( .A(B[733]), .B(A[733]), .Z(n594) );
  XOR U892 ( .A(A[732]), .B(n595), .Z(O[732]) );
  AND U893 ( .A(S), .B(n596), .Z(n595) );
  XOR U894 ( .A(B[732]), .B(A[732]), .Z(n596) );
  XOR U895 ( .A(A[731]), .B(n597), .Z(O[731]) );
  AND U896 ( .A(S), .B(n598), .Z(n597) );
  XOR U897 ( .A(B[731]), .B(A[731]), .Z(n598) );
  XOR U898 ( .A(A[730]), .B(n599), .Z(O[730]) );
  AND U899 ( .A(S), .B(n600), .Z(n599) );
  XOR U900 ( .A(B[730]), .B(A[730]), .Z(n600) );
  XOR U901 ( .A(A[72]), .B(n601), .Z(O[72]) );
  AND U902 ( .A(S), .B(n602), .Z(n601) );
  XOR U903 ( .A(B[72]), .B(A[72]), .Z(n602) );
  XOR U904 ( .A(A[729]), .B(n603), .Z(O[729]) );
  AND U905 ( .A(S), .B(n604), .Z(n603) );
  XOR U906 ( .A(B[729]), .B(A[729]), .Z(n604) );
  XOR U907 ( .A(A[728]), .B(n605), .Z(O[728]) );
  AND U908 ( .A(S), .B(n606), .Z(n605) );
  XOR U909 ( .A(B[728]), .B(A[728]), .Z(n606) );
  XOR U910 ( .A(A[727]), .B(n607), .Z(O[727]) );
  AND U911 ( .A(S), .B(n608), .Z(n607) );
  XOR U912 ( .A(B[727]), .B(A[727]), .Z(n608) );
  XOR U913 ( .A(A[726]), .B(n609), .Z(O[726]) );
  AND U914 ( .A(S), .B(n610), .Z(n609) );
  XOR U915 ( .A(B[726]), .B(A[726]), .Z(n610) );
  XOR U916 ( .A(A[725]), .B(n611), .Z(O[725]) );
  AND U917 ( .A(S), .B(n612), .Z(n611) );
  XOR U918 ( .A(B[725]), .B(A[725]), .Z(n612) );
  XOR U919 ( .A(A[724]), .B(n613), .Z(O[724]) );
  AND U920 ( .A(S), .B(n614), .Z(n613) );
  XOR U921 ( .A(B[724]), .B(A[724]), .Z(n614) );
  XOR U922 ( .A(A[723]), .B(n615), .Z(O[723]) );
  AND U923 ( .A(S), .B(n616), .Z(n615) );
  XOR U924 ( .A(B[723]), .B(A[723]), .Z(n616) );
  XOR U925 ( .A(A[722]), .B(n617), .Z(O[722]) );
  AND U926 ( .A(S), .B(n618), .Z(n617) );
  XOR U927 ( .A(B[722]), .B(A[722]), .Z(n618) );
  XOR U928 ( .A(A[721]), .B(n619), .Z(O[721]) );
  AND U929 ( .A(S), .B(n620), .Z(n619) );
  XOR U930 ( .A(B[721]), .B(A[721]), .Z(n620) );
  XOR U931 ( .A(A[720]), .B(n621), .Z(O[720]) );
  AND U932 ( .A(S), .B(n622), .Z(n621) );
  XOR U933 ( .A(B[720]), .B(A[720]), .Z(n622) );
  XOR U934 ( .A(A[71]), .B(n623), .Z(O[71]) );
  AND U935 ( .A(S), .B(n624), .Z(n623) );
  XOR U936 ( .A(B[71]), .B(A[71]), .Z(n624) );
  XOR U937 ( .A(A[719]), .B(n625), .Z(O[719]) );
  AND U938 ( .A(S), .B(n626), .Z(n625) );
  XOR U939 ( .A(B[719]), .B(A[719]), .Z(n626) );
  XOR U940 ( .A(A[718]), .B(n627), .Z(O[718]) );
  AND U941 ( .A(S), .B(n628), .Z(n627) );
  XOR U942 ( .A(B[718]), .B(A[718]), .Z(n628) );
  XOR U943 ( .A(A[717]), .B(n629), .Z(O[717]) );
  AND U944 ( .A(S), .B(n630), .Z(n629) );
  XOR U945 ( .A(B[717]), .B(A[717]), .Z(n630) );
  XOR U946 ( .A(A[716]), .B(n631), .Z(O[716]) );
  AND U947 ( .A(S), .B(n632), .Z(n631) );
  XOR U948 ( .A(B[716]), .B(A[716]), .Z(n632) );
  XOR U949 ( .A(A[715]), .B(n633), .Z(O[715]) );
  AND U950 ( .A(S), .B(n634), .Z(n633) );
  XOR U951 ( .A(B[715]), .B(A[715]), .Z(n634) );
  XOR U952 ( .A(A[714]), .B(n635), .Z(O[714]) );
  AND U953 ( .A(S), .B(n636), .Z(n635) );
  XOR U954 ( .A(B[714]), .B(A[714]), .Z(n636) );
  XOR U955 ( .A(A[713]), .B(n637), .Z(O[713]) );
  AND U956 ( .A(S), .B(n638), .Z(n637) );
  XOR U957 ( .A(B[713]), .B(A[713]), .Z(n638) );
  XOR U958 ( .A(A[712]), .B(n639), .Z(O[712]) );
  AND U959 ( .A(S), .B(n640), .Z(n639) );
  XOR U960 ( .A(B[712]), .B(A[712]), .Z(n640) );
  XOR U961 ( .A(A[711]), .B(n641), .Z(O[711]) );
  AND U962 ( .A(S), .B(n642), .Z(n641) );
  XOR U963 ( .A(B[711]), .B(A[711]), .Z(n642) );
  XOR U964 ( .A(A[710]), .B(n643), .Z(O[710]) );
  AND U965 ( .A(S), .B(n644), .Z(n643) );
  XOR U966 ( .A(B[710]), .B(A[710]), .Z(n644) );
  XOR U967 ( .A(A[70]), .B(n645), .Z(O[70]) );
  AND U968 ( .A(S), .B(n646), .Z(n645) );
  XOR U969 ( .A(B[70]), .B(A[70]), .Z(n646) );
  XOR U970 ( .A(A[709]), .B(n647), .Z(O[709]) );
  AND U971 ( .A(S), .B(n648), .Z(n647) );
  XOR U972 ( .A(B[709]), .B(A[709]), .Z(n648) );
  XOR U973 ( .A(A[708]), .B(n649), .Z(O[708]) );
  AND U974 ( .A(S), .B(n650), .Z(n649) );
  XOR U975 ( .A(B[708]), .B(A[708]), .Z(n650) );
  XOR U976 ( .A(A[707]), .B(n651), .Z(O[707]) );
  AND U977 ( .A(S), .B(n652), .Z(n651) );
  XOR U978 ( .A(B[707]), .B(A[707]), .Z(n652) );
  XOR U979 ( .A(A[706]), .B(n653), .Z(O[706]) );
  AND U980 ( .A(S), .B(n654), .Z(n653) );
  XOR U981 ( .A(B[706]), .B(A[706]), .Z(n654) );
  XOR U982 ( .A(A[705]), .B(n655), .Z(O[705]) );
  AND U983 ( .A(S), .B(n656), .Z(n655) );
  XOR U984 ( .A(B[705]), .B(A[705]), .Z(n656) );
  XOR U985 ( .A(A[704]), .B(n657), .Z(O[704]) );
  AND U986 ( .A(S), .B(n658), .Z(n657) );
  XOR U987 ( .A(B[704]), .B(A[704]), .Z(n658) );
  XOR U988 ( .A(A[703]), .B(n659), .Z(O[703]) );
  AND U989 ( .A(S), .B(n660), .Z(n659) );
  XOR U990 ( .A(B[703]), .B(A[703]), .Z(n660) );
  XOR U991 ( .A(A[702]), .B(n661), .Z(O[702]) );
  AND U992 ( .A(S), .B(n662), .Z(n661) );
  XOR U993 ( .A(B[702]), .B(A[702]), .Z(n662) );
  XOR U994 ( .A(A[701]), .B(n663), .Z(O[701]) );
  AND U995 ( .A(S), .B(n664), .Z(n663) );
  XOR U996 ( .A(B[701]), .B(A[701]), .Z(n664) );
  XOR U997 ( .A(A[700]), .B(n665), .Z(O[700]) );
  AND U998 ( .A(S), .B(n666), .Z(n665) );
  XOR U999 ( .A(B[700]), .B(A[700]), .Z(n666) );
  XOR U1000 ( .A(A[6]), .B(n667), .Z(O[6]) );
  AND U1001 ( .A(S), .B(n668), .Z(n667) );
  XOR U1002 ( .A(B[6]), .B(A[6]), .Z(n668) );
  XOR U1003 ( .A(A[69]), .B(n669), .Z(O[69]) );
  AND U1004 ( .A(S), .B(n670), .Z(n669) );
  XOR U1005 ( .A(B[69]), .B(A[69]), .Z(n670) );
  XOR U1006 ( .A(A[699]), .B(n671), .Z(O[699]) );
  AND U1007 ( .A(S), .B(n672), .Z(n671) );
  XOR U1008 ( .A(B[699]), .B(A[699]), .Z(n672) );
  XOR U1009 ( .A(A[698]), .B(n673), .Z(O[698]) );
  AND U1010 ( .A(S), .B(n674), .Z(n673) );
  XOR U1011 ( .A(B[698]), .B(A[698]), .Z(n674) );
  XOR U1012 ( .A(A[697]), .B(n675), .Z(O[697]) );
  AND U1013 ( .A(S), .B(n676), .Z(n675) );
  XOR U1014 ( .A(B[697]), .B(A[697]), .Z(n676) );
  XOR U1015 ( .A(A[696]), .B(n677), .Z(O[696]) );
  AND U1016 ( .A(S), .B(n678), .Z(n677) );
  XOR U1017 ( .A(B[696]), .B(A[696]), .Z(n678) );
  XOR U1018 ( .A(A[695]), .B(n679), .Z(O[695]) );
  AND U1019 ( .A(S), .B(n680), .Z(n679) );
  XOR U1020 ( .A(B[695]), .B(A[695]), .Z(n680) );
  XOR U1021 ( .A(A[694]), .B(n681), .Z(O[694]) );
  AND U1022 ( .A(S), .B(n682), .Z(n681) );
  XOR U1023 ( .A(B[694]), .B(A[694]), .Z(n682) );
  XOR U1024 ( .A(A[693]), .B(n683), .Z(O[693]) );
  AND U1025 ( .A(S), .B(n684), .Z(n683) );
  XOR U1026 ( .A(B[693]), .B(A[693]), .Z(n684) );
  XOR U1027 ( .A(A[692]), .B(n685), .Z(O[692]) );
  AND U1028 ( .A(S), .B(n686), .Z(n685) );
  XOR U1029 ( .A(B[692]), .B(A[692]), .Z(n686) );
  XOR U1030 ( .A(A[691]), .B(n687), .Z(O[691]) );
  AND U1031 ( .A(S), .B(n688), .Z(n687) );
  XOR U1032 ( .A(B[691]), .B(A[691]), .Z(n688) );
  XOR U1033 ( .A(A[690]), .B(n689), .Z(O[690]) );
  AND U1034 ( .A(S), .B(n690), .Z(n689) );
  XOR U1035 ( .A(B[690]), .B(A[690]), .Z(n690) );
  XOR U1036 ( .A(A[68]), .B(n691), .Z(O[68]) );
  AND U1037 ( .A(S), .B(n692), .Z(n691) );
  XOR U1038 ( .A(B[68]), .B(A[68]), .Z(n692) );
  XOR U1039 ( .A(A[689]), .B(n693), .Z(O[689]) );
  AND U1040 ( .A(S), .B(n694), .Z(n693) );
  XOR U1041 ( .A(B[689]), .B(A[689]), .Z(n694) );
  XOR U1042 ( .A(A[688]), .B(n695), .Z(O[688]) );
  AND U1043 ( .A(S), .B(n696), .Z(n695) );
  XOR U1044 ( .A(B[688]), .B(A[688]), .Z(n696) );
  XOR U1045 ( .A(A[687]), .B(n697), .Z(O[687]) );
  AND U1046 ( .A(S), .B(n698), .Z(n697) );
  XOR U1047 ( .A(B[687]), .B(A[687]), .Z(n698) );
  XOR U1048 ( .A(A[686]), .B(n699), .Z(O[686]) );
  AND U1049 ( .A(S), .B(n700), .Z(n699) );
  XOR U1050 ( .A(B[686]), .B(A[686]), .Z(n700) );
  XOR U1051 ( .A(A[685]), .B(n701), .Z(O[685]) );
  AND U1052 ( .A(S), .B(n702), .Z(n701) );
  XOR U1053 ( .A(B[685]), .B(A[685]), .Z(n702) );
  XOR U1054 ( .A(A[684]), .B(n703), .Z(O[684]) );
  AND U1055 ( .A(S), .B(n704), .Z(n703) );
  XOR U1056 ( .A(B[684]), .B(A[684]), .Z(n704) );
  XOR U1057 ( .A(A[683]), .B(n705), .Z(O[683]) );
  AND U1058 ( .A(S), .B(n706), .Z(n705) );
  XOR U1059 ( .A(B[683]), .B(A[683]), .Z(n706) );
  XOR U1060 ( .A(A[682]), .B(n707), .Z(O[682]) );
  AND U1061 ( .A(S), .B(n708), .Z(n707) );
  XOR U1062 ( .A(B[682]), .B(A[682]), .Z(n708) );
  XOR U1063 ( .A(A[681]), .B(n709), .Z(O[681]) );
  AND U1064 ( .A(S), .B(n710), .Z(n709) );
  XOR U1065 ( .A(B[681]), .B(A[681]), .Z(n710) );
  XOR U1066 ( .A(A[680]), .B(n711), .Z(O[680]) );
  AND U1067 ( .A(S), .B(n712), .Z(n711) );
  XOR U1068 ( .A(B[680]), .B(A[680]), .Z(n712) );
  XOR U1069 ( .A(A[67]), .B(n713), .Z(O[67]) );
  AND U1070 ( .A(S), .B(n714), .Z(n713) );
  XOR U1071 ( .A(B[67]), .B(A[67]), .Z(n714) );
  XOR U1072 ( .A(A[679]), .B(n715), .Z(O[679]) );
  AND U1073 ( .A(S), .B(n716), .Z(n715) );
  XOR U1074 ( .A(B[679]), .B(A[679]), .Z(n716) );
  XOR U1075 ( .A(A[678]), .B(n717), .Z(O[678]) );
  AND U1076 ( .A(S), .B(n718), .Z(n717) );
  XOR U1077 ( .A(B[678]), .B(A[678]), .Z(n718) );
  XOR U1078 ( .A(A[677]), .B(n719), .Z(O[677]) );
  AND U1079 ( .A(S), .B(n720), .Z(n719) );
  XOR U1080 ( .A(B[677]), .B(A[677]), .Z(n720) );
  XOR U1081 ( .A(A[676]), .B(n721), .Z(O[676]) );
  AND U1082 ( .A(S), .B(n722), .Z(n721) );
  XOR U1083 ( .A(B[676]), .B(A[676]), .Z(n722) );
  XOR U1084 ( .A(A[675]), .B(n723), .Z(O[675]) );
  AND U1085 ( .A(S), .B(n724), .Z(n723) );
  XOR U1086 ( .A(B[675]), .B(A[675]), .Z(n724) );
  XOR U1087 ( .A(A[674]), .B(n725), .Z(O[674]) );
  AND U1088 ( .A(S), .B(n726), .Z(n725) );
  XOR U1089 ( .A(B[674]), .B(A[674]), .Z(n726) );
  XOR U1090 ( .A(A[673]), .B(n727), .Z(O[673]) );
  AND U1091 ( .A(S), .B(n728), .Z(n727) );
  XOR U1092 ( .A(B[673]), .B(A[673]), .Z(n728) );
  XOR U1093 ( .A(A[672]), .B(n729), .Z(O[672]) );
  AND U1094 ( .A(S), .B(n730), .Z(n729) );
  XOR U1095 ( .A(B[672]), .B(A[672]), .Z(n730) );
  XOR U1096 ( .A(A[671]), .B(n731), .Z(O[671]) );
  AND U1097 ( .A(S), .B(n732), .Z(n731) );
  XOR U1098 ( .A(B[671]), .B(A[671]), .Z(n732) );
  XOR U1099 ( .A(A[670]), .B(n733), .Z(O[670]) );
  AND U1100 ( .A(S), .B(n734), .Z(n733) );
  XOR U1101 ( .A(B[670]), .B(A[670]), .Z(n734) );
  XOR U1102 ( .A(A[66]), .B(n735), .Z(O[66]) );
  AND U1103 ( .A(S), .B(n736), .Z(n735) );
  XOR U1104 ( .A(B[66]), .B(A[66]), .Z(n736) );
  XOR U1105 ( .A(A[669]), .B(n737), .Z(O[669]) );
  AND U1106 ( .A(S), .B(n738), .Z(n737) );
  XOR U1107 ( .A(B[669]), .B(A[669]), .Z(n738) );
  XOR U1108 ( .A(A[668]), .B(n739), .Z(O[668]) );
  AND U1109 ( .A(S), .B(n740), .Z(n739) );
  XOR U1110 ( .A(B[668]), .B(A[668]), .Z(n740) );
  XOR U1111 ( .A(A[667]), .B(n741), .Z(O[667]) );
  AND U1112 ( .A(S), .B(n742), .Z(n741) );
  XOR U1113 ( .A(B[667]), .B(A[667]), .Z(n742) );
  XOR U1114 ( .A(A[666]), .B(n743), .Z(O[666]) );
  AND U1115 ( .A(S), .B(n744), .Z(n743) );
  XOR U1116 ( .A(B[666]), .B(A[666]), .Z(n744) );
  XOR U1117 ( .A(A[665]), .B(n745), .Z(O[665]) );
  AND U1118 ( .A(S), .B(n746), .Z(n745) );
  XOR U1119 ( .A(B[665]), .B(A[665]), .Z(n746) );
  XOR U1120 ( .A(A[664]), .B(n747), .Z(O[664]) );
  AND U1121 ( .A(S), .B(n748), .Z(n747) );
  XOR U1122 ( .A(B[664]), .B(A[664]), .Z(n748) );
  XOR U1123 ( .A(A[663]), .B(n749), .Z(O[663]) );
  AND U1124 ( .A(S), .B(n750), .Z(n749) );
  XOR U1125 ( .A(B[663]), .B(A[663]), .Z(n750) );
  XOR U1126 ( .A(A[662]), .B(n751), .Z(O[662]) );
  AND U1127 ( .A(S), .B(n752), .Z(n751) );
  XOR U1128 ( .A(B[662]), .B(A[662]), .Z(n752) );
  XOR U1129 ( .A(A[661]), .B(n753), .Z(O[661]) );
  AND U1130 ( .A(S), .B(n754), .Z(n753) );
  XOR U1131 ( .A(B[661]), .B(A[661]), .Z(n754) );
  XOR U1132 ( .A(A[660]), .B(n755), .Z(O[660]) );
  AND U1133 ( .A(S), .B(n756), .Z(n755) );
  XOR U1134 ( .A(B[660]), .B(A[660]), .Z(n756) );
  XOR U1135 ( .A(A[65]), .B(n757), .Z(O[65]) );
  AND U1136 ( .A(S), .B(n758), .Z(n757) );
  XOR U1137 ( .A(B[65]), .B(A[65]), .Z(n758) );
  XOR U1138 ( .A(A[659]), .B(n759), .Z(O[659]) );
  AND U1139 ( .A(S), .B(n760), .Z(n759) );
  XOR U1140 ( .A(B[659]), .B(A[659]), .Z(n760) );
  XOR U1141 ( .A(A[658]), .B(n761), .Z(O[658]) );
  AND U1142 ( .A(S), .B(n762), .Z(n761) );
  XOR U1143 ( .A(B[658]), .B(A[658]), .Z(n762) );
  XOR U1144 ( .A(A[657]), .B(n763), .Z(O[657]) );
  AND U1145 ( .A(S), .B(n764), .Z(n763) );
  XOR U1146 ( .A(B[657]), .B(A[657]), .Z(n764) );
  XOR U1147 ( .A(A[656]), .B(n765), .Z(O[656]) );
  AND U1148 ( .A(S), .B(n766), .Z(n765) );
  XOR U1149 ( .A(B[656]), .B(A[656]), .Z(n766) );
  XOR U1150 ( .A(A[655]), .B(n767), .Z(O[655]) );
  AND U1151 ( .A(S), .B(n768), .Z(n767) );
  XOR U1152 ( .A(B[655]), .B(A[655]), .Z(n768) );
  XOR U1153 ( .A(A[654]), .B(n769), .Z(O[654]) );
  AND U1154 ( .A(S), .B(n770), .Z(n769) );
  XOR U1155 ( .A(B[654]), .B(A[654]), .Z(n770) );
  XOR U1156 ( .A(A[653]), .B(n771), .Z(O[653]) );
  AND U1157 ( .A(S), .B(n772), .Z(n771) );
  XOR U1158 ( .A(B[653]), .B(A[653]), .Z(n772) );
  XOR U1159 ( .A(A[652]), .B(n773), .Z(O[652]) );
  AND U1160 ( .A(S), .B(n774), .Z(n773) );
  XOR U1161 ( .A(B[652]), .B(A[652]), .Z(n774) );
  XOR U1162 ( .A(A[651]), .B(n775), .Z(O[651]) );
  AND U1163 ( .A(S), .B(n776), .Z(n775) );
  XOR U1164 ( .A(B[651]), .B(A[651]), .Z(n776) );
  XOR U1165 ( .A(A[650]), .B(n777), .Z(O[650]) );
  AND U1166 ( .A(S), .B(n778), .Z(n777) );
  XOR U1167 ( .A(B[650]), .B(A[650]), .Z(n778) );
  XOR U1168 ( .A(A[64]), .B(n779), .Z(O[64]) );
  AND U1169 ( .A(S), .B(n780), .Z(n779) );
  XOR U1170 ( .A(B[64]), .B(A[64]), .Z(n780) );
  XOR U1171 ( .A(A[649]), .B(n781), .Z(O[649]) );
  AND U1172 ( .A(S), .B(n782), .Z(n781) );
  XOR U1173 ( .A(B[649]), .B(A[649]), .Z(n782) );
  XOR U1174 ( .A(A[648]), .B(n783), .Z(O[648]) );
  AND U1175 ( .A(S), .B(n784), .Z(n783) );
  XOR U1176 ( .A(B[648]), .B(A[648]), .Z(n784) );
  XOR U1177 ( .A(A[647]), .B(n785), .Z(O[647]) );
  AND U1178 ( .A(S), .B(n786), .Z(n785) );
  XOR U1179 ( .A(B[647]), .B(A[647]), .Z(n786) );
  XOR U1180 ( .A(A[646]), .B(n787), .Z(O[646]) );
  AND U1181 ( .A(S), .B(n788), .Z(n787) );
  XOR U1182 ( .A(B[646]), .B(A[646]), .Z(n788) );
  XOR U1183 ( .A(A[645]), .B(n789), .Z(O[645]) );
  AND U1184 ( .A(S), .B(n790), .Z(n789) );
  XOR U1185 ( .A(B[645]), .B(A[645]), .Z(n790) );
  XOR U1186 ( .A(A[644]), .B(n791), .Z(O[644]) );
  AND U1187 ( .A(S), .B(n792), .Z(n791) );
  XOR U1188 ( .A(B[644]), .B(A[644]), .Z(n792) );
  XOR U1189 ( .A(A[643]), .B(n793), .Z(O[643]) );
  AND U1190 ( .A(S), .B(n794), .Z(n793) );
  XOR U1191 ( .A(B[643]), .B(A[643]), .Z(n794) );
  XOR U1192 ( .A(A[642]), .B(n795), .Z(O[642]) );
  AND U1193 ( .A(S), .B(n796), .Z(n795) );
  XOR U1194 ( .A(B[642]), .B(A[642]), .Z(n796) );
  XOR U1195 ( .A(A[641]), .B(n797), .Z(O[641]) );
  AND U1196 ( .A(S), .B(n798), .Z(n797) );
  XOR U1197 ( .A(B[641]), .B(A[641]), .Z(n798) );
  XOR U1198 ( .A(A[640]), .B(n799), .Z(O[640]) );
  AND U1199 ( .A(S), .B(n800), .Z(n799) );
  XOR U1200 ( .A(B[640]), .B(A[640]), .Z(n800) );
  XOR U1201 ( .A(A[63]), .B(n801), .Z(O[63]) );
  AND U1202 ( .A(S), .B(n802), .Z(n801) );
  XOR U1203 ( .A(B[63]), .B(A[63]), .Z(n802) );
  XOR U1204 ( .A(A[639]), .B(n803), .Z(O[639]) );
  AND U1205 ( .A(S), .B(n804), .Z(n803) );
  XOR U1206 ( .A(B[639]), .B(A[639]), .Z(n804) );
  XOR U1207 ( .A(A[638]), .B(n805), .Z(O[638]) );
  AND U1208 ( .A(S), .B(n806), .Z(n805) );
  XOR U1209 ( .A(B[638]), .B(A[638]), .Z(n806) );
  XOR U1210 ( .A(A[637]), .B(n807), .Z(O[637]) );
  AND U1211 ( .A(S), .B(n808), .Z(n807) );
  XOR U1212 ( .A(B[637]), .B(A[637]), .Z(n808) );
  XOR U1213 ( .A(A[636]), .B(n809), .Z(O[636]) );
  AND U1214 ( .A(S), .B(n810), .Z(n809) );
  XOR U1215 ( .A(B[636]), .B(A[636]), .Z(n810) );
  XOR U1216 ( .A(A[635]), .B(n811), .Z(O[635]) );
  AND U1217 ( .A(S), .B(n812), .Z(n811) );
  XOR U1218 ( .A(B[635]), .B(A[635]), .Z(n812) );
  XOR U1219 ( .A(A[634]), .B(n813), .Z(O[634]) );
  AND U1220 ( .A(S), .B(n814), .Z(n813) );
  XOR U1221 ( .A(B[634]), .B(A[634]), .Z(n814) );
  XOR U1222 ( .A(A[633]), .B(n815), .Z(O[633]) );
  AND U1223 ( .A(S), .B(n816), .Z(n815) );
  XOR U1224 ( .A(B[633]), .B(A[633]), .Z(n816) );
  XOR U1225 ( .A(A[632]), .B(n817), .Z(O[632]) );
  AND U1226 ( .A(S), .B(n818), .Z(n817) );
  XOR U1227 ( .A(B[632]), .B(A[632]), .Z(n818) );
  XOR U1228 ( .A(A[631]), .B(n819), .Z(O[631]) );
  AND U1229 ( .A(S), .B(n820), .Z(n819) );
  XOR U1230 ( .A(B[631]), .B(A[631]), .Z(n820) );
  XOR U1231 ( .A(A[630]), .B(n821), .Z(O[630]) );
  AND U1232 ( .A(S), .B(n822), .Z(n821) );
  XOR U1233 ( .A(B[630]), .B(A[630]), .Z(n822) );
  XOR U1234 ( .A(A[62]), .B(n823), .Z(O[62]) );
  AND U1235 ( .A(S), .B(n824), .Z(n823) );
  XOR U1236 ( .A(B[62]), .B(A[62]), .Z(n824) );
  XOR U1237 ( .A(A[629]), .B(n825), .Z(O[629]) );
  AND U1238 ( .A(S), .B(n826), .Z(n825) );
  XOR U1239 ( .A(B[629]), .B(A[629]), .Z(n826) );
  XOR U1240 ( .A(A[628]), .B(n827), .Z(O[628]) );
  AND U1241 ( .A(S), .B(n828), .Z(n827) );
  XOR U1242 ( .A(B[628]), .B(A[628]), .Z(n828) );
  XOR U1243 ( .A(A[627]), .B(n829), .Z(O[627]) );
  AND U1244 ( .A(S), .B(n830), .Z(n829) );
  XOR U1245 ( .A(B[627]), .B(A[627]), .Z(n830) );
  XOR U1246 ( .A(A[626]), .B(n831), .Z(O[626]) );
  AND U1247 ( .A(S), .B(n832), .Z(n831) );
  XOR U1248 ( .A(B[626]), .B(A[626]), .Z(n832) );
  XOR U1249 ( .A(A[625]), .B(n833), .Z(O[625]) );
  AND U1250 ( .A(S), .B(n834), .Z(n833) );
  XOR U1251 ( .A(B[625]), .B(A[625]), .Z(n834) );
  XOR U1252 ( .A(A[624]), .B(n835), .Z(O[624]) );
  AND U1253 ( .A(S), .B(n836), .Z(n835) );
  XOR U1254 ( .A(B[624]), .B(A[624]), .Z(n836) );
  XOR U1255 ( .A(A[623]), .B(n837), .Z(O[623]) );
  AND U1256 ( .A(S), .B(n838), .Z(n837) );
  XOR U1257 ( .A(B[623]), .B(A[623]), .Z(n838) );
  XOR U1258 ( .A(A[622]), .B(n839), .Z(O[622]) );
  AND U1259 ( .A(S), .B(n840), .Z(n839) );
  XOR U1260 ( .A(B[622]), .B(A[622]), .Z(n840) );
  XOR U1261 ( .A(A[621]), .B(n841), .Z(O[621]) );
  AND U1262 ( .A(S), .B(n842), .Z(n841) );
  XOR U1263 ( .A(B[621]), .B(A[621]), .Z(n842) );
  XOR U1264 ( .A(A[620]), .B(n843), .Z(O[620]) );
  AND U1265 ( .A(S), .B(n844), .Z(n843) );
  XOR U1266 ( .A(B[620]), .B(A[620]), .Z(n844) );
  XOR U1267 ( .A(A[61]), .B(n845), .Z(O[61]) );
  AND U1268 ( .A(S), .B(n846), .Z(n845) );
  XOR U1269 ( .A(B[61]), .B(A[61]), .Z(n846) );
  XOR U1270 ( .A(A[619]), .B(n847), .Z(O[619]) );
  AND U1271 ( .A(S), .B(n848), .Z(n847) );
  XOR U1272 ( .A(B[619]), .B(A[619]), .Z(n848) );
  XOR U1273 ( .A(A[618]), .B(n849), .Z(O[618]) );
  AND U1274 ( .A(S), .B(n850), .Z(n849) );
  XOR U1275 ( .A(B[618]), .B(A[618]), .Z(n850) );
  XOR U1276 ( .A(A[617]), .B(n851), .Z(O[617]) );
  AND U1277 ( .A(S), .B(n852), .Z(n851) );
  XOR U1278 ( .A(B[617]), .B(A[617]), .Z(n852) );
  XOR U1279 ( .A(A[616]), .B(n853), .Z(O[616]) );
  AND U1280 ( .A(S), .B(n854), .Z(n853) );
  XOR U1281 ( .A(B[616]), .B(A[616]), .Z(n854) );
  XOR U1282 ( .A(A[615]), .B(n855), .Z(O[615]) );
  AND U1283 ( .A(S), .B(n856), .Z(n855) );
  XOR U1284 ( .A(B[615]), .B(A[615]), .Z(n856) );
  XOR U1285 ( .A(A[614]), .B(n857), .Z(O[614]) );
  AND U1286 ( .A(S), .B(n858), .Z(n857) );
  XOR U1287 ( .A(B[614]), .B(A[614]), .Z(n858) );
  XOR U1288 ( .A(A[613]), .B(n859), .Z(O[613]) );
  AND U1289 ( .A(S), .B(n860), .Z(n859) );
  XOR U1290 ( .A(B[613]), .B(A[613]), .Z(n860) );
  XOR U1291 ( .A(A[612]), .B(n861), .Z(O[612]) );
  AND U1292 ( .A(S), .B(n862), .Z(n861) );
  XOR U1293 ( .A(B[612]), .B(A[612]), .Z(n862) );
  XOR U1294 ( .A(A[611]), .B(n863), .Z(O[611]) );
  AND U1295 ( .A(S), .B(n864), .Z(n863) );
  XOR U1296 ( .A(B[611]), .B(A[611]), .Z(n864) );
  XOR U1297 ( .A(A[610]), .B(n865), .Z(O[610]) );
  AND U1298 ( .A(S), .B(n866), .Z(n865) );
  XOR U1299 ( .A(B[610]), .B(A[610]), .Z(n866) );
  XOR U1300 ( .A(A[60]), .B(n867), .Z(O[60]) );
  AND U1301 ( .A(S), .B(n868), .Z(n867) );
  XOR U1302 ( .A(B[60]), .B(A[60]), .Z(n868) );
  XOR U1303 ( .A(A[609]), .B(n869), .Z(O[609]) );
  AND U1304 ( .A(S), .B(n870), .Z(n869) );
  XOR U1305 ( .A(B[609]), .B(A[609]), .Z(n870) );
  XOR U1306 ( .A(A[608]), .B(n871), .Z(O[608]) );
  AND U1307 ( .A(S), .B(n872), .Z(n871) );
  XOR U1308 ( .A(B[608]), .B(A[608]), .Z(n872) );
  XOR U1309 ( .A(A[607]), .B(n873), .Z(O[607]) );
  AND U1310 ( .A(S), .B(n874), .Z(n873) );
  XOR U1311 ( .A(B[607]), .B(A[607]), .Z(n874) );
  XOR U1312 ( .A(A[606]), .B(n875), .Z(O[606]) );
  AND U1313 ( .A(S), .B(n876), .Z(n875) );
  XOR U1314 ( .A(B[606]), .B(A[606]), .Z(n876) );
  XOR U1315 ( .A(A[605]), .B(n877), .Z(O[605]) );
  AND U1316 ( .A(S), .B(n878), .Z(n877) );
  XOR U1317 ( .A(B[605]), .B(A[605]), .Z(n878) );
  XOR U1318 ( .A(A[604]), .B(n879), .Z(O[604]) );
  AND U1319 ( .A(S), .B(n880), .Z(n879) );
  XOR U1320 ( .A(B[604]), .B(A[604]), .Z(n880) );
  XOR U1321 ( .A(A[603]), .B(n881), .Z(O[603]) );
  AND U1322 ( .A(S), .B(n882), .Z(n881) );
  XOR U1323 ( .A(B[603]), .B(A[603]), .Z(n882) );
  XOR U1324 ( .A(A[602]), .B(n883), .Z(O[602]) );
  AND U1325 ( .A(S), .B(n884), .Z(n883) );
  XOR U1326 ( .A(B[602]), .B(A[602]), .Z(n884) );
  XOR U1327 ( .A(A[601]), .B(n885), .Z(O[601]) );
  AND U1328 ( .A(S), .B(n886), .Z(n885) );
  XOR U1329 ( .A(B[601]), .B(A[601]), .Z(n886) );
  XOR U1330 ( .A(A[600]), .B(n887), .Z(O[600]) );
  AND U1331 ( .A(S), .B(n888), .Z(n887) );
  XOR U1332 ( .A(B[600]), .B(A[600]), .Z(n888) );
  XOR U1333 ( .A(A[5]), .B(n889), .Z(O[5]) );
  AND U1334 ( .A(S), .B(n890), .Z(n889) );
  XOR U1335 ( .A(B[5]), .B(A[5]), .Z(n890) );
  XOR U1336 ( .A(A[59]), .B(n891), .Z(O[59]) );
  AND U1337 ( .A(S), .B(n892), .Z(n891) );
  XOR U1338 ( .A(B[59]), .B(A[59]), .Z(n892) );
  XOR U1339 ( .A(A[599]), .B(n893), .Z(O[599]) );
  AND U1340 ( .A(S), .B(n894), .Z(n893) );
  XOR U1341 ( .A(B[599]), .B(A[599]), .Z(n894) );
  XOR U1342 ( .A(A[598]), .B(n895), .Z(O[598]) );
  AND U1343 ( .A(S), .B(n896), .Z(n895) );
  XOR U1344 ( .A(B[598]), .B(A[598]), .Z(n896) );
  XOR U1345 ( .A(A[597]), .B(n897), .Z(O[597]) );
  AND U1346 ( .A(S), .B(n898), .Z(n897) );
  XOR U1347 ( .A(B[597]), .B(A[597]), .Z(n898) );
  XOR U1348 ( .A(A[596]), .B(n899), .Z(O[596]) );
  AND U1349 ( .A(S), .B(n900), .Z(n899) );
  XOR U1350 ( .A(B[596]), .B(A[596]), .Z(n900) );
  XOR U1351 ( .A(A[595]), .B(n901), .Z(O[595]) );
  AND U1352 ( .A(S), .B(n902), .Z(n901) );
  XOR U1353 ( .A(B[595]), .B(A[595]), .Z(n902) );
  XOR U1354 ( .A(A[594]), .B(n903), .Z(O[594]) );
  AND U1355 ( .A(S), .B(n904), .Z(n903) );
  XOR U1356 ( .A(B[594]), .B(A[594]), .Z(n904) );
  XOR U1357 ( .A(A[593]), .B(n905), .Z(O[593]) );
  AND U1358 ( .A(S), .B(n906), .Z(n905) );
  XOR U1359 ( .A(B[593]), .B(A[593]), .Z(n906) );
  XOR U1360 ( .A(A[592]), .B(n907), .Z(O[592]) );
  AND U1361 ( .A(S), .B(n908), .Z(n907) );
  XOR U1362 ( .A(B[592]), .B(A[592]), .Z(n908) );
  XOR U1363 ( .A(A[591]), .B(n909), .Z(O[591]) );
  AND U1364 ( .A(S), .B(n910), .Z(n909) );
  XOR U1365 ( .A(B[591]), .B(A[591]), .Z(n910) );
  XOR U1366 ( .A(A[590]), .B(n911), .Z(O[590]) );
  AND U1367 ( .A(S), .B(n912), .Z(n911) );
  XOR U1368 ( .A(B[590]), .B(A[590]), .Z(n912) );
  XOR U1369 ( .A(A[58]), .B(n913), .Z(O[58]) );
  AND U1370 ( .A(S), .B(n914), .Z(n913) );
  XOR U1371 ( .A(B[58]), .B(A[58]), .Z(n914) );
  XOR U1372 ( .A(A[589]), .B(n915), .Z(O[589]) );
  AND U1373 ( .A(S), .B(n916), .Z(n915) );
  XOR U1374 ( .A(B[589]), .B(A[589]), .Z(n916) );
  XOR U1375 ( .A(A[588]), .B(n917), .Z(O[588]) );
  AND U1376 ( .A(S), .B(n918), .Z(n917) );
  XOR U1377 ( .A(B[588]), .B(A[588]), .Z(n918) );
  XOR U1378 ( .A(A[587]), .B(n919), .Z(O[587]) );
  AND U1379 ( .A(S), .B(n920), .Z(n919) );
  XOR U1380 ( .A(B[587]), .B(A[587]), .Z(n920) );
  XOR U1381 ( .A(A[586]), .B(n921), .Z(O[586]) );
  AND U1382 ( .A(S), .B(n922), .Z(n921) );
  XOR U1383 ( .A(B[586]), .B(A[586]), .Z(n922) );
  XOR U1384 ( .A(A[585]), .B(n923), .Z(O[585]) );
  AND U1385 ( .A(S), .B(n924), .Z(n923) );
  XOR U1386 ( .A(B[585]), .B(A[585]), .Z(n924) );
  XOR U1387 ( .A(A[584]), .B(n925), .Z(O[584]) );
  AND U1388 ( .A(S), .B(n926), .Z(n925) );
  XOR U1389 ( .A(B[584]), .B(A[584]), .Z(n926) );
  XOR U1390 ( .A(A[583]), .B(n927), .Z(O[583]) );
  AND U1391 ( .A(S), .B(n928), .Z(n927) );
  XOR U1392 ( .A(B[583]), .B(A[583]), .Z(n928) );
  XOR U1393 ( .A(A[582]), .B(n929), .Z(O[582]) );
  AND U1394 ( .A(S), .B(n930), .Z(n929) );
  XOR U1395 ( .A(B[582]), .B(A[582]), .Z(n930) );
  XOR U1396 ( .A(A[581]), .B(n931), .Z(O[581]) );
  AND U1397 ( .A(S), .B(n932), .Z(n931) );
  XOR U1398 ( .A(B[581]), .B(A[581]), .Z(n932) );
  XOR U1399 ( .A(A[580]), .B(n933), .Z(O[580]) );
  AND U1400 ( .A(S), .B(n934), .Z(n933) );
  XOR U1401 ( .A(B[580]), .B(A[580]), .Z(n934) );
  XOR U1402 ( .A(A[57]), .B(n935), .Z(O[57]) );
  AND U1403 ( .A(S), .B(n936), .Z(n935) );
  XOR U1404 ( .A(B[57]), .B(A[57]), .Z(n936) );
  XOR U1405 ( .A(A[579]), .B(n937), .Z(O[579]) );
  AND U1406 ( .A(S), .B(n938), .Z(n937) );
  XOR U1407 ( .A(B[579]), .B(A[579]), .Z(n938) );
  XOR U1408 ( .A(A[578]), .B(n939), .Z(O[578]) );
  AND U1409 ( .A(S), .B(n940), .Z(n939) );
  XOR U1410 ( .A(B[578]), .B(A[578]), .Z(n940) );
  XOR U1411 ( .A(A[577]), .B(n941), .Z(O[577]) );
  AND U1412 ( .A(S), .B(n942), .Z(n941) );
  XOR U1413 ( .A(B[577]), .B(A[577]), .Z(n942) );
  XOR U1414 ( .A(A[576]), .B(n943), .Z(O[576]) );
  AND U1415 ( .A(S), .B(n944), .Z(n943) );
  XOR U1416 ( .A(B[576]), .B(A[576]), .Z(n944) );
  XOR U1417 ( .A(A[575]), .B(n945), .Z(O[575]) );
  AND U1418 ( .A(S), .B(n946), .Z(n945) );
  XOR U1419 ( .A(B[575]), .B(A[575]), .Z(n946) );
  XOR U1420 ( .A(A[574]), .B(n947), .Z(O[574]) );
  AND U1421 ( .A(S), .B(n948), .Z(n947) );
  XOR U1422 ( .A(B[574]), .B(A[574]), .Z(n948) );
  XOR U1423 ( .A(A[573]), .B(n949), .Z(O[573]) );
  AND U1424 ( .A(S), .B(n950), .Z(n949) );
  XOR U1425 ( .A(B[573]), .B(A[573]), .Z(n950) );
  XOR U1426 ( .A(A[572]), .B(n951), .Z(O[572]) );
  AND U1427 ( .A(S), .B(n952), .Z(n951) );
  XOR U1428 ( .A(B[572]), .B(A[572]), .Z(n952) );
  XOR U1429 ( .A(A[571]), .B(n953), .Z(O[571]) );
  AND U1430 ( .A(S), .B(n954), .Z(n953) );
  XOR U1431 ( .A(B[571]), .B(A[571]), .Z(n954) );
  XOR U1432 ( .A(A[570]), .B(n955), .Z(O[570]) );
  AND U1433 ( .A(S), .B(n956), .Z(n955) );
  XOR U1434 ( .A(B[570]), .B(A[570]), .Z(n956) );
  XOR U1435 ( .A(A[56]), .B(n957), .Z(O[56]) );
  AND U1436 ( .A(S), .B(n958), .Z(n957) );
  XOR U1437 ( .A(B[56]), .B(A[56]), .Z(n958) );
  XOR U1438 ( .A(A[569]), .B(n959), .Z(O[569]) );
  AND U1439 ( .A(S), .B(n960), .Z(n959) );
  XOR U1440 ( .A(B[569]), .B(A[569]), .Z(n960) );
  XOR U1441 ( .A(A[568]), .B(n961), .Z(O[568]) );
  AND U1442 ( .A(S), .B(n962), .Z(n961) );
  XOR U1443 ( .A(B[568]), .B(A[568]), .Z(n962) );
  XOR U1444 ( .A(A[567]), .B(n963), .Z(O[567]) );
  AND U1445 ( .A(S), .B(n964), .Z(n963) );
  XOR U1446 ( .A(B[567]), .B(A[567]), .Z(n964) );
  XOR U1447 ( .A(A[566]), .B(n965), .Z(O[566]) );
  AND U1448 ( .A(S), .B(n966), .Z(n965) );
  XOR U1449 ( .A(B[566]), .B(A[566]), .Z(n966) );
  XOR U1450 ( .A(A[565]), .B(n967), .Z(O[565]) );
  AND U1451 ( .A(S), .B(n968), .Z(n967) );
  XOR U1452 ( .A(B[565]), .B(A[565]), .Z(n968) );
  XOR U1453 ( .A(A[564]), .B(n969), .Z(O[564]) );
  AND U1454 ( .A(S), .B(n970), .Z(n969) );
  XOR U1455 ( .A(B[564]), .B(A[564]), .Z(n970) );
  XOR U1456 ( .A(A[563]), .B(n971), .Z(O[563]) );
  AND U1457 ( .A(S), .B(n972), .Z(n971) );
  XOR U1458 ( .A(B[563]), .B(A[563]), .Z(n972) );
  XOR U1459 ( .A(A[562]), .B(n973), .Z(O[562]) );
  AND U1460 ( .A(S), .B(n974), .Z(n973) );
  XOR U1461 ( .A(B[562]), .B(A[562]), .Z(n974) );
  XOR U1462 ( .A(A[561]), .B(n975), .Z(O[561]) );
  AND U1463 ( .A(S), .B(n976), .Z(n975) );
  XOR U1464 ( .A(B[561]), .B(A[561]), .Z(n976) );
  XOR U1465 ( .A(A[560]), .B(n977), .Z(O[560]) );
  AND U1466 ( .A(S), .B(n978), .Z(n977) );
  XOR U1467 ( .A(B[560]), .B(A[560]), .Z(n978) );
  XOR U1468 ( .A(A[55]), .B(n979), .Z(O[55]) );
  AND U1469 ( .A(S), .B(n980), .Z(n979) );
  XOR U1470 ( .A(B[55]), .B(A[55]), .Z(n980) );
  XOR U1471 ( .A(A[559]), .B(n981), .Z(O[559]) );
  AND U1472 ( .A(S), .B(n982), .Z(n981) );
  XOR U1473 ( .A(B[559]), .B(A[559]), .Z(n982) );
  XOR U1474 ( .A(A[558]), .B(n983), .Z(O[558]) );
  AND U1475 ( .A(S), .B(n984), .Z(n983) );
  XOR U1476 ( .A(B[558]), .B(A[558]), .Z(n984) );
  XOR U1477 ( .A(A[557]), .B(n985), .Z(O[557]) );
  AND U1478 ( .A(S), .B(n986), .Z(n985) );
  XOR U1479 ( .A(B[557]), .B(A[557]), .Z(n986) );
  XOR U1480 ( .A(A[556]), .B(n987), .Z(O[556]) );
  AND U1481 ( .A(S), .B(n988), .Z(n987) );
  XOR U1482 ( .A(B[556]), .B(A[556]), .Z(n988) );
  XOR U1483 ( .A(A[555]), .B(n989), .Z(O[555]) );
  AND U1484 ( .A(S), .B(n990), .Z(n989) );
  XOR U1485 ( .A(B[555]), .B(A[555]), .Z(n990) );
  XOR U1486 ( .A(A[554]), .B(n991), .Z(O[554]) );
  AND U1487 ( .A(S), .B(n992), .Z(n991) );
  XOR U1488 ( .A(B[554]), .B(A[554]), .Z(n992) );
  XOR U1489 ( .A(A[553]), .B(n993), .Z(O[553]) );
  AND U1490 ( .A(S), .B(n994), .Z(n993) );
  XOR U1491 ( .A(B[553]), .B(A[553]), .Z(n994) );
  XOR U1492 ( .A(A[552]), .B(n995), .Z(O[552]) );
  AND U1493 ( .A(S), .B(n996), .Z(n995) );
  XOR U1494 ( .A(B[552]), .B(A[552]), .Z(n996) );
  XOR U1495 ( .A(A[551]), .B(n997), .Z(O[551]) );
  AND U1496 ( .A(S), .B(n998), .Z(n997) );
  XOR U1497 ( .A(B[551]), .B(A[551]), .Z(n998) );
  XOR U1498 ( .A(A[550]), .B(n999), .Z(O[550]) );
  AND U1499 ( .A(S), .B(n1000), .Z(n999) );
  XOR U1500 ( .A(B[550]), .B(A[550]), .Z(n1000) );
  XOR U1501 ( .A(A[54]), .B(n1001), .Z(O[54]) );
  AND U1502 ( .A(S), .B(n1002), .Z(n1001) );
  XOR U1503 ( .A(B[54]), .B(A[54]), .Z(n1002) );
  XOR U1504 ( .A(A[549]), .B(n1003), .Z(O[549]) );
  AND U1505 ( .A(S), .B(n1004), .Z(n1003) );
  XOR U1506 ( .A(B[549]), .B(A[549]), .Z(n1004) );
  XOR U1507 ( .A(A[548]), .B(n1005), .Z(O[548]) );
  AND U1508 ( .A(S), .B(n1006), .Z(n1005) );
  XOR U1509 ( .A(B[548]), .B(A[548]), .Z(n1006) );
  XOR U1510 ( .A(A[547]), .B(n1007), .Z(O[547]) );
  AND U1511 ( .A(S), .B(n1008), .Z(n1007) );
  XOR U1512 ( .A(B[547]), .B(A[547]), .Z(n1008) );
  XOR U1513 ( .A(A[546]), .B(n1009), .Z(O[546]) );
  AND U1514 ( .A(S), .B(n1010), .Z(n1009) );
  XOR U1515 ( .A(B[546]), .B(A[546]), .Z(n1010) );
  XOR U1516 ( .A(A[545]), .B(n1011), .Z(O[545]) );
  AND U1517 ( .A(S), .B(n1012), .Z(n1011) );
  XOR U1518 ( .A(B[545]), .B(A[545]), .Z(n1012) );
  XOR U1519 ( .A(A[544]), .B(n1013), .Z(O[544]) );
  AND U1520 ( .A(S), .B(n1014), .Z(n1013) );
  XOR U1521 ( .A(B[544]), .B(A[544]), .Z(n1014) );
  XOR U1522 ( .A(A[543]), .B(n1015), .Z(O[543]) );
  AND U1523 ( .A(S), .B(n1016), .Z(n1015) );
  XOR U1524 ( .A(B[543]), .B(A[543]), .Z(n1016) );
  XOR U1525 ( .A(A[542]), .B(n1017), .Z(O[542]) );
  AND U1526 ( .A(S), .B(n1018), .Z(n1017) );
  XOR U1527 ( .A(B[542]), .B(A[542]), .Z(n1018) );
  XOR U1528 ( .A(A[541]), .B(n1019), .Z(O[541]) );
  AND U1529 ( .A(S), .B(n1020), .Z(n1019) );
  XOR U1530 ( .A(B[541]), .B(A[541]), .Z(n1020) );
  XOR U1531 ( .A(A[540]), .B(n1021), .Z(O[540]) );
  AND U1532 ( .A(S), .B(n1022), .Z(n1021) );
  XOR U1533 ( .A(B[540]), .B(A[540]), .Z(n1022) );
  XOR U1534 ( .A(A[53]), .B(n1023), .Z(O[53]) );
  AND U1535 ( .A(S), .B(n1024), .Z(n1023) );
  XOR U1536 ( .A(B[53]), .B(A[53]), .Z(n1024) );
  XOR U1537 ( .A(A[539]), .B(n1025), .Z(O[539]) );
  AND U1538 ( .A(S), .B(n1026), .Z(n1025) );
  XOR U1539 ( .A(B[539]), .B(A[539]), .Z(n1026) );
  XOR U1540 ( .A(A[538]), .B(n1027), .Z(O[538]) );
  AND U1541 ( .A(S), .B(n1028), .Z(n1027) );
  XOR U1542 ( .A(B[538]), .B(A[538]), .Z(n1028) );
  XOR U1543 ( .A(A[537]), .B(n1029), .Z(O[537]) );
  AND U1544 ( .A(S), .B(n1030), .Z(n1029) );
  XOR U1545 ( .A(B[537]), .B(A[537]), .Z(n1030) );
  XOR U1546 ( .A(A[536]), .B(n1031), .Z(O[536]) );
  AND U1547 ( .A(S), .B(n1032), .Z(n1031) );
  XOR U1548 ( .A(B[536]), .B(A[536]), .Z(n1032) );
  XOR U1549 ( .A(A[535]), .B(n1033), .Z(O[535]) );
  AND U1550 ( .A(S), .B(n1034), .Z(n1033) );
  XOR U1551 ( .A(B[535]), .B(A[535]), .Z(n1034) );
  XOR U1552 ( .A(A[534]), .B(n1035), .Z(O[534]) );
  AND U1553 ( .A(S), .B(n1036), .Z(n1035) );
  XOR U1554 ( .A(B[534]), .B(A[534]), .Z(n1036) );
  XOR U1555 ( .A(A[533]), .B(n1037), .Z(O[533]) );
  AND U1556 ( .A(S), .B(n1038), .Z(n1037) );
  XOR U1557 ( .A(B[533]), .B(A[533]), .Z(n1038) );
  XOR U1558 ( .A(A[532]), .B(n1039), .Z(O[532]) );
  AND U1559 ( .A(S), .B(n1040), .Z(n1039) );
  XOR U1560 ( .A(B[532]), .B(A[532]), .Z(n1040) );
  XOR U1561 ( .A(A[531]), .B(n1041), .Z(O[531]) );
  AND U1562 ( .A(S), .B(n1042), .Z(n1041) );
  XOR U1563 ( .A(B[531]), .B(A[531]), .Z(n1042) );
  XOR U1564 ( .A(A[530]), .B(n1043), .Z(O[530]) );
  AND U1565 ( .A(S), .B(n1044), .Z(n1043) );
  XOR U1566 ( .A(B[530]), .B(A[530]), .Z(n1044) );
  XOR U1567 ( .A(A[52]), .B(n1045), .Z(O[52]) );
  AND U1568 ( .A(S), .B(n1046), .Z(n1045) );
  XOR U1569 ( .A(B[52]), .B(A[52]), .Z(n1046) );
  XOR U1570 ( .A(A[529]), .B(n1047), .Z(O[529]) );
  AND U1571 ( .A(S), .B(n1048), .Z(n1047) );
  XOR U1572 ( .A(B[529]), .B(A[529]), .Z(n1048) );
  XOR U1573 ( .A(A[528]), .B(n1049), .Z(O[528]) );
  AND U1574 ( .A(S), .B(n1050), .Z(n1049) );
  XOR U1575 ( .A(B[528]), .B(A[528]), .Z(n1050) );
  XOR U1576 ( .A(A[527]), .B(n1051), .Z(O[527]) );
  AND U1577 ( .A(S), .B(n1052), .Z(n1051) );
  XOR U1578 ( .A(B[527]), .B(A[527]), .Z(n1052) );
  XOR U1579 ( .A(A[526]), .B(n1053), .Z(O[526]) );
  AND U1580 ( .A(S), .B(n1054), .Z(n1053) );
  XOR U1581 ( .A(B[526]), .B(A[526]), .Z(n1054) );
  XOR U1582 ( .A(A[525]), .B(n1055), .Z(O[525]) );
  AND U1583 ( .A(S), .B(n1056), .Z(n1055) );
  XOR U1584 ( .A(B[525]), .B(A[525]), .Z(n1056) );
  XOR U1585 ( .A(A[524]), .B(n1057), .Z(O[524]) );
  AND U1586 ( .A(S), .B(n1058), .Z(n1057) );
  XOR U1587 ( .A(B[524]), .B(A[524]), .Z(n1058) );
  XOR U1588 ( .A(A[523]), .B(n1059), .Z(O[523]) );
  AND U1589 ( .A(S), .B(n1060), .Z(n1059) );
  XOR U1590 ( .A(B[523]), .B(A[523]), .Z(n1060) );
  XOR U1591 ( .A(A[522]), .B(n1061), .Z(O[522]) );
  AND U1592 ( .A(S), .B(n1062), .Z(n1061) );
  XOR U1593 ( .A(B[522]), .B(A[522]), .Z(n1062) );
  XOR U1594 ( .A(A[521]), .B(n1063), .Z(O[521]) );
  AND U1595 ( .A(S), .B(n1064), .Z(n1063) );
  XOR U1596 ( .A(B[521]), .B(A[521]), .Z(n1064) );
  XOR U1597 ( .A(A[520]), .B(n1065), .Z(O[520]) );
  AND U1598 ( .A(S), .B(n1066), .Z(n1065) );
  XOR U1599 ( .A(B[520]), .B(A[520]), .Z(n1066) );
  XOR U1600 ( .A(A[51]), .B(n1067), .Z(O[51]) );
  AND U1601 ( .A(S), .B(n1068), .Z(n1067) );
  XOR U1602 ( .A(B[51]), .B(A[51]), .Z(n1068) );
  XOR U1603 ( .A(A[519]), .B(n1069), .Z(O[519]) );
  AND U1604 ( .A(S), .B(n1070), .Z(n1069) );
  XOR U1605 ( .A(B[519]), .B(A[519]), .Z(n1070) );
  XOR U1606 ( .A(A[518]), .B(n1071), .Z(O[518]) );
  AND U1607 ( .A(S), .B(n1072), .Z(n1071) );
  XOR U1608 ( .A(B[518]), .B(A[518]), .Z(n1072) );
  XOR U1609 ( .A(A[517]), .B(n1073), .Z(O[517]) );
  AND U1610 ( .A(S), .B(n1074), .Z(n1073) );
  XOR U1611 ( .A(B[517]), .B(A[517]), .Z(n1074) );
  XOR U1612 ( .A(A[516]), .B(n1075), .Z(O[516]) );
  AND U1613 ( .A(S), .B(n1076), .Z(n1075) );
  XOR U1614 ( .A(B[516]), .B(A[516]), .Z(n1076) );
  XOR U1615 ( .A(A[515]), .B(n1077), .Z(O[515]) );
  AND U1616 ( .A(S), .B(n1078), .Z(n1077) );
  XOR U1617 ( .A(B[515]), .B(A[515]), .Z(n1078) );
  XOR U1618 ( .A(A[514]), .B(n1079), .Z(O[514]) );
  AND U1619 ( .A(S), .B(n1080), .Z(n1079) );
  XOR U1620 ( .A(B[514]), .B(A[514]), .Z(n1080) );
  XOR U1621 ( .A(A[513]), .B(n1081), .Z(O[513]) );
  AND U1622 ( .A(S), .B(n1082), .Z(n1081) );
  XOR U1623 ( .A(B[513]), .B(A[513]), .Z(n1082) );
  XOR U1624 ( .A(A[512]), .B(n1083), .Z(O[512]) );
  AND U1625 ( .A(S), .B(n1084), .Z(n1083) );
  XOR U1626 ( .A(B[512]), .B(A[512]), .Z(n1084) );
  XOR U1627 ( .A(A[511]), .B(n1085), .Z(O[511]) );
  AND U1628 ( .A(S), .B(n1086), .Z(n1085) );
  XOR U1629 ( .A(B[511]), .B(A[511]), .Z(n1086) );
  XOR U1630 ( .A(A[510]), .B(n1087), .Z(O[510]) );
  AND U1631 ( .A(S), .B(n1088), .Z(n1087) );
  XOR U1632 ( .A(B[510]), .B(A[510]), .Z(n1088) );
  XOR U1633 ( .A(A[50]), .B(n1089), .Z(O[50]) );
  AND U1634 ( .A(S), .B(n1090), .Z(n1089) );
  XOR U1635 ( .A(B[50]), .B(A[50]), .Z(n1090) );
  XOR U1636 ( .A(A[509]), .B(n1091), .Z(O[509]) );
  AND U1637 ( .A(S), .B(n1092), .Z(n1091) );
  XOR U1638 ( .A(B[509]), .B(A[509]), .Z(n1092) );
  XOR U1639 ( .A(A[508]), .B(n1093), .Z(O[508]) );
  AND U1640 ( .A(S), .B(n1094), .Z(n1093) );
  XOR U1641 ( .A(B[508]), .B(A[508]), .Z(n1094) );
  XOR U1642 ( .A(A[507]), .B(n1095), .Z(O[507]) );
  AND U1643 ( .A(S), .B(n1096), .Z(n1095) );
  XOR U1644 ( .A(B[507]), .B(A[507]), .Z(n1096) );
  XOR U1645 ( .A(A[506]), .B(n1097), .Z(O[506]) );
  AND U1646 ( .A(S), .B(n1098), .Z(n1097) );
  XOR U1647 ( .A(B[506]), .B(A[506]), .Z(n1098) );
  XOR U1648 ( .A(A[505]), .B(n1099), .Z(O[505]) );
  AND U1649 ( .A(S), .B(n1100), .Z(n1099) );
  XOR U1650 ( .A(B[505]), .B(A[505]), .Z(n1100) );
  XOR U1651 ( .A(A[504]), .B(n1101), .Z(O[504]) );
  AND U1652 ( .A(S), .B(n1102), .Z(n1101) );
  XOR U1653 ( .A(B[504]), .B(A[504]), .Z(n1102) );
  XOR U1654 ( .A(A[503]), .B(n1103), .Z(O[503]) );
  AND U1655 ( .A(S), .B(n1104), .Z(n1103) );
  XOR U1656 ( .A(B[503]), .B(A[503]), .Z(n1104) );
  XOR U1657 ( .A(A[502]), .B(n1105), .Z(O[502]) );
  AND U1658 ( .A(S), .B(n1106), .Z(n1105) );
  XOR U1659 ( .A(B[502]), .B(A[502]), .Z(n1106) );
  XOR U1660 ( .A(A[501]), .B(n1107), .Z(O[501]) );
  AND U1661 ( .A(S), .B(n1108), .Z(n1107) );
  XOR U1662 ( .A(B[501]), .B(A[501]), .Z(n1108) );
  XOR U1663 ( .A(A[500]), .B(n1109), .Z(O[500]) );
  AND U1664 ( .A(S), .B(n1110), .Z(n1109) );
  XOR U1665 ( .A(B[500]), .B(A[500]), .Z(n1110) );
  XOR U1666 ( .A(A[4]), .B(n1111), .Z(O[4]) );
  AND U1667 ( .A(S), .B(n1112), .Z(n1111) );
  XOR U1668 ( .A(B[4]), .B(A[4]), .Z(n1112) );
  XOR U1669 ( .A(A[49]), .B(n1113), .Z(O[49]) );
  AND U1670 ( .A(S), .B(n1114), .Z(n1113) );
  XOR U1671 ( .A(B[49]), .B(A[49]), .Z(n1114) );
  XOR U1672 ( .A(A[499]), .B(n1115), .Z(O[499]) );
  AND U1673 ( .A(S), .B(n1116), .Z(n1115) );
  XOR U1674 ( .A(B[499]), .B(A[499]), .Z(n1116) );
  XOR U1675 ( .A(A[498]), .B(n1117), .Z(O[498]) );
  AND U1676 ( .A(S), .B(n1118), .Z(n1117) );
  XOR U1677 ( .A(B[498]), .B(A[498]), .Z(n1118) );
  XOR U1678 ( .A(A[497]), .B(n1119), .Z(O[497]) );
  AND U1679 ( .A(S), .B(n1120), .Z(n1119) );
  XOR U1680 ( .A(B[497]), .B(A[497]), .Z(n1120) );
  XOR U1681 ( .A(A[496]), .B(n1121), .Z(O[496]) );
  AND U1682 ( .A(S), .B(n1122), .Z(n1121) );
  XOR U1683 ( .A(B[496]), .B(A[496]), .Z(n1122) );
  XOR U1684 ( .A(A[495]), .B(n1123), .Z(O[495]) );
  AND U1685 ( .A(S), .B(n1124), .Z(n1123) );
  XOR U1686 ( .A(B[495]), .B(A[495]), .Z(n1124) );
  XOR U1687 ( .A(A[494]), .B(n1125), .Z(O[494]) );
  AND U1688 ( .A(S), .B(n1126), .Z(n1125) );
  XOR U1689 ( .A(B[494]), .B(A[494]), .Z(n1126) );
  XOR U1690 ( .A(A[493]), .B(n1127), .Z(O[493]) );
  AND U1691 ( .A(S), .B(n1128), .Z(n1127) );
  XOR U1692 ( .A(B[493]), .B(A[493]), .Z(n1128) );
  XOR U1693 ( .A(A[492]), .B(n1129), .Z(O[492]) );
  AND U1694 ( .A(S), .B(n1130), .Z(n1129) );
  XOR U1695 ( .A(B[492]), .B(A[492]), .Z(n1130) );
  XOR U1696 ( .A(A[491]), .B(n1131), .Z(O[491]) );
  AND U1697 ( .A(S), .B(n1132), .Z(n1131) );
  XOR U1698 ( .A(B[491]), .B(A[491]), .Z(n1132) );
  XOR U1699 ( .A(A[490]), .B(n1133), .Z(O[490]) );
  AND U1700 ( .A(S), .B(n1134), .Z(n1133) );
  XOR U1701 ( .A(B[490]), .B(A[490]), .Z(n1134) );
  XOR U1702 ( .A(A[48]), .B(n1135), .Z(O[48]) );
  AND U1703 ( .A(S), .B(n1136), .Z(n1135) );
  XOR U1704 ( .A(B[48]), .B(A[48]), .Z(n1136) );
  XOR U1705 ( .A(A[489]), .B(n1137), .Z(O[489]) );
  AND U1706 ( .A(S), .B(n1138), .Z(n1137) );
  XOR U1707 ( .A(B[489]), .B(A[489]), .Z(n1138) );
  XOR U1708 ( .A(A[488]), .B(n1139), .Z(O[488]) );
  AND U1709 ( .A(S), .B(n1140), .Z(n1139) );
  XOR U1710 ( .A(B[488]), .B(A[488]), .Z(n1140) );
  XOR U1711 ( .A(A[487]), .B(n1141), .Z(O[487]) );
  AND U1712 ( .A(S), .B(n1142), .Z(n1141) );
  XOR U1713 ( .A(B[487]), .B(A[487]), .Z(n1142) );
  XOR U1714 ( .A(A[486]), .B(n1143), .Z(O[486]) );
  AND U1715 ( .A(S), .B(n1144), .Z(n1143) );
  XOR U1716 ( .A(B[486]), .B(A[486]), .Z(n1144) );
  XOR U1717 ( .A(A[485]), .B(n1145), .Z(O[485]) );
  AND U1718 ( .A(S), .B(n1146), .Z(n1145) );
  XOR U1719 ( .A(B[485]), .B(A[485]), .Z(n1146) );
  XOR U1720 ( .A(A[484]), .B(n1147), .Z(O[484]) );
  AND U1721 ( .A(S), .B(n1148), .Z(n1147) );
  XOR U1722 ( .A(B[484]), .B(A[484]), .Z(n1148) );
  XOR U1723 ( .A(A[483]), .B(n1149), .Z(O[483]) );
  AND U1724 ( .A(S), .B(n1150), .Z(n1149) );
  XOR U1725 ( .A(B[483]), .B(A[483]), .Z(n1150) );
  XOR U1726 ( .A(A[482]), .B(n1151), .Z(O[482]) );
  AND U1727 ( .A(S), .B(n1152), .Z(n1151) );
  XOR U1728 ( .A(B[482]), .B(A[482]), .Z(n1152) );
  XOR U1729 ( .A(A[481]), .B(n1153), .Z(O[481]) );
  AND U1730 ( .A(S), .B(n1154), .Z(n1153) );
  XOR U1731 ( .A(B[481]), .B(A[481]), .Z(n1154) );
  XOR U1732 ( .A(A[480]), .B(n1155), .Z(O[480]) );
  AND U1733 ( .A(S), .B(n1156), .Z(n1155) );
  XOR U1734 ( .A(B[480]), .B(A[480]), .Z(n1156) );
  XOR U1735 ( .A(A[47]), .B(n1157), .Z(O[47]) );
  AND U1736 ( .A(S), .B(n1158), .Z(n1157) );
  XOR U1737 ( .A(B[47]), .B(A[47]), .Z(n1158) );
  XOR U1738 ( .A(A[479]), .B(n1159), .Z(O[479]) );
  AND U1739 ( .A(S), .B(n1160), .Z(n1159) );
  XOR U1740 ( .A(B[479]), .B(A[479]), .Z(n1160) );
  XOR U1741 ( .A(A[478]), .B(n1161), .Z(O[478]) );
  AND U1742 ( .A(S), .B(n1162), .Z(n1161) );
  XOR U1743 ( .A(B[478]), .B(A[478]), .Z(n1162) );
  XOR U1744 ( .A(A[477]), .B(n1163), .Z(O[477]) );
  AND U1745 ( .A(S), .B(n1164), .Z(n1163) );
  XOR U1746 ( .A(B[477]), .B(A[477]), .Z(n1164) );
  XOR U1747 ( .A(A[476]), .B(n1165), .Z(O[476]) );
  AND U1748 ( .A(S), .B(n1166), .Z(n1165) );
  XOR U1749 ( .A(B[476]), .B(A[476]), .Z(n1166) );
  XOR U1750 ( .A(A[475]), .B(n1167), .Z(O[475]) );
  AND U1751 ( .A(S), .B(n1168), .Z(n1167) );
  XOR U1752 ( .A(B[475]), .B(A[475]), .Z(n1168) );
  XOR U1753 ( .A(A[474]), .B(n1169), .Z(O[474]) );
  AND U1754 ( .A(S), .B(n1170), .Z(n1169) );
  XOR U1755 ( .A(B[474]), .B(A[474]), .Z(n1170) );
  XOR U1756 ( .A(A[473]), .B(n1171), .Z(O[473]) );
  AND U1757 ( .A(S), .B(n1172), .Z(n1171) );
  XOR U1758 ( .A(B[473]), .B(A[473]), .Z(n1172) );
  XOR U1759 ( .A(A[472]), .B(n1173), .Z(O[472]) );
  AND U1760 ( .A(S), .B(n1174), .Z(n1173) );
  XOR U1761 ( .A(B[472]), .B(A[472]), .Z(n1174) );
  XOR U1762 ( .A(A[471]), .B(n1175), .Z(O[471]) );
  AND U1763 ( .A(S), .B(n1176), .Z(n1175) );
  XOR U1764 ( .A(B[471]), .B(A[471]), .Z(n1176) );
  XOR U1765 ( .A(A[470]), .B(n1177), .Z(O[470]) );
  AND U1766 ( .A(S), .B(n1178), .Z(n1177) );
  XOR U1767 ( .A(B[470]), .B(A[470]), .Z(n1178) );
  XOR U1768 ( .A(A[46]), .B(n1179), .Z(O[46]) );
  AND U1769 ( .A(S), .B(n1180), .Z(n1179) );
  XOR U1770 ( .A(B[46]), .B(A[46]), .Z(n1180) );
  XOR U1771 ( .A(A[469]), .B(n1181), .Z(O[469]) );
  AND U1772 ( .A(S), .B(n1182), .Z(n1181) );
  XOR U1773 ( .A(B[469]), .B(A[469]), .Z(n1182) );
  XOR U1774 ( .A(A[468]), .B(n1183), .Z(O[468]) );
  AND U1775 ( .A(S), .B(n1184), .Z(n1183) );
  XOR U1776 ( .A(B[468]), .B(A[468]), .Z(n1184) );
  XOR U1777 ( .A(A[467]), .B(n1185), .Z(O[467]) );
  AND U1778 ( .A(S), .B(n1186), .Z(n1185) );
  XOR U1779 ( .A(B[467]), .B(A[467]), .Z(n1186) );
  XOR U1780 ( .A(A[466]), .B(n1187), .Z(O[466]) );
  AND U1781 ( .A(S), .B(n1188), .Z(n1187) );
  XOR U1782 ( .A(B[466]), .B(A[466]), .Z(n1188) );
  XOR U1783 ( .A(A[465]), .B(n1189), .Z(O[465]) );
  AND U1784 ( .A(S), .B(n1190), .Z(n1189) );
  XOR U1785 ( .A(B[465]), .B(A[465]), .Z(n1190) );
  XOR U1786 ( .A(A[464]), .B(n1191), .Z(O[464]) );
  AND U1787 ( .A(S), .B(n1192), .Z(n1191) );
  XOR U1788 ( .A(B[464]), .B(A[464]), .Z(n1192) );
  XOR U1789 ( .A(A[463]), .B(n1193), .Z(O[463]) );
  AND U1790 ( .A(S), .B(n1194), .Z(n1193) );
  XOR U1791 ( .A(B[463]), .B(A[463]), .Z(n1194) );
  XOR U1792 ( .A(A[462]), .B(n1195), .Z(O[462]) );
  AND U1793 ( .A(S), .B(n1196), .Z(n1195) );
  XOR U1794 ( .A(B[462]), .B(A[462]), .Z(n1196) );
  XOR U1795 ( .A(A[461]), .B(n1197), .Z(O[461]) );
  AND U1796 ( .A(S), .B(n1198), .Z(n1197) );
  XOR U1797 ( .A(B[461]), .B(A[461]), .Z(n1198) );
  XOR U1798 ( .A(A[460]), .B(n1199), .Z(O[460]) );
  AND U1799 ( .A(S), .B(n1200), .Z(n1199) );
  XOR U1800 ( .A(B[460]), .B(A[460]), .Z(n1200) );
  XOR U1801 ( .A(A[45]), .B(n1201), .Z(O[45]) );
  AND U1802 ( .A(S), .B(n1202), .Z(n1201) );
  XOR U1803 ( .A(B[45]), .B(A[45]), .Z(n1202) );
  XOR U1804 ( .A(A[459]), .B(n1203), .Z(O[459]) );
  AND U1805 ( .A(S), .B(n1204), .Z(n1203) );
  XOR U1806 ( .A(B[459]), .B(A[459]), .Z(n1204) );
  XOR U1807 ( .A(A[458]), .B(n1205), .Z(O[458]) );
  AND U1808 ( .A(S), .B(n1206), .Z(n1205) );
  XOR U1809 ( .A(B[458]), .B(A[458]), .Z(n1206) );
  XOR U1810 ( .A(A[457]), .B(n1207), .Z(O[457]) );
  AND U1811 ( .A(S), .B(n1208), .Z(n1207) );
  XOR U1812 ( .A(B[457]), .B(A[457]), .Z(n1208) );
  XOR U1813 ( .A(A[456]), .B(n1209), .Z(O[456]) );
  AND U1814 ( .A(S), .B(n1210), .Z(n1209) );
  XOR U1815 ( .A(B[456]), .B(A[456]), .Z(n1210) );
  XOR U1816 ( .A(A[455]), .B(n1211), .Z(O[455]) );
  AND U1817 ( .A(S), .B(n1212), .Z(n1211) );
  XOR U1818 ( .A(B[455]), .B(A[455]), .Z(n1212) );
  XOR U1819 ( .A(A[454]), .B(n1213), .Z(O[454]) );
  AND U1820 ( .A(S), .B(n1214), .Z(n1213) );
  XOR U1821 ( .A(B[454]), .B(A[454]), .Z(n1214) );
  XOR U1822 ( .A(A[453]), .B(n1215), .Z(O[453]) );
  AND U1823 ( .A(S), .B(n1216), .Z(n1215) );
  XOR U1824 ( .A(B[453]), .B(A[453]), .Z(n1216) );
  XOR U1825 ( .A(A[452]), .B(n1217), .Z(O[452]) );
  AND U1826 ( .A(S), .B(n1218), .Z(n1217) );
  XOR U1827 ( .A(B[452]), .B(A[452]), .Z(n1218) );
  XOR U1828 ( .A(A[451]), .B(n1219), .Z(O[451]) );
  AND U1829 ( .A(S), .B(n1220), .Z(n1219) );
  XOR U1830 ( .A(B[451]), .B(A[451]), .Z(n1220) );
  XOR U1831 ( .A(A[450]), .B(n1221), .Z(O[450]) );
  AND U1832 ( .A(S), .B(n1222), .Z(n1221) );
  XOR U1833 ( .A(B[450]), .B(A[450]), .Z(n1222) );
  XOR U1834 ( .A(A[44]), .B(n1223), .Z(O[44]) );
  AND U1835 ( .A(S), .B(n1224), .Z(n1223) );
  XOR U1836 ( .A(B[44]), .B(A[44]), .Z(n1224) );
  XOR U1837 ( .A(A[449]), .B(n1225), .Z(O[449]) );
  AND U1838 ( .A(S), .B(n1226), .Z(n1225) );
  XOR U1839 ( .A(B[449]), .B(A[449]), .Z(n1226) );
  XOR U1840 ( .A(A[448]), .B(n1227), .Z(O[448]) );
  AND U1841 ( .A(S), .B(n1228), .Z(n1227) );
  XOR U1842 ( .A(B[448]), .B(A[448]), .Z(n1228) );
  XOR U1843 ( .A(A[447]), .B(n1229), .Z(O[447]) );
  AND U1844 ( .A(S), .B(n1230), .Z(n1229) );
  XOR U1845 ( .A(B[447]), .B(A[447]), .Z(n1230) );
  XOR U1846 ( .A(A[446]), .B(n1231), .Z(O[446]) );
  AND U1847 ( .A(S), .B(n1232), .Z(n1231) );
  XOR U1848 ( .A(B[446]), .B(A[446]), .Z(n1232) );
  XOR U1849 ( .A(A[445]), .B(n1233), .Z(O[445]) );
  AND U1850 ( .A(S), .B(n1234), .Z(n1233) );
  XOR U1851 ( .A(B[445]), .B(A[445]), .Z(n1234) );
  XOR U1852 ( .A(A[444]), .B(n1235), .Z(O[444]) );
  AND U1853 ( .A(S), .B(n1236), .Z(n1235) );
  XOR U1854 ( .A(B[444]), .B(A[444]), .Z(n1236) );
  XOR U1855 ( .A(A[443]), .B(n1237), .Z(O[443]) );
  AND U1856 ( .A(S), .B(n1238), .Z(n1237) );
  XOR U1857 ( .A(B[443]), .B(A[443]), .Z(n1238) );
  XOR U1858 ( .A(A[442]), .B(n1239), .Z(O[442]) );
  AND U1859 ( .A(S), .B(n1240), .Z(n1239) );
  XOR U1860 ( .A(B[442]), .B(A[442]), .Z(n1240) );
  XOR U1861 ( .A(A[441]), .B(n1241), .Z(O[441]) );
  AND U1862 ( .A(S), .B(n1242), .Z(n1241) );
  XOR U1863 ( .A(B[441]), .B(A[441]), .Z(n1242) );
  XOR U1864 ( .A(A[440]), .B(n1243), .Z(O[440]) );
  AND U1865 ( .A(S), .B(n1244), .Z(n1243) );
  XOR U1866 ( .A(B[440]), .B(A[440]), .Z(n1244) );
  XOR U1867 ( .A(A[43]), .B(n1245), .Z(O[43]) );
  AND U1868 ( .A(S), .B(n1246), .Z(n1245) );
  XOR U1869 ( .A(B[43]), .B(A[43]), .Z(n1246) );
  XOR U1870 ( .A(A[439]), .B(n1247), .Z(O[439]) );
  AND U1871 ( .A(S), .B(n1248), .Z(n1247) );
  XOR U1872 ( .A(B[439]), .B(A[439]), .Z(n1248) );
  XOR U1873 ( .A(A[438]), .B(n1249), .Z(O[438]) );
  AND U1874 ( .A(S), .B(n1250), .Z(n1249) );
  XOR U1875 ( .A(B[438]), .B(A[438]), .Z(n1250) );
  XOR U1876 ( .A(A[437]), .B(n1251), .Z(O[437]) );
  AND U1877 ( .A(S), .B(n1252), .Z(n1251) );
  XOR U1878 ( .A(B[437]), .B(A[437]), .Z(n1252) );
  XOR U1879 ( .A(A[436]), .B(n1253), .Z(O[436]) );
  AND U1880 ( .A(S), .B(n1254), .Z(n1253) );
  XOR U1881 ( .A(B[436]), .B(A[436]), .Z(n1254) );
  XOR U1882 ( .A(A[435]), .B(n1255), .Z(O[435]) );
  AND U1883 ( .A(S), .B(n1256), .Z(n1255) );
  XOR U1884 ( .A(B[435]), .B(A[435]), .Z(n1256) );
  XOR U1885 ( .A(A[434]), .B(n1257), .Z(O[434]) );
  AND U1886 ( .A(S), .B(n1258), .Z(n1257) );
  XOR U1887 ( .A(B[434]), .B(A[434]), .Z(n1258) );
  XOR U1888 ( .A(A[433]), .B(n1259), .Z(O[433]) );
  AND U1889 ( .A(S), .B(n1260), .Z(n1259) );
  XOR U1890 ( .A(B[433]), .B(A[433]), .Z(n1260) );
  XOR U1891 ( .A(A[432]), .B(n1261), .Z(O[432]) );
  AND U1892 ( .A(S), .B(n1262), .Z(n1261) );
  XOR U1893 ( .A(B[432]), .B(A[432]), .Z(n1262) );
  XOR U1894 ( .A(A[431]), .B(n1263), .Z(O[431]) );
  AND U1895 ( .A(S), .B(n1264), .Z(n1263) );
  XOR U1896 ( .A(B[431]), .B(A[431]), .Z(n1264) );
  XOR U1897 ( .A(A[430]), .B(n1265), .Z(O[430]) );
  AND U1898 ( .A(S), .B(n1266), .Z(n1265) );
  XOR U1899 ( .A(B[430]), .B(A[430]), .Z(n1266) );
  XOR U1900 ( .A(A[42]), .B(n1267), .Z(O[42]) );
  AND U1901 ( .A(S), .B(n1268), .Z(n1267) );
  XOR U1902 ( .A(B[42]), .B(A[42]), .Z(n1268) );
  XOR U1903 ( .A(A[429]), .B(n1269), .Z(O[429]) );
  AND U1904 ( .A(S), .B(n1270), .Z(n1269) );
  XOR U1905 ( .A(B[429]), .B(A[429]), .Z(n1270) );
  XOR U1906 ( .A(A[428]), .B(n1271), .Z(O[428]) );
  AND U1907 ( .A(S), .B(n1272), .Z(n1271) );
  XOR U1908 ( .A(B[428]), .B(A[428]), .Z(n1272) );
  XOR U1909 ( .A(A[427]), .B(n1273), .Z(O[427]) );
  AND U1910 ( .A(S), .B(n1274), .Z(n1273) );
  XOR U1911 ( .A(B[427]), .B(A[427]), .Z(n1274) );
  XOR U1912 ( .A(A[426]), .B(n1275), .Z(O[426]) );
  AND U1913 ( .A(S), .B(n1276), .Z(n1275) );
  XOR U1914 ( .A(B[426]), .B(A[426]), .Z(n1276) );
  XOR U1915 ( .A(A[425]), .B(n1277), .Z(O[425]) );
  AND U1916 ( .A(S), .B(n1278), .Z(n1277) );
  XOR U1917 ( .A(B[425]), .B(A[425]), .Z(n1278) );
  XOR U1918 ( .A(A[424]), .B(n1279), .Z(O[424]) );
  AND U1919 ( .A(S), .B(n1280), .Z(n1279) );
  XOR U1920 ( .A(B[424]), .B(A[424]), .Z(n1280) );
  XOR U1921 ( .A(A[423]), .B(n1281), .Z(O[423]) );
  AND U1922 ( .A(S), .B(n1282), .Z(n1281) );
  XOR U1923 ( .A(B[423]), .B(A[423]), .Z(n1282) );
  XOR U1924 ( .A(A[422]), .B(n1283), .Z(O[422]) );
  AND U1925 ( .A(S), .B(n1284), .Z(n1283) );
  XOR U1926 ( .A(B[422]), .B(A[422]), .Z(n1284) );
  XOR U1927 ( .A(A[421]), .B(n1285), .Z(O[421]) );
  AND U1928 ( .A(S), .B(n1286), .Z(n1285) );
  XOR U1929 ( .A(B[421]), .B(A[421]), .Z(n1286) );
  XOR U1930 ( .A(A[420]), .B(n1287), .Z(O[420]) );
  AND U1931 ( .A(S), .B(n1288), .Z(n1287) );
  XOR U1932 ( .A(B[420]), .B(A[420]), .Z(n1288) );
  XOR U1933 ( .A(A[41]), .B(n1289), .Z(O[41]) );
  AND U1934 ( .A(S), .B(n1290), .Z(n1289) );
  XOR U1935 ( .A(B[41]), .B(A[41]), .Z(n1290) );
  XOR U1936 ( .A(A[419]), .B(n1291), .Z(O[419]) );
  AND U1937 ( .A(S), .B(n1292), .Z(n1291) );
  XOR U1938 ( .A(B[419]), .B(A[419]), .Z(n1292) );
  XOR U1939 ( .A(A[418]), .B(n1293), .Z(O[418]) );
  AND U1940 ( .A(S), .B(n1294), .Z(n1293) );
  XOR U1941 ( .A(B[418]), .B(A[418]), .Z(n1294) );
  XOR U1942 ( .A(A[417]), .B(n1295), .Z(O[417]) );
  AND U1943 ( .A(S), .B(n1296), .Z(n1295) );
  XOR U1944 ( .A(B[417]), .B(A[417]), .Z(n1296) );
  XOR U1945 ( .A(A[416]), .B(n1297), .Z(O[416]) );
  AND U1946 ( .A(S), .B(n1298), .Z(n1297) );
  XOR U1947 ( .A(B[416]), .B(A[416]), .Z(n1298) );
  XOR U1948 ( .A(A[415]), .B(n1299), .Z(O[415]) );
  AND U1949 ( .A(S), .B(n1300), .Z(n1299) );
  XOR U1950 ( .A(B[415]), .B(A[415]), .Z(n1300) );
  XOR U1951 ( .A(A[414]), .B(n1301), .Z(O[414]) );
  AND U1952 ( .A(S), .B(n1302), .Z(n1301) );
  XOR U1953 ( .A(B[414]), .B(A[414]), .Z(n1302) );
  XOR U1954 ( .A(A[413]), .B(n1303), .Z(O[413]) );
  AND U1955 ( .A(S), .B(n1304), .Z(n1303) );
  XOR U1956 ( .A(B[413]), .B(A[413]), .Z(n1304) );
  XOR U1957 ( .A(A[412]), .B(n1305), .Z(O[412]) );
  AND U1958 ( .A(S), .B(n1306), .Z(n1305) );
  XOR U1959 ( .A(B[412]), .B(A[412]), .Z(n1306) );
  XOR U1960 ( .A(A[411]), .B(n1307), .Z(O[411]) );
  AND U1961 ( .A(S), .B(n1308), .Z(n1307) );
  XOR U1962 ( .A(B[411]), .B(A[411]), .Z(n1308) );
  XOR U1963 ( .A(A[410]), .B(n1309), .Z(O[410]) );
  AND U1964 ( .A(S), .B(n1310), .Z(n1309) );
  XOR U1965 ( .A(B[410]), .B(A[410]), .Z(n1310) );
  XOR U1966 ( .A(A[40]), .B(n1311), .Z(O[40]) );
  AND U1967 ( .A(S), .B(n1312), .Z(n1311) );
  XOR U1968 ( .A(B[40]), .B(A[40]), .Z(n1312) );
  XOR U1969 ( .A(A[409]), .B(n1313), .Z(O[409]) );
  AND U1970 ( .A(S), .B(n1314), .Z(n1313) );
  XOR U1971 ( .A(B[409]), .B(A[409]), .Z(n1314) );
  XOR U1972 ( .A(A[408]), .B(n1315), .Z(O[408]) );
  AND U1973 ( .A(S), .B(n1316), .Z(n1315) );
  XOR U1974 ( .A(B[408]), .B(A[408]), .Z(n1316) );
  XOR U1975 ( .A(A[407]), .B(n1317), .Z(O[407]) );
  AND U1976 ( .A(S), .B(n1318), .Z(n1317) );
  XOR U1977 ( .A(B[407]), .B(A[407]), .Z(n1318) );
  XOR U1978 ( .A(A[406]), .B(n1319), .Z(O[406]) );
  AND U1979 ( .A(S), .B(n1320), .Z(n1319) );
  XOR U1980 ( .A(B[406]), .B(A[406]), .Z(n1320) );
  XOR U1981 ( .A(A[405]), .B(n1321), .Z(O[405]) );
  AND U1982 ( .A(S), .B(n1322), .Z(n1321) );
  XOR U1983 ( .A(B[405]), .B(A[405]), .Z(n1322) );
  XOR U1984 ( .A(A[404]), .B(n1323), .Z(O[404]) );
  AND U1985 ( .A(S), .B(n1324), .Z(n1323) );
  XOR U1986 ( .A(B[404]), .B(A[404]), .Z(n1324) );
  XOR U1987 ( .A(A[403]), .B(n1325), .Z(O[403]) );
  AND U1988 ( .A(S), .B(n1326), .Z(n1325) );
  XOR U1989 ( .A(B[403]), .B(A[403]), .Z(n1326) );
  XOR U1990 ( .A(A[402]), .B(n1327), .Z(O[402]) );
  AND U1991 ( .A(S), .B(n1328), .Z(n1327) );
  XOR U1992 ( .A(B[402]), .B(A[402]), .Z(n1328) );
  XOR U1993 ( .A(A[401]), .B(n1329), .Z(O[401]) );
  AND U1994 ( .A(S), .B(n1330), .Z(n1329) );
  XOR U1995 ( .A(B[401]), .B(A[401]), .Z(n1330) );
  XOR U1996 ( .A(A[400]), .B(n1331), .Z(O[400]) );
  AND U1997 ( .A(S), .B(n1332), .Z(n1331) );
  XOR U1998 ( .A(B[400]), .B(A[400]), .Z(n1332) );
  XOR U1999 ( .A(A[3]), .B(n1333), .Z(O[3]) );
  AND U2000 ( .A(S), .B(n1334), .Z(n1333) );
  XOR U2001 ( .A(B[3]), .B(A[3]), .Z(n1334) );
  XOR U2002 ( .A(A[39]), .B(n1335), .Z(O[39]) );
  AND U2003 ( .A(S), .B(n1336), .Z(n1335) );
  XOR U2004 ( .A(B[39]), .B(A[39]), .Z(n1336) );
  XOR U2005 ( .A(A[399]), .B(n1337), .Z(O[399]) );
  AND U2006 ( .A(S), .B(n1338), .Z(n1337) );
  XOR U2007 ( .A(B[399]), .B(A[399]), .Z(n1338) );
  XOR U2008 ( .A(A[398]), .B(n1339), .Z(O[398]) );
  AND U2009 ( .A(S), .B(n1340), .Z(n1339) );
  XOR U2010 ( .A(B[398]), .B(A[398]), .Z(n1340) );
  XOR U2011 ( .A(A[397]), .B(n1341), .Z(O[397]) );
  AND U2012 ( .A(S), .B(n1342), .Z(n1341) );
  XOR U2013 ( .A(B[397]), .B(A[397]), .Z(n1342) );
  XOR U2014 ( .A(A[396]), .B(n1343), .Z(O[396]) );
  AND U2015 ( .A(S), .B(n1344), .Z(n1343) );
  XOR U2016 ( .A(B[396]), .B(A[396]), .Z(n1344) );
  XOR U2017 ( .A(A[395]), .B(n1345), .Z(O[395]) );
  AND U2018 ( .A(S), .B(n1346), .Z(n1345) );
  XOR U2019 ( .A(B[395]), .B(A[395]), .Z(n1346) );
  XOR U2020 ( .A(A[394]), .B(n1347), .Z(O[394]) );
  AND U2021 ( .A(S), .B(n1348), .Z(n1347) );
  XOR U2022 ( .A(B[394]), .B(A[394]), .Z(n1348) );
  XOR U2023 ( .A(A[393]), .B(n1349), .Z(O[393]) );
  AND U2024 ( .A(S), .B(n1350), .Z(n1349) );
  XOR U2025 ( .A(B[393]), .B(A[393]), .Z(n1350) );
  XOR U2026 ( .A(A[392]), .B(n1351), .Z(O[392]) );
  AND U2027 ( .A(S), .B(n1352), .Z(n1351) );
  XOR U2028 ( .A(B[392]), .B(A[392]), .Z(n1352) );
  XOR U2029 ( .A(A[391]), .B(n1353), .Z(O[391]) );
  AND U2030 ( .A(S), .B(n1354), .Z(n1353) );
  XOR U2031 ( .A(B[391]), .B(A[391]), .Z(n1354) );
  XOR U2032 ( .A(A[390]), .B(n1355), .Z(O[390]) );
  AND U2033 ( .A(S), .B(n1356), .Z(n1355) );
  XOR U2034 ( .A(B[390]), .B(A[390]), .Z(n1356) );
  XOR U2035 ( .A(A[38]), .B(n1357), .Z(O[38]) );
  AND U2036 ( .A(S), .B(n1358), .Z(n1357) );
  XOR U2037 ( .A(B[38]), .B(A[38]), .Z(n1358) );
  XOR U2038 ( .A(A[389]), .B(n1359), .Z(O[389]) );
  AND U2039 ( .A(S), .B(n1360), .Z(n1359) );
  XOR U2040 ( .A(B[389]), .B(A[389]), .Z(n1360) );
  XOR U2041 ( .A(A[388]), .B(n1361), .Z(O[388]) );
  AND U2042 ( .A(S), .B(n1362), .Z(n1361) );
  XOR U2043 ( .A(B[388]), .B(A[388]), .Z(n1362) );
  XOR U2044 ( .A(A[387]), .B(n1363), .Z(O[387]) );
  AND U2045 ( .A(S), .B(n1364), .Z(n1363) );
  XOR U2046 ( .A(B[387]), .B(A[387]), .Z(n1364) );
  XOR U2047 ( .A(A[386]), .B(n1365), .Z(O[386]) );
  AND U2048 ( .A(S), .B(n1366), .Z(n1365) );
  XOR U2049 ( .A(B[386]), .B(A[386]), .Z(n1366) );
  XOR U2050 ( .A(A[385]), .B(n1367), .Z(O[385]) );
  AND U2051 ( .A(S), .B(n1368), .Z(n1367) );
  XOR U2052 ( .A(B[385]), .B(A[385]), .Z(n1368) );
  XOR U2053 ( .A(A[384]), .B(n1369), .Z(O[384]) );
  AND U2054 ( .A(S), .B(n1370), .Z(n1369) );
  XOR U2055 ( .A(B[384]), .B(A[384]), .Z(n1370) );
  XOR U2056 ( .A(A[383]), .B(n1371), .Z(O[383]) );
  AND U2057 ( .A(S), .B(n1372), .Z(n1371) );
  XOR U2058 ( .A(B[383]), .B(A[383]), .Z(n1372) );
  XOR U2059 ( .A(A[382]), .B(n1373), .Z(O[382]) );
  AND U2060 ( .A(S), .B(n1374), .Z(n1373) );
  XOR U2061 ( .A(B[382]), .B(A[382]), .Z(n1374) );
  XOR U2062 ( .A(A[381]), .B(n1375), .Z(O[381]) );
  AND U2063 ( .A(S), .B(n1376), .Z(n1375) );
  XOR U2064 ( .A(B[381]), .B(A[381]), .Z(n1376) );
  XOR U2065 ( .A(A[380]), .B(n1377), .Z(O[380]) );
  AND U2066 ( .A(S), .B(n1378), .Z(n1377) );
  XOR U2067 ( .A(B[380]), .B(A[380]), .Z(n1378) );
  XOR U2068 ( .A(A[37]), .B(n1379), .Z(O[37]) );
  AND U2069 ( .A(S), .B(n1380), .Z(n1379) );
  XOR U2070 ( .A(B[37]), .B(A[37]), .Z(n1380) );
  XOR U2071 ( .A(A[379]), .B(n1381), .Z(O[379]) );
  AND U2072 ( .A(S), .B(n1382), .Z(n1381) );
  XOR U2073 ( .A(B[379]), .B(A[379]), .Z(n1382) );
  XOR U2074 ( .A(A[378]), .B(n1383), .Z(O[378]) );
  AND U2075 ( .A(S), .B(n1384), .Z(n1383) );
  XOR U2076 ( .A(B[378]), .B(A[378]), .Z(n1384) );
  XOR U2077 ( .A(A[377]), .B(n1385), .Z(O[377]) );
  AND U2078 ( .A(S), .B(n1386), .Z(n1385) );
  XOR U2079 ( .A(B[377]), .B(A[377]), .Z(n1386) );
  XOR U2080 ( .A(A[376]), .B(n1387), .Z(O[376]) );
  AND U2081 ( .A(S), .B(n1388), .Z(n1387) );
  XOR U2082 ( .A(B[376]), .B(A[376]), .Z(n1388) );
  XOR U2083 ( .A(A[375]), .B(n1389), .Z(O[375]) );
  AND U2084 ( .A(S), .B(n1390), .Z(n1389) );
  XOR U2085 ( .A(B[375]), .B(A[375]), .Z(n1390) );
  XOR U2086 ( .A(A[374]), .B(n1391), .Z(O[374]) );
  AND U2087 ( .A(S), .B(n1392), .Z(n1391) );
  XOR U2088 ( .A(B[374]), .B(A[374]), .Z(n1392) );
  XOR U2089 ( .A(A[373]), .B(n1393), .Z(O[373]) );
  AND U2090 ( .A(S), .B(n1394), .Z(n1393) );
  XOR U2091 ( .A(B[373]), .B(A[373]), .Z(n1394) );
  XOR U2092 ( .A(A[372]), .B(n1395), .Z(O[372]) );
  AND U2093 ( .A(S), .B(n1396), .Z(n1395) );
  XOR U2094 ( .A(B[372]), .B(A[372]), .Z(n1396) );
  XOR U2095 ( .A(A[371]), .B(n1397), .Z(O[371]) );
  AND U2096 ( .A(S), .B(n1398), .Z(n1397) );
  XOR U2097 ( .A(B[371]), .B(A[371]), .Z(n1398) );
  XOR U2098 ( .A(A[370]), .B(n1399), .Z(O[370]) );
  AND U2099 ( .A(S), .B(n1400), .Z(n1399) );
  XOR U2100 ( .A(B[370]), .B(A[370]), .Z(n1400) );
  XOR U2101 ( .A(A[36]), .B(n1401), .Z(O[36]) );
  AND U2102 ( .A(S), .B(n1402), .Z(n1401) );
  XOR U2103 ( .A(B[36]), .B(A[36]), .Z(n1402) );
  XOR U2104 ( .A(A[369]), .B(n1403), .Z(O[369]) );
  AND U2105 ( .A(S), .B(n1404), .Z(n1403) );
  XOR U2106 ( .A(B[369]), .B(A[369]), .Z(n1404) );
  XOR U2107 ( .A(A[368]), .B(n1405), .Z(O[368]) );
  AND U2108 ( .A(S), .B(n1406), .Z(n1405) );
  XOR U2109 ( .A(B[368]), .B(A[368]), .Z(n1406) );
  XOR U2110 ( .A(A[367]), .B(n1407), .Z(O[367]) );
  AND U2111 ( .A(S), .B(n1408), .Z(n1407) );
  XOR U2112 ( .A(B[367]), .B(A[367]), .Z(n1408) );
  XOR U2113 ( .A(A[366]), .B(n1409), .Z(O[366]) );
  AND U2114 ( .A(S), .B(n1410), .Z(n1409) );
  XOR U2115 ( .A(B[366]), .B(A[366]), .Z(n1410) );
  XOR U2116 ( .A(A[365]), .B(n1411), .Z(O[365]) );
  AND U2117 ( .A(S), .B(n1412), .Z(n1411) );
  XOR U2118 ( .A(B[365]), .B(A[365]), .Z(n1412) );
  XOR U2119 ( .A(A[364]), .B(n1413), .Z(O[364]) );
  AND U2120 ( .A(S), .B(n1414), .Z(n1413) );
  XOR U2121 ( .A(B[364]), .B(A[364]), .Z(n1414) );
  XOR U2122 ( .A(A[363]), .B(n1415), .Z(O[363]) );
  AND U2123 ( .A(S), .B(n1416), .Z(n1415) );
  XOR U2124 ( .A(B[363]), .B(A[363]), .Z(n1416) );
  XOR U2125 ( .A(A[362]), .B(n1417), .Z(O[362]) );
  AND U2126 ( .A(S), .B(n1418), .Z(n1417) );
  XOR U2127 ( .A(B[362]), .B(A[362]), .Z(n1418) );
  XOR U2128 ( .A(A[361]), .B(n1419), .Z(O[361]) );
  AND U2129 ( .A(S), .B(n1420), .Z(n1419) );
  XOR U2130 ( .A(B[361]), .B(A[361]), .Z(n1420) );
  XOR U2131 ( .A(A[360]), .B(n1421), .Z(O[360]) );
  AND U2132 ( .A(S), .B(n1422), .Z(n1421) );
  XOR U2133 ( .A(B[360]), .B(A[360]), .Z(n1422) );
  XOR U2134 ( .A(A[35]), .B(n1423), .Z(O[35]) );
  AND U2135 ( .A(S), .B(n1424), .Z(n1423) );
  XOR U2136 ( .A(B[35]), .B(A[35]), .Z(n1424) );
  XOR U2137 ( .A(A[359]), .B(n1425), .Z(O[359]) );
  AND U2138 ( .A(S), .B(n1426), .Z(n1425) );
  XOR U2139 ( .A(B[359]), .B(A[359]), .Z(n1426) );
  XOR U2140 ( .A(A[358]), .B(n1427), .Z(O[358]) );
  AND U2141 ( .A(S), .B(n1428), .Z(n1427) );
  XOR U2142 ( .A(B[358]), .B(A[358]), .Z(n1428) );
  XOR U2143 ( .A(A[357]), .B(n1429), .Z(O[357]) );
  AND U2144 ( .A(S), .B(n1430), .Z(n1429) );
  XOR U2145 ( .A(B[357]), .B(A[357]), .Z(n1430) );
  XOR U2146 ( .A(A[356]), .B(n1431), .Z(O[356]) );
  AND U2147 ( .A(S), .B(n1432), .Z(n1431) );
  XOR U2148 ( .A(B[356]), .B(A[356]), .Z(n1432) );
  XOR U2149 ( .A(A[355]), .B(n1433), .Z(O[355]) );
  AND U2150 ( .A(S), .B(n1434), .Z(n1433) );
  XOR U2151 ( .A(B[355]), .B(A[355]), .Z(n1434) );
  XOR U2152 ( .A(A[354]), .B(n1435), .Z(O[354]) );
  AND U2153 ( .A(S), .B(n1436), .Z(n1435) );
  XOR U2154 ( .A(B[354]), .B(A[354]), .Z(n1436) );
  XOR U2155 ( .A(A[353]), .B(n1437), .Z(O[353]) );
  AND U2156 ( .A(S), .B(n1438), .Z(n1437) );
  XOR U2157 ( .A(B[353]), .B(A[353]), .Z(n1438) );
  XOR U2158 ( .A(A[352]), .B(n1439), .Z(O[352]) );
  AND U2159 ( .A(S), .B(n1440), .Z(n1439) );
  XOR U2160 ( .A(B[352]), .B(A[352]), .Z(n1440) );
  XOR U2161 ( .A(A[351]), .B(n1441), .Z(O[351]) );
  AND U2162 ( .A(S), .B(n1442), .Z(n1441) );
  XOR U2163 ( .A(B[351]), .B(A[351]), .Z(n1442) );
  XOR U2164 ( .A(A[350]), .B(n1443), .Z(O[350]) );
  AND U2165 ( .A(S), .B(n1444), .Z(n1443) );
  XOR U2166 ( .A(B[350]), .B(A[350]), .Z(n1444) );
  XOR U2167 ( .A(A[34]), .B(n1445), .Z(O[34]) );
  AND U2168 ( .A(S), .B(n1446), .Z(n1445) );
  XOR U2169 ( .A(B[34]), .B(A[34]), .Z(n1446) );
  XOR U2170 ( .A(A[349]), .B(n1447), .Z(O[349]) );
  AND U2171 ( .A(S), .B(n1448), .Z(n1447) );
  XOR U2172 ( .A(B[349]), .B(A[349]), .Z(n1448) );
  XOR U2173 ( .A(A[348]), .B(n1449), .Z(O[348]) );
  AND U2174 ( .A(S), .B(n1450), .Z(n1449) );
  XOR U2175 ( .A(B[348]), .B(A[348]), .Z(n1450) );
  XOR U2176 ( .A(A[347]), .B(n1451), .Z(O[347]) );
  AND U2177 ( .A(S), .B(n1452), .Z(n1451) );
  XOR U2178 ( .A(B[347]), .B(A[347]), .Z(n1452) );
  XOR U2179 ( .A(A[346]), .B(n1453), .Z(O[346]) );
  AND U2180 ( .A(S), .B(n1454), .Z(n1453) );
  XOR U2181 ( .A(B[346]), .B(A[346]), .Z(n1454) );
  XOR U2182 ( .A(A[345]), .B(n1455), .Z(O[345]) );
  AND U2183 ( .A(S), .B(n1456), .Z(n1455) );
  XOR U2184 ( .A(B[345]), .B(A[345]), .Z(n1456) );
  XOR U2185 ( .A(A[344]), .B(n1457), .Z(O[344]) );
  AND U2186 ( .A(S), .B(n1458), .Z(n1457) );
  XOR U2187 ( .A(B[344]), .B(A[344]), .Z(n1458) );
  XOR U2188 ( .A(A[343]), .B(n1459), .Z(O[343]) );
  AND U2189 ( .A(S), .B(n1460), .Z(n1459) );
  XOR U2190 ( .A(B[343]), .B(A[343]), .Z(n1460) );
  XOR U2191 ( .A(A[342]), .B(n1461), .Z(O[342]) );
  AND U2192 ( .A(S), .B(n1462), .Z(n1461) );
  XOR U2193 ( .A(B[342]), .B(A[342]), .Z(n1462) );
  XOR U2194 ( .A(A[341]), .B(n1463), .Z(O[341]) );
  AND U2195 ( .A(S), .B(n1464), .Z(n1463) );
  XOR U2196 ( .A(B[341]), .B(A[341]), .Z(n1464) );
  XOR U2197 ( .A(A[340]), .B(n1465), .Z(O[340]) );
  AND U2198 ( .A(S), .B(n1466), .Z(n1465) );
  XOR U2199 ( .A(B[340]), .B(A[340]), .Z(n1466) );
  XOR U2200 ( .A(A[33]), .B(n1467), .Z(O[33]) );
  AND U2201 ( .A(S), .B(n1468), .Z(n1467) );
  XOR U2202 ( .A(B[33]), .B(A[33]), .Z(n1468) );
  XOR U2203 ( .A(A[339]), .B(n1469), .Z(O[339]) );
  AND U2204 ( .A(S), .B(n1470), .Z(n1469) );
  XOR U2205 ( .A(B[339]), .B(A[339]), .Z(n1470) );
  XOR U2206 ( .A(A[338]), .B(n1471), .Z(O[338]) );
  AND U2207 ( .A(S), .B(n1472), .Z(n1471) );
  XOR U2208 ( .A(B[338]), .B(A[338]), .Z(n1472) );
  XOR U2209 ( .A(A[337]), .B(n1473), .Z(O[337]) );
  AND U2210 ( .A(S), .B(n1474), .Z(n1473) );
  XOR U2211 ( .A(B[337]), .B(A[337]), .Z(n1474) );
  XOR U2212 ( .A(A[336]), .B(n1475), .Z(O[336]) );
  AND U2213 ( .A(S), .B(n1476), .Z(n1475) );
  XOR U2214 ( .A(B[336]), .B(A[336]), .Z(n1476) );
  XOR U2215 ( .A(A[335]), .B(n1477), .Z(O[335]) );
  AND U2216 ( .A(S), .B(n1478), .Z(n1477) );
  XOR U2217 ( .A(B[335]), .B(A[335]), .Z(n1478) );
  XOR U2218 ( .A(A[334]), .B(n1479), .Z(O[334]) );
  AND U2219 ( .A(S), .B(n1480), .Z(n1479) );
  XOR U2220 ( .A(B[334]), .B(A[334]), .Z(n1480) );
  XOR U2221 ( .A(A[333]), .B(n1481), .Z(O[333]) );
  AND U2222 ( .A(S), .B(n1482), .Z(n1481) );
  XOR U2223 ( .A(B[333]), .B(A[333]), .Z(n1482) );
  XOR U2224 ( .A(A[332]), .B(n1483), .Z(O[332]) );
  AND U2225 ( .A(S), .B(n1484), .Z(n1483) );
  XOR U2226 ( .A(B[332]), .B(A[332]), .Z(n1484) );
  XOR U2227 ( .A(A[331]), .B(n1485), .Z(O[331]) );
  AND U2228 ( .A(S), .B(n1486), .Z(n1485) );
  XOR U2229 ( .A(B[331]), .B(A[331]), .Z(n1486) );
  XOR U2230 ( .A(A[330]), .B(n1487), .Z(O[330]) );
  AND U2231 ( .A(S), .B(n1488), .Z(n1487) );
  XOR U2232 ( .A(B[330]), .B(A[330]), .Z(n1488) );
  XOR U2233 ( .A(A[32]), .B(n1489), .Z(O[32]) );
  AND U2234 ( .A(S), .B(n1490), .Z(n1489) );
  XOR U2235 ( .A(B[32]), .B(A[32]), .Z(n1490) );
  XOR U2236 ( .A(A[329]), .B(n1491), .Z(O[329]) );
  AND U2237 ( .A(S), .B(n1492), .Z(n1491) );
  XOR U2238 ( .A(B[329]), .B(A[329]), .Z(n1492) );
  XOR U2239 ( .A(A[328]), .B(n1493), .Z(O[328]) );
  AND U2240 ( .A(S), .B(n1494), .Z(n1493) );
  XOR U2241 ( .A(B[328]), .B(A[328]), .Z(n1494) );
  XOR U2242 ( .A(A[327]), .B(n1495), .Z(O[327]) );
  AND U2243 ( .A(S), .B(n1496), .Z(n1495) );
  XOR U2244 ( .A(B[327]), .B(A[327]), .Z(n1496) );
  XOR U2245 ( .A(A[326]), .B(n1497), .Z(O[326]) );
  AND U2246 ( .A(S), .B(n1498), .Z(n1497) );
  XOR U2247 ( .A(B[326]), .B(A[326]), .Z(n1498) );
  XOR U2248 ( .A(A[325]), .B(n1499), .Z(O[325]) );
  AND U2249 ( .A(S), .B(n1500), .Z(n1499) );
  XOR U2250 ( .A(B[325]), .B(A[325]), .Z(n1500) );
  XOR U2251 ( .A(A[324]), .B(n1501), .Z(O[324]) );
  AND U2252 ( .A(S), .B(n1502), .Z(n1501) );
  XOR U2253 ( .A(B[324]), .B(A[324]), .Z(n1502) );
  XOR U2254 ( .A(A[323]), .B(n1503), .Z(O[323]) );
  AND U2255 ( .A(S), .B(n1504), .Z(n1503) );
  XOR U2256 ( .A(B[323]), .B(A[323]), .Z(n1504) );
  XOR U2257 ( .A(A[322]), .B(n1505), .Z(O[322]) );
  AND U2258 ( .A(S), .B(n1506), .Z(n1505) );
  XOR U2259 ( .A(B[322]), .B(A[322]), .Z(n1506) );
  XOR U2260 ( .A(A[321]), .B(n1507), .Z(O[321]) );
  AND U2261 ( .A(S), .B(n1508), .Z(n1507) );
  XOR U2262 ( .A(B[321]), .B(A[321]), .Z(n1508) );
  XOR U2263 ( .A(A[320]), .B(n1509), .Z(O[320]) );
  AND U2264 ( .A(S), .B(n1510), .Z(n1509) );
  XOR U2265 ( .A(B[320]), .B(A[320]), .Z(n1510) );
  XOR U2266 ( .A(A[31]), .B(n1511), .Z(O[31]) );
  AND U2267 ( .A(S), .B(n1512), .Z(n1511) );
  XOR U2268 ( .A(B[31]), .B(A[31]), .Z(n1512) );
  XOR U2269 ( .A(A[319]), .B(n1513), .Z(O[319]) );
  AND U2270 ( .A(S), .B(n1514), .Z(n1513) );
  XOR U2271 ( .A(B[319]), .B(A[319]), .Z(n1514) );
  XOR U2272 ( .A(A[318]), .B(n1515), .Z(O[318]) );
  AND U2273 ( .A(S), .B(n1516), .Z(n1515) );
  XOR U2274 ( .A(B[318]), .B(A[318]), .Z(n1516) );
  XOR U2275 ( .A(A[317]), .B(n1517), .Z(O[317]) );
  AND U2276 ( .A(S), .B(n1518), .Z(n1517) );
  XOR U2277 ( .A(B[317]), .B(A[317]), .Z(n1518) );
  XOR U2278 ( .A(A[316]), .B(n1519), .Z(O[316]) );
  AND U2279 ( .A(S), .B(n1520), .Z(n1519) );
  XOR U2280 ( .A(B[316]), .B(A[316]), .Z(n1520) );
  XOR U2281 ( .A(A[315]), .B(n1521), .Z(O[315]) );
  AND U2282 ( .A(S), .B(n1522), .Z(n1521) );
  XOR U2283 ( .A(B[315]), .B(A[315]), .Z(n1522) );
  XOR U2284 ( .A(A[314]), .B(n1523), .Z(O[314]) );
  AND U2285 ( .A(S), .B(n1524), .Z(n1523) );
  XOR U2286 ( .A(B[314]), .B(A[314]), .Z(n1524) );
  XOR U2287 ( .A(A[313]), .B(n1525), .Z(O[313]) );
  AND U2288 ( .A(S), .B(n1526), .Z(n1525) );
  XOR U2289 ( .A(B[313]), .B(A[313]), .Z(n1526) );
  XOR U2290 ( .A(A[312]), .B(n1527), .Z(O[312]) );
  AND U2291 ( .A(S), .B(n1528), .Z(n1527) );
  XOR U2292 ( .A(B[312]), .B(A[312]), .Z(n1528) );
  XOR U2293 ( .A(A[311]), .B(n1529), .Z(O[311]) );
  AND U2294 ( .A(S), .B(n1530), .Z(n1529) );
  XOR U2295 ( .A(B[311]), .B(A[311]), .Z(n1530) );
  XOR U2296 ( .A(A[310]), .B(n1531), .Z(O[310]) );
  AND U2297 ( .A(S), .B(n1532), .Z(n1531) );
  XOR U2298 ( .A(B[310]), .B(A[310]), .Z(n1532) );
  XOR U2299 ( .A(A[30]), .B(n1533), .Z(O[30]) );
  AND U2300 ( .A(S), .B(n1534), .Z(n1533) );
  XOR U2301 ( .A(B[30]), .B(A[30]), .Z(n1534) );
  XOR U2302 ( .A(A[309]), .B(n1535), .Z(O[309]) );
  AND U2303 ( .A(S), .B(n1536), .Z(n1535) );
  XOR U2304 ( .A(B[309]), .B(A[309]), .Z(n1536) );
  XOR U2305 ( .A(A[308]), .B(n1537), .Z(O[308]) );
  AND U2306 ( .A(S), .B(n1538), .Z(n1537) );
  XOR U2307 ( .A(B[308]), .B(A[308]), .Z(n1538) );
  XOR U2308 ( .A(A[307]), .B(n1539), .Z(O[307]) );
  AND U2309 ( .A(S), .B(n1540), .Z(n1539) );
  XOR U2310 ( .A(B[307]), .B(A[307]), .Z(n1540) );
  XOR U2311 ( .A(A[306]), .B(n1541), .Z(O[306]) );
  AND U2312 ( .A(S), .B(n1542), .Z(n1541) );
  XOR U2313 ( .A(B[306]), .B(A[306]), .Z(n1542) );
  XOR U2314 ( .A(A[305]), .B(n1543), .Z(O[305]) );
  AND U2315 ( .A(S), .B(n1544), .Z(n1543) );
  XOR U2316 ( .A(B[305]), .B(A[305]), .Z(n1544) );
  XOR U2317 ( .A(A[304]), .B(n1545), .Z(O[304]) );
  AND U2318 ( .A(S), .B(n1546), .Z(n1545) );
  XOR U2319 ( .A(B[304]), .B(A[304]), .Z(n1546) );
  XOR U2320 ( .A(A[303]), .B(n1547), .Z(O[303]) );
  AND U2321 ( .A(S), .B(n1548), .Z(n1547) );
  XOR U2322 ( .A(B[303]), .B(A[303]), .Z(n1548) );
  XOR U2323 ( .A(A[302]), .B(n1549), .Z(O[302]) );
  AND U2324 ( .A(S), .B(n1550), .Z(n1549) );
  XOR U2325 ( .A(B[302]), .B(A[302]), .Z(n1550) );
  XOR U2326 ( .A(A[301]), .B(n1551), .Z(O[301]) );
  AND U2327 ( .A(S), .B(n1552), .Z(n1551) );
  XOR U2328 ( .A(B[301]), .B(A[301]), .Z(n1552) );
  XOR U2329 ( .A(A[300]), .B(n1553), .Z(O[300]) );
  AND U2330 ( .A(S), .B(n1554), .Z(n1553) );
  XOR U2331 ( .A(B[300]), .B(A[300]), .Z(n1554) );
  XOR U2332 ( .A(A[2]), .B(n1555), .Z(O[2]) );
  AND U2333 ( .A(S), .B(n1556), .Z(n1555) );
  XOR U2334 ( .A(B[2]), .B(A[2]), .Z(n1556) );
  XOR U2335 ( .A(A[29]), .B(n1557), .Z(O[29]) );
  AND U2336 ( .A(S), .B(n1558), .Z(n1557) );
  XOR U2337 ( .A(B[29]), .B(A[29]), .Z(n1558) );
  XOR U2338 ( .A(A[299]), .B(n1559), .Z(O[299]) );
  AND U2339 ( .A(S), .B(n1560), .Z(n1559) );
  XOR U2340 ( .A(B[299]), .B(A[299]), .Z(n1560) );
  XOR U2341 ( .A(A[298]), .B(n1561), .Z(O[298]) );
  AND U2342 ( .A(S), .B(n1562), .Z(n1561) );
  XOR U2343 ( .A(B[298]), .B(A[298]), .Z(n1562) );
  XOR U2344 ( .A(A[297]), .B(n1563), .Z(O[297]) );
  AND U2345 ( .A(S), .B(n1564), .Z(n1563) );
  XOR U2346 ( .A(B[297]), .B(A[297]), .Z(n1564) );
  XOR U2347 ( .A(A[296]), .B(n1565), .Z(O[296]) );
  AND U2348 ( .A(S), .B(n1566), .Z(n1565) );
  XOR U2349 ( .A(B[296]), .B(A[296]), .Z(n1566) );
  XOR U2350 ( .A(A[295]), .B(n1567), .Z(O[295]) );
  AND U2351 ( .A(S), .B(n1568), .Z(n1567) );
  XOR U2352 ( .A(B[295]), .B(A[295]), .Z(n1568) );
  XOR U2353 ( .A(A[294]), .B(n1569), .Z(O[294]) );
  AND U2354 ( .A(S), .B(n1570), .Z(n1569) );
  XOR U2355 ( .A(B[294]), .B(A[294]), .Z(n1570) );
  XOR U2356 ( .A(A[293]), .B(n1571), .Z(O[293]) );
  AND U2357 ( .A(S), .B(n1572), .Z(n1571) );
  XOR U2358 ( .A(B[293]), .B(A[293]), .Z(n1572) );
  XOR U2359 ( .A(A[292]), .B(n1573), .Z(O[292]) );
  AND U2360 ( .A(S), .B(n1574), .Z(n1573) );
  XOR U2361 ( .A(B[292]), .B(A[292]), .Z(n1574) );
  XOR U2362 ( .A(A[291]), .B(n1575), .Z(O[291]) );
  AND U2363 ( .A(S), .B(n1576), .Z(n1575) );
  XOR U2364 ( .A(B[291]), .B(A[291]), .Z(n1576) );
  XOR U2365 ( .A(A[290]), .B(n1577), .Z(O[290]) );
  AND U2366 ( .A(S), .B(n1578), .Z(n1577) );
  XOR U2367 ( .A(B[290]), .B(A[290]), .Z(n1578) );
  XOR U2368 ( .A(A[28]), .B(n1579), .Z(O[28]) );
  AND U2369 ( .A(S), .B(n1580), .Z(n1579) );
  XOR U2370 ( .A(B[28]), .B(A[28]), .Z(n1580) );
  XOR U2371 ( .A(A[289]), .B(n1581), .Z(O[289]) );
  AND U2372 ( .A(S), .B(n1582), .Z(n1581) );
  XOR U2373 ( .A(B[289]), .B(A[289]), .Z(n1582) );
  XOR U2374 ( .A(A[288]), .B(n1583), .Z(O[288]) );
  AND U2375 ( .A(S), .B(n1584), .Z(n1583) );
  XOR U2376 ( .A(B[288]), .B(A[288]), .Z(n1584) );
  XOR U2377 ( .A(A[287]), .B(n1585), .Z(O[287]) );
  AND U2378 ( .A(S), .B(n1586), .Z(n1585) );
  XOR U2379 ( .A(B[287]), .B(A[287]), .Z(n1586) );
  XOR U2380 ( .A(A[286]), .B(n1587), .Z(O[286]) );
  AND U2381 ( .A(S), .B(n1588), .Z(n1587) );
  XOR U2382 ( .A(B[286]), .B(A[286]), .Z(n1588) );
  XOR U2383 ( .A(A[285]), .B(n1589), .Z(O[285]) );
  AND U2384 ( .A(S), .B(n1590), .Z(n1589) );
  XOR U2385 ( .A(B[285]), .B(A[285]), .Z(n1590) );
  XOR U2386 ( .A(A[284]), .B(n1591), .Z(O[284]) );
  AND U2387 ( .A(S), .B(n1592), .Z(n1591) );
  XOR U2388 ( .A(B[284]), .B(A[284]), .Z(n1592) );
  XOR U2389 ( .A(A[283]), .B(n1593), .Z(O[283]) );
  AND U2390 ( .A(S), .B(n1594), .Z(n1593) );
  XOR U2391 ( .A(B[283]), .B(A[283]), .Z(n1594) );
  XOR U2392 ( .A(A[282]), .B(n1595), .Z(O[282]) );
  AND U2393 ( .A(S), .B(n1596), .Z(n1595) );
  XOR U2394 ( .A(B[282]), .B(A[282]), .Z(n1596) );
  XOR U2395 ( .A(A[281]), .B(n1597), .Z(O[281]) );
  AND U2396 ( .A(S), .B(n1598), .Z(n1597) );
  XOR U2397 ( .A(B[281]), .B(A[281]), .Z(n1598) );
  XOR U2398 ( .A(A[280]), .B(n1599), .Z(O[280]) );
  AND U2399 ( .A(S), .B(n1600), .Z(n1599) );
  XOR U2400 ( .A(B[280]), .B(A[280]), .Z(n1600) );
  XOR U2401 ( .A(A[27]), .B(n1601), .Z(O[27]) );
  AND U2402 ( .A(S), .B(n1602), .Z(n1601) );
  XOR U2403 ( .A(B[27]), .B(A[27]), .Z(n1602) );
  XOR U2404 ( .A(A[279]), .B(n1603), .Z(O[279]) );
  AND U2405 ( .A(S), .B(n1604), .Z(n1603) );
  XOR U2406 ( .A(B[279]), .B(A[279]), .Z(n1604) );
  XOR U2407 ( .A(A[278]), .B(n1605), .Z(O[278]) );
  AND U2408 ( .A(S), .B(n1606), .Z(n1605) );
  XOR U2409 ( .A(B[278]), .B(A[278]), .Z(n1606) );
  XOR U2410 ( .A(A[277]), .B(n1607), .Z(O[277]) );
  AND U2411 ( .A(S), .B(n1608), .Z(n1607) );
  XOR U2412 ( .A(B[277]), .B(A[277]), .Z(n1608) );
  XOR U2413 ( .A(A[276]), .B(n1609), .Z(O[276]) );
  AND U2414 ( .A(S), .B(n1610), .Z(n1609) );
  XOR U2415 ( .A(B[276]), .B(A[276]), .Z(n1610) );
  XOR U2416 ( .A(A[275]), .B(n1611), .Z(O[275]) );
  AND U2417 ( .A(S), .B(n1612), .Z(n1611) );
  XOR U2418 ( .A(B[275]), .B(A[275]), .Z(n1612) );
  XOR U2419 ( .A(A[274]), .B(n1613), .Z(O[274]) );
  AND U2420 ( .A(S), .B(n1614), .Z(n1613) );
  XOR U2421 ( .A(B[274]), .B(A[274]), .Z(n1614) );
  XOR U2422 ( .A(A[273]), .B(n1615), .Z(O[273]) );
  AND U2423 ( .A(S), .B(n1616), .Z(n1615) );
  XOR U2424 ( .A(B[273]), .B(A[273]), .Z(n1616) );
  XOR U2425 ( .A(A[272]), .B(n1617), .Z(O[272]) );
  AND U2426 ( .A(S), .B(n1618), .Z(n1617) );
  XOR U2427 ( .A(B[272]), .B(A[272]), .Z(n1618) );
  XOR U2428 ( .A(A[271]), .B(n1619), .Z(O[271]) );
  AND U2429 ( .A(S), .B(n1620), .Z(n1619) );
  XOR U2430 ( .A(B[271]), .B(A[271]), .Z(n1620) );
  XOR U2431 ( .A(A[270]), .B(n1621), .Z(O[270]) );
  AND U2432 ( .A(S), .B(n1622), .Z(n1621) );
  XOR U2433 ( .A(B[270]), .B(A[270]), .Z(n1622) );
  XOR U2434 ( .A(A[26]), .B(n1623), .Z(O[26]) );
  AND U2435 ( .A(S), .B(n1624), .Z(n1623) );
  XOR U2436 ( .A(B[26]), .B(A[26]), .Z(n1624) );
  XOR U2437 ( .A(A[269]), .B(n1625), .Z(O[269]) );
  AND U2438 ( .A(S), .B(n1626), .Z(n1625) );
  XOR U2439 ( .A(B[269]), .B(A[269]), .Z(n1626) );
  XOR U2440 ( .A(A[268]), .B(n1627), .Z(O[268]) );
  AND U2441 ( .A(S), .B(n1628), .Z(n1627) );
  XOR U2442 ( .A(B[268]), .B(A[268]), .Z(n1628) );
  XOR U2443 ( .A(A[267]), .B(n1629), .Z(O[267]) );
  AND U2444 ( .A(S), .B(n1630), .Z(n1629) );
  XOR U2445 ( .A(B[267]), .B(A[267]), .Z(n1630) );
  XOR U2446 ( .A(A[266]), .B(n1631), .Z(O[266]) );
  AND U2447 ( .A(S), .B(n1632), .Z(n1631) );
  XOR U2448 ( .A(B[266]), .B(A[266]), .Z(n1632) );
  XOR U2449 ( .A(A[265]), .B(n1633), .Z(O[265]) );
  AND U2450 ( .A(S), .B(n1634), .Z(n1633) );
  XOR U2451 ( .A(B[265]), .B(A[265]), .Z(n1634) );
  XOR U2452 ( .A(A[264]), .B(n1635), .Z(O[264]) );
  AND U2453 ( .A(S), .B(n1636), .Z(n1635) );
  XOR U2454 ( .A(B[264]), .B(A[264]), .Z(n1636) );
  XOR U2455 ( .A(A[263]), .B(n1637), .Z(O[263]) );
  AND U2456 ( .A(S), .B(n1638), .Z(n1637) );
  XOR U2457 ( .A(B[263]), .B(A[263]), .Z(n1638) );
  XOR U2458 ( .A(A[262]), .B(n1639), .Z(O[262]) );
  AND U2459 ( .A(S), .B(n1640), .Z(n1639) );
  XOR U2460 ( .A(B[262]), .B(A[262]), .Z(n1640) );
  XOR U2461 ( .A(A[261]), .B(n1641), .Z(O[261]) );
  AND U2462 ( .A(S), .B(n1642), .Z(n1641) );
  XOR U2463 ( .A(B[261]), .B(A[261]), .Z(n1642) );
  XOR U2464 ( .A(A[260]), .B(n1643), .Z(O[260]) );
  AND U2465 ( .A(S), .B(n1644), .Z(n1643) );
  XOR U2466 ( .A(B[260]), .B(A[260]), .Z(n1644) );
  XOR U2467 ( .A(A[25]), .B(n1645), .Z(O[25]) );
  AND U2468 ( .A(S), .B(n1646), .Z(n1645) );
  XOR U2469 ( .A(B[25]), .B(A[25]), .Z(n1646) );
  XOR U2470 ( .A(A[259]), .B(n1647), .Z(O[259]) );
  AND U2471 ( .A(S), .B(n1648), .Z(n1647) );
  XOR U2472 ( .A(B[259]), .B(A[259]), .Z(n1648) );
  XOR U2473 ( .A(A[258]), .B(n1649), .Z(O[258]) );
  AND U2474 ( .A(S), .B(n1650), .Z(n1649) );
  XOR U2475 ( .A(B[258]), .B(A[258]), .Z(n1650) );
  XOR U2476 ( .A(A[257]), .B(n1651), .Z(O[257]) );
  AND U2477 ( .A(S), .B(n1652), .Z(n1651) );
  XOR U2478 ( .A(B[257]), .B(A[257]), .Z(n1652) );
  XOR U2479 ( .A(A[256]), .B(n1653), .Z(O[256]) );
  AND U2480 ( .A(S), .B(n1654), .Z(n1653) );
  XOR U2481 ( .A(B[256]), .B(A[256]), .Z(n1654) );
  XOR U2482 ( .A(A[255]), .B(n1655), .Z(O[255]) );
  AND U2483 ( .A(S), .B(n1656), .Z(n1655) );
  XOR U2484 ( .A(B[255]), .B(A[255]), .Z(n1656) );
  XOR U2485 ( .A(A[254]), .B(n1657), .Z(O[254]) );
  AND U2486 ( .A(S), .B(n1658), .Z(n1657) );
  XOR U2487 ( .A(B[254]), .B(A[254]), .Z(n1658) );
  XOR U2488 ( .A(A[253]), .B(n1659), .Z(O[253]) );
  AND U2489 ( .A(S), .B(n1660), .Z(n1659) );
  XOR U2490 ( .A(B[253]), .B(A[253]), .Z(n1660) );
  XOR U2491 ( .A(A[252]), .B(n1661), .Z(O[252]) );
  AND U2492 ( .A(S), .B(n1662), .Z(n1661) );
  XOR U2493 ( .A(B[252]), .B(A[252]), .Z(n1662) );
  XOR U2494 ( .A(A[251]), .B(n1663), .Z(O[251]) );
  AND U2495 ( .A(S), .B(n1664), .Z(n1663) );
  XOR U2496 ( .A(B[251]), .B(A[251]), .Z(n1664) );
  XOR U2497 ( .A(A[250]), .B(n1665), .Z(O[250]) );
  AND U2498 ( .A(S), .B(n1666), .Z(n1665) );
  XOR U2499 ( .A(B[250]), .B(A[250]), .Z(n1666) );
  XOR U2500 ( .A(A[24]), .B(n1667), .Z(O[24]) );
  AND U2501 ( .A(S), .B(n1668), .Z(n1667) );
  XOR U2502 ( .A(B[24]), .B(A[24]), .Z(n1668) );
  XOR U2503 ( .A(A[249]), .B(n1669), .Z(O[249]) );
  AND U2504 ( .A(S), .B(n1670), .Z(n1669) );
  XOR U2505 ( .A(B[249]), .B(A[249]), .Z(n1670) );
  XOR U2506 ( .A(A[248]), .B(n1671), .Z(O[248]) );
  AND U2507 ( .A(S), .B(n1672), .Z(n1671) );
  XOR U2508 ( .A(B[248]), .B(A[248]), .Z(n1672) );
  XOR U2509 ( .A(A[247]), .B(n1673), .Z(O[247]) );
  AND U2510 ( .A(S), .B(n1674), .Z(n1673) );
  XOR U2511 ( .A(B[247]), .B(A[247]), .Z(n1674) );
  XOR U2512 ( .A(A[246]), .B(n1675), .Z(O[246]) );
  AND U2513 ( .A(S), .B(n1676), .Z(n1675) );
  XOR U2514 ( .A(B[246]), .B(A[246]), .Z(n1676) );
  XOR U2515 ( .A(A[245]), .B(n1677), .Z(O[245]) );
  AND U2516 ( .A(S), .B(n1678), .Z(n1677) );
  XOR U2517 ( .A(B[245]), .B(A[245]), .Z(n1678) );
  XOR U2518 ( .A(A[244]), .B(n1679), .Z(O[244]) );
  AND U2519 ( .A(S), .B(n1680), .Z(n1679) );
  XOR U2520 ( .A(B[244]), .B(A[244]), .Z(n1680) );
  XOR U2521 ( .A(A[243]), .B(n1681), .Z(O[243]) );
  AND U2522 ( .A(S), .B(n1682), .Z(n1681) );
  XOR U2523 ( .A(B[243]), .B(A[243]), .Z(n1682) );
  XOR U2524 ( .A(A[242]), .B(n1683), .Z(O[242]) );
  AND U2525 ( .A(S), .B(n1684), .Z(n1683) );
  XOR U2526 ( .A(B[242]), .B(A[242]), .Z(n1684) );
  XOR U2527 ( .A(A[241]), .B(n1685), .Z(O[241]) );
  AND U2528 ( .A(S), .B(n1686), .Z(n1685) );
  XOR U2529 ( .A(B[241]), .B(A[241]), .Z(n1686) );
  XOR U2530 ( .A(A[240]), .B(n1687), .Z(O[240]) );
  AND U2531 ( .A(S), .B(n1688), .Z(n1687) );
  XOR U2532 ( .A(B[240]), .B(A[240]), .Z(n1688) );
  XOR U2533 ( .A(A[23]), .B(n1689), .Z(O[23]) );
  AND U2534 ( .A(S), .B(n1690), .Z(n1689) );
  XOR U2535 ( .A(B[23]), .B(A[23]), .Z(n1690) );
  XOR U2536 ( .A(A[239]), .B(n1691), .Z(O[239]) );
  AND U2537 ( .A(S), .B(n1692), .Z(n1691) );
  XOR U2538 ( .A(B[239]), .B(A[239]), .Z(n1692) );
  XOR U2539 ( .A(A[238]), .B(n1693), .Z(O[238]) );
  AND U2540 ( .A(S), .B(n1694), .Z(n1693) );
  XOR U2541 ( .A(B[238]), .B(A[238]), .Z(n1694) );
  XOR U2542 ( .A(A[237]), .B(n1695), .Z(O[237]) );
  AND U2543 ( .A(S), .B(n1696), .Z(n1695) );
  XOR U2544 ( .A(B[237]), .B(A[237]), .Z(n1696) );
  XOR U2545 ( .A(A[236]), .B(n1697), .Z(O[236]) );
  AND U2546 ( .A(S), .B(n1698), .Z(n1697) );
  XOR U2547 ( .A(B[236]), .B(A[236]), .Z(n1698) );
  XOR U2548 ( .A(A[235]), .B(n1699), .Z(O[235]) );
  AND U2549 ( .A(S), .B(n1700), .Z(n1699) );
  XOR U2550 ( .A(B[235]), .B(A[235]), .Z(n1700) );
  XOR U2551 ( .A(A[234]), .B(n1701), .Z(O[234]) );
  AND U2552 ( .A(S), .B(n1702), .Z(n1701) );
  XOR U2553 ( .A(B[234]), .B(A[234]), .Z(n1702) );
  XOR U2554 ( .A(A[233]), .B(n1703), .Z(O[233]) );
  AND U2555 ( .A(S), .B(n1704), .Z(n1703) );
  XOR U2556 ( .A(B[233]), .B(A[233]), .Z(n1704) );
  XOR U2557 ( .A(A[232]), .B(n1705), .Z(O[232]) );
  AND U2558 ( .A(S), .B(n1706), .Z(n1705) );
  XOR U2559 ( .A(B[232]), .B(A[232]), .Z(n1706) );
  XOR U2560 ( .A(A[231]), .B(n1707), .Z(O[231]) );
  AND U2561 ( .A(S), .B(n1708), .Z(n1707) );
  XOR U2562 ( .A(B[231]), .B(A[231]), .Z(n1708) );
  XOR U2563 ( .A(A[230]), .B(n1709), .Z(O[230]) );
  AND U2564 ( .A(S), .B(n1710), .Z(n1709) );
  XOR U2565 ( .A(B[230]), .B(A[230]), .Z(n1710) );
  XOR U2566 ( .A(A[22]), .B(n1711), .Z(O[22]) );
  AND U2567 ( .A(S), .B(n1712), .Z(n1711) );
  XOR U2568 ( .A(B[22]), .B(A[22]), .Z(n1712) );
  XOR U2569 ( .A(A[229]), .B(n1713), .Z(O[229]) );
  AND U2570 ( .A(S), .B(n1714), .Z(n1713) );
  XOR U2571 ( .A(B[229]), .B(A[229]), .Z(n1714) );
  XOR U2572 ( .A(A[228]), .B(n1715), .Z(O[228]) );
  AND U2573 ( .A(S), .B(n1716), .Z(n1715) );
  XOR U2574 ( .A(B[228]), .B(A[228]), .Z(n1716) );
  XOR U2575 ( .A(A[227]), .B(n1717), .Z(O[227]) );
  AND U2576 ( .A(S), .B(n1718), .Z(n1717) );
  XOR U2577 ( .A(B[227]), .B(A[227]), .Z(n1718) );
  XOR U2578 ( .A(A[226]), .B(n1719), .Z(O[226]) );
  AND U2579 ( .A(S), .B(n1720), .Z(n1719) );
  XOR U2580 ( .A(B[226]), .B(A[226]), .Z(n1720) );
  XOR U2581 ( .A(A[225]), .B(n1721), .Z(O[225]) );
  AND U2582 ( .A(S), .B(n1722), .Z(n1721) );
  XOR U2583 ( .A(B[225]), .B(A[225]), .Z(n1722) );
  XOR U2584 ( .A(A[224]), .B(n1723), .Z(O[224]) );
  AND U2585 ( .A(S), .B(n1724), .Z(n1723) );
  XOR U2586 ( .A(B[224]), .B(A[224]), .Z(n1724) );
  XOR U2587 ( .A(A[223]), .B(n1725), .Z(O[223]) );
  AND U2588 ( .A(S), .B(n1726), .Z(n1725) );
  XOR U2589 ( .A(B[223]), .B(A[223]), .Z(n1726) );
  XOR U2590 ( .A(A[222]), .B(n1727), .Z(O[222]) );
  AND U2591 ( .A(S), .B(n1728), .Z(n1727) );
  XOR U2592 ( .A(B[222]), .B(A[222]), .Z(n1728) );
  XOR U2593 ( .A(A[221]), .B(n1729), .Z(O[221]) );
  AND U2594 ( .A(S), .B(n1730), .Z(n1729) );
  XOR U2595 ( .A(B[221]), .B(A[221]), .Z(n1730) );
  XOR U2596 ( .A(A[220]), .B(n1731), .Z(O[220]) );
  AND U2597 ( .A(S), .B(n1732), .Z(n1731) );
  XOR U2598 ( .A(B[220]), .B(A[220]), .Z(n1732) );
  XOR U2599 ( .A(A[21]), .B(n1733), .Z(O[21]) );
  AND U2600 ( .A(S), .B(n1734), .Z(n1733) );
  XOR U2601 ( .A(B[21]), .B(A[21]), .Z(n1734) );
  XOR U2602 ( .A(A[219]), .B(n1735), .Z(O[219]) );
  AND U2603 ( .A(S), .B(n1736), .Z(n1735) );
  XOR U2604 ( .A(B[219]), .B(A[219]), .Z(n1736) );
  XOR U2605 ( .A(A[218]), .B(n1737), .Z(O[218]) );
  AND U2606 ( .A(S), .B(n1738), .Z(n1737) );
  XOR U2607 ( .A(B[218]), .B(A[218]), .Z(n1738) );
  XOR U2608 ( .A(A[217]), .B(n1739), .Z(O[217]) );
  AND U2609 ( .A(S), .B(n1740), .Z(n1739) );
  XOR U2610 ( .A(B[217]), .B(A[217]), .Z(n1740) );
  XOR U2611 ( .A(A[216]), .B(n1741), .Z(O[216]) );
  AND U2612 ( .A(S), .B(n1742), .Z(n1741) );
  XOR U2613 ( .A(B[216]), .B(A[216]), .Z(n1742) );
  XOR U2614 ( .A(A[215]), .B(n1743), .Z(O[215]) );
  AND U2615 ( .A(S), .B(n1744), .Z(n1743) );
  XOR U2616 ( .A(B[215]), .B(A[215]), .Z(n1744) );
  XOR U2617 ( .A(A[214]), .B(n1745), .Z(O[214]) );
  AND U2618 ( .A(S), .B(n1746), .Z(n1745) );
  XOR U2619 ( .A(B[214]), .B(A[214]), .Z(n1746) );
  XOR U2620 ( .A(A[213]), .B(n1747), .Z(O[213]) );
  AND U2621 ( .A(S), .B(n1748), .Z(n1747) );
  XOR U2622 ( .A(B[213]), .B(A[213]), .Z(n1748) );
  XOR U2623 ( .A(A[212]), .B(n1749), .Z(O[212]) );
  AND U2624 ( .A(S), .B(n1750), .Z(n1749) );
  XOR U2625 ( .A(B[212]), .B(A[212]), .Z(n1750) );
  XOR U2626 ( .A(A[211]), .B(n1751), .Z(O[211]) );
  AND U2627 ( .A(S), .B(n1752), .Z(n1751) );
  XOR U2628 ( .A(B[211]), .B(A[211]), .Z(n1752) );
  XOR U2629 ( .A(A[210]), .B(n1753), .Z(O[210]) );
  AND U2630 ( .A(S), .B(n1754), .Z(n1753) );
  XOR U2631 ( .A(B[210]), .B(A[210]), .Z(n1754) );
  XOR U2632 ( .A(A[20]), .B(n1755), .Z(O[20]) );
  AND U2633 ( .A(S), .B(n1756), .Z(n1755) );
  XOR U2634 ( .A(B[20]), .B(A[20]), .Z(n1756) );
  XOR U2635 ( .A(A[209]), .B(n1757), .Z(O[209]) );
  AND U2636 ( .A(S), .B(n1758), .Z(n1757) );
  XOR U2637 ( .A(B[209]), .B(A[209]), .Z(n1758) );
  XOR U2638 ( .A(A[208]), .B(n1759), .Z(O[208]) );
  AND U2639 ( .A(S), .B(n1760), .Z(n1759) );
  XOR U2640 ( .A(B[208]), .B(A[208]), .Z(n1760) );
  XOR U2641 ( .A(A[207]), .B(n1761), .Z(O[207]) );
  AND U2642 ( .A(S), .B(n1762), .Z(n1761) );
  XOR U2643 ( .A(B[207]), .B(A[207]), .Z(n1762) );
  XOR U2644 ( .A(A[206]), .B(n1763), .Z(O[206]) );
  AND U2645 ( .A(S), .B(n1764), .Z(n1763) );
  XOR U2646 ( .A(B[206]), .B(A[206]), .Z(n1764) );
  XOR U2647 ( .A(A[205]), .B(n1765), .Z(O[205]) );
  AND U2648 ( .A(S), .B(n1766), .Z(n1765) );
  XOR U2649 ( .A(B[205]), .B(A[205]), .Z(n1766) );
  XOR U2650 ( .A(A[204]), .B(n1767), .Z(O[204]) );
  AND U2651 ( .A(S), .B(n1768), .Z(n1767) );
  XOR U2652 ( .A(B[204]), .B(A[204]), .Z(n1768) );
  XOR U2653 ( .A(A[203]), .B(n1769), .Z(O[203]) );
  AND U2654 ( .A(S), .B(n1770), .Z(n1769) );
  XOR U2655 ( .A(B[203]), .B(A[203]), .Z(n1770) );
  XOR U2656 ( .A(A[202]), .B(n1771), .Z(O[202]) );
  AND U2657 ( .A(S), .B(n1772), .Z(n1771) );
  XOR U2658 ( .A(B[202]), .B(A[202]), .Z(n1772) );
  XOR U2659 ( .A(A[201]), .B(n1773), .Z(O[201]) );
  AND U2660 ( .A(S), .B(n1774), .Z(n1773) );
  XOR U2661 ( .A(B[201]), .B(A[201]), .Z(n1774) );
  XOR U2662 ( .A(A[200]), .B(n1775), .Z(O[200]) );
  AND U2663 ( .A(S), .B(n1776), .Z(n1775) );
  XOR U2664 ( .A(B[200]), .B(A[200]), .Z(n1776) );
  XOR U2665 ( .A(A[1]), .B(n1777), .Z(O[1]) );
  AND U2666 ( .A(S), .B(n1778), .Z(n1777) );
  XOR U2667 ( .A(B[1]), .B(A[1]), .Z(n1778) );
  XOR U2668 ( .A(A[19]), .B(n1779), .Z(O[19]) );
  AND U2669 ( .A(S), .B(n1780), .Z(n1779) );
  XOR U2670 ( .A(B[19]), .B(A[19]), .Z(n1780) );
  XOR U2671 ( .A(A[199]), .B(n1781), .Z(O[199]) );
  AND U2672 ( .A(S), .B(n1782), .Z(n1781) );
  XOR U2673 ( .A(B[199]), .B(A[199]), .Z(n1782) );
  XOR U2674 ( .A(A[198]), .B(n1783), .Z(O[198]) );
  AND U2675 ( .A(S), .B(n1784), .Z(n1783) );
  XOR U2676 ( .A(B[198]), .B(A[198]), .Z(n1784) );
  XOR U2677 ( .A(A[197]), .B(n1785), .Z(O[197]) );
  AND U2678 ( .A(S), .B(n1786), .Z(n1785) );
  XOR U2679 ( .A(B[197]), .B(A[197]), .Z(n1786) );
  XOR U2680 ( .A(A[196]), .B(n1787), .Z(O[196]) );
  AND U2681 ( .A(S), .B(n1788), .Z(n1787) );
  XOR U2682 ( .A(B[196]), .B(A[196]), .Z(n1788) );
  XOR U2683 ( .A(A[195]), .B(n1789), .Z(O[195]) );
  AND U2684 ( .A(S), .B(n1790), .Z(n1789) );
  XOR U2685 ( .A(B[195]), .B(A[195]), .Z(n1790) );
  XOR U2686 ( .A(A[194]), .B(n1791), .Z(O[194]) );
  AND U2687 ( .A(S), .B(n1792), .Z(n1791) );
  XOR U2688 ( .A(B[194]), .B(A[194]), .Z(n1792) );
  XOR U2689 ( .A(A[193]), .B(n1793), .Z(O[193]) );
  AND U2690 ( .A(S), .B(n1794), .Z(n1793) );
  XOR U2691 ( .A(B[193]), .B(A[193]), .Z(n1794) );
  XOR U2692 ( .A(A[192]), .B(n1795), .Z(O[192]) );
  AND U2693 ( .A(S), .B(n1796), .Z(n1795) );
  XOR U2694 ( .A(B[192]), .B(A[192]), .Z(n1796) );
  XOR U2695 ( .A(A[191]), .B(n1797), .Z(O[191]) );
  AND U2696 ( .A(S), .B(n1798), .Z(n1797) );
  XOR U2697 ( .A(B[191]), .B(A[191]), .Z(n1798) );
  XOR U2698 ( .A(A[190]), .B(n1799), .Z(O[190]) );
  AND U2699 ( .A(S), .B(n1800), .Z(n1799) );
  XOR U2700 ( .A(B[190]), .B(A[190]), .Z(n1800) );
  XOR U2701 ( .A(A[18]), .B(n1801), .Z(O[18]) );
  AND U2702 ( .A(S), .B(n1802), .Z(n1801) );
  XOR U2703 ( .A(B[18]), .B(A[18]), .Z(n1802) );
  XOR U2704 ( .A(A[189]), .B(n1803), .Z(O[189]) );
  AND U2705 ( .A(S), .B(n1804), .Z(n1803) );
  XOR U2706 ( .A(B[189]), .B(A[189]), .Z(n1804) );
  XOR U2707 ( .A(A[188]), .B(n1805), .Z(O[188]) );
  AND U2708 ( .A(S), .B(n1806), .Z(n1805) );
  XOR U2709 ( .A(B[188]), .B(A[188]), .Z(n1806) );
  XOR U2710 ( .A(A[187]), .B(n1807), .Z(O[187]) );
  AND U2711 ( .A(S), .B(n1808), .Z(n1807) );
  XOR U2712 ( .A(B[187]), .B(A[187]), .Z(n1808) );
  XOR U2713 ( .A(A[186]), .B(n1809), .Z(O[186]) );
  AND U2714 ( .A(S), .B(n1810), .Z(n1809) );
  XOR U2715 ( .A(B[186]), .B(A[186]), .Z(n1810) );
  XOR U2716 ( .A(A[185]), .B(n1811), .Z(O[185]) );
  AND U2717 ( .A(S), .B(n1812), .Z(n1811) );
  XOR U2718 ( .A(B[185]), .B(A[185]), .Z(n1812) );
  XOR U2719 ( .A(A[184]), .B(n1813), .Z(O[184]) );
  AND U2720 ( .A(S), .B(n1814), .Z(n1813) );
  XOR U2721 ( .A(B[184]), .B(A[184]), .Z(n1814) );
  XOR U2722 ( .A(A[183]), .B(n1815), .Z(O[183]) );
  AND U2723 ( .A(S), .B(n1816), .Z(n1815) );
  XOR U2724 ( .A(B[183]), .B(A[183]), .Z(n1816) );
  XOR U2725 ( .A(A[182]), .B(n1817), .Z(O[182]) );
  AND U2726 ( .A(S), .B(n1818), .Z(n1817) );
  XOR U2727 ( .A(B[182]), .B(A[182]), .Z(n1818) );
  XOR U2728 ( .A(A[181]), .B(n1819), .Z(O[181]) );
  AND U2729 ( .A(S), .B(n1820), .Z(n1819) );
  XOR U2730 ( .A(B[181]), .B(A[181]), .Z(n1820) );
  XOR U2731 ( .A(A[180]), .B(n1821), .Z(O[180]) );
  AND U2732 ( .A(S), .B(n1822), .Z(n1821) );
  XOR U2733 ( .A(B[180]), .B(A[180]), .Z(n1822) );
  XOR U2734 ( .A(A[17]), .B(n1823), .Z(O[17]) );
  AND U2735 ( .A(S), .B(n1824), .Z(n1823) );
  XOR U2736 ( .A(B[17]), .B(A[17]), .Z(n1824) );
  XOR U2737 ( .A(A[179]), .B(n1825), .Z(O[179]) );
  AND U2738 ( .A(S), .B(n1826), .Z(n1825) );
  XOR U2739 ( .A(B[179]), .B(A[179]), .Z(n1826) );
  XOR U2740 ( .A(A[178]), .B(n1827), .Z(O[178]) );
  AND U2741 ( .A(S), .B(n1828), .Z(n1827) );
  XOR U2742 ( .A(B[178]), .B(A[178]), .Z(n1828) );
  XOR U2743 ( .A(A[177]), .B(n1829), .Z(O[177]) );
  AND U2744 ( .A(S), .B(n1830), .Z(n1829) );
  XOR U2745 ( .A(B[177]), .B(A[177]), .Z(n1830) );
  XOR U2746 ( .A(A[176]), .B(n1831), .Z(O[176]) );
  AND U2747 ( .A(S), .B(n1832), .Z(n1831) );
  XOR U2748 ( .A(B[176]), .B(A[176]), .Z(n1832) );
  XOR U2749 ( .A(A[175]), .B(n1833), .Z(O[175]) );
  AND U2750 ( .A(S), .B(n1834), .Z(n1833) );
  XOR U2751 ( .A(B[175]), .B(A[175]), .Z(n1834) );
  XOR U2752 ( .A(A[174]), .B(n1835), .Z(O[174]) );
  AND U2753 ( .A(S), .B(n1836), .Z(n1835) );
  XOR U2754 ( .A(B[174]), .B(A[174]), .Z(n1836) );
  XOR U2755 ( .A(A[173]), .B(n1837), .Z(O[173]) );
  AND U2756 ( .A(S), .B(n1838), .Z(n1837) );
  XOR U2757 ( .A(B[173]), .B(A[173]), .Z(n1838) );
  XOR U2758 ( .A(A[172]), .B(n1839), .Z(O[172]) );
  AND U2759 ( .A(S), .B(n1840), .Z(n1839) );
  XOR U2760 ( .A(B[172]), .B(A[172]), .Z(n1840) );
  XOR U2761 ( .A(A[171]), .B(n1841), .Z(O[171]) );
  AND U2762 ( .A(S), .B(n1842), .Z(n1841) );
  XOR U2763 ( .A(B[171]), .B(A[171]), .Z(n1842) );
  XOR U2764 ( .A(A[170]), .B(n1843), .Z(O[170]) );
  AND U2765 ( .A(S), .B(n1844), .Z(n1843) );
  XOR U2766 ( .A(B[170]), .B(A[170]), .Z(n1844) );
  XOR U2767 ( .A(A[16]), .B(n1845), .Z(O[16]) );
  AND U2768 ( .A(S), .B(n1846), .Z(n1845) );
  XOR U2769 ( .A(B[16]), .B(A[16]), .Z(n1846) );
  XOR U2770 ( .A(A[169]), .B(n1847), .Z(O[169]) );
  AND U2771 ( .A(S), .B(n1848), .Z(n1847) );
  XOR U2772 ( .A(B[169]), .B(A[169]), .Z(n1848) );
  XOR U2773 ( .A(A[168]), .B(n1849), .Z(O[168]) );
  AND U2774 ( .A(S), .B(n1850), .Z(n1849) );
  XOR U2775 ( .A(B[168]), .B(A[168]), .Z(n1850) );
  XOR U2776 ( .A(A[167]), .B(n1851), .Z(O[167]) );
  AND U2777 ( .A(S), .B(n1852), .Z(n1851) );
  XOR U2778 ( .A(B[167]), .B(A[167]), .Z(n1852) );
  XOR U2779 ( .A(A[166]), .B(n1853), .Z(O[166]) );
  AND U2780 ( .A(S), .B(n1854), .Z(n1853) );
  XOR U2781 ( .A(B[166]), .B(A[166]), .Z(n1854) );
  XOR U2782 ( .A(A[165]), .B(n1855), .Z(O[165]) );
  AND U2783 ( .A(S), .B(n1856), .Z(n1855) );
  XOR U2784 ( .A(B[165]), .B(A[165]), .Z(n1856) );
  XOR U2785 ( .A(A[164]), .B(n1857), .Z(O[164]) );
  AND U2786 ( .A(S), .B(n1858), .Z(n1857) );
  XOR U2787 ( .A(B[164]), .B(A[164]), .Z(n1858) );
  XOR U2788 ( .A(A[163]), .B(n1859), .Z(O[163]) );
  AND U2789 ( .A(S), .B(n1860), .Z(n1859) );
  XOR U2790 ( .A(B[163]), .B(A[163]), .Z(n1860) );
  XOR U2791 ( .A(A[162]), .B(n1861), .Z(O[162]) );
  AND U2792 ( .A(S), .B(n1862), .Z(n1861) );
  XOR U2793 ( .A(B[162]), .B(A[162]), .Z(n1862) );
  XOR U2794 ( .A(A[161]), .B(n1863), .Z(O[161]) );
  AND U2795 ( .A(S), .B(n1864), .Z(n1863) );
  XOR U2796 ( .A(B[161]), .B(A[161]), .Z(n1864) );
  XOR U2797 ( .A(A[160]), .B(n1865), .Z(O[160]) );
  AND U2798 ( .A(S), .B(n1866), .Z(n1865) );
  XOR U2799 ( .A(B[160]), .B(A[160]), .Z(n1866) );
  XOR U2800 ( .A(A[15]), .B(n1867), .Z(O[15]) );
  AND U2801 ( .A(S), .B(n1868), .Z(n1867) );
  XOR U2802 ( .A(B[15]), .B(A[15]), .Z(n1868) );
  XOR U2803 ( .A(A[159]), .B(n1869), .Z(O[159]) );
  AND U2804 ( .A(S), .B(n1870), .Z(n1869) );
  XOR U2805 ( .A(B[159]), .B(A[159]), .Z(n1870) );
  XOR U2806 ( .A(A[158]), .B(n1871), .Z(O[158]) );
  AND U2807 ( .A(S), .B(n1872), .Z(n1871) );
  XOR U2808 ( .A(B[158]), .B(A[158]), .Z(n1872) );
  XOR U2809 ( .A(A[157]), .B(n1873), .Z(O[157]) );
  AND U2810 ( .A(S), .B(n1874), .Z(n1873) );
  XOR U2811 ( .A(B[157]), .B(A[157]), .Z(n1874) );
  XOR U2812 ( .A(A[156]), .B(n1875), .Z(O[156]) );
  AND U2813 ( .A(S), .B(n1876), .Z(n1875) );
  XOR U2814 ( .A(B[156]), .B(A[156]), .Z(n1876) );
  XOR U2815 ( .A(A[155]), .B(n1877), .Z(O[155]) );
  AND U2816 ( .A(S), .B(n1878), .Z(n1877) );
  XOR U2817 ( .A(B[155]), .B(A[155]), .Z(n1878) );
  XOR U2818 ( .A(A[154]), .B(n1879), .Z(O[154]) );
  AND U2819 ( .A(S), .B(n1880), .Z(n1879) );
  XOR U2820 ( .A(B[154]), .B(A[154]), .Z(n1880) );
  XOR U2821 ( .A(A[153]), .B(n1881), .Z(O[153]) );
  AND U2822 ( .A(S), .B(n1882), .Z(n1881) );
  XOR U2823 ( .A(B[153]), .B(A[153]), .Z(n1882) );
  XOR U2824 ( .A(A[152]), .B(n1883), .Z(O[152]) );
  AND U2825 ( .A(S), .B(n1884), .Z(n1883) );
  XOR U2826 ( .A(B[152]), .B(A[152]), .Z(n1884) );
  XOR U2827 ( .A(A[151]), .B(n1885), .Z(O[151]) );
  AND U2828 ( .A(S), .B(n1886), .Z(n1885) );
  XOR U2829 ( .A(B[151]), .B(A[151]), .Z(n1886) );
  XOR U2830 ( .A(A[150]), .B(n1887), .Z(O[150]) );
  AND U2831 ( .A(S), .B(n1888), .Z(n1887) );
  XOR U2832 ( .A(B[150]), .B(A[150]), .Z(n1888) );
  XOR U2833 ( .A(A[14]), .B(n1889), .Z(O[14]) );
  AND U2834 ( .A(S), .B(n1890), .Z(n1889) );
  XOR U2835 ( .A(B[14]), .B(A[14]), .Z(n1890) );
  XOR U2836 ( .A(A[149]), .B(n1891), .Z(O[149]) );
  AND U2837 ( .A(S), .B(n1892), .Z(n1891) );
  XOR U2838 ( .A(B[149]), .B(A[149]), .Z(n1892) );
  XOR U2839 ( .A(A[148]), .B(n1893), .Z(O[148]) );
  AND U2840 ( .A(S), .B(n1894), .Z(n1893) );
  XOR U2841 ( .A(B[148]), .B(A[148]), .Z(n1894) );
  XOR U2842 ( .A(A[147]), .B(n1895), .Z(O[147]) );
  AND U2843 ( .A(S), .B(n1896), .Z(n1895) );
  XOR U2844 ( .A(B[147]), .B(A[147]), .Z(n1896) );
  XOR U2845 ( .A(A[146]), .B(n1897), .Z(O[146]) );
  AND U2846 ( .A(S), .B(n1898), .Z(n1897) );
  XOR U2847 ( .A(B[146]), .B(A[146]), .Z(n1898) );
  XOR U2848 ( .A(A[145]), .B(n1899), .Z(O[145]) );
  AND U2849 ( .A(S), .B(n1900), .Z(n1899) );
  XOR U2850 ( .A(B[145]), .B(A[145]), .Z(n1900) );
  XOR U2851 ( .A(A[144]), .B(n1901), .Z(O[144]) );
  AND U2852 ( .A(S), .B(n1902), .Z(n1901) );
  XOR U2853 ( .A(B[144]), .B(A[144]), .Z(n1902) );
  XOR U2854 ( .A(A[143]), .B(n1903), .Z(O[143]) );
  AND U2855 ( .A(S), .B(n1904), .Z(n1903) );
  XOR U2856 ( .A(B[143]), .B(A[143]), .Z(n1904) );
  XOR U2857 ( .A(A[142]), .B(n1905), .Z(O[142]) );
  AND U2858 ( .A(S), .B(n1906), .Z(n1905) );
  XOR U2859 ( .A(B[142]), .B(A[142]), .Z(n1906) );
  XOR U2860 ( .A(A[141]), .B(n1907), .Z(O[141]) );
  AND U2861 ( .A(S), .B(n1908), .Z(n1907) );
  XOR U2862 ( .A(B[141]), .B(A[141]), .Z(n1908) );
  XOR U2863 ( .A(A[140]), .B(n1909), .Z(O[140]) );
  AND U2864 ( .A(S), .B(n1910), .Z(n1909) );
  XOR U2865 ( .A(B[140]), .B(A[140]), .Z(n1910) );
  XOR U2866 ( .A(A[13]), .B(n1911), .Z(O[13]) );
  AND U2867 ( .A(S), .B(n1912), .Z(n1911) );
  XOR U2868 ( .A(B[13]), .B(A[13]), .Z(n1912) );
  XOR U2869 ( .A(A[139]), .B(n1913), .Z(O[139]) );
  AND U2870 ( .A(S), .B(n1914), .Z(n1913) );
  XOR U2871 ( .A(B[139]), .B(A[139]), .Z(n1914) );
  XOR U2872 ( .A(A[138]), .B(n1915), .Z(O[138]) );
  AND U2873 ( .A(S), .B(n1916), .Z(n1915) );
  XOR U2874 ( .A(B[138]), .B(A[138]), .Z(n1916) );
  XOR U2875 ( .A(A[137]), .B(n1917), .Z(O[137]) );
  AND U2876 ( .A(S), .B(n1918), .Z(n1917) );
  XOR U2877 ( .A(B[137]), .B(A[137]), .Z(n1918) );
  XOR U2878 ( .A(A[136]), .B(n1919), .Z(O[136]) );
  AND U2879 ( .A(S), .B(n1920), .Z(n1919) );
  XOR U2880 ( .A(B[136]), .B(A[136]), .Z(n1920) );
  XOR U2881 ( .A(A[135]), .B(n1921), .Z(O[135]) );
  AND U2882 ( .A(S), .B(n1922), .Z(n1921) );
  XOR U2883 ( .A(B[135]), .B(A[135]), .Z(n1922) );
  XOR U2884 ( .A(A[134]), .B(n1923), .Z(O[134]) );
  AND U2885 ( .A(S), .B(n1924), .Z(n1923) );
  XOR U2886 ( .A(B[134]), .B(A[134]), .Z(n1924) );
  XOR U2887 ( .A(A[133]), .B(n1925), .Z(O[133]) );
  AND U2888 ( .A(S), .B(n1926), .Z(n1925) );
  XOR U2889 ( .A(B[133]), .B(A[133]), .Z(n1926) );
  XOR U2890 ( .A(A[132]), .B(n1927), .Z(O[132]) );
  AND U2891 ( .A(S), .B(n1928), .Z(n1927) );
  XOR U2892 ( .A(B[132]), .B(A[132]), .Z(n1928) );
  XOR U2893 ( .A(A[131]), .B(n1929), .Z(O[131]) );
  AND U2894 ( .A(S), .B(n1930), .Z(n1929) );
  XOR U2895 ( .A(B[131]), .B(A[131]), .Z(n1930) );
  XOR U2896 ( .A(A[130]), .B(n1931), .Z(O[130]) );
  AND U2897 ( .A(S), .B(n1932), .Z(n1931) );
  XOR U2898 ( .A(B[130]), .B(A[130]), .Z(n1932) );
  XOR U2899 ( .A(A[12]), .B(n1933), .Z(O[12]) );
  AND U2900 ( .A(S), .B(n1934), .Z(n1933) );
  XOR U2901 ( .A(B[12]), .B(A[12]), .Z(n1934) );
  XOR U2902 ( .A(A[129]), .B(n1935), .Z(O[129]) );
  AND U2903 ( .A(S), .B(n1936), .Z(n1935) );
  XOR U2904 ( .A(B[129]), .B(A[129]), .Z(n1936) );
  XOR U2905 ( .A(A[128]), .B(n1937), .Z(O[128]) );
  AND U2906 ( .A(S), .B(n1938), .Z(n1937) );
  XOR U2907 ( .A(B[128]), .B(A[128]), .Z(n1938) );
  XOR U2908 ( .A(A[127]), .B(n1939), .Z(O[127]) );
  AND U2909 ( .A(S), .B(n1940), .Z(n1939) );
  XOR U2910 ( .A(B[127]), .B(A[127]), .Z(n1940) );
  XOR U2911 ( .A(A[126]), .B(n1941), .Z(O[126]) );
  AND U2912 ( .A(S), .B(n1942), .Z(n1941) );
  XOR U2913 ( .A(B[126]), .B(A[126]), .Z(n1942) );
  XOR U2914 ( .A(A[125]), .B(n1943), .Z(O[125]) );
  AND U2915 ( .A(S), .B(n1944), .Z(n1943) );
  XOR U2916 ( .A(B[125]), .B(A[125]), .Z(n1944) );
  XOR U2917 ( .A(A[124]), .B(n1945), .Z(O[124]) );
  AND U2918 ( .A(S), .B(n1946), .Z(n1945) );
  XOR U2919 ( .A(B[124]), .B(A[124]), .Z(n1946) );
  XOR U2920 ( .A(A[123]), .B(n1947), .Z(O[123]) );
  AND U2921 ( .A(S), .B(n1948), .Z(n1947) );
  XOR U2922 ( .A(B[123]), .B(A[123]), .Z(n1948) );
  XOR U2923 ( .A(A[122]), .B(n1949), .Z(O[122]) );
  AND U2924 ( .A(S), .B(n1950), .Z(n1949) );
  XOR U2925 ( .A(B[122]), .B(A[122]), .Z(n1950) );
  XOR U2926 ( .A(A[121]), .B(n1951), .Z(O[121]) );
  AND U2927 ( .A(S), .B(n1952), .Z(n1951) );
  XOR U2928 ( .A(B[121]), .B(A[121]), .Z(n1952) );
  XOR U2929 ( .A(A[120]), .B(n1953), .Z(O[120]) );
  AND U2930 ( .A(S), .B(n1954), .Z(n1953) );
  XOR U2931 ( .A(B[120]), .B(A[120]), .Z(n1954) );
  XOR U2932 ( .A(A[11]), .B(n1955), .Z(O[11]) );
  AND U2933 ( .A(S), .B(n1956), .Z(n1955) );
  XOR U2934 ( .A(B[11]), .B(A[11]), .Z(n1956) );
  XOR U2935 ( .A(A[119]), .B(n1957), .Z(O[119]) );
  AND U2936 ( .A(S), .B(n1958), .Z(n1957) );
  XOR U2937 ( .A(B[119]), .B(A[119]), .Z(n1958) );
  XOR U2938 ( .A(A[118]), .B(n1959), .Z(O[118]) );
  AND U2939 ( .A(S), .B(n1960), .Z(n1959) );
  XOR U2940 ( .A(B[118]), .B(A[118]), .Z(n1960) );
  XOR U2941 ( .A(A[117]), .B(n1961), .Z(O[117]) );
  AND U2942 ( .A(S), .B(n1962), .Z(n1961) );
  XOR U2943 ( .A(B[117]), .B(A[117]), .Z(n1962) );
  XOR U2944 ( .A(A[116]), .B(n1963), .Z(O[116]) );
  AND U2945 ( .A(S), .B(n1964), .Z(n1963) );
  XOR U2946 ( .A(B[116]), .B(A[116]), .Z(n1964) );
  XOR U2947 ( .A(A[115]), .B(n1965), .Z(O[115]) );
  AND U2948 ( .A(S), .B(n1966), .Z(n1965) );
  XOR U2949 ( .A(B[115]), .B(A[115]), .Z(n1966) );
  XOR U2950 ( .A(A[114]), .B(n1967), .Z(O[114]) );
  AND U2951 ( .A(S), .B(n1968), .Z(n1967) );
  XOR U2952 ( .A(B[114]), .B(A[114]), .Z(n1968) );
  XOR U2953 ( .A(A[113]), .B(n1969), .Z(O[113]) );
  AND U2954 ( .A(S), .B(n1970), .Z(n1969) );
  XOR U2955 ( .A(B[113]), .B(A[113]), .Z(n1970) );
  XOR U2956 ( .A(A[112]), .B(n1971), .Z(O[112]) );
  AND U2957 ( .A(S), .B(n1972), .Z(n1971) );
  XOR U2958 ( .A(B[112]), .B(A[112]), .Z(n1972) );
  XOR U2959 ( .A(A[111]), .B(n1973), .Z(O[111]) );
  AND U2960 ( .A(S), .B(n1974), .Z(n1973) );
  XOR U2961 ( .A(B[111]), .B(A[111]), .Z(n1974) );
  XOR U2962 ( .A(A[110]), .B(n1975), .Z(O[110]) );
  AND U2963 ( .A(S), .B(n1976), .Z(n1975) );
  XOR U2964 ( .A(B[110]), .B(A[110]), .Z(n1976) );
  XOR U2965 ( .A(A[10]), .B(n1977), .Z(O[10]) );
  AND U2966 ( .A(S), .B(n1978), .Z(n1977) );
  XOR U2967 ( .A(B[10]), .B(A[10]), .Z(n1978) );
  XOR U2968 ( .A(A[109]), .B(n1979), .Z(O[109]) );
  AND U2969 ( .A(S), .B(n1980), .Z(n1979) );
  XOR U2970 ( .A(B[109]), .B(A[109]), .Z(n1980) );
  XOR U2971 ( .A(A[108]), .B(n1981), .Z(O[108]) );
  AND U2972 ( .A(S), .B(n1982), .Z(n1981) );
  XOR U2973 ( .A(B[108]), .B(A[108]), .Z(n1982) );
  XOR U2974 ( .A(A[107]), .B(n1983), .Z(O[107]) );
  AND U2975 ( .A(S), .B(n1984), .Z(n1983) );
  XOR U2976 ( .A(B[107]), .B(A[107]), .Z(n1984) );
  XOR U2977 ( .A(A[106]), .B(n1985), .Z(O[106]) );
  AND U2978 ( .A(S), .B(n1986), .Z(n1985) );
  XOR U2979 ( .A(B[106]), .B(A[106]), .Z(n1986) );
  XOR U2980 ( .A(A[105]), .B(n1987), .Z(O[105]) );
  AND U2981 ( .A(S), .B(n1988), .Z(n1987) );
  XOR U2982 ( .A(B[105]), .B(A[105]), .Z(n1988) );
  XOR U2983 ( .A(A[104]), .B(n1989), .Z(O[104]) );
  AND U2984 ( .A(S), .B(n1990), .Z(n1989) );
  XOR U2985 ( .A(B[104]), .B(A[104]), .Z(n1990) );
  XOR U2986 ( .A(A[103]), .B(n1991), .Z(O[103]) );
  AND U2987 ( .A(S), .B(n1992), .Z(n1991) );
  XOR U2988 ( .A(B[103]), .B(A[103]), .Z(n1992) );
  XOR U2989 ( .A(A[102]), .B(n1993), .Z(O[102]) );
  AND U2990 ( .A(S), .B(n1994), .Z(n1993) );
  XOR U2991 ( .A(B[102]), .B(A[102]), .Z(n1994) );
  XOR U2992 ( .A(A[1023]), .B(n1995), .Z(O[1023]) );
  AND U2993 ( .A(S), .B(n1996), .Z(n1995) );
  XOR U2994 ( .A(B[1023]), .B(A[1023]), .Z(n1996) );
  XOR U2995 ( .A(A[1022]), .B(n1997), .Z(O[1022]) );
  AND U2996 ( .A(S), .B(n1998), .Z(n1997) );
  XOR U2997 ( .A(B[1022]), .B(A[1022]), .Z(n1998) );
  XOR U2998 ( .A(A[1021]), .B(n1999), .Z(O[1021]) );
  AND U2999 ( .A(S), .B(n2000), .Z(n1999) );
  XOR U3000 ( .A(B[1021]), .B(A[1021]), .Z(n2000) );
  XOR U3001 ( .A(A[1020]), .B(n2001), .Z(O[1020]) );
  AND U3002 ( .A(S), .B(n2002), .Z(n2001) );
  XOR U3003 ( .A(B[1020]), .B(A[1020]), .Z(n2002) );
  XOR U3004 ( .A(A[101]), .B(n2003), .Z(O[101]) );
  AND U3005 ( .A(S), .B(n2004), .Z(n2003) );
  XOR U3006 ( .A(B[101]), .B(A[101]), .Z(n2004) );
  XOR U3007 ( .A(A[1019]), .B(n2005), .Z(O[1019]) );
  AND U3008 ( .A(S), .B(n2006), .Z(n2005) );
  XOR U3009 ( .A(B[1019]), .B(A[1019]), .Z(n2006) );
  XOR U3010 ( .A(A[1018]), .B(n2007), .Z(O[1018]) );
  AND U3011 ( .A(S), .B(n2008), .Z(n2007) );
  XOR U3012 ( .A(B[1018]), .B(A[1018]), .Z(n2008) );
  XOR U3013 ( .A(A[1017]), .B(n2009), .Z(O[1017]) );
  AND U3014 ( .A(S), .B(n2010), .Z(n2009) );
  XOR U3015 ( .A(B[1017]), .B(A[1017]), .Z(n2010) );
  XOR U3016 ( .A(A[1016]), .B(n2011), .Z(O[1016]) );
  AND U3017 ( .A(S), .B(n2012), .Z(n2011) );
  XOR U3018 ( .A(B[1016]), .B(A[1016]), .Z(n2012) );
  XOR U3019 ( .A(A[1015]), .B(n2013), .Z(O[1015]) );
  AND U3020 ( .A(S), .B(n2014), .Z(n2013) );
  XOR U3021 ( .A(B[1015]), .B(A[1015]), .Z(n2014) );
  XOR U3022 ( .A(A[1014]), .B(n2015), .Z(O[1014]) );
  AND U3023 ( .A(S), .B(n2016), .Z(n2015) );
  XOR U3024 ( .A(B[1014]), .B(A[1014]), .Z(n2016) );
  XOR U3025 ( .A(A[1013]), .B(n2017), .Z(O[1013]) );
  AND U3026 ( .A(S), .B(n2018), .Z(n2017) );
  XOR U3027 ( .A(B[1013]), .B(A[1013]), .Z(n2018) );
  XOR U3028 ( .A(A[1012]), .B(n2019), .Z(O[1012]) );
  AND U3029 ( .A(S), .B(n2020), .Z(n2019) );
  XOR U3030 ( .A(B[1012]), .B(A[1012]), .Z(n2020) );
  XOR U3031 ( .A(A[1011]), .B(n2021), .Z(O[1011]) );
  AND U3032 ( .A(S), .B(n2022), .Z(n2021) );
  XOR U3033 ( .A(B[1011]), .B(A[1011]), .Z(n2022) );
  XOR U3034 ( .A(A[1010]), .B(n2023), .Z(O[1010]) );
  AND U3035 ( .A(S), .B(n2024), .Z(n2023) );
  XOR U3036 ( .A(B[1010]), .B(A[1010]), .Z(n2024) );
  XOR U3037 ( .A(A[100]), .B(n2025), .Z(O[100]) );
  AND U3038 ( .A(S), .B(n2026), .Z(n2025) );
  XOR U3039 ( .A(B[100]), .B(A[100]), .Z(n2026) );
  XOR U3040 ( .A(A[1009]), .B(n2027), .Z(O[1009]) );
  AND U3041 ( .A(S), .B(n2028), .Z(n2027) );
  XOR U3042 ( .A(B[1009]), .B(A[1009]), .Z(n2028) );
  XOR U3043 ( .A(A[1008]), .B(n2029), .Z(O[1008]) );
  AND U3044 ( .A(S), .B(n2030), .Z(n2029) );
  XOR U3045 ( .A(B[1008]), .B(A[1008]), .Z(n2030) );
  XOR U3046 ( .A(A[1007]), .B(n2031), .Z(O[1007]) );
  AND U3047 ( .A(S), .B(n2032), .Z(n2031) );
  XOR U3048 ( .A(B[1007]), .B(A[1007]), .Z(n2032) );
  XOR U3049 ( .A(A[1006]), .B(n2033), .Z(O[1006]) );
  AND U3050 ( .A(S), .B(n2034), .Z(n2033) );
  XOR U3051 ( .A(B[1006]), .B(A[1006]), .Z(n2034) );
  XOR U3052 ( .A(A[1005]), .B(n2035), .Z(O[1005]) );
  AND U3053 ( .A(S), .B(n2036), .Z(n2035) );
  XOR U3054 ( .A(B[1005]), .B(A[1005]), .Z(n2036) );
  XOR U3055 ( .A(A[1004]), .B(n2037), .Z(O[1004]) );
  AND U3056 ( .A(S), .B(n2038), .Z(n2037) );
  XOR U3057 ( .A(B[1004]), .B(A[1004]), .Z(n2038) );
  XOR U3058 ( .A(A[1003]), .B(n2039), .Z(O[1003]) );
  AND U3059 ( .A(S), .B(n2040), .Z(n2039) );
  XOR U3060 ( .A(B[1003]), .B(A[1003]), .Z(n2040) );
  XOR U3061 ( .A(A[1002]), .B(n2041), .Z(O[1002]) );
  AND U3062 ( .A(S), .B(n2042), .Z(n2041) );
  XOR U3063 ( .A(B[1002]), .B(A[1002]), .Z(n2042) );
  XOR U3064 ( .A(A[1001]), .B(n2043), .Z(O[1001]) );
  AND U3065 ( .A(S), .B(n2044), .Z(n2043) );
  XOR U3066 ( .A(B[1001]), .B(A[1001]), .Z(n2044) );
  XOR U3067 ( .A(A[1000]), .B(n2045), .Z(O[1000]) );
  AND U3068 ( .A(S), .B(n2046), .Z(n2045) );
  XOR U3069 ( .A(B[1000]), .B(A[1000]), .Z(n2046) );
  XOR U3070 ( .A(A[0]), .B(n2047), .Z(O[0]) );
  AND U3071 ( .A(S), .B(n2048), .Z(n2047) );
  XOR U3072 ( .A(B[0]), .B(A[0]), .Z(n2048) );
endmodule


module MUX_N1026_0 ( A, B, S, O );
  input [1025:0] A;
  input [1025:0] B;
  output [1025:0] O;
  input S;


  ANDN U1 ( .B(A[9]), .A(S), .Z(O[9]) );
  ANDN U2 ( .B(A[99]), .A(S), .Z(O[99]) );
  ANDN U3 ( .B(A[999]), .A(S), .Z(O[999]) );
  ANDN U4 ( .B(A[998]), .A(S), .Z(O[998]) );
  ANDN U5 ( .B(A[997]), .A(S), .Z(O[997]) );
  ANDN U6 ( .B(A[996]), .A(S), .Z(O[996]) );
  ANDN U7 ( .B(A[995]), .A(S), .Z(O[995]) );
  ANDN U8 ( .B(A[994]), .A(S), .Z(O[994]) );
  ANDN U9 ( .B(A[993]), .A(S), .Z(O[993]) );
  ANDN U10 ( .B(A[992]), .A(S), .Z(O[992]) );
  ANDN U11 ( .B(A[991]), .A(S), .Z(O[991]) );
  ANDN U12 ( .B(A[990]), .A(S), .Z(O[990]) );
  ANDN U13 ( .B(A[98]), .A(S), .Z(O[98]) );
  ANDN U14 ( .B(A[989]), .A(S), .Z(O[989]) );
  ANDN U15 ( .B(A[988]), .A(S), .Z(O[988]) );
  ANDN U16 ( .B(A[987]), .A(S), .Z(O[987]) );
  ANDN U17 ( .B(A[986]), .A(S), .Z(O[986]) );
  ANDN U18 ( .B(A[985]), .A(S), .Z(O[985]) );
  ANDN U19 ( .B(A[984]), .A(S), .Z(O[984]) );
  ANDN U20 ( .B(A[983]), .A(S), .Z(O[983]) );
  ANDN U21 ( .B(A[982]), .A(S), .Z(O[982]) );
  ANDN U22 ( .B(A[981]), .A(S), .Z(O[981]) );
  ANDN U23 ( .B(A[980]), .A(S), .Z(O[980]) );
  ANDN U24 ( .B(A[97]), .A(S), .Z(O[97]) );
  ANDN U25 ( .B(A[979]), .A(S), .Z(O[979]) );
  ANDN U26 ( .B(A[978]), .A(S), .Z(O[978]) );
  ANDN U27 ( .B(A[977]), .A(S), .Z(O[977]) );
  ANDN U28 ( .B(A[976]), .A(S), .Z(O[976]) );
  ANDN U29 ( .B(A[975]), .A(S), .Z(O[975]) );
  ANDN U30 ( .B(A[974]), .A(S), .Z(O[974]) );
  ANDN U31 ( .B(A[973]), .A(S), .Z(O[973]) );
  ANDN U32 ( .B(A[972]), .A(S), .Z(O[972]) );
  ANDN U33 ( .B(A[971]), .A(S), .Z(O[971]) );
  ANDN U34 ( .B(A[970]), .A(S), .Z(O[970]) );
  ANDN U35 ( .B(A[96]), .A(S), .Z(O[96]) );
  ANDN U36 ( .B(A[969]), .A(S), .Z(O[969]) );
  ANDN U37 ( .B(A[968]), .A(S), .Z(O[968]) );
  ANDN U38 ( .B(A[967]), .A(S), .Z(O[967]) );
  ANDN U39 ( .B(A[966]), .A(S), .Z(O[966]) );
  ANDN U40 ( .B(A[965]), .A(S), .Z(O[965]) );
  ANDN U41 ( .B(A[964]), .A(S), .Z(O[964]) );
  ANDN U42 ( .B(A[963]), .A(S), .Z(O[963]) );
  ANDN U43 ( .B(A[962]), .A(S), .Z(O[962]) );
  ANDN U44 ( .B(A[961]), .A(S), .Z(O[961]) );
  ANDN U45 ( .B(A[960]), .A(S), .Z(O[960]) );
  ANDN U46 ( .B(A[95]), .A(S), .Z(O[95]) );
  ANDN U47 ( .B(A[959]), .A(S), .Z(O[959]) );
  ANDN U48 ( .B(A[958]), .A(S), .Z(O[958]) );
  ANDN U49 ( .B(A[957]), .A(S), .Z(O[957]) );
  ANDN U50 ( .B(A[956]), .A(S), .Z(O[956]) );
  ANDN U51 ( .B(A[955]), .A(S), .Z(O[955]) );
  ANDN U52 ( .B(A[954]), .A(S), .Z(O[954]) );
  ANDN U53 ( .B(A[953]), .A(S), .Z(O[953]) );
  ANDN U54 ( .B(A[952]), .A(S), .Z(O[952]) );
  ANDN U55 ( .B(A[951]), .A(S), .Z(O[951]) );
  ANDN U56 ( .B(A[950]), .A(S), .Z(O[950]) );
  ANDN U57 ( .B(A[94]), .A(S), .Z(O[94]) );
  ANDN U58 ( .B(A[949]), .A(S), .Z(O[949]) );
  ANDN U59 ( .B(A[948]), .A(S), .Z(O[948]) );
  ANDN U60 ( .B(A[947]), .A(S), .Z(O[947]) );
  ANDN U61 ( .B(A[946]), .A(S), .Z(O[946]) );
  ANDN U62 ( .B(A[945]), .A(S), .Z(O[945]) );
  ANDN U63 ( .B(A[944]), .A(S), .Z(O[944]) );
  ANDN U64 ( .B(A[943]), .A(S), .Z(O[943]) );
  ANDN U65 ( .B(A[942]), .A(S), .Z(O[942]) );
  ANDN U66 ( .B(A[941]), .A(S), .Z(O[941]) );
  ANDN U67 ( .B(A[940]), .A(S), .Z(O[940]) );
  ANDN U68 ( .B(A[93]), .A(S), .Z(O[93]) );
  ANDN U69 ( .B(A[939]), .A(S), .Z(O[939]) );
  ANDN U70 ( .B(A[938]), .A(S), .Z(O[938]) );
  ANDN U71 ( .B(A[937]), .A(S), .Z(O[937]) );
  ANDN U72 ( .B(A[936]), .A(S), .Z(O[936]) );
  ANDN U73 ( .B(A[935]), .A(S), .Z(O[935]) );
  ANDN U74 ( .B(A[934]), .A(S), .Z(O[934]) );
  ANDN U75 ( .B(A[933]), .A(S), .Z(O[933]) );
  ANDN U76 ( .B(A[932]), .A(S), .Z(O[932]) );
  ANDN U77 ( .B(A[931]), .A(S), .Z(O[931]) );
  ANDN U78 ( .B(A[930]), .A(S), .Z(O[930]) );
  ANDN U79 ( .B(A[92]), .A(S), .Z(O[92]) );
  ANDN U80 ( .B(A[929]), .A(S), .Z(O[929]) );
  ANDN U81 ( .B(A[928]), .A(S), .Z(O[928]) );
  ANDN U82 ( .B(A[927]), .A(S), .Z(O[927]) );
  ANDN U83 ( .B(A[926]), .A(S), .Z(O[926]) );
  ANDN U84 ( .B(A[925]), .A(S), .Z(O[925]) );
  ANDN U85 ( .B(A[924]), .A(S), .Z(O[924]) );
  ANDN U86 ( .B(A[923]), .A(S), .Z(O[923]) );
  ANDN U87 ( .B(A[922]), .A(S), .Z(O[922]) );
  ANDN U88 ( .B(A[921]), .A(S), .Z(O[921]) );
  ANDN U89 ( .B(A[920]), .A(S), .Z(O[920]) );
  ANDN U90 ( .B(A[91]), .A(S), .Z(O[91]) );
  ANDN U91 ( .B(A[919]), .A(S), .Z(O[919]) );
  ANDN U92 ( .B(A[918]), .A(S), .Z(O[918]) );
  ANDN U93 ( .B(A[917]), .A(S), .Z(O[917]) );
  ANDN U94 ( .B(A[916]), .A(S), .Z(O[916]) );
  ANDN U95 ( .B(A[915]), .A(S), .Z(O[915]) );
  ANDN U96 ( .B(A[914]), .A(S), .Z(O[914]) );
  ANDN U97 ( .B(A[913]), .A(S), .Z(O[913]) );
  ANDN U98 ( .B(A[912]), .A(S), .Z(O[912]) );
  ANDN U99 ( .B(A[911]), .A(S), .Z(O[911]) );
  ANDN U100 ( .B(A[910]), .A(S), .Z(O[910]) );
  ANDN U101 ( .B(A[90]), .A(S), .Z(O[90]) );
  ANDN U102 ( .B(A[909]), .A(S), .Z(O[909]) );
  ANDN U103 ( .B(A[908]), .A(S), .Z(O[908]) );
  ANDN U104 ( .B(A[907]), .A(S), .Z(O[907]) );
  ANDN U105 ( .B(A[906]), .A(S), .Z(O[906]) );
  ANDN U106 ( .B(A[905]), .A(S), .Z(O[905]) );
  ANDN U107 ( .B(A[904]), .A(S), .Z(O[904]) );
  ANDN U108 ( .B(A[903]), .A(S), .Z(O[903]) );
  ANDN U109 ( .B(A[902]), .A(S), .Z(O[902]) );
  ANDN U110 ( .B(A[901]), .A(S), .Z(O[901]) );
  ANDN U111 ( .B(A[900]), .A(S), .Z(O[900]) );
  ANDN U112 ( .B(A[8]), .A(S), .Z(O[8]) );
  ANDN U113 ( .B(A[89]), .A(S), .Z(O[89]) );
  ANDN U114 ( .B(A[899]), .A(S), .Z(O[899]) );
  ANDN U115 ( .B(A[898]), .A(S), .Z(O[898]) );
  ANDN U116 ( .B(A[897]), .A(S), .Z(O[897]) );
  ANDN U117 ( .B(A[896]), .A(S), .Z(O[896]) );
  ANDN U118 ( .B(A[895]), .A(S), .Z(O[895]) );
  ANDN U119 ( .B(A[894]), .A(S), .Z(O[894]) );
  ANDN U120 ( .B(A[893]), .A(S), .Z(O[893]) );
  ANDN U121 ( .B(A[892]), .A(S), .Z(O[892]) );
  ANDN U122 ( .B(A[891]), .A(S), .Z(O[891]) );
  ANDN U123 ( .B(A[890]), .A(S), .Z(O[890]) );
  ANDN U124 ( .B(A[88]), .A(S), .Z(O[88]) );
  ANDN U125 ( .B(A[889]), .A(S), .Z(O[889]) );
  ANDN U126 ( .B(A[888]), .A(S), .Z(O[888]) );
  ANDN U127 ( .B(A[887]), .A(S), .Z(O[887]) );
  ANDN U128 ( .B(A[886]), .A(S), .Z(O[886]) );
  ANDN U129 ( .B(A[885]), .A(S), .Z(O[885]) );
  ANDN U130 ( .B(A[884]), .A(S), .Z(O[884]) );
  ANDN U131 ( .B(A[883]), .A(S), .Z(O[883]) );
  ANDN U132 ( .B(A[882]), .A(S), .Z(O[882]) );
  ANDN U133 ( .B(A[881]), .A(S), .Z(O[881]) );
  ANDN U134 ( .B(A[880]), .A(S), .Z(O[880]) );
  ANDN U135 ( .B(A[87]), .A(S), .Z(O[87]) );
  ANDN U136 ( .B(A[879]), .A(S), .Z(O[879]) );
  ANDN U137 ( .B(A[878]), .A(S), .Z(O[878]) );
  ANDN U138 ( .B(A[877]), .A(S), .Z(O[877]) );
  ANDN U139 ( .B(A[876]), .A(S), .Z(O[876]) );
  ANDN U140 ( .B(A[875]), .A(S), .Z(O[875]) );
  ANDN U141 ( .B(A[874]), .A(S), .Z(O[874]) );
  ANDN U142 ( .B(A[873]), .A(S), .Z(O[873]) );
  ANDN U143 ( .B(A[872]), .A(S), .Z(O[872]) );
  ANDN U144 ( .B(A[871]), .A(S), .Z(O[871]) );
  ANDN U145 ( .B(A[870]), .A(S), .Z(O[870]) );
  ANDN U146 ( .B(A[86]), .A(S), .Z(O[86]) );
  ANDN U147 ( .B(A[869]), .A(S), .Z(O[869]) );
  ANDN U148 ( .B(A[868]), .A(S), .Z(O[868]) );
  ANDN U149 ( .B(A[867]), .A(S), .Z(O[867]) );
  ANDN U150 ( .B(A[866]), .A(S), .Z(O[866]) );
  ANDN U151 ( .B(A[865]), .A(S), .Z(O[865]) );
  ANDN U152 ( .B(A[864]), .A(S), .Z(O[864]) );
  ANDN U153 ( .B(A[863]), .A(S), .Z(O[863]) );
  ANDN U154 ( .B(A[862]), .A(S), .Z(O[862]) );
  ANDN U155 ( .B(A[861]), .A(S), .Z(O[861]) );
  ANDN U156 ( .B(A[860]), .A(S), .Z(O[860]) );
  ANDN U157 ( .B(A[85]), .A(S), .Z(O[85]) );
  ANDN U158 ( .B(A[859]), .A(S), .Z(O[859]) );
  ANDN U159 ( .B(A[858]), .A(S), .Z(O[858]) );
  ANDN U160 ( .B(A[857]), .A(S), .Z(O[857]) );
  ANDN U161 ( .B(A[856]), .A(S), .Z(O[856]) );
  ANDN U162 ( .B(A[855]), .A(S), .Z(O[855]) );
  ANDN U163 ( .B(A[854]), .A(S), .Z(O[854]) );
  ANDN U164 ( .B(A[853]), .A(S), .Z(O[853]) );
  ANDN U165 ( .B(A[852]), .A(S), .Z(O[852]) );
  ANDN U166 ( .B(A[851]), .A(S), .Z(O[851]) );
  ANDN U167 ( .B(A[850]), .A(S), .Z(O[850]) );
  ANDN U168 ( .B(A[84]), .A(S), .Z(O[84]) );
  ANDN U169 ( .B(A[849]), .A(S), .Z(O[849]) );
  ANDN U170 ( .B(A[848]), .A(S), .Z(O[848]) );
  ANDN U171 ( .B(A[847]), .A(S), .Z(O[847]) );
  ANDN U172 ( .B(A[846]), .A(S), .Z(O[846]) );
  ANDN U173 ( .B(A[845]), .A(S), .Z(O[845]) );
  ANDN U174 ( .B(A[844]), .A(S), .Z(O[844]) );
  ANDN U175 ( .B(A[843]), .A(S), .Z(O[843]) );
  ANDN U176 ( .B(A[842]), .A(S), .Z(O[842]) );
  ANDN U177 ( .B(A[841]), .A(S), .Z(O[841]) );
  ANDN U178 ( .B(A[840]), .A(S), .Z(O[840]) );
  ANDN U179 ( .B(A[83]), .A(S), .Z(O[83]) );
  ANDN U180 ( .B(A[839]), .A(S), .Z(O[839]) );
  ANDN U181 ( .B(A[838]), .A(S), .Z(O[838]) );
  ANDN U182 ( .B(A[837]), .A(S), .Z(O[837]) );
  ANDN U183 ( .B(A[836]), .A(S), .Z(O[836]) );
  ANDN U184 ( .B(A[835]), .A(S), .Z(O[835]) );
  ANDN U185 ( .B(A[834]), .A(S), .Z(O[834]) );
  ANDN U186 ( .B(A[833]), .A(S), .Z(O[833]) );
  ANDN U187 ( .B(A[832]), .A(S), .Z(O[832]) );
  ANDN U188 ( .B(A[831]), .A(S), .Z(O[831]) );
  ANDN U189 ( .B(A[830]), .A(S), .Z(O[830]) );
  ANDN U190 ( .B(A[82]), .A(S), .Z(O[82]) );
  ANDN U191 ( .B(A[829]), .A(S), .Z(O[829]) );
  ANDN U192 ( .B(A[828]), .A(S), .Z(O[828]) );
  ANDN U193 ( .B(A[827]), .A(S), .Z(O[827]) );
  ANDN U194 ( .B(A[826]), .A(S), .Z(O[826]) );
  ANDN U195 ( .B(A[825]), .A(S), .Z(O[825]) );
  ANDN U196 ( .B(A[824]), .A(S), .Z(O[824]) );
  ANDN U197 ( .B(A[823]), .A(S), .Z(O[823]) );
  ANDN U198 ( .B(A[822]), .A(S), .Z(O[822]) );
  ANDN U199 ( .B(A[821]), .A(S), .Z(O[821]) );
  ANDN U200 ( .B(A[820]), .A(S), .Z(O[820]) );
  ANDN U201 ( .B(A[81]), .A(S), .Z(O[81]) );
  ANDN U202 ( .B(A[819]), .A(S), .Z(O[819]) );
  ANDN U203 ( .B(A[818]), .A(S), .Z(O[818]) );
  ANDN U204 ( .B(A[817]), .A(S), .Z(O[817]) );
  ANDN U205 ( .B(A[816]), .A(S), .Z(O[816]) );
  ANDN U206 ( .B(A[815]), .A(S), .Z(O[815]) );
  ANDN U207 ( .B(A[814]), .A(S), .Z(O[814]) );
  ANDN U208 ( .B(A[813]), .A(S), .Z(O[813]) );
  ANDN U209 ( .B(A[812]), .A(S), .Z(O[812]) );
  ANDN U210 ( .B(A[811]), .A(S), .Z(O[811]) );
  ANDN U211 ( .B(A[810]), .A(S), .Z(O[810]) );
  ANDN U212 ( .B(A[80]), .A(S), .Z(O[80]) );
  ANDN U213 ( .B(A[809]), .A(S), .Z(O[809]) );
  ANDN U214 ( .B(A[808]), .A(S), .Z(O[808]) );
  ANDN U215 ( .B(A[807]), .A(S), .Z(O[807]) );
  ANDN U216 ( .B(A[806]), .A(S), .Z(O[806]) );
  ANDN U217 ( .B(A[805]), .A(S), .Z(O[805]) );
  ANDN U218 ( .B(A[804]), .A(S), .Z(O[804]) );
  ANDN U219 ( .B(A[803]), .A(S), .Z(O[803]) );
  ANDN U220 ( .B(A[802]), .A(S), .Z(O[802]) );
  ANDN U221 ( .B(A[801]), .A(S), .Z(O[801]) );
  ANDN U222 ( .B(A[800]), .A(S), .Z(O[800]) );
  ANDN U223 ( .B(A[7]), .A(S), .Z(O[7]) );
  ANDN U224 ( .B(A[79]), .A(S), .Z(O[79]) );
  ANDN U225 ( .B(A[799]), .A(S), .Z(O[799]) );
  ANDN U226 ( .B(A[798]), .A(S), .Z(O[798]) );
  ANDN U227 ( .B(A[797]), .A(S), .Z(O[797]) );
  ANDN U228 ( .B(A[796]), .A(S), .Z(O[796]) );
  ANDN U229 ( .B(A[795]), .A(S), .Z(O[795]) );
  ANDN U230 ( .B(A[794]), .A(S), .Z(O[794]) );
  ANDN U231 ( .B(A[793]), .A(S), .Z(O[793]) );
  ANDN U232 ( .B(A[792]), .A(S), .Z(O[792]) );
  ANDN U233 ( .B(A[791]), .A(S), .Z(O[791]) );
  ANDN U234 ( .B(A[790]), .A(S), .Z(O[790]) );
  ANDN U235 ( .B(A[78]), .A(S), .Z(O[78]) );
  ANDN U236 ( .B(A[789]), .A(S), .Z(O[789]) );
  ANDN U237 ( .B(A[788]), .A(S), .Z(O[788]) );
  ANDN U238 ( .B(A[787]), .A(S), .Z(O[787]) );
  ANDN U239 ( .B(A[786]), .A(S), .Z(O[786]) );
  ANDN U240 ( .B(A[785]), .A(S), .Z(O[785]) );
  ANDN U241 ( .B(A[784]), .A(S), .Z(O[784]) );
  ANDN U242 ( .B(A[783]), .A(S), .Z(O[783]) );
  ANDN U243 ( .B(A[782]), .A(S), .Z(O[782]) );
  ANDN U244 ( .B(A[781]), .A(S), .Z(O[781]) );
  ANDN U245 ( .B(A[780]), .A(S), .Z(O[780]) );
  ANDN U246 ( .B(A[77]), .A(S), .Z(O[77]) );
  ANDN U247 ( .B(A[779]), .A(S), .Z(O[779]) );
  ANDN U248 ( .B(A[778]), .A(S), .Z(O[778]) );
  ANDN U249 ( .B(A[777]), .A(S), .Z(O[777]) );
  ANDN U250 ( .B(A[776]), .A(S), .Z(O[776]) );
  ANDN U251 ( .B(A[775]), .A(S), .Z(O[775]) );
  ANDN U252 ( .B(A[774]), .A(S), .Z(O[774]) );
  ANDN U253 ( .B(A[773]), .A(S), .Z(O[773]) );
  ANDN U254 ( .B(A[772]), .A(S), .Z(O[772]) );
  ANDN U255 ( .B(A[771]), .A(S), .Z(O[771]) );
  ANDN U256 ( .B(A[770]), .A(S), .Z(O[770]) );
  ANDN U257 ( .B(A[76]), .A(S), .Z(O[76]) );
  ANDN U258 ( .B(A[769]), .A(S), .Z(O[769]) );
  ANDN U259 ( .B(A[768]), .A(S), .Z(O[768]) );
  ANDN U260 ( .B(A[767]), .A(S), .Z(O[767]) );
  ANDN U261 ( .B(A[766]), .A(S), .Z(O[766]) );
  ANDN U262 ( .B(A[765]), .A(S), .Z(O[765]) );
  ANDN U263 ( .B(A[764]), .A(S), .Z(O[764]) );
  ANDN U264 ( .B(A[763]), .A(S), .Z(O[763]) );
  ANDN U265 ( .B(A[762]), .A(S), .Z(O[762]) );
  ANDN U266 ( .B(A[761]), .A(S), .Z(O[761]) );
  ANDN U267 ( .B(A[760]), .A(S), .Z(O[760]) );
  ANDN U268 ( .B(A[75]), .A(S), .Z(O[75]) );
  ANDN U269 ( .B(A[759]), .A(S), .Z(O[759]) );
  ANDN U270 ( .B(A[758]), .A(S), .Z(O[758]) );
  ANDN U271 ( .B(A[757]), .A(S), .Z(O[757]) );
  ANDN U272 ( .B(A[756]), .A(S), .Z(O[756]) );
  ANDN U273 ( .B(A[755]), .A(S), .Z(O[755]) );
  ANDN U274 ( .B(A[754]), .A(S), .Z(O[754]) );
  ANDN U275 ( .B(A[753]), .A(S), .Z(O[753]) );
  ANDN U276 ( .B(A[752]), .A(S), .Z(O[752]) );
  ANDN U277 ( .B(A[751]), .A(S), .Z(O[751]) );
  ANDN U278 ( .B(A[750]), .A(S), .Z(O[750]) );
  ANDN U279 ( .B(A[74]), .A(S), .Z(O[74]) );
  ANDN U280 ( .B(A[749]), .A(S), .Z(O[749]) );
  ANDN U281 ( .B(A[748]), .A(S), .Z(O[748]) );
  ANDN U282 ( .B(A[747]), .A(S), .Z(O[747]) );
  ANDN U283 ( .B(A[746]), .A(S), .Z(O[746]) );
  ANDN U284 ( .B(A[745]), .A(S), .Z(O[745]) );
  ANDN U285 ( .B(A[744]), .A(S), .Z(O[744]) );
  ANDN U286 ( .B(A[743]), .A(S), .Z(O[743]) );
  ANDN U287 ( .B(A[742]), .A(S), .Z(O[742]) );
  ANDN U288 ( .B(A[741]), .A(S), .Z(O[741]) );
  ANDN U289 ( .B(A[740]), .A(S), .Z(O[740]) );
  ANDN U290 ( .B(A[73]), .A(S), .Z(O[73]) );
  ANDN U291 ( .B(A[739]), .A(S), .Z(O[739]) );
  ANDN U292 ( .B(A[738]), .A(S), .Z(O[738]) );
  ANDN U293 ( .B(A[737]), .A(S), .Z(O[737]) );
  ANDN U294 ( .B(A[736]), .A(S), .Z(O[736]) );
  ANDN U295 ( .B(A[735]), .A(S), .Z(O[735]) );
  ANDN U296 ( .B(A[734]), .A(S), .Z(O[734]) );
  ANDN U297 ( .B(A[733]), .A(S), .Z(O[733]) );
  ANDN U298 ( .B(A[732]), .A(S), .Z(O[732]) );
  ANDN U299 ( .B(A[731]), .A(S), .Z(O[731]) );
  ANDN U300 ( .B(A[730]), .A(S), .Z(O[730]) );
  ANDN U301 ( .B(A[72]), .A(S), .Z(O[72]) );
  ANDN U302 ( .B(A[729]), .A(S), .Z(O[729]) );
  ANDN U303 ( .B(A[728]), .A(S), .Z(O[728]) );
  ANDN U304 ( .B(A[727]), .A(S), .Z(O[727]) );
  ANDN U305 ( .B(A[726]), .A(S), .Z(O[726]) );
  ANDN U306 ( .B(A[725]), .A(S), .Z(O[725]) );
  ANDN U307 ( .B(A[724]), .A(S), .Z(O[724]) );
  ANDN U308 ( .B(A[723]), .A(S), .Z(O[723]) );
  ANDN U309 ( .B(A[722]), .A(S), .Z(O[722]) );
  ANDN U310 ( .B(A[721]), .A(S), .Z(O[721]) );
  ANDN U311 ( .B(A[720]), .A(S), .Z(O[720]) );
  ANDN U312 ( .B(A[71]), .A(S), .Z(O[71]) );
  ANDN U313 ( .B(A[719]), .A(S), .Z(O[719]) );
  ANDN U314 ( .B(A[718]), .A(S), .Z(O[718]) );
  ANDN U315 ( .B(A[717]), .A(S), .Z(O[717]) );
  ANDN U316 ( .B(A[716]), .A(S), .Z(O[716]) );
  ANDN U317 ( .B(A[715]), .A(S), .Z(O[715]) );
  ANDN U318 ( .B(A[714]), .A(S), .Z(O[714]) );
  ANDN U319 ( .B(A[713]), .A(S), .Z(O[713]) );
  ANDN U320 ( .B(A[712]), .A(S), .Z(O[712]) );
  ANDN U321 ( .B(A[711]), .A(S), .Z(O[711]) );
  ANDN U322 ( .B(A[710]), .A(S), .Z(O[710]) );
  ANDN U323 ( .B(A[70]), .A(S), .Z(O[70]) );
  ANDN U324 ( .B(A[709]), .A(S), .Z(O[709]) );
  ANDN U325 ( .B(A[708]), .A(S), .Z(O[708]) );
  ANDN U326 ( .B(A[707]), .A(S), .Z(O[707]) );
  ANDN U327 ( .B(A[706]), .A(S), .Z(O[706]) );
  ANDN U328 ( .B(A[705]), .A(S), .Z(O[705]) );
  ANDN U329 ( .B(A[704]), .A(S), .Z(O[704]) );
  ANDN U330 ( .B(A[703]), .A(S), .Z(O[703]) );
  ANDN U331 ( .B(A[702]), .A(S), .Z(O[702]) );
  ANDN U332 ( .B(A[701]), .A(S), .Z(O[701]) );
  ANDN U333 ( .B(A[700]), .A(S), .Z(O[700]) );
  ANDN U334 ( .B(A[6]), .A(S), .Z(O[6]) );
  ANDN U335 ( .B(A[69]), .A(S), .Z(O[69]) );
  ANDN U336 ( .B(A[699]), .A(S), .Z(O[699]) );
  ANDN U337 ( .B(A[698]), .A(S), .Z(O[698]) );
  ANDN U338 ( .B(A[697]), .A(S), .Z(O[697]) );
  ANDN U339 ( .B(A[696]), .A(S), .Z(O[696]) );
  ANDN U340 ( .B(A[695]), .A(S), .Z(O[695]) );
  ANDN U341 ( .B(A[694]), .A(S), .Z(O[694]) );
  ANDN U342 ( .B(A[693]), .A(S), .Z(O[693]) );
  ANDN U343 ( .B(A[692]), .A(S), .Z(O[692]) );
  ANDN U344 ( .B(A[691]), .A(S), .Z(O[691]) );
  ANDN U345 ( .B(A[690]), .A(S), .Z(O[690]) );
  ANDN U346 ( .B(A[68]), .A(S), .Z(O[68]) );
  ANDN U347 ( .B(A[689]), .A(S), .Z(O[689]) );
  ANDN U348 ( .B(A[688]), .A(S), .Z(O[688]) );
  ANDN U349 ( .B(A[687]), .A(S), .Z(O[687]) );
  ANDN U350 ( .B(A[686]), .A(S), .Z(O[686]) );
  ANDN U351 ( .B(A[685]), .A(S), .Z(O[685]) );
  ANDN U352 ( .B(A[684]), .A(S), .Z(O[684]) );
  ANDN U353 ( .B(A[683]), .A(S), .Z(O[683]) );
  ANDN U354 ( .B(A[682]), .A(S), .Z(O[682]) );
  ANDN U355 ( .B(A[681]), .A(S), .Z(O[681]) );
  ANDN U356 ( .B(A[680]), .A(S), .Z(O[680]) );
  ANDN U357 ( .B(A[67]), .A(S), .Z(O[67]) );
  ANDN U358 ( .B(A[679]), .A(S), .Z(O[679]) );
  ANDN U359 ( .B(A[678]), .A(S), .Z(O[678]) );
  ANDN U360 ( .B(A[677]), .A(S), .Z(O[677]) );
  ANDN U361 ( .B(A[676]), .A(S), .Z(O[676]) );
  ANDN U362 ( .B(A[675]), .A(S), .Z(O[675]) );
  ANDN U363 ( .B(A[674]), .A(S), .Z(O[674]) );
  ANDN U364 ( .B(A[673]), .A(S), .Z(O[673]) );
  ANDN U365 ( .B(A[672]), .A(S), .Z(O[672]) );
  ANDN U366 ( .B(A[671]), .A(S), .Z(O[671]) );
  ANDN U367 ( .B(A[670]), .A(S), .Z(O[670]) );
  ANDN U368 ( .B(A[66]), .A(S), .Z(O[66]) );
  ANDN U369 ( .B(A[669]), .A(S), .Z(O[669]) );
  ANDN U370 ( .B(A[668]), .A(S), .Z(O[668]) );
  ANDN U371 ( .B(A[667]), .A(S), .Z(O[667]) );
  ANDN U372 ( .B(A[666]), .A(S), .Z(O[666]) );
  ANDN U373 ( .B(A[665]), .A(S), .Z(O[665]) );
  ANDN U374 ( .B(A[664]), .A(S), .Z(O[664]) );
  ANDN U375 ( .B(A[663]), .A(S), .Z(O[663]) );
  ANDN U376 ( .B(A[662]), .A(S), .Z(O[662]) );
  ANDN U377 ( .B(A[661]), .A(S), .Z(O[661]) );
  ANDN U378 ( .B(A[660]), .A(S), .Z(O[660]) );
  ANDN U379 ( .B(A[65]), .A(S), .Z(O[65]) );
  ANDN U380 ( .B(A[659]), .A(S), .Z(O[659]) );
  ANDN U381 ( .B(A[658]), .A(S), .Z(O[658]) );
  ANDN U382 ( .B(A[657]), .A(S), .Z(O[657]) );
  ANDN U383 ( .B(A[656]), .A(S), .Z(O[656]) );
  ANDN U384 ( .B(A[655]), .A(S), .Z(O[655]) );
  ANDN U385 ( .B(A[654]), .A(S), .Z(O[654]) );
  ANDN U386 ( .B(A[653]), .A(S), .Z(O[653]) );
  ANDN U387 ( .B(A[652]), .A(S), .Z(O[652]) );
  ANDN U388 ( .B(A[651]), .A(S), .Z(O[651]) );
  ANDN U389 ( .B(A[650]), .A(S), .Z(O[650]) );
  ANDN U390 ( .B(A[64]), .A(S), .Z(O[64]) );
  ANDN U391 ( .B(A[649]), .A(S), .Z(O[649]) );
  ANDN U392 ( .B(A[648]), .A(S), .Z(O[648]) );
  ANDN U393 ( .B(A[647]), .A(S), .Z(O[647]) );
  ANDN U394 ( .B(A[646]), .A(S), .Z(O[646]) );
  ANDN U395 ( .B(A[645]), .A(S), .Z(O[645]) );
  ANDN U396 ( .B(A[644]), .A(S), .Z(O[644]) );
  ANDN U397 ( .B(A[643]), .A(S), .Z(O[643]) );
  ANDN U398 ( .B(A[642]), .A(S), .Z(O[642]) );
  ANDN U399 ( .B(A[641]), .A(S), .Z(O[641]) );
  ANDN U400 ( .B(A[640]), .A(S), .Z(O[640]) );
  ANDN U401 ( .B(A[63]), .A(S), .Z(O[63]) );
  ANDN U402 ( .B(A[639]), .A(S), .Z(O[639]) );
  ANDN U403 ( .B(A[638]), .A(S), .Z(O[638]) );
  ANDN U404 ( .B(A[637]), .A(S), .Z(O[637]) );
  ANDN U405 ( .B(A[636]), .A(S), .Z(O[636]) );
  ANDN U406 ( .B(A[635]), .A(S), .Z(O[635]) );
  ANDN U407 ( .B(A[634]), .A(S), .Z(O[634]) );
  ANDN U408 ( .B(A[633]), .A(S), .Z(O[633]) );
  ANDN U409 ( .B(A[632]), .A(S), .Z(O[632]) );
  ANDN U410 ( .B(A[631]), .A(S), .Z(O[631]) );
  ANDN U411 ( .B(A[630]), .A(S), .Z(O[630]) );
  ANDN U412 ( .B(A[62]), .A(S), .Z(O[62]) );
  ANDN U413 ( .B(A[629]), .A(S), .Z(O[629]) );
  ANDN U414 ( .B(A[628]), .A(S), .Z(O[628]) );
  ANDN U415 ( .B(A[627]), .A(S), .Z(O[627]) );
  ANDN U416 ( .B(A[626]), .A(S), .Z(O[626]) );
  ANDN U417 ( .B(A[625]), .A(S), .Z(O[625]) );
  ANDN U418 ( .B(A[624]), .A(S), .Z(O[624]) );
  ANDN U419 ( .B(A[623]), .A(S), .Z(O[623]) );
  ANDN U420 ( .B(A[622]), .A(S), .Z(O[622]) );
  ANDN U421 ( .B(A[621]), .A(S), .Z(O[621]) );
  ANDN U422 ( .B(A[620]), .A(S), .Z(O[620]) );
  ANDN U423 ( .B(A[61]), .A(S), .Z(O[61]) );
  ANDN U424 ( .B(A[619]), .A(S), .Z(O[619]) );
  ANDN U425 ( .B(A[618]), .A(S), .Z(O[618]) );
  ANDN U426 ( .B(A[617]), .A(S), .Z(O[617]) );
  ANDN U427 ( .B(A[616]), .A(S), .Z(O[616]) );
  ANDN U428 ( .B(A[615]), .A(S), .Z(O[615]) );
  ANDN U429 ( .B(A[614]), .A(S), .Z(O[614]) );
  ANDN U430 ( .B(A[613]), .A(S), .Z(O[613]) );
  ANDN U431 ( .B(A[612]), .A(S), .Z(O[612]) );
  ANDN U432 ( .B(A[611]), .A(S), .Z(O[611]) );
  ANDN U433 ( .B(A[610]), .A(S), .Z(O[610]) );
  ANDN U434 ( .B(A[60]), .A(S), .Z(O[60]) );
  ANDN U435 ( .B(A[609]), .A(S), .Z(O[609]) );
  ANDN U436 ( .B(A[608]), .A(S), .Z(O[608]) );
  ANDN U437 ( .B(A[607]), .A(S), .Z(O[607]) );
  ANDN U438 ( .B(A[606]), .A(S), .Z(O[606]) );
  ANDN U439 ( .B(A[605]), .A(S), .Z(O[605]) );
  ANDN U440 ( .B(A[604]), .A(S), .Z(O[604]) );
  ANDN U441 ( .B(A[603]), .A(S), .Z(O[603]) );
  ANDN U442 ( .B(A[602]), .A(S), .Z(O[602]) );
  ANDN U443 ( .B(A[601]), .A(S), .Z(O[601]) );
  ANDN U444 ( .B(A[600]), .A(S), .Z(O[600]) );
  ANDN U445 ( .B(A[5]), .A(S), .Z(O[5]) );
  ANDN U446 ( .B(A[59]), .A(S), .Z(O[59]) );
  ANDN U447 ( .B(A[599]), .A(S), .Z(O[599]) );
  ANDN U448 ( .B(A[598]), .A(S), .Z(O[598]) );
  ANDN U449 ( .B(A[597]), .A(S), .Z(O[597]) );
  ANDN U450 ( .B(A[596]), .A(S), .Z(O[596]) );
  ANDN U451 ( .B(A[595]), .A(S), .Z(O[595]) );
  ANDN U452 ( .B(A[594]), .A(S), .Z(O[594]) );
  ANDN U453 ( .B(A[593]), .A(S), .Z(O[593]) );
  ANDN U454 ( .B(A[592]), .A(S), .Z(O[592]) );
  ANDN U455 ( .B(A[591]), .A(S), .Z(O[591]) );
  ANDN U456 ( .B(A[590]), .A(S), .Z(O[590]) );
  ANDN U457 ( .B(A[58]), .A(S), .Z(O[58]) );
  ANDN U458 ( .B(A[589]), .A(S), .Z(O[589]) );
  ANDN U459 ( .B(A[588]), .A(S), .Z(O[588]) );
  ANDN U460 ( .B(A[587]), .A(S), .Z(O[587]) );
  ANDN U461 ( .B(A[586]), .A(S), .Z(O[586]) );
  ANDN U462 ( .B(A[585]), .A(S), .Z(O[585]) );
  ANDN U463 ( .B(A[584]), .A(S), .Z(O[584]) );
  ANDN U464 ( .B(A[583]), .A(S), .Z(O[583]) );
  ANDN U465 ( .B(A[582]), .A(S), .Z(O[582]) );
  ANDN U466 ( .B(A[581]), .A(S), .Z(O[581]) );
  ANDN U467 ( .B(A[580]), .A(S), .Z(O[580]) );
  ANDN U468 ( .B(A[57]), .A(S), .Z(O[57]) );
  ANDN U469 ( .B(A[579]), .A(S), .Z(O[579]) );
  ANDN U470 ( .B(A[578]), .A(S), .Z(O[578]) );
  ANDN U471 ( .B(A[577]), .A(S), .Z(O[577]) );
  ANDN U472 ( .B(A[576]), .A(S), .Z(O[576]) );
  ANDN U473 ( .B(A[575]), .A(S), .Z(O[575]) );
  ANDN U474 ( .B(A[574]), .A(S), .Z(O[574]) );
  ANDN U475 ( .B(A[573]), .A(S), .Z(O[573]) );
  ANDN U476 ( .B(A[572]), .A(S), .Z(O[572]) );
  ANDN U477 ( .B(A[571]), .A(S), .Z(O[571]) );
  ANDN U478 ( .B(A[570]), .A(S), .Z(O[570]) );
  ANDN U479 ( .B(A[56]), .A(S), .Z(O[56]) );
  ANDN U480 ( .B(A[569]), .A(S), .Z(O[569]) );
  ANDN U481 ( .B(A[568]), .A(S), .Z(O[568]) );
  ANDN U482 ( .B(A[567]), .A(S), .Z(O[567]) );
  ANDN U483 ( .B(A[566]), .A(S), .Z(O[566]) );
  ANDN U484 ( .B(A[565]), .A(S), .Z(O[565]) );
  ANDN U485 ( .B(A[564]), .A(S), .Z(O[564]) );
  ANDN U486 ( .B(A[563]), .A(S), .Z(O[563]) );
  ANDN U487 ( .B(A[562]), .A(S), .Z(O[562]) );
  ANDN U488 ( .B(A[561]), .A(S), .Z(O[561]) );
  ANDN U489 ( .B(A[560]), .A(S), .Z(O[560]) );
  ANDN U490 ( .B(A[55]), .A(S), .Z(O[55]) );
  ANDN U491 ( .B(A[559]), .A(S), .Z(O[559]) );
  ANDN U492 ( .B(A[558]), .A(S), .Z(O[558]) );
  ANDN U493 ( .B(A[557]), .A(S), .Z(O[557]) );
  ANDN U494 ( .B(A[556]), .A(S), .Z(O[556]) );
  ANDN U495 ( .B(A[555]), .A(S), .Z(O[555]) );
  ANDN U496 ( .B(A[554]), .A(S), .Z(O[554]) );
  ANDN U497 ( .B(A[553]), .A(S), .Z(O[553]) );
  ANDN U498 ( .B(A[552]), .A(S), .Z(O[552]) );
  ANDN U499 ( .B(A[551]), .A(S), .Z(O[551]) );
  ANDN U500 ( .B(A[550]), .A(S), .Z(O[550]) );
  ANDN U501 ( .B(A[54]), .A(S), .Z(O[54]) );
  ANDN U502 ( .B(A[549]), .A(S), .Z(O[549]) );
  ANDN U503 ( .B(A[548]), .A(S), .Z(O[548]) );
  ANDN U504 ( .B(A[547]), .A(S), .Z(O[547]) );
  ANDN U505 ( .B(A[546]), .A(S), .Z(O[546]) );
  ANDN U506 ( .B(A[545]), .A(S), .Z(O[545]) );
  ANDN U507 ( .B(A[544]), .A(S), .Z(O[544]) );
  ANDN U508 ( .B(A[543]), .A(S), .Z(O[543]) );
  ANDN U509 ( .B(A[542]), .A(S), .Z(O[542]) );
  ANDN U510 ( .B(A[541]), .A(S), .Z(O[541]) );
  ANDN U511 ( .B(A[540]), .A(S), .Z(O[540]) );
  ANDN U512 ( .B(A[53]), .A(S), .Z(O[53]) );
  ANDN U513 ( .B(A[539]), .A(S), .Z(O[539]) );
  ANDN U514 ( .B(A[538]), .A(S), .Z(O[538]) );
  ANDN U515 ( .B(A[537]), .A(S), .Z(O[537]) );
  ANDN U516 ( .B(A[536]), .A(S), .Z(O[536]) );
  ANDN U517 ( .B(A[535]), .A(S), .Z(O[535]) );
  ANDN U518 ( .B(A[534]), .A(S), .Z(O[534]) );
  ANDN U519 ( .B(A[533]), .A(S), .Z(O[533]) );
  ANDN U520 ( .B(A[532]), .A(S), .Z(O[532]) );
  ANDN U521 ( .B(A[531]), .A(S), .Z(O[531]) );
  ANDN U522 ( .B(A[530]), .A(S), .Z(O[530]) );
  ANDN U523 ( .B(A[52]), .A(S), .Z(O[52]) );
  ANDN U524 ( .B(A[529]), .A(S), .Z(O[529]) );
  ANDN U525 ( .B(A[528]), .A(S), .Z(O[528]) );
  ANDN U526 ( .B(A[527]), .A(S), .Z(O[527]) );
  ANDN U527 ( .B(A[526]), .A(S), .Z(O[526]) );
  ANDN U528 ( .B(A[525]), .A(S), .Z(O[525]) );
  ANDN U529 ( .B(A[524]), .A(S), .Z(O[524]) );
  ANDN U530 ( .B(A[523]), .A(S), .Z(O[523]) );
  ANDN U531 ( .B(A[522]), .A(S), .Z(O[522]) );
  ANDN U532 ( .B(A[521]), .A(S), .Z(O[521]) );
  ANDN U533 ( .B(A[520]), .A(S), .Z(O[520]) );
  ANDN U534 ( .B(A[51]), .A(S), .Z(O[51]) );
  ANDN U535 ( .B(A[519]), .A(S), .Z(O[519]) );
  ANDN U536 ( .B(A[518]), .A(S), .Z(O[518]) );
  ANDN U537 ( .B(A[517]), .A(S), .Z(O[517]) );
  ANDN U538 ( .B(A[516]), .A(S), .Z(O[516]) );
  ANDN U539 ( .B(A[515]), .A(S), .Z(O[515]) );
  ANDN U540 ( .B(A[514]), .A(S), .Z(O[514]) );
  ANDN U541 ( .B(A[513]), .A(S), .Z(O[513]) );
  ANDN U542 ( .B(A[512]), .A(S), .Z(O[512]) );
  ANDN U543 ( .B(A[511]), .A(S), .Z(O[511]) );
  ANDN U544 ( .B(A[510]), .A(S), .Z(O[510]) );
  ANDN U545 ( .B(A[50]), .A(S), .Z(O[50]) );
  ANDN U546 ( .B(A[509]), .A(S), .Z(O[509]) );
  ANDN U547 ( .B(A[508]), .A(S), .Z(O[508]) );
  ANDN U548 ( .B(A[507]), .A(S), .Z(O[507]) );
  ANDN U549 ( .B(A[506]), .A(S), .Z(O[506]) );
  ANDN U550 ( .B(A[505]), .A(S), .Z(O[505]) );
  ANDN U551 ( .B(A[504]), .A(S), .Z(O[504]) );
  ANDN U552 ( .B(A[503]), .A(S), .Z(O[503]) );
  ANDN U553 ( .B(A[502]), .A(S), .Z(O[502]) );
  ANDN U554 ( .B(A[501]), .A(S), .Z(O[501]) );
  ANDN U555 ( .B(A[500]), .A(S), .Z(O[500]) );
  ANDN U556 ( .B(A[4]), .A(S), .Z(O[4]) );
  ANDN U557 ( .B(A[49]), .A(S), .Z(O[49]) );
  ANDN U558 ( .B(A[499]), .A(S), .Z(O[499]) );
  ANDN U559 ( .B(A[498]), .A(S), .Z(O[498]) );
  ANDN U560 ( .B(A[497]), .A(S), .Z(O[497]) );
  ANDN U561 ( .B(A[496]), .A(S), .Z(O[496]) );
  ANDN U562 ( .B(A[495]), .A(S), .Z(O[495]) );
  ANDN U563 ( .B(A[494]), .A(S), .Z(O[494]) );
  ANDN U564 ( .B(A[493]), .A(S), .Z(O[493]) );
  ANDN U565 ( .B(A[492]), .A(S), .Z(O[492]) );
  ANDN U566 ( .B(A[491]), .A(S), .Z(O[491]) );
  ANDN U567 ( .B(A[490]), .A(S), .Z(O[490]) );
  ANDN U568 ( .B(A[48]), .A(S), .Z(O[48]) );
  ANDN U569 ( .B(A[489]), .A(S), .Z(O[489]) );
  ANDN U570 ( .B(A[488]), .A(S), .Z(O[488]) );
  ANDN U571 ( .B(A[487]), .A(S), .Z(O[487]) );
  ANDN U572 ( .B(A[486]), .A(S), .Z(O[486]) );
  ANDN U573 ( .B(A[485]), .A(S), .Z(O[485]) );
  ANDN U574 ( .B(A[484]), .A(S), .Z(O[484]) );
  ANDN U575 ( .B(A[483]), .A(S), .Z(O[483]) );
  ANDN U576 ( .B(A[482]), .A(S), .Z(O[482]) );
  ANDN U577 ( .B(A[481]), .A(S), .Z(O[481]) );
  ANDN U578 ( .B(A[480]), .A(S), .Z(O[480]) );
  ANDN U579 ( .B(A[47]), .A(S), .Z(O[47]) );
  ANDN U580 ( .B(A[479]), .A(S), .Z(O[479]) );
  ANDN U581 ( .B(A[478]), .A(S), .Z(O[478]) );
  ANDN U582 ( .B(A[477]), .A(S), .Z(O[477]) );
  ANDN U583 ( .B(A[476]), .A(S), .Z(O[476]) );
  ANDN U584 ( .B(A[475]), .A(S), .Z(O[475]) );
  ANDN U585 ( .B(A[474]), .A(S), .Z(O[474]) );
  ANDN U586 ( .B(A[473]), .A(S), .Z(O[473]) );
  ANDN U587 ( .B(A[472]), .A(S), .Z(O[472]) );
  ANDN U588 ( .B(A[471]), .A(S), .Z(O[471]) );
  ANDN U589 ( .B(A[470]), .A(S), .Z(O[470]) );
  ANDN U590 ( .B(A[46]), .A(S), .Z(O[46]) );
  ANDN U591 ( .B(A[469]), .A(S), .Z(O[469]) );
  ANDN U592 ( .B(A[468]), .A(S), .Z(O[468]) );
  ANDN U593 ( .B(A[467]), .A(S), .Z(O[467]) );
  ANDN U594 ( .B(A[466]), .A(S), .Z(O[466]) );
  ANDN U595 ( .B(A[465]), .A(S), .Z(O[465]) );
  ANDN U596 ( .B(A[464]), .A(S), .Z(O[464]) );
  ANDN U597 ( .B(A[463]), .A(S), .Z(O[463]) );
  ANDN U598 ( .B(A[462]), .A(S), .Z(O[462]) );
  ANDN U599 ( .B(A[461]), .A(S), .Z(O[461]) );
  ANDN U600 ( .B(A[460]), .A(S), .Z(O[460]) );
  ANDN U601 ( .B(A[45]), .A(S), .Z(O[45]) );
  ANDN U602 ( .B(A[459]), .A(S), .Z(O[459]) );
  ANDN U603 ( .B(A[458]), .A(S), .Z(O[458]) );
  ANDN U604 ( .B(A[457]), .A(S), .Z(O[457]) );
  ANDN U605 ( .B(A[456]), .A(S), .Z(O[456]) );
  ANDN U606 ( .B(A[455]), .A(S), .Z(O[455]) );
  ANDN U607 ( .B(A[454]), .A(S), .Z(O[454]) );
  ANDN U608 ( .B(A[453]), .A(S), .Z(O[453]) );
  ANDN U609 ( .B(A[452]), .A(S), .Z(O[452]) );
  ANDN U610 ( .B(A[451]), .A(S), .Z(O[451]) );
  ANDN U611 ( .B(A[450]), .A(S), .Z(O[450]) );
  ANDN U612 ( .B(A[44]), .A(S), .Z(O[44]) );
  ANDN U613 ( .B(A[449]), .A(S), .Z(O[449]) );
  ANDN U614 ( .B(A[448]), .A(S), .Z(O[448]) );
  ANDN U615 ( .B(A[447]), .A(S), .Z(O[447]) );
  ANDN U616 ( .B(A[446]), .A(S), .Z(O[446]) );
  ANDN U617 ( .B(A[445]), .A(S), .Z(O[445]) );
  ANDN U618 ( .B(A[444]), .A(S), .Z(O[444]) );
  ANDN U619 ( .B(A[443]), .A(S), .Z(O[443]) );
  ANDN U620 ( .B(A[442]), .A(S), .Z(O[442]) );
  ANDN U621 ( .B(A[441]), .A(S), .Z(O[441]) );
  ANDN U622 ( .B(A[440]), .A(S), .Z(O[440]) );
  ANDN U623 ( .B(A[43]), .A(S), .Z(O[43]) );
  ANDN U624 ( .B(A[439]), .A(S), .Z(O[439]) );
  ANDN U625 ( .B(A[438]), .A(S), .Z(O[438]) );
  ANDN U626 ( .B(A[437]), .A(S), .Z(O[437]) );
  ANDN U627 ( .B(A[436]), .A(S), .Z(O[436]) );
  ANDN U628 ( .B(A[435]), .A(S), .Z(O[435]) );
  ANDN U629 ( .B(A[434]), .A(S), .Z(O[434]) );
  ANDN U630 ( .B(A[433]), .A(S), .Z(O[433]) );
  ANDN U631 ( .B(A[432]), .A(S), .Z(O[432]) );
  ANDN U632 ( .B(A[431]), .A(S), .Z(O[431]) );
  ANDN U633 ( .B(A[430]), .A(S), .Z(O[430]) );
  ANDN U634 ( .B(A[42]), .A(S), .Z(O[42]) );
  ANDN U635 ( .B(A[429]), .A(S), .Z(O[429]) );
  ANDN U636 ( .B(A[428]), .A(S), .Z(O[428]) );
  ANDN U637 ( .B(A[427]), .A(S), .Z(O[427]) );
  ANDN U638 ( .B(A[426]), .A(S), .Z(O[426]) );
  ANDN U639 ( .B(A[425]), .A(S), .Z(O[425]) );
  ANDN U640 ( .B(A[424]), .A(S), .Z(O[424]) );
  ANDN U641 ( .B(A[423]), .A(S), .Z(O[423]) );
  ANDN U642 ( .B(A[422]), .A(S), .Z(O[422]) );
  ANDN U643 ( .B(A[421]), .A(S), .Z(O[421]) );
  ANDN U644 ( .B(A[420]), .A(S), .Z(O[420]) );
  ANDN U645 ( .B(A[41]), .A(S), .Z(O[41]) );
  ANDN U646 ( .B(A[419]), .A(S), .Z(O[419]) );
  ANDN U647 ( .B(A[418]), .A(S), .Z(O[418]) );
  ANDN U648 ( .B(A[417]), .A(S), .Z(O[417]) );
  ANDN U649 ( .B(A[416]), .A(S), .Z(O[416]) );
  ANDN U650 ( .B(A[415]), .A(S), .Z(O[415]) );
  ANDN U651 ( .B(A[414]), .A(S), .Z(O[414]) );
  ANDN U652 ( .B(A[413]), .A(S), .Z(O[413]) );
  ANDN U653 ( .B(A[412]), .A(S), .Z(O[412]) );
  ANDN U654 ( .B(A[411]), .A(S), .Z(O[411]) );
  ANDN U655 ( .B(A[410]), .A(S), .Z(O[410]) );
  ANDN U656 ( .B(A[40]), .A(S), .Z(O[40]) );
  ANDN U657 ( .B(A[409]), .A(S), .Z(O[409]) );
  ANDN U658 ( .B(A[408]), .A(S), .Z(O[408]) );
  ANDN U659 ( .B(A[407]), .A(S), .Z(O[407]) );
  ANDN U660 ( .B(A[406]), .A(S), .Z(O[406]) );
  ANDN U661 ( .B(A[405]), .A(S), .Z(O[405]) );
  ANDN U662 ( .B(A[404]), .A(S), .Z(O[404]) );
  ANDN U663 ( .B(A[403]), .A(S), .Z(O[403]) );
  ANDN U664 ( .B(A[402]), .A(S), .Z(O[402]) );
  ANDN U665 ( .B(A[401]), .A(S), .Z(O[401]) );
  ANDN U666 ( .B(A[400]), .A(S), .Z(O[400]) );
  ANDN U667 ( .B(A[3]), .A(S), .Z(O[3]) );
  ANDN U668 ( .B(A[39]), .A(S), .Z(O[39]) );
  ANDN U669 ( .B(A[399]), .A(S), .Z(O[399]) );
  ANDN U670 ( .B(A[398]), .A(S), .Z(O[398]) );
  ANDN U671 ( .B(A[397]), .A(S), .Z(O[397]) );
  ANDN U672 ( .B(A[396]), .A(S), .Z(O[396]) );
  ANDN U673 ( .B(A[395]), .A(S), .Z(O[395]) );
  ANDN U674 ( .B(A[394]), .A(S), .Z(O[394]) );
  ANDN U675 ( .B(A[393]), .A(S), .Z(O[393]) );
  ANDN U676 ( .B(A[392]), .A(S), .Z(O[392]) );
  ANDN U677 ( .B(A[391]), .A(S), .Z(O[391]) );
  ANDN U678 ( .B(A[390]), .A(S), .Z(O[390]) );
  ANDN U679 ( .B(A[38]), .A(S), .Z(O[38]) );
  ANDN U680 ( .B(A[389]), .A(S), .Z(O[389]) );
  ANDN U681 ( .B(A[388]), .A(S), .Z(O[388]) );
  ANDN U682 ( .B(A[387]), .A(S), .Z(O[387]) );
  ANDN U683 ( .B(A[386]), .A(S), .Z(O[386]) );
  ANDN U684 ( .B(A[385]), .A(S), .Z(O[385]) );
  ANDN U685 ( .B(A[384]), .A(S), .Z(O[384]) );
  ANDN U686 ( .B(A[383]), .A(S), .Z(O[383]) );
  ANDN U687 ( .B(A[382]), .A(S), .Z(O[382]) );
  ANDN U688 ( .B(A[381]), .A(S), .Z(O[381]) );
  ANDN U689 ( .B(A[380]), .A(S), .Z(O[380]) );
  ANDN U690 ( .B(A[37]), .A(S), .Z(O[37]) );
  ANDN U691 ( .B(A[379]), .A(S), .Z(O[379]) );
  ANDN U692 ( .B(A[378]), .A(S), .Z(O[378]) );
  ANDN U693 ( .B(A[377]), .A(S), .Z(O[377]) );
  ANDN U694 ( .B(A[376]), .A(S), .Z(O[376]) );
  ANDN U695 ( .B(A[375]), .A(S), .Z(O[375]) );
  ANDN U696 ( .B(A[374]), .A(S), .Z(O[374]) );
  ANDN U697 ( .B(A[373]), .A(S), .Z(O[373]) );
  ANDN U698 ( .B(A[372]), .A(S), .Z(O[372]) );
  ANDN U699 ( .B(A[371]), .A(S), .Z(O[371]) );
  ANDN U700 ( .B(A[370]), .A(S), .Z(O[370]) );
  ANDN U701 ( .B(A[36]), .A(S), .Z(O[36]) );
  ANDN U702 ( .B(A[369]), .A(S), .Z(O[369]) );
  ANDN U703 ( .B(A[368]), .A(S), .Z(O[368]) );
  ANDN U704 ( .B(A[367]), .A(S), .Z(O[367]) );
  ANDN U705 ( .B(A[366]), .A(S), .Z(O[366]) );
  ANDN U706 ( .B(A[365]), .A(S), .Z(O[365]) );
  ANDN U707 ( .B(A[364]), .A(S), .Z(O[364]) );
  ANDN U708 ( .B(A[363]), .A(S), .Z(O[363]) );
  ANDN U709 ( .B(A[362]), .A(S), .Z(O[362]) );
  ANDN U710 ( .B(A[361]), .A(S), .Z(O[361]) );
  ANDN U711 ( .B(A[360]), .A(S), .Z(O[360]) );
  ANDN U712 ( .B(A[35]), .A(S), .Z(O[35]) );
  ANDN U713 ( .B(A[359]), .A(S), .Z(O[359]) );
  ANDN U714 ( .B(A[358]), .A(S), .Z(O[358]) );
  ANDN U715 ( .B(A[357]), .A(S), .Z(O[357]) );
  ANDN U716 ( .B(A[356]), .A(S), .Z(O[356]) );
  ANDN U717 ( .B(A[355]), .A(S), .Z(O[355]) );
  ANDN U718 ( .B(A[354]), .A(S), .Z(O[354]) );
  ANDN U719 ( .B(A[353]), .A(S), .Z(O[353]) );
  ANDN U720 ( .B(A[352]), .A(S), .Z(O[352]) );
  ANDN U721 ( .B(A[351]), .A(S), .Z(O[351]) );
  ANDN U722 ( .B(A[350]), .A(S), .Z(O[350]) );
  ANDN U723 ( .B(A[34]), .A(S), .Z(O[34]) );
  ANDN U724 ( .B(A[349]), .A(S), .Z(O[349]) );
  ANDN U725 ( .B(A[348]), .A(S), .Z(O[348]) );
  ANDN U726 ( .B(A[347]), .A(S), .Z(O[347]) );
  ANDN U727 ( .B(A[346]), .A(S), .Z(O[346]) );
  ANDN U728 ( .B(A[345]), .A(S), .Z(O[345]) );
  ANDN U729 ( .B(A[344]), .A(S), .Z(O[344]) );
  ANDN U730 ( .B(A[343]), .A(S), .Z(O[343]) );
  ANDN U731 ( .B(A[342]), .A(S), .Z(O[342]) );
  ANDN U732 ( .B(A[341]), .A(S), .Z(O[341]) );
  ANDN U733 ( .B(A[340]), .A(S), .Z(O[340]) );
  ANDN U734 ( .B(A[33]), .A(S), .Z(O[33]) );
  ANDN U735 ( .B(A[339]), .A(S), .Z(O[339]) );
  ANDN U736 ( .B(A[338]), .A(S), .Z(O[338]) );
  ANDN U737 ( .B(A[337]), .A(S), .Z(O[337]) );
  ANDN U738 ( .B(A[336]), .A(S), .Z(O[336]) );
  ANDN U739 ( .B(A[335]), .A(S), .Z(O[335]) );
  ANDN U740 ( .B(A[334]), .A(S), .Z(O[334]) );
  ANDN U741 ( .B(A[333]), .A(S), .Z(O[333]) );
  ANDN U742 ( .B(A[332]), .A(S), .Z(O[332]) );
  ANDN U743 ( .B(A[331]), .A(S), .Z(O[331]) );
  ANDN U744 ( .B(A[330]), .A(S), .Z(O[330]) );
  ANDN U745 ( .B(A[32]), .A(S), .Z(O[32]) );
  ANDN U746 ( .B(A[329]), .A(S), .Z(O[329]) );
  ANDN U747 ( .B(A[328]), .A(S), .Z(O[328]) );
  ANDN U748 ( .B(A[327]), .A(S), .Z(O[327]) );
  ANDN U749 ( .B(A[326]), .A(S), .Z(O[326]) );
  ANDN U750 ( .B(A[325]), .A(S), .Z(O[325]) );
  ANDN U751 ( .B(A[324]), .A(S), .Z(O[324]) );
  ANDN U752 ( .B(A[323]), .A(S), .Z(O[323]) );
  ANDN U753 ( .B(A[322]), .A(S), .Z(O[322]) );
  ANDN U754 ( .B(A[321]), .A(S), .Z(O[321]) );
  ANDN U755 ( .B(A[320]), .A(S), .Z(O[320]) );
  ANDN U756 ( .B(A[31]), .A(S), .Z(O[31]) );
  ANDN U757 ( .B(A[319]), .A(S), .Z(O[319]) );
  ANDN U758 ( .B(A[318]), .A(S), .Z(O[318]) );
  ANDN U759 ( .B(A[317]), .A(S), .Z(O[317]) );
  ANDN U760 ( .B(A[316]), .A(S), .Z(O[316]) );
  ANDN U761 ( .B(A[315]), .A(S), .Z(O[315]) );
  ANDN U762 ( .B(A[314]), .A(S), .Z(O[314]) );
  ANDN U763 ( .B(A[313]), .A(S), .Z(O[313]) );
  ANDN U764 ( .B(A[312]), .A(S), .Z(O[312]) );
  ANDN U765 ( .B(A[311]), .A(S), .Z(O[311]) );
  ANDN U766 ( .B(A[310]), .A(S), .Z(O[310]) );
  ANDN U767 ( .B(A[30]), .A(S), .Z(O[30]) );
  ANDN U768 ( .B(A[309]), .A(S), .Z(O[309]) );
  ANDN U769 ( .B(A[308]), .A(S), .Z(O[308]) );
  ANDN U770 ( .B(A[307]), .A(S), .Z(O[307]) );
  ANDN U771 ( .B(A[306]), .A(S), .Z(O[306]) );
  ANDN U772 ( .B(A[305]), .A(S), .Z(O[305]) );
  ANDN U773 ( .B(A[304]), .A(S), .Z(O[304]) );
  ANDN U774 ( .B(A[303]), .A(S), .Z(O[303]) );
  ANDN U775 ( .B(A[302]), .A(S), .Z(O[302]) );
  ANDN U776 ( .B(A[301]), .A(S), .Z(O[301]) );
  ANDN U777 ( .B(A[300]), .A(S), .Z(O[300]) );
  ANDN U778 ( .B(A[2]), .A(S), .Z(O[2]) );
  ANDN U779 ( .B(A[29]), .A(S), .Z(O[29]) );
  ANDN U780 ( .B(A[299]), .A(S), .Z(O[299]) );
  ANDN U781 ( .B(A[298]), .A(S), .Z(O[298]) );
  ANDN U782 ( .B(A[297]), .A(S), .Z(O[297]) );
  ANDN U783 ( .B(A[296]), .A(S), .Z(O[296]) );
  ANDN U784 ( .B(A[295]), .A(S), .Z(O[295]) );
  ANDN U785 ( .B(A[294]), .A(S), .Z(O[294]) );
  ANDN U786 ( .B(A[293]), .A(S), .Z(O[293]) );
  ANDN U787 ( .B(A[292]), .A(S), .Z(O[292]) );
  ANDN U788 ( .B(A[291]), .A(S), .Z(O[291]) );
  ANDN U789 ( .B(A[290]), .A(S), .Z(O[290]) );
  ANDN U790 ( .B(A[28]), .A(S), .Z(O[28]) );
  ANDN U791 ( .B(A[289]), .A(S), .Z(O[289]) );
  ANDN U792 ( .B(A[288]), .A(S), .Z(O[288]) );
  ANDN U793 ( .B(A[287]), .A(S), .Z(O[287]) );
  ANDN U794 ( .B(A[286]), .A(S), .Z(O[286]) );
  ANDN U795 ( .B(A[285]), .A(S), .Z(O[285]) );
  ANDN U796 ( .B(A[284]), .A(S), .Z(O[284]) );
  ANDN U797 ( .B(A[283]), .A(S), .Z(O[283]) );
  ANDN U798 ( .B(A[282]), .A(S), .Z(O[282]) );
  ANDN U799 ( .B(A[281]), .A(S), .Z(O[281]) );
  ANDN U800 ( .B(A[280]), .A(S), .Z(O[280]) );
  ANDN U801 ( .B(A[27]), .A(S), .Z(O[27]) );
  ANDN U802 ( .B(A[279]), .A(S), .Z(O[279]) );
  ANDN U803 ( .B(A[278]), .A(S), .Z(O[278]) );
  ANDN U804 ( .B(A[277]), .A(S), .Z(O[277]) );
  ANDN U805 ( .B(A[276]), .A(S), .Z(O[276]) );
  ANDN U806 ( .B(A[275]), .A(S), .Z(O[275]) );
  ANDN U807 ( .B(A[274]), .A(S), .Z(O[274]) );
  ANDN U808 ( .B(A[273]), .A(S), .Z(O[273]) );
  ANDN U809 ( .B(A[272]), .A(S), .Z(O[272]) );
  ANDN U810 ( .B(A[271]), .A(S), .Z(O[271]) );
  ANDN U811 ( .B(A[270]), .A(S), .Z(O[270]) );
  ANDN U812 ( .B(A[26]), .A(S), .Z(O[26]) );
  ANDN U813 ( .B(A[269]), .A(S), .Z(O[269]) );
  ANDN U814 ( .B(A[268]), .A(S), .Z(O[268]) );
  ANDN U815 ( .B(A[267]), .A(S), .Z(O[267]) );
  ANDN U816 ( .B(A[266]), .A(S), .Z(O[266]) );
  ANDN U817 ( .B(A[265]), .A(S), .Z(O[265]) );
  ANDN U818 ( .B(A[264]), .A(S), .Z(O[264]) );
  ANDN U819 ( .B(A[263]), .A(S), .Z(O[263]) );
  ANDN U820 ( .B(A[262]), .A(S), .Z(O[262]) );
  ANDN U821 ( .B(A[261]), .A(S), .Z(O[261]) );
  ANDN U822 ( .B(A[260]), .A(S), .Z(O[260]) );
  ANDN U823 ( .B(A[25]), .A(S), .Z(O[25]) );
  ANDN U824 ( .B(A[259]), .A(S), .Z(O[259]) );
  ANDN U825 ( .B(A[258]), .A(S), .Z(O[258]) );
  ANDN U826 ( .B(A[257]), .A(S), .Z(O[257]) );
  ANDN U827 ( .B(A[256]), .A(S), .Z(O[256]) );
  ANDN U828 ( .B(A[255]), .A(S), .Z(O[255]) );
  ANDN U829 ( .B(A[254]), .A(S), .Z(O[254]) );
  ANDN U830 ( .B(A[253]), .A(S), .Z(O[253]) );
  ANDN U831 ( .B(A[252]), .A(S), .Z(O[252]) );
  ANDN U832 ( .B(A[251]), .A(S), .Z(O[251]) );
  ANDN U833 ( .B(A[250]), .A(S), .Z(O[250]) );
  ANDN U834 ( .B(A[24]), .A(S), .Z(O[24]) );
  ANDN U835 ( .B(A[249]), .A(S), .Z(O[249]) );
  ANDN U836 ( .B(A[248]), .A(S), .Z(O[248]) );
  ANDN U837 ( .B(A[247]), .A(S), .Z(O[247]) );
  ANDN U838 ( .B(A[246]), .A(S), .Z(O[246]) );
  ANDN U839 ( .B(A[245]), .A(S), .Z(O[245]) );
  ANDN U840 ( .B(A[244]), .A(S), .Z(O[244]) );
  ANDN U841 ( .B(A[243]), .A(S), .Z(O[243]) );
  ANDN U842 ( .B(A[242]), .A(S), .Z(O[242]) );
  ANDN U843 ( .B(A[241]), .A(S), .Z(O[241]) );
  ANDN U844 ( .B(A[240]), .A(S), .Z(O[240]) );
  ANDN U845 ( .B(A[23]), .A(S), .Z(O[23]) );
  ANDN U846 ( .B(A[239]), .A(S), .Z(O[239]) );
  ANDN U847 ( .B(A[238]), .A(S), .Z(O[238]) );
  ANDN U848 ( .B(A[237]), .A(S), .Z(O[237]) );
  ANDN U849 ( .B(A[236]), .A(S), .Z(O[236]) );
  ANDN U850 ( .B(A[235]), .A(S), .Z(O[235]) );
  ANDN U851 ( .B(A[234]), .A(S), .Z(O[234]) );
  ANDN U852 ( .B(A[233]), .A(S), .Z(O[233]) );
  ANDN U853 ( .B(A[232]), .A(S), .Z(O[232]) );
  ANDN U854 ( .B(A[231]), .A(S), .Z(O[231]) );
  ANDN U855 ( .B(A[230]), .A(S), .Z(O[230]) );
  ANDN U856 ( .B(A[22]), .A(S), .Z(O[22]) );
  ANDN U857 ( .B(A[229]), .A(S), .Z(O[229]) );
  ANDN U858 ( .B(A[228]), .A(S), .Z(O[228]) );
  ANDN U859 ( .B(A[227]), .A(S), .Z(O[227]) );
  ANDN U860 ( .B(A[226]), .A(S), .Z(O[226]) );
  ANDN U861 ( .B(A[225]), .A(S), .Z(O[225]) );
  ANDN U862 ( .B(A[224]), .A(S), .Z(O[224]) );
  ANDN U863 ( .B(A[223]), .A(S), .Z(O[223]) );
  ANDN U864 ( .B(A[222]), .A(S), .Z(O[222]) );
  ANDN U865 ( .B(A[221]), .A(S), .Z(O[221]) );
  ANDN U866 ( .B(A[220]), .A(S), .Z(O[220]) );
  ANDN U867 ( .B(A[21]), .A(S), .Z(O[21]) );
  ANDN U868 ( .B(A[219]), .A(S), .Z(O[219]) );
  ANDN U869 ( .B(A[218]), .A(S), .Z(O[218]) );
  ANDN U870 ( .B(A[217]), .A(S), .Z(O[217]) );
  ANDN U871 ( .B(A[216]), .A(S), .Z(O[216]) );
  ANDN U872 ( .B(A[215]), .A(S), .Z(O[215]) );
  ANDN U873 ( .B(A[214]), .A(S), .Z(O[214]) );
  ANDN U874 ( .B(A[213]), .A(S), .Z(O[213]) );
  ANDN U875 ( .B(A[212]), .A(S), .Z(O[212]) );
  ANDN U876 ( .B(A[211]), .A(S), .Z(O[211]) );
  ANDN U877 ( .B(A[210]), .A(S), .Z(O[210]) );
  ANDN U878 ( .B(A[20]), .A(S), .Z(O[20]) );
  ANDN U879 ( .B(A[209]), .A(S), .Z(O[209]) );
  ANDN U880 ( .B(A[208]), .A(S), .Z(O[208]) );
  ANDN U881 ( .B(A[207]), .A(S), .Z(O[207]) );
  ANDN U882 ( .B(A[206]), .A(S), .Z(O[206]) );
  ANDN U883 ( .B(A[205]), .A(S), .Z(O[205]) );
  ANDN U884 ( .B(A[204]), .A(S), .Z(O[204]) );
  ANDN U885 ( .B(A[203]), .A(S), .Z(O[203]) );
  ANDN U886 ( .B(A[202]), .A(S), .Z(O[202]) );
  ANDN U887 ( .B(A[201]), .A(S), .Z(O[201]) );
  ANDN U888 ( .B(A[200]), .A(S), .Z(O[200]) );
  ANDN U889 ( .B(A[1]), .A(S), .Z(O[1]) );
  ANDN U890 ( .B(A[19]), .A(S), .Z(O[19]) );
  ANDN U891 ( .B(A[199]), .A(S), .Z(O[199]) );
  ANDN U892 ( .B(A[198]), .A(S), .Z(O[198]) );
  ANDN U893 ( .B(A[197]), .A(S), .Z(O[197]) );
  ANDN U894 ( .B(A[196]), .A(S), .Z(O[196]) );
  ANDN U895 ( .B(A[195]), .A(S), .Z(O[195]) );
  ANDN U896 ( .B(A[194]), .A(S), .Z(O[194]) );
  ANDN U897 ( .B(A[193]), .A(S), .Z(O[193]) );
  ANDN U898 ( .B(A[192]), .A(S), .Z(O[192]) );
  ANDN U899 ( .B(A[191]), .A(S), .Z(O[191]) );
  ANDN U900 ( .B(A[190]), .A(S), .Z(O[190]) );
  ANDN U901 ( .B(A[18]), .A(S), .Z(O[18]) );
  ANDN U902 ( .B(A[189]), .A(S), .Z(O[189]) );
  ANDN U903 ( .B(A[188]), .A(S), .Z(O[188]) );
  ANDN U904 ( .B(A[187]), .A(S), .Z(O[187]) );
  ANDN U905 ( .B(A[186]), .A(S), .Z(O[186]) );
  ANDN U906 ( .B(A[185]), .A(S), .Z(O[185]) );
  ANDN U907 ( .B(A[184]), .A(S), .Z(O[184]) );
  ANDN U908 ( .B(A[183]), .A(S), .Z(O[183]) );
  ANDN U909 ( .B(A[182]), .A(S), .Z(O[182]) );
  ANDN U910 ( .B(A[181]), .A(S), .Z(O[181]) );
  ANDN U911 ( .B(A[180]), .A(S), .Z(O[180]) );
  ANDN U912 ( .B(A[17]), .A(S), .Z(O[17]) );
  ANDN U913 ( .B(A[179]), .A(S), .Z(O[179]) );
  ANDN U914 ( .B(A[178]), .A(S), .Z(O[178]) );
  ANDN U915 ( .B(A[177]), .A(S), .Z(O[177]) );
  ANDN U916 ( .B(A[176]), .A(S), .Z(O[176]) );
  ANDN U917 ( .B(A[175]), .A(S), .Z(O[175]) );
  ANDN U918 ( .B(A[174]), .A(S), .Z(O[174]) );
  ANDN U919 ( .B(A[173]), .A(S), .Z(O[173]) );
  ANDN U920 ( .B(A[172]), .A(S), .Z(O[172]) );
  ANDN U921 ( .B(A[171]), .A(S), .Z(O[171]) );
  ANDN U922 ( .B(A[170]), .A(S), .Z(O[170]) );
  ANDN U923 ( .B(A[16]), .A(S), .Z(O[16]) );
  ANDN U924 ( .B(A[169]), .A(S), .Z(O[169]) );
  ANDN U925 ( .B(A[168]), .A(S), .Z(O[168]) );
  ANDN U926 ( .B(A[167]), .A(S), .Z(O[167]) );
  ANDN U927 ( .B(A[166]), .A(S), .Z(O[166]) );
  ANDN U928 ( .B(A[165]), .A(S), .Z(O[165]) );
  ANDN U929 ( .B(A[164]), .A(S), .Z(O[164]) );
  ANDN U930 ( .B(A[163]), .A(S), .Z(O[163]) );
  ANDN U931 ( .B(A[162]), .A(S), .Z(O[162]) );
  ANDN U932 ( .B(A[161]), .A(S), .Z(O[161]) );
  ANDN U933 ( .B(A[160]), .A(S), .Z(O[160]) );
  ANDN U934 ( .B(A[15]), .A(S), .Z(O[15]) );
  ANDN U935 ( .B(A[159]), .A(S), .Z(O[159]) );
  ANDN U936 ( .B(A[158]), .A(S), .Z(O[158]) );
  ANDN U937 ( .B(A[157]), .A(S), .Z(O[157]) );
  ANDN U938 ( .B(A[156]), .A(S), .Z(O[156]) );
  ANDN U939 ( .B(A[155]), .A(S), .Z(O[155]) );
  ANDN U940 ( .B(A[154]), .A(S), .Z(O[154]) );
  ANDN U941 ( .B(A[153]), .A(S), .Z(O[153]) );
  ANDN U942 ( .B(A[152]), .A(S), .Z(O[152]) );
  ANDN U943 ( .B(A[151]), .A(S), .Z(O[151]) );
  ANDN U944 ( .B(A[150]), .A(S), .Z(O[150]) );
  ANDN U945 ( .B(A[14]), .A(S), .Z(O[14]) );
  ANDN U946 ( .B(A[149]), .A(S), .Z(O[149]) );
  ANDN U947 ( .B(A[148]), .A(S), .Z(O[148]) );
  ANDN U948 ( .B(A[147]), .A(S), .Z(O[147]) );
  ANDN U949 ( .B(A[146]), .A(S), .Z(O[146]) );
  ANDN U950 ( .B(A[145]), .A(S), .Z(O[145]) );
  ANDN U951 ( .B(A[144]), .A(S), .Z(O[144]) );
  ANDN U952 ( .B(A[143]), .A(S), .Z(O[143]) );
  ANDN U953 ( .B(A[142]), .A(S), .Z(O[142]) );
  ANDN U954 ( .B(A[141]), .A(S), .Z(O[141]) );
  ANDN U955 ( .B(A[140]), .A(S), .Z(O[140]) );
  ANDN U956 ( .B(A[13]), .A(S), .Z(O[13]) );
  ANDN U957 ( .B(A[139]), .A(S), .Z(O[139]) );
  ANDN U958 ( .B(A[138]), .A(S), .Z(O[138]) );
  ANDN U959 ( .B(A[137]), .A(S), .Z(O[137]) );
  ANDN U960 ( .B(A[136]), .A(S), .Z(O[136]) );
  ANDN U961 ( .B(A[135]), .A(S), .Z(O[135]) );
  ANDN U962 ( .B(A[134]), .A(S), .Z(O[134]) );
  ANDN U963 ( .B(A[133]), .A(S), .Z(O[133]) );
  ANDN U964 ( .B(A[132]), .A(S), .Z(O[132]) );
  ANDN U965 ( .B(A[131]), .A(S), .Z(O[131]) );
  ANDN U966 ( .B(A[130]), .A(S), .Z(O[130]) );
  ANDN U967 ( .B(A[12]), .A(S), .Z(O[12]) );
  ANDN U968 ( .B(A[129]), .A(S), .Z(O[129]) );
  ANDN U969 ( .B(A[128]), .A(S), .Z(O[128]) );
  ANDN U970 ( .B(A[127]), .A(S), .Z(O[127]) );
  ANDN U971 ( .B(A[126]), .A(S), .Z(O[126]) );
  ANDN U972 ( .B(A[125]), .A(S), .Z(O[125]) );
  ANDN U973 ( .B(A[124]), .A(S), .Z(O[124]) );
  ANDN U974 ( .B(A[123]), .A(S), .Z(O[123]) );
  ANDN U975 ( .B(A[122]), .A(S), .Z(O[122]) );
  ANDN U976 ( .B(A[121]), .A(S), .Z(O[121]) );
  ANDN U977 ( .B(A[120]), .A(S), .Z(O[120]) );
  ANDN U978 ( .B(A[11]), .A(S), .Z(O[11]) );
  ANDN U979 ( .B(A[119]), .A(S), .Z(O[119]) );
  ANDN U980 ( .B(A[118]), .A(S), .Z(O[118]) );
  ANDN U981 ( .B(A[117]), .A(S), .Z(O[117]) );
  ANDN U982 ( .B(A[116]), .A(S), .Z(O[116]) );
  ANDN U983 ( .B(A[115]), .A(S), .Z(O[115]) );
  ANDN U984 ( .B(A[114]), .A(S), .Z(O[114]) );
  ANDN U985 ( .B(A[113]), .A(S), .Z(O[113]) );
  ANDN U986 ( .B(A[112]), .A(S), .Z(O[112]) );
  ANDN U987 ( .B(A[111]), .A(S), .Z(O[111]) );
  ANDN U988 ( .B(A[110]), .A(S), .Z(O[110]) );
  ANDN U989 ( .B(A[10]), .A(S), .Z(O[10]) );
  ANDN U990 ( .B(A[109]), .A(S), .Z(O[109]) );
  ANDN U991 ( .B(A[108]), .A(S), .Z(O[108]) );
  ANDN U992 ( .B(A[107]), .A(S), .Z(O[107]) );
  ANDN U993 ( .B(A[106]), .A(S), .Z(O[106]) );
  ANDN U994 ( .B(A[105]), .A(S), .Z(O[105]) );
  ANDN U995 ( .B(A[104]), .A(S), .Z(O[104]) );
  ANDN U996 ( .B(A[103]), .A(S), .Z(O[103]) );
  ANDN U997 ( .B(A[102]), .A(S), .Z(O[102]) );
  ANDN U998 ( .B(A[1023]), .A(S), .Z(O[1023]) );
  ANDN U999 ( .B(A[1022]), .A(S), .Z(O[1022]) );
  ANDN U1000 ( .B(A[1021]), .A(S), .Z(O[1021]) );
  ANDN U1001 ( .B(A[1020]), .A(S), .Z(O[1020]) );
  ANDN U1002 ( .B(A[101]), .A(S), .Z(O[101]) );
  ANDN U1003 ( .B(A[1019]), .A(S), .Z(O[1019]) );
  ANDN U1004 ( .B(A[1018]), .A(S), .Z(O[1018]) );
  ANDN U1005 ( .B(A[1017]), .A(S), .Z(O[1017]) );
  ANDN U1006 ( .B(A[1016]), .A(S), .Z(O[1016]) );
  ANDN U1007 ( .B(A[1015]), .A(S), .Z(O[1015]) );
  ANDN U1008 ( .B(A[1014]), .A(S), .Z(O[1014]) );
  ANDN U1009 ( .B(A[1013]), .A(S), .Z(O[1013]) );
  ANDN U1010 ( .B(A[1012]), .A(S), .Z(O[1012]) );
  ANDN U1011 ( .B(A[1011]), .A(S), .Z(O[1011]) );
  ANDN U1012 ( .B(A[1010]), .A(S), .Z(O[1010]) );
  ANDN U1013 ( .B(A[100]), .A(S), .Z(O[100]) );
  ANDN U1014 ( .B(A[1009]), .A(S), .Z(O[1009]) );
  ANDN U1015 ( .B(A[1008]), .A(S), .Z(O[1008]) );
  ANDN U1016 ( .B(A[1007]), .A(S), .Z(O[1007]) );
  ANDN U1017 ( .B(A[1006]), .A(S), .Z(O[1006]) );
  ANDN U1018 ( .B(A[1005]), .A(S), .Z(O[1005]) );
  ANDN U1019 ( .B(A[1004]), .A(S), .Z(O[1004]) );
  ANDN U1020 ( .B(A[1003]), .A(S), .Z(O[1003]) );
  ANDN U1021 ( .B(A[1002]), .A(S), .Z(O[1002]) );
  ANDN U1022 ( .B(A[1001]), .A(S), .Z(O[1001]) );
  ANDN U1023 ( .B(A[1000]), .A(S), .Z(O[1000]) );
  ANDN U1024 ( .B(A[0]), .A(S), .Z(O[0]) );
endmodule


module FA_6437 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_15679 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(CI), .B(A), .Z(S) );
endmodule


module FA_15680 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  ANDN U1 ( .B(CI), .A(S), .Z(CO) );
  XOR U2 ( .A(A), .B(CI), .Z(S) );
endmodule


module FA_15681 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15682 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15683 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15684 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15685 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15686 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15687 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15688 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15689 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15690 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15691 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15692 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15693 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15694 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15695 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15696 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15697 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15698 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15699 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15700 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15701 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15702 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15703 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15704 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15705 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15706 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15707 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15708 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15709 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15710 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15711 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15712 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15713 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15714 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15715 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15716 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15717 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15718 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15719 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15720 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15721 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15722 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15723 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15724 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15725 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15726 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15727 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15728 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15729 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15730 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15731 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15732 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15733 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15734 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15735 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15736 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15737 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15738 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15739 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15740 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15741 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15742 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15743 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15744 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15745 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15746 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15747 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15748 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15749 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15750 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15751 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15752 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15753 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15754 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15755 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15756 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15757 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15758 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15759 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15760 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15761 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15762 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15763 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15764 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15765 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15766 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15767 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15768 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15769 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15770 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15771 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15772 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15773 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15774 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15775 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15776 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15777 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15778 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15779 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15780 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15781 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15782 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15783 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15784 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15785 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15786 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15787 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15788 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15789 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15790 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15791 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15792 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15793 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15794 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15795 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15796 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15797 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15798 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15799 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15800 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15801 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15802 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15803 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15804 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15805 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15806 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15807 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15808 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15809 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15810 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15811 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15812 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15813 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15814 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15815 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15816 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15817 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15818 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15819 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15820 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15821 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15822 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15823 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15824 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15825 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15826 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15827 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15828 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15829 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15830 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15831 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15832 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15833 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15834 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15835 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15836 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15837 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15838 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15839 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15840 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15841 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15842 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15843 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15844 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15845 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15846 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15847 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15848 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15849 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15850 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15851 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15852 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15853 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15854 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15855 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15856 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15857 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15858 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15859 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15860 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15861 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15862 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15863 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15864 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15865 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15866 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15867 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15868 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15869 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15870 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15871 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15872 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15873 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15874 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15875 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15876 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15877 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15878 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15879 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15880 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15881 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15882 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15883 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15884 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15885 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15886 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15887 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15888 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15889 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15890 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15891 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15892 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15893 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15894 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15895 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15896 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15897 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15898 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15899 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15900 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15901 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15902 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15903 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15904 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15905 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15906 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15907 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15908 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15909 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15910 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15911 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15912 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15913 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15914 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15915 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15916 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15917 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15918 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15919 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15920 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15921 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15922 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15923 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15924 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15925 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15926 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15927 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15928 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15929 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15930 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15931 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15932 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15933 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15934 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15935 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15936 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15937 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15938 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15939 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15940 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15941 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15942 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15943 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15944 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15945 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15946 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15947 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15948 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15949 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15950 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15951 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15952 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15953 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15954 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15955 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15956 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15957 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15958 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15959 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15960 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15961 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15962 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15963 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15964 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15965 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15966 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15967 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15968 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15969 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15970 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15971 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15972 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15973 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15974 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15975 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15976 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15977 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15978 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15979 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15980 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15981 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15982 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15983 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15984 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15985 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15986 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15987 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15988 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15989 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15990 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15991 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15992 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15993 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15994 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15995 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15996 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15997 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15998 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15999 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16000 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16001 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16002 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16003 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16004 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16005 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16006 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16007 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16008 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16009 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16010 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16011 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16012 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16013 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16014 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16015 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16016 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16017 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16018 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16019 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16020 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16021 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16022 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16023 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16024 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16025 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16026 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16027 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16028 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16029 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16030 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16031 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16032 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16033 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16034 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16035 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16036 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16037 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16038 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16039 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16040 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16041 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16042 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16043 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16044 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16045 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16046 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16047 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16048 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16049 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16050 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16051 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16052 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16053 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16054 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16055 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16056 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16057 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16058 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16059 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16060 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16061 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16062 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16063 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16064 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16065 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16066 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16067 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16068 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16069 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16070 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16071 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16072 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16073 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16074 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16075 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16076 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16077 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16078 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16079 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16080 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16081 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16082 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16083 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16084 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16085 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16086 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16087 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16088 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16089 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16090 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16091 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16092 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16093 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16094 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16095 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16096 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16097 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16098 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16099 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16100 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16101 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16102 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16103 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16104 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16105 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16106 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16107 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16108 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16109 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16110 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16111 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16112 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16113 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16114 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16115 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16116 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16117 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16118 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16119 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16120 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16121 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16122 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16123 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16124 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16125 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16126 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16127 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16128 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16129 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16130 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16131 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16132 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16133 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16134 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16135 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16136 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16137 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16138 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16139 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16140 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16141 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16142 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16143 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16144 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16145 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16146 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16147 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16148 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16149 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16150 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16151 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16152 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16153 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16154 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16155 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16156 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16157 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16158 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16159 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16160 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16161 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16162 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16163 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16164 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16165 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16166 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16167 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16168 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16169 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16170 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16171 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16172 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16173 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16174 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16175 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16176 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16177 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16178 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16179 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16180 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16181 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16182 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16183 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16184 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16185 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16186 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16187 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16188 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16189 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16190 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16191 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16192 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16193 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16194 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16195 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16196 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16197 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16198 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16199 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16200 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16201 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16202 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16203 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16204 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16205 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16206 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16207 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16208 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16209 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16210 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16211 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16212 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16213 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16214 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16215 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16216 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16217 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16218 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16219 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16220 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16221 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16222 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16223 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16224 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16225 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16226 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16227 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16228 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16229 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16230 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16231 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16232 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16233 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16234 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16235 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16236 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16237 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16238 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16239 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16240 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16241 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16242 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16243 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16244 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16245 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16246 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16247 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16248 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16249 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16250 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16251 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16252 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16253 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16254 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16255 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16256 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16257 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16258 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16259 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16260 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16261 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16262 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16263 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16264 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16265 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16266 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16267 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16268 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16269 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16270 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16271 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16272 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16273 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16274 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16275 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16276 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16277 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16278 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16279 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16280 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16281 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16282 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16283 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16284 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16285 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16286 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16287 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16288 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16289 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16290 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16291 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16292 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16293 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16294 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16295 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16296 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16297 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16298 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16299 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16300 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16301 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16302 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16303 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16304 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16305 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16306 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16307 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16308 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16309 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16310 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16311 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16312 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16313 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16314 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16315 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16316 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16317 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16318 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16319 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16320 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16321 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16322 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16323 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16324 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16325 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16326 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16327 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16328 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16329 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16330 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16331 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16332 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16333 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16334 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16335 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16336 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16337 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16338 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16339 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16340 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16341 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16342 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16343 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16344 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16345 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16346 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16347 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16348 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16349 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16350 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16351 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16352 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16353 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16354 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16355 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16356 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16357 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16358 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16359 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16360 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16361 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16362 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16363 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16364 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16365 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16366 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16367 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16368 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16369 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16370 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16371 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16372 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16373 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16374 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16375 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16376 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16377 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16378 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16379 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16380 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16381 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16382 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16383 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16384 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16385 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16386 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16387 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16388 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16389 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16390 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16391 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16392 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16393 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16394 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16395 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16396 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16397 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16398 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16399 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16400 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16401 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16402 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16403 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16404 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16405 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16406 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16407 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16408 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16409 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16410 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16411 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16412 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16413 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16414 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16415 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16416 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16417 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16418 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16419 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16420 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16421 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16422 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16423 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16424 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16425 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16426 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16427 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16428 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16429 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16430 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16431 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16432 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16433 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16434 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16435 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16436 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16437 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16438 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16439 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16440 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16441 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16442 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16443 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16444 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16445 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16446 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16447 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16448 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16449 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16450 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16451 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16452 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16453 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16454 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16455 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16456 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16457 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16458 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16459 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16460 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16461 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16462 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16463 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16464 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16465 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16466 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16467 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16468 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16469 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16470 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16471 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16472 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16473 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16474 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16475 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16476 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16477 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16478 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16479 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16480 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16481 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16482 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16483 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16484 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16485 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16486 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16487 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16488 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16489 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16490 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16491 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16492 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16493 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16494 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16495 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16496 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16497 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16498 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16499 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16500 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16501 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16502 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16503 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16504 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16505 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16506 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16507 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16508 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16509 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16510 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16511 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16512 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16513 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16514 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16515 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16516 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16517 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16518 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16519 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16520 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16521 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16522 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16523 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16524 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16525 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16526 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16527 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16528 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16529 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16530 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16531 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16532 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16533 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16534 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16535 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16536 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16537 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16538 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16539 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16540 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16541 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16542 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16543 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16544 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16545 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16546 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16547 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16548 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16549 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16550 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16551 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16552 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16553 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16554 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16555 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16556 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16557 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16558 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16559 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16560 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16561 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16562 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16563 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16564 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16565 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16566 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16567 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16568 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16569 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16570 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16571 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16572 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16573 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16574 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16575 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16576 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16577 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16578 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16579 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16580 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16581 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16582 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16583 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16584 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16585 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16586 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16587 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16588 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16589 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16590 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16591 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16592 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16593 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16594 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16595 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16596 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16597 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16598 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16599 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16600 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16601 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16602 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16603 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16604 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16605 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16606 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16607 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16608 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16609 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16610 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16611 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16612 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16613 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16614 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16615 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16616 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16617 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16618 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16619 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16620 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16621 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16622 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16623 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16624 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16625 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16626 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16627 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16628 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16629 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16630 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16631 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16632 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16633 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16634 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16635 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16636 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16637 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16638 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16639 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16640 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16641 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16642 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16643 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16644 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16645 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16646 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16647 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16648 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16649 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16650 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16651 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16652 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16653 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16654 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16655 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16656 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16657 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16658 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16659 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16660 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16661 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16662 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16663 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16664 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16665 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16666 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16667 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16668 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16669 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16670 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16671 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16672 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16673 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16674 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16675 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16676 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16677 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16678 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16679 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16680 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16681 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16682 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16683 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16684 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16685 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16686 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16687 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16688 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16689 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16690 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16691 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16692 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16693 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16694 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16695 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16696 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16697 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16698 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16699 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16700 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16701 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16702 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16703 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module ADD_N1026 ( A, B, CI, S, CO );
  input [1025:0] A;
  input [1025:0] B;
  output [1025:0] S;
  input CI;
  output CO;

  wire   [1025:1] C;

  FA_6437 \FA_INST_0[0].FA_INST_1[0].FA_  ( .A(1'b0), .B(B[0]), .CI(1'b0), .S(
        S[0]) );
  FA_16703 \FA_INST_0[0].FA_INST_1[1].FA_  ( .A(A[1]), .B(B[1]), .CI(1'b0), 
        .S(S[1]), .CO(C[2]) );
  FA_16702 \FA_INST_0[0].FA_INST_1[2].FA_  ( .A(A[2]), .B(B[2]), .CI(C[2]), 
        .S(S[2]), .CO(C[3]) );
  FA_16701 \FA_INST_0[0].FA_INST_1[3].FA_  ( .A(A[3]), .B(B[3]), .CI(C[3]), 
        .S(S[3]), .CO(C[4]) );
  FA_16700 \FA_INST_0[0].FA_INST_1[4].FA_  ( .A(A[4]), .B(B[4]), .CI(C[4]), 
        .S(S[4]), .CO(C[5]) );
  FA_16699 \FA_INST_0[0].FA_INST_1[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), 
        .S(S[5]), .CO(C[6]) );
  FA_16698 \FA_INST_0[0].FA_INST_1[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), 
        .S(S[6]), .CO(C[7]) );
  FA_16697 \FA_INST_0[0].FA_INST_1[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), 
        .S(S[7]), .CO(C[8]) );
  FA_16696 \FA_INST_0[0].FA_INST_1[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), 
        .S(S[8]), .CO(C[9]) );
  FA_16695 \FA_INST_0[0].FA_INST_1[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), 
        .S(S[9]), .CO(C[10]) );
  FA_16694 \FA_INST_0[0].FA_INST_1[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), 
        .S(S[10]), .CO(C[11]) );
  FA_16693 \FA_INST_0[0].FA_INST_1[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), 
        .S(S[11]), .CO(C[12]) );
  FA_16692 \FA_INST_0[0].FA_INST_1[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), 
        .S(S[12]), .CO(C[13]) );
  FA_16691 \FA_INST_0[0].FA_INST_1[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), 
        .S(S[13]), .CO(C[14]) );
  FA_16690 \FA_INST_0[0].FA_INST_1[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), 
        .S(S[14]), .CO(C[15]) );
  FA_16689 \FA_INST_0[0].FA_INST_1[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), 
        .S(S[15]), .CO(C[16]) );
  FA_16688 \FA_INST_0[0].FA_INST_1[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), 
        .S(S[16]), .CO(C[17]) );
  FA_16687 \FA_INST_0[0].FA_INST_1[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), 
        .S(S[17]), .CO(C[18]) );
  FA_16686 \FA_INST_0[0].FA_INST_1[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), 
        .S(S[18]), .CO(C[19]) );
  FA_16685 \FA_INST_0[0].FA_INST_1[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), 
        .S(S[19]), .CO(C[20]) );
  FA_16684 \FA_INST_0[0].FA_INST_1[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), 
        .S(S[20]), .CO(C[21]) );
  FA_16683 \FA_INST_0[0].FA_INST_1[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), 
        .S(S[21]), .CO(C[22]) );
  FA_16682 \FA_INST_0[0].FA_INST_1[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), 
        .S(S[22]), .CO(C[23]) );
  FA_16681 \FA_INST_0[0].FA_INST_1[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), 
        .S(S[23]), .CO(C[24]) );
  FA_16680 \FA_INST_0[0].FA_INST_1[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), 
        .S(S[24]), .CO(C[25]) );
  FA_16679 \FA_INST_0[0].FA_INST_1[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), 
        .S(S[25]), .CO(C[26]) );
  FA_16678 \FA_INST_0[0].FA_INST_1[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), 
        .S(S[26]), .CO(C[27]) );
  FA_16677 \FA_INST_0[0].FA_INST_1[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), 
        .S(S[27]), .CO(C[28]) );
  FA_16676 \FA_INST_0[0].FA_INST_1[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), 
        .S(S[28]), .CO(C[29]) );
  FA_16675 \FA_INST_0[0].FA_INST_1[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), 
        .S(S[29]), .CO(C[30]) );
  FA_16674 \FA_INST_0[0].FA_INST_1[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), 
        .S(S[30]), .CO(C[31]) );
  FA_16673 \FA_INST_0[0].FA_INST_1[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), 
        .S(S[31]), .CO(C[32]) );
  FA_16672 \FA_INST_0[0].FA_INST_1[32].FA_  ( .A(A[32]), .B(B[32]), .CI(C[32]), 
        .S(S[32]), .CO(C[33]) );
  FA_16671 \FA_INST_0[0].FA_INST_1[33].FA_  ( .A(A[33]), .B(B[33]), .CI(C[33]), 
        .S(S[33]), .CO(C[34]) );
  FA_16670 \FA_INST_0[0].FA_INST_1[34].FA_  ( .A(A[34]), .B(B[34]), .CI(C[34]), 
        .S(S[34]), .CO(C[35]) );
  FA_16669 \FA_INST_0[0].FA_INST_1[35].FA_  ( .A(A[35]), .B(B[35]), .CI(C[35]), 
        .S(S[35]), .CO(C[36]) );
  FA_16668 \FA_INST_0[0].FA_INST_1[36].FA_  ( .A(A[36]), .B(B[36]), .CI(C[36]), 
        .S(S[36]), .CO(C[37]) );
  FA_16667 \FA_INST_0[0].FA_INST_1[37].FA_  ( .A(A[37]), .B(B[37]), .CI(C[37]), 
        .S(S[37]), .CO(C[38]) );
  FA_16666 \FA_INST_0[0].FA_INST_1[38].FA_  ( .A(A[38]), .B(B[38]), .CI(C[38]), 
        .S(S[38]), .CO(C[39]) );
  FA_16665 \FA_INST_0[0].FA_INST_1[39].FA_  ( .A(A[39]), .B(B[39]), .CI(C[39]), 
        .S(S[39]), .CO(C[40]) );
  FA_16664 \FA_INST_0[0].FA_INST_1[40].FA_  ( .A(A[40]), .B(B[40]), .CI(C[40]), 
        .S(S[40]), .CO(C[41]) );
  FA_16663 \FA_INST_0[0].FA_INST_1[41].FA_  ( .A(A[41]), .B(B[41]), .CI(C[41]), 
        .S(S[41]), .CO(C[42]) );
  FA_16662 \FA_INST_0[0].FA_INST_1[42].FA_  ( .A(A[42]), .B(B[42]), .CI(C[42]), 
        .S(S[42]), .CO(C[43]) );
  FA_16661 \FA_INST_0[0].FA_INST_1[43].FA_  ( .A(A[43]), .B(B[43]), .CI(C[43]), 
        .S(S[43]), .CO(C[44]) );
  FA_16660 \FA_INST_0[0].FA_INST_1[44].FA_  ( .A(A[44]), .B(B[44]), .CI(C[44]), 
        .S(S[44]), .CO(C[45]) );
  FA_16659 \FA_INST_0[0].FA_INST_1[45].FA_  ( .A(A[45]), .B(B[45]), .CI(C[45]), 
        .S(S[45]), .CO(C[46]) );
  FA_16658 \FA_INST_0[0].FA_INST_1[46].FA_  ( .A(A[46]), .B(B[46]), .CI(C[46]), 
        .S(S[46]), .CO(C[47]) );
  FA_16657 \FA_INST_0[0].FA_INST_1[47].FA_  ( .A(A[47]), .B(B[47]), .CI(C[47]), 
        .S(S[47]), .CO(C[48]) );
  FA_16656 \FA_INST_0[0].FA_INST_1[48].FA_  ( .A(A[48]), .B(B[48]), .CI(C[48]), 
        .S(S[48]), .CO(C[49]) );
  FA_16655 \FA_INST_0[0].FA_INST_1[49].FA_  ( .A(A[49]), .B(B[49]), .CI(C[49]), 
        .S(S[49]), .CO(C[50]) );
  FA_16654 \FA_INST_0[0].FA_INST_1[50].FA_  ( .A(A[50]), .B(B[50]), .CI(C[50]), 
        .S(S[50]), .CO(C[51]) );
  FA_16653 \FA_INST_0[0].FA_INST_1[51].FA_  ( .A(A[51]), .B(B[51]), .CI(C[51]), 
        .S(S[51]), .CO(C[52]) );
  FA_16652 \FA_INST_0[0].FA_INST_1[52].FA_  ( .A(A[52]), .B(B[52]), .CI(C[52]), 
        .S(S[52]), .CO(C[53]) );
  FA_16651 \FA_INST_0[0].FA_INST_1[53].FA_  ( .A(A[53]), .B(B[53]), .CI(C[53]), 
        .S(S[53]), .CO(C[54]) );
  FA_16650 \FA_INST_0[0].FA_INST_1[54].FA_  ( .A(A[54]), .B(B[54]), .CI(C[54]), 
        .S(S[54]), .CO(C[55]) );
  FA_16649 \FA_INST_0[0].FA_INST_1[55].FA_  ( .A(A[55]), .B(B[55]), .CI(C[55]), 
        .S(S[55]), .CO(C[56]) );
  FA_16648 \FA_INST_0[0].FA_INST_1[56].FA_  ( .A(A[56]), .B(B[56]), .CI(C[56]), 
        .S(S[56]), .CO(C[57]) );
  FA_16647 \FA_INST_0[0].FA_INST_1[57].FA_  ( .A(A[57]), .B(B[57]), .CI(C[57]), 
        .S(S[57]), .CO(C[58]) );
  FA_16646 \FA_INST_0[0].FA_INST_1[58].FA_  ( .A(A[58]), .B(B[58]), .CI(C[58]), 
        .S(S[58]), .CO(C[59]) );
  FA_16645 \FA_INST_0[0].FA_INST_1[59].FA_  ( .A(A[59]), .B(B[59]), .CI(C[59]), 
        .S(S[59]), .CO(C[60]) );
  FA_16644 \FA_INST_0[0].FA_INST_1[60].FA_  ( .A(A[60]), .B(B[60]), .CI(C[60]), 
        .S(S[60]), .CO(C[61]) );
  FA_16643 \FA_INST_0[0].FA_INST_1[61].FA_  ( .A(A[61]), .B(B[61]), .CI(C[61]), 
        .S(S[61]), .CO(C[62]) );
  FA_16642 \FA_INST_0[0].FA_INST_1[62].FA_  ( .A(A[62]), .B(B[62]), .CI(C[62]), 
        .S(S[62]), .CO(C[63]) );
  FA_16641 \FA_INST_0[0].FA_INST_1[63].FA_  ( .A(A[63]), .B(B[63]), .CI(C[63]), 
        .S(S[63]), .CO(C[64]) );
  FA_16640 \FA_INST_0[0].FA_INST_1[64].FA_  ( .A(A[64]), .B(B[64]), .CI(C[64]), 
        .S(S[64]), .CO(C[65]) );
  FA_16639 \FA_INST_0[0].FA_INST_1[65].FA_  ( .A(A[65]), .B(B[65]), .CI(C[65]), 
        .S(S[65]), .CO(C[66]) );
  FA_16638 \FA_INST_0[0].FA_INST_1[66].FA_  ( .A(A[66]), .B(B[66]), .CI(C[66]), 
        .S(S[66]), .CO(C[67]) );
  FA_16637 \FA_INST_0[0].FA_INST_1[67].FA_  ( .A(A[67]), .B(B[67]), .CI(C[67]), 
        .S(S[67]), .CO(C[68]) );
  FA_16636 \FA_INST_0[0].FA_INST_1[68].FA_  ( .A(A[68]), .B(B[68]), .CI(C[68]), 
        .S(S[68]), .CO(C[69]) );
  FA_16635 \FA_INST_0[0].FA_INST_1[69].FA_  ( .A(A[69]), .B(B[69]), .CI(C[69]), 
        .S(S[69]), .CO(C[70]) );
  FA_16634 \FA_INST_0[0].FA_INST_1[70].FA_  ( .A(A[70]), .B(B[70]), .CI(C[70]), 
        .S(S[70]), .CO(C[71]) );
  FA_16633 \FA_INST_0[0].FA_INST_1[71].FA_  ( .A(A[71]), .B(B[71]), .CI(C[71]), 
        .S(S[71]), .CO(C[72]) );
  FA_16632 \FA_INST_0[0].FA_INST_1[72].FA_  ( .A(A[72]), .B(B[72]), .CI(C[72]), 
        .S(S[72]), .CO(C[73]) );
  FA_16631 \FA_INST_0[0].FA_INST_1[73].FA_  ( .A(A[73]), .B(B[73]), .CI(C[73]), 
        .S(S[73]), .CO(C[74]) );
  FA_16630 \FA_INST_0[0].FA_INST_1[74].FA_  ( .A(A[74]), .B(B[74]), .CI(C[74]), 
        .S(S[74]), .CO(C[75]) );
  FA_16629 \FA_INST_0[0].FA_INST_1[75].FA_  ( .A(A[75]), .B(B[75]), .CI(C[75]), 
        .S(S[75]), .CO(C[76]) );
  FA_16628 \FA_INST_0[0].FA_INST_1[76].FA_  ( .A(A[76]), .B(B[76]), .CI(C[76]), 
        .S(S[76]), .CO(C[77]) );
  FA_16627 \FA_INST_0[0].FA_INST_1[77].FA_  ( .A(A[77]), .B(B[77]), .CI(C[77]), 
        .S(S[77]), .CO(C[78]) );
  FA_16626 \FA_INST_0[0].FA_INST_1[78].FA_  ( .A(A[78]), .B(B[78]), .CI(C[78]), 
        .S(S[78]), .CO(C[79]) );
  FA_16625 \FA_INST_0[0].FA_INST_1[79].FA_  ( .A(A[79]), .B(B[79]), .CI(C[79]), 
        .S(S[79]), .CO(C[80]) );
  FA_16624 \FA_INST_0[0].FA_INST_1[80].FA_  ( .A(A[80]), .B(B[80]), .CI(C[80]), 
        .S(S[80]), .CO(C[81]) );
  FA_16623 \FA_INST_0[0].FA_INST_1[81].FA_  ( .A(A[81]), .B(B[81]), .CI(C[81]), 
        .S(S[81]), .CO(C[82]) );
  FA_16622 \FA_INST_0[0].FA_INST_1[82].FA_  ( .A(A[82]), .B(B[82]), .CI(C[82]), 
        .S(S[82]), .CO(C[83]) );
  FA_16621 \FA_INST_0[0].FA_INST_1[83].FA_  ( .A(A[83]), .B(B[83]), .CI(C[83]), 
        .S(S[83]), .CO(C[84]) );
  FA_16620 \FA_INST_0[0].FA_INST_1[84].FA_  ( .A(A[84]), .B(B[84]), .CI(C[84]), 
        .S(S[84]), .CO(C[85]) );
  FA_16619 \FA_INST_0[0].FA_INST_1[85].FA_  ( .A(A[85]), .B(B[85]), .CI(C[85]), 
        .S(S[85]), .CO(C[86]) );
  FA_16618 \FA_INST_0[0].FA_INST_1[86].FA_  ( .A(A[86]), .B(B[86]), .CI(C[86]), 
        .S(S[86]), .CO(C[87]) );
  FA_16617 \FA_INST_0[0].FA_INST_1[87].FA_  ( .A(A[87]), .B(B[87]), .CI(C[87]), 
        .S(S[87]), .CO(C[88]) );
  FA_16616 \FA_INST_0[0].FA_INST_1[88].FA_  ( .A(A[88]), .B(B[88]), .CI(C[88]), 
        .S(S[88]), .CO(C[89]) );
  FA_16615 \FA_INST_0[0].FA_INST_1[89].FA_  ( .A(A[89]), .B(B[89]), .CI(C[89]), 
        .S(S[89]), .CO(C[90]) );
  FA_16614 \FA_INST_0[0].FA_INST_1[90].FA_  ( .A(A[90]), .B(B[90]), .CI(C[90]), 
        .S(S[90]), .CO(C[91]) );
  FA_16613 \FA_INST_0[0].FA_INST_1[91].FA_  ( .A(A[91]), .B(B[91]), .CI(C[91]), 
        .S(S[91]), .CO(C[92]) );
  FA_16612 \FA_INST_0[0].FA_INST_1[92].FA_  ( .A(A[92]), .B(B[92]), .CI(C[92]), 
        .S(S[92]), .CO(C[93]) );
  FA_16611 \FA_INST_0[0].FA_INST_1[93].FA_  ( .A(A[93]), .B(B[93]), .CI(C[93]), 
        .S(S[93]), .CO(C[94]) );
  FA_16610 \FA_INST_0[0].FA_INST_1[94].FA_  ( .A(A[94]), .B(B[94]), .CI(C[94]), 
        .S(S[94]), .CO(C[95]) );
  FA_16609 \FA_INST_0[0].FA_INST_1[95].FA_  ( .A(A[95]), .B(B[95]), .CI(C[95]), 
        .S(S[95]), .CO(C[96]) );
  FA_16608 \FA_INST_0[0].FA_INST_1[96].FA_  ( .A(A[96]), .B(B[96]), .CI(C[96]), 
        .S(S[96]), .CO(C[97]) );
  FA_16607 \FA_INST_0[0].FA_INST_1[97].FA_  ( .A(A[97]), .B(B[97]), .CI(C[97]), 
        .S(S[97]), .CO(C[98]) );
  FA_16606 \FA_INST_0[0].FA_INST_1[98].FA_  ( .A(A[98]), .B(B[98]), .CI(C[98]), 
        .S(S[98]), .CO(C[99]) );
  FA_16605 \FA_INST_0[0].FA_INST_1[99].FA_  ( .A(A[99]), .B(B[99]), .CI(C[99]), 
        .S(S[99]), .CO(C[100]) );
  FA_16604 \FA_INST_0[0].FA_INST_1[100].FA_  ( .A(A[100]), .B(B[100]), .CI(
        C[100]), .S(S[100]), .CO(C[101]) );
  FA_16603 \FA_INST_0[0].FA_INST_1[101].FA_  ( .A(A[101]), .B(B[101]), .CI(
        C[101]), .S(S[101]), .CO(C[102]) );
  FA_16602 \FA_INST_0[0].FA_INST_1[102].FA_  ( .A(A[102]), .B(B[102]), .CI(
        C[102]), .S(S[102]), .CO(C[103]) );
  FA_16601 \FA_INST_0[0].FA_INST_1[103].FA_  ( .A(A[103]), .B(B[103]), .CI(
        C[103]), .S(S[103]), .CO(C[104]) );
  FA_16600 \FA_INST_0[0].FA_INST_1[104].FA_  ( .A(A[104]), .B(B[104]), .CI(
        C[104]), .S(S[104]), .CO(C[105]) );
  FA_16599 \FA_INST_0[0].FA_INST_1[105].FA_  ( .A(A[105]), .B(B[105]), .CI(
        C[105]), .S(S[105]), .CO(C[106]) );
  FA_16598 \FA_INST_0[0].FA_INST_1[106].FA_  ( .A(A[106]), .B(B[106]), .CI(
        C[106]), .S(S[106]), .CO(C[107]) );
  FA_16597 \FA_INST_0[0].FA_INST_1[107].FA_  ( .A(A[107]), .B(B[107]), .CI(
        C[107]), .S(S[107]), .CO(C[108]) );
  FA_16596 \FA_INST_0[0].FA_INST_1[108].FA_  ( .A(A[108]), .B(B[108]), .CI(
        C[108]), .S(S[108]), .CO(C[109]) );
  FA_16595 \FA_INST_0[0].FA_INST_1[109].FA_  ( .A(A[109]), .B(B[109]), .CI(
        C[109]), .S(S[109]), .CO(C[110]) );
  FA_16594 \FA_INST_0[0].FA_INST_1[110].FA_  ( .A(A[110]), .B(B[110]), .CI(
        C[110]), .S(S[110]), .CO(C[111]) );
  FA_16593 \FA_INST_0[0].FA_INST_1[111].FA_  ( .A(A[111]), .B(B[111]), .CI(
        C[111]), .S(S[111]), .CO(C[112]) );
  FA_16592 \FA_INST_0[0].FA_INST_1[112].FA_  ( .A(A[112]), .B(B[112]), .CI(
        C[112]), .S(S[112]), .CO(C[113]) );
  FA_16591 \FA_INST_0[0].FA_INST_1[113].FA_  ( .A(A[113]), .B(B[113]), .CI(
        C[113]), .S(S[113]), .CO(C[114]) );
  FA_16590 \FA_INST_0[0].FA_INST_1[114].FA_  ( .A(A[114]), .B(B[114]), .CI(
        C[114]), .S(S[114]), .CO(C[115]) );
  FA_16589 \FA_INST_0[0].FA_INST_1[115].FA_  ( .A(A[115]), .B(B[115]), .CI(
        C[115]), .S(S[115]), .CO(C[116]) );
  FA_16588 \FA_INST_0[0].FA_INST_1[116].FA_  ( .A(A[116]), .B(B[116]), .CI(
        C[116]), .S(S[116]), .CO(C[117]) );
  FA_16587 \FA_INST_0[0].FA_INST_1[117].FA_  ( .A(A[117]), .B(B[117]), .CI(
        C[117]), .S(S[117]), .CO(C[118]) );
  FA_16586 \FA_INST_0[0].FA_INST_1[118].FA_  ( .A(A[118]), .B(B[118]), .CI(
        C[118]), .S(S[118]), .CO(C[119]) );
  FA_16585 \FA_INST_0[0].FA_INST_1[119].FA_  ( .A(A[119]), .B(B[119]), .CI(
        C[119]), .S(S[119]), .CO(C[120]) );
  FA_16584 \FA_INST_0[0].FA_INST_1[120].FA_  ( .A(A[120]), .B(B[120]), .CI(
        C[120]), .S(S[120]), .CO(C[121]) );
  FA_16583 \FA_INST_0[0].FA_INST_1[121].FA_  ( .A(A[121]), .B(B[121]), .CI(
        C[121]), .S(S[121]), .CO(C[122]) );
  FA_16582 \FA_INST_0[0].FA_INST_1[122].FA_  ( .A(A[122]), .B(B[122]), .CI(
        C[122]), .S(S[122]), .CO(C[123]) );
  FA_16581 \FA_INST_0[0].FA_INST_1[123].FA_  ( .A(A[123]), .B(B[123]), .CI(
        C[123]), .S(S[123]), .CO(C[124]) );
  FA_16580 \FA_INST_0[0].FA_INST_1[124].FA_  ( .A(A[124]), .B(B[124]), .CI(
        C[124]), .S(S[124]), .CO(C[125]) );
  FA_16579 \FA_INST_0[0].FA_INST_1[125].FA_  ( .A(A[125]), .B(B[125]), .CI(
        C[125]), .S(S[125]), .CO(C[126]) );
  FA_16578 \FA_INST_0[0].FA_INST_1[126].FA_  ( .A(A[126]), .B(B[126]), .CI(
        C[126]), .S(S[126]), .CO(C[127]) );
  FA_16577 \FA_INST_0[0].FA_INST_1[127].FA_  ( .A(A[127]), .B(B[127]), .CI(
        C[127]), .S(S[127]), .CO(C[128]) );
  FA_16576 \FA_INST_0[0].FA_INST_1[128].FA_  ( .A(A[128]), .B(B[128]), .CI(
        C[128]), .S(S[128]), .CO(C[129]) );
  FA_16575 \FA_INST_0[0].FA_INST_1[129].FA_  ( .A(A[129]), .B(B[129]), .CI(
        C[129]), .S(S[129]), .CO(C[130]) );
  FA_16574 \FA_INST_0[0].FA_INST_1[130].FA_  ( .A(A[130]), .B(B[130]), .CI(
        C[130]), .S(S[130]), .CO(C[131]) );
  FA_16573 \FA_INST_0[0].FA_INST_1[131].FA_  ( .A(A[131]), .B(B[131]), .CI(
        C[131]), .S(S[131]), .CO(C[132]) );
  FA_16572 \FA_INST_0[0].FA_INST_1[132].FA_  ( .A(A[132]), .B(B[132]), .CI(
        C[132]), .S(S[132]), .CO(C[133]) );
  FA_16571 \FA_INST_0[0].FA_INST_1[133].FA_  ( .A(A[133]), .B(B[133]), .CI(
        C[133]), .S(S[133]), .CO(C[134]) );
  FA_16570 \FA_INST_0[0].FA_INST_1[134].FA_  ( .A(A[134]), .B(B[134]), .CI(
        C[134]), .S(S[134]), .CO(C[135]) );
  FA_16569 \FA_INST_0[0].FA_INST_1[135].FA_  ( .A(A[135]), .B(B[135]), .CI(
        C[135]), .S(S[135]), .CO(C[136]) );
  FA_16568 \FA_INST_0[0].FA_INST_1[136].FA_  ( .A(A[136]), .B(B[136]), .CI(
        C[136]), .S(S[136]), .CO(C[137]) );
  FA_16567 \FA_INST_0[0].FA_INST_1[137].FA_  ( .A(A[137]), .B(B[137]), .CI(
        C[137]), .S(S[137]), .CO(C[138]) );
  FA_16566 \FA_INST_0[0].FA_INST_1[138].FA_  ( .A(A[138]), .B(B[138]), .CI(
        C[138]), .S(S[138]), .CO(C[139]) );
  FA_16565 \FA_INST_0[0].FA_INST_1[139].FA_  ( .A(A[139]), .B(B[139]), .CI(
        C[139]), .S(S[139]), .CO(C[140]) );
  FA_16564 \FA_INST_0[0].FA_INST_1[140].FA_  ( .A(A[140]), .B(B[140]), .CI(
        C[140]), .S(S[140]), .CO(C[141]) );
  FA_16563 \FA_INST_0[0].FA_INST_1[141].FA_  ( .A(A[141]), .B(B[141]), .CI(
        C[141]), .S(S[141]), .CO(C[142]) );
  FA_16562 \FA_INST_0[0].FA_INST_1[142].FA_  ( .A(A[142]), .B(B[142]), .CI(
        C[142]), .S(S[142]), .CO(C[143]) );
  FA_16561 \FA_INST_0[0].FA_INST_1[143].FA_  ( .A(A[143]), .B(B[143]), .CI(
        C[143]), .S(S[143]), .CO(C[144]) );
  FA_16560 \FA_INST_0[0].FA_INST_1[144].FA_  ( .A(A[144]), .B(B[144]), .CI(
        C[144]), .S(S[144]), .CO(C[145]) );
  FA_16559 \FA_INST_0[0].FA_INST_1[145].FA_  ( .A(A[145]), .B(B[145]), .CI(
        C[145]), .S(S[145]), .CO(C[146]) );
  FA_16558 \FA_INST_0[0].FA_INST_1[146].FA_  ( .A(A[146]), .B(B[146]), .CI(
        C[146]), .S(S[146]), .CO(C[147]) );
  FA_16557 \FA_INST_0[0].FA_INST_1[147].FA_  ( .A(A[147]), .B(B[147]), .CI(
        C[147]), .S(S[147]), .CO(C[148]) );
  FA_16556 \FA_INST_0[0].FA_INST_1[148].FA_  ( .A(A[148]), .B(B[148]), .CI(
        C[148]), .S(S[148]), .CO(C[149]) );
  FA_16555 \FA_INST_0[0].FA_INST_1[149].FA_  ( .A(A[149]), .B(B[149]), .CI(
        C[149]), .S(S[149]), .CO(C[150]) );
  FA_16554 \FA_INST_0[0].FA_INST_1[150].FA_  ( .A(A[150]), .B(B[150]), .CI(
        C[150]), .S(S[150]), .CO(C[151]) );
  FA_16553 \FA_INST_0[0].FA_INST_1[151].FA_  ( .A(A[151]), .B(B[151]), .CI(
        C[151]), .S(S[151]), .CO(C[152]) );
  FA_16552 \FA_INST_0[0].FA_INST_1[152].FA_  ( .A(A[152]), .B(B[152]), .CI(
        C[152]), .S(S[152]), .CO(C[153]) );
  FA_16551 \FA_INST_0[0].FA_INST_1[153].FA_  ( .A(A[153]), .B(B[153]), .CI(
        C[153]), .S(S[153]), .CO(C[154]) );
  FA_16550 \FA_INST_0[0].FA_INST_1[154].FA_  ( .A(A[154]), .B(B[154]), .CI(
        C[154]), .S(S[154]), .CO(C[155]) );
  FA_16549 \FA_INST_0[0].FA_INST_1[155].FA_  ( .A(A[155]), .B(B[155]), .CI(
        C[155]), .S(S[155]), .CO(C[156]) );
  FA_16548 \FA_INST_0[0].FA_INST_1[156].FA_  ( .A(A[156]), .B(B[156]), .CI(
        C[156]), .S(S[156]), .CO(C[157]) );
  FA_16547 \FA_INST_0[0].FA_INST_1[157].FA_  ( .A(A[157]), .B(B[157]), .CI(
        C[157]), .S(S[157]), .CO(C[158]) );
  FA_16546 \FA_INST_0[0].FA_INST_1[158].FA_  ( .A(A[158]), .B(B[158]), .CI(
        C[158]), .S(S[158]), .CO(C[159]) );
  FA_16545 \FA_INST_0[0].FA_INST_1[159].FA_  ( .A(A[159]), .B(B[159]), .CI(
        C[159]), .S(S[159]), .CO(C[160]) );
  FA_16544 \FA_INST_0[0].FA_INST_1[160].FA_  ( .A(A[160]), .B(B[160]), .CI(
        C[160]), .S(S[160]), .CO(C[161]) );
  FA_16543 \FA_INST_0[0].FA_INST_1[161].FA_  ( .A(A[161]), .B(B[161]), .CI(
        C[161]), .S(S[161]), .CO(C[162]) );
  FA_16542 \FA_INST_0[0].FA_INST_1[162].FA_  ( .A(A[162]), .B(B[162]), .CI(
        C[162]), .S(S[162]), .CO(C[163]) );
  FA_16541 \FA_INST_0[0].FA_INST_1[163].FA_  ( .A(A[163]), .B(B[163]), .CI(
        C[163]), .S(S[163]), .CO(C[164]) );
  FA_16540 \FA_INST_0[0].FA_INST_1[164].FA_  ( .A(A[164]), .B(B[164]), .CI(
        C[164]), .S(S[164]), .CO(C[165]) );
  FA_16539 \FA_INST_0[0].FA_INST_1[165].FA_  ( .A(A[165]), .B(B[165]), .CI(
        C[165]), .S(S[165]), .CO(C[166]) );
  FA_16538 \FA_INST_0[0].FA_INST_1[166].FA_  ( .A(A[166]), .B(B[166]), .CI(
        C[166]), .S(S[166]), .CO(C[167]) );
  FA_16537 \FA_INST_0[0].FA_INST_1[167].FA_  ( .A(A[167]), .B(B[167]), .CI(
        C[167]), .S(S[167]), .CO(C[168]) );
  FA_16536 \FA_INST_0[0].FA_INST_1[168].FA_  ( .A(A[168]), .B(B[168]), .CI(
        C[168]), .S(S[168]), .CO(C[169]) );
  FA_16535 \FA_INST_0[0].FA_INST_1[169].FA_  ( .A(A[169]), .B(B[169]), .CI(
        C[169]), .S(S[169]), .CO(C[170]) );
  FA_16534 \FA_INST_0[0].FA_INST_1[170].FA_  ( .A(A[170]), .B(B[170]), .CI(
        C[170]), .S(S[170]), .CO(C[171]) );
  FA_16533 \FA_INST_0[0].FA_INST_1[171].FA_  ( .A(A[171]), .B(B[171]), .CI(
        C[171]), .S(S[171]), .CO(C[172]) );
  FA_16532 \FA_INST_0[0].FA_INST_1[172].FA_  ( .A(A[172]), .B(B[172]), .CI(
        C[172]), .S(S[172]), .CO(C[173]) );
  FA_16531 \FA_INST_0[0].FA_INST_1[173].FA_  ( .A(A[173]), .B(B[173]), .CI(
        C[173]), .S(S[173]), .CO(C[174]) );
  FA_16530 \FA_INST_0[0].FA_INST_1[174].FA_  ( .A(A[174]), .B(B[174]), .CI(
        C[174]), .S(S[174]), .CO(C[175]) );
  FA_16529 \FA_INST_0[0].FA_INST_1[175].FA_  ( .A(A[175]), .B(B[175]), .CI(
        C[175]), .S(S[175]), .CO(C[176]) );
  FA_16528 \FA_INST_0[0].FA_INST_1[176].FA_  ( .A(A[176]), .B(B[176]), .CI(
        C[176]), .S(S[176]), .CO(C[177]) );
  FA_16527 \FA_INST_0[0].FA_INST_1[177].FA_  ( .A(A[177]), .B(B[177]), .CI(
        C[177]), .S(S[177]), .CO(C[178]) );
  FA_16526 \FA_INST_0[0].FA_INST_1[178].FA_  ( .A(A[178]), .B(B[178]), .CI(
        C[178]), .S(S[178]), .CO(C[179]) );
  FA_16525 \FA_INST_0[0].FA_INST_1[179].FA_  ( .A(A[179]), .B(B[179]), .CI(
        C[179]), .S(S[179]), .CO(C[180]) );
  FA_16524 \FA_INST_0[0].FA_INST_1[180].FA_  ( .A(A[180]), .B(B[180]), .CI(
        C[180]), .S(S[180]), .CO(C[181]) );
  FA_16523 \FA_INST_0[0].FA_INST_1[181].FA_  ( .A(A[181]), .B(B[181]), .CI(
        C[181]), .S(S[181]), .CO(C[182]) );
  FA_16522 \FA_INST_0[0].FA_INST_1[182].FA_  ( .A(A[182]), .B(B[182]), .CI(
        C[182]), .S(S[182]), .CO(C[183]) );
  FA_16521 \FA_INST_0[0].FA_INST_1[183].FA_  ( .A(A[183]), .B(B[183]), .CI(
        C[183]), .S(S[183]), .CO(C[184]) );
  FA_16520 \FA_INST_0[0].FA_INST_1[184].FA_  ( .A(A[184]), .B(B[184]), .CI(
        C[184]), .S(S[184]), .CO(C[185]) );
  FA_16519 \FA_INST_0[0].FA_INST_1[185].FA_  ( .A(A[185]), .B(B[185]), .CI(
        C[185]), .S(S[185]), .CO(C[186]) );
  FA_16518 \FA_INST_0[0].FA_INST_1[186].FA_  ( .A(A[186]), .B(B[186]), .CI(
        C[186]), .S(S[186]), .CO(C[187]) );
  FA_16517 \FA_INST_0[0].FA_INST_1[187].FA_  ( .A(A[187]), .B(B[187]), .CI(
        C[187]), .S(S[187]), .CO(C[188]) );
  FA_16516 \FA_INST_0[0].FA_INST_1[188].FA_  ( .A(A[188]), .B(B[188]), .CI(
        C[188]), .S(S[188]), .CO(C[189]) );
  FA_16515 \FA_INST_0[0].FA_INST_1[189].FA_  ( .A(A[189]), .B(B[189]), .CI(
        C[189]), .S(S[189]), .CO(C[190]) );
  FA_16514 \FA_INST_0[0].FA_INST_1[190].FA_  ( .A(A[190]), .B(B[190]), .CI(
        C[190]), .S(S[190]), .CO(C[191]) );
  FA_16513 \FA_INST_0[0].FA_INST_1[191].FA_  ( .A(A[191]), .B(B[191]), .CI(
        C[191]), .S(S[191]), .CO(C[192]) );
  FA_16512 \FA_INST_0[0].FA_INST_1[192].FA_  ( .A(A[192]), .B(B[192]), .CI(
        C[192]), .S(S[192]), .CO(C[193]) );
  FA_16511 \FA_INST_0[0].FA_INST_1[193].FA_  ( .A(A[193]), .B(B[193]), .CI(
        C[193]), .S(S[193]), .CO(C[194]) );
  FA_16510 \FA_INST_0[0].FA_INST_1[194].FA_  ( .A(A[194]), .B(B[194]), .CI(
        C[194]), .S(S[194]), .CO(C[195]) );
  FA_16509 \FA_INST_0[0].FA_INST_1[195].FA_  ( .A(A[195]), .B(B[195]), .CI(
        C[195]), .S(S[195]), .CO(C[196]) );
  FA_16508 \FA_INST_0[0].FA_INST_1[196].FA_  ( .A(A[196]), .B(B[196]), .CI(
        C[196]), .S(S[196]), .CO(C[197]) );
  FA_16507 \FA_INST_0[0].FA_INST_1[197].FA_  ( .A(A[197]), .B(B[197]), .CI(
        C[197]), .S(S[197]), .CO(C[198]) );
  FA_16506 \FA_INST_0[0].FA_INST_1[198].FA_  ( .A(A[198]), .B(B[198]), .CI(
        C[198]), .S(S[198]), .CO(C[199]) );
  FA_16505 \FA_INST_0[0].FA_INST_1[199].FA_  ( .A(A[199]), .B(B[199]), .CI(
        C[199]), .S(S[199]), .CO(C[200]) );
  FA_16504 \FA_INST_0[0].FA_INST_1[200].FA_  ( .A(A[200]), .B(B[200]), .CI(
        C[200]), .S(S[200]), .CO(C[201]) );
  FA_16503 \FA_INST_0[0].FA_INST_1[201].FA_  ( .A(A[201]), .B(B[201]), .CI(
        C[201]), .S(S[201]), .CO(C[202]) );
  FA_16502 \FA_INST_0[0].FA_INST_1[202].FA_  ( .A(A[202]), .B(B[202]), .CI(
        C[202]), .S(S[202]), .CO(C[203]) );
  FA_16501 \FA_INST_0[0].FA_INST_1[203].FA_  ( .A(A[203]), .B(B[203]), .CI(
        C[203]), .S(S[203]), .CO(C[204]) );
  FA_16500 \FA_INST_0[0].FA_INST_1[204].FA_  ( .A(A[204]), .B(B[204]), .CI(
        C[204]), .S(S[204]), .CO(C[205]) );
  FA_16499 \FA_INST_0[0].FA_INST_1[205].FA_  ( .A(A[205]), .B(B[205]), .CI(
        C[205]), .S(S[205]), .CO(C[206]) );
  FA_16498 \FA_INST_0[0].FA_INST_1[206].FA_  ( .A(A[206]), .B(B[206]), .CI(
        C[206]), .S(S[206]), .CO(C[207]) );
  FA_16497 \FA_INST_0[0].FA_INST_1[207].FA_  ( .A(A[207]), .B(B[207]), .CI(
        C[207]), .S(S[207]), .CO(C[208]) );
  FA_16496 \FA_INST_0[0].FA_INST_1[208].FA_  ( .A(A[208]), .B(B[208]), .CI(
        C[208]), .S(S[208]), .CO(C[209]) );
  FA_16495 \FA_INST_0[0].FA_INST_1[209].FA_  ( .A(A[209]), .B(B[209]), .CI(
        C[209]), .S(S[209]), .CO(C[210]) );
  FA_16494 \FA_INST_0[0].FA_INST_1[210].FA_  ( .A(A[210]), .B(B[210]), .CI(
        C[210]), .S(S[210]), .CO(C[211]) );
  FA_16493 \FA_INST_0[0].FA_INST_1[211].FA_  ( .A(A[211]), .B(B[211]), .CI(
        C[211]), .S(S[211]), .CO(C[212]) );
  FA_16492 \FA_INST_0[0].FA_INST_1[212].FA_  ( .A(A[212]), .B(B[212]), .CI(
        C[212]), .S(S[212]), .CO(C[213]) );
  FA_16491 \FA_INST_0[0].FA_INST_1[213].FA_  ( .A(A[213]), .B(B[213]), .CI(
        C[213]), .S(S[213]), .CO(C[214]) );
  FA_16490 \FA_INST_0[0].FA_INST_1[214].FA_  ( .A(A[214]), .B(B[214]), .CI(
        C[214]), .S(S[214]), .CO(C[215]) );
  FA_16489 \FA_INST_0[0].FA_INST_1[215].FA_  ( .A(A[215]), .B(B[215]), .CI(
        C[215]), .S(S[215]), .CO(C[216]) );
  FA_16488 \FA_INST_0[0].FA_INST_1[216].FA_  ( .A(A[216]), .B(B[216]), .CI(
        C[216]), .S(S[216]), .CO(C[217]) );
  FA_16487 \FA_INST_0[0].FA_INST_1[217].FA_  ( .A(A[217]), .B(B[217]), .CI(
        C[217]), .S(S[217]), .CO(C[218]) );
  FA_16486 \FA_INST_0[0].FA_INST_1[218].FA_  ( .A(A[218]), .B(B[218]), .CI(
        C[218]), .S(S[218]), .CO(C[219]) );
  FA_16485 \FA_INST_0[0].FA_INST_1[219].FA_  ( .A(A[219]), .B(B[219]), .CI(
        C[219]), .S(S[219]), .CO(C[220]) );
  FA_16484 \FA_INST_0[0].FA_INST_1[220].FA_  ( .A(A[220]), .B(B[220]), .CI(
        C[220]), .S(S[220]), .CO(C[221]) );
  FA_16483 \FA_INST_0[0].FA_INST_1[221].FA_  ( .A(A[221]), .B(B[221]), .CI(
        C[221]), .S(S[221]), .CO(C[222]) );
  FA_16482 \FA_INST_0[0].FA_INST_1[222].FA_  ( .A(A[222]), .B(B[222]), .CI(
        C[222]), .S(S[222]), .CO(C[223]) );
  FA_16481 \FA_INST_0[0].FA_INST_1[223].FA_  ( .A(A[223]), .B(B[223]), .CI(
        C[223]), .S(S[223]), .CO(C[224]) );
  FA_16480 \FA_INST_0[0].FA_INST_1[224].FA_  ( .A(A[224]), .B(B[224]), .CI(
        C[224]), .S(S[224]), .CO(C[225]) );
  FA_16479 \FA_INST_0[0].FA_INST_1[225].FA_  ( .A(A[225]), .B(B[225]), .CI(
        C[225]), .S(S[225]), .CO(C[226]) );
  FA_16478 \FA_INST_0[0].FA_INST_1[226].FA_  ( .A(A[226]), .B(B[226]), .CI(
        C[226]), .S(S[226]), .CO(C[227]) );
  FA_16477 \FA_INST_0[0].FA_INST_1[227].FA_  ( .A(A[227]), .B(B[227]), .CI(
        C[227]), .S(S[227]), .CO(C[228]) );
  FA_16476 \FA_INST_0[0].FA_INST_1[228].FA_  ( .A(A[228]), .B(B[228]), .CI(
        C[228]), .S(S[228]), .CO(C[229]) );
  FA_16475 \FA_INST_0[0].FA_INST_1[229].FA_  ( .A(A[229]), .B(B[229]), .CI(
        C[229]), .S(S[229]), .CO(C[230]) );
  FA_16474 \FA_INST_0[0].FA_INST_1[230].FA_  ( .A(A[230]), .B(B[230]), .CI(
        C[230]), .S(S[230]), .CO(C[231]) );
  FA_16473 \FA_INST_0[0].FA_INST_1[231].FA_  ( .A(A[231]), .B(B[231]), .CI(
        C[231]), .S(S[231]), .CO(C[232]) );
  FA_16472 \FA_INST_0[0].FA_INST_1[232].FA_  ( .A(A[232]), .B(B[232]), .CI(
        C[232]), .S(S[232]), .CO(C[233]) );
  FA_16471 \FA_INST_0[0].FA_INST_1[233].FA_  ( .A(A[233]), .B(B[233]), .CI(
        C[233]), .S(S[233]), .CO(C[234]) );
  FA_16470 \FA_INST_0[0].FA_INST_1[234].FA_  ( .A(A[234]), .B(B[234]), .CI(
        C[234]), .S(S[234]), .CO(C[235]) );
  FA_16469 \FA_INST_0[0].FA_INST_1[235].FA_  ( .A(A[235]), .B(B[235]), .CI(
        C[235]), .S(S[235]), .CO(C[236]) );
  FA_16468 \FA_INST_0[0].FA_INST_1[236].FA_  ( .A(A[236]), .B(B[236]), .CI(
        C[236]), .S(S[236]), .CO(C[237]) );
  FA_16467 \FA_INST_0[0].FA_INST_1[237].FA_  ( .A(A[237]), .B(B[237]), .CI(
        C[237]), .S(S[237]), .CO(C[238]) );
  FA_16466 \FA_INST_0[0].FA_INST_1[238].FA_  ( .A(A[238]), .B(B[238]), .CI(
        C[238]), .S(S[238]), .CO(C[239]) );
  FA_16465 \FA_INST_0[0].FA_INST_1[239].FA_  ( .A(A[239]), .B(B[239]), .CI(
        C[239]), .S(S[239]), .CO(C[240]) );
  FA_16464 \FA_INST_0[0].FA_INST_1[240].FA_  ( .A(A[240]), .B(B[240]), .CI(
        C[240]), .S(S[240]), .CO(C[241]) );
  FA_16463 \FA_INST_0[0].FA_INST_1[241].FA_  ( .A(A[241]), .B(B[241]), .CI(
        C[241]), .S(S[241]), .CO(C[242]) );
  FA_16462 \FA_INST_0[0].FA_INST_1[242].FA_  ( .A(A[242]), .B(B[242]), .CI(
        C[242]), .S(S[242]), .CO(C[243]) );
  FA_16461 \FA_INST_0[0].FA_INST_1[243].FA_  ( .A(A[243]), .B(B[243]), .CI(
        C[243]), .S(S[243]), .CO(C[244]) );
  FA_16460 \FA_INST_0[0].FA_INST_1[244].FA_  ( .A(A[244]), .B(B[244]), .CI(
        C[244]), .S(S[244]), .CO(C[245]) );
  FA_16459 \FA_INST_0[0].FA_INST_1[245].FA_  ( .A(A[245]), .B(B[245]), .CI(
        C[245]), .S(S[245]), .CO(C[246]) );
  FA_16458 \FA_INST_0[0].FA_INST_1[246].FA_  ( .A(A[246]), .B(B[246]), .CI(
        C[246]), .S(S[246]), .CO(C[247]) );
  FA_16457 \FA_INST_0[0].FA_INST_1[247].FA_  ( .A(A[247]), .B(B[247]), .CI(
        C[247]), .S(S[247]), .CO(C[248]) );
  FA_16456 \FA_INST_0[0].FA_INST_1[248].FA_  ( .A(A[248]), .B(B[248]), .CI(
        C[248]), .S(S[248]), .CO(C[249]) );
  FA_16455 \FA_INST_0[0].FA_INST_1[249].FA_  ( .A(A[249]), .B(B[249]), .CI(
        C[249]), .S(S[249]), .CO(C[250]) );
  FA_16454 \FA_INST_0[0].FA_INST_1[250].FA_  ( .A(A[250]), .B(B[250]), .CI(
        C[250]), .S(S[250]), .CO(C[251]) );
  FA_16453 \FA_INST_0[0].FA_INST_1[251].FA_  ( .A(A[251]), .B(B[251]), .CI(
        C[251]), .S(S[251]), .CO(C[252]) );
  FA_16452 \FA_INST_0[0].FA_INST_1[252].FA_  ( .A(A[252]), .B(B[252]), .CI(
        C[252]), .S(S[252]), .CO(C[253]) );
  FA_16451 \FA_INST_0[0].FA_INST_1[253].FA_  ( .A(A[253]), .B(B[253]), .CI(
        C[253]), .S(S[253]), .CO(C[254]) );
  FA_16450 \FA_INST_0[0].FA_INST_1[254].FA_  ( .A(A[254]), .B(B[254]), .CI(
        C[254]), .S(S[254]), .CO(C[255]) );
  FA_16449 \FA_INST_0[0].FA_INST_1[255].FA_  ( .A(A[255]), .B(B[255]), .CI(
        C[255]), .S(S[255]), .CO(C[256]) );
  FA_16448 \FA_INST_0[0].FA_INST_1[256].FA_  ( .A(A[256]), .B(B[256]), .CI(
        C[256]), .S(S[256]), .CO(C[257]) );
  FA_16447 \FA_INST_0[0].FA_INST_1[257].FA_  ( .A(A[257]), .B(B[257]), .CI(
        C[257]), .S(S[257]), .CO(C[258]) );
  FA_16446 \FA_INST_0[0].FA_INST_1[258].FA_  ( .A(A[258]), .B(B[258]), .CI(
        C[258]), .S(S[258]), .CO(C[259]) );
  FA_16445 \FA_INST_0[0].FA_INST_1[259].FA_  ( .A(A[259]), .B(B[259]), .CI(
        C[259]), .S(S[259]), .CO(C[260]) );
  FA_16444 \FA_INST_0[0].FA_INST_1[260].FA_  ( .A(A[260]), .B(B[260]), .CI(
        C[260]), .S(S[260]), .CO(C[261]) );
  FA_16443 \FA_INST_0[0].FA_INST_1[261].FA_  ( .A(A[261]), .B(B[261]), .CI(
        C[261]), .S(S[261]), .CO(C[262]) );
  FA_16442 \FA_INST_0[0].FA_INST_1[262].FA_  ( .A(A[262]), .B(B[262]), .CI(
        C[262]), .S(S[262]), .CO(C[263]) );
  FA_16441 \FA_INST_0[0].FA_INST_1[263].FA_  ( .A(A[263]), .B(B[263]), .CI(
        C[263]), .S(S[263]), .CO(C[264]) );
  FA_16440 \FA_INST_0[0].FA_INST_1[264].FA_  ( .A(A[264]), .B(B[264]), .CI(
        C[264]), .S(S[264]), .CO(C[265]) );
  FA_16439 \FA_INST_0[0].FA_INST_1[265].FA_  ( .A(A[265]), .B(B[265]), .CI(
        C[265]), .S(S[265]), .CO(C[266]) );
  FA_16438 \FA_INST_0[0].FA_INST_1[266].FA_  ( .A(A[266]), .B(B[266]), .CI(
        C[266]), .S(S[266]), .CO(C[267]) );
  FA_16437 \FA_INST_0[0].FA_INST_1[267].FA_  ( .A(A[267]), .B(B[267]), .CI(
        C[267]), .S(S[267]), .CO(C[268]) );
  FA_16436 \FA_INST_0[0].FA_INST_1[268].FA_  ( .A(A[268]), .B(B[268]), .CI(
        C[268]), .S(S[268]), .CO(C[269]) );
  FA_16435 \FA_INST_0[0].FA_INST_1[269].FA_  ( .A(A[269]), .B(B[269]), .CI(
        C[269]), .S(S[269]), .CO(C[270]) );
  FA_16434 \FA_INST_0[0].FA_INST_1[270].FA_  ( .A(A[270]), .B(B[270]), .CI(
        C[270]), .S(S[270]), .CO(C[271]) );
  FA_16433 \FA_INST_0[0].FA_INST_1[271].FA_  ( .A(A[271]), .B(B[271]), .CI(
        C[271]), .S(S[271]), .CO(C[272]) );
  FA_16432 \FA_INST_0[0].FA_INST_1[272].FA_  ( .A(A[272]), .B(B[272]), .CI(
        C[272]), .S(S[272]), .CO(C[273]) );
  FA_16431 \FA_INST_0[0].FA_INST_1[273].FA_  ( .A(A[273]), .B(B[273]), .CI(
        C[273]), .S(S[273]), .CO(C[274]) );
  FA_16430 \FA_INST_0[0].FA_INST_1[274].FA_  ( .A(A[274]), .B(B[274]), .CI(
        C[274]), .S(S[274]), .CO(C[275]) );
  FA_16429 \FA_INST_0[0].FA_INST_1[275].FA_  ( .A(A[275]), .B(B[275]), .CI(
        C[275]), .S(S[275]), .CO(C[276]) );
  FA_16428 \FA_INST_0[0].FA_INST_1[276].FA_  ( .A(A[276]), .B(B[276]), .CI(
        C[276]), .S(S[276]), .CO(C[277]) );
  FA_16427 \FA_INST_0[0].FA_INST_1[277].FA_  ( .A(A[277]), .B(B[277]), .CI(
        C[277]), .S(S[277]), .CO(C[278]) );
  FA_16426 \FA_INST_0[0].FA_INST_1[278].FA_  ( .A(A[278]), .B(B[278]), .CI(
        C[278]), .S(S[278]), .CO(C[279]) );
  FA_16425 \FA_INST_0[0].FA_INST_1[279].FA_  ( .A(A[279]), .B(B[279]), .CI(
        C[279]), .S(S[279]), .CO(C[280]) );
  FA_16424 \FA_INST_0[0].FA_INST_1[280].FA_  ( .A(A[280]), .B(B[280]), .CI(
        C[280]), .S(S[280]), .CO(C[281]) );
  FA_16423 \FA_INST_0[0].FA_INST_1[281].FA_  ( .A(A[281]), .B(B[281]), .CI(
        C[281]), .S(S[281]), .CO(C[282]) );
  FA_16422 \FA_INST_0[0].FA_INST_1[282].FA_  ( .A(A[282]), .B(B[282]), .CI(
        C[282]), .S(S[282]), .CO(C[283]) );
  FA_16421 \FA_INST_0[0].FA_INST_1[283].FA_  ( .A(A[283]), .B(B[283]), .CI(
        C[283]), .S(S[283]), .CO(C[284]) );
  FA_16420 \FA_INST_0[0].FA_INST_1[284].FA_  ( .A(A[284]), .B(B[284]), .CI(
        C[284]), .S(S[284]), .CO(C[285]) );
  FA_16419 \FA_INST_0[0].FA_INST_1[285].FA_  ( .A(A[285]), .B(B[285]), .CI(
        C[285]), .S(S[285]), .CO(C[286]) );
  FA_16418 \FA_INST_0[0].FA_INST_1[286].FA_  ( .A(A[286]), .B(B[286]), .CI(
        C[286]), .S(S[286]), .CO(C[287]) );
  FA_16417 \FA_INST_0[0].FA_INST_1[287].FA_  ( .A(A[287]), .B(B[287]), .CI(
        C[287]), .S(S[287]), .CO(C[288]) );
  FA_16416 \FA_INST_0[0].FA_INST_1[288].FA_  ( .A(A[288]), .B(B[288]), .CI(
        C[288]), .S(S[288]), .CO(C[289]) );
  FA_16415 \FA_INST_0[0].FA_INST_1[289].FA_  ( .A(A[289]), .B(B[289]), .CI(
        C[289]), .S(S[289]), .CO(C[290]) );
  FA_16414 \FA_INST_0[0].FA_INST_1[290].FA_  ( .A(A[290]), .B(B[290]), .CI(
        C[290]), .S(S[290]), .CO(C[291]) );
  FA_16413 \FA_INST_0[0].FA_INST_1[291].FA_  ( .A(A[291]), .B(B[291]), .CI(
        C[291]), .S(S[291]), .CO(C[292]) );
  FA_16412 \FA_INST_0[0].FA_INST_1[292].FA_  ( .A(A[292]), .B(B[292]), .CI(
        C[292]), .S(S[292]), .CO(C[293]) );
  FA_16411 \FA_INST_0[0].FA_INST_1[293].FA_  ( .A(A[293]), .B(B[293]), .CI(
        C[293]), .S(S[293]), .CO(C[294]) );
  FA_16410 \FA_INST_0[0].FA_INST_1[294].FA_  ( .A(A[294]), .B(B[294]), .CI(
        C[294]), .S(S[294]), .CO(C[295]) );
  FA_16409 \FA_INST_0[0].FA_INST_1[295].FA_  ( .A(A[295]), .B(B[295]), .CI(
        C[295]), .S(S[295]), .CO(C[296]) );
  FA_16408 \FA_INST_0[0].FA_INST_1[296].FA_  ( .A(A[296]), .B(B[296]), .CI(
        C[296]), .S(S[296]), .CO(C[297]) );
  FA_16407 \FA_INST_0[0].FA_INST_1[297].FA_  ( .A(A[297]), .B(B[297]), .CI(
        C[297]), .S(S[297]), .CO(C[298]) );
  FA_16406 \FA_INST_0[0].FA_INST_1[298].FA_  ( .A(A[298]), .B(B[298]), .CI(
        C[298]), .S(S[298]), .CO(C[299]) );
  FA_16405 \FA_INST_0[0].FA_INST_1[299].FA_  ( .A(A[299]), .B(B[299]), .CI(
        C[299]), .S(S[299]), .CO(C[300]) );
  FA_16404 \FA_INST_0[0].FA_INST_1[300].FA_  ( .A(A[300]), .B(B[300]), .CI(
        C[300]), .S(S[300]), .CO(C[301]) );
  FA_16403 \FA_INST_0[0].FA_INST_1[301].FA_  ( .A(A[301]), .B(B[301]), .CI(
        C[301]), .S(S[301]), .CO(C[302]) );
  FA_16402 \FA_INST_0[0].FA_INST_1[302].FA_  ( .A(A[302]), .B(B[302]), .CI(
        C[302]), .S(S[302]), .CO(C[303]) );
  FA_16401 \FA_INST_0[0].FA_INST_1[303].FA_  ( .A(A[303]), .B(B[303]), .CI(
        C[303]), .S(S[303]), .CO(C[304]) );
  FA_16400 \FA_INST_0[0].FA_INST_1[304].FA_  ( .A(A[304]), .B(B[304]), .CI(
        C[304]), .S(S[304]), .CO(C[305]) );
  FA_16399 \FA_INST_0[0].FA_INST_1[305].FA_  ( .A(A[305]), .B(B[305]), .CI(
        C[305]), .S(S[305]), .CO(C[306]) );
  FA_16398 \FA_INST_0[0].FA_INST_1[306].FA_  ( .A(A[306]), .B(B[306]), .CI(
        C[306]), .S(S[306]), .CO(C[307]) );
  FA_16397 \FA_INST_0[0].FA_INST_1[307].FA_  ( .A(A[307]), .B(B[307]), .CI(
        C[307]), .S(S[307]), .CO(C[308]) );
  FA_16396 \FA_INST_0[0].FA_INST_1[308].FA_  ( .A(A[308]), .B(B[308]), .CI(
        C[308]), .S(S[308]), .CO(C[309]) );
  FA_16395 \FA_INST_0[0].FA_INST_1[309].FA_  ( .A(A[309]), .B(B[309]), .CI(
        C[309]), .S(S[309]), .CO(C[310]) );
  FA_16394 \FA_INST_0[0].FA_INST_1[310].FA_  ( .A(A[310]), .B(B[310]), .CI(
        C[310]), .S(S[310]), .CO(C[311]) );
  FA_16393 \FA_INST_0[0].FA_INST_1[311].FA_  ( .A(A[311]), .B(B[311]), .CI(
        C[311]), .S(S[311]), .CO(C[312]) );
  FA_16392 \FA_INST_0[0].FA_INST_1[312].FA_  ( .A(A[312]), .B(B[312]), .CI(
        C[312]), .S(S[312]), .CO(C[313]) );
  FA_16391 \FA_INST_0[0].FA_INST_1[313].FA_  ( .A(A[313]), .B(B[313]), .CI(
        C[313]), .S(S[313]), .CO(C[314]) );
  FA_16390 \FA_INST_0[0].FA_INST_1[314].FA_  ( .A(A[314]), .B(B[314]), .CI(
        C[314]), .S(S[314]), .CO(C[315]) );
  FA_16389 \FA_INST_0[0].FA_INST_1[315].FA_  ( .A(A[315]), .B(B[315]), .CI(
        C[315]), .S(S[315]), .CO(C[316]) );
  FA_16388 \FA_INST_0[0].FA_INST_1[316].FA_  ( .A(A[316]), .B(B[316]), .CI(
        C[316]), .S(S[316]), .CO(C[317]) );
  FA_16387 \FA_INST_0[0].FA_INST_1[317].FA_  ( .A(A[317]), .B(B[317]), .CI(
        C[317]), .S(S[317]), .CO(C[318]) );
  FA_16386 \FA_INST_0[0].FA_INST_1[318].FA_  ( .A(A[318]), .B(B[318]), .CI(
        C[318]), .S(S[318]), .CO(C[319]) );
  FA_16385 \FA_INST_0[0].FA_INST_1[319].FA_  ( .A(A[319]), .B(B[319]), .CI(
        C[319]), .S(S[319]), .CO(C[320]) );
  FA_16384 \FA_INST_0[0].FA_INST_1[320].FA_  ( .A(A[320]), .B(B[320]), .CI(
        C[320]), .S(S[320]), .CO(C[321]) );
  FA_16383 \FA_INST_0[0].FA_INST_1[321].FA_  ( .A(A[321]), .B(B[321]), .CI(
        C[321]), .S(S[321]), .CO(C[322]) );
  FA_16382 \FA_INST_0[0].FA_INST_1[322].FA_  ( .A(A[322]), .B(B[322]), .CI(
        C[322]), .S(S[322]), .CO(C[323]) );
  FA_16381 \FA_INST_0[0].FA_INST_1[323].FA_  ( .A(A[323]), .B(B[323]), .CI(
        C[323]), .S(S[323]), .CO(C[324]) );
  FA_16380 \FA_INST_0[0].FA_INST_1[324].FA_  ( .A(A[324]), .B(B[324]), .CI(
        C[324]), .S(S[324]), .CO(C[325]) );
  FA_16379 \FA_INST_0[0].FA_INST_1[325].FA_  ( .A(A[325]), .B(B[325]), .CI(
        C[325]), .S(S[325]), .CO(C[326]) );
  FA_16378 \FA_INST_0[0].FA_INST_1[326].FA_  ( .A(A[326]), .B(B[326]), .CI(
        C[326]), .S(S[326]), .CO(C[327]) );
  FA_16377 \FA_INST_0[0].FA_INST_1[327].FA_  ( .A(A[327]), .B(B[327]), .CI(
        C[327]), .S(S[327]), .CO(C[328]) );
  FA_16376 \FA_INST_0[0].FA_INST_1[328].FA_  ( .A(A[328]), .B(B[328]), .CI(
        C[328]), .S(S[328]), .CO(C[329]) );
  FA_16375 \FA_INST_0[0].FA_INST_1[329].FA_  ( .A(A[329]), .B(B[329]), .CI(
        C[329]), .S(S[329]), .CO(C[330]) );
  FA_16374 \FA_INST_0[0].FA_INST_1[330].FA_  ( .A(A[330]), .B(B[330]), .CI(
        C[330]), .S(S[330]), .CO(C[331]) );
  FA_16373 \FA_INST_0[0].FA_INST_1[331].FA_  ( .A(A[331]), .B(B[331]), .CI(
        C[331]), .S(S[331]), .CO(C[332]) );
  FA_16372 \FA_INST_0[0].FA_INST_1[332].FA_  ( .A(A[332]), .B(B[332]), .CI(
        C[332]), .S(S[332]), .CO(C[333]) );
  FA_16371 \FA_INST_0[0].FA_INST_1[333].FA_  ( .A(A[333]), .B(B[333]), .CI(
        C[333]), .S(S[333]), .CO(C[334]) );
  FA_16370 \FA_INST_0[0].FA_INST_1[334].FA_  ( .A(A[334]), .B(B[334]), .CI(
        C[334]), .S(S[334]), .CO(C[335]) );
  FA_16369 \FA_INST_0[0].FA_INST_1[335].FA_  ( .A(A[335]), .B(B[335]), .CI(
        C[335]), .S(S[335]), .CO(C[336]) );
  FA_16368 \FA_INST_0[0].FA_INST_1[336].FA_  ( .A(A[336]), .B(B[336]), .CI(
        C[336]), .S(S[336]), .CO(C[337]) );
  FA_16367 \FA_INST_0[0].FA_INST_1[337].FA_  ( .A(A[337]), .B(B[337]), .CI(
        C[337]), .S(S[337]), .CO(C[338]) );
  FA_16366 \FA_INST_0[0].FA_INST_1[338].FA_  ( .A(A[338]), .B(B[338]), .CI(
        C[338]), .S(S[338]), .CO(C[339]) );
  FA_16365 \FA_INST_0[0].FA_INST_1[339].FA_  ( .A(A[339]), .B(B[339]), .CI(
        C[339]), .S(S[339]), .CO(C[340]) );
  FA_16364 \FA_INST_0[0].FA_INST_1[340].FA_  ( .A(A[340]), .B(B[340]), .CI(
        C[340]), .S(S[340]), .CO(C[341]) );
  FA_16363 \FA_INST_0[0].FA_INST_1[341].FA_  ( .A(A[341]), .B(B[341]), .CI(
        C[341]), .S(S[341]), .CO(C[342]) );
  FA_16362 \FA_INST_0[0].FA_INST_1[342].FA_  ( .A(A[342]), .B(B[342]), .CI(
        C[342]), .S(S[342]), .CO(C[343]) );
  FA_16361 \FA_INST_0[0].FA_INST_1[343].FA_  ( .A(A[343]), .B(B[343]), .CI(
        C[343]), .S(S[343]), .CO(C[344]) );
  FA_16360 \FA_INST_0[0].FA_INST_1[344].FA_  ( .A(A[344]), .B(B[344]), .CI(
        C[344]), .S(S[344]), .CO(C[345]) );
  FA_16359 \FA_INST_0[0].FA_INST_1[345].FA_  ( .A(A[345]), .B(B[345]), .CI(
        C[345]), .S(S[345]), .CO(C[346]) );
  FA_16358 \FA_INST_0[0].FA_INST_1[346].FA_  ( .A(A[346]), .B(B[346]), .CI(
        C[346]), .S(S[346]), .CO(C[347]) );
  FA_16357 \FA_INST_0[0].FA_INST_1[347].FA_  ( .A(A[347]), .B(B[347]), .CI(
        C[347]), .S(S[347]), .CO(C[348]) );
  FA_16356 \FA_INST_0[0].FA_INST_1[348].FA_  ( .A(A[348]), .B(B[348]), .CI(
        C[348]), .S(S[348]), .CO(C[349]) );
  FA_16355 \FA_INST_0[0].FA_INST_1[349].FA_  ( .A(A[349]), .B(B[349]), .CI(
        C[349]), .S(S[349]), .CO(C[350]) );
  FA_16354 \FA_INST_0[0].FA_INST_1[350].FA_  ( .A(A[350]), .B(B[350]), .CI(
        C[350]), .S(S[350]), .CO(C[351]) );
  FA_16353 \FA_INST_0[0].FA_INST_1[351].FA_  ( .A(A[351]), .B(B[351]), .CI(
        C[351]), .S(S[351]), .CO(C[352]) );
  FA_16352 \FA_INST_0[0].FA_INST_1[352].FA_  ( .A(A[352]), .B(B[352]), .CI(
        C[352]), .S(S[352]), .CO(C[353]) );
  FA_16351 \FA_INST_0[0].FA_INST_1[353].FA_  ( .A(A[353]), .B(B[353]), .CI(
        C[353]), .S(S[353]), .CO(C[354]) );
  FA_16350 \FA_INST_0[0].FA_INST_1[354].FA_  ( .A(A[354]), .B(B[354]), .CI(
        C[354]), .S(S[354]), .CO(C[355]) );
  FA_16349 \FA_INST_0[0].FA_INST_1[355].FA_  ( .A(A[355]), .B(B[355]), .CI(
        C[355]), .S(S[355]), .CO(C[356]) );
  FA_16348 \FA_INST_0[0].FA_INST_1[356].FA_  ( .A(A[356]), .B(B[356]), .CI(
        C[356]), .S(S[356]), .CO(C[357]) );
  FA_16347 \FA_INST_0[0].FA_INST_1[357].FA_  ( .A(A[357]), .B(B[357]), .CI(
        C[357]), .S(S[357]), .CO(C[358]) );
  FA_16346 \FA_INST_0[0].FA_INST_1[358].FA_  ( .A(A[358]), .B(B[358]), .CI(
        C[358]), .S(S[358]), .CO(C[359]) );
  FA_16345 \FA_INST_0[0].FA_INST_1[359].FA_  ( .A(A[359]), .B(B[359]), .CI(
        C[359]), .S(S[359]), .CO(C[360]) );
  FA_16344 \FA_INST_0[0].FA_INST_1[360].FA_  ( .A(A[360]), .B(B[360]), .CI(
        C[360]), .S(S[360]), .CO(C[361]) );
  FA_16343 \FA_INST_0[0].FA_INST_1[361].FA_  ( .A(A[361]), .B(B[361]), .CI(
        C[361]), .S(S[361]), .CO(C[362]) );
  FA_16342 \FA_INST_0[0].FA_INST_1[362].FA_  ( .A(A[362]), .B(B[362]), .CI(
        C[362]), .S(S[362]), .CO(C[363]) );
  FA_16341 \FA_INST_0[0].FA_INST_1[363].FA_  ( .A(A[363]), .B(B[363]), .CI(
        C[363]), .S(S[363]), .CO(C[364]) );
  FA_16340 \FA_INST_0[0].FA_INST_1[364].FA_  ( .A(A[364]), .B(B[364]), .CI(
        C[364]), .S(S[364]), .CO(C[365]) );
  FA_16339 \FA_INST_0[0].FA_INST_1[365].FA_  ( .A(A[365]), .B(B[365]), .CI(
        C[365]), .S(S[365]), .CO(C[366]) );
  FA_16338 \FA_INST_0[0].FA_INST_1[366].FA_  ( .A(A[366]), .B(B[366]), .CI(
        C[366]), .S(S[366]), .CO(C[367]) );
  FA_16337 \FA_INST_0[0].FA_INST_1[367].FA_  ( .A(A[367]), .B(B[367]), .CI(
        C[367]), .S(S[367]), .CO(C[368]) );
  FA_16336 \FA_INST_0[0].FA_INST_1[368].FA_  ( .A(A[368]), .B(B[368]), .CI(
        C[368]), .S(S[368]), .CO(C[369]) );
  FA_16335 \FA_INST_0[0].FA_INST_1[369].FA_  ( .A(A[369]), .B(B[369]), .CI(
        C[369]), .S(S[369]), .CO(C[370]) );
  FA_16334 \FA_INST_0[0].FA_INST_1[370].FA_  ( .A(A[370]), .B(B[370]), .CI(
        C[370]), .S(S[370]), .CO(C[371]) );
  FA_16333 \FA_INST_0[0].FA_INST_1[371].FA_  ( .A(A[371]), .B(B[371]), .CI(
        C[371]), .S(S[371]), .CO(C[372]) );
  FA_16332 \FA_INST_0[0].FA_INST_1[372].FA_  ( .A(A[372]), .B(B[372]), .CI(
        C[372]), .S(S[372]), .CO(C[373]) );
  FA_16331 \FA_INST_0[0].FA_INST_1[373].FA_  ( .A(A[373]), .B(B[373]), .CI(
        C[373]), .S(S[373]), .CO(C[374]) );
  FA_16330 \FA_INST_0[0].FA_INST_1[374].FA_  ( .A(A[374]), .B(B[374]), .CI(
        C[374]), .S(S[374]), .CO(C[375]) );
  FA_16329 \FA_INST_0[0].FA_INST_1[375].FA_  ( .A(A[375]), .B(B[375]), .CI(
        C[375]), .S(S[375]), .CO(C[376]) );
  FA_16328 \FA_INST_0[0].FA_INST_1[376].FA_  ( .A(A[376]), .B(B[376]), .CI(
        C[376]), .S(S[376]), .CO(C[377]) );
  FA_16327 \FA_INST_0[0].FA_INST_1[377].FA_  ( .A(A[377]), .B(B[377]), .CI(
        C[377]), .S(S[377]), .CO(C[378]) );
  FA_16326 \FA_INST_0[0].FA_INST_1[378].FA_  ( .A(A[378]), .B(B[378]), .CI(
        C[378]), .S(S[378]), .CO(C[379]) );
  FA_16325 \FA_INST_0[0].FA_INST_1[379].FA_  ( .A(A[379]), .B(B[379]), .CI(
        C[379]), .S(S[379]), .CO(C[380]) );
  FA_16324 \FA_INST_0[0].FA_INST_1[380].FA_  ( .A(A[380]), .B(B[380]), .CI(
        C[380]), .S(S[380]), .CO(C[381]) );
  FA_16323 \FA_INST_0[0].FA_INST_1[381].FA_  ( .A(A[381]), .B(B[381]), .CI(
        C[381]), .S(S[381]), .CO(C[382]) );
  FA_16322 \FA_INST_0[0].FA_INST_1[382].FA_  ( .A(A[382]), .B(B[382]), .CI(
        C[382]), .S(S[382]), .CO(C[383]) );
  FA_16321 \FA_INST_0[0].FA_INST_1[383].FA_  ( .A(A[383]), .B(B[383]), .CI(
        C[383]), .S(S[383]), .CO(C[384]) );
  FA_16320 \FA_INST_0[0].FA_INST_1[384].FA_  ( .A(A[384]), .B(B[384]), .CI(
        C[384]), .S(S[384]), .CO(C[385]) );
  FA_16319 \FA_INST_0[0].FA_INST_1[385].FA_  ( .A(A[385]), .B(B[385]), .CI(
        C[385]), .S(S[385]), .CO(C[386]) );
  FA_16318 \FA_INST_0[0].FA_INST_1[386].FA_  ( .A(A[386]), .B(B[386]), .CI(
        C[386]), .S(S[386]), .CO(C[387]) );
  FA_16317 \FA_INST_0[0].FA_INST_1[387].FA_  ( .A(A[387]), .B(B[387]), .CI(
        C[387]), .S(S[387]), .CO(C[388]) );
  FA_16316 \FA_INST_0[0].FA_INST_1[388].FA_  ( .A(A[388]), .B(B[388]), .CI(
        C[388]), .S(S[388]), .CO(C[389]) );
  FA_16315 \FA_INST_0[0].FA_INST_1[389].FA_  ( .A(A[389]), .B(B[389]), .CI(
        C[389]), .S(S[389]), .CO(C[390]) );
  FA_16314 \FA_INST_0[0].FA_INST_1[390].FA_  ( .A(A[390]), .B(B[390]), .CI(
        C[390]), .S(S[390]), .CO(C[391]) );
  FA_16313 \FA_INST_0[0].FA_INST_1[391].FA_  ( .A(A[391]), .B(B[391]), .CI(
        C[391]), .S(S[391]), .CO(C[392]) );
  FA_16312 \FA_INST_0[0].FA_INST_1[392].FA_  ( .A(A[392]), .B(B[392]), .CI(
        C[392]), .S(S[392]), .CO(C[393]) );
  FA_16311 \FA_INST_0[0].FA_INST_1[393].FA_  ( .A(A[393]), .B(B[393]), .CI(
        C[393]), .S(S[393]), .CO(C[394]) );
  FA_16310 \FA_INST_0[0].FA_INST_1[394].FA_  ( .A(A[394]), .B(B[394]), .CI(
        C[394]), .S(S[394]), .CO(C[395]) );
  FA_16309 \FA_INST_0[0].FA_INST_1[395].FA_  ( .A(A[395]), .B(B[395]), .CI(
        C[395]), .S(S[395]), .CO(C[396]) );
  FA_16308 \FA_INST_0[0].FA_INST_1[396].FA_  ( .A(A[396]), .B(B[396]), .CI(
        C[396]), .S(S[396]), .CO(C[397]) );
  FA_16307 \FA_INST_0[0].FA_INST_1[397].FA_  ( .A(A[397]), .B(B[397]), .CI(
        C[397]), .S(S[397]), .CO(C[398]) );
  FA_16306 \FA_INST_0[0].FA_INST_1[398].FA_  ( .A(A[398]), .B(B[398]), .CI(
        C[398]), .S(S[398]), .CO(C[399]) );
  FA_16305 \FA_INST_0[0].FA_INST_1[399].FA_  ( .A(A[399]), .B(B[399]), .CI(
        C[399]), .S(S[399]), .CO(C[400]) );
  FA_16304 \FA_INST_0[0].FA_INST_1[400].FA_  ( .A(A[400]), .B(B[400]), .CI(
        C[400]), .S(S[400]), .CO(C[401]) );
  FA_16303 \FA_INST_0[0].FA_INST_1[401].FA_  ( .A(A[401]), .B(B[401]), .CI(
        C[401]), .S(S[401]), .CO(C[402]) );
  FA_16302 \FA_INST_0[0].FA_INST_1[402].FA_  ( .A(A[402]), .B(B[402]), .CI(
        C[402]), .S(S[402]), .CO(C[403]) );
  FA_16301 \FA_INST_0[0].FA_INST_1[403].FA_  ( .A(A[403]), .B(B[403]), .CI(
        C[403]), .S(S[403]), .CO(C[404]) );
  FA_16300 \FA_INST_0[0].FA_INST_1[404].FA_  ( .A(A[404]), .B(B[404]), .CI(
        C[404]), .S(S[404]), .CO(C[405]) );
  FA_16299 \FA_INST_0[0].FA_INST_1[405].FA_  ( .A(A[405]), .B(B[405]), .CI(
        C[405]), .S(S[405]), .CO(C[406]) );
  FA_16298 \FA_INST_0[0].FA_INST_1[406].FA_  ( .A(A[406]), .B(B[406]), .CI(
        C[406]), .S(S[406]), .CO(C[407]) );
  FA_16297 \FA_INST_0[0].FA_INST_1[407].FA_  ( .A(A[407]), .B(B[407]), .CI(
        C[407]), .S(S[407]), .CO(C[408]) );
  FA_16296 \FA_INST_0[0].FA_INST_1[408].FA_  ( .A(A[408]), .B(B[408]), .CI(
        C[408]), .S(S[408]), .CO(C[409]) );
  FA_16295 \FA_INST_0[0].FA_INST_1[409].FA_  ( .A(A[409]), .B(B[409]), .CI(
        C[409]), .S(S[409]), .CO(C[410]) );
  FA_16294 \FA_INST_0[0].FA_INST_1[410].FA_  ( .A(A[410]), .B(B[410]), .CI(
        C[410]), .S(S[410]), .CO(C[411]) );
  FA_16293 \FA_INST_0[0].FA_INST_1[411].FA_  ( .A(A[411]), .B(B[411]), .CI(
        C[411]), .S(S[411]), .CO(C[412]) );
  FA_16292 \FA_INST_0[0].FA_INST_1[412].FA_  ( .A(A[412]), .B(B[412]), .CI(
        C[412]), .S(S[412]), .CO(C[413]) );
  FA_16291 \FA_INST_0[0].FA_INST_1[413].FA_  ( .A(A[413]), .B(B[413]), .CI(
        C[413]), .S(S[413]), .CO(C[414]) );
  FA_16290 \FA_INST_0[0].FA_INST_1[414].FA_  ( .A(A[414]), .B(B[414]), .CI(
        C[414]), .S(S[414]), .CO(C[415]) );
  FA_16289 \FA_INST_0[0].FA_INST_1[415].FA_  ( .A(A[415]), .B(B[415]), .CI(
        C[415]), .S(S[415]), .CO(C[416]) );
  FA_16288 \FA_INST_0[0].FA_INST_1[416].FA_  ( .A(A[416]), .B(B[416]), .CI(
        C[416]), .S(S[416]), .CO(C[417]) );
  FA_16287 \FA_INST_0[0].FA_INST_1[417].FA_  ( .A(A[417]), .B(B[417]), .CI(
        C[417]), .S(S[417]), .CO(C[418]) );
  FA_16286 \FA_INST_0[0].FA_INST_1[418].FA_  ( .A(A[418]), .B(B[418]), .CI(
        C[418]), .S(S[418]), .CO(C[419]) );
  FA_16285 \FA_INST_0[0].FA_INST_1[419].FA_  ( .A(A[419]), .B(B[419]), .CI(
        C[419]), .S(S[419]), .CO(C[420]) );
  FA_16284 \FA_INST_0[0].FA_INST_1[420].FA_  ( .A(A[420]), .B(B[420]), .CI(
        C[420]), .S(S[420]), .CO(C[421]) );
  FA_16283 \FA_INST_0[0].FA_INST_1[421].FA_  ( .A(A[421]), .B(B[421]), .CI(
        C[421]), .S(S[421]), .CO(C[422]) );
  FA_16282 \FA_INST_0[0].FA_INST_1[422].FA_  ( .A(A[422]), .B(B[422]), .CI(
        C[422]), .S(S[422]), .CO(C[423]) );
  FA_16281 \FA_INST_0[0].FA_INST_1[423].FA_  ( .A(A[423]), .B(B[423]), .CI(
        C[423]), .S(S[423]), .CO(C[424]) );
  FA_16280 \FA_INST_0[0].FA_INST_1[424].FA_  ( .A(A[424]), .B(B[424]), .CI(
        C[424]), .S(S[424]), .CO(C[425]) );
  FA_16279 \FA_INST_0[0].FA_INST_1[425].FA_  ( .A(A[425]), .B(B[425]), .CI(
        C[425]), .S(S[425]), .CO(C[426]) );
  FA_16278 \FA_INST_0[0].FA_INST_1[426].FA_  ( .A(A[426]), .B(B[426]), .CI(
        C[426]), .S(S[426]), .CO(C[427]) );
  FA_16277 \FA_INST_0[0].FA_INST_1[427].FA_  ( .A(A[427]), .B(B[427]), .CI(
        C[427]), .S(S[427]), .CO(C[428]) );
  FA_16276 \FA_INST_0[0].FA_INST_1[428].FA_  ( .A(A[428]), .B(B[428]), .CI(
        C[428]), .S(S[428]), .CO(C[429]) );
  FA_16275 \FA_INST_0[0].FA_INST_1[429].FA_  ( .A(A[429]), .B(B[429]), .CI(
        C[429]), .S(S[429]), .CO(C[430]) );
  FA_16274 \FA_INST_0[0].FA_INST_1[430].FA_  ( .A(A[430]), .B(B[430]), .CI(
        C[430]), .S(S[430]), .CO(C[431]) );
  FA_16273 \FA_INST_0[0].FA_INST_1[431].FA_  ( .A(A[431]), .B(B[431]), .CI(
        C[431]), .S(S[431]), .CO(C[432]) );
  FA_16272 \FA_INST_0[0].FA_INST_1[432].FA_  ( .A(A[432]), .B(B[432]), .CI(
        C[432]), .S(S[432]), .CO(C[433]) );
  FA_16271 \FA_INST_0[0].FA_INST_1[433].FA_  ( .A(A[433]), .B(B[433]), .CI(
        C[433]), .S(S[433]), .CO(C[434]) );
  FA_16270 \FA_INST_0[0].FA_INST_1[434].FA_  ( .A(A[434]), .B(B[434]), .CI(
        C[434]), .S(S[434]), .CO(C[435]) );
  FA_16269 \FA_INST_0[0].FA_INST_1[435].FA_  ( .A(A[435]), .B(B[435]), .CI(
        C[435]), .S(S[435]), .CO(C[436]) );
  FA_16268 \FA_INST_0[0].FA_INST_1[436].FA_  ( .A(A[436]), .B(B[436]), .CI(
        C[436]), .S(S[436]), .CO(C[437]) );
  FA_16267 \FA_INST_0[0].FA_INST_1[437].FA_  ( .A(A[437]), .B(B[437]), .CI(
        C[437]), .S(S[437]), .CO(C[438]) );
  FA_16266 \FA_INST_0[0].FA_INST_1[438].FA_  ( .A(A[438]), .B(B[438]), .CI(
        C[438]), .S(S[438]), .CO(C[439]) );
  FA_16265 \FA_INST_0[0].FA_INST_1[439].FA_  ( .A(A[439]), .B(B[439]), .CI(
        C[439]), .S(S[439]), .CO(C[440]) );
  FA_16264 \FA_INST_0[0].FA_INST_1[440].FA_  ( .A(A[440]), .B(B[440]), .CI(
        C[440]), .S(S[440]), .CO(C[441]) );
  FA_16263 \FA_INST_0[0].FA_INST_1[441].FA_  ( .A(A[441]), .B(B[441]), .CI(
        C[441]), .S(S[441]), .CO(C[442]) );
  FA_16262 \FA_INST_0[0].FA_INST_1[442].FA_  ( .A(A[442]), .B(B[442]), .CI(
        C[442]), .S(S[442]), .CO(C[443]) );
  FA_16261 \FA_INST_0[0].FA_INST_1[443].FA_  ( .A(A[443]), .B(B[443]), .CI(
        C[443]), .S(S[443]), .CO(C[444]) );
  FA_16260 \FA_INST_0[0].FA_INST_1[444].FA_  ( .A(A[444]), .B(B[444]), .CI(
        C[444]), .S(S[444]), .CO(C[445]) );
  FA_16259 \FA_INST_0[0].FA_INST_1[445].FA_  ( .A(A[445]), .B(B[445]), .CI(
        C[445]), .S(S[445]), .CO(C[446]) );
  FA_16258 \FA_INST_0[0].FA_INST_1[446].FA_  ( .A(A[446]), .B(B[446]), .CI(
        C[446]), .S(S[446]), .CO(C[447]) );
  FA_16257 \FA_INST_0[0].FA_INST_1[447].FA_  ( .A(A[447]), .B(B[447]), .CI(
        C[447]), .S(S[447]), .CO(C[448]) );
  FA_16256 \FA_INST_0[0].FA_INST_1[448].FA_  ( .A(A[448]), .B(B[448]), .CI(
        C[448]), .S(S[448]), .CO(C[449]) );
  FA_16255 \FA_INST_0[0].FA_INST_1[449].FA_  ( .A(A[449]), .B(B[449]), .CI(
        C[449]), .S(S[449]), .CO(C[450]) );
  FA_16254 \FA_INST_0[0].FA_INST_1[450].FA_  ( .A(A[450]), .B(B[450]), .CI(
        C[450]), .S(S[450]), .CO(C[451]) );
  FA_16253 \FA_INST_0[0].FA_INST_1[451].FA_  ( .A(A[451]), .B(B[451]), .CI(
        C[451]), .S(S[451]), .CO(C[452]) );
  FA_16252 \FA_INST_0[0].FA_INST_1[452].FA_  ( .A(A[452]), .B(B[452]), .CI(
        C[452]), .S(S[452]), .CO(C[453]) );
  FA_16251 \FA_INST_0[0].FA_INST_1[453].FA_  ( .A(A[453]), .B(B[453]), .CI(
        C[453]), .S(S[453]), .CO(C[454]) );
  FA_16250 \FA_INST_0[0].FA_INST_1[454].FA_  ( .A(A[454]), .B(B[454]), .CI(
        C[454]), .S(S[454]), .CO(C[455]) );
  FA_16249 \FA_INST_0[0].FA_INST_1[455].FA_  ( .A(A[455]), .B(B[455]), .CI(
        C[455]), .S(S[455]), .CO(C[456]) );
  FA_16248 \FA_INST_0[0].FA_INST_1[456].FA_  ( .A(A[456]), .B(B[456]), .CI(
        C[456]), .S(S[456]), .CO(C[457]) );
  FA_16247 \FA_INST_0[0].FA_INST_1[457].FA_  ( .A(A[457]), .B(B[457]), .CI(
        C[457]), .S(S[457]), .CO(C[458]) );
  FA_16246 \FA_INST_0[0].FA_INST_1[458].FA_  ( .A(A[458]), .B(B[458]), .CI(
        C[458]), .S(S[458]), .CO(C[459]) );
  FA_16245 \FA_INST_0[0].FA_INST_1[459].FA_  ( .A(A[459]), .B(B[459]), .CI(
        C[459]), .S(S[459]), .CO(C[460]) );
  FA_16244 \FA_INST_0[0].FA_INST_1[460].FA_  ( .A(A[460]), .B(B[460]), .CI(
        C[460]), .S(S[460]), .CO(C[461]) );
  FA_16243 \FA_INST_0[0].FA_INST_1[461].FA_  ( .A(A[461]), .B(B[461]), .CI(
        C[461]), .S(S[461]), .CO(C[462]) );
  FA_16242 \FA_INST_0[0].FA_INST_1[462].FA_  ( .A(A[462]), .B(B[462]), .CI(
        C[462]), .S(S[462]), .CO(C[463]) );
  FA_16241 \FA_INST_0[0].FA_INST_1[463].FA_  ( .A(A[463]), .B(B[463]), .CI(
        C[463]), .S(S[463]), .CO(C[464]) );
  FA_16240 \FA_INST_0[0].FA_INST_1[464].FA_  ( .A(A[464]), .B(B[464]), .CI(
        C[464]), .S(S[464]), .CO(C[465]) );
  FA_16239 \FA_INST_0[0].FA_INST_1[465].FA_  ( .A(A[465]), .B(B[465]), .CI(
        C[465]), .S(S[465]), .CO(C[466]) );
  FA_16238 \FA_INST_0[0].FA_INST_1[466].FA_  ( .A(A[466]), .B(B[466]), .CI(
        C[466]), .S(S[466]), .CO(C[467]) );
  FA_16237 \FA_INST_0[0].FA_INST_1[467].FA_  ( .A(A[467]), .B(B[467]), .CI(
        C[467]), .S(S[467]), .CO(C[468]) );
  FA_16236 \FA_INST_0[0].FA_INST_1[468].FA_  ( .A(A[468]), .B(B[468]), .CI(
        C[468]), .S(S[468]), .CO(C[469]) );
  FA_16235 \FA_INST_0[0].FA_INST_1[469].FA_  ( .A(A[469]), .B(B[469]), .CI(
        C[469]), .S(S[469]), .CO(C[470]) );
  FA_16234 \FA_INST_0[0].FA_INST_1[470].FA_  ( .A(A[470]), .B(B[470]), .CI(
        C[470]), .S(S[470]), .CO(C[471]) );
  FA_16233 \FA_INST_0[0].FA_INST_1[471].FA_  ( .A(A[471]), .B(B[471]), .CI(
        C[471]), .S(S[471]), .CO(C[472]) );
  FA_16232 \FA_INST_0[0].FA_INST_1[472].FA_  ( .A(A[472]), .B(B[472]), .CI(
        C[472]), .S(S[472]), .CO(C[473]) );
  FA_16231 \FA_INST_0[0].FA_INST_1[473].FA_  ( .A(A[473]), .B(B[473]), .CI(
        C[473]), .S(S[473]), .CO(C[474]) );
  FA_16230 \FA_INST_0[0].FA_INST_1[474].FA_  ( .A(A[474]), .B(B[474]), .CI(
        C[474]), .S(S[474]), .CO(C[475]) );
  FA_16229 \FA_INST_0[0].FA_INST_1[475].FA_  ( .A(A[475]), .B(B[475]), .CI(
        C[475]), .S(S[475]), .CO(C[476]) );
  FA_16228 \FA_INST_0[0].FA_INST_1[476].FA_  ( .A(A[476]), .B(B[476]), .CI(
        C[476]), .S(S[476]), .CO(C[477]) );
  FA_16227 \FA_INST_0[0].FA_INST_1[477].FA_  ( .A(A[477]), .B(B[477]), .CI(
        C[477]), .S(S[477]), .CO(C[478]) );
  FA_16226 \FA_INST_0[0].FA_INST_1[478].FA_  ( .A(A[478]), .B(B[478]), .CI(
        C[478]), .S(S[478]), .CO(C[479]) );
  FA_16225 \FA_INST_0[0].FA_INST_1[479].FA_  ( .A(A[479]), .B(B[479]), .CI(
        C[479]), .S(S[479]), .CO(C[480]) );
  FA_16224 \FA_INST_0[0].FA_INST_1[480].FA_  ( .A(A[480]), .B(B[480]), .CI(
        C[480]), .S(S[480]), .CO(C[481]) );
  FA_16223 \FA_INST_0[0].FA_INST_1[481].FA_  ( .A(A[481]), .B(B[481]), .CI(
        C[481]), .S(S[481]), .CO(C[482]) );
  FA_16222 \FA_INST_0[0].FA_INST_1[482].FA_  ( .A(A[482]), .B(B[482]), .CI(
        C[482]), .S(S[482]), .CO(C[483]) );
  FA_16221 \FA_INST_0[0].FA_INST_1[483].FA_  ( .A(A[483]), .B(B[483]), .CI(
        C[483]), .S(S[483]), .CO(C[484]) );
  FA_16220 \FA_INST_0[0].FA_INST_1[484].FA_  ( .A(A[484]), .B(B[484]), .CI(
        C[484]), .S(S[484]), .CO(C[485]) );
  FA_16219 \FA_INST_0[0].FA_INST_1[485].FA_  ( .A(A[485]), .B(B[485]), .CI(
        C[485]), .S(S[485]), .CO(C[486]) );
  FA_16218 \FA_INST_0[0].FA_INST_1[486].FA_  ( .A(A[486]), .B(B[486]), .CI(
        C[486]), .S(S[486]), .CO(C[487]) );
  FA_16217 \FA_INST_0[0].FA_INST_1[487].FA_  ( .A(A[487]), .B(B[487]), .CI(
        C[487]), .S(S[487]), .CO(C[488]) );
  FA_16216 \FA_INST_0[0].FA_INST_1[488].FA_  ( .A(A[488]), .B(B[488]), .CI(
        C[488]), .S(S[488]), .CO(C[489]) );
  FA_16215 \FA_INST_0[0].FA_INST_1[489].FA_  ( .A(A[489]), .B(B[489]), .CI(
        C[489]), .S(S[489]), .CO(C[490]) );
  FA_16214 \FA_INST_0[0].FA_INST_1[490].FA_  ( .A(A[490]), .B(B[490]), .CI(
        C[490]), .S(S[490]), .CO(C[491]) );
  FA_16213 \FA_INST_0[0].FA_INST_1[491].FA_  ( .A(A[491]), .B(B[491]), .CI(
        C[491]), .S(S[491]), .CO(C[492]) );
  FA_16212 \FA_INST_0[0].FA_INST_1[492].FA_  ( .A(A[492]), .B(B[492]), .CI(
        C[492]), .S(S[492]), .CO(C[493]) );
  FA_16211 \FA_INST_0[0].FA_INST_1[493].FA_  ( .A(A[493]), .B(B[493]), .CI(
        C[493]), .S(S[493]), .CO(C[494]) );
  FA_16210 \FA_INST_0[0].FA_INST_1[494].FA_  ( .A(A[494]), .B(B[494]), .CI(
        C[494]), .S(S[494]), .CO(C[495]) );
  FA_16209 \FA_INST_0[0].FA_INST_1[495].FA_  ( .A(A[495]), .B(B[495]), .CI(
        C[495]), .S(S[495]), .CO(C[496]) );
  FA_16208 \FA_INST_0[0].FA_INST_1[496].FA_  ( .A(A[496]), .B(B[496]), .CI(
        C[496]), .S(S[496]), .CO(C[497]) );
  FA_16207 \FA_INST_0[0].FA_INST_1[497].FA_  ( .A(A[497]), .B(B[497]), .CI(
        C[497]), .S(S[497]), .CO(C[498]) );
  FA_16206 \FA_INST_0[0].FA_INST_1[498].FA_  ( .A(A[498]), .B(B[498]), .CI(
        C[498]), .S(S[498]), .CO(C[499]) );
  FA_16205 \FA_INST_0[0].FA_INST_1[499].FA_  ( .A(A[499]), .B(B[499]), .CI(
        C[499]), .S(S[499]), .CO(C[500]) );
  FA_16204 \FA_INST_0[0].FA_INST_1[500].FA_  ( .A(A[500]), .B(B[500]), .CI(
        C[500]), .S(S[500]), .CO(C[501]) );
  FA_16203 \FA_INST_0[0].FA_INST_1[501].FA_  ( .A(A[501]), .B(B[501]), .CI(
        C[501]), .S(S[501]), .CO(C[502]) );
  FA_16202 \FA_INST_0[0].FA_INST_1[502].FA_  ( .A(A[502]), .B(B[502]), .CI(
        C[502]), .S(S[502]), .CO(C[503]) );
  FA_16201 \FA_INST_0[0].FA_INST_1[503].FA_  ( .A(A[503]), .B(B[503]), .CI(
        C[503]), .S(S[503]), .CO(C[504]) );
  FA_16200 \FA_INST_0[0].FA_INST_1[504].FA_  ( .A(A[504]), .B(B[504]), .CI(
        C[504]), .S(S[504]), .CO(C[505]) );
  FA_16199 \FA_INST_0[0].FA_INST_1[505].FA_  ( .A(A[505]), .B(B[505]), .CI(
        C[505]), .S(S[505]), .CO(C[506]) );
  FA_16198 \FA_INST_0[0].FA_INST_1[506].FA_  ( .A(A[506]), .B(B[506]), .CI(
        C[506]), .S(S[506]), .CO(C[507]) );
  FA_16197 \FA_INST_0[0].FA_INST_1[507].FA_  ( .A(A[507]), .B(B[507]), .CI(
        C[507]), .S(S[507]), .CO(C[508]) );
  FA_16196 \FA_INST_0[0].FA_INST_1[508].FA_  ( .A(A[508]), .B(B[508]), .CI(
        C[508]), .S(S[508]), .CO(C[509]) );
  FA_16195 \FA_INST_0[0].FA_INST_1[509].FA_  ( .A(A[509]), .B(B[509]), .CI(
        C[509]), .S(S[509]), .CO(C[510]) );
  FA_16194 \FA_INST_0[0].FA_INST_1[510].FA_  ( .A(A[510]), .B(B[510]), .CI(
        C[510]), .S(S[510]), .CO(C[511]) );
  FA_16193 \FA_INST_0[0].FA_INST_1[511].FA_  ( .A(A[511]), .B(B[511]), .CI(
        C[511]), .S(S[511]), .CO(C[512]) );
  FA_16192 \FA_INST_0[1].FA_INST_1[0].FA_  ( .A(A[512]), .B(B[512]), .CI(
        C[512]), .S(S[512]), .CO(C[513]) );
  FA_16191 \FA_INST_0[1].FA_INST_1[1].FA_  ( .A(A[513]), .B(B[513]), .CI(
        C[513]), .S(S[513]), .CO(C[514]) );
  FA_16190 \FA_INST_0[1].FA_INST_1[2].FA_  ( .A(A[514]), .B(B[514]), .CI(
        C[514]), .S(S[514]), .CO(C[515]) );
  FA_16189 \FA_INST_0[1].FA_INST_1[3].FA_  ( .A(A[515]), .B(B[515]), .CI(
        C[515]), .S(S[515]), .CO(C[516]) );
  FA_16188 \FA_INST_0[1].FA_INST_1[4].FA_  ( .A(A[516]), .B(B[516]), .CI(
        C[516]), .S(S[516]), .CO(C[517]) );
  FA_16187 \FA_INST_0[1].FA_INST_1[5].FA_  ( .A(A[517]), .B(B[517]), .CI(
        C[517]), .S(S[517]), .CO(C[518]) );
  FA_16186 \FA_INST_0[1].FA_INST_1[6].FA_  ( .A(A[518]), .B(B[518]), .CI(
        C[518]), .S(S[518]), .CO(C[519]) );
  FA_16185 \FA_INST_0[1].FA_INST_1[7].FA_  ( .A(A[519]), .B(B[519]), .CI(
        C[519]), .S(S[519]), .CO(C[520]) );
  FA_16184 \FA_INST_0[1].FA_INST_1[8].FA_  ( .A(A[520]), .B(B[520]), .CI(
        C[520]), .S(S[520]), .CO(C[521]) );
  FA_16183 \FA_INST_0[1].FA_INST_1[9].FA_  ( .A(A[521]), .B(B[521]), .CI(
        C[521]), .S(S[521]), .CO(C[522]) );
  FA_16182 \FA_INST_0[1].FA_INST_1[10].FA_  ( .A(A[522]), .B(B[522]), .CI(
        C[522]), .S(S[522]), .CO(C[523]) );
  FA_16181 \FA_INST_0[1].FA_INST_1[11].FA_  ( .A(A[523]), .B(B[523]), .CI(
        C[523]), .S(S[523]), .CO(C[524]) );
  FA_16180 \FA_INST_0[1].FA_INST_1[12].FA_  ( .A(A[524]), .B(B[524]), .CI(
        C[524]), .S(S[524]), .CO(C[525]) );
  FA_16179 \FA_INST_0[1].FA_INST_1[13].FA_  ( .A(A[525]), .B(B[525]), .CI(
        C[525]), .S(S[525]), .CO(C[526]) );
  FA_16178 \FA_INST_0[1].FA_INST_1[14].FA_  ( .A(A[526]), .B(B[526]), .CI(
        C[526]), .S(S[526]), .CO(C[527]) );
  FA_16177 \FA_INST_0[1].FA_INST_1[15].FA_  ( .A(A[527]), .B(B[527]), .CI(
        C[527]), .S(S[527]), .CO(C[528]) );
  FA_16176 \FA_INST_0[1].FA_INST_1[16].FA_  ( .A(A[528]), .B(B[528]), .CI(
        C[528]), .S(S[528]), .CO(C[529]) );
  FA_16175 \FA_INST_0[1].FA_INST_1[17].FA_  ( .A(A[529]), .B(B[529]), .CI(
        C[529]), .S(S[529]), .CO(C[530]) );
  FA_16174 \FA_INST_0[1].FA_INST_1[18].FA_  ( .A(A[530]), .B(B[530]), .CI(
        C[530]), .S(S[530]), .CO(C[531]) );
  FA_16173 \FA_INST_0[1].FA_INST_1[19].FA_  ( .A(A[531]), .B(B[531]), .CI(
        C[531]), .S(S[531]), .CO(C[532]) );
  FA_16172 \FA_INST_0[1].FA_INST_1[20].FA_  ( .A(A[532]), .B(B[532]), .CI(
        C[532]), .S(S[532]), .CO(C[533]) );
  FA_16171 \FA_INST_0[1].FA_INST_1[21].FA_  ( .A(A[533]), .B(B[533]), .CI(
        C[533]), .S(S[533]), .CO(C[534]) );
  FA_16170 \FA_INST_0[1].FA_INST_1[22].FA_  ( .A(A[534]), .B(B[534]), .CI(
        C[534]), .S(S[534]), .CO(C[535]) );
  FA_16169 \FA_INST_0[1].FA_INST_1[23].FA_  ( .A(A[535]), .B(B[535]), .CI(
        C[535]), .S(S[535]), .CO(C[536]) );
  FA_16168 \FA_INST_0[1].FA_INST_1[24].FA_  ( .A(A[536]), .B(B[536]), .CI(
        C[536]), .S(S[536]), .CO(C[537]) );
  FA_16167 \FA_INST_0[1].FA_INST_1[25].FA_  ( .A(A[537]), .B(B[537]), .CI(
        C[537]), .S(S[537]), .CO(C[538]) );
  FA_16166 \FA_INST_0[1].FA_INST_1[26].FA_  ( .A(A[538]), .B(B[538]), .CI(
        C[538]), .S(S[538]), .CO(C[539]) );
  FA_16165 \FA_INST_0[1].FA_INST_1[27].FA_  ( .A(A[539]), .B(B[539]), .CI(
        C[539]), .S(S[539]), .CO(C[540]) );
  FA_16164 \FA_INST_0[1].FA_INST_1[28].FA_  ( .A(A[540]), .B(B[540]), .CI(
        C[540]), .S(S[540]), .CO(C[541]) );
  FA_16163 \FA_INST_0[1].FA_INST_1[29].FA_  ( .A(A[541]), .B(B[541]), .CI(
        C[541]), .S(S[541]), .CO(C[542]) );
  FA_16162 \FA_INST_0[1].FA_INST_1[30].FA_  ( .A(A[542]), .B(B[542]), .CI(
        C[542]), .S(S[542]), .CO(C[543]) );
  FA_16161 \FA_INST_0[1].FA_INST_1[31].FA_  ( .A(A[543]), .B(B[543]), .CI(
        C[543]), .S(S[543]), .CO(C[544]) );
  FA_16160 \FA_INST_0[1].FA_INST_1[32].FA_  ( .A(A[544]), .B(B[544]), .CI(
        C[544]), .S(S[544]), .CO(C[545]) );
  FA_16159 \FA_INST_0[1].FA_INST_1[33].FA_  ( .A(A[545]), .B(B[545]), .CI(
        C[545]), .S(S[545]), .CO(C[546]) );
  FA_16158 \FA_INST_0[1].FA_INST_1[34].FA_  ( .A(A[546]), .B(B[546]), .CI(
        C[546]), .S(S[546]), .CO(C[547]) );
  FA_16157 \FA_INST_0[1].FA_INST_1[35].FA_  ( .A(A[547]), .B(B[547]), .CI(
        C[547]), .S(S[547]), .CO(C[548]) );
  FA_16156 \FA_INST_0[1].FA_INST_1[36].FA_  ( .A(A[548]), .B(B[548]), .CI(
        C[548]), .S(S[548]), .CO(C[549]) );
  FA_16155 \FA_INST_0[1].FA_INST_1[37].FA_  ( .A(A[549]), .B(B[549]), .CI(
        C[549]), .S(S[549]), .CO(C[550]) );
  FA_16154 \FA_INST_0[1].FA_INST_1[38].FA_  ( .A(A[550]), .B(B[550]), .CI(
        C[550]), .S(S[550]), .CO(C[551]) );
  FA_16153 \FA_INST_0[1].FA_INST_1[39].FA_  ( .A(A[551]), .B(B[551]), .CI(
        C[551]), .S(S[551]), .CO(C[552]) );
  FA_16152 \FA_INST_0[1].FA_INST_1[40].FA_  ( .A(A[552]), .B(B[552]), .CI(
        C[552]), .S(S[552]), .CO(C[553]) );
  FA_16151 \FA_INST_0[1].FA_INST_1[41].FA_  ( .A(A[553]), .B(B[553]), .CI(
        C[553]), .S(S[553]), .CO(C[554]) );
  FA_16150 \FA_INST_0[1].FA_INST_1[42].FA_  ( .A(A[554]), .B(B[554]), .CI(
        C[554]), .S(S[554]), .CO(C[555]) );
  FA_16149 \FA_INST_0[1].FA_INST_1[43].FA_  ( .A(A[555]), .B(B[555]), .CI(
        C[555]), .S(S[555]), .CO(C[556]) );
  FA_16148 \FA_INST_0[1].FA_INST_1[44].FA_  ( .A(A[556]), .B(B[556]), .CI(
        C[556]), .S(S[556]), .CO(C[557]) );
  FA_16147 \FA_INST_0[1].FA_INST_1[45].FA_  ( .A(A[557]), .B(B[557]), .CI(
        C[557]), .S(S[557]), .CO(C[558]) );
  FA_16146 \FA_INST_0[1].FA_INST_1[46].FA_  ( .A(A[558]), .B(B[558]), .CI(
        C[558]), .S(S[558]), .CO(C[559]) );
  FA_16145 \FA_INST_0[1].FA_INST_1[47].FA_  ( .A(A[559]), .B(B[559]), .CI(
        C[559]), .S(S[559]), .CO(C[560]) );
  FA_16144 \FA_INST_0[1].FA_INST_1[48].FA_  ( .A(A[560]), .B(B[560]), .CI(
        C[560]), .S(S[560]), .CO(C[561]) );
  FA_16143 \FA_INST_0[1].FA_INST_1[49].FA_  ( .A(A[561]), .B(B[561]), .CI(
        C[561]), .S(S[561]), .CO(C[562]) );
  FA_16142 \FA_INST_0[1].FA_INST_1[50].FA_  ( .A(A[562]), .B(B[562]), .CI(
        C[562]), .S(S[562]), .CO(C[563]) );
  FA_16141 \FA_INST_0[1].FA_INST_1[51].FA_  ( .A(A[563]), .B(B[563]), .CI(
        C[563]), .S(S[563]), .CO(C[564]) );
  FA_16140 \FA_INST_0[1].FA_INST_1[52].FA_  ( .A(A[564]), .B(B[564]), .CI(
        C[564]), .S(S[564]), .CO(C[565]) );
  FA_16139 \FA_INST_0[1].FA_INST_1[53].FA_  ( .A(A[565]), .B(B[565]), .CI(
        C[565]), .S(S[565]), .CO(C[566]) );
  FA_16138 \FA_INST_0[1].FA_INST_1[54].FA_  ( .A(A[566]), .B(B[566]), .CI(
        C[566]), .S(S[566]), .CO(C[567]) );
  FA_16137 \FA_INST_0[1].FA_INST_1[55].FA_  ( .A(A[567]), .B(B[567]), .CI(
        C[567]), .S(S[567]), .CO(C[568]) );
  FA_16136 \FA_INST_0[1].FA_INST_1[56].FA_  ( .A(A[568]), .B(B[568]), .CI(
        C[568]), .S(S[568]), .CO(C[569]) );
  FA_16135 \FA_INST_0[1].FA_INST_1[57].FA_  ( .A(A[569]), .B(B[569]), .CI(
        C[569]), .S(S[569]), .CO(C[570]) );
  FA_16134 \FA_INST_0[1].FA_INST_1[58].FA_  ( .A(A[570]), .B(B[570]), .CI(
        C[570]), .S(S[570]), .CO(C[571]) );
  FA_16133 \FA_INST_0[1].FA_INST_1[59].FA_  ( .A(A[571]), .B(B[571]), .CI(
        C[571]), .S(S[571]), .CO(C[572]) );
  FA_16132 \FA_INST_0[1].FA_INST_1[60].FA_  ( .A(A[572]), .B(B[572]), .CI(
        C[572]), .S(S[572]), .CO(C[573]) );
  FA_16131 \FA_INST_0[1].FA_INST_1[61].FA_  ( .A(A[573]), .B(B[573]), .CI(
        C[573]), .S(S[573]), .CO(C[574]) );
  FA_16130 \FA_INST_0[1].FA_INST_1[62].FA_  ( .A(A[574]), .B(B[574]), .CI(
        C[574]), .S(S[574]), .CO(C[575]) );
  FA_16129 \FA_INST_0[1].FA_INST_1[63].FA_  ( .A(A[575]), .B(B[575]), .CI(
        C[575]), .S(S[575]), .CO(C[576]) );
  FA_16128 \FA_INST_0[1].FA_INST_1[64].FA_  ( .A(A[576]), .B(B[576]), .CI(
        C[576]), .S(S[576]), .CO(C[577]) );
  FA_16127 \FA_INST_0[1].FA_INST_1[65].FA_  ( .A(A[577]), .B(B[577]), .CI(
        C[577]), .S(S[577]), .CO(C[578]) );
  FA_16126 \FA_INST_0[1].FA_INST_1[66].FA_  ( .A(A[578]), .B(B[578]), .CI(
        C[578]), .S(S[578]), .CO(C[579]) );
  FA_16125 \FA_INST_0[1].FA_INST_1[67].FA_  ( .A(A[579]), .B(B[579]), .CI(
        C[579]), .S(S[579]), .CO(C[580]) );
  FA_16124 \FA_INST_0[1].FA_INST_1[68].FA_  ( .A(A[580]), .B(B[580]), .CI(
        C[580]), .S(S[580]), .CO(C[581]) );
  FA_16123 \FA_INST_0[1].FA_INST_1[69].FA_  ( .A(A[581]), .B(B[581]), .CI(
        C[581]), .S(S[581]), .CO(C[582]) );
  FA_16122 \FA_INST_0[1].FA_INST_1[70].FA_  ( .A(A[582]), .B(B[582]), .CI(
        C[582]), .S(S[582]), .CO(C[583]) );
  FA_16121 \FA_INST_0[1].FA_INST_1[71].FA_  ( .A(A[583]), .B(B[583]), .CI(
        C[583]), .S(S[583]), .CO(C[584]) );
  FA_16120 \FA_INST_0[1].FA_INST_1[72].FA_  ( .A(A[584]), .B(B[584]), .CI(
        C[584]), .S(S[584]), .CO(C[585]) );
  FA_16119 \FA_INST_0[1].FA_INST_1[73].FA_  ( .A(A[585]), .B(B[585]), .CI(
        C[585]), .S(S[585]), .CO(C[586]) );
  FA_16118 \FA_INST_0[1].FA_INST_1[74].FA_  ( .A(A[586]), .B(B[586]), .CI(
        C[586]), .S(S[586]), .CO(C[587]) );
  FA_16117 \FA_INST_0[1].FA_INST_1[75].FA_  ( .A(A[587]), .B(B[587]), .CI(
        C[587]), .S(S[587]), .CO(C[588]) );
  FA_16116 \FA_INST_0[1].FA_INST_1[76].FA_  ( .A(A[588]), .B(B[588]), .CI(
        C[588]), .S(S[588]), .CO(C[589]) );
  FA_16115 \FA_INST_0[1].FA_INST_1[77].FA_  ( .A(A[589]), .B(B[589]), .CI(
        C[589]), .S(S[589]), .CO(C[590]) );
  FA_16114 \FA_INST_0[1].FA_INST_1[78].FA_  ( .A(A[590]), .B(B[590]), .CI(
        C[590]), .S(S[590]), .CO(C[591]) );
  FA_16113 \FA_INST_0[1].FA_INST_1[79].FA_  ( .A(A[591]), .B(B[591]), .CI(
        C[591]), .S(S[591]), .CO(C[592]) );
  FA_16112 \FA_INST_0[1].FA_INST_1[80].FA_  ( .A(A[592]), .B(B[592]), .CI(
        C[592]), .S(S[592]), .CO(C[593]) );
  FA_16111 \FA_INST_0[1].FA_INST_1[81].FA_  ( .A(A[593]), .B(B[593]), .CI(
        C[593]), .S(S[593]), .CO(C[594]) );
  FA_16110 \FA_INST_0[1].FA_INST_1[82].FA_  ( .A(A[594]), .B(B[594]), .CI(
        C[594]), .S(S[594]), .CO(C[595]) );
  FA_16109 \FA_INST_0[1].FA_INST_1[83].FA_  ( .A(A[595]), .B(B[595]), .CI(
        C[595]), .S(S[595]), .CO(C[596]) );
  FA_16108 \FA_INST_0[1].FA_INST_1[84].FA_  ( .A(A[596]), .B(B[596]), .CI(
        C[596]), .S(S[596]), .CO(C[597]) );
  FA_16107 \FA_INST_0[1].FA_INST_1[85].FA_  ( .A(A[597]), .B(B[597]), .CI(
        C[597]), .S(S[597]), .CO(C[598]) );
  FA_16106 \FA_INST_0[1].FA_INST_1[86].FA_  ( .A(A[598]), .B(B[598]), .CI(
        C[598]), .S(S[598]), .CO(C[599]) );
  FA_16105 \FA_INST_0[1].FA_INST_1[87].FA_  ( .A(A[599]), .B(B[599]), .CI(
        C[599]), .S(S[599]), .CO(C[600]) );
  FA_16104 \FA_INST_0[1].FA_INST_1[88].FA_  ( .A(A[600]), .B(B[600]), .CI(
        C[600]), .S(S[600]), .CO(C[601]) );
  FA_16103 \FA_INST_0[1].FA_INST_1[89].FA_  ( .A(A[601]), .B(B[601]), .CI(
        C[601]), .S(S[601]), .CO(C[602]) );
  FA_16102 \FA_INST_0[1].FA_INST_1[90].FA_  ( .A(A[602]), .B(B[602]), .CI(
        C[602]), .S(S[602]), .CO(C[603]) );
  FA_16101 \FA_INST_0[1].FA_INST_1[91].FA_  ( .A(A[603]), .B(B[603]), .CI(
        C[603]), .S(S[603]), .CO(C[604]) );
  FA_16100 \FA_INST_0[1].FA_INST_1[92].FA_  ( .A(A[604]), .B(B[604]), .CI(
        C[604]), .S(S[604]), .CO(C[605]) );
  FA_16099 \FA_INST_0[1].FA_INST_1[93].FA_  ( .A(A[605]), .B(B[605]), .CI(
        C[605]), .S(S[605]), .CO(C[606]) );
  FA_16098 \FA_INST_0[1].FA_INST_1[94].FA_  ( .A(A[606]), .B(B[606]), .CI(
        C[606]), .S(S[606]), .CO(C[607]) );
  FA_16097 \FA_INST_0[1].FA_INST_1[95].FA_  ( .A(A[607]), .B(B[607]), .CI(
        C[607]), .S(S[607]), .CO(C[608]) );
  FA_16096 \FA_INST_0[1].FA_INST_1[96].FA_  ( .A(A[608]), .B(B[608]), .CI(
        C[608]), .S(S[608]), .CO(C[609]) );
  FA_16095 \FA_INST_0[1].FA_INST_1[97].FA_  ( .A(A[609]), .B(B[609]), .CI(
        C[609]), .S(S[609]), .CO(C[610]) );
  FA_16094 \FA_INST_0[1].FA_INST_1[98].FA_  ( .A(A[610]), .B(B[610]), .CI(
        C[610]), .S(S[610]), .CO(C[611]) );
  FA_16093 \FA_INST_0[1].FA_INST_1[99].FA_  ( .A(A[611]), .B(B[611]), .CI(
        C[611]), .S(S[611]), .CO(C[612]) );
  FA_16092 \FA_INST_0[1].FA_INST_1[100].FA_  ( .A(A[612]), .B(B[612]), .CI(
        C[612]), .S(S[612]), .CO(C[613]) );
  FA_16091 \FA_INST_0[1].FA_INST_1[101].FA_  ( .A(A[613]), .B(B[613]), .CI(
        C[613]), .S(S[613]), .CO(C[614]) );
  FA_16090 \FA_INST_0[1].FA_INST_1[102].FA_  ( .A(A[614]), .B(B[614]), .CI(
        C[614]), .S(S[614]), .CO(C[615]) );
  FA_16089 \FA_INST_0[1].FA_INST_1[103].FA_  ( .A(A[615]), .B(B[615]), .CI(
        C[615]), .S(S[615]), .CO(C[616]) );
  FA_16088 \FA_INST_0[1].FA_INST_1[104].FA_  ( .A(A[616]), .B(B[616]), .CI(
        C[616]), .S(S[616]), .CO(C[617]) );
  FA_16087 \FA_INST_0[1].FA_INST_1[105].FA_  ( .A(A[617]), .B(B[617]), .CI(
        C[617]), .S(S[617]), .CO(C[618]) );
  FA_16086 \FA_INST_0[1].FA_INST_1[106].FA_  ( .A(A[618]), .B(B[618]), .CI(
        C[618]), .S(S[618]), .CO(C[619]) );
  FA_16085 \FA_INST_0[1].FA_INST_1[107].FA_  ( .A(A[619]), .B(B[619]), .CI(
        C[619]), .S(S[619]), .CO(C[620]) );
  FA_16084 \FA_INST_0[1].FA_INST_1[108].FA_  ( .A(A[620]), .B(B[620]), .CI(
        C[620]), .S(S[620]), .CO(C[621]) );
  FA_16083 \FA_INST_0[1].FA_INST_1[109].FA_  ( .A(A[621]), .B(B[621]), .CI(
        C[621]), .S(S[621]), .CO(C[622]) );
  FA_16082 \FA_INST_0[1].FA_INST_1[110].FA_  ( .A(A[622]), .B(B[622]), .CI(
        C[622]), .S(S[622]), .CO(C[623]) );
  FA_16081 \FA_INST_0[1].FA_INST_1[111].FA_  ( .A(A[623]), .B(B[623]), .CI(
        C[623]), .S(S[623]), .CO(C[624]) );
  FA_16080 \FA_INST_0[1].FA_INST_1[112].FA_  ( .A(A[624]), .B(B[624]), .CI(
        C[624]), .S(S[624]), .CO(C[625]) );
  FA_16079 \FA_INST_0[1].FA_INST_1[113].FA_  ( .A(A[625]), .B(B[625]), .CI(
        C[625]), .S(S[625]), .CO(C[626]) );
  FA_16078 \FA_INST_0[1].FA_INST_1[114].FA_  ( .A(A[626]), .B(B[626]), .CI(
        C[626]), .S(S[626]), .CO(C[627]) );
  FA_16077 \FA_INST_0[1].FA_INST_1[115].FA_  ( .A(A[627]), .B(B[627]), .CI(
        C[627]), .S(S[627]), .CO(C[628]) );
  FA_16076 \FA_INST_0[1].FA_INST_1[116].FA_  ( .A(A[628]), .B(B[628]), .CI(
        C[628]), .S(S[628]), .CO(C[629]) );
  FA_16075 \FA_INST_0[1].FA_INST_1[117].FA_  ( .A(A[629]), .B(B[629]), .CI(
        C[629]), .S(S[629]), .CO(C[630]) );
  FA_16074 \FA_INST_0[1].FA_INST_1[118].FA_  ( .A(A[630]), .B(B[630]), .CI(
        C[630]), .S(S[630]), .CO(C[631]) );
  FA_16073 \FA_INST_0[1].FA_INST_1[119].FA_  ( .A(A[631]), .B(B[631]), .CI(
        C[631]), .S(S[631]), .CO(C[632]) );
  FA_16072 \FA_INST_0[1].FA_INST_1[120].FA_  ( .A(A[632]), .B(B[632]), .CI(
        C[632]), .S(S[632]), .CO(C[633]) );
  FA_16071 \FA_INST_0[1].FA_INST_1[121].FA_  ( .A(A[633]), .B(B[633]), .CI(
        C[633]), .S(S[633]), .CO(C[634]) );
  FA_16070 \FA_INST_0[1].FA_INST_1[122].FA_  ( .A(A[634]), .B(B[634]), .CI(
        C[634]), .S(S[634]), .CO(C[635]) );
  FA_16069 \FA_INST_0[1].FA_INST_1[123].FA_  ( .A(A[635]), .B(B[635]), .CI(
        C[635]), .S(S[635]), .CO(C[636]) );
  FA_16068 \FA_INST_0[1].FA_INST_1[124].FA_  ( .A(A[636]), .B(B[636]), .CI(
        C[636]), .S(S[636]), .CO(C[637]) );
  FA_16067 \FA_INST_0[1].FA_INST_1[125].FA_  ( .A(A[637]), .B(B[637]), .CI(
        C[637]), .S(S[637]), .CO(C[638]) );
  FA_16066 \FA_INST_0[1].FA_INST_1[126].FA_  ( .A(A[638]), .B(B[638]), .CI(
        C[638]), .S(S[638]), .CO(C[639]) );
  FA_16065 \FA_INST_0[1].FA_INST_1[127].FA_  ( .A(A[639]), .B(B[639]), .CI(
        C[639]), .S(S[639]), .CO(C[640]) );
  FA_16064 \FA_INST_0[1].FA_INST_1[128].FA_  ( .A(A[640]), .B(B[640]), .CI(
        C[640]), .S(S[640]), .CO(C[641]) );
  FA_16063 \FA_INST_0[1].FA_INST_1[129].FA_  ( .A(A[641]), .B(B[641]), .CI(
        C[641]), .S(S[641]), .CO(C[642]) );
  FA_16062 \FA_INST_0[1].FA_INST_1[130].FA_  ( .A(A[642]), .B(B[642]), .CI(
        C[642]), .S(S[642]), .CO(C[643]) );
  FA_16061 \FA_INST_0[1].FA_INST_1[131].FA_  ( .A(A[643]), .B(B[643]), .CI(
        C[643]), .S(S[643]), .CO(C[644]) );
  FA_16060 \FA_INST_0[1].FA_INST_1[132].FA_  ( .A(A[644]), .B(B[644]), .CI(
        C[644]), .S(S[644]), .CO(C[645]) );
  FA_16059 \FA_INST_0[1].FA_INST_1[133].FA_  ( .A(A[645]), .B(B[645]), .CI(
        C[645]), .S(S[645]), .CO(C[646]) );
  FA_16058 \FA_INST_0[1].FA_INST_1[134].FA_  ( .A(A[646]), .B(B[646]), .CI(
        C[646]), .S(S[646]), .CO(C[647]) );
  FA_16057 \FA_INST_0[1].FA_INST_1[135].FA_  ( .A(A[647]), .B(B[647]), .CI(
        C[647]), .S(S[647]), .CO(C[648]) );
  FA_16056 \FA_INST_0[1].FA_INST_1[136].FA_  ( .A(A[648]), .B(B[648]), .CI(
        C[648]), .S(S[648]), .CO(C[649]) );
  FA_16055 \FA_INST_0[1].FA_INST_1[137].FA_  ( .A(A[649]), .B(B[649]), .CI(
        C[649]), .S(S[649]), .CO(C[650]) );
  FA_16054 \FA_INST_0[1].FA_INST_1[138].FA_  ( .A(A[650]), .B(B[650]), .CI(
        C[650]), .S(S[650]), .CO(C[651]) );
  FA_16053 \FA_INST_0[1].FA_INST_1[139].FA_  ( .A(A[651]), .B(B[651]), .CI(
        C[651]), .S(S[651]), .CO(C[652]) );
  FA_16052 \FA_INST_0[1].FA_INST_1[140].FA_  ( .A(A[652]), .B(B[652]), .CI(
        C[652]), .S(S[652]), .CO(C[653]) );
  FA_16051 \FA_INST_0[1].FA_INST_1[141].FA_  ( .A(A[653]), .B(B[653]), .CI(
        C[653]), .S(S[653]), .CO(C[654]) );
  FA_16050 \FA_INST_0[1].FA_INST_1[142].FA_  ( .A(A[654]), .B(B[654]), .CI(
        C[654]), .S(S[654]), .CO(C[655]) );
  FA_16049 \FA_INST_0[1].FA_INST_1[143].FA_  ( .A(A[655]), .B(B[655]), .CI(
        C[655]), .S(S[655]), .CO(C[656]) );
  FA_16048 \FA_INST_0[1].FA_INST_1[144].FA_  ( .A(A[656]), .B(B[656]), .CI(
        C[656]), .S(S[656]), .CO(C[657]) );
  FA_16047 \FA_INST_0[1].FA_INST_1[145].FA_  ( .A(A[657]), .B(B[657]), .CI(
        C[657]), .S(S[657]), .CO(C[658]) );
  FA_16046 \FA_INST_0[1].FA_INST_1[146].FA_  ( .A(A[658]), .B(B[658]), .CI(
        C[658]), .S(S[658]), .CO(C[659]) );
  FA_16045 \FA_INST_0[1].FA_INST_1[147].FA_  ( .A(A[659]), .B(B[659]), .CI(
        C[659]), .S(S[659]), .CO(C[660]) );
  FA_16044 \FA_INST_0[1].FA_INST_1[148].FA_  ( .A(A[660]), .B(B[660]), .CI(
        C[660]), .S(S[660]), .CO(C[661]) );
  FA_16043 \FA_INST_0[1].FA_INST_1[149].FA_  ( .A(A[661]), .B(B[661]), .CI(
        C[661]), .S(S[661]), .CO(C[662]) );
  FA_16042 \FA_INST_0[1].FA_INST_1[150].FA_  ( .A(A[662]), .B(B[662]), .CI(
        C[662]), .S(S[662]), .CO(C[663]) );
  FA_16041 \FA_INST_0[1].FA_INST_1[151].FA_  ( .A(A[663]), .B(B[663]), .CI(
        C[663]), .S(S[663]), .CO(C[664]) );
  FA_16040 \FA_INST_0[1].FA_INST_1[152].FA_  ( .A(A[664]), .B(B[664]), .CI(
        C[664]), .S(S[664]), .CO(C[665]) );
  FA_16039 \FA_INST_0[1].FA_INST_1[153].FA_  ( .A(A[665]), .B(B[665]), .CI(
        C[665]), .S(S[665]), .CO(C[666]) );
  FA_16038 \FA_INST_0[1].FA_INST_1[154].FA_  ( .A(A[666]), .B(B[666]), .CI(
        C[666]), .S(S[666]), .CO(C[667]) );
  FA_16037 \FA_INST_0[1].FA_INST_1[155].FA_  ( .A(A[667]), .B(B[667]), .CI(
        C[667]), .S(S[667]), .CO(C[668]) );
  FA_16036 \FA_INST_0[1].FA_INST_1[156].FA_  ( .A(A[668]), .B(B[668]), .CI(
        C[668]), .S(S[668]), .CO(C[669]) );
  FA_16035 \FA_INST_0[1].FA_INST_1[157].FA_  ( .A(A[669]), .B(B[669]), .CI(
        C[669]), .S(S[669]), .CO(C[670]) );
  FA_16034 \FA_INST_0[1].FA_INST_1[158].FA_  ( .A(A[670]), .B(B[670]), .CI(
        C[670]), .S(S[670]), .CO(C[671]) );
  FA_16033 \FA_INST_0[1].FA_INST_1[159].FA_  ( .A(A[671]), .B(B[671]), .CI(
        C[671]), .S(S[671]), .CO(C[672]) );
  FA_16032 \FA_INST_0[1].FA_INST_1[160].FA_  ( .A(A[672]), .B(B[672]), .CI(
        C[672]), .S(S[672]), .CO(C[673]) );
  FA_16031 \FA_INST_0[1].FA_INST_1[161].FA_  ( .A(A[673]), .B(B[673]), .CI(
        C[673]), .S(S[673]), .CO(C[674]) );
  FA_16030 \FA_INST_0[1].FA_INST_1[162].FA_  ( .A(A[674]), .B(B[674]), .CI(
        C[674]), .S(S[674]), .CO(C[675]) );
  FA_16029 \FA_INST_0[1].FA_INST_1[163].FA_  ( .A(A[675]), .B(B[675]), .CI(
        C[675]), .S(S[675]), .CO(C[676]) );
  FA_16028 \FA_INST_0[1].FA_INST_1[164].FA_  ( .A(A[676]), .B(B[676]), .CI(
        C[676]), .S(S[676]), .CO(C[677]) );
  FA_16027 \FA_INST_0[1].FA_INST_1[165].FA_  ( .A(A[677]), .B(B[677]), .CI(
        C[677]), .S(S[677]), .CO(C[678]) );
  FA_16026 \FA_INST_0[1].FA_INST_1[166].FA_  ( .A(A[678]), .B(B[678]), .CI(
        C[678]), .S(S[678]), .CO(C[679]) );
  FA_16025 \FA_INST_0[1].FA_INST_1[167].FA_  ( .A(A[679]), .B(B[679]), .CI(
        C[679]), .S(S[679]), .CO(C[680]) );
  FA_16024 \FA_INST_0[1].FA_INST_1[168].FA_  ( .A(A[680]), .B(B[680]), .CI(
        C[680]), .S(S[680]), .CO(C[681]) );
  FA_16023 \FA_INST_0[1].FA_INST_1[169].FA_  ( .A(A[681]), .B(B[681]), .CI(
        C[681]), .S(S[681]), .CO(C[682]) );
  FA_16022 \FA_INST_0[1].FA_INST_1[170].FA_  ( .A(A[682]), .B(B[682]), .CI(
        C[682]), .S(S[682]), .CO(C[683]) );
  FA_16021 \FA_INST_0[1].FA_INST_1[171].FA_  ( .A(A[683]), .B(B[683]), .CI(
        C[683]), .S(S[683]), .CO(C[684]) );
  FA_16020 \FA_INST_0[1].FA_INST_1[172].FA_  ( .A(A[684]), .B(B[684]), .CI(
        C[684]), .S(S[684]), .CO(C[685]) );
  FA_16019 \FA_INST_0[1].FA_INST_1[173].FA_  ( .A(A[685]), .B(B[685]), .CI(
        C[685]), .S(S[685]), .CO(C[686]) );
  FA_16018 \FA_INST_0[1].FA_INST_1[174].FA_  ( .A(A[686]), .B(B[686]), .CI(
        C[686]), .S(S[686]), .CO(C[687]) );
  FA_16017 \FA_INST_0[1].FA_INST_1[175].FA_  ( .A(A[687]), .B(B[687]), .CI(
        C[687]), .S(S[687]), .CO(C[688]) );
  FA_16016 \FA_INST_0[1].FA_INST_1[176].FA_  ( .A(A[688]), .B(B[688]), .CI(
        C[688]), .S(S[688]), .CO(C[689]) );
  FA_16015 \FA_INST_0[1].FA_INST_1[177].FA_  ( .A(A[689]), .B(B[689]), .CI(
        C[689]), .S(S[689]), .CO(C[690]) );
  FA_16014 \FA_INST_0[1].FA_INST_1[178].FA_  ( .A(A[690]), .B(B[690]), .CI(
        C[690]), .S(S[690]), .CO(C[691]) );
  FA_16013 \FA_INST_0[1].FA_INST_1[179].FA_  ( .A(A[691]), .B(B[691]), .CI(
        C[691]), .S(S[691]), .CO(C[692]) );
  FA_16012 \FA_INST_0[1].FA_INST_1[180].FA_  ( .A(A[692]), .B(B[692]), .CI(
        C[692]), .S(S[692]), .CO(C[693]) );
  FA_16011 \FA_INST_0[1].FA_INST_1[181].FA_  ( .A(A[693]), .B(B[693]), .CI(
        C[693]), .S(S[693]), .CO(C[694]) );
  FA_16010 \FA_INST_0[1].FA_INST_1[182].FA_  ( .A(A[694]), .B(B[694]), .CI(
        C[694]), .S(S[694]), .CO(C[695]) );
  FA_16009 \FA_INST_0[1].FA_INST_1[183].FA_  ( .A(A[695]), .B(B[695]), .CI(
        C[695]), .S(S[695]), .CO(C[696]) );
  FA_16008 \FA_INST_0[1].FA_INST_1[184].FA_  ( .A(A[696]), .B(B[696]), .CI(
        C[696]), .S(S[696]), .CO(C[697]) );
  FA_16007 \FA_INST_0[1].FA_INST_1[185].FA_  ( .A(A[697]), .B(B[697]), .CI(
        C[697]), .S(S[697]), .CO(C[698]) );
  FA_16006 \FA_INST_0[1].FA_INST_1[186].FA_  ( .A(A[698]), .B(B[698]), .CI(
        C[698]), .S(S[698]), .CO(C[699]) );
  FA_16005 \FA_INST_0[1].FA_INST_1[187].FA_  ( .A(A[699]), .B(B[699]), .CI(
        C[699]), .S(S[699]), .CO(C[700]) );
  FA_16004 \FA_INST_0[1].FA_INST_1[188].FA_  ( .A(A[700]), .B(B[700]), .CI(
        C[700]), .S(S[700]), .CO(C[701]) );
  FA_16003 \FA_INST_0[1].FA_INST_1[189].FA_  ( .A(A[701]), .B(B[701]), .CI(
        C[701]), .S(S[701]), .CO(C[702]) );
  FA_16002 \FA_INST_0[1].FA_INST_1[190].FA_  ( .A(A[702]), .B(B[702]), .CI(
        C[702]), .S(S[702]), .CO(C[703]) );
  FA_16001 \FA_INST_0[1].FA_INST_1[191].FA_  ( .A(A[703]), .B(B[703]), .CI(
        C[703]), .S(S[703]), .CO(C[704]) );
  FA_16000 \FA_INST_0[1].FA_INST_1[192].FA_  ( .A(A[704]), .B(B[704]), .CI(
        C[704]), .S(S[704]), .CO(C[705]) );
  FA_15999 \FA_INST_0[1].FA_INST_1[193].FA_  ( .A(A[705]), .B(B[705]), .CI(
        C[705]), .S(S[705]), .CO(C[706]) );
  FA_15998 \FA_INST_0[1].FA_INST_1[194].FA_  ( .A(A[706]), .B(B[706]), .CI(
        C[706]), .S(S[706]), .CO(C[707]) );
  FA_15997 \FA_INST_0[1].FA_INST_1[195].FA_  ( .A(A[707]), .B(B[707]), .CI(
        C[707]), .S(S[707]), .CO(C[708]) );
  FA_15996 \FA_INST_0[1].FA_INST_1[196].FA_  ( .A(A[708]), .B(B[708]), .CI(
        C[708]), .S(S[708]), .CO(C[709]) );
  FA_15995 \FA_INST_0[1].FA_INST_1[197].FA_  ( .A(A[709]), .B(B[709]), .CI(
        C[709]), .S(S[709]), .CO(C[710]) );
  FA_15994 \FA_INST_0[1].FA_INST_1[198].FA_  ( .A(A[710]), .B(B[710]), .CI(
        C[710]), .S(S[710]), .CO(C[711]) );
  FA_15993 \FA_INST_0[1].FA_INST_1[199].FA_  ( .A(A[711]), .B(B[711]), .CI(
        C[711]), .S(S[711]), .CO(C[712]) );
  FA_15992 \FA_INST_0[1].FA_INST_1[200].FA_  ( .A(A[712]), .B(B[712]), .CI(
        C[712]), .S(S[712]), .CO(C[713]) );
  FA_15991 \FA_INST_0[1].FA_INST_1[201].FA_  ( .A(A[713]), .B(B[713]), .CI(
        C[713]), .S(S[713]), .CO(C[714]) );
  FA_15990 \FA_INST_0[1].FA_INST_1[202].FA_  ( .A(A[714]), .B(B[714]), .CI(
        C[714]), .S(S[714]), .CO(C[715]) );
  FA_15989 \FA_INST_0[1].FA_INST_1[203].FA_  ( .A(A[715]), .B(B[715]), .CI(
        C[715]), .S(S[715]), .CO(C[716]) );
  FA_15988 \FA_INST_0[1].FA_INST_1[204].FA_  ( .A(A[716]), .B(B[716]), .CI(
        C[716]), .S(S[716]), .CO(C[717]) );
  FA_15987 \FA_INST_0[1].FA_INST_1[205].FA_  ( .A(A[717]), .B(B[717]), .CI(
        C[717]), .S(S[717]), .CO(C[718]) );
  FA_15986 \FA_INST_0[1].FA_INST_1[206].FA_  ( .A(A[718]), .B(B[718]), .CI(
        C[718]), .S(S[718]), .CO(C[719]) );
  FA_15985 \FA_INST_0[1].FA_INST_1[207].FA_  ( .A(A[719]), .B(B[719]), .CI(
        C[719]), .S(S[719]), .CO(C[720]) );
  FA_15984 \FA_INST_0[1].FA_INST_1[208].FA_  ( .A(A[720]), .B(B[720]), .CI(
        C[720]), .S(S[720]), .CO(C[721]) );
  FA_15983 \FA_INST_0[1].FA_INST_1[209].FA_  ( .A(A[721]), .B(B[721]), .CI(
        C[721]), .S(S[721]), .CO(C[722]) );
  FA_15982 \FA_INST_0[1].FA_INST_1[210].FA_  ( .A(A[722]), .B(B[722]), .CI(
        C[722]), .S(S[722]), .CO(C[723]) );
  FA_15981 \FA_INST_0[1].FA_INST_1[211].FA_  ( .A(A[723]), .B(B[723]), .CI(
        C[723]), .S(S[723]), .CO(C[724]) );
  FA_15980 \FA_INST_0[1].FA_INST_1[212].FA_  ( .A(A[724]), .B(B[724]), .CI(
        C[724]), .S(S[724]), .CO(C[725]) );
  FA_15979 \FA_INST_0[1].FA_INST_1[213].FA_  ( .A(A[725]), .B(B[725]), .CI(
        C[725]), .S(S[725]), .CO(C[726]) );
  FA_15978 \FA_INST_0[1].FA_INST_1[214].FA_  ( .A(A[726]), .B(B[726]), .CI(
        C[726]), .S(S[726]), .CO(C[727]) );
  FA_15977 \FA_INST_0[1].FA_INST_1[215].FA_  ( .A(A[727]), .B(B[727]), .CI(
        C[727]), .S(S[727]), .CO(C[728]) );
  FA_15976 \FA_INST_0[1].FA_INST_1[216].FA_  ( .A(A[728]), .B(B[728]), .CI(
        C[728]), .S(S[728]), .CO(C[729]) );
  FA_15975 \FA_INST_0[1].FA_INST_1[217].FA_  ( .A(A[729]), .B(B[729]), .CI(
        C[729]), .S(S[729]), .CO(C[730]) );
  FA_15974 \FA_INST_0[1].FA_INST_1[218].FA_  ( .A(A[730]), .B(B[730]), .CI(
        C[730]), .S(S[730]), .CO(C[731]) );
  FA_15973 \FA_INST_0[1].FA_INST_1[219].FA_  ( .A(A[731]), .B(B[731]), .CI(
        C[731]), .S(S[731]), .CO(C[732]) );
  FA_15972 \FA_INST_0[1].FA_INST_1[220].FA_  ( .A(A[732]), .B(B[732]), .CI(
        C[732]), .S(S[732]), .CO(C[733]) );
  FA_15971 \FA_INST_0[1].FA_INST_1[221].FA_  ( .A(A[733]), .B(B[733]), .CI(
        C[733]), .S(S[733]), .CO(C[734]) );
  FA_15970 \FA_INST_0[1].FA_INST_1[222].FA_  ( .A(A[734]), .B(B[734]), .CI(
        C[734]), .S(S[734]), .CO(C[735]) );
  FA_15969 \FA_INST_0[1].FA_INST_1[223].FA_  ( .A(A[735]), .B(B[735]), .CI(
        C[735]), .S(S[735]), .CO(C[736]) );
  FA_15968 \FA_INST_0[1].FA_INST_1[224].FA_  ( .A(A[736]), .B(B[736]), .CI(
        C[736]), .S(S[736]), .CO(C[737]) );
  FA_15967 \FA_INST_0[1].FA_INST_1[225].FA_  ( .A(A[737]), .B(B[737]), .CI(
        C[737]), .S(S[737]), .CO(C[738]) );
  FA_15966 \FA_INST_0[1].FA_INST_1[226].FA_  ( .A(A[738]), .B(B[738]), .CI(
        C[738]), .S(S[738]), .CO(C[739]) );
  FA_15965 \FA_INST_0[1].FA_INST_1[227].FA_  ( .A(A[739]), .B(B[739]), .CI(
        C[739]), .S(S[739]), .CO(C[740]) );
  FA_15964 \FA_INST_0[1].FA_INST_1[228].FA_  ( .A(A[740]), .B(B[740]), .CI(
        C[740]), .S(S[740]), .CO(C[741]) );
  FA_15963 \FA_INST_0[1].FA_INST_1[229].FA_  ( .A(A[741]), .B(B[741]), .CI(
        C[741]), .S(S[741]), .CO(C[742]) );
  FA_15962 \FA_INST_0[1].FA_INST_1[230].FA_  ( .A(A[742]), .B(B[742]), .CI(
        C[742]), .S(S[742]), .CO(C[743]) );
  FA_15961 \FA_INST_0[1].FA_INST_1[231].FA_  ( .A(A[743]), .B(B[743]), .CI(
        C[743]), .S(S[743]), .CO(C[744]) );
  FA_15960 \FA_INST_0[1].FA_INST_1[232].FA_  ( .A(A[744]), .B(B[744]), .CI(
        C[744]), .S(S[744]), .CO(C[745]) );
  FA_15959 \FA_INST_0[1].FA_INST_1[233].FA_  ( .A(A[745]), .B(B[745]), .CI(
        C[745]), .S(S[745]), .CO(C[746]) );
  FA_15958 \FA_INST_0[1].FA_INST_1[234].FA_  ( .A(A[746]), .B(B[746]), .CI(
        C[746]), .S(S[746]), .CO(C[747]) );
  FA_15957 \FA_INST_0[1].FA_INST_1[235].FA_  ( .A(A[747]), .B(B[747]), .CI(
        C[747]), .S(S[747]), .CO(C[748]) );
  FA_15956 \FA_INST_0[1].FA_INST_1[236].FA_  ( .A(A[748]), .B(B[748]), .CI(
        C[748]), .S(S[748]), .CO(C[749]) );
  FA_15955 \FA_INST_0[1].FA_INST_1[237].FA_  ( .A(A[749]), .B(B[749]), .CI(
        C[749]), .S(S[749]), .CO(C[750]) );
  FA_15954 \FA_INST_0[1].FA_INST_1[238].FA_  ( .A(A[750]), .B(B[750]), .CI(
        C[750]), .S(S[750]), .CO(C[751]) );
  FA_15953 \FA_INST_0[1].FA_INST_1[239].FA_  ( .A(A[751]), .B(B[751]), .CI(
        C[751]), .S(S[751]), .CO(C[752]) );
  FA_15952 \FA_INST_0[1].FA_INST_1[240].FA_  ( .A(A[752]), .B(B[752]), .CI(
        C[752]), .S(S[752]), .CO(C[753]) );
  FA_15951 \FA_INST_0[1].FA_INST_1[241].FA_  ( .A(A[753]), .B(B[753]), .CI(
        C[753]), .S(S[753]), .CO(C[754]) );
  FA_15950 \FA_INST_0[1].FA_INST_1[242].FA_  ( .A(A[754]), .B(B[754]), .CI(
        C[754]), .S(S[754]), .CO(C[755]) );
  FA_15949 \FA_INST_0[1].FA_INST_1[243].FA_  ( .A(A[755]), .B(B[755]), .CI(
        C[755]), .S(S[755]), .CO(C[756]) );
  FA_15948 \FA_INST_0[1].FA_INST_1[244].FA_  ( .A(A[756]), .B(B[756]), .CI(
        C[756]), .S(S[756]), .CO(C[757]) );
  FA_15947 \FA_INST_0[1].FA_INST_1[245].FA_  ( .A(A[757]), .B(B[757]), .CI(
        C[757]), .S(S[757]), .CO(C[758]) );
  FA_15946 \FA_INST_0[1].FA_INST_1[246].FA_  ( .A(A[758]), .B(B[758]), .CI(
        C[758]), .S(S[758]), .CO(C[759]) );
  FA_15945 \FA_INST_0[1].FA_INST_1[247].FA_  ( .A(A[759]), .B(B[759]), .CI(
        C[759]), .S(S[759]), .CO(C[760]) );
  FA_15944 \FA_INST_0[1].FA_INST_1[248].FA_  ( .A(A[760]), .B(B[760]), .CI(
        C[760]), .S(S[760]), .CO(C[761]) );
  FA_15943 \FA_INST_0[1].FA_INST_1[249].FA_  ( .A(A[761]), .B(B[761]), .CI(
        C[761]), .S(S[761]), .CO(C[762]) );
  FA_15942 \FA_INST_0[1].FA_INST_1[250].FA_  ( .A(A[762]), .B(B[762]), .CI(
        C[762]), .S(S[762]), .CO(C[763]) );
  FA_15941 \FA_INST_0[1].FA_INST_1[251].FA_  ( .A(A[763]), .B(B[763]), .CI(
        C[763]), .S(S[763]), .CO(C[764]) );
  FA_15940 \FA_INST_0[1].FA_INST_1[252].FA_  ( .A(A[764]), .B(B[764]), .CI(
        C[764]), .S(S[764]), .CO(C[765]) );
  FA_15939 \FA_INST_0[1].FA_INST_1[253].FA_  ( .A(A[765]), .B(B[765]), .CI(
        C[765]), .S(S[765]), .CO(C[766]) );
  FA_15938 \FA_INST_0[1].FA_INST_1[254].FA_  ( .A(A[766]), .B(B[766]), .CI(
        C[766]), .S(S[766]), .CO(C[767]) );
  FA_15937 \FA_INST_0[1].FA_INST_1[255].FA_  ( .A(A[767]), .B(B[767]), .CI(
        C[767]), .S(S[767]), .CO(C[768]) );
  FA_15936 \FA_INST_0[1].FA_INST_1[256].FA_  ( .A(A[768]), .B(B[768]), .CI(
        C[768]), .S(S[768]), .CO(C[769]) );
  FA_15935 \FA_INST_0[1].FA_INST_1[257].FA_  ( .A(A[769]), .B(B[769]), .CI(
        C[769]), .S(S[769]), .CO(C[770]) );
  FA_15934 \FA_INST_0[1].FA_INST_1[258].FA_  ( .A(A[770]), .B(B[770]), .CI(
        C[770]), .S(S[770]), .CO(C[771]) );
  FA_15933 \FA_INST_0[1].FA_INST_1[259].FA_  ( .A(A[771]), .B(B[771]), .CI(
        C[771]), .S(S[771]), .CO(C[772]) );
  FA_15932 \FA_INST_0[1].FA_INST_1[260].FA_  ( .A(A[772]), .B(B[772]), .CI(
        C[772]), .S(S[772]), .CO(C[773]) );
  FA_15931 \FA_INST_0[1].FA_INST_1[261].FA_  ( .A(A[773]), .B(B[773]), .CI(
        C[773]), .S(S[773]), .CO(C[774]) );
  FA_15930 \FA_INST_0[1].FA_INST_1[262].FA_  ( .A(A[774]), .B(B[774]), .CI(
        C[774]), .S(S[774]), .CO(C[775]) );
  FA_15929 \FA_INST_0[1].FA_INST_1[263].FA_  ( .A(A[775]), .B(B[775]), .CI(
        C[775]), .S(S[775]), .CO(C[776]) );
  FA_15928 \FA_INST_0[1].FA_INST_1[264].FA_  ( .A(A[776]), .B(B[776]), .CI(
        C[776]), .S(S[776]), .CO(C[777]) );
  FA_15927 \FA_INST_0[1].FA_INST_1[265].FA_  ( .A(A[777]), .B(B[777]), .CI(
        C[777]), .S(S[777]), .CO(C[778]) );
  FA_15926 \FA_INST_0[1].FA_INST_1[266].FA_  ( .A(A[778]), .B(B[778]), .CI(
        C[778]), .S(S[778]), .CO(C[779]) );
  FA_15925 \FA_INST_0[1].FA_INST_1[267].FA_  ( .A(A[779]), .B(B[779]), .CI(
        C[779]), .S(S[779]), .CO(C[780]) );
  FA_15924 \FA_INST_0[1].FA_INST_1[268].FA_  ( .A(A[780]), .B(B[780]), .CI(
        C[780]), .S(S[780]), .CO(C[781]) );
  FA_15923 \FA_INST_0[1].FA_INST_1[269].FA_  ( .A(A[781]), .B(B[781]), .CI(
        C[781]), .S(S[781]), .CO(C[782]) );
  FA_15922 \FA_INST_0[1].FA_INST_1[270].FA_  ( .A(A[782]), .B(B[782]), .CI(
        C[782]), .S(S[782]), .CO(C[783]) );
  FA_15921 \FA_INST_0[1].FA_INST_1[271].FA_  ( .A(A[783]), .B(B[783]), .CI(
        C[783]), .S(S[783]), .CO(C[784]) );
  FA_15920 \FA_INST_0[1].FA_INST_1[272].FA_  ( .A(A[784]), .B(B[784]), .CI(
        C[784]), .S(S[784]), .CO(C[785]) );
  FA_15919 \FA_INST_0[1].FA_INST_1[273].FA_  ( .A(A[785]), .B(B[785]), .CI(
        C[785]), .S(S[785]), .CO(C[786]) );
  FA_15918 \FA_INST_0[1].FA_INST_1[274].FA_  ( .A(A[786]), .B(B[786]), .CI(
        C[786]), .S(S[786]), .CO(C[787]) );
  FA_15917 \FA_INST_0[1].FA_INST_1[275].FA_  ( .A(A[787]), .B(B[787]), .CI(
        C[787]), .S(S[787]), .CO(C[788]) );
  FA_15916 \FA_INST_0[1].FA_INST_1[276].FA_  ( .A(A[788]), .B(B[788]), .CI(
        C[788]), .S(S[788]), .CO(C[789]) );
  FA_15915 \FA_INST_0[1].FA_INST_1[277].FA_  ( .A(A[789]), .B(B[789]), .CI(
        C[789]), .S(S[789]), .CO(C[790]) );
  FA_15914 \FA_INST_0[1].FA_INST_1[278].FA_  ( .A(A[790]), .B(B[790]), .CI(
        C[790]), .S(S[790]), .CO(C[791]) );
  FA_15913 \FA_INST_0[1].FA_INST_1[279].FA_  ( .A(A[791]), .B(B[791]), .CI(
        C[791]), .S(S[791]), .CO(C[792]) );
  FA_15912 \FA_INST_0[1].FA_INST_1[280].FA_  ( .A(A[792]), .B(B[792]), .CI(
        C[792]), .S(S[792]), .CO(C[793]) );
  FA_15911 \FA_INST_0[1].FA_INST_1[281].FA_  ( .A(A[793]), .B(B[793]), .CI(
        C[793]), .S(S[793]), .CO(C[794]) );
  FA_15910 \FA_INST_0[1].FA_INST_1[282].FA_  ( .A(A[794]), .B(B[794]), .CI(
        C[794]), .S(S[794]), .CO(C[795]) );
  FA_15909 \FA_INST_0[1].FA_INST_1[283].FA_  ( .A(A[795]), .B(B[795]), .CI(
        C[795]), .S(S[795]), .CO(C[796]) );
  FA_15908 \FA_INST_0[1].FA_INST_1[284].FA_  ( .A(A[796]), .B(B[796]), .CI(
        C[796]), .S(S[796]), .CO(C[797]) );
  FA_15907 \FA_INST_0[1].FA_INST_1[285].FA_  ( .A(A[797]), .B(B[797]), .CI(
        C[797]), .S(S[797]), .CO(C[798]) );
  FA_15906 \FA_INST_0[1].FA_INST_1[286].FA_  ( .A(A[798]), .B(B[798]), .CI(
        C[798]), .S(S[798]), .CO(C[799]) );
  FA_15905 \FA_INST_0[1].FA_INST_1[287].FA_  ( .A(A[799]), .B(B[799]), .CI(
        C[799]), .S(S[799]), .CO(C[800]) );
  FA_15904 \FA_INST_0[1].FA_INST_1[288].FA_  ( .A(A[800]), .B(B[800]), .CI(
        C[800]), .S(S[800]), .CO(C[801]) );
  FA_15903 \FA_INST_0[1].FA_INST_1[289].FA_  ( .A(A[801]), .B(B[801]), .CI(
        C[801]), .S(S[801]), .CO(C[802]) );
  FA_15902 \FA_INST_0[1].FA_INST_1[290].FA_  ( .A(A[802]), .B(B[802]), .CI(
        C[802]), .S(S[802]), .CO(C[803]) );
  FA_15901 \FA_INST_0[1].FA_INST_1[291].FA_  ( .A(A[803]), .B(B[803]), .CI(
        C[803]), .S(S[803]), .CO(C[804]) );
  FA_15900 \FA_INST_0[1].FA_INST_1[292].FA_  ( .A(A[804]), .B(B[804]), .CI(
        C[804]), .S(S[804]), .CO(C[805]) );
  FA_15899 \FA_INST_0[1].FA_INST_1[293].FA_  ( .A(A[805]), .B(B[805]), .CI(
        C[805]), .S(S[805]), .CO(C[806]) );
  FA_15898 \FA_INST_0[1].FA_INST_1[294].FA_  ( .A(A[806]), .B(B[806]), .CI(
        C[806]), .S(S[806]), .CO(C[807]) );
  FA_15897 \FA_INST_0[1].FA_INST_1[295].FA_  ( .A(A[807]), .B(B[807]), .CI(
        C[807]), .S(S[807]), .CO(C[808]) );
  FA_15896 \FA_INST_0[1].FA_INST_1[296].FA_  ( .A(A[808]), .B(B[808]), .CI(
        C[808]), .S(S[808]), .CO(C[809]) );
  FA_15895 \FA_INST_0[1].FA_INST_1[297].FA_  ( .A(A[809]), .B(B[809]), .CI(
        C[809]), .S(S[809]), .CO(C[810]) );
  FA_15894 \FA_INST_0[1].FA_INST_1[298].FA_  ( .A(A[810]), .B(B[810]), .CI(
        C[810]), .S(S[810]), .CO(C[811]) );
  FA_15893 \FA_INST_0[1].FA_INST_1[299].FA_  ( .A(A[811]), .B(B[811]), .CI(
        C[811]), .S(S[811]), .CO(C[812]) );
  FA_15892 \FA_INST_0[1].FA_INST_1[300].FA_  ( .A(A[812]), .B(B[812]), .CI(
        C[812]), .S(S[812]), .CO(C[813]) );
  FA_15891 \FA_INST_0[1].FA_INST_1[301].FA_  ( .A(A[813]), .B(B[813]), .CI(
        C[813]), .S(S[813]), .CO(C[814]) );
  FA_15890 \FA_INST_0[1].FA_INST_1[302].FA_  ( .A(A[814]), .B(B[814]), .CI(
        C[814]), .S(S[814]), .CO(C[815]) );
  FA_15889 \FA_INST_0[1].FA_INST_1[303].FA_  ( .A(A[815]), .B(B[815]), .CI(
        C[815]), .S(S[815]), .CO(C[816]) );
  FA_15888 \FA_INST_0[1].FA_INST_1[304].FA_  ( .A(A[816]), .B(B[816]), .CI(
        C[816]), .S(S[816]), .CO(C[817]) );
  FA_15887 \FA_INST_0[1].FA_INST_1[305].FA_  ( .A(A[817]), .B(B[817]), .CI(
        C[817]), .S(S[817]), .CO(C[818]) );
  FA_15886 \FA_INST_0[1].FA_INST_1[306].FA_  ( .A(A[818]), .B(B[818]), .CI(
        C[818]), .S(S[818]), .CO(C[819]) );
  FA_15885 \FA_INST_0[1].FA_INST_1[307].FA_  ( .A(A[819]), .B(B[819]), .CI(
        C[819]), .S(S[819]), .CO(C[820]) );
  FA_15884 \FA_INST_0[1].FA_INST_1[308].FA_  ( .A(A[820]), .B(B[820]), .CI(
        C[820]), .S(S[820]), .CO(C[821]) );
  FA_15883 \FA_INST_0[1].FA_INST_1[309].FA_  ( .A(A[821]), .B(B[821]), .CI(
        C[821]), .S(S[821]), .CO(C[822]) );
  FA_15882 \FA_INST_0[1].FA_INST_1[310].FA_  ( .A(A[822]), .B(B[822]), .CI(
        C[822]), .S(S[822]), .CO(C[823]) );
  FA_15881 \FA_INST_0[1].FA_INST_1[311].FA_  ( .A(A[823]), .B(B[823]), .CI(
        C[823]), .S(S[823]), .CO(C[824]) );
  FA_15880 \FA_INST_0[1].FA_INST_1[312].FA_  ( .A(A[824]), .B(B[824]), .CI(
        C[824]), .S(S[824]), .CO(C[825]) );
  FA_15879 \FA_INST_0[1].FA_INST_1[313].FA_  ( .A(A[825]), .B(B[825]), .CI(
        C[825]), .S(S[825]), .CO(C[826]) );
  FA_15878 \FA_INST_0[1].FA_INST_1[314].FA_  ( .A(A[826]), .B(B[826]), .CI(
        C[826]), .S(S[826]), .CO(C[827]) );
  FA_15877 \FA_INST_0[1].FA_INST_1[315].FA_  ( .A(A[827]), .B(B[827]), .CI(
        C[827]), .S(S[827]), .CO(C[828]) );
  FA_15876 \FA_INST_0[1].FA_INST_1[316].FA_  ( .A(A[828]), .B(B[828]), .CI(
        C[828]), .S(S[828]), .CO(C[829]) );
  FA_15875 \FA_INST_0[1].FA_INST_1[317].FA_  ( .A(A[829]), .B(B[829]), .CI(
        C[829]), .S(S[829]), .CO(C[830]) );
  FA_15874 \FA_INST_0[1].FA_INST_1[318].FA_  ( .A(A[830]), .B(B[830]), .CI(
        C[830]), .S(S[830]), .CO(C[831]) );
  FA_15873 \FA_INST_0[1].FA_INST_1[319].FA_  ( .A(A[831]), .B(B[831]), .CI(
        C[831]), .S(S[831]), .CO(C[832]) );
  FA_15872 \FA_INST_0[1].FA_INST_1[320].FA_  ( .A(A[832]), .B(B[832]), .CI(
        C[832]), .S(S[832]), .CO(C[833]) );
  FA_15871 \FA_INST_0[1].FA_INST_1[321].FA_  ( .A(A[833]), .B(B[833]), .CI(
        C[833]), .S(S[833]), .CO(C[834]) );
  FA_15870 \FA_INST_0[1].FA_INST_1[322].FA_  ( .A(A[834]), .B(B[834]), .CI(
        C[834]), .S(S[834]), .CO(C[835]) );
  FA_15869 \FA_INST_0[1].FA_INST_1[323].FA_  ( .A(A[835]), .B(B[835]), .CI(
        C[835]), .S(S[835]), .CO(C[836]) );
  FA_15868 \FA_INST_0[1].FA_INST_1[324].FA_  ( .A(A[836]), .B(B[836]), .CI(
        C[836]), .S(S[836]), .CO(C[837]) );
  FA_15867 \FA_INST_0[1].FA_INST_1[325].FA_  ( .A(A[837]), .B(B[837]), .CI(
        C[837]), .S(S[837]), .CO(C[838]) );
  FA_15866 \FA_INST_0[1].FA_INST_1[326].FA_  ( .A(A[838]), .B(B[838]), .CI(
        C[838]), .S(S[838]), .CO(C[839]) );
  FA_15865 \FA_INST_0[1].FA_INST_1[327].FA_  ( .A(A[839]), .B(B[839]), .CI(
        C[839]), .S(S[839]), .CO(C[840]) );
  FA_15864 \FA_INST_0[1].FA_INST_1[328].FA_  ( .A(A[840]), .B(B[840]), .CI(
        C[840]), .S(S[840]), .CO(C[841]) );
  FA_15863 \FA_INST_0[1].FA_INST_1[329].FA_  ( .A(A[841]), .B(B[841]), .CI(
        C[841]), .S(S[841]), .CO(C[842]) );
  FA_15862 \FA_INST_0[1].FA_INST_1[330].FA_  ( .A(A[842]), .B(B[842]), .CI(
        C[842]), .S(S[842]), .CO(C[843]) );
  FA_15861 \FA_INST_0[1].FA_INST_1[331].FA_  ( .A(A[843]), .B(B[843]), .CI(
        C[843]), .S(S[843]), .CO(C[844]) );
  FA_15860 \FA_INST_0[1].FA_INST_1[332].FA_  ( .A(A[844]), .B(B[844]), .CI(
        C[844]), .S(S[844]), .CO(C[845]) );
  FA_15859 \FA_INST_0[1].FA_INST_1[333].FA_  ( .A(A[845]), .B(B[845]), .CI(
        C[845]), .S(S[845]), .CO(C[846]) );
  FA_15858 \FA_INST_0[1].FA_INST_1[334].FA_  ( .A(A[846]), .B(B[846]), .CI(
        C[846]), .S(S[846]), .CO(C[847]) );
  FA_15857 \FA_INST_0[1].FA_INST_1[335].FA_  ( .A(A[847]), .B(B[847]), .CI(
        C[847]), .S(S[847]), .CO(C[848]) );
  FA_15856 \FA_INST_0[1].FA_INST_1[336].FA_  ( .A(A[848]), .B(B[848]), .CI(
        C[848]), .S(S[848]), .CO(C[849]) );
  FA_15855 \FA_INST_0[1].FA_INST_1[337].FA_  ( .A(A[849]), .B(B[849]), .CI(
        C[849]), .S(S[849]), .CO(C[850]) );
  FA_15854 \FA_INST_0[1].FA_INST_1[338].FA_  ( .A(A[850]), .B(B[850]), .CI(
        C[850]), .S(S[850]), .CO(C[851]) );
  FA_15853 \FA_INST_0[1].FA_INST_1[339].FA_  ( .A(A[851]), .B(B[851]), .CI(
        C[851]), .S(S[851]), .CO(C[852]) );
  FA_15852 \FA_INST_0[1].FA_INST_1[340].FA_  ( .A(A[852]), .B(B[852]), .CI(
        C[852]), .S(S[852]), .CO(C[853]) );
  FA_15851 \FA_INST_0[1].FA_INST_1[341].FA_  ( .A(A[853]), .B(B[853]), .CI(
        C[853]), .S(S[853]), .CO(C[854]) );
  FA_15850 \FA_INST_0[1].FA_INST_1[342].FA_  ( .A(A[854]), .B(B[854]), .CI(
        C[854]), .S(S[854]), .CO(C[855]) );
  FA_15849 \FA_INST_0[1].FA_INST_1[343].FA_  ( .A(A[855]), .B(B[855]), .CI(
        C[855]), .S(S[855]), .CO(C[856]) );
  FA_15848 \FA_INST_0[1].FA_INST_1[344].FA_  ( .A(A[856]), .B(B[856]), .CI(
        C[856]), .S(S[856]), .CO(C[857]) );
  FA_15847 \FA_INST_0[1].FA_INST_1[345].FA_  ( .A(A[857]), .B(B[857]), .CI(
        C[857]), .S(S[857]), .CO(C[858]) );
  FA_15846 \FA_INST_0[1].FA_INST_1[346].FA_  ( .A(A[858]), .B(B[858]), .CI(
        C[858]), .S(S[858]), .CO(C[859]) );
  FA_15845 \FA_INST_0[1].FA_INST_1[347].FA_  ( .A(A[859]), .B(B[859]), .CI(
        C[859]), .S(S[859]), .CO(C[860]) );
  FA_15844 \FA_INST_0[1].FA_INST_1[348].FA_  ( .A(A[860]), .B(B[860]), .CI(
        C[860]), .S(S[860]), .CO(C[861]) );
  FA_15843 \FA_INST_0[1].FA_INST_1[349].FA_  ( .A(A[861]), .B(B[861]), .CI(
        C[861]), .S(S[861]), .CO(C[862]) );
  FA_15842 \FA_INST_0[1].FA_INST_1[350].FA_  ( .A(A[862]), .B(B[862]), .CI(
        C[862]), .S(S[862]), .CO(C[863]) );
  FA_15841 \FA_INST_0[1].FA_INST_1[351].FA_  ( .A(A[863]), .B(B[863]), .CI(
        C[863]), .S(S[863]), .CO(C[864]) );
  FA_15840 \FA_INST_0[1].FA_INST_1[352].FA_  ( .A(A[864]), .B(B[864]), .CI(
        C[864]), .S(S[864]), .CO(C[865]) );
  FA_15839 \FA_INST_0[1].FA_INST_1[353].FA_  ( .A(A[865]), .B(B[865]), .CI(
        C[865]), .S(S[865]), .CO(C[866]) );
  FA_15838 \FA_INST_0[1].FA_INST_1[354].FA_  ( .A(A[866]), .B(B[866]), .CI(
        C[866]), .S(S[866]), .CO(C[867]) );
  FA_15837 \FA_INST_0[1].FA_INST_1[355].FA_  ( .A(A[867]), .B(B[867]), .CI(
        C[867]), .S(S[867]), .CO(C[868]) );
  FA_15836 \FA_INST_0[1].FA_INST_1[356].FA_  ( .A(A[868]), .B(B[868]), .CI(
        C[868]), .S(S[868]), .CO(C[869]) );
  FA_15835 \FA_INST_0[1].FA_INST_1[357].FA_  ( .A(A[869]), .B(B[869]), .CI(
        C[869]), .S(S[869]), .CO(C[870]) );
  FA_15834 \FA_INST_0[1].FA_INST_1[358].FA_  ( .A(A[870]), .B(B[870]), .CI(
        C[870]), .S(S[870]), .CO(C[871]) );
  FA_15833 \FA_INST_0[1].FA_INST_1[359].FA_  ( .A(A[871]), .B(B[871]), .CI(
        C[871]), .S(S[871]), .CO(C[872]) );
  FA_15832 \FA_INST_0[1].FA_INST_1[360].FA_  ( .A(A[872]), .B(B[872]), .CI(
        C[872]), .S(S[872]), .CO(C[873]) );
  FA_15831 \FA_INST_0[1].FA_INST_1[361].FA_  ( .A(A[873]), .B(B[873]), .CI(
        C[873]), .S(S[873]), .CO(C[874]) );
  FA_15830 \FA_INST_0[1].FA_INST_1[362].FA_  ( .A(A[874]), .B(B[874]), .CI(
        C[874]), .S(S[874]), .CO(C[875]) );
  FA_15829 \FA_INST_0[1].FA_INST_1[363].FA_  ( .A(A[875]), .B(B[875]), .CI(
        C[875]), .S(S[875]), .CO(C[876]) );
  FA_15828 \FA_INST_0[1].FA_INST_1[364].FA_  ( .A(A[876]), .B(B[876]), .CI(
        C[876]), .S(S[876]), .CO(C[877]) );
  FA_15827 \FA_INST_0[1].FA_INST_1[365].FA_  ( .A(A[877]), .B(B[877]), .CI(
        C[877]), .S(S[877]), .CO(C[878]) );
  FA_15826 \FA_INST_0[1].FA_INST_1[366].FA_  ( .A(A[878]), .B(B[878]), .CI(
        C[878]), .S(S[878]), .CO(C[879]) );
  FA_15825 \FA_INST_0[1].FA_INST_1[367].FA_  ( .A(A[879]), .B(B[879]), .CI(
        C[879]), .S(S[879]), .CO(C[880]) );
  FA_15824 \FA_INST_0[1].FA_INST_1[368].FA_  ( .A(A[880]), .B(B[880]), .CI(
        C[880]), .S(S[880]), .CO(C[881]) );
  FA_15823 \FA_INST_0[1].FA_INST_1[369].FA_  ( .A(A[881]), .B(B[881]), .CI(
        C[881]), .S(S[881]), .CO(C[882]) );
  FA_15822 \FA_INST_0[1].FA_INST_1[370].FA_  ( .A(A[882]), .B(B[882]), .CI(
        C[882]), .S(S[882]), .CO(C[883]) );
  FA_15821 \FA_INST_0[1].FA_INST_1[371].FA_  ( .A(A[883]), .B(B[883]), .CI(
        C[883]), .S(S[883]), .CO(C[884]) );
  FA_15820 \FA_INST_0[1].FA_INST_1[372].FA_  ( .A(A[884]), .B(B[884]), .CI(
        C[884]), .S(S[884]), .CO(C[885]) );
  FA_15819 \FA_INST_0[1].FA_INST_1[373].FA_  ( .A(A[885]), .B(B[885]), .CI(
        C[885]), .S(S[885]), .CO(C[886]) );
  FA_15818 \FA_INST_0[1].FA_INST_1[374].FA_  ( .A(A[886]), .B(B[886]), .CI(
        C[886]), .S(S[886]), .CO(C[887]) );
  FA_15817 \FA_INST_0[1].FA_INST_1[375].FA_  ( .A(A[887]), .B(B[887]), .CI(
        C[887]), .S(S[887]), .CO(C[888]) );
  FA_15816 \FA_INST_0[1].FA_INST_1[376].FA_  ( .A(A[888]), .B(B[888]), .CI(
        C[888]), .S(S[888]), .CO(C[889]) );
  FA_15815 \FA_INST_0[1].FA_INST_1[377].FA_  ( .A(A[889]), .B(B[889]), .CI(
        C[889]), .S(S[889]), .CO(C[890]) );
  FA_15814 \FA_INST_0[1].FA_INST_1[378].FA_  ( .A(A[890]), .B(B[890]), .CI(
        C[890]), .S(S[890]), .CO(C[891]) );
  FA_15813 \FA_INST_0[1].FA_INST_1[379].FA_  ( .A(A[891]), .B(B[891]), .CI(
        C[891]), .S(S[891]), .CO(C[892]) );
  FA_15812 \FA_INST_0[1].FA_INST_1[380].FA_  ( .A(A[892]), .B(B[892]), .CI(
        C[892]), .S(S[892]), .CO(C[893]) );
  FA_15811 \FA_INST_0[1].FA_INST_1[381].FA_  ( .A(A[893]), .B(B[893]), .CI(
        C[893]), .S(S[893]), .CO(C[894]) );
  FA_15810 \FA_INST_0[1].FA_INST_1[382].FA_  ( .A(A[894]), .B(B[894]), .CI(
        C[894]), .S(S[894]), .CO(C[895]) );
  FA_15809 \FA_INST_0[1].FA_INST_1[383].FA_  ( .A(A[895]), .B(B[895]), .CI(
        C[895]), .S(S[895]), .CO(C[896]) );
  FA_15808 \FA_INST_0[1].FA_INST_1[384].FA_  ( .A(A[896]), .B(B[896]), .CI(
        C[896]), .S(S[896]), .CO(C[897]) );
  FA_15807 \FA_INST_0[1].FA_INST_1[385].FA_  ( .A(A[897]), .B(B[897]), .CI(
        C[897]), .S(S[897]), .CO(C[898]) );
  FA_15806 \FA_INST_0[1].FA_INST_1[386].FA_  ( .A(A[898]), .B(B[898]), .CI(
        C[898]), .S(S[898]), .CO(C[899]) );
  FA_15805 \FA_INST_0[1].FA_INST_1[387].FA_  ( .A(A[899]), .B(B[899]), .CI(
        C[899]), .S(S[899]), .CO(C[900]) );
  FA_15804 \FA_INST_0[1].FA_INST_1[388].FA_  ( .A(A[900]), .B(B[900]), .CI(
        C[900]), .S(S[900]), .CO(C[901]) );
  FA_15803 \FA_INST_0[1].FA_INST_1[389].FA_  ( .A(A[901]), .B(B[901]), .CI(
        C[901]), .S(S[901]), .CO(C[902]) );
  FA_15802 \FA_INST_0[1].FA_INST_1[390].FA_  ( .A(A[902]), .B(B[902]), .CI(
        C[902]), .S(S[902]), .CO(C[903]) );
  FA_15801 \FA_INST_0[1].FA_INST_1[391].FA_  ( .A(A[903]), .B(B[903]), .CI(
        C[903]), .S(S[903]), .CO(C[904]) );
  FA_15800 \FA_INST_0[1].FA_INST_1[392].FA_  ( .A(A[904]), .B(B[904]), .CI(
        C[904]), .S(S[904]), .CO(C[905]) );
  FA_15799 \FA_INST_0[1].FA_INST_1[393].FA_  ( .A(A[905]), .B(B[905]), .CI(
        C[905]), .S(S[905]), .CO(C[906]) );
  FA_15798 \FA_INST_0[1].FA_INST_1[394].FA_  ( .A(A[906]), .B(B[906]), .CI(
        C[906]), .S(S[906]), .CO(C[907]) );
  FA_15797 \FA_INST_0[1].FA_INST_1[395].FA_  ( .A(A[907]), .B(B[907]), .CI(
        C[907]), .S(S[907]), .CO(C[908]) );
  FA_15796 \FA_INST_0[1].FA_INST_1[396].FA_  ( .A(A[908]), .B(B[908]), .CI(
        C[908]), .S(S[908]), .CO(C[909]) );
  FA_15795 \FA_INST_0[1].FA_INST_1[397].FA_  ( .A(A[909]), .B(B[909]), .CI(
        C[909]), .S(S[909]), .CO(C[910]) );
  FA_15794 \FA_INST_0[1].FA_INST_1[398].FA_  ( .A(A[910]), .B(B[910]), .CI(
        C[910]), .S(S[910]), .CO(C[911]) );
  FA_15793 \FA_INST_0[1].FA_INST_1[399].FA_  ( .A(A[911]), .B(B[911]), .CI(
        C[911]), .S(S[911]), .CO(C[912]) );
  FA_15792 \FA_INST_0[1].FA_INST_1[400].FA_  ( .A(A[912]), .B(B[912]), .CI(
        C[912]), .S(S[912]), .CO(C[913]) );
  FA_15791 \FA_INST_0[1].FA_INST_1[401].FA_  ( .A(A[913]), .B(B[913]), .CI(
        C[913]), .S(S[913]), .CO(C[914]) );
  FA_15790 \FA_INST_0[1].FA_INST_1[402].FA_  ( .A(A[914]), .B(B[914]), .CI(
        C[914]), .S(S[914]), .CO(C[915]) );
  FA_15789 \FA_INST_0[1].FA_INST_1[403].FA_  ( .A(A[915]), .B(B[915]), .CI(
        C[915]), .S(S[915]), .CO(C[916]) );
  FA_15788 \FA_INST_0[1].FA_INST_1[404].FA_  ( .A(A[916]), .B(B[916]), .CI(
        C[916]), .S(S[916]), .CO(C[917]) );
  FA_15787 \FA_INST_0[1].FA_INST_1[405].FA_  ( .A(A[917]), .B(B[917]), .CI(
        C[917]), .S(S[917]), .CO(C[918]) );
  FA_15786 \FA_INST_0[1].FA_INST_1[406].FA_  ( .A(A[918]), .B(B[918]), .CI(
        C[918]), .S(S[918]), .CO(C[919]) );
  FA_15785 \FA_INST_0[1].FA_INST_1[407].FA_  ( .A(A[919]), .B(B[919]), .CI(
        C[919]), .S(S[919]), .CO(C[920]) );
  FA_15784 \FA_INST_0[1].FA_INST_1[408].FA_  ( .A(A[920]), .B(B[920]), .CI(
        C[920]), .S(S[920]), .CO(C[921]) );
  FA_15783 \FA_INST_0[1].FA_INST_1[409].FA_  ( .A(A[921]), .B(B[921]), .CI(
        C[921]), .S(S[921]), .CO(C[922]) );
  FA_15782 \FA_INST_0[1].FA_INST_1[410].FA_  ( .A(A[922]), .B(B[922]), .CI(
        C[922]), .S(S[922]), .CO(C[923]) );
  FA_15781 \FA_INST_0[1].FA_INST_1[411].FA_  ( .A(A[923]), .B(B[923]), .CI(
        C[923]), .S(S[923]), .CO(C[924]) );
  FA_15780 \FA_INST_0[1].FA_INST_1[412].FA_  ( .A(A[924]), .B(B[924]), .CI(
        C[924]), .S(S[924]), .CO(C[925]) );
  FA_15779 \FA_INST_0[1].FA_INST_1[413].FA_  ( .A(A[925]), .B(B[925]), .CI(
        C[925]), .S(S[925]), .CO(C[926]) );
  FA_15778 \FA_INST_0[1].FA_INST_1[414].FA_  ( .A(A[926]), .B(B[926]), .CI(
        C[926]), .S(S[926]), .CO(C[927]) );
  FA_15777 \FA_INST_0[1].FA_INST_1[415].FA_  ( .A(A[927]), .B(B[927]), .CI(
        C[927]), .S(S[927]), .CO(C[928]) );
  FA_15776 \FA_INST_0[1].FA_INST_1[416].FA_  ( .A(A[928]), .B(B[928]), .CI(
        C[928]), .S(S[928]), .CO(C[929]) );
  FA_15775 \FA_INST_0[1].FA_INST_1[417].FA_  ( .A(A[929]), .B(B[929]), .CI(
        C[929]), .S(S[929]), .CO(C[930]) );
  FA_15774 \FA_INST_0[1].FA_INST_1[418].FA_  ( .A(A[930]), .B(B[930]), .CI(
        C[930]), .S(S[930]), .CO(C[931]) );
  FA_15773 \FA_INST_0[1].FA_INST_1[419].FA_  ( .A(A[931]), .B(B[931]), .CI(
        C[931]), .S(S[931]), .CO(C[932]) );
  FA_15772 \FA_INST_0[1].FA_INST_1[420].FA_  ( .A(A[932]), .B(B[932]), .CI(
        C[932]), .S(S[932]), .CO(C[933]) );
  FA_15771 \FA_INST_0[1].FA_INST_1[421].FA_  ( .A(A[933]), .B(B[933]), .CI(
        C[933]), .S(S[933]), .CO(C[934]) );
  FA_15770 \FA_INST_0[1].FA_INST_1[422].FA_  ( .A(A[934]), .B(B[934]), .CI(
        C[934]), .S(S[934]), .CO(C[935]) );
  FA_15769 \FA_INST_0[1].FA_INST_1[423].FA_  ( .A(A[935]), .B(B[935]), .CI(
        C[935]), .S(S[935]), .CO(C[936]) );
  FA_15768 \FA_INST_0[1].FA_INST_1[424].FA_  ( .A(A[936]), .B(B[936]), .CI(
        C[936]), .S(S[936]), .CO(C[937]) );
  FA_15767 \FA_INST_0[1].FA_INST_1[425].FA_  ( .A(A[937]), .B(B[937]), .CI(
        C[937]), .S(S[937]), .CO(C[938]) );
  FA_15766 \FA_INST_0[1].FA_INST_1[426].FA_  ( .A(A[938]), .B(B[938]), .CI(
        C[938]), .S(S[938]), .CO(C[939]) );
  FA_15765 \FA_INST_0[1].FA_INST_1[427].FA_  ( .A(A[939]), .B(B[939]), .CI(
        C[939]), .S(S[939]), .CO(C[940]) );
  FA_15764 \FA_INST_0[1].FA_INST_1[428].FA_  ( .A(A[940]), .B(B[940]), .CI(
        C[940]), .S(S[940]), .CO(C[941]) );
  FA_15763 \FA_INST_0[1].FA_INST_1[429].FA_  ( .A(A[941]), .B(B[941]), .CI(
        C[941]), .S(S[941]), .CO(C[942]) );
  FA_15762 \FA_INST_0[1].FA_INST_1[430].FA_  ( .A(A[942]), .B(B[942]), .CI(
        C[942]), .S(S[942]), .CO(C[943]) );
  FA_15761 \FA_INST_0[1].FA_INST_1[431].FA_  ( .A(A[943]), .B(B[943]), .CI(
        C[943]), .S(S[943]), .CO(C[944]) );
  FA_15760 \FA_INST_0[1].FA_INST_1[432].FA_  ( .A(A[944]), .B(B[944]), .CI(
        C[944]), .S(S[944]), .CO(C[945]) );
  FA_15759 \FA_INST_0[1].FA_INST_1[433].FA_  ( .A(A[945]), .B(B[945]), .CI(
        C[945]), .S(S[945]), .CO(C[946]) );
  FA_15758 \FA_INST_0[1].FA_INST_1[434].FA_  ( .A(A[946]), .B(B[946]), .CI(
        C[946]), .S(S[946]), .CO(C[947]) );
  FA_15757 \FA_INST_0[1].FA_INST_1[435].FA_  ( .A(A[947]), .B(B[947]), .CI(
        C[947]), .S(S[947]), .CO(C[948]) );
  FA_15756 \FA_INST_0[1].FA_INST_1[436].FA_  ( .A(A[948]), .B(B[948]), .CI(
        C[948]), .S(S[948]), .CO(C[949]) );
  FA_15755 \FA_INST_0[1].FA_INST_1[437].FA_  ( .A(A[949]), .B(B[949]), .CI(
        C[949]), .S(S[949]), .CO(C[950]) );
  FA_15754 \FA_INST_0[1].FA_INST_1[438].FA_  ( .A(A[950]), .B(B[950]), .CI(
        C[950]), .S(S[950]), .CO(C[951]) );
  FA_15753 \FA_INST_0[1].FA_INST_1[439].FA_  ( .A(A[951]), .B(B[951]), .CI(
        C[951]), .S(S[951]), .CO(C[952]) );
  FA_15752 \FA_INST_0[1].FA_INST_1[440].FA_  ( .A(A[952]), .B(B[952]), .CI(
        C[952]), .S(S[952]), .CO(C[953]) );
  FA_15751 \FA_INST_0[1].FA_INST_1[441].FA_  ( .A(A[953]), .B(B[953]), .CI(
        C[953]), .S(S[953]), .CO(C[954]) );
  FA_15750 \FA_INST_0[1].FA_INST_1[442].FA_  ( .A(A[954]), .B(B[954]), .CI(
        C[954]), .S(S[954]), .CO(C[955]) );
  FA_15749 \FA_INST_0[1].FA_INST_1[443].FA_  ( .A(A[955]), .B(B[955]), .CI(
        C[955]), .S(S[955]), .CO(C[956]) );
  FA_15748 \FA_INST_0[1].FA_INST_1[444].FA_  ( .A(A[956]), .B(B[956]), .CI(
        C[956]), .S(S[956]), .CO(C[957]) );
  FA_15747 \FA_INST_0[1].FA_INST_1[445].FA_  ( .A(A[957]), .B(B[957]), .CI(
        C[957]), .S(S[957]), .CO(C[958]) );
  FA_15746 \FA_INST_0[1].FA_INST_1[446].FA_  ( .A(A[958]), .B(B[958]), .CI(
        C[958]), .S(S[958]), .CO(C[959]) );
  FA_15745 \FA_INST_0[1].FA_INST_1[447].FA_  ( .A(A[959]), .B(B[959]), .CI(
        C[959]), .S(S[959]), .CO(C[960]) );
  FA_15744 \FA_INST_0[1].FA_INST_1[448].FA_  ( .A(A[960]), .B(B[960]), .CI(
        C[960]), .S(S[960]), .CO(C[961]) );
  FA_15743 \FA_INST_0[1].FA_INST_1[449].FA_  ( .A(A[961]), .B(B[961]), .CI(
        C[961]), .S(S[961]), .CO(C[962]) );
  FA_15742 \FA_INST_0[1].FA_INST_1[450].FA_  ( .A(A[962]), .B(B[962]), .CI(
        C[962]), .S(S[962]), .CO(C[963]) );
  FA_15741 \FA_INST_0[1].FA_INST_1[451].FA_  ( .A(A[963]), .B(B[963]), .CI(
        C[963]), .S(S[963]), .CO(C[964]) );
  FA_15740 \FA_INST_0[1].FA_INST_1[452].FA_  ( .A(A[964]), .B(B[964]), .CI(
        C[964]), .S(S[964]), .CO(C[965]) );
  FA_15739 \FA_INST_0[1].FA_INST_1[453].FA_  ( .A(A[965]), .B(B[965]), .CI(
        C[965]), .S(S[965]), .CO(C[966]) );
  FA_15738 \FA_INST_0[1].FA_INST_1[454].FA_  ( .A(A[966]), .B(B[966]), .CI(
        C[966]), .S(S[966]), .CO(C[967]) );
  FA_15737 \FA_INST_0[1].FA_INST_1[455].FA_  ( .A(A[967]), .B(B[967]), .CI(
        C[967]), .S(S[967]), .CO(C[968]) );
  FA_15736 \FA_INST_0[1].FA_INST_1[456].FA_  ( .A(A[968]), .B(B[968]), .CI(
        C[968]), .S(S[968]), .CO(C[969]) );
  FA_15735 \FA_INST_0[1].FA_INST_1[457].FA_  ( .A(A[969]), .B(B[969]), .CI(
        C[969]), .S(S[969]), .CO(C[970]) );
  FA_15734 \FA_INST_0[1].FA_INST_1[458].FA_  ( .A(A[970]), .B(B[970]), .CI(
        C[970]), .S(S[970]), .CO(C[971]) );
  FA_15733 \FA_INST_0[1].FA_INST_1[459].FA_  ( .A(A[971]), .B(B[971]), .CI(
        C[971]), .S(S[971]), .CO(C[972]) );
  FA_15732 \FA_INST_0[1].FA_INST_1[460].FA_  ( .A(A[972]), .B(B[972]), .CI(
        C[972]), .S(S[972]), .CO(C[973]) );
  FA_15731 \FA_INST_0[1].FA_INST_1[461].FA_  ( .A(A[973]), .B(B[973]), .CI(
        C[973]), .S(S[973]), .CO(C[974]) );
  FA_15730 \FA_INST_0[1].FA_INST_1[462].FA_  ( .A(A[974]), .B(B[974]), .CI(
        C[974]), .S(S[974]), .CO(C[975]) );
  FA_15729 \FA_INST_0[1].FA_INST_1[463].FA_  ( .A(A[975]), .B(B[975]), .CI(
        C[975]), .S(S[975]), .CO(C[976]) );
  FA_15728 \FA_INST_0[1].FA_INST_1[464].FA_  ( .A(A[976]), .B(B[976]), .CI(
        C[976]), .S(S[976]), .CO(C[977]) );
  FA_15727 \FA_INST_0[1].FA_INST_1[465].FA_  ( .A(A[977]), .B(B[977]), .CI(
        C[977]), .S(S[977]), .CO(C[978]) );
  FA_15726 \FA_INST_0[1].FA_INST_1[466].FA_  ( .A(A[978]), .B(B[978]), .CI(
        C[978]), .S(S[978]), .CO(C[979]) );
  FA_15725 \FA_INST_0[1].FA_INST_1[467].FA_  ( .A(A[979]), .B(B[979]), .CI(
        C[979]), .S(S[979]), .CO(C[980]) );
  FA_15724 \FA_INST_0[1].FA_INST_1[468].FA_  ( .A(A[980]), .B(B[980]), .CI(
        C[980]), .S(S[980]), .CO(C[981]) );
  FA_15723 \FA_INST_0[1].FA_INST_1[469].FA_  ( .A(A[981]), .B(B[981]), .CI(
        C[981]), .S(S[981]), .CO(C[982]) );
  FA_15722 \FA_INST_0[1].FA_INST_1[470].FA_  ( .A(A[982]), .B(B[982]), .CI(
        C[982]), .S(S[982]), .CO(C[983]) );
  FA_15721 \FA_INST_0[1].FA_INST_1[471].FA_  ( .A(A[983]), .B(B[983]), .CI(
        C[983]), .S(S[983]), .CO(C[984]) );
  FA_15720 \FA_INST_0[1].FA_INST_1[472].FA_  ( .A(A[984]), .B(B[984]), .CI(
        C[984]), .S(S[984]), .CO(C[985]) );
  FA_15719 \FA_INST_0[1].FA_INST_1[473].FA_  ( .A(A[985]), .B(B[985]), .CI(
        C[985]), .S(S[985]), .CO(C[986]) );
  FA_15718 \FA_INST_0[1].FA_INST_1[474].FA_  ( .A(A[986]), .B(B[986]), .CI(
        C[986]), .S(S[986]), .CO(C[987]) );
  FA_15717 \FA_INST_0[1].FA_INST_1[475].FA_  ( .A(A[987]), .B(B[987]), .CI(
        C[987]), .S(S[987]), .CO(C[988]) );
  FA_15716 \FA_INST_0[1].FA_INST_1[476].FA_  ( .A(A[988]), .B(B[988]), .CI(
        C[988]), .S(S[988]), .CO(C[989]) );
  FA_15715 \FA_INST_0[1].FA_INST_1[477].FA_  ( .A(A[989]), .B(B[989]), .CI(
        C[989]), .S(S[989]), .CO(C[990]) );
  FA_15714 \FA_INST_0[1].FA_INST_1[478].FA_  ( .A(A[990]), .B(B[990]), .CI(
        C[990]), .S(S[990]), .CO(C[991]) );
  FA_15713 \FA_INST_0[1].FA_INST_1[479].FA_  ( .A(A[991]), .B(B[991]), .CI(
        C[991]), .S(S[991]), .CO(C[992]) );
  FA_15712 \FA_INST_0[1].FA_INST_1[480].FA_  ( .A(A[992]), .B(B[992]), .CI(
        C[992]), .S(S[992]), .CO(C[993]) );
  FA_15711 \FA_INST_0[1].FA_INST_1[481].FA_  ( .A(A[993]), .B(B[993]), .CI(
        C[993]), .S(S[993]), .CO(C[994]) );
  FA_15710 \FA_INST_0[1].FA_INST_1[482].FA_  ( .A(A[994]), .B(B[994]), .CI(
        C[994]), .S(S[994]), .CO(C[995]) );
  FA_15709 \FA_INST_0[1].FA_INST_1[483].FA_  ( .A(A[995]), .B(B[995]), .CI(
        C[995]), .S(S[995]), .CO(C[996]) );
  FA_15708 \FA_INST_0[1].FA_INST_1[484].FA_  ( .A(A[996]), .B(B[996]), .CI(
        C[996]), .S(S[996]), .CO(C[997]) );
  FA_15707 \FA_INST_0[1].FA_INST_1[485].FA_  ( .A(A[997]), .B(B[997]), .CI(
        C[997]), .S(S[997]), .CO(C[998]) );
  FA_15706 \FA_INST_0[1].FA_INST_1[486].FA_  ( .A(A[998]), .B(B[998]), .CI(
        C[998]), .S(S[998]), .CO(C[999]) );
  FA_15705 \FA_INST_0[1].FA_INST_1[487].FA_  ( .A(A[999]), .B(B[999]), .CI(
        C[999]), .S(S[999]), .CO(C[1000]) );
  FA_15704 \FA_INST_0[1].FA_INST_1[488].FA_  ( .A(A[1000]), .B(B[1000]), .CI(
        C[1000]), .S(S[1000]), .CO(C[1001]) );
  FA_15703 \FA_INST_0[1].FA_INST_1[489].FA_  ( .A(A[1001]), .B(B[1001]), .CI(
        C[1001]), .S(S[1001]), .CO(C[1002]) );
  FA_15702 \FA_INST_0[1].FA_INST_1[490].FA_  ( .A(A[1002]), .B(B[1002]), .CI(
        C[1002]), .S(S[1002]), .CO(C[1003]) );
  FA_15701 \FA_INST_0[1].FA_INST_1[491].FA_  ( .A(A[1003]), .B(B[1003]), .CI(
        C[1003]), .S(S[1003]), .CO(C[1004]) );
  FA_15700 \FA_INST_0[1].FA_INST_1[492].FA_  ( .A(A[1004]), .B(B[1004]), .CI(
        C[1004]), .S(S[1004]), .CO(C[1005]) );
  FA_15699 \FA_INST_0[1].FA_INST_1[493].FA_  ( .A(A[1005]), .B(B[1005]), .CI(
        C[1005]), .S(S[1005]), .CO(C[1006]) );
  FA_15698 \FA_INST_0[1].FA_INST_1[494].FA_  ( .A(A[1006]), .B(B[1006]), .CI(
        C[1006]), .S(S[1006]), .CO(C[1007]) );
  FA_15697 \FA_INST_0[1].FA_INST_1[495].FA_  ( .A(A[1007]), .B(B[1007]), .CI(
        C[1007]), .S(S[1007]), .CO(C[1008]) );
  FA_15696 \FA_INST_0[1].FA_INST_1[496].FA_  ( .A(A[1008]), .B(B[1008]), .CI(
        C[1008]), .S(S[1008]), .CO(C[1009]) );
  FA_15695 \FA_INST_0[1].FA_INST_1[497].FA_  ( .A(A[1009]), .B(B[1009]), .CI(
        C[1009]), .S(S[1009]), .CO(C[1010]) );
  FA_15694 \FA_INST_0[1].FA_INST_1[498].FA_  ( .A(A[1010]), .B(B[1010]), .CI(
        C[1010]), .S(S[1010]), .CO(C[1011]) );
  FA_15693 \FA_INST_0[1].FA_INST_1[499].FA_  ( .A(A[1011]), .B(B[1011]), .CI(
        C[1011]), .S(S[1011]), .CO(C[1012]) );
  FA_15692 \FA_INST_0[1].FA_INST_1[500].FA_  ( .A(A[1012]), .B(B[1012]), .CI(
        C[1012]), .S(S[1012]), .CO(C[1013]) );
  FA_15691 \FA_INST_0[1].FA_INST_1[501].FA_  ( .A(A[1013]), .B(B[1013]), .CI(
        C[1013]), .S(S[1013]), .CO(C[1014]) );
  FA_15690 \FA_INST_0[1].FA_INST_1[502].FA_  ( .A(A[1014]), .B(B[1014]), .CI(
        C[1014]), .S(S[1014]), .CO(C[1015]) );
  FA_15689 \FA_INST_0[1].FA_INST_1[503].FA_  ( .A(A[1015]), .B(B[1015]), .CI(
        C[1015]), .S(S[1015]), .CO(C[1016]) );
  FA_15688 \FA_INST_0[1].FA_INST_1[504].FA_  ( .A(A[1016]), .B(B[1016]), .CI(
        C[1016]), .S(S[1016]), .CO(C[1017]) );
  FA_15687 \FA_INST_0[1].FA_INST_1[505].FA_  ( .A(A[1017]), .B(B[1017]), .CI(
        C[1017]), .S(S[1017]), .CO(C[1018]) );
  FA_15686 \FA_INST_0[1].FA_INST_1[506].FA_  ( .A(A[1018]), .B(B[1018]), .CI(
        C[1018]), .S(S[1018]), .CO(C[1019]) );
  FA_15685 \FA_INST_0[1].FA_INST_1[507].FA_  ( .A(A[1019]), .B(B[1019]), .CI(
        C[1019]), .S(S[1019]), .CO(C[1020]) );
  FA_15684 \FA_INST_0[1].FA_INST_1[508].FA_  ( .A(A[1020]), .B(B[1020]), .CI(
        C[1020]), .S(S[1020]), .CO(C[1021]) );
  FA_15683 \FA_INST_0[1].FA_INST_1[509].FA_  ( .A(A[1021]), .B(B[1021]), .CI(
        C[1021]), .S(S[1021]), .CO(C[1022]) );
  FA_15682 \FA_INST_0[1].FA_INST_1[510].FA_  ( .A(A[1022]), .B(B[1022]), .CI(
        C[1022]), .S(S[1022]), .CO(C[1023]) );
  FA_15681 \FA_INST_0[1].FA_INST_1[511].FA_  ( .A(A[1023]), .B(B[1023]), .CI(
        C[1023]), .S(S[1023]), .CO(C[1024]) );
  FA_15680 \FA_INST_1[1024].FA_  ( .A(A[1024]), .B(1'b0), .CI(C[1024]), .S(
        S[1024]), .CO(C[1025]) );
  FA_15679 \FA_INST_1[1025].FA_  ( .A(A[1025]), .B(1'b0), .CI(C[1025]), .S(
        S[1025]) );
endmodule


module FA_14653 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  OR U1 ( .A(CI), .B(A), .Z(CO) );
endmodule


module FA_14654 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  OR U1 ( .A(CI), .B(A), .Z(CO) );
endmodule


module FA_14655 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14656 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14657 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14658 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14659 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14660 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14661 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14662 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14663 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14664 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14665 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14666 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14667 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14668 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14669 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14670 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14671 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14672 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14673 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14674 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14675 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14676 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14677 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14678 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14679 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14680 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14681 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14682 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14683 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14684 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14685 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14686 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14687 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14688 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14689 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14690 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14691 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14692 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14693 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14694 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14695 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14696 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14697 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14698 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14699 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14700 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14701 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14702 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14703 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14704 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14705 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14706 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14707 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14708 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14709 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14710 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14711 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14712 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14713 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14714 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14715 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14716 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14717 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14718 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14719 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14720 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14721 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14722 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14723 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14724 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14725 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14726 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14727 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14728 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14729 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14730 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14731 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14732 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14733 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14734 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14735 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14736 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14737 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14738 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14739 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14740 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14741 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14742 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14743 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14744 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14745 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14746 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14747 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14748 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14749 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14750 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14751 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14752 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14753 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14754 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14755 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14756 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14757 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14758 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14759 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14760 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14761 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14762 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14763 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14764 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14765 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14766 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14767 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14768 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14769 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14770 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14771 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14772 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14773 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14774 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14775 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14776 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14777 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14778 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14779 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14780 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14781 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14782 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14783 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14784 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14785 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14786 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14787 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14788 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14789 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14790 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14791 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14792 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14793 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14794 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14795 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14796 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14797 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14798 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14799 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14800 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14801 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14802 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14803 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14804 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14805 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14806 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14807 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14808 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14809 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14810 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14811 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14812 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14813 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14814 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14815 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14816 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14817 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14818 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14819 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14820 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14821 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14822 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14823 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14824 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14825 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14826 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14827 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14828 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14829 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14830 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14831 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14832 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14833 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14834 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14835 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14836 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14837 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14838 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14839 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14840 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14841 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14842 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14843 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14844 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14845 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14846 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14847 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14848 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14849 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14850 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14851 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14852 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14853 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14854 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14855 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14856 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14857 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14858 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14859 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14860 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14861 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14862 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14863 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14864 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14865 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14866 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14867 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14868 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14869 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14870 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14871 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14872 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14873 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14874 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14875 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14876 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14877 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14878 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14879 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14880 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14881 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14882 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14883 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14884 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14885 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14886 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14887 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14888 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14889 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14890 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14891 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14892 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14893 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14894 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14895 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14896 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14897 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14898 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14899 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14900 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14901 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14902 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14903 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14904 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14905 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14906 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14907 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14908 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14909 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14910 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14911 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14912 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14913 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14914 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14915 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14916 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14917 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14918 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14919 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14920 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14921 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14922 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14923 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14924 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14925 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14926 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14927 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14928 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14929 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14930 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14931 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14932 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14933 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14934 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14935 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14936 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14937 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14938 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14939 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14940 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14941 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14942 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14943 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14944 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14945 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14946 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14947 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14948 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14949 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14950 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14951 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14952 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14953 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14954 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14955 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14956 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14957 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14958 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14959 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14960 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14961 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14962 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14963 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14964 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14965 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14966 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14967 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14968 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14969 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14970 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14971 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14972 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14973 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14974 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14975 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14976 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14977 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14978 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14979 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14980 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14981 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14982 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14983 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14984 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14985 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14986 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14987 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14988 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14989 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14990 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14991 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14992 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14993 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14994 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14995 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14996 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14997 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14998 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_14999 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15000 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15001 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15002 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15003 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15004 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15005 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15006 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15007 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15008 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15009 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15010 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15011 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15012 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15013 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15014 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15015 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15016 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15017 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15018 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15019 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15020 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15021 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15022 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15023 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15024 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15025 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15026 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15027 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15028 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15029 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15030 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15031 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15032 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15033 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15034 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15035 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15036 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15037 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15038 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15039 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15040 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15041 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15042 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15043 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15044 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15045 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15046 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15047 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15048 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15049 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15050 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15051 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15052 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15053 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15054 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15055 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15056 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15057 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15058 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15059 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15060 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15061 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15062 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15063 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15064 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15065 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15066 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15067 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15068 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15069 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15070 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15071 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15072 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15073 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15074 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15075 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15076 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15077 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15078 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15079 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15080 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15081 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15082 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15083 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15084 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15085 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15086 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15087 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15088 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15089 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15090 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15091 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15092 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15093 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15094 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15095 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15096 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15097 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15098 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15099 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15100 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15101 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15102 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15103 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15104 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15105 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15106 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15107 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15108 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15109 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15110 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15111 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15112 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15113 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15114 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15115 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15116 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15117 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15118 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15119 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15120 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15121 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15122 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15123 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15124 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15125 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15126 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15127 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15128 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15129 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15130 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15131 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15132 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15133 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15134 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15135 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15136 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15137 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15138 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15139 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15140 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15141 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15142 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15143 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15144 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15145 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15146 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15147 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15148 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15149 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15150 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15151 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15152 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15153 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15154 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15155 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15156 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15157 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15158 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15159 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15160 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15161 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15162 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15163 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15164 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15165 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15166 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15167 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15168 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15169 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15170 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15171 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15172 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15173 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15174 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15175 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15176 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15177 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15178 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15179 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15180 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15181 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15182 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15183 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15184 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15185 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15186 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15187 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15188 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15189 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15190 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15191 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15192 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15193 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15194 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15195 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15196 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15197 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15198 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15199 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15200 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15201 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15202 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15203 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15204 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15205 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15206 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15207 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15208 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15209 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15210 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15211 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15212 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15213 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15214 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15215 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15216 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15217 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15218 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15219 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15220 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15221 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15222 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15223 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15224 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15225 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15226 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15227 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15228 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15229 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15230 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15231 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15232 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15233 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15234 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15235 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15236 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15237 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15238 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15239 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15240 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15241 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15242 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15243 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15244 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15245 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15246 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15247 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15248 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15249 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15250 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15251 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15252 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15253 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15254 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15255 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15256 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15257 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15258 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15259 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15260 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15261 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15262 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15263 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15264 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15265 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15266 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15267 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15268 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15269 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15270 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15271 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15272 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15273 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15274 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15275 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15276 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15277 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15278 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15279 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15280 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15281 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15282 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15283 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15284 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15285 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15286 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15287 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15288 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15289 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15290 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15291 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15292 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15293 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15294 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15295 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15296 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15297 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15298 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15299 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15300 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15301 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15302 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15303 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15304 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15305 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15306 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15307 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15308 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15309 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15310 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15311 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15312 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15313 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15314 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15315 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15316 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15317 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15318 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15319 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15320 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15321 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15322 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15323 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15324 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15325 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15326 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15327 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15328 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15329 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15330 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15331 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15332 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15333 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15334 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15335 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15336 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15337 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15338 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15339 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15340 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15341 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15342 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15343 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15344 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15345 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15346 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15347 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15348 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15349 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15350 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15351 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15352 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15353 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15354 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15355 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15356 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15357 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15358 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15359 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15360 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15361 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15362 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15363 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15364 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15365 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15366 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15367 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15368 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15369 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15370 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15371 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15372 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15373 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15374 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15375 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15376 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15377 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15378 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15379 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15380 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15381 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15382 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15383 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15384 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15385 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15386 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15387 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15388 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15389 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15390 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15391 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15392 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15393 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15394 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15395 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15396 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15397 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15398 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15399 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15400 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15401 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15402 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15403 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15404 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15405 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15406 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15407 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15408 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15409 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15410 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15411 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15412 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15413 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15414 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15415 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15416 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15417 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15418 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15419 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15420 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15421 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15422 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15423 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15424 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15425 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15426 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15427 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15428 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15429 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15430 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15431 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15432 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15433 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15434 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15435 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15436 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15437 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15438 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15439 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15440 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15441 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15442 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15443 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15444 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15445 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15446 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15447 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15448 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15449 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15450 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15451 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15452 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15453 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15454 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15455 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15456 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15457 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15458 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15459 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15460 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15461 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15462 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15463 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15464 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15465 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15466 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15467 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15468 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15469 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15470 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15471 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15472 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15473 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15474 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15475 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15476 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15477 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15478 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15479 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15480 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15481 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15482 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15483 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15484 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15485 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15486 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15487 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15488 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15489 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15490 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15491 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15492 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15493 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15494 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15495 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15496 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15497 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15498 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15499 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15500 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15501 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15502 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15503 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15504 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15505 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15506 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15507 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15508 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15509 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15510 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15511 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15512 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15513 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15514 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15515 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15516 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15517 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15518 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15519 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15520 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15521 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15522 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15523 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15524 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15525 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15526 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15527 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15528 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15529 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15530 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15531 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15532 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15533 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15534 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15535 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15536 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15537 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15538 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15539 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15540 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15541 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15542 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15543 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15544 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15545 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15546 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15547 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15548 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15549 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15550 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15551 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15552 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15553 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15554 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15555 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15556 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15557 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15558 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15559 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15560 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15561 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15562 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15563 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15564 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15565 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15566 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15567 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15568 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15569 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15570 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15571 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15572 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15573 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15574 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15575 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15576 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15577 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15578 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15579 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15580 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15581 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15582 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15583 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15584 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15585 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15586 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15587 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15588 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15589 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15590 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15591 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15592 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15593 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15594 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15595 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15596 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15597 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15598 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15599 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15600 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15601 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15602 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15603 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15604 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15605 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15606 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15607 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15608 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15609 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15610 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15611 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15612 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15613 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15614 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15615 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15616 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15617 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15618 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15619 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15620 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15621 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15622 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15623 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15624 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15625 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15626 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15627 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15628 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15629 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15630 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15631 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15632 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15633 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15634 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15635 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15636 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15637 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15638 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15639 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15640 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15641 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15642 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15643 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15644 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15645 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15646 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15647 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15648 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15649 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15650 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15651 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15652 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15653 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15654 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15655 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15656 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15657 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15658 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15659 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15660 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15661 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15662 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15663 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15664 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15665 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15666 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15667 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15668 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15669 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15670 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15671 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15672 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15673 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15674 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15675 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15676 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15677 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_15678 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  OR U1 ( .A(B), .B(A), .Z(CO) );
endmodule


module COMP_N1026_0 ( A, B, O );
  input [1025:0] A;
  input [1025:0] B;
  output O;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026;
  wire   [1025:1] C;

  FA_15678 \FA_INST_0[0].FA_INST_1[0].FA_  ( .A(A[0]), .B(n1026), .CI(1'b1), 
        .CO(C[1]) );
  FA_15677 \FA_INST_0[0].FA_INST_1[1].FA_  ( .A(A[1]), .B(n1025), .CI(C[1]), 
        .CO(C[2]) );
  FA_15676 \FA_INST_0[0].FA_INST_1[2].FA_  ( .A(A[2]), .B(n1024), .CI(C[2]), 
        .CO(C[3]) );
  FA_15675 \FA_INST_0[0].FA_INST_1[3].FA_  ( .A(A[3]), .B(n1023), .CI(C[3]), 
        .CO(C[4]) );
  FA_15674 \FA_INST_0[0].FA_INST_1[4].FA_  ( .A(A[4]), .B(n1022), .CI(C[4]), 
        .CO(C[5]) );
  FA_15673 \FA_INST_0[0].FA_INST_1[5].FA_  ( .A(A[5]), .B(n1021), .CI(C[5]), 
        .CO(C[6]) );
  FA_15672 \FA_INST_0[0].FA_INST_1[6].FA_  ( .A(A[6]), .B(n1020), .CI(C[6]), 
        .CO(C[7]) );
  FA_15671 \FA_INST_0[0].FA_INST_1[7].FA_  ( .A(A[7]), .B(n1019), .CI(C[7]), 
        .CO(C[8]) );
  FA_15670 \FA_INST_0[0].FA_INST_1[8].FA_  ( .A(A[8]), .B(n1018), .CI(C[8]), 
        .CO(C[9]) );
  FA_15669 \FA_INST_0[0].FA_INST_1[9].FA_  ( .A(A[9]), .B(n1017), .CI(C[9]), 
        .CO(C[10]) );
  FA_15668 \FA_INST_0[0].FA_INST_1[10].FA_  ( .A(A[10]), .B(n1016), .CI(C[10]), 
        .CO(C[11]) );
  FA_15667 \FA_INST_0[0].FA_INST_1[11].FA_  ( .A(A[11]), .B(n1015), .CI(C[11]), 
        .CO(C[12]) );
  FA_15666 \FA_INST_0[0].FA_INST_1[12].FA_  ( .A(A[12]), .B(n1014), .CI(C[12]), 
        .CO(C[13]) );
  FA_15665 \FA_INST_0[0].FA_INST_1[13].FA_  ( .A(A[13]), .B(n1013), .CI(C[13]), 
        .CO(C[14]) );
  FA_15664 \FA_INST_0[0].FA_INST_1[14].FA_  ( .A(A[14]), .B(n1012), .CI(C[14]), 
        .CO(C[15]) );
  FA_15663 \FA_INST_0[0].FA_INST_1[15].FA_  ( .A(A[15]), .B(n1011), .CI(C[15]), 
        .CO(C[16]) );
  FA_15662 \FA_INST_0[0].FA_INST_1[16].FA_  ( .A(A[16]), .B(n1010), .CI(C[16]), 
        .CO(C[17]) );
  FA_15661 \FA_INST_0[0].FA_INST_1[17].FA_  ( .A(A[17]), .B(n1009), .CI(C[17]), 
        .CO(C[18]) );
  FA_15660 \FA_INST_0[0].FA_INST_1[18].FA_  ( .A(A[18]), .B(n1008), .CI(C[18]), 
        .CO(C[19]) );
  FA_15659 \FA_INST_0[0].FA_INST_1[19].FA_  ( .A(A[19]), .B(n1007), .CI(C[19]), 
        .CO(C[20]) );
  FA_15658 \FA_INST_0[0].FA_INST_1[20].FA_  ( .A(A[20]), .B(n1006), .CI(C[20]), 
        .CO(C[21]) );
  FA_15657 \FA_INST_0[0].FA_INST_1[21].FA_  ( .A(A[21]), .B(n1005), .CI(C[21]), 
        .CO(C[22]) );
  FA_15656 \FA_INST_0[0].FA_INST_1[22].FA_  ( .A(A[22]), .B(n1004), .CI(C[22]), 
        .CO(C[23]) );
  FA_15655 \FA_INST_0[0].FA_INST_1[23].FA_  ( .A(A[23]), .B(n1003), .CI(C[23]), 
        .CO(C[24]) );
  FA_15654 \FA_INST_0[0].FA_INST_1[24].FA_  ( .A(A[24]), .B(n1002), .CI(C[24]), 
        .CO(C[25]) );
  FA_15653 \FA_INST_0[0].FA_INST_1[25].FA_  ( .A(A[25]), .B(n1001), .CI(C[25]), 
        .CO(C[26]) );
  FA_15652 \FA_INST_0[0].FA_INST_1[26].FA_  ( .A(A[26]), .B(n1000), .CI(C[26]), 
        .CO(C[27]) );
  FA_15651 \FA_INST_0[0].FA_INST_1[27].FA_  ( .A(A[27]), .B(n999), .CI(C[27]), 
        .CO(C[28]) );
  FA_15650 \FA_INST_0[0].FA_INST_1[28].FA_  ( .A(A[28]), .B(n998), .CI(C[28]), 
        .CO(C[29]) );
  FA_15649 \FA_INST_0[0].FA_INST_1[29].FA_  ( .A(A[29]), .B(n997), .CI(C[29]), 
        .CO(C[30]) );
  FA_15648 \FA_INST_0[0].FA_INST_1[30].FA_  ( .A(A[30]), .B(n996), .CI(C[30]), 
        .CO(C[31]) );
  FA_15647 \FA_INST_0[0].FA_INST_1[31].FA_  ( .A(A[31]), .B(n995), .CI(C[31]), 
        .CO(C[32]) );
  FA_15646 \FA_INST_0[0].FA_INST_1[32].FA_  ( .A(A[32]), .B(n994), .CI(C[32]), 
        .CO(C[33]) );
  FA_15645 \FA_INST_0[0].FA_INST_1[33].FA_  ( .A(A[33]), .B(n993), .CI(C[33]), 
        .CO(C[34]) );
  FA_15644 \FA_INST_0[0].FA_INST_1[34].FA_  ( .A(A[34]), .B(n992), .CI(C[34]), 
        .CO(C[35]) );
  FA_15643 \FA_INST_0[0].FA_INST_1[35].FA_  ( .A(A[35]), .B(n991), .CI(C[35]), 
        .CO(C[36]) );
  FA_15642 \FA_INST_0[0].FA_INST_1[36].FA_  ( .A(A[36]), .B(n990), .CI(C[36]), 
        .CO(C[37]) );
  FA_15641 \FA_INST_0[0].FA_INST_1[37].FA_  ( .A(A[37]), .B(n989), .CI(C[37]), 
        .CO(C[38]) );
  FA_15640 \FA_INST_0[0].FA_INST_1[38].FA_  ( .A(A[38]), .B(n988), .CI(C[38]), 
        .CO(C[39]) );
  FA_15639 \FA_INST_0[0].FA_INST_1[39].FA_  ( .A(A[39]), .B(n987), .CI(C[39]), 
        .CO(C[40]) );
  FA_15638 \FA_INST_0[0].FA_INST_1[40].FA_  ( .A(A[40]), .B(n986), .CI(C[40]), 
        .CO(C[41]) );
  FA_15637 \FA_INST_0[0].FA_INST_1[41].FA_  ( .A(A[41]), .B(n985), .CI(C[41]), 
        .CO(C[42]) );
  FA_15636 \FA_INST_0[0].FA_INST_1[42].FA_  ( .A(A[42]), .B(n984), .CI(C[42]), 
        .CO(C[43]) );
  FA_15635 \FA_INST_0[0].FA_INST_1[43].FA_  ( .A(A[43]), .B(n983), .CI(C[43]), 
        .CO(C[44]) );
  FA_15634 \FA_INST_0[0].FA_INST_1[44].FA_  ( .A(A[44]), .B(n982), .CI(C[44]), 
        .CO(C[45]) );
  FA_15633 \FA_INST_0[0].FA_INST_1[45].FA_  ( .A(A[45]), .B(n981), .CI(C[45]), 
        .CO(C[46]) );
  FA_15632 \FA_INST_0[0].FA_INST_1[46].FA_  ( .A(A[46]), .B(n980), .CI(C[46]), 
        .CO(C[47]) );
  FA_15631 \FA_INST_0[0].FA_INST_1[47].FA_  ( .A(A[47]), .B(n979), .CI(C[47]), 
        .CO(C[48]) );
  FA_15630 \FA_INST_0[0].FA_INST_1[48].FA_  ( .A(A[48]), .B(n978), .CI(C[48]), 
        .CO(C[49]) );
  FA_15629 \FA_INST_0[0].FA_INST_1[49].FA_  ( .A(A[49]), .B(n977), .CI(C[49]), 
        .CO(C[50]) );
  FA_15628 \FA_INST_0[0].FA_INST_1[50].FA_  ( .A(A[50]), .B(n976), .CI(C[50]), 
        .CO(C[51]) );
  FA_15627 \FA_INST_0[0].FA_INST_1[51].FA_  ( .A(A[51]), .B(n975), .CI(C[51]), 
        .CO(C[52]) );
  FA_15626 \FA_INST_0[0].FA_INST_1[52].FA_  ( .A(A[52]), .B(n974), .CI(C[52]), 
        .CO(C[53]) );
  FA_15625 \FA_INST_0[0].FA_INST_1[53].FA_  ( .A(A[53]), .B(n973), .CI(C[53]), 
        .CO(C[54]) );
  FA_15624 \FA_INST_0[0].FA_INST_1[54].FA_  ( .A(A[54]), .B(n972), .CI(C[54]), 
        .CO(C[55]) );
  FA_15623 \FA_INST_0[0].FA_INST_1[55].FA_  ( .A(A[55]), .B(n971), .CI(C[55]), 
        .CO(C[56]) );
  FA_15622 \FA_INST_0[0].FA_INST_1[56].FA_  ( .A(A[56]), .B(n970), .CI(C[56]), 
        .CO(C[57]) );
  FA_15621 \FA_INST_0[0].FA_INST_1[57].FA_  ( .A(A[57]), .B(n969), .CI(C[57]), 
        .CO(C[58]) );
  FA_15620 \FA_INST_0[0].FA_INST_1[58].FA_  ( .A(A[58]), .B(n968), .CI(C[58]), 
        .CO(C[59]) );
  FA_15619 \FA_INST_0[0].FA_INST_1[59].FA_  ( .A(A[59]), .B(n967), .CI(C[59]), 
        .CO(C[60]) );
  FA_15618 \FA_INST_0[0].FA_INST_1[60].FA_  ( .A(A[60]), .B(n966), .CI(C[60]), 
        .CO(C[61]) );
  FA_15617 \FA_INST_0[0].FA_INST_1[61].FA_  ( .A(A[61]), .B(n965), .CI(C[61]), 
        .CO(C[62]) );
  FA_15616 \FA_INST_0[0].FA_INST_1[62].FA_  ( .A(A[62]), .B(n964), .CI(C[62]), 
        .CO(C[63]) );
  FA_15615 \FA_INST_0[0].FA_INST_1[63].FA_  ( .A(A[63]), .B(n963), .CI(C[63]), 
        .CO(C[64]) );
  FA_15614 \FA_INST_0[0].FA_INST_1[64].FA_  ( .A(A[64]), .B(n962), .CI(C[64]), 
        .CO(C[65]) );
  FA_15613 \FA_INST_0[0].FA_INST_1[65].FA_  ( .A(A[65]), .B(n961), .CI(C[65]), 
        .CO(C[66]) );
  FA_15612 \FA_INST_0[0].FA_INST_1[66].FA_  ( .A(A[66]), .B(n960), .CI(C[66]), 
        .CO(C[67]) );
  FA_15611 \FA_INST_0[0].FA_INST_1[67].FA_  ( .A(A[67]), .B(n959), .CI(C[67]), 
        .CO(C[68]) );
  FA_15610 \FA_INST_0[0].FA_INST_1[68].FA_  ( .A(A[68]), .B(n958), .CI(C[68]), 
        .CO(C[69]) );
  FA_15609 \FA_INST_0[0].FA_INST_1[69].FA_  ( .A(A[69]), .B(n957), .CI(C[69]), 
        .CO(C[70]) );
  FA_15608 \FA_INST_0[0].FA_INST_1[70].FA_  ( .A(A[70]), .B(n956), .CI(C[70]), 
        .CO(C[71]) );
  FA_15607 \FA_INST_0[0].FA_INST_1[71].FA_  ( .A(A[71]), .B(n955), .CI(C[71]), 
        .CO(C[72]) );
  FA_15606 \FA_INST_0[0].FA_INST_1[72].FA_  ( .A(A[72]), .B(n954), .CI(C[72]), 
        .CO(C[73]) );
  FA_15605 \FA_INST_0[0].FA_INST_1[73].FA_  ( .A(A[73]), .B(n953), .CI(C[73]), 
        .CO(C[74]) );
  FA_15604 \FA_INST_0[0].FA_INST_1[74].FA_  ( .A(A[74]), .B(n952), .CI(C[74]), 
        .CO(C[75]) );
  FA_15603 \FA_INST_0[0].FA_INST_1[75].FA_  ( .A(A[75]), .B(n951), .CI(C[75]), 
        .CO(C[76]) );
  FA_15602 \FA_INST_0[0].FA_INST_1[76].FA_  ( .A(A[76]), .B(n950), .CI(C[76]), 
        .CO(C[77]) );
  FA_15601 \FA_INST_0[0].FA_INST_1[77].FA_  ( .A(A[77]), .B(n949), .CI(C[77]), 
        .CO(C[78]) );
  FA_15600 \FA_INST_0[0].FA_INST_1[78].FA_  ( .A(A[78]), .B(n948), .CI(C[78]), 
        .CO(C[79]) );
  FA_15599 \FA_INST_0[0].FA_INST_1[79].FA_  ( .A(A[79]), .B(n947), .CI(C[79]), 
        .CO(C[80]) );
  FA_15598 \FA_INST_0[0].FA_INST_1[80].FA_  ( .A(A[80]), .B(n946), .CI(C[80]), 
        .CO(C[81]) );
  FA_15597 \FA_INST_0[0].FA_INST_1[81].FA_  ( .A(A[81]), .B(n945), .CI(C[81]), 
        .CO(C[82]) );
  FA_15596 \FA_INST_0[0].FA_INST_1[82].FA_  ( .A(A[82]), .B(n944), .CI(C[82]), 
        .CO(C[83]) );
  FA_15595 \FA_INST_0[0].FA_INST_1[83].FA_  ( .A(A[83]), .B(n943), .CI(C[83]), 
        .CO(C[84]) );
  FA_15594 \FA_INST_0[0].FA_INST_1[84].FA_  ( .A(A[84]), .B(n942), .CI(C[84]), 
        .CO(C[85]) );
  FA_15593 \FA_INST_0[0].FA_INST_1[85].FA_  ( .A(A[85]), .B(n941), .CI(C[85]), 
        .CO(C[86]) );
  FA_15592 \FA_INST_0[0].FA_INST_1[86].FA_  ( .A(A[86]), .B(n940), .CI(C[86]), 
        .CO(C[87]) );
  FA_15591 \FA_INST_0[0].FA_INST_1[87].FA_  ( .A(A[87]), .B(n939), .CI(C[87]), 
        .CO(C[88]) );
  FA_15590 \FA_INST_0[0].FA_INST_1[88].FA_  ( .A(A[88]), .B(n938), .CI(C[88]), 
        .CO(C[89]) );
  FA_15589 \FA_INST_0[0].FA_INST_1[89].FA_  ( .A(A[89]), .B(n937), .CI(C[89]), 
        .CO(C[90]) );
  FA_15588 \FA_INST_0[0].FA_INST_1[90].FA_  ( .A(A[90]), .B(n936), .CI(C[90]), 
        .CO(C[91]) );
  FA_15587 \FA_INST_0[0].FA_INST_1[91].FA_  ( .A(A[91]), .B(n935), .CI(C[91]), 
        .CO(C[92]) );
  FA_15586 \FA_INST_0[0].FA_INST_1[92].FA_  ( .A(A[92]), .B(n934), .CI(C[92]), 
        .CO(C[93]) );
  FA_15585 \FA_INST_0[0].FA_INST_1[93].FA_  ( .A(A[93]), .B(n933), .CI(C[93]), 
        .CO(C[94]) );
  FA_15584 \FA_INST_0[0].FA_INST_1[94].FA_  ( .A(A[94]), .B(n932), .CI(C[94]), 
        .CO(C[95]) );
  FA_15583 \FA_INST_0[0].FA_INST_1[95].FA_  ( .A(A[95]), .B(n931), .CI(C[95]), 
        .CO(C[96]) );
  FA_15582 \FA_INST_0[0].FA_INST_1[96].FA_  ( .A(A[96]), .B(n930), .CI(C[96]), 
        .CO(C[97]) );
  FA_15581 \FA_INST_0[0].FA_INST_1[97].FA_  ( .A(A[97]), .B(n929), .CI(C[97]), 
        .CO(C[98]) );
  FA_15580 \FA_INST_0[0].FA_INST_1[98].FA_  ( .A(A[98]), .B(n928), .CI(C[98]), 
        .CO(C[99]) );
  FA_15579 \FA_INST_0[0].FA_INST_1[99].FA_  ( .A(A[99]), .B(n927), .CI(C[99]), 
        .CO(C[100]) );
  FA_15578 \FA_INST_0[0].FA_INST_1[100].FA_  ( .A(A[100]), .B(n926), .CI(
        C[100]), .CO(C[101]) );
  FA_15577 \FA_INST_0[0].FA_INST_1[101].FA_  ( .A(A[101]), .B(n925), .CI(
        C[101]), .CO(C[102]) );
  FA_15576 \FA_INST_0[0].FA_INST_1[102].FA_  ( .A(A[102]), .B(n924), .CI(
        C[102]), .CO(C[103]) );
  FA_15575 \FA_INST_0[0].FA_INST_1[103].FA_  ( .A(A[103]), .B(n923), .CI(
        C[103]), .CO(C[104]) );
  FA_15574 \FA_INST_0[0].FA_INST_1[104].FA_  ( .A(A[104]), .B(n922), .CI(
        C[104]), .CO(C[105]) );
  FA_15573 \FA_INST_0[0].FA_INST_1[105].FA_  ( .A(A[105]), .B(n921), .CI(
        C[105]), .CO(C[106]) );
  FA_15572 \FA_INST_0[0].FA_INST_1[106].FA_  ( .A(A[106]), .B(n920), .CI(
        C[106]), .CO(C[107]) );
  FA_15571 \FA_INST_0[0].FA_INST_1[107].FA_  ( .A(A[107]), .B(n919), .CI(
        C[107]), .CO(C[108]) );
  FA_15570 \FA_INST_0[0].FA_INST_1[108].FA_  ( .A(A[108]), .B(n918), .CI(
        C[108]), .CO(C[109]) );
  FA_15569 \FA_INST_0[0].FA_INST_1[109].FA_  ( .A(A[109]), .B(n917), .CI(
        C[109]), .CO(C[110]) );
  FA_15568 \FA_INST_0[0].FA_INST_1[110].FA_  ( .A(A[110]), .B(n916), .CI(
        C[110]), .CO(C[111]) );
  FA_15567 \FA_INST_0[0].FA_INST_1[111].FA_  ( .A(A[111]), .B(n915), .CI(
        C[111]), .CO(C[112]) );
  FA_15566 \FA_INST_0[0].FA_INST_1[112].FA_  ( .A(A[112]), .B(n914), .CI(
        C[112]), .CO(C[113]) );
  FA_15565 \FA_INST_0[0].FA_INST_1[113].FA_  ( .A(A[113]), .B(n913), .CI(
        C[113]), .CO(C[114]) );
  FA_15564 \FA_INST_0[0].FA_INST_1[114].FA_  ( .A(A[114]), .B(n912), .CI(
        C[114]), .CO(C[115]) );
  FA_15563 \FA_INST_0[0].FA_INST_1[115].FA_  ( .A(A[115]), .B(n911), .CI(
        C[115]), .CO(C[116]) );
  FA_15562 \FA_INST_0[0].FA_INST_1[116].FA_  ( .A(A[116]), .B(n910), .CI(
        C[116]), .CO(C[117]) );
  FA_15561 \FA_INST_0[0].FA_INST_1[117].FA_  ( .A(A[117]), .B(n909), .CI(
        C[117]), .CO(C[118]) );
  FA_15560 \FA_INST_0[0].FA_INST_1[118].FA_  ( .A(A[118]), .B(n908), .CI(
        C[118]), .CO(C[119]) );
  FA_15559 \FA_INST_0[0].FA_INST_1[119].FA_  ( .A(A[119]), .B(n907), .CI(
        C[119]), .CO(C[120]) );
  FA_15558 \FA_INST_0[0].FA_INST_1[120].FA_  ( .A(A[120]), .B(n906), .CI(
        C[120]), .CO(C[121]) );
  FA_15557 \FA_INST_0[0].FA_INST_1[121].FA_  ( .A(A[121]), .B(n905), .CI(
        C[121]), .CO(C[122]) );
  FA_15556 \FA_INST_0[0].FA_INST_1[122].FA_  ( .A(A[122]), .B(n904), .CI(
        C[122]), .CO(C[123]) );
  FA_15555 \FA_INST_0[0].FA_INST_1[123].FA_  ( .A(A[123]), .B(n903), .CI(
        C[123]), .CO(C[124]) );
  FA_15554 \FA_INST_0[0].FA_INST_1[124].FA_  ( .A(A[124]), .B(n902), .CI(
        C[124]), .CO(C[125]) );
  FA_15553 \FA_INST_0[0].FA_INST_1[125].FA_  ( .A(A[125]), .B(n901), .CI(
        C[125]), .CO(C[126]) );
  FA_15552 \FA_INST_0[0].FA_INST_1[126].FA_  ( .A(A[126]), .B(n900), .CI(
        C[126]), .CO(C[127]) );
  FA_15551 \FA_INST_0[0].FA_INST_1[127].FA_  ( .A(A[127]), .B(n899), .CI(
        C[127]), .CO(C[128]) );
  FA_15550 \FA_INST_0[0].FA_INST_1[128].FA_  ( .A(A[128]), .B(n898), .CI(
        C[128]), .CO(C[129]) );
  FA_15549 \FA_INST_0[0].FA_INST_1[129].FA_  ( .A(A[129]), .B(n897), .CI(
        C[129]), .CO(C[130]) );
  FA_15548 \FA_INST_0[0].FA_INST_1[130].FA_  ( .A(A[130]), .B(n896), .CI(
        C[130]), .CO(C[131]) );
  FA_15547 \FA_INST_0[0].FA_INST_1[131].FA_  ( .A(A[131]), .B(n895), .CI(
        C[131]), .CO(C[132]) );
  FA_15546 \FA_INST_0[0].FA_INST_1[132].FA_  ( .A(A[132]), .B(n894), .CI(
        C[132]), .CO(C[133]) );
  FA_15545 \FA_INST_0[0].FA_INST_1[133].FA_  ( .A(A[133]), .B(n893), .CI(
        C[133]), .CO(C[134]) );
  FA_15544 \FA_INST_0[0].FA_INST_1[134].FA_  ( .A(A[134]), .B(n892), .CI(
        C[134]), .CO(C[135]) );
  FA_15543 \FA_INST_0[0].FA_INST_1[135].FA_  ( .A(A[135]), .B(n891), .CI(
        C[135]), .CO(C[136]) );
  FA_15542 \FA_INST_0[0].FA_INST_1[136].FA_  ( .A(A[136]), .B(n890), .CI(
        C[136]), .CO(C[137]) );
  FA_15541 \FA_INST_0[0].FA_INST_1[137].FA_  ( .A(A[137]), .B(n889), .CI(
        C[137]), .CO(C[138]) );
  FA_15540 \FA_INST_0[0].FA_INST_1[138].FA_  ( .A(A[138]), .B(n888), .CI(
        C[138]), .CO(C[139]) );
  FA_15539 \FA_INST_0[0].FA_INST_1[139].FA_  ( .A(A[139]), .B(n887), .CI(
        C[139]), .CO(C[140]) );
  FA_15538 \FA_INST_0[0].FA_INST_1[140].FA_  ( .A(A[140]), .B(n886), .CI(
        C[140]), .CO(C[141]) );
  FA_15537 \FA_INST_0[0].FA_INST_1[141].FA_  ( .A(A[141]), .B(n885), .CI(
        C[141]), .CO(C[142]) );
  FA_15536 \FA_INST_0[0].FA_INST_1[142].FA_  ( .A(A[142]), .B(n884), .CI(
        C[142]), .CO(C[143]) );
  FA_15535 \FA_INST_0[0].FA_INST_1[143].FA_  ( .A(A[143]), .B(n883), .CI(
        C[143]), .CO(C[144]) );
  FA_15534 \FA_INST_0[0].FA_INST_1[144].FA_  ( .A(A[144]), .B(n882), .CI(
        C[144]), .CO(C[145]) );
  FA_15533 \FA_INST_0[0].FA_INST_1[145].FA_  ( .A(A[145]), .B(n881), .CI(
        C[145]), .CO(C[146]) );
  FA_15532 \FA_INST_0[0].FA_INST_1[146].FA_  ( .A(A[146]), .B(n880), .CI(
        C[146]), .CO(C[147]) );
  FA_15531 \FA_INST_0[0].FA_INST_1[147].FA_  ( .A(A[147]), .B(n879), .CI(
        C[147]), .CO(C[148]) );
  FA_15530 \FA_INST_0[0].FA_INST_1[148].FA_  ( .A(A[148]), .B(n878), .CI(
        C[148]), .CO(C[149]) );
  FA_15529 \FA_INST_0[0].FA_INST_1[149].FA_  ( .A(A[149]), .B(n877), .CI(
        C[149]), .CO(C[150]) );
  FA_15528 \FA_INST_0[0].FA_INST_1[150].FA_  ( .A(A[150]), .B(n876), .CI(
        C[150]), .CO(C[151]) );
  FA_15527 \FA_INST_0[0].FA_INST_1[151].FA_  ( .A(A[151]), .B(n875), .CI(
        C[151]), .CO(C[152]) );
  FA_15526 \FA_INST_0[0].FA_INST_1[152].FA_  ( .A(A[152]), .B(n874), .CI(
        C[152]), .CO(C[153]) );
  FA_15525 \FA_INST_0[0].FA_INST_1[153].FA_  ( .A(A[153]), .B(n873), .CI(
        C[153]), .CO(C[154]) );
  FA_15524 \FA_INST_0[0].FA_INST_1[154].FA_  ( .A(A[154]), .B(n872), .CI(
        C[154]), .CO(C[155]) );
  FA_15523 \FA_INST_0[0].FA_INST_1[155].FA_  ( .A(A[155]), .B(n871), .CI(
        C[155]), .CO(C[156]) );
  FA_15522 \FA_INST_0[0].FA_INST_1[156].FA_  ( .A(A[156]), .B(n870), .CI(
        C[156]), .CO(C[157]) );
  FA_15521 \FA_INST_0[0].FA_INST_1[157].FA_  ( .A(A[157]), .B(n869), .CI(
        C[157]), .CO(C[158]) );
  FA_15520 \FA_INST_0[0].FA_INST_1[158].FA_  ( .A(A[158]), .B(n868), .CI(
        C[158]), .CO(C[159]) );
  FA_15519 \FA_INST_0[0].FA_INST_1[159].FA_  ( .A(A[159]), .B(n867), .CI(
        C[159]), .CO(C[160]) );
  FA_15518 \FA_INST_0[0].FA_INST_1[160].FA_  ( .A(A[160]), .B(n866), .CI(
        C[160]), .CO(C[161]) );
  FA_15517 \FA_INST_0[0].FA_INST_1[161].FA_  ( .A(A[161]), .B(n865), .CI(
        C[161]), .CO(C[162]) );
  FA_15516 \FA_INST_0[0].FA_INST_1[162].FA_  ( .A(A[162]), .B(n864), .CI(
        C[162]), .CO(C[163]) );
  FA_15515 \FA_INST_0[0].FA_INST_1[163].FA_  ( .A(A[163]), .B(n863), .CI(
        C[163]), .CO(C[164]) );
  FA_15514 \FA_INST_0[0].FA_INST_1[164].FA_  ( .A(A[164]), .B(n862), .CI(
        C[164]), .CO(C[165]) );
  FA_15513 \FA_INST_0[0].FA_INST_1[165].FA_  ( .A(A[165]), .B(n861), .CI(
        C[165]), .CO(C[166]) );
  FA_15512 \FA_INST_0[0].FA_INST_1[166].FA_  ( .A(A[166]), .B(n860), .CI(
        C[166]), .CO(C[167]) );
  FA_15511 \FA_INST_0[0].FA_INST_1[167].FA_  ( .A(A[167]), .B(n859), .CI(
        C[167]), .CO(C[168]) );
  FA_15510 \FA_INST_0[0].FA_INST_1[168].FA_  ( .A(A[168]), .B(n858), .CI(
        C[168]), .CO(C[169]) );
  FA_15509 \FA_INST_0[0].FA_INST_1[169].FA_  ( .A(A[169]), .B(n857), .CI(
        C[169]), .CO(C[170]) );
  FA_15508 \FA_INST_0[0].FA_INST_1[170].FA_  ( .A(A[170]), .B(n856), .CI(
        C[170]), .CO(C[171]) );
  FA_15507 \FA_INST_0[0].FA_INST_1[171].FA_  ( .A(A[171]), .B(n855), .CI(
        C[171]), .CO(C[172]) );
  FA_15506 \FA_INST_0[0].FA_INST_1[172].FA_  ( .A(A[172]), .B(n854), .CI(
        C[172]), .CO(C[173]) );
  FA_15505 \FA_INST_0[0].FA_INST_1[173].FA_  ( .A(A[173]), .B(n853), .CI(
        C[173]), .CO(C[174]) );
  FA_15504 \FA_INST_0[0].FA_INST_1[174].FA_  ( .A(A[174]), .B(n852), .CI(
        C[174]), .CO(C[175]) );
  FA_15503 \FA_INST_0[0].FA_INST_1[175].FA_  ( .A(A[175]), .B(n851), .CI(
        C[175]), .CO(C[176]) );
  FA_15502 \FA_INST_0[0].FA_INST_1[176].FA_  ( .A(A[176]), .B(n850), .CI(
        C[176]), .CO(C[177]) );
  FA_15501 \FA_INST_0[0].FA_INST_1[177].FA_  ( .A(A[177]), .B(n849), .CI(
        C[177]), .CO(C[178]) );
  FA_15500 \FA_INST_0[0].FA_INST_1[178].FA_  ( .A(A[178]), .B(n848), .CI(
        C[178]), .CO(C[179]) );
  FA_15499 \FA_INST_0[0].FA_INST_1[179].FA_  ( .A(A[179]), .B(n847), .CI(
        C[179]), .CO(C[180]) );
  FA_15498 \FA_INST_0[0].FA_INST_1[180].FA_  ( .A(A[180]), .B(n846), .CI(
        C[180]), .CO(C[181]) );
  FA_15497 \FA_INST_0[0].FA_INST_1[181].FA_  ( .A(A[181]), .B(n845), .CI(
        C[181]), .CO(C[182]) );
  FA_15496 \FA_INST_0[0].FA_INST_1[182].FA_  ( .A(A[182]), .B(n844), .CI(
        C[182]), .CO(C[183]) );
  FA_15495 \FA_INST_0[0].FA_INST_1[183].FA_  ( .A(A[183]), .B(n843), .CI(
        C[183]), .CO(C[184]) );
  FA_15494 \FA_INST_0[0].FA_INST_1[184].FA_  ( .A(A[184]), .B(n842), .CI(
        C[184]), .CO(C[185]) );
  FA_15493 \FA_INST_0[0].FA_INST_1[185].FA_  ( .A(A[185]), .B(n841), .CI(
        C[185]), .CO(C[186]) );
  FA_15492 \FA_INST_0[0].FA_INST_1[186].FA_  ( .A(A[186]), .B(n840), .CI(
        C[186]), .CO(C[187]) );
  FA_15491 \FA_INST_0[0].FA_INST_1[187].FA_  ( .A(A[187]), .B(n839), .CI(
        C[187]), .CO(C[188]) );
  FA_15490 \FA_INST_0[0].FA_INST_1[188].FA_  ( .A(A[188]), .B(n838), .CI(
        C[188]), .CO(C[189]) );
  FA_15489 \FA_INST_0[0].FA_INST_1[189].FA_  ( .A(A[189]), .B(n837), .CI(
        C[189]), .CO(C[190]) );
  FA_15488 \FA_INST_0[0].FA_INST_1[190].FA_  ( .A(A[190]), .B(n836), .CI(
        C[190]), .CO(C[191]) );
  FA_15487 \FA_INST_0[0].FA_INST_1[191].FA_  ( .A(A[191]), .B(n835), .CI(
        C[191]), .CO(C[192]) );
  FA_15486 \FA_INST_0[0].FA_INST_1[192].FA_  ( .A(A[192]), .B(n834), .CI(
        C[192]), .CO(C[193]) );
  FA_15485 \FA_INST_0[0].FA_INST_1[193].FA_  ( .A(A[193]), .B(n833), .CI(
        C[193]), .CO(C[194]) );
  FA_15484 \FA_INST_0[0].FA_INST_1[194].FA_  ( .A(A[194]), .B(n832), .CI(
        C[194]), .CO(C[195]) );
  FA_15483 \FA_INST_0[0].FA_INST_1[195].FA_  ( .A(A[195]), .B(n831), .CI(
        C[195]), .CO(C[196]) );
  FA_15482 \FA_INST_0[0].FA_INST_1[196].FA_  ( .A(A[196]), .B(n830), .CI(
        C[196]), .CO(C[197]) );
  FA_15481 \FA_INST_0[0].FA_INST_1[197].FA_  ( .A(A[197]), .B(n829), .CI(
        C[197]), .CO(C[198]) );
  FA_15480 \FA_INST_0[0].FA_INST_1[198].FA_  ( .A(A[198]), .B(n828), .CI(
        C[198]), .CO(C[199]) );
  FA_15479 \FA_INST_0[0].FA_INST_1[199].FA_  ( .A(A[199]), .B(n827), .CI(
        C[199]), .CO(C[200]) );
  FA_15478 \FA_INST_0[0].FA_INST_1[200].FA_  ( .A(A[200]), .B(n826), .CI(
        C[200]), .CO(C[201]) );
  FA_15477 \FA_INST_0[0].FA_INST_1[201].FA_  ( .A(A[201]), .B(n825), .CI(
        C[201]), .CO(C[202]) );
  FA_15476 \FA_INST_0[0].FA_INST_1[202].FA_  ( .A(A[202]), .B(n824), .CI(
        C[202]), .CO(C[203]) );
  FA_15475 \FA_INST_0[0].FA_INST_1[203].FA_  ( .A(A[203]), .B(n823), .CI(
        C[203]), .CO(C[204]) );
  FA_15474 \FA_INST_0[0].FA_INST_1[204].FA_  ( .A(A[204]), .B(n822), .CI(
        C[204]), .CO(C[205]) );
  FA_15473 \FA_INST_0[0].FA_INST_1[205].FA_  ( .A(A[205]), .B(n821), .CI(
        C[205]), .CO(C[206]) );
  FA_15472 \FA_INST_0[0].FA_INST_1[206].FA_  ( .A(A[206]), .B(n820), .CI(
        C[206]), .CO(C[207]) );
  FA_15471 \FA_INST_0[0].FA_INST_1[207].FA_  ( .A(A[207]), .B(n819), .CI(
        C[207]), .CO(C[208]) );
  FA_15470 \FA_INST_0[0].FA_INST_1[208].FA_  ( .A(A[208]), .B(n818), .CI(
        C[208]), .CO(C[209]) );
  FA_15469 \FA_INST_0[0].FA_INST_1[209].FA_  ( .A(A[209]), .B(n817), .CI(
        C[209]), .CO(C[210]) );
  FA_15468 \FA_INST_0[0].FA_INST_1[210].FA_  ( .A(A[210]), .B(n816), .CI(
        C[210]), .CO(C[211]) );
  FA_15467 \FA_INST_0[0].FA_INST_1[211].FA_  ( .A(A[211]), .B(n815), .CI(
        C[211]), .CO(C[212]) );
  FA_15466 \FA_INST_0[0].FA_INST_1[212].FA_  ( .A(A[212]), .B(n814), .CI(
        C[212]), .CO(C[213]) );
  FA_15465 \FA_INST_0[0].FA_INST_1[213].FA_  ( .A(A[213]), .B(n813), .CI(
        C[213]), .CO(C[214]) );
  FA_15464 \FA_INST_0[0].FA_INST_1[214].FA_  ( .A(A[214]), .B(n812), .CI(
        C[214]), .CO(C[215]) );
  FA_15463 \FA_INST_0[0].FA_INST_1[215].FA_  ( .A(A[215]), .B(n811), .CI(
        C[215]), .CO(C[216]) );
  FA_15462 \FA_INST_0[0].FA_INST_1[216].FA_  ( .A(A[216]), .B(n810), .CI(
        C[216]), .CO(C[217]) );
  FA_15461 \FA_INST_0[0].FA_INST_1[217].FA_  ( .A(A[217]), .B(n809), .CI(
        C[217]), .CO(C[218]) );
  FA_15460 \FA_INST_0[0].FA_INST_1[218].FA_  ( .A(A[218]), .B(n808), .CI(
        C[218]), .CO(C[219]) );
  FA_15459 \FA_INST_0[0].FA_INST_1[219].FA_  ( .A(A[219]), .B(n807), .CI(
        C[219]), .CO(C[220]) );
  FA_15458 \FA_INST_0[0].FA_INST_1[220].FA_  ( .A(A[220]), .B(n806), .CI(
        C[220]), .CO(C[221]) );
  FA_15457 \FA_INST_0[0].FA_INST_1[221].FA_  ( .A(A[221]), .B(n805), .CI(
        C[221]), .CO(C[222]) );
  FA_15456 \FA_INST_0[0].FA_INST_1[222].FA_  ( .A(A[222]), .B(n804), .CI(
        C[222]), .CO(C[223]) );
  FA_15455 \FA_INST_0[0].FA_INST_1[223].FA_  ( .A(A[223]), .B(n803), .CI(
        C[223]), .CO(C[224]) );
  FA_15454 \FA_INST_0[0].FA_INST_1[224].FA_  ( .A(A[224]), .B(n802), .CI(
        C[224]), .CO(C[225]) );
  FA_15453 \FA_INST_0[0].FA_INST_1[225].FA_  ( .A(A[225]), .B(n801), .CI(
        C[225]), .CO(C[226]) );
  FA_15452 \FA_INST_0[0].FA_INST_1[226].FA_  ( .A(A[226]), .B(n800), .CI(
        C[226]), .CO(C[227]) );
  FA_15451 \FA_INST_0[0].FA_INST_1[227].FA_  ( .A(A[227]), .B(n799), .CI(
        C[227]), .CO(C[228]) );
  FA_15450 \FA_INST_0[0].FA_INST_1[228].FA_  ( .A(A[228]), .B(n798), .CI(
        C[228]), .CO(C[229]) );
  FA_15449 \FA_INST_0[0].FA_INST_1[229].FA_  ( .A(A[229]), .B(n797), .CI(
        C[229]), .CO(C[230]) );
  FA_15448 \FA_INST_0[0].FA_INST_1[230].FA_  ( .A(A[230]), .B(n796), .CI(
        C[230]), .CO(C[231]) );
  FA_15447 \FA_INST_0[0].FA_INST_1[231].FA_  ( .A(A[231]), .B(n795), .CI(
        C[231]), .CO(C[232]) );
  FA_15446 \FA_INST_0[0].FA_INST_1[232].FA_  ( .A(A[232]), .B(n794), .CI(
        C[232]), .CO(C[233]) );
  FA_15445 \FA_INST_0[0].FA_INST_1[233].FA_  ( .A(A[233]), .B(n793), .CI(
        C[233]), .CO(C[234]) );
  FA_15444 \FA_INST_0[0].FA_INST_1[234].FA_  ( .A(A[234]), .B(n792), .CI(
        C[234]), .CO(C[235]) );
  FA_15443 \FA_INST_0[0].FA_INST_1[235].FA_  ( .A(A[235]), .B(n791), .CI(
        C[235]), .CO(C[236]) );
  FA_15442 \FA_INST_0[0].FA_INST_1[236].FA_  ( .A(A[236]), .B(n790), .CI(
        C[236]), .CO(C[237]) );
  FA_15441 \FA_INST_0[0].FA_INST_1[237].FA_  ( .A(A[237]), .B(n789), .CI(
        C[237]), .CO(C[238]) );
  FA_15440 \FA_INST_0[0].FA_INST_1[238].FA_  ( .A(A[238]), .B(n788), .CI(
        C[238]), .CO(C[239]) );
  FA_15439 \FA_INST_0[0].FA_INST_1[239].FA_  ( .A(A[239]), .B(n787), .CI(
        C[239]), .CO(C[240]) );
  FA_15438 \FA_INST_0[0].FA_INST_1[240].FA_  ( .A(A[240]), .B(n786), .CI(
        C[240]), .CO(C[241]) );
  FA_15437 \FA_INST_0[0].FA_INST_1[241].FA_  ( .A(A[241]), .B(n785), .CI(
        C[241]), .CO(C[242]) );
  FA_15436 \FA_INST_0[0].FA_INST_1[242].FA_  ( .A(A[242]), .B(n784), .CI(
        C[242]), .CO(C[243]) );
  FA_15435 \FA_INST_0[0].FA_INST_1[243].FA_  ( .A(A[243]), .B(n783), .CI(
        C[243]), .CO(C[244]) );
  FA_15434 \FA_INST_0[0].FA_INST_1[244].FA_  ( .A(A[244]), .B(n782), .CI(
        C[244]), .CO(C[245]) );
  FA_15433 \FA_INST_0[0].FA_INST_1[245].FA_  ( .A(A[245]), .B(n781), .CI(
        C[245]), .CO(C[246]) );
  FA_15432 \FA_INST_0[0].FA_INST_1[246].FA_  ( .A(A[246]), .B(n780), .CI(
        C[246]), .CO(C[247]) );
  FA_15431 \FA_INST_0[0].FA_INST_1[247].FA_  ( .A(A[247]), .B(n779), .CI(
        C[247]), .CO(C[248]) );
  FA_15430 \FA_INST_0[0].FA_INST_1[248].FA_  ( .A(A[248]), .B(n778), .CI(
        C[248]), .CO(C[249]) );
  FA_15429 \FA_INST_0[0].FA_INST_1[249].FA_  ( .A(A[249]), .B(n777), .CI(
        C[249]), .CO(C[250]) );
  FA_15428 \FA_INST_0[0].FA_INST_1[250].FA_  ( .A(A[250]), .B(n776), .CI(
        C[250]), .CO(C[251]) );
  FA_15427 \FA_INST_0[0].FA_INST_1[251].FA_  ( .A(A[251]), .B(n775), .CI(
        C[251]), .CO(C[252]) );
  FA_15426 \FA_INST_0[0].FA_INST_1[252].FA_  ( .A(A[252]), .B(n774), .CI(
        C[252]), .CO(C[253]) );
  FA_15425 \FA_INST_0[0].FA_INST_1[253].FA_  ( .A(A[253]), .B(n773), .CI(
        C[253]), .CO(C[254]) );
  FA_15424 \FA_INST_0[0].FA_INST_1[254].FA_  ( .A(A[254]), .B(n772), .CI(
        C[254]), .CO(C[255]) );
  FA_15423 \FA_INST_0[0].FA_INST_1[255].FA_  ( .A(A[255]), .B(n771), .CI(
        C[255]), .CO(C[256]) );
  FA_15422 \FA_INST_0[0].FA_INST_1[256].FA_  ( .A(A[256]), .B(n770), .CI(
        C[256]), .CO(C[257]) );
  FA_15421 \FA_INST_0[0].FA_INST_1[257].FA_  ( .A(A[257]), .B(n769), .CI(
        C[257]), .CO(C[258]) );
  FA_15420 \FA_INST_0[0].FA_INST_1[258].FA_  ( .A(A[258]), .B(n768), .CI(
        C[258]), .CO(C[259]) );
  FA_15419 \FA_INST_0[0].FA_INST_1[259].FA_  ( .A(A[259]), .B(n767), .CI(
        C[259]), .CO(C[260]) );
  FA_15418 \FA_INST_0[0].FA_INST_1[260].FA_  ( .A(A[260]), .B(n766), .CI(
        C[260]), .CO(C[261]) );
  FA_15417 \FA_INST_0[0].FA_INST_1[261].FA_  ( .A(A[261]), .B(n765), .CI(
        C[261]), .CO(C[262]) );
  FA_15416 \FA_INST_0[0].FA_INST_1[262].FA_  ( .A(A[262]), .B(n764), .CI(
        C[262]), .CO(C[263]) );
  FA_15415 \FA_INST_0[0].FA_INST_1[263].FA_  ( .A(A[263]), .B(n763), .CI(
        C[263]), .CO(C[264]) );
  FA_15414 \FA_INST_0[0].FA_INST_1[264].FA_  ( .A(A[264]), .B(n762), .CI(
        C[264]), .CO(C[265]) );
  FA_15413 \FA_INST_0[0].FA_INST_1[265].FA_  ( .A(A[265]), .B(n761), .CI(
        C[265]), .CO(C[266]) );
  FA_15412 \FA_INST_0[0].FA_INST_1[266].FA_  ( .A(A[266]), .B(n760), .CI(
        C[266]), .CO(C[267]) );
  FA_15411 \FA_INST_0[0].FA_INST_1[267].FA_  ( .A(A[267]), .B(n759), .CI(
        C[267]), .CO(C[268]) );
  FA_15410 \FA_INST_0[0].FA_INST_1[268].FA_  ( .A(A[268]), .B(n758), .CI(
        C[268]), .CO(C[269]) );
  FA_15409 \FA_INST_0[0].FA_INST_1[269].FA_  ( .A(A[269]), .B(n757), .CI(
        C[269]), .CO(C[270]) );
  FA_15408 \FA_INST_0[0].FA_INST_1[270].FA_  ( .A(A[270]), .B(n756), .CI(
        C[270]), .CO(C[271]) );
  FA_15407 \FA_INST_0[0].FA_INST_1[271].FA_  ( .A(A[271]), .B(n755), .CI(
        C[271]), .CO(C[272]) );
  FA_15406 \FA_INST_0[0].FA_INST_1[272].FA_  ( .A(A[272]), .B(n754), .CI(
        C[272]), .CO(C[273]) );
  FA_15405 \FA_INST_0[0].FA_INST_1[273].FA_  ( .A(A[273]), .B(n753), .CI(
        C[273]), .CO(C[274]) );
  FA_15404 \FA_INST_0[0].FA_INST_1[274].FA_  ( .A(A[274]), .B(n752), .CI(
        C[274]), .CO(C[275]) );
  FA_15403 \FA_INST_0[0].FA_INST_1[275].FA_  ( .A(A[275]), .B(n751), .CI(
        C[275]), .CO(C[276]) );
  FA_15402 \FA_INST_0[0].FA_INST_1[276].FA_  ( .A(A[276]), .B(n750), .CI(
        C[276]), .CO(C[277]) );
  FA_15401 \FA_INST_0[0].FA_INST_1[277].FA_  ( .A(A[277]), .B(n749), .CI(
        C[277]), .CO(C[278]) );
  FA_15400 \FA_INST_0[0].FA_INST_1[278].FA_  ( .A(A[278]), .B(n748), .CI(
        C[278]), .CO(C[279]) );
  FA_15399 \FA_INST_0[0].FA_INST_1[279].FA_  ( .A(A[279]), .B(n747), .CI(
        C[279]), .CO(C[280]) );
  FA_15398 \FA_INST_0[0].FA_INST_1[280].FA_  ( .A(A[280]), .B(n746), .CI(
        C[280]), .CO(C[281]) );
  FA_15397 \FA_INST_0[0].FA_INST_1[281].FA_  ( .A(A[281]), .B(n745), .CI(
        C[281]), .CO(C[282]) );
  FA_15396 \FA_INST_0[0].FA_INST_1[282].FA_  ( .A(A[282]), .B(n744), .CI(
        C[282]), .CO(C[283]) );
  FA_15395 \FA_INST_0[0].FA_INST_1[283].FA_  ( .A(A[283]), .B(n743), .CI(
        C[283]), .CO(C[284]) );
  FA_15394 \FA_INST_0[0].FA_INST_1[284].FA_  ( .A(A[284]), .B(n742), .CI(
        C[284]), .CO(C[285]) );
  FA_15393 \FA_INST_0[0].FA_INST_1[285].FA_  ( .A(A[285]), .B(n741), .CI(
        C[285]), .CO(C[286]) );
  FA_15392 \FA_INST_0[0].FA_INST_1[286].FA_  ( .A(A[286]), .B(n740), .CI(
        C[286]), .CO(C[287]) );
  FA_15391 \FA_INST_0[0].FA_INST_1[287].FA_  ( .A(A[287]), .B(n739), .CI(
        C[287]), .CO(C[288]) );
  FA_15390 \FA_INST_0[0].FA_INST_1[288].FA_  ( .A(A[288]), .B(n738), .CI(
        C[288]), .CO(C[289]) );
  FA_15389 \FA_INST_0[0].FA_INST_1[289].FA_  ( .A(A[289]), .B(n737), .CI(
        C[289]), .CO(C[290]) );
  FA_15388 \FA_INST_0[0].FA_INST_1[290].FA_  ( .A(A[290]), .B(n736), .CI(
        C[290]), .CO(C[291]) );
  FA_15387 \FA_INST_0[0].FA_INST_1[291].FA_  ( .A(A[291]), .B(n735), .CI(
        C[291]), .CO(C[292]) );
  FA_15386 \FA_INST_0[0].FA_INST_1[292].FA_  ( .A(A[292]), .B(n734), .CI(
        C[292]), .CO(C[293]) );
  FA_15385 \FA_INST_0[0].FA_INST_1[293].FA_  ( .A(A[293]), .B(n733), .CI(
        C[293]), .CO(C[294]) );
  FA_15384 \FA_INST_0[0].FA_INST_1[294].FA_  ( .A(A[294]), .B(n732), .CI(
        C[294]), .CO(C[295]) );
  FA_15383 \FA_INST_0[0].FA_INST_1[295].FA_  ( .A(A[295]), .B(n731), .CI(
        C[295]), .CO(C[296]) );
  FA_15382 \FA_INST_0[0].FA_INST_1[296].FA_  ( .A(A[296]), .B(n730), .CI(
        C[296]), .CO(C[297]) );
  FA_15381 \FA_INST_0[0].FA_INST_1[297].FA_  ( .A(A[297]), .B(n729), .CI(
        C[297]), .CO(C[298]) );
  FA_15380 \FA_INST_0[0].FA_INST_1[298].FA_  ( .A(A[298]), .B(n728), .CI(
        C[298]), .CO(C[299]) );
  FA_15379 \FA_INST_0[0].FA_INST_1[299].FA_  ( .A(A[299]), .B(n727), .CI(
        C[299]), .CO(C[300]) );
  FA_15378 \FA_INST_0[0].FA_INST_1[300].FA_  ( .A(A[300]), .B(n726), .CI(
        C[300]), .CO(C[301]) );
  FA_15377 \FA_INST_0[0].FA_INST_1[301].FA_  ( .A(A[301]), .B(n725), .CI(
        C[301]), .CO(C[302]) );
  FA_15376 \FA_INST_0[0].FA_INST_1[302].FA_  ( .A(A[302]), .B(n724), .CI(
        C[302]), .CO(C[303]) );
  FA_15375 \FA_INST_0[0].FA_INST_1[303].FA_  ( .A(A[303]), .B(n723), .CI(
        C[303]), .CO(C[304]) );
  FA_15374 \FA_INST_0[0].FA_INST_1[304].FA_  ( .A(A[304]), .B(n722), .CI(
        C[304]), .CO(C[305]) );
  FA_15373 \FA_INST_0[0].FA_INST_1[305].FA_  ( .A(A[305]), .B(n721), .CI(
        C[305]), .CO(C[306]) );
  FA_15372 \FA_INST_0[0].FA_INST_1[306].FA_  ( .A(A[306]), .B(n720), .CI(
        C[306]), .CO(C[307]) );
  FA_15371 \FA_INST_0[0].FA_INST_1[307].FA_  ( .A(A[307]), .B(n719), .CI(
        C[307]), .CO(C[308]) );
  FA_15370 \FA_INST_0[0].FA_INST_1[308].FA_  ( .A(A[308]), .B(n718), .CI(
        C[308]), .CO(C[309]) );
  FA_15369 \FA_INST_0[0].FA_INST_1[309].FA_  ( .A(A[309]), .B(n717), .CI(
        C[309]), .CO(C[310]) );
  FA_15368 \FA_INST_0[0].FA_INST_1[310].FA_  ( .A(A[310]), .B(n716), .CI(
        C[310]), .CO(C[311]) );
  FA_15367 \FA_INST_0[0].FA_INST_1[311].FA_  ( .A(A[311]), .B(n715), .CI(
        C[311]), .CO(C[312]) );
  FA_15366 \FA_INST_0[0].FA_INST_1[312].FA_  ( .A(A[312]), .B(n714), .CI(
        C[312]), .CO(C[313]) );
  FA_15365 \FA_INST_0[0].FA_INST_1[313].FA_  ( .A(A[313]), .B(n713), .CI(
        C[313]), .CO(C[314]) );
  FA_15364 \FA_INST_0[0].FA_INST_1[314].FA_  ( .A(A[314]), .B(n712), .CI(
        C[314]), .CO(C[315]) );
  FA_15363 \FA_INST_0[0].FA_INST_1[315].FA_  ( .A(A[315]), .B(n711), .CI(
        C[315]), .CO(C[316]) );
  FA_15362 \FA_INST_0[0].FA_INST_1[316].FA_  ( .A(A[316]), .B(n710), .CI(
        C[316]), .CO(C[317]) );
  FA_15361 \FA_INST_0[0].FA_INST_1[317].FA_  ( .A(A[317]), .B(n709), .CI(
        C[317]), .CO(C[318]) );
  FA_15360 \FA_INST_0[0].FA_INST_1[318].FA_  ( .A(A[318]), .B(n708), .CI(
        C[318]), .CO(C[319]) );
  FA_15359 \FA_INST_0[0].FA_INST_1[319].FA_  ( .A(A[319]), .B(n707), .CI(
        C[319]), .CO(C[320]) );
  FA_15358 \FA_INST_0[0].FA_INST_1[320].FA_  ( .A(A[320]), .B(n706), .CI(
        C[320]), .CO(C[321]) );
  FA_15357 \FA_INST_0[0].FA_INST_1[321].FA_  ( .A(A[321]), .B(n705), .CI(
        C[321]), .CO(C[322]) );
  FA_15356 \FA_INST_0[0].FA_INST_1[322].FA_  ( .A(A[322]), .B(n704), .CI(
        C[322]), .CO(C[323]) );
  FA_15355 \FA_INST_0[0].FA_INST_1[323].FA_  ( .A(A[323]), .B(n703), .CI(
        C[323]), .CO(C[324]) );
  FA_15354 \FA_INST_0[0].FA_INST_1[324].FA_  ( .A(A[324]), .B(n702), .CI(
        C[324]), .CO(C[325]) );
  FA_15353 \FA_INST_0[0].FA_INST_1[325].FA_  ( .A(A[325]), .B(n701), .CI(
        C[325]), .CO(C[326]) );
  FA_15352 \FA_INST_0[0].FA_INST_1[326].FA_  ( .A(A[326]), .B(n700), .CI(
        C[326]), .CO(C[327]) );
  FA_15351 \FA_INST_0[0].FA_INST_1[327].FA_  ( .A(A[327]), .B(n699), .CI(
        C[327]), .CO(C[328]) );
  FA_15350 \FA_INST_0[0].FA_INST_1[328].FA_  ( .A(A[328]), .B(n698), .CI(
        C[328]), .CO(C[329]) );
  FA_15349 \FA_INST_0[0].FA_INST_1[329].FA_  ( .A(A[329]), .B(n697), .CI(
        C[329]), .CO(C[330]) );
  FA_15348 \FA_INST_0[0].FA_INST_1[330].FA_  ( .A(A[330]), .B(n696), .CI(
        C[330]), .CO(C[331]) );
  FA_15347 \FA_INST_0[0].FA_INST_1[331].FA_  ( .A(A[331]), .B(n695), .CI(
        C[331]), .CO(C[332]) );
  FA_15346 \FA_INST_0[0].FA_INST_1[332].FA_  ( .A(A[332]), .B(n694), .CI(
        C[332]), .CO(C[333]) );
  FA_15345 \FA_INST_0[0].FA_INST_1[333].FA_  ( .A(A[333]), .B(n693), .CI(
        C[333]), .CO(C[334]) );
  FA_15344 \FA_INST_0[0].FA_INST_1[334].FA_  ( .A(A[334]), .B(n692), .CI(
        C[334]), .CO(C[335]) );
  FA_15343 \FA_INST_0[0].FA_INST_1[335].FA_  ( .A(A[335]), .B(n691), .CI(
        C[335]), .CO(C[336]) );
  FA_15342 \FA_INST_0[0].FA_INST_1[336].FA_  ( .A(A[336]), .B(n690), .CI(
        C[336]), .CO(C[337]) );
  FA_15341 \FA_INST_0[0].FA_INST_1[337].FA_  ( .A(A[337]), .B(n689), .CI(
        C[337]), .CO(C[338]) );
  FA_15340 \FA_INST_0[0].FA_INST_1[338].FA_  ( .A(A[338]), .B(n688), .CI(
        C[338]), .CO(C[339]) );
  FA_15339 \FA_INST_0[0].FA_INST_1[339].FA_  ( .A(A[339]), .B(n687), .CI(
        C[339]), .CO(C[340]) );
  FA_15338 \FA_INST_0[0].FA_INST_1[340].FA_  ( .A(A[340]), .B(n686), .CI(
        C[340]), .CO(C[341]) );
  FA_15337 \FA_INST_0[0].FA_INST_1[341].FA_  ( .A(A[341]), .B(n685), .CI(
        C[341]), .CO(C[342]) );
  FA_15336 \FA_INST_0[0].FA_INST_1[342].FA_  ( .A(A[342]), .B(n684), .CI(
        C[342]), .CO(C[343]) );
  FA_15335 \FA_INST_0[0].FA_INST_1[343].FA_  ( .A(A[343]), .B(n683), .CI(
        C[343]), .CO(C[344]) );
  FA_15334 \FA_INST_0[0].FA_INST_1[344].FA_  ( .A(A[344]), .B(n682), .CI(
        C[344]), .CO(C[345]) );
  FA_15333 \FA_INST_0[0].FA_INST_1[345].FA_  ( .A(A[345]), .B(n681), .CI(
        C[345]), .CO(C[346]) );
  FA_15332 \FA_INST_0[0].FA_INST_1[346].FA_  ( .A(A[346]), .B(n680), .CI(
        C[346]), .CO(C[347]) );
  FA_15331 \FA_INST_0[0].FA_INST_1[347].FA_  ( .A(A[347]), .B(n679), .CI(
        C[347]), .CO(C[348]) );
  FA_15330 \FA_INST_0[0].FA_INST_1[348].FA_  ( .A(A[348]), .B(n678), .CI(
        C[348]), .CO(C[349]) );
  FA_15329 \FA_INST_0[0].FA_INST_1[349].FA_  ( .A(A[349]), .B(n677), .CI(
        C[349]), .CO(C[350]) );
  FA_15328 \FA_INST_0[0].FA_INST_1[350].FA_  ( .A(A[350]), .B(n676), .CI(
        C[350]), .CO(C[351]) );
  FA_15327 \FA_INST_0[0].FA_INST_1[351].FA_  ( .A(A[351]), .B(n675), .CI(
        C[351]), .CO(C[352]) );
  FA_15326 \FA_INST_0[0].FA_INST_1[352].FA_  ( .A(A[352]), .B(n674), .CI(
        C[352]), .CO(C[353]) );
  FA_15325 \FA_INST_0[0].FA_INST_1[353].FA_  ( .A(A[353]), .B(n673), .CI(
        C[353]), .CO(C[354]) );
  FA_15324 \FA_INST_0[0].FA_INST_1[354].FA_  ( .A(A[354]), .B(n672), .CI(
        C[354]), .CO(C[355]) );
  FA_15323 \FA_INST_0[0].FA_INST_1[355].FA_  ( .A(A[355]), .B(n671), .CI(
        C[355]), .CO(C[356]) );
  FA_15322 \FA_INST_0[0].FA_INST_1[356].FA_  ( .A(A[356]), .B(n670), .CI(
        C[356]), .CO(C[357]) );
  FA_15321 \FA_INST_0[0].FA_INST_1[357].FA_  ( .A(A[357]), .B(n669), .CI(
        C[357]), .CO(C[358]) );
  FA_15320 \FA_INST_0[0].FA_INST_1[358].FA_  ( .A(A[358]), .B(n668), .CI(
        C[358]), .CO(C[359]) );
  FA_15319 \FA_INST_0[0].FA_INST_1[359].FA_  ( .A(A[359]), .B(n667), .CI(
        C[359]), .CO(C[360]) );
  FA_15318 \FA_INST_0[0].FA_INST_1[360].FA_  ( .A(A[360]), .B(n666), .CI(
        C[360]), .CO(C[361]) );
  FA_15317 \FA_INST_0[0].FA_INST_1[361].FA_  ( .A(A[361]), .B(n665), .CI(
        C[361]), .CO(C[362]) );
  FA_15316 \FA_INST_0[0].FA_INST_1[362].FA_  ( .A(A[362]), .B(n664), .CI(
        C[362]), .CO(C[363]) );
  FA_15315 \FA_INST_0[0].FA_INST_1[363].FA_  ( .A(A[363]), .B(n663), .CI(
        C[363]), .CO(C[364]) );
  FA_15314 \FA_INST_0[0].FA_INST_1[364].FA_  ( .A(A[364]), .B(n662), .CI(
        C[364]), .CO(C[365]) );
  FA_15313 \FA_INST_0[0].FA_INST_1[365].FA_  ( .A(A[365]), .B(n661), .CI(
        C[365]), .CO(C[366]) );
  FA_15312 \FA_INST_0[0].FA_INST_1[366].FA_  ( .A(A[366]), .B(n660), .CI(
        C[366]), .CO(C[367]) );
  FA_15311 \FA_INST_0[0].FA_INST_1[367].FA_  ( .A(A[367]), .B(n659), .CI(
        C[367]), .CO(C[368]) );
  FA_15310 \FA_INST_0[0].FA_INST_1[368].FA_  ( .A(A[368]), .B(n658), .CI(
        C[368]), .CO(C[369]) );
  FA_15309 \FA_INST_0[0].FA_INST_1[369].FA_  ( .A(A[369]), .B(n657), .CI(
        C[369]), .CO(C[370]) );
  FA_15308 \FA_INST_0[0].FA_INST_1[370].FA_  ( .A(A[370]), .B(n656), .CI(
        C[370]), .CO(C[371]) );
  FA_15307 \FA_INST_0[0].FA_INST_1[371].FA_  ( .A(A[371]), .B(n655), .CI(
        C[371]), .CO(C[372]) );
  FA_15306 \FA_INST_0[0].FA_INST_1[372].FA_  ( .A(A[372]), .B(n654), .CI(
        C[372]), .CO(C[373]) );
  FA_15305 \FA_INST_0[0].FA_INST_1[373].FA_  ( .A(A[373]), .B(n653), .CI(
        C[373]), .CO(C[374]) );
  FA_15304 \FA_INST_0[0].FA_INST_1[374].FA_  ( .A(A[374]), .B(n652), .CI(
        C[374]), .CO(C[375]) );
  FA_15303 \FA_INST_0[0].FA_INST_1[375].FA_  ( .A(A[375]), .B(n651), .CI(
        C[375]), .CO(C[376]) );
  FA_15302 \FA_INST_0[0].FA_INST_1[376].FA_  ( .A(A[376]), .B(n650), .CI(
        C[376]), .CO(C[377]) );
  FA_15301 \FA_INST_0[0].FA_INST_1[377].FA_  ( .A(A[377]), .B(n649), .CI(
        C[377]), .CO(C[378]) );
  FA_15300 \FA_INST_0[0].FA_INST_1[378].FA_  ( .A(A[378]), .B(n648), .CI(
        C[378]), .CO(C[379]) );
  FA_15299 \FA_INST_0[0].FA_INST_1[379].FA_  ( .A(A[379]), .B(n647), .CI(
        C[379]), .CO(C[380]) );
  FA_15298 \FA_INST_0[0].FA_INST_1[380].FA_  ( .A(A[380]), .B(n646), .CI(
        C[380]), .CO(C[381]) );
  FA_15297 \FA_INST_0[0].FA_INST_1[381].FA_  ( .A(A[381]), .B(n645), .CI(
        C[381]), .CO(C[382]) );
  FA_15296 \FA_INST_0[0].FA_INST_1[382].FA_  ( .A(A[382]), .B(n644), .CI(
        C[382]), .CO(C[383]) );
  FA_15295 \FA_INST_0[0].FA_INST_1[383].FA_  ( .A(A[383]), .B(n643), .CI(
        C[383]), .CO(C[384]) );
  FA_15294 \FA_INST_0[0].FA_INST_1[384].FA_  ( .A(A[384]), .B(n642), .CI(
        C[384]), .CO(C[385]) );
  FA_15293 \FA_INST_0[0].FA_INST_1[385].FA_  ( .A(A[385]), .B(n641), .CI(
        C[385]), .CO(C[386]) );
  FA_15292 \FA_INST_0[0].FA_INST_1[386].FA_  ( .A(A[386]), .B(n640), .CI(
        C[386]), .CO(C[387]) );
  FA_15291 \FA_INST_0[0].FA_INST_1[387].FA_  ( .A(A[387]), .B(n639), .CI(
        C[387]), .CO(C[388]) );
  FA_15290 \FA_INST_0[0].FA_INST_1[388].FA_  ( .A(A[388]), .B(n638), .CI(
        C[388]), .CO(C[389]) );
  FA_15289 \FA_INST_0[0].FA_INST_1[389].FA_  ( .A(A[389]), .B(n637), .CI(
        C[389]), .CO(C[390]) );
  FA_15288 \FA_INST_0[0].FA_INST_1[390].FA_  ( .A(A[390]), .B(n636), .CI(
        C[390]), .CO(C[391]) );
  FA_15287 \FA_INST_0[0].FA_INST_1[391].FA_  ( .A(A[391]), .B(n635), .CI(
        C[391]), .CO(C[392]) );
  FA_15286 \FA_INST_0[0].FA_INST_1[392].FA_  ( .A(A[392]), .B(n634), .CI(
        C[392]), .CO(C[393]) );
  FA_15285 \FA_INST_0[0].FA_INST_1[393].FA_  ( .A(A[393]), .B(n633), .CI(
        C[393]), .CO(C[394]) );
  FA_15284 \FA_INST_0[0].FA_INST_1[394].FA_  ( .A(A[394]), .B(n632), .CI(
        C[394]), .CO(C[395]) );
  FA_15283 \FA_INST_0[0].FA_INST_1[395].FA_  ( .A(A[395]), .B(n631), .CI(
        C[395]), .CO(C[396]) );
  FA_15282 \FA_INST_0[0].FA_INST_1[396].FA_  ( .A(A[396]), .B(n630), .CI(
        C[396]), .CO(C[397]) );
  FA_15281 \FA_INST_0[0].FA_INST_1[397].FA_  ( .A(A[397]), .B(n629), .CI(
        C[397]), .CO(C[398]) );
  FA_15280 \FA_INST_0[0].FA_INST_1[398].FA_  ( .A(A[398]), .B(n628), .CI(
        C[398]), .CO(C[399]) );
  FA_15279 \FA_INST_0[0].FA_INST_1[399].FA_  ( .A(A[399]), .B(n627), .CI(
        C[399]), .CO(C[400]) );
  FA_15278 \FA_INST_0[0].FA_INST_1[400].FA_  ( .A(A[400]), .B(n626), .CI(
        C[400]), .CO(C[401]) );
  FA_15277 \FA_INST_0[0].FA_INST_1[401].FA_  ( .A(A[401]), .B(n625), .CI(
        C[401]), .CO(C[402]) );
  FA_15276 \FA_INST_0[0].FA_INST_1[402].FA_  ( .A(A[402]), .B(n624), .CI(
        C[402]), .CO(C[403]) );
  FA_15275 \FA_INST_0[0].FA_INST_1[403].FA_  ( .A(A[403]), .B(n623), .CI(
        C[403]), .CO(C[404]) );
  FA_15274 \FA_INST_0[0].FA_INST_1[404].FA_  ( .A(A[404]), .B(n622), .CI(
        C[404]), .CO(C[405]) );
  FA_15273 \FA_INST_0[0].FA_INST_1[405].FA_  ( .A(A[405]), .B(n621), .CI(
        C[405]), .CO(C[406]) );
  FA_15272 \FA_INST_0[0].FA_INST_1[406].FA_  ( .A(A[406]), .B(n620), .CI(
        C[406]), .CO(C[407]) );
  FA_15271 \FA_INST_0[0].FA_INST_1[407].FA_  ( .A(A[407]), .B(n619), .CI(
        C[407]), .CO(C[408]) );
  FA_15270 \FA_INST_0[0].FA_INST_1[408].FA_  ( .A(A[408]), .B(n618), .CI(
        C[408]), .CO(C[409]) );
  FA_15269 \FA_INST_0[0].FA_INST_1[409].FA_  ( .A(A[409]), .B(n617), .CI(
        C[409]), .CO(C[410]) );
  FA_15268 \FA_INST_0[0].FA_INST_1[410].FA_  ( .A(A[410]), .B(n616), .CI(
        C[410]), .CO(C[411]) );
  FA_15267 \FA_INST_0[0].FA_INST_1[411].FA_  ( .A(A[411]), .B(n615), .CI(
        C[411]), .CO(C[412]) );
  FA_15266 \FA_INST_0[0].FA_INST_1[412].FA_  ( .A(A[412]), .B(n614), .CI(
        C[412]), .CO(C[413]) );
  FA_15265 \FA_INST_0[0].FA_INST_1[413].FA_  ( .A(A[413]), .B(n613), .CI(
        C[413]), .CO(C[414]) );
  FA_15264 \FA_INST_0[0].FA_INST_1[414].FA_  ( .A(A[414]), .B(n612), .CI(
        C[414]), .CO(C[415]) );
  FA_15263 \FA_INST_0[0].FA_INST_1[415].FA_  ( .A(A[415]), .B(n611), .CI(
        C[415]), .CO(C[416]) );
  FA_15262 \FA_INST_0[0].FA_INST_1[416].FA_  ( .A(A[416]), .B(n610), .CI(
        C[416]), .CO(C[417]) );
  FA_15261 \FA_INST_0[0].FA_INST_1[417].FA_  ( .A(A[417]), .B(n609), .CI(
        C[417]), .CO(C[418]) );
  FA_15260 \FA_INST_0[0].FA_INST_1[418].FA_  ( .A(A[418]), .B(n608), .CI(
        C[418]), .CO(C[419]) );
  FA_15259 \FA_INST_0[0].FA_INST_1[419].FA_  ( .A(A[419]), .B(n607), .CI(
        C[419]), .CO(C[420]) );
  FA_15258 \FA_INST_0[0].FA_INST_1[420].FA_  ( .A(A[420]), .B(n606), .CI(
        C[420]), .CO(C[421]) );
  FA_15257 \FA_INST_0[0].FA_INST_1[421].FA_  ( .A(A[421]), .B(n605), .CI(
        C[421]), .CO(C[422]) );
  FA_15256 \FA_INST_0[0].FA_INST_1[422].FA_  ( .A(A[422]), .B(n604), .CI(
        C[422]), .CO(C[423]) );
  FA_15255 \FA_INST_0[0].FA_INST_1[423].FA_  ( .A(A[423]), .B(n603), .CI(
        C[423]), .CO(C[424]) );
  FA_15254 \FA_INST_0[0].FA_INST_1[424].FA_  ( .A(A[424]), .B(n602), .CI(
        C[424]), .CO(C[425]) );
  FA_15253 \FA_INST_0[0].FA_INST_1[425].FA_  ( .A(A[425]), .B(n601), .CI(
        C[425]), .CO(C[426]) );
  FA_15252 \FA_INST_0[0].FA_INST_1[426].FA_  ( .A(A[426]), .B(n600), .CI(
        C[426]), .CO(C[427]) );
  FA_15251 \FA_INST_0[0].FA_INST_1[427].FA_  ( .A(A[427]), .B(n599), .CI(
        C[427]), .CO(C[428]) );
  FA_15250 \FA_INST_0[0].FA_INST_1[428].FA_  ( .A(A[428]), .B(n598), .CI(
        C[428]), .CO(C[429]) );
  FA_15249 \FA_INST_0[0].FA_INST_1[429].FA_  ( .A(A[429]), .B(n597), .CI(
        C[429]), .CO(C[430]) );
  FA_15248 \FA_INST_0[0].FA_INST_1[430].FA_  ( .A(A[430]), .B(n596), .CI(
        C[430]), .CO(C[431]) );
  FA_15247 \FA_INST_0[0].FA_INST_1[431].FA_  ( .A(A[431]), .B(n595), .CI(
        C[431]), .CO(C[432]) );
  FA_15246 \FA_INST_0[0].FA_INST_1[432].FA_  ( .A(A[432]), .B(n594), .CI(
        C[432]), .CO(C[433]) );
  FA_15245 \FA_INST_0[0].FA_INST_1[433].FA_  ( .A(A[433]), .B(n593), .CI(
        C[433]), .CO(C[434]) );
  FA_15244 \FA_INST_0[0].FA_INST_1[434].FA_  ( .A(A[434]), .B(n592), .CI(
        C[434]), .CO(C[435]) );
  FA_15243 \FA_INST_0[0].FA_INST_1[435].FA_  ( .A(A[435]), .B(n591), .CI(
        C[435]), .CO(C[436]) );
  FA_15242 \FA_INST_0[0].FA_INST_1[436].FA_  ( .A(A[436]), .B(n590), .CI(
        C[436]), .CO(C[437]) );
  FA_15241 \FA_INST_0[0].FA_INST_1[437].FA_  ( .A(A[437]), .B(n589), .CI(
        C[437]), .CO(C[438]) );
  FA_15240 \FA_INST_0[0].FA_INST_1[438].FA_  ( .A(A[438]), .B(n588), .CI(
        C[438]), .CO(C[439]) );
  FA_15239 \FA_INST_0[0].FA_INST_1[439].FA_  ( .A(A[439]), .B(n587), .CI(
        C[439]), .CO(C[440]) );
  FA_15238 \FA_INST_0[0].FA_INST_1[440].FA_  ( .A(A[440]), .B(n586), .CI(
        C[440]), .CO(C[441]) );
  FA_15237 \FA_INST_0[0].FA_INST_1[441].FA_  ( .A(A[441]), .B(n585), .CI(
        C[441]), .CO(C[442]) );
  FA_15236 \FA_INST_0[0].FA_INST_1[442].FA_  ( .A(A[442]), .B(n584), .CI(
        C[442]), .CO(C[443]) );
  FA_15235 \FA_INST_0[0].FA_INST_1[443].FA_  ( .A(A[443]), .B(n583), .CI(
        C[443]), .CO(C[444]) );
  FA_15234 \FA_INST_0[0].FA_INST_1[444].FA_  ( .A(A[444]), .B(n582), .CI(
        C[444]), .CO(C[445]) );
  FA_15233 \FA_INST_0[0].FA_INST_1[445].FA_  ( .A(A[445]), .B(n581), .CI(
        C[445]), .CO(C[446]) );
  FA_15232 \FA_INST_0[0].FA_INST_1[446].FA_  ( .A(A[446]), .B(n580), .CI(
        C[446]), .CO(C[447]) );
  FA_15231 \FA_INST_0[0].FA_INST_1[447].FA_  ( .A(A[447]), .B(n579), .CI(
        C[447]), .CO(C[448]) );
  FA_15230 \FA_INST_0[0].FA_INST_1[448].FA_  ( .A(A[448]), .B(n578), .CI(
        C[448]), .CO(C[449]) );
  FA_15229 \FA_INST_0[0].FA_INST_1[449].FA_  ( .A(A[449]), .B(n577), .CI(
        C[449]), .CO(C[450]) );
  FA_15228 \FA_INST_0[0].FA_INST_1[450].FA_  ( .A(A[450]), .B(n576), .CI(
        C[450]), .CO(C[451]) );
  FA_15227 \FA_INST_0[0].FA_INST_1[451].FA_  ( .A(A[451]), .B(n575), .CI(
        C[451]), .CO(C[452]) );
  FA_15226 \FA_INST_0[0].FA_INST_1[452].FA_  ( .A(A[452]), .B(n574), .CI(
        C[452]), .CO(C[453]) );
  FA_15225 \FA_INST_0[0].FA_INST_1[453].FA_  ( .A(A[453]), .B(n573), .CI(
        C[453]), .CO(C[454]) );
  FA_15224 \FA_INST_0[0].FA_INST_1[454].FA_  ( .A(A[454]), .B(n572), .CI(
        C[454]), .CO(C[455]) );
  FA_15223 \FA_INST_0[0].FA_INST_1[455].FA_  ( .A(A[455]), .B(n571), .CI(
        C[455]), .CO(C[456]) );
  FA_15222 \FA_INST_0[0].FA_INST_1[456].FA_  ( .A(A[456]), .B(n570), .CI(
        C[456]), .CO(C[457]) );
  FA_15221 \FA_INST_0[0].FA_INST_1[457].FA_  ( .A(A[457]), .B(n569), .CI(
        C[457]), .CO(C[458]) );
  FA_15220 \FA_INST_0[0].FA_INST_1[458].FA_  ( .A(A[458]), .B(n568), .CI(
        C[458]), .CO(C[459]) );
  FA_15219 \FA_INST_0[0].FA_INST_1[459].FA_  ( .A(A[459]), .B(n567), .CI(
        C[459]), .CO(C[460]) );
  FA_15218 \FA_INST_0[0].FA_INST_1[460].FA_  ( .A(A[460]), .B(n566), .CI(
        C[460]), .CO(C[461]) );
  FA_15217 \FA_INST_0[0].FA_INST_1[461].FA_  ( .A(A[461]), .B(n565), .CI(
        C[461]), .CO(C[462]) );
  FA_15216 \FA_INST_0[0].FA_INST_1[462].FA_  ( .A(A[462]), .B(n564), .CI(
        C[462]), .CO(C[463]) );
  FA_15215 \FA_INST_0[0].FA_INST_1[463].FA_  ( .A(A[463]), .B(n563), .CI(
        C[463]), .CO(C[464]) );
  FA_15214 \FA_INST_0[0].FA_INST_1[464].FA_  ( .A(A[464]), .B(n562), .CI(
        C[464]), .CO(C[465]) );
  FA_15213 \FA_INST_0[0].FA_INST_1[465].FA_  ( .A(A[465]), .B(n561), .CI(
        C[465]), .CO(C[466]) );
  FA_15212 \FA_INST_0[0].FA_INST_1[466].FA_  ( .A(A[466]), .B(n560), .CI(
        C[466]), .CO(C[467]) );
  FA_15211 \FA_INST_0[0].FA_INST_1[467].FA_  ( .A(A[467]), .B(n559), .CI(
        C[467]), .CO(C[468]) );
  FA_15210 \FA_INST_0[0].FA_INST_1[468].FA_  ( .A(A[468]), .B(n558), .CI(
        C[468]), .CO(C[469]) );
  FA_15209 \FA_INST_0[0].FA_INST_1[469].FA_  ( .A(A[469]), .B(n557), .CI(
        C[469]), .CO(C[470]) );
  FA_15208 \FA_INST_0[0].FA_INST_1[470].FA_  ( .A(A[470]), .B(n556), .CI(
        C[470]), .CO(C[471]) );
  FA_15207 \FA_INST_0[0].FA_INST_1[471].FA_  ( .A(A[471]), .B(n555), .CI(
        C[471]), .CO(C[472]) );
  FA_15206 \FA_INST_0[0].FA_INST_1[472].FA_  ( .A(A[472]), .B(n554), .CI(
        C[472]), .CO(C[473]) );
  FA_15205 \FA_INST_0[0].FA_INST_1[473].FA_  ( .A(A[473]), .B(n553), .CI(
        C[473]), .CO(C[474]) );
  FA_15204 \FA_INST_0[0].FA_INST_1[474].FA_  ( .A(A[474]), .B(n552), .CI(
        C[474]), .CO(C[475]) );
  FA_15203 \FA_INST_0[0].FA_INST_1[475].FA_  ( .A(A[475]), .B(n551), .CI(
        C[475]), .CO(C[476]) );
  FA_15202 \FA_INST_0[0].FA_INST_1[476].FA_  ( .A(A[476]), .B(n550), .CI(
        C[476]), .CO(C[477]) );
  FA_15201 \FA_INST_0[0].FA_INST_1[477].FA_  ( .A(A[477]), .B(n549), .CI(
        C[477]), .CO(C[478]) );
  FA_15200 \FA_INST_0[0].FA_INST_1[478].FA_  ( .A(A[478]), .B(n548), .CI(
        C[478]), .CO(C[479]) );
  FA_15199 \FA_INST_0[0].FA_INST_1[479].FA_  ( .A(A[479]), .B(n547), .CI(
        C[479]), .CO(C[480]) );
  FA_15198 \FA_INST_0[0].FA_INST_1[480].FA_  ( .A(A[480]), .B(n546), .CI(
        C[480]), .CO(C[481]) );
  FA_15197 \FA_INST_0[0].FA_INST_1[481].FA_  ( .A(A[481]), .B(n545), .CI(
        C[481]), .CO(C[482]) );
  FA_15196 \FA_INST_0[0].FA_INST_1[482].FA_  ( .A(A[482]), .B(n544), .CI(
        C[482]), .CO(C[483]) );
  FA_15195 \FA_INST_0[0].FA_INST_1[483].FA_  ( .A(A[483]), .B(n543), .CI(
        C[483]), .CO(C[484]) );
  FA_15194 \FA_INST_0[0].FA_INST_1[484].FA_  ( .A(A[484]), .B(n542), .CI(
        C[484]), .CO(C[485]) );
  FA_15193 \FA_INST_0[0].FA_INST_1[485].FA_  ( .A(A[485]), .B(n541), .CI(
        C[485]), .CO(C[486]) );
  FA_15192 \FA_INST_0[0].FA_INST_1[486].FA_  ( .A(A[486]), .B(n540), .CI(
        C[486]), .CO(C[487]) );
  FA_15191 \FA_INST_0[0].FA_INST_1[487].FA_  ( .A(A[487]), .B(n539), .CI(
        C[487]), .CO(C[488]) );
  FA_15190 \FA_INST_0[0].FA_INST_1[488].FA_  ( .A(A[488]), .B(n538), .CI(
        C[488]), .CO(C[489]) );
  FA_15189 \FA_INST_0[0].FA_INST_1[489].FA_  ( .A(A[489]), .B(n537), .CI(
        C[489]), .CO(C[490]) );
  FA_15188 \FA_INST_0[0].FA_INST_1[490].FA_  ( .A(A[490]), .B(n536), .CI(
        C[490]), .CO(C[491]) );
  FA_15187 \FA_INST_0[0].FA_INST_1[491].FA_  ( .A(A[491]), .B(n535), .CI(
        C[491]), .CO(C[492]) );
  FA_15186 \FA_INST_0[0].FA_INST_1[492].FA_  ( .A(A[492]), .B(n534), .CI(
        C[492]), .CO(C[493]) );
  FA_15185 \FA_INST_0[0].FA_INST_1[493].FA_  ( .A(A[493]), .B(n533), .CI(
        C[493]), .CO(C[494]) );
  FA_15184 \FA_INST_0[0].FA_INST_1[494].FA_  ( .A(A[494]), .B(n532), .CI(
        C[494]), .CO(C[495]) );
  FA_15183 \FA_INST_0[0].FA_INST_1[495].FA_  ( .A(A[495]), .B(n531), .CI(
        C[495]), .CO(C[496]) );
  FA_15182 \FA_INST_0[0].FA_INST_1[496].FA_  ( .A(A[496]), .B(n530), .CI(
        C[496]), .CO(C[497]) );
  FA_15181 \FA_INST_0[0].FA_INST_1[497].FA_  ( .A(A[497]), .B(n529), .CI(
        C[497]), .CO(C[498]) );
  FA_15180 \FA_INST_0[0].FA_INST_1[498].FA_  ( .A(A[498]), .B(n528), .CI(
        C[498]), .CO(C[499]) );
  FA_15179 \FA_INST_0[0].FA_INST_1[499].FA_  ( .A(A[499]), .B(n527), .CI(
        C[499]), .CO(C[500]) );
  FA_15178 \FA_INST_0[0].FA_INST_1[500].FA_  ( .A(A[500]), .B(n526), .CI(
        C[500]), .CO(C[501]) );
  FA_15177 \FA_INST_0[0].FA_INST_1[501].FA_  ( .A(A[501]), .B(n525), .CI(
        C[501]), .CO(C[502]) );
  FA_15176 \FA_INST_0[0].FA_INST_1[502].FA_  ( .A(A[502]), .B(n524), .CI(
        C[502]), .CO(C[503]) );
  FA_15175 \FA_INST_0[0].FA_INST_1[503].FA_  ( .A(A[503]), .B(n523), .CI(
        C[503]), .CO(C[504]) );
  FA_15174 \FA_INST_0[0].FA_INST_1[504].FA_  ( .A(A[504]), .B(n522), .CI(
        C[504]), .CO(C[505]) );
  FA_15173 \FA_INST_0[0].FA_INST_1[505].FA_  ( .A(A[505]), .B(n521), .CI(
        C[505]), .CO(C[506]) );
  FA_15172 \FA_INST_0[0].FA_INST_1[506].FA_  ( .A(A[506]), .B(n520), .CI(
        C[506]), .CO(C[507]) );
  FA_15171 \FA_INST_0[0].FA_INST_1[507].FA_  ( .A(A[507]), .B(n519), .CI(
        C[507]), .CO(C[508]) );
  FA_15170 \FA_INST_0[0].FA_INST_1[508].FA_  ( .A(A[508]), .B(n518), .CI(
        C[508]), .CO(C[509]) );
  FA_15169 \FA_INST_0[0].FA_INST_1[509].FA_  ( .A(A[509]), .B(n517), .CI(
        C[509]), .CO(C[510]) );
  FA_15168 \FA_INST_0[0].FA_INST_1[510].FA_  ( .A(A[510]), .B(n516), .CI(
        C[510]), .CO(C[511]) );
  FA_15167 \FA_INST_0[0].FA_INST_1[511].FA_  ( .A(A[511]), .B(n515), .CI(
        C[511]), .CO(C[512]) );
  FA_15166 \FA_INST_0[1].FA_INST_1[0].FA_  ( .A(A[512]), .B(n514), .CI(C[512]), 
        .CO(C[513]) );
  FA_15165 \FA_INST_0[1].FA_INST_1[1].FA_  ( .A(A[513]), .B(n513), .CI(C[513]), 
        .CO(C[514]) );
  FA_15164 \FA_INST_0[1].FA_INST_1[2].FA_  ( .A(A[514]), .B(n512), .CI(C[514]), 
        .CO(C[515]) );
  FA_15163 \FA_INST_0[1].FA_INST_1[3].FA_  ( .A(A[515]), .B(n511), .CI(C[515]), 
        .CO(C[516]) );
  FA_15162 \FA_INST_0[1].FA_INST_1[4].FA_  ( .A(A[516]), .B(n510), .CI(C[516]), 
        .CO(C[517]) );
  FA_15161 \FA_INST_0[1].FA_INST_1[5].FA_  ( .A(A[517]), .B(n509), .CI(C[517]), 
        .CO(C[518]) );
  FA_15160 \FA_INST_0[1].FA_INST_1[6].FA_  ( .A(A[518]), .B(n508), .CI(C[518]), 
        .CO(C[519]) );
  FA_15159 \FA_INST_0[1].FA_INST_1[7].FA_  ( .A(A[519]), .B(n507), .CI(C[519]), 
        .CO(C[520]) );
  FA_15158 \FA_INST_0[1].FA_INST_1[8].FA_  ( .A(A[520]), .B(n506), .CI(C[520]), 
        .CO(C[521]) );
  FA_15157 \FA_INST_0[1].FA_INST_1[9].FA_  ( .A(A[521]), .B(n505), .CI(C[521]), 
        .CO(C[522]) );
  FA_15156 \FA_INST_0[1].FA_INST_1[10].FA_  ( .A(A[522]), .B(n504), .CI(C[522]), .CO(C[523]) );
  FA_15155 \FA_INST_0[1].FA_INST_1[11].FA_  ( .A(A[523]), .B(n503), .CI(C[523]), .CO(C[524]) );
  FA_15154 \FA_INST_0[1].FA_INST_1[12].FA_  ( .A(A[524]), .B(n502), .CI(C[524]), .CO(C[525]) );
  FA_15153 \FA_INST_0[1].FA_INST_1[13].FA_  ( .A(A[525]), .B(n501), .CI(C[525]), .CO(C[526]) );
  FA_15152 \FA_INST_0[1].FA_INST_1[14].FA_  ( .A(A[526]), .B(n500), .CI(C[526]), .CO(C[527]) );
  FA_15151 \FA_INST_0[1].FA_INST_1[15].FA_  ( .A(A[527]), .B(n499), .CI(C[527]), .CO(C[528]) );
  FA_15150 \FA_INST_0[1].FA_INST_1[16].FA_  ( .A(A[528]), .B(n498), .CI(C[528]), .CO(C[529]) );
  FA_15149 \FA_INST_0[1].FA_INST_1[17].FA_  ( .A(A[529]), .B(n497), .CI(C[529]), .CO(C[530]) );
  FA_15148 \FA_INST_0[1].FA_INST_1[18].FA_  ( .A(A[530]), .B(n496), .CI(C[530]), .CO(C[531]) );
  FA_15147 \FA_INST_0[1].FA_INST_1[19].FA_  ( .A(A[531]), .B(n495), .CI(C[531]), .CO(C[532]) );
  FA_15146 \FA_INST_0[1].FA_INST_1[20].FA_  ( .A(A[532]), .B(n494), .CI(C[532]), .CO(C[533]) );
  FA_15145 \FA_INST_0[1].FA_INST_1[21].FA_  ( .A(A[533]), .B(n493), .CI(C[533]), .CO(C[534]) );
  FA_15144 \FA_INST_0[1].FA_INST_1[22].FA_  ( .A(A[534]), .B(n492), .CI(C[534]), .CO(C[535]) );
  FA_15143 \FA_INST_0[1].FA_INST_1[23].FA_  ( .A(A[535]), .B(n491), .CI(C[535]), .CO(C[536]) );
  FA_15142 \FA_INST_0[1].FA_INST_1[24].FA_  ( .A(A[536]), .B(n490), .CI(C[536]), .CO(C[537]) );
  FA_15141 \FA_INST_0[1].FA_INST_1[25].FA_  ( .A(A[537]), .B(n489), .CI(C[537]), .CO(C[538]) );
  FA_15140 \FA_INST_0[1].FA_INST_1[26].FA_  ( .A(A[538]), .B(n488), .CI(C[538]), .CO(C[539]) );
  FA_15139 \FA_INST_0[1].FA_INST_1[27].FA_  ( .A(A[539]), .B(n487), .CI(C[539]), .CO(C[540]) );
  FA_15138 \FA_INST_0[1].FA_INST_1[28].FA_  ( .A(A[540]), .B(n486), .CI(C[540]), .CO(C[541]) );
  FA_15137 \FA_INST_0[1].FA_INST_1[29].FA_  ( .A(A[541]), .B(n485), .CI(C[541]), .CO(C[542]) );
  FA_15136 \FA_INST_0[1].FA_INST_1[30].FA_  ( .A(A[542]), .B(n484), .CI(C[542]), .CO(C[543]) );
  FA_15135 \FA_INST_0[1].FA_INST_1[31].FA_  ( .A(A[543]), .B(n483), .CI(C[543]), .CO(C[544]) );
  FA_15134 \FA_INST_0[1].FA_INST_1[32].FA_  ( .A(A[544]), .B(n482), .CI(C[544]), .CO(C[545]) );
  FA_15133 \FA_INST_0[1].FA_INST_1[33].FA_  ( .A(A[545]), .B(n481), .CI(C[545]), .CO(C[546]) );
  FA_15132 \FA_INST_0[1].FA_INST_1[34].FA_  ( .A(A[546]), .B(n480), .CI(C[546]), .CO(C[547]) );
  FA_15131 \FA_INST_0[1].FA_INST_1[35].FA_  ( .A(A[547]), .B(n479), .CI(C[547]), .CO(C[548]) );
  FA_15130 \FA_INST_0[1].FA_INST_1[36].FA_  ( .A(A[548]), .B(n478), .CI(C[548]), .CO(C[549]) );
  FA_15129 \FA_INST_0[1].FA_INST_1[37].FA_  ( .A(A[549]), .B(n477), .CI(C[549]), .CO(C[550]) );
  FA_15128 \FA_INST_0[1].FA_INST_1[38].FA_  ( .A(A[550]), .B(n476), .CI(C[550]), .CO(C[551]) );
  FA_15127 \FA_INST_0[1].FA_INST_1[39].FA_  ( .A(A[551]), .B(n475), .CI(C[551]), .CO(C[552]) );
  FA_15126 \FA_INST_0[1].FA_INST_1[40].FA_  ( .A(A[552]), .B(n474), .CI(C[552]), .CO(C[553]) );
  FA_15125 \FA_INST_0[1].FA_INST_1[41].FA_  ( .A(A[553]), .B(n473), .CI(C[553]), .CO(C[554]) );
  FA_15124 \FA_INST_0[1].FA_INST_1[42].FA_  ( .A(A[554]), .B(n472), .CI(C[554]), .CO(C[555]) );
  FA_15123 \FA_INST_0[1].FA_INST_1[43].FA_  ( .A(A[555]), .B(n471), .CI(C[555]), .CO(C[556]) );
  FA_15122 \FA_INST_0[1].FA_INST_1[44].FA_  ( .A(A[556]), .B(n470), .CI(C[556]), .CO(C[557]) );
  FA_15121 \FA_INST_0[1].FA_INST_1[45].FA_  ( .A(A[557]), .B(n469), .CI(C[557]), .CO(C[558]) );
  FA_15120 \FA_INST_0[1].FA_INST_1[46].FA_  ( .A(A[558]), .B(n468), .CI(C[558]), .CO(C[559]) );
  FA_15119 \FA_INST_0[1].FA_INST_1[47].FA_  ( .A(A[559]), .B(n467), .CI(C[559]), .CO(C[560]) );
  FA_15118 \FA_INST_0[1].FA_INST_1[48].FA_  ( .A(A[560]), .B(n466), .CI(C[560]), .CO(C[561]) );
  FA_15117 \FA_INST_0[1].FA_INST_1[49].FA_  ( .A(A[561]), .B(n465), .CI(C[561]), .CO(C[562]) );
  FA_15116 \FA_INST_0[1].FA_INST_1[50].FA_  ( .A(A[562]), .B(n464), .CI(C[562]), .CO(C[563]) );
  FA_15115 \FA_INST_0[1].FA_INST_1[51].FA_  ( .A(A[563]), .B(n463), .CI(C[563]), .CO(C[564]) );
  FA_15114 \FA_INST_0[1].FA_INST_1[52].FA_  ( .A(A[564]), .B(n462), .CI(C[564]), .CO(C[565]) );
  FA_15113 \FA_INST_0[1].FA_INST_1[53].FA_  ( .A(A[565]), .B(n461), .CI(C[565]), .CO(C[566]) );
  FA_15112 \FA_INST_0[1].FA_INST_1[54].FA_  ( .A(A[566]), .B(n460), .CI(C[566]), .CO(C[567]) );
  FA_15111 \FA_INST_0[1].FA_INST_1[55].FA_  ( .A(A[567]), .B(n459), .CI(C[567]), .CO(C[568]) );
  FA_15110 \FA_INST_0[1].FA_INST_1[56].FA_  ( .A(A[568]), .B(n458), .CI(C[568]), .CO(C[569]) );
  FA_15109 \FA_INST_0[1].FA_INST_1[57].FA_  ( .A(A[569]), .B(n457), .CI(C[569]), .CO(C[570]) );
  FA_15108 \FA_INST_0[1].FA_INST_1[58].FA_  ( .A(A[570]), .B(n456), .CI(C[570]), .CO(C[571]) );
  FA_15107 \FA_INST_0[1].FA_INST_1[59].FA_  ( .A(A[571]), .B(n455), .CI(C[571]), .CO(C[572]) );
  FA_15106 \FA_INST_0[1].FA_INST_1[60].FA_  ( .A(A[572]), .B(n454), .CI(C[572]), .CO(C[573]) );
  FA_15105 \FA_INST_0[1].FA_INST_1[61].FA_  ( .A(A[573]), .B(n453), .CI(C[573]), .CO(C[574]) );
  FA_15104 \FA_INST_0[1].FA_INST_1[62].FA_  ( .A(A[574]), .B(n452), .CI(C[574]), .CO(C[575]) );
  FA_15103 \FA_INST_0[1].FA_INST_1[63].FA_  ( .A(A[575]), .B(n451), .CI(C[575]), .CO(C[576]) );
  FA_15102 \FA_INST_0[1].FA_INST_1[64].FA_  ( .A(A[576]), .B(n450), .CI(C[576]), .CO(C[577]) );
  FA_15101 \FA_INST_0[1].FA_INST_1[65].FA_  ( .A(A[577]), .B(n449), .CI(C[577]), .CO(C[578]) );
  FA_15100 \FA_INST_0[1].FA_INST_1[66].FA_  ( .A(A[578]), .B(n448), .CI(C[578]), .CO(C[579]) );
  FA_15099 \FA_INST_0[1].FA_INST_1[67].FA_  ( .A(A[579]), .B(n447), .CI(C[579]), .CO(C[580]) );
  FA_15098 \FA_INST_0[1].FA_INST_1[68].FA_  ( .A(A[580]), .B(n446), .CI(C[580]), .CO(C[581]) );
  FA_15097 \FA_INST_0[1].FA_INST_1[69].FA_  ( .A(A[581]), .B(n445), .CI(C[581]), .CO(C[582]) );
  FA_15096 \FA_INST_0[1].FA_INST_1[70].FA_  ( .A(A[582]), .B(n444), .CI(C[582]), .CO(C[583]) );
  FA_15095 \FA_INST_0[1].FA_INST_1[71].FA_  ( .A(A[583]), .B(n443), .CI(C[583]), .CO(C[584]) );
  FA_15094 \FA_INST_0[1].FA_INST_1[72].FA_  ( .A(A[584]), .B(n442), .CI(C[584]), .CO(C[585]) );
  FA_15093 \FA_INST_0[1].FA_INST_1[73].FA_  ( .A(A[585]), .B(n441), .CI(C[585]), .CO(C[586]) );
  FA_15092 \FA_INST_0[1].FA_INST_1[74].FA_  ( .A(A[586]), .B(n440), .CI(C[586]), .CO(C[587]) );
  FA_15091 \FA_INST_0[1].FA_INST_1[75].FA_  ( .A(A[587]), .B(n439), .CI(C[587]), .CO(C[588]) );
  FA_15090 \FA_INST_0[1].FA_INST_1[76].FA_  ( .A(A[588]), .B(n438), .CI(C[588]), .CO(C[589]) );
  FA_15089 \FA_INST_0[1].FA_INST_1[77].FA_  ( .A(A[589]), .B(n437), .CI(C[589]), .CO(C[590]) );
  FA_15088 \FA_INST_0[1].FA_INST_1[78].FA_  ( .A(A[590]), .B(n436), .CI(C[590]), .CO(C[591]) );
  FA_15087 \FA_INST_0[1].FA_INST_1[79].FA_  ( .A(A[591]), .B(n435), .CI(C[591]), .CO(C[592]) );
  FA_15086 \FA_INST_0[1].FA_INST_1[80].FA_  ( .A(A[592]), .B(n434), .CI(C[592]), .CO(C[593]) );
  FA_15085 \FA_INST_0[1].FA_INST_1[81].FA_  ( .A(A[593]), .B(n433), .CI(C[593]), .CO(C[594]) );
  FA_15084 \FA_INST_0[1].FA_INST_1[82].FA_  ( .A(A[594]), .B(n432), .CI(C[594]), .CO(C[595]) );
  FA_15083 \FA_INST_0[1].FA_INST_1[83].FA_  ( .A(A[595]), .B(n431), .CI(C[595]), .CO(C[596]) );
  FA_15082 \FA_INST_0[1].FA_INST_1[84].FA_  ( .A(A[596]), .B(n430), .CI(C[596]), .CO(C[597]) );
  FA_15081 \FA_INST_0[1].FA_INST_1[85].FA_  ( .A(A[597]), .B(n429), .CI(C[597]), .CO(C[598]) );
  FA_15080 \FA_INST_0[1].FA_INST_1[86].FA_  ( .A(A[598]), .B(n428), .CI(C[598]), .CO(C[599]) );
  FA_15079 \FA_INST_0[1].FA_INST_1[87].FA_  ( .A(A[599]), .B(n427), .CI(C[599]), .CO(C[600]) );
  FA_15078 \FA_INST_0[1].FA_INST_1[88].FA_  ( .A(A[600]), .B(n426), .CI(C[600]), .CO(C[601]) );
  FA_15077 \FA_INST_0[1].FA_INST_1[89].FA_  ( .A(A[601]), .B(n425), .CI(C[601]), .CO(C[602]) );
  FA_15076 \FA_INST_0[1].FA_INST_1[90].FA_  ( .A(A[602]), .B(n424), .CI(C[602]), .CO(C[603]) );
  FA_15075 \FA_INST_0[1].FA_INST_1[91].FA_  ( .A(A[603]), .B(n423), .CI(C[603]), .CO(C[604]) );
  FA_15074 \FA_INST_0[1].FA_INST_1[92].FA_  ( .A(A[604]), .B(n422), .CI(C[604]), .CO(C[605]) );
  FA_15073 \FA_INST_0[1].FA_INST_1[93].FA_  ( .A(A[605]), .B(n421), .CI(C[605]), .CO(C[606]) );
  FA_15072 \FA_INST_0[1].FA_INST_1[94].FA_  ( .A(A[606]), .B(n420), .CI(C[606]), .CO(C[607]) );
  FA_15071 \FA_INST_0[1].FA_INST_1[95].FA_  ( .A(A[607]), .B(n419), .CI(C[607]), .CO(C[608]) );
  FA_15070 \FA_INST_0[1].FA_INST_1[96].FA_  ( .A(A[608]), .B(n418), .CI(C[608]), .CO(C[609]) );
  FA_15069 \FA_INST_0[1].FA_INST_1[97].FA_  ( .A(A[609]), .B(n417), .CI(C[609]), .CO(C[610]) );
  FA_15068 \FA_INST_0[1].FA_INST_1[98].FA_  ( .A(A[610]), .B(n416), .CI(C[610]), .CO(C[611]) );
  FA_15067 \FA_INST_0[1].FA_INST_1[99].FA_  ( .A(A[611]), .B(n415), .CI(C[611]), .CO(C[612]) );
  FA_15066 \FA_INST_0[1].FA_INST_1[100].FA_  ( .A(A[612]), .B(n414), .CI(
        C[612]), .CO(C[613]) );
  FA_15065 \FA_INST_0[1].FA_INST_1[101].FA_  ( .A(A[613]), .B(n413), .CI(
        C[613]), .CO(C[614]) );
  FA_15064 \FA_INST_0[1].FA_INST_1[102].FA_  ( .A(A[614]), .B(n412), .CI(
        C[614]), .CO(C[615]) );
  FA_15063 \FA_INST_0[1].FA_INST_1[103].FA_  ( .A(A[615]), .B(n411), .CI(
        C[615]), .CO(C[616]) );
  FA_15062 \FA_INST_0[1].FA_INST_1[104].FA_  ( .A(A[616]), .B(n410), .CI(
        C[616]), .CO(C[617]) );
  FA_15061 \FA_INST_0[1].FA_INST_1[105].FA_  ( .A(A[617]), .B(n409), .CI(
        C[617]), .CO(C[618]) );
  FA_15060 \FA_INST_0[1].FA_INST_1[106].FA_  ( .A(A[618]), .B(n408), .CI(
        C[618]), .CO(C[619]) );
  FA_15059 \FA_INST_0[1].FA_INST_1[107].FA_  ( .A(A[619]), .B(n407), .CI(
        C[619]), .CO(C[620]) );
  FA_15058 \FA_INST_0[1].FA_INST_1[108].FA_  ( .A(A[620]), .B(n406), .CI(
        C[620]), .CO(C[621]) );
  FA_15057 \FA_INST_0[1].FA_INST_1[109].FA_  ( .A(A[621]), .B(n405), .CI(
        C[621]), .CO(C[622]) );
  FA_15056 \FA_INST_0[1].FA_INST_1[110].FA_  ( .A(A[622]), .B(n404), .CI(
        C[622]), .CO(C[623]) );
  FA_15055 \FA_INST_0[1].FA_INST_1[111].FA_  ( .A(A[623]), .B(n403), .CI(
        C[623]), .CO(C[624]) );
  FA_15054 \FA_INST_0[1].FA_INST_1[112].FA_  ( .A(A[624]), .B(n402), .CI(
        C[624]), .CO(C[625]) );
  FA_15053 \FA_INST_0[1].FA_INST_1[113].FA_  ( .A(A[625]), .B(n401), .CI(
        C[625]), .CO(C[626]) );
  FA_15052 \FA_INST_0[1].FA_INST_1[114].FA_  ( .A(A[626]), .B(n400), .CI(
        C[626]), .CO(C[627]) );
  FA_15051 \FA_INST_0[1].FA_INST_1[115].FA_  ( .A(A[627]), .B(n399), .CI(
        C[627]), .CO(C[628]) );
  FA_15050 \FA_INST_0[1].FA_INST_1[116].FA_  ( .A(A[628]), .B(n398), .CI(
        C[628]), .CO(C[629]) );
  FA_15049 \FA_INST_0[1].FA_INST_1[117].FA_  ( .A(A[629]), .B(n397), .CI(
        C[629]), .CO(C[630]) );
  FA_15048 \FA_INST_0[1].FA_INST_1[118].FA_  ( .A(A[630]), .B(n396), .CI(
        C[630]), .CO(C[631]) );
  FA_15047 \FA_INST_0[1].FA_INST_1[119].FA_  ( .A(A[631]), .B(n395), .CI(
        C[631]), .CO(C[632]) );
  FA_15046 \FA_INST_0[1].FA_INST_1[120].FA_  ( .A(A[632]), .B(n394), .CI(
        C[632]), .CO(C[633]) );
  FA_15045 \FA_INST_0[1].FA_INST_1[121].FA_  ( .A(A[633]), .B(n393), .CI(
        C[633]), .CO(C[634]) );
  FA_15044 \FA_INST_0[1].FA_INST_1[122].FA_  ( .A(A[634]), .B(n392), .CI(
        C[634]), .CO(C[635]) );
  FA_15043 \FA_INST_0[1].FA_INST_1[123].FA_  ( .A(A[635]), .B(n391), .CI(
        C[635]), .CO(C[636]) );
  FA_15042 \FA_INST_0[1].FA_INST_1[124].FA_  ( .A(A[636]), .B(n390), .CI(
        C[636]), .CO(C[637]) );
  FA_15041 \FA_INST_0[1].FA_INST_1[125].FA_  ( .A(A[637]), .B(n389), .CI(
        C[637]), .CO(C[638]) );
  FA_15040 \FA_INST_0[1].FA_INST_1[126].FA_  ( .A(A[638]), .B(n388), .CI(
        C[638]), .CO(C[639]) );
  FA_15039 \FA_INST_0[1].FA_INST_1[127].FA_  ( .A(A[639]), .B(n387), .CI(
        C[639]), .CO(C[640]) );
  FA_15038 \FA_INST_0[1].FA_INST_1[128].FA_  ( .A(A[640]), .B(n386), .CI(
        C[640]), .CO(C[641]) );
  FA_15037 \FA_INST_0[1].FA_INST_1[129].FA_  ( .A(A[641]), .B(n385), .CI(
        C[641]), .CO(C[642]) );
  FA_15036 \FA_INST_0[1].FA_INST_1[130].FA_  ( .A(A[642]), .B(n384), .CI(
        C[642]), .CO(C[643]) );
  FA_15035 \FA_INST_0[1].FA_INST_1[131].FA_  ( .A(A[643]), .B(n383), .CI(
        C[643]), .CO(C[644]) );
  FA_15034 \FA_INST_0[1].FA_INST_1[132].FA_  ( .A(A[644]), .B(n382), .CI(
        C[644]), .CO(C[645]) );
  FA_15033 \FA_INST_0[1].FA_INST_1[133].FA_  ( .A(A[645]), .B(n381), .CI(
        C[645]), .CO(C[646]) );
  FA_15032 \FA_INST_0[1].FA_INST_1[134].FA_  ( .A(A[646]), .B(n380), .CI(
        C[646]), .CO(C[647]) );
  FA_15031 \FA_INST_0[1].FA_INST_1[135].FA_  ( .A(A[647]), .B(n379), .CI(
        C[647]), .CO(C[648]) );
  FA_15030 \FA_INST_0[1].FA_INST_1[136].FA_  ( .A(A[648]), .B(n378), .CI(
        C[648]), .CO(C[649]) );
  FA_15029 \FA_INST_0[1].FA_INST_1[137].FA_  ( .A(A[649]), .B(n377), .CI(
        C[649]), .CO(C[650]) );
  FA_15028 \FA_INST_0[1].FA_INST_1[138].FA_  ( .A(A[650]), .B(n376), .CI(
        C[650]), .CO(C[651]) );
  FA_15027 \FA_INST_0[1].FA_INST_1[139].FA_  ( .A(A[651]), .B(n375), .CI(
        C[651]), .CO(C[652]) );
  FA_15026 \FA_INST_0[1].FA_INST_1[140].FA_  ( .A(A[652]), .B(n374), .CI(
        C[652]), .CO(C[653]) );
  FA_15025 \FA_INST_0[1].FA_INST_1[141].FA_  ( .A(A[653]), .B(n373), .CI(
        C[653]), .CO(C[654]) );
  FA_15024 \FA_INST_0[1].FA_INST_1[142].FA_  ( .A(A[654]), .B(n372), .CI(
        C[654]), .CO(C[655]) );
  FA_15023 \FA_INST_0[1].FA_INST_1[143].FA_  ( .A(A[655]), .B(n371), .CI(
        C[655]), .CO(C[656]) );
  FA_15022 \FA_INST_0[1].FA_INST_1[144].FA_  ( .A(A[656]), .B(n370), .CI(
        C[656]), .CO(C[657]) );
  FA_15021 \FA_INST_0[1].FA_INST_1[145].FA_  ( .A(A[657]), .B(n369), .CI(
        C[657]), .CO(C[658]) );
  FA_15020 \FA_INST_0[1].FA_INST_1[146].FA_  ( .A(A[658]), .B(n368), .CI(
        C[658]), .CO(C[659]) );
  FA_15019 \FA_INST_0[1].FA_INST_1[147].FA_  ( .A(A[659]), .B(n367), .CI(
        C[659]), .CO(C[660]) );
  FA_15018 \FA_INST_0[1].FA_INST_1[148].FA_  ( .A(A[660]), .B(n366), .CI(
        C[660]), .CO(C[661]) );
  FA_15017 \FA_INST_0[1].FA_INST_1[149].FA_  ( .A(A[661]), .B(n365), .CI(
        C[661]), .CO(C[662]) );
  FA_15016 \FA_INST_0[1].FA_INST_1[150].FA_  ( .A(A[662]), .B(n364), .CI(
        C[662]), .CO(C[663]) );
  FA_15015 \FA_INST_0[1].FA_INST_1[151].FA_  ( .A(A[663]), .B(n363), .CI(
        C[663]), .CO(C[664]) );
  FA_15014 \FA_INST_0[1].FA_INST_1[152].FA_  ( .A(A[664]), .B(n362), .CI(
        C[664]), .CO(C[665]) );
  FA_15013 \FA_INST_0[1].FA_INST_1[153].FA_  ( .A(A[665]), .B(n361), .CI(
        C[665]), .CO(C[666]) );
  FA_15012 \FA_INST_0[1].FA_INST_1[154].FA_  ( .A(A[666]), .B(n360), .CI(
        C[666]), .CO(C[667]) );
  FA_15011 \FA_INST_0[1].FA_INST_1[155].FA_  ( .A(A[667]), .B(n359), .CI(
        C[667]), .CO(C[668]) );
  FA_15010 \FA_INST_0[1].FA_INST_1[156].FA_  ( .A(A[668]), .B(n358), .CI(
        C[668]), .CO(C[669]) );
  FA_15009 \FA_INST_0[1].FA_INST_1[157].FA_  ( .A(A[669]), .B(n357), .CI(
        C[669]), .CO(C[670]) );
  FA_15008 \FA_INST_0[1].FA_INST_1[158].FA_  ( .A(A[670]), .B(n356), .CI(
        C[670]), .CO(C[671]) );
  FA_15007 \FA_INST_0[1].FA_INST_1[159].FA_  ( .A(A[671]), .B(n355), .CI(
        C[671]), .CO(C[672]) );
  FA_15006 \FA_INST_0[1].FA_INST_1[160].FA_  ( .A(A[672]), .B(n354), .CI(
        C[672]), .CO(C[673]) );
  FA_15005 \FA_INST_0[1].FA_INST_1[161].FA_  ( .A(A[673]), .B(n353), .CI(
        C[673]), .CO(C[674]) );
  FA_15004 \FA_INST_0[1].FA_INST_1[162].FA_  ( .A(A[674]), .B(n352), .CI(
        C[674]), .CO(C[675]) );
  FA_15003 \FA_INST_0[1].FA_INST_1[163].FA_  ( .A(A[675]), .B(n351), .CI(
        C[675]), .CO(C[676]) );
  FA_15002 \FA_INST_0[1].FA_INST_1[164].FA_  ( .A(A[676]), .B(n350), .CI(
        C[676]), .CO(C[677]) );
  FA_15001 \FA_INST_0[1].FA_INST_1[165].FA_  ( .A(A[677]), .B(n349), .CI(
        C[677]), .CO(C[678]) );
  FA_15000 \FA_INST_0[1].FA_INST_1[166].FA_  ( .A(A[678]), .B(n348), .CI(
        C[678]), .CO(C[679]) );
  FA_14999 \FA_INST_0[1].FA_INST_1[167].FA_  ( .A(A[679]), .B(n347), .CI(
        C[679]), .CO(C[680]) );
  FA_14998 \FA_INST_0[1].FA_INST_1[168].FA_  ( .A(A[680]), .B(n346), .CI(
        C[680]), .CO(C[681]) );
  FA_14997 \FA_INST_0[1].FA_INST_1[169].FA_  ( .A(A[681]), .B(n345), .CI(
        C[681]), .CO(C[682]) );
  FA_14996 \FA_INST_0[1].FA_INST_1[170].FA_  ( .A(A[682]), .B(n344), .CI(
        C[682]), .CO(C[683]) );
  FA_14995 \FA_INST_0[1].FA_INST_1[171].FA_  ( .A(A[683]), .B(n343), .CI(
        C[683]), .CO(C[684]) );
  FA_14994 \FA_INST_0[1].FA_INST_1[172].FA_  ( .A(A[684]), .B(n342), .CI(
        C[684]), .CO(C[685]) );
  FA_14993 \FA_INST_0[1].FA_INST_1[173].FA_  ( .A(A[685]), .B(n341), .CI(
        C[685]), .CO(C[686]) );
  FA_14992 \FA_INST_0[1].FA_INST_1[174].FA_  ( .A(A[686]), .B(n340), .CI(
        C[686]), .CO(C[687]) );
  FA_14991 \FA_INST_0[1].FA_INST_1[175].FA_  ( .A(A[687]), .B(n339), .CI(
        C[687]), .CO(C[688]) );
  FA_14990 \FA_INST_0[1].FA_INST_1[176].FA_  ( .A(A[688]), .B(n338), .CI(
        C[688]), .CO(C[689]) );
  FA_14989 \FA_INST_0[1].FA_INST_1[177].FA_  ( .A(A[689]), .B(n337), .CI(
        C[689]), .CO(C[690]) );
  FA_14988 \FA_INST_0[1].FA_INST_1[178].FA_  ( .A(A[690]), .B(n336), .CI(
        C[690]), .CO(C[691]) );
  FA_14987 \FA_INST_0[1].FA_INST_1[179].FA_  ( .A(A[691]), .B(n335), .CI(
        C[691]), .CO(C[692]) );
  FA_14986 \FA_INST_0[1].FA_INST_1[180].FA_  ( .A(A[692]), .B(n334), .CI(
        C[692]), .CO(C[693]) );
  FA_14985 \FA_INST_0[1].FA_INST_1[181].FA_  ( .A(A[693]), .B(n333), .CI(
        C[693]), .CO(C[694]) );
  FA_14984 \FA_INST_0[1].FA_INST_1[182].FA_  ( .A(A[694]), .B(n332), .CI(
        C[694]), .CO(C[695]) );
  FA_14983 \FA_INST_0[1].FA_INST_1[183].FA_  ( .A(A[695]), .B(n331), .CI(
        C[695]), .CO(C[696]) );
  FA_14982 \FA_INST_0[1].FA_INST_1[184].FA_  ( .A(A[696]), .B(n330), .CI(
        C[696]), .CO(C[697]) );
  FA_14981 \FA_INST_0[1].FA_INST_1[185].FA_  ( .A(A[697]), .B(n329), .CI(
        C[697]), .CO(C[698]) );
  FA_14980 \FA_INST_0[1].FA_INST_1[186].FA_  ( .A(A[698]), .B(n328), .CI(
        C[698]), .CO(C[699]) );
  FA_14979 \FA_INST_0[1].FA_INST_1[187].FA_  ( .A(A[699]), .B(n327), .CI(
        C[699]), .CO(C[700]) );
  FA_14978 \FA_INST_0[1].FA_INST_1[188].FA_  ( .A(A[700]), .B(n326), .CI(
        C[700]), .CO(C[701]) );
  FA_14977 \FA_INST_0[1].FA_INST_1[189].FA_  ( .A(A[701]), .B(n325), .CI(
        C[701]), .CO(C[702]) );
  FA_14976 \FA_INST_0[1].FA_INST_1[190].FA_  ( .A(A[702]), .B(n324), .CI(
        C[702]), .CO(C[703]) );
  FA_14975 \FA_INST_0[1].FA_INST_1[191].FA_  ( .A(A[703]), .B(n323), .CI(
        C[703]), .CO(C[704]) );
  FA_14974 \FA_INST_0[1].FA_INST_1[192].FA_  ( .A(A[704]), .B(n322), .CI(
        C[704]), .CO(C[705]) );
  FA_14973 \FA_INST_0[1].FA_INST_1[193].FA_  ( .A(A[705]), .B(n321), .CI(
        C[705]), .CO(C[706]) );
  FA_14972 \FA_INST_0[1].FA_INST_1[194].FA_  ( .A(A[706]), .B(n320), .CI(
        C[706]), .CO(C[707]) );
  FA_14971 \FA_INST_0[1].FA_INST_1[195].FA_  ( .A(A[707]), .B(n319), .CI(
        C[707]), .CO(C[708]) );
  FA_14970 \FA_INST_0[1].FA_INST_1[196].FA_  ( .A(A[708]), .B(n318), .CI(
        C[708]), .CO(C[709]) );
  FA_14969 \FA_INST_0[1].FA_INST_1[197].FA_  ( .A(A[709]), .B(n317), .CI(
        C[709]), .CO(C[710]) );
  FA_14968 \FA_INST_0[1].FA_INST_1[198].FA_  ( .A(A[710]), .B(n316), .CI(
        C[710]), .CO(C[711]) );
  FA_14967 \FA_INST_0[1].FA_INST_1[199].FA_  ( .A(A[711]), .B(n315), .CI(
        C[711]), .CO(C[712]) );
  FA_14966 \FA_INST_0[1].FA_INST_1[200].FA_  ( .A(A[712]), .B(n314), .CI(
        C[712]), .CO(C[713]) );
  FA_14965 \FA_INST_0[1].FA_INST_1[201].FA_  ( .A(A[713]), .B(n313), .CI(
        C[713]), .CO(C[714]) );
  FA_14964 \FA_INST_0[1].FA_INST_1[202].FA_  ( .A(A[714]), .B(n312), .CI(
        C[714]), .CO(C[715]) );
  FA_14963 \FA_INST_0[1].FA_INST_1[203].FA_  ( .A(A[715]), .B(n311), .CI(
        C[715]), .CO(C[716]) );
  FA_14962 \FA_INST_0[1].FA_INST_1[204].FA_  ( .A(A[716]), .B(n310), .CI(
        C[716]), .CO(C[717]) );
  FA_14961 \FA_INST_0[1].FA_INST_1[205].FA_  ( .A(A[717]), .B(n309), .CI(
        C[717]), .CO(C[718]) );
  FA_14960 \FA_INST_0[1].FA_INST_1[206].FA_  ( .A(A[718]), .B(n308), .CI(
        C[718]), .CO(C[719]) );
  FA_14959 \FA_INST_0[1].FA_INST_1[207].FA_  ( .A(A[719]), .B(n307), .CI(
        C[719]), .CO(C[720]) );
  FA_14958 \FA_INST_0[1].FA_INST_1[208].FA_  ( .A(A[720]), .B(n306), .CI(
        C[720]), .CO(C[721]) );
  FA_14957 \FA_INST_0[1].FA_INST_1[209].FA_  ( .A(A[721]), .B(n305), .CI(
        C[721]), .CO(C[722]) );
  FA_14956 \FA_INST_0[1].FA_INST_1[210].FA_  ( .A(A[722]), .B(n304), .CI(
        C[722]), .CO(C[723]) );
  FA_14955 \FA_INST_0[1].FA_INST_1[211].FA_  ( .A(A[723]), .B(n303), .CI(
        C[723]), .CO(C[724]) );
  FA_14954 \FA_INST_0[1].FA_INST_1[212].FA_  ( .A(A[724]), .B(n302), .CI(
        C[724]), .CO(C[725]) );
  FA_14953 \FA_INST_0[1].FA_INST_1[213].FA_  ( .A(A[725]), .B(n301), .CI(
        C[725]), .CO(C[726]) );
  FA_14952 \FA_INST_0[1].FA_INST_1[214].FA_  ( .A(A[726]), .B(n300), .CI(
        C[726]), .CO(C[727]) );
  FA_14951 \FA_INST_0[1].FA_INST_1[215].FA_  ( .A(A[727]), .B(n299), .CI(
        C[727]), .CO(C[728]) );
  FA_14950 \FA_INST_0[1].FA_INST_1[216].FA_  ( .A(A[728]), .B(n298), .CI(
        C[728]), .CO(C[729]) );
  FA_14949 \FA_INST_0[1].FA_INST_1[217].FA_  ( .A(A[729]), .B(n297), .CI(
        C[729]), .CO(C[730]) );
  FA_14948 \FA_INST_0[1].FA_INST_1[218].FA_  ( .A(A[730]), .B(n296), .CI(
        C[730]), .CO(C[731]) );
  FA_14947 \FA_INST_0[1].FA_INST_1[219].FA_  ( .A(A[731]), .B(n295), .CI(
        C[731]), .CO(C[732]) );
  FA_14946 \FA_INST_0[1].FA_INST_1[220].FA_  ( .A(A[732]), .B(n294), .CI(
        C[732]), .CO(C[733]) );
  FA_14945 \FA_INST_0[1].FA_INST_1[221].FA_  ( .A(A[733]), .B(n293), .CI(
        C[733]), .CO(C[734]) );
  FA_14944 \FA_INST_0[1].FA_INST_1[222].FA_  ( .A(A[734]), .B(n292), .CI(
        C[734]), .CO(C[735]) );
  FA_14943 \FA_INST_0[1].FA_INST_1[223].FA_  ( .A(A[735]), .B(n291), .CI(
        C[735]), .CO(C[736]) );
  FA_14942 \FA_INST_0[1].FA_INST_1[224].FA_  ( .A(A[736]), .B(n290), .CI(
        C[736]), .CO(C[737]) );
  FA_14941 \FA_INST_0[1].FA_INST_1[225].FA_  ( .A(A[737]), .B(n289), .CI(
        C[737]), .CO(C[738]) );
  FA_14940 \FA_INST_0[1].FA_INST_1[226].FA_  ( .A(A[738]), .B(n288), .CI(
        C[738]), .CO(C[739]) );
  FA_14939 \FA_INST_0[1].FA_INST_1[227].FA_  ( .A(A[739]), .B(n287), .CI(
        C[739]), .CO(C[740]) );
  FA_14938 \FA_INST_0[1].FA_INST_1[228].FA_  ( .A(A[740]), .B(n286), .CI(
        C[740]), .CO(C[741]) );
  FA_14937 \FA_INST_0[1].FA_INST_1[229].FA_  ( .A(A[741]), .B(n285), .CI(
        C[741]), .CO(C[742]) );
  FA_14936 \FA_INST_0[1].FA_INST_1[230].FA_  ( .A(A[742]), .B(n284), .CI(
        C[742]), .CO(C[743]) );
  FA_14935 \FA_INST_0[1].FA_INST_1[231].FA_  ( .A(A[743]), .B(n283), .CI(
        C[743]), .CO(C[744]) );
  FA_14934 \FA_INST_0[1].FA_INST_1[232].FA_  ( .A(A[744]), .B(n282), .CI(
        C[744]), .CO(C[745]) );
  FA_14933 \FA_INST_0[1].FA_INST_1[233].FA_  ( .A(A[745]), .B(n281), .CI(
        C[745]), .CO(C[746]) );
  FA_14932 \FA_INST_0[1].FA_INST_1[234].FA_  ( .A(A[746]), .B(n280), .CI(
        C[746]), .CO(C[747]) );
  FA_14931 \FA_INST_0[1].FA_INST_1[235].FA_  ( .A(A[747]), .B(n279), .CI(
        C[747]), .CO(C[748]) );
  FA_14930 \FA_INST_0[1].FA_INST_1[236].FA_  ( .A(A[748]), .B(n278), .CI(
        C[748]), .CO(C[749]) );
  FA_14929 \FA_INST_0[1].FA_INST_1[237].FA_  ( .A(A[749]), .B(n277), .CI(
        C[749]), .CO(C[750]) );
  FA_14928 \FA_INST_0[1].FA_INST_1[238].FA_  ( .A(A[750]), .B(n276), .CI(
        C[750]), .CO(C[751]) );
  FA_14927 \FA_INST_0[1].FA_INST_1[239].FA_  ( .A(A[751]), .B(n275), .CI(
        C[751]), .CO(C[752]) );
  FA_14926 \FA_INST_0[1].FA_INST_1[240].FA_  ( .A(A[752]), .B(n274), .CI(
        C[752]), .CO(C[753]) );
  FA_14925 \FA_INST_0[1].FA_INST_1[241].FA_  ( .A(A[753]), .B(n273), .CI(
        C[753]), .CO(C[754]) );
  FA_14924 \FA_INST_0[1].FA_INST_1[242].FA_  ( .A(A[754]), .B(n272), .CI(
        C[754]), .CO(C[755]) );
  FA_14923 \FA_INST_0[1].FA_INST_1[243].FA_  ( .A(A[755]), .B(n271), .CI(
        C[755]), .CO(C[756]) );
  FA_14922 \FA_INST_0[1].FA_INST_1[244].FA_  ( .A(A[756]), .B(n270), .CI(
        C[756]), .CO(C[757]) );
  FA_14921 \FA_INST_0[1].FA_INST_1[245].FA_  ( .A(A[757]), .B(n269), .CI(
        C[757]), .CO(C[758]) );
  FA_14920 \FA_INST_0[1].FA_INST_1[246].FA_  ( .A(A[758]), .B(n268), .CI(
        C[758]), .CO(C[759]) );
  FA_14919 \FA_INST_0[1].FA_INST_1[247].FA_  ( .A(A[759]), .B(n267), .CI(
        C[759]), .CO(C[760]) );
  FA_14918 \FA_INST_0[1].FA_INST_1[248].FA_  ( .A(A[760]), .B(n266), .CI(
        C[760]), .CO(C[761]) );
  FA_14917 \FA_INST_0[1].FA_INST_1[249].FA_  ( .A(A[761]), .B(n265), .CI(
        C[761]), .CO(C[762]) );
  FA_14916 \FA_INST_0[1].FA_INST_1[250].FA_  ( .A(A[762]), .B(n264), .CI(
        C[762]), .CO(C[763]) );
  FA_14915 \FA_INST_0[1].FA_INST_1[251].FA_  ( .A(A[763]), .B(n263), .CI(
        C[763]), .CO(C[764]) );
  FA_14914 \FA_INST_0[1].FA_INST_1[252].FA_  ( .A(A[764]), .B(n262), .CI(
        C[764]), .CO(C[765]) );
  FA_14913 \FA_INST_0[1].FA_INST_1[253].FA_  ( .A(A[765]), .B(n261), .CI(
        C[765]), .CO(C[766]) );
  FA_14912 \FA_INST_0[1].FA_INST_1[254].FA_  ( .A(A[766]), .B(n260), .CI(
        C[766]), .CO(C[767]) );
  FA_14911 \FA_INST_0[1].FA_INST_1[255].FA_  ( .A(A[767]), .B(n259), .CI(
        C[767]), .CO(C[768]) );
  FA_14910 \FA_INST_0[1].FA_INST_1[256].FA_  ( .A(A[768]), .B(n258), .CI(
        C[768]), .CO(C[769]) );
  FA_14909 \FA_INST_0[1].FA_INST_1[257].FA_  ( .A(A[769]), .B(n257), .CI(
        C[769]), .CO(C[770]) );
  FA_14908 \FA_INST_0[1].FA_INST_1[258].FA_  ( .A(A[770]), .B(n256), .CI(
        C[770]), .CO(C[771]) );
  FA_14907 \FA_INST_0[1].FA_INST_1[259].FA_  ( .A(A[771]), .B(n255), .CI(
        C[771]), .CO(C[772]) );
  FA_14906 \FA_INST_0[1].FA_INST_1[260].FA_  ( .A(A[772]), .B(n254), .CI(
        C[772]), .CO(C[773]) );
  FA_14905 \FA_INST_0[1].FA_INST_1[261].FA_  ( .A(A[773]), .B(n253), .CI(
        C[773]), .CO(C[774]) );
  FA_14904 \FA_INST_0[1].FA_INST_1[262].FA_  ( .A(A[774]), .B(n252), .CI(
        C[774]), .CO(C[775]) );
  FA_14903 \FA_INST_0[1].FA_INST_1[263].FA_  ( .A(A[775]), .B(n251), .CI(
        C[775]), .CO(C[776]) );
  FA_14902 \FA_INST_0[1].FA_INST_1[264].FA_  ( .A(A[776]), .B(n250), .CI(
        C[776]), .CO(C[777]) );
  FA_14901 \FA_INST_0[1].FA_INST_1[265].FA_  ( .A(A[777]), .B(n249), .CI(
        C[777]), .CO(C[778]) );
  FA_14900 \FA_INST_0[1].FA_INST_1[266].FA_  ( .A(A[778]), .B(n248), .CI(
        C[778]), .CO(C[779]) );
  FA_14899 \FA_INST_0[1].FA_INST_1[267].FA_  ( .A(A[779]), .B(n247), .CI(
        C[779]), .CO(C[780]) );
  FA_14898 \FA_INST_0[1].FA_INST_1[268].FA_  ( .A(A[780]), .B(n246), .CI(
        C[780]), .CO(C[781]) );
  FA_14897 \FA_INST_0[1].FA_INST_1[269].FA_  ( .A(A[781]), .B(n245), .CI(
        C[781]), .CO(C[782]) );
  FA_14896 \FA_INST_0[1].FA_INST_1[270].FA_  ( .A(A[782]), .B(n244), .CI(
        C[782]), .CO(C[783]) );
  FA_14895 \FA_INST_0[1].FA_INST_1[271].FA_  ( .A(A[783]), .B(n243), .CI(
        C[783]), .CO(C[784]) );
  FA_14894 \FA_INST_0[1].FA_INST_1[272].FA_  ( .A(A[784]), .B(n242), .CI(
        C[784]), .CO(C[785]) );
  FA_14893 \FA_INST_0[1].FA_INST_1[273].FA_  ( .A(A[785]), .B(n241), .CI(
        C[785]), .CO(C[786]) );
  FA_14892 \FA_INST_0[1].FA_INST_1[274].FA_  ( .A(A[786]), .B(n240), .CI(
        C[786]), .CO(C[787]) );
  FA_14891 \FA_INST_0[1].FA_INST_1[275].FA_  ( .A(A[787]), .B(n239), .CI(
        C[787]), .CO(C[788]) );
  FA_14890 \FA_INST_0[1].FA_INST_1[276].FA_  ( .A(A[788]), .B(n238), .CI(
        C[788]), .CO(C[789]) );
  FA_14889 \FA_INST_0[1].FA_INST_1[277].FA_  ( .A(A[789]), .B(n237), .CI(
        C[789]), .CO(C[790]) );
  FA_14888 \FA_INST_0[1].FA_INST_1[278].FA_  ( .A(A[790]), .B(n236), .CI(
        C[790]), .CO(C[791]) );
  FA_14887 \FA_INST_0[1].FA_INST_1[279].FA_  ( .A(A[791]), .B(n235), .CI(
        C[791]), .CO(C[792]) );
  FA_14886 \FA_INST_0[1].FA_INST_1[280].FA_  ( .A(A[792]), .B(n234), .CI(
        C[792]), .CO(C[793]) );
  FA_14885 \FA_INST_0[1].FA_INST_1[281].FA_  ( .A(A[793]), .B(n233), .CI(
        C[793]), .CO(C[794]) );
  FA_14884 \FA_INST_0[1].FA_INST_1[282].FA_  ( .A(A[794]), .B(n232), .CI(
        C[794]), .CO(C[795]) );
  FA_14883 \FA_INST_0[1].FA_INST_1[283].FA_  ( .A(A[795]), .B(n231), .CI(
        C[795]), .CO(C[796]) );
  FA_14882 \FA_INST_0[1].FA_INST_1[284].FA_  ( .A(A[796]), .B(n230), .CI(
        C[796]), .CO(C[797]) );
  FA_14881 \FA_INST_0[1].FA_INST_1[285].FA_  ( .A(A[797]), .B(n229), .CI(
        C[797]), .CO(C[798]) );
  FA_14880 \FA_INST_0[1].FA_INST_1[286].FA_  ( .A(A[798]), .B(n228), .CI(
        C[798]), .CO(C[799]) );
  FA_14879 \FA_INST_0[1].FA_INST_1[287].FA_  ( .A(A[799]), .B(n227), .CI(
        C[799]), .CO(C[800]) );
  FA_14878 \FA_INST_0[1].FA_INST_1[288].FA_  ( .A(A[800]), .B(n226), .CI(
        C[800]), .CO(C[801]) );
  FA_14877 \FA_INST_0[1].FA_INST_1[289].FA_  ( .A(A[801]), .B(n225), .CI(
        C[801]), .CO(C[802]) );
  FA_14876 \FA_INST_0[1].FA_INST_1[290].FA_  ( .A(A[802]), .B(n224), .CI(
        C[802]), .CO(C[803]) );
  FA_14875 \FA_INST_0[1].FA_INST_1[291].FA_  ( .A(A[803]), .B(n223), .CI(
        C[803]), .CO(C[804]) );
  FA_14874 \FA_INST_0[1].FA_INST_1[292].FA_  ( .A(A[804]), .B(n222), .CI(
        C[804]), .CO(C[805]) );
  FA_14873 \FA_INST_0[1].FA_INST_1[293].FA_  ( .A(A[805]), .B(n221), .CI(
        C[805]), .CO(C[806]) );
  FA_14872 \FA_INST_0[1].FA_INST_1[294].FA_  ( .A(A[806]), .B(n220), .CI(
        C[806]), .CO(C[807]) );
  FA_14871 \FA_INST_0[1].FA_INST_1[295].FA_  ( .A(A[807]), .B(n219), .CI(
        C[807]), .CO(C[808]) );
  FA_14870 \FA_INST_0[1].FA_INST_1[296].FA_  ( .A(A[808]), .B(n218), .CI(
        C[808]), .CO(C[809]) );
  FA_14869 \FA_INST_0[1].FA_INST_1[297].FA_  ( .A(A[809]), .B(n217), .CI(
        C[809]), .CO(C[810]) );
  FA_14868 \FA_INST_0[1].FA_INST_1[298].FA_  ( .A(A[810]), .B(n216), .CI(
        C[810]), .CO(C[811]) );
  FA_14867 \FA_INST_0[1].FA_INST_1[299].FA_  ( .A(A[811]), .B(n215), .CI(
        C[811]), .CO(C[812]) );
  FA_14866 \FA_INST_0[1].FA_INST_1[300].FA_  ( .A(A[812]), .B(n214), .CI(
        C[812]), .CO(C[813]) );
  FA_14865 \FA_INST_0[1].FA_INST_1[301].FA_  ( .A(A[813]), .B(n213), .CI(
        C[813]), .CO(C[814]) );
  FA_14864 \FA_INST_0[1].FA_INST_1[302].FA_  ( .A(A[814]), .B(n212), .CI(
        C[814]), .CO(C[815]) );
  FA_14863 \FA_INST_0[1].FA_INST_1[303].FA_  ( .A(A[815]), .B(n211), .CI(
        C[815]), .CO(C[816]) );
  FA_14862 \FA_INST_0[1].FA_INST_1[304].FA_  ( .A(A[816]), .B(n210), .CI(
        C[816]), .CO(C[817]) );
  FA_14861 \FA_INST_0[1].FA_INST_1[305].FA_  ( .A(A[817]), .B(n209), .CI(
        C[817]), .CO(C[818]) );
  FA_14860 \FA_INST_0[1].FA_INST_1[306].FA_  ( .A(A[818]), .B(n208), .CI(
        C[818]), .CO(C[819]) );
  FA_14859 \FA_INST_0[1].FA_INST_1[307].FA_  ( .A(A[819]), .B(n207), .CI(
        C[819]), .CO(C[820]) );
  FA_14858 \FA_INST_0[1].FA_INST_1[308].FA_  ( .A(A[820]), .B(n206), .CI(
        C[820]), .CO(C[821]) );
  FA_14857 \FA_INST_0[1].FA_INST_1[309].FA_  ( .A(A[821]), .B(n205), .CI(
        C[821]), .CO(C[822]) );
  FA_14856 \FA_INST_0[1].FA_INST_1[310].FA_  ( .A(A[822]), .B(n204), .CI(
        C[822]), .CO(C[823]) );
  FA_14855 \FA_INST_0[1].FA_INST_1[311].FA_  ( .A(A[823]), .B(n203), .CI(
        C[823]), .CO(C[824]) );
  FA_14854 \FA_INST_0[1].FA_INST_1[312].FA_  ( .A(A[824]), .B(n202), .CI(
        C[824]), .CO(C[825]) );
  FA_14853 \FA_INST_0[1].FA_INST_1[313].FA_  ( .A(A[825]), .B(n201), .CI(
        C[825]), .CO(C[826]) );
  FA_14852 \FA_INST_0[1].FA_INST_1[314].FA_  ( .A(A[826]), .B(n200), .CI(
        C[826]), .CO(C[827]) );
  FA_14851 \FA_INST_0[1].FA_INST_1[315].FA_  ( .A(A[827]), .B(n199), .CI(
        C[827]), .CO(C[828]) );
  FA_14850 \FA_INST_0[1].FA_INST_1[316].FA_  ( .A(A[828]), .B(n198), .CI(
        C[828]), .CO(C[829]) );
  FA_14849 \FA_INST_0[1].FA_INST_1[317].FA_  ( .A(A[829]), .B(n197), .CI(
        C[829]), .CO(C[830]) );
  FA_14848 \FA_INST_0[1].FA_INST_1[318].FA_  ( .A(A[830]), .B(n196), .CI(
        C[830]), .CO(C[831]) );
  FA_14847 \FA_INST_0[1].FA_INST_1[319].FA_  ( .A(A[831]), .B(n195), .CI(
        C[831]), .CO(C[832]) );
  FA_14846 \FA_INST_0[1].FA_INST_1[320].FA_  ( .A(A[832]), .B(n194), .CI(
        C[832]), .CO(C[833]) );
  FA_14845 \FA_INST_0[1].FA_INST_1[321].FA_  ( .A(A[833]), .B(n193), .CI(
        C[833]), .CO(C[834]) );
  FA_14844 \FA_INST_0[1].FA_INST_1[322].FA_  ( .A(A[834]), .B(n192), .CI(
        C[834]), .CO(C[835]) );
  FA_14843 \FA_INST_0[1].FA_INST_1[323].FA_  ( .A(A[835]), .B(n191), .CI(
        C[835]), .CO(C[836]) );
  FA_14842 \FA_INST_0[1].FA_INST_1[324].FA_  ( .A(A[836]), .B(n190), .CI(
        C[836]), .CO(C[837]) );
  FA_14841 \FA_INST_0[1].FA_INST_1[325].FA_  ( .A(A[837]), .B(n189), .CI(
        C[837]), .CO(C[838]) );
  FA_14840 \FA_INST_0[1].FA_INST_1[326].FA_  ( .A(A[838]), .B(n188), .CI(
        C[838]), .CO(C[839]) );
  FA_14839 \FA_INST_0[1].FA_INST_1[327].FA_  ( .A(A[839]), .B(n187), .CI(
        C[839]), .CO(C[840]) );
  FA_14838 \FA_INST_0[1].FA_INST_1[328].FA_  ( .A(A[840]), .B(n186), .CI(
        C[840]), .CO(C[841]) );
  FA_14837 \FA_INST_0[1].FA_INST_1[329].FA_  ( .A(A[841]), .B(n185), .CI(
        C[841]), .CO(C[842]) );
  FA_14836 \FA_INST_0[1].FA_INST_1[330].FA_  ( .A(A[842]), .B(n184), .CI(
        C[842]), .CO(C[843]) );
  FA_14835 \FA_INST_0[1].FA_INST_1[331].FA_  ( .A(A[843]), .B(n183), .CI(
        C[843]), .CO(C[844]) );
  FA_14834 \FA_INST_0[1].FA_INST_1[332].FA_  ( .A(A[844]), .B(n182), .CI(
        C[844]), .CO(C[845]) );
  FA_14833 \FA_INST_0[1].FA_INST_1[333].FA_  ( .A(A[845]), .B(n181), .CI(
        C[845]), .CO(C[846]) );
  FA_14832 \FA_INST_0[1].FA_INST_1[334].FA_  ( .A(A[846]), .B(n180), .CI(
        C[846]), .CO(C[847]) );
  FA_14831 \FA_INST_0[1].FA_INST_1[335].FA_  ( .A(A[847]), .B(n179), .CI(
        C[847]), .CO(C[848]) );
  FA_14830 \FA_INST_0[1].FA_INST_1[336].FA_  ( .A(A[848]), .B(n178), .CI(
        C[848]), .CO(C[849]) );
  FA_14829 \FA_INST_0[1].FA_INST_1[337].FA_  ( .A(A[849]), .B(n177), .CI(
        C[849]), .CO(C[850]) );
  FA_14828 \FA_INST_0[1].FA_INST_1[338].FA_  ( .A(A[850]), .B(n176), .CI(
        C[850]), .CO(C[851]) );
  FA_14827 \FA_INST_0[1].FA_INST_1[339].FA_  ( .A(A[851]), .B(n175), .CI(
        C[851]), .CO(C[852]) );
  FA_14826 \FA_INST_0[1].FA_INST_1[340].FA_  ( .A(A[852]), .B(n174), .CI(
        C[852]), .CO(C[853]) );
  FA_14825 \FA_INST_0[1].FA_INST_1[341].FA_  ( .A(A[853]), .B(n173), .CI(
        C[853]), .CO(C[854]) );
  FA_14824 \FA_INST_0[1].FA_INST_1[342].FA_  ( .A(A[854]), .B(n172), .CI(
        C[854]), .CO(C[855]) );
  FA_14823 \FA_INST_0[1].FA_INST_1[343].FA_  ( .A(A[855]), .B(n171), .CI(
        C[855]), .CO(C[856]) );
  FA_14822 \FA_INST_0[1].FA_INST_1[344].FA_  ( .A(A[856]), .B(n170), .CI(
        C[856]), .CO(C[857]) );
  FA_14821 \FA_INST_0[1].FA_INST_1[345].FA_  ( .A(A[857]), .B(n169), .CI(
        C[857]), .CO(C[858]) );
  FA_14820 \FA_INST_0[1].FA_INST_1[346].FA_  ( .A(A[858]), .B(n168), .CI(
        C[858]), .CO(C[859]) );
  FA_14819 \FA_INST_0[1].FA_INST_1[347].FA_  ( .A(A[859]), .B(n167), .CI(
        C[859]), .CO(C[860]) );
  FA_14818 \FA_INST_0[1].FA_INST_1[348].FA_  ( .A(A[860]), .B(n166), .CI(
        C[860]), .CO(C[861]) );
  FA_14817 \FA_INST_0[1].FA_INST_1[349].FA_  ( .A(A[861]), .B(n165), .CI(
        C[861]), .CO(C[862]) );
  FA_14816 \FA_INST_0[1].FA_INST_1[350].FA_  ( .A(A[862]), .B(n164), .CI(
        C[862]), .CO(C[863]) );
  FA_14815 \FA_INST_0[1].FA_INST_1[351].FA_  ( .A(A[863]), .B(n163), .CI(
        C[863]), .CO(C[864]) );
  FA_14814 \FA_INST_0[1].FA_INST_1[352].FA_  ( .A(A[864]), .B(n162), .CI(
        C[864]), .CO(C[865]) );
  FA_14813 \FA_INST_0[1].FA_INST_1[353].FA_  ( .A(A[865]), .B(n161), .CI(
        C[865]), .CO(C[866]) );
  FA_14812 \FA_INST_0[1].FA_INST_1[354].FA_  ( .A(A[866]), .B(n160), .CI(
        C[866]), .CO(C[867]) );
  FA_14811 \FA_INST_0[1].FA_INST_1[355].FA_  ( .A(A[867]), .B(n159), .CI(
        C[867]), .CO(C[868]) );
  FA_14810 \FA_INST_0[1].FA_INST_1[356].FA_  ( .A(A[868]), .B(n158), .CI(
        C[868]), .CO(C[869]) );
  FA_14809 \FA_INST_0[1].FA_INST_1[357].FA_  ( .A(A[869]), .B(n157), .CI(
        C[869]), .CO(C[870]) );
  FA_14808 \FA_INST_0[1].FA_INST_1[358].FA_  ( .A(A[870]), .B(n156), .CI(
        C[870]), .CO(C[871]) );
  FA_14807 \FA_INST_0[1].FA_INST_1[359].FA_  ( .A(A[871]), .B(n155), .CI(
        C[871]), .CO(C[872]) );
  FA_14806 \FA_INST_0[1].FA_INST_1[360].FA_  ( .A(A[872]), .B(n154), .CI(
        C[872]), .CO(C[873]) );
  FA_14805 \FA_INST_0[1].FA_INST_1[361].FA_  ( .A(A[873]), .B(n153), .CI(
        C[873]), .CO(C[874]) );
  FA_14804 \FA_INST_0[1].FA_INST_1[362].FA_  ( .A(A[874]), .B(n152), .CI(
        C[874]), .CO(C[875]) );
  FA_14803 \FA_INST_0[1].FA_INST_1[363].FA_  ( .A(A[875]), .B(n151), .CI(
        C[875]), .CO(C[876]) );
  FA_14802 \FA_INST_0[1].FA_INST_1[364].FA_  ( .A(A[876]), .B(n150), .CI(
        C[876]), .CO(C[877]) );
  FA_14801 \FA_INST_0[1].FA_INST_1[365].FA_  ( .A(A[877]), .B(n149), .CI(
        C[877]), .CO(C[878]) );
  FA_14800 \FA_INST_0[1].FA_INST_1[366].FA_  ( .A(A[878]), .B(n148), .CI(
        C[878]), .CO(C[879]) );
  FA_14799 \FA_INST_0[1].FA_INST_1[367].FA_  ( .A(A[879]), .B(n147), .CI(
        C[879]), .CO(C[880]) );
  FA_14798 \FA_INST_0[1].FA_INST_1[368].FA_  ( .A(A[880]), .B(n146), .CI(
        C[880]), .CO(C[881]) );
  FA_14797 \FA_INST_0[1].FA_INST_1[369].FA_  ( .A(A[881]), .B(n145), .CI(
        C[881]), .CO(C[882]) );
  FA_14796 \FA_INST_0[1].FA_INST_1[370].FA_  ( .A(A[882]), .B(n144), .CI(
        C[882]), .CO(C[883]) );
  FA_14795 \FA_INST_0[1].FA_INST_1[371].FA_  ( .A(A[883]), .B(n143), .CI(
        C[883]), .CO(C[884]) );
  FA_14794 \FA_INST_0[1].FA_INST_1[372].FA_  ( .A(A[884]), .B(n142), .CI(
        C[884]), .CO(C[885]) );
  FA_14793 \FA_INST_0[1].FA_INST_1[373].FA_  ( .A(A[885]), .B(n141), .CI(
        C[885]), .CO(C[886]) );
  FA_14792 \FA_INST_0[1].FA_INST_1[374].FA_  ( .A(A[886]), .B(n140), .CI(
        C[886]), .CO(C[887]) );
  FA_14791 \FA_INST_0[1].FA_INST_1[375].FA_  ( .A(A[887]), .B(n139), .CI(
        C[887]), .CO(C[888]) );
  FA_14790 \FA_INST_0[1].FA_INST_1[376].FA_  ( .A(A[888]), .B(n138), .CI(
        C[888]), .CO(C[889]) );
  FA_14789 \FA_INST_0[1].FA_INST_1[377].FA_  ( .A(A[889]), .B(n137), .CI(
        C[889]), .CO(C[890]) );
  FA_14788 \FA_INST_0[1].FA_INST_1[378].FA_  ( .A(A[890]), .B(n136), .CI(
        C[890]), .CO(C[891]) );
  FA_14787 \FA_INST_0[1].FA_INST_1[379].FA_  ( .A(A[891]), .B(n135), .CI(
        C[891]), .CO(C[892]) );
  FA_14786 \FA_INST_0[1].FA_INST_1[380].FA_  ( .A(A[892]), .B(n134), .CI(
        C[892]), .CO(C[893]) );
  FA_14785 \FA_INST_0[1].FA_INST_1[381].FA_  ( .A(A[893]), .B(n133), .CI(
        C[893]), .CO(C[894]) );
  FA_14784 \FA_INST_0[1].FA_INST_1[382].FA_  ( .A(A[894]), .B(n132), .CI(
        C[894]), .CO(C[895]) );
  FA_14783 \FA_INST_0[1].FA_INST_1[383].FA_  ( .A(A[895]), .B(n131), .CI(
        C[895]), .CO(C[896]) );
  FA_14782 \FA_INST_0[1].FA_INST_1[384].FA_  ( .A(A[896]), .B(n130), .CI(
        C[896]), .CO(C[897]) );
  FA_14781 \FA_INST_0[1].FA_INST_1[385].FA_  ( .A(A[897]), .B(n129), .CI(
        C[897]), .CO(C[898]) );
  FA_14780 \FA_INST_0[1].FA_INST_1[386].FA_  ( .A(A[898]), .B(n128), .CI(
        C[898]), .CO(C[899]) );
  FA_14779 \FA_INST_0[1].FA_INST_1[387].FA_  ( .A(A[899]), .B(n127), .CI(
        C[899]), .CO(C[900]) );
  FA_14778 \FA_INST_0[1].FA_INST_1[388].FA_  ( .A(A[900]), .B(n126), .CI(
        C[900]), .CO(C[901]) );
  FA_14777 \FA_INST_0[1].FA_INST_1[389].FA_  ( .A(A[901]), .B(n125), .CI(
        C[901]), .CO(C[902]) );
  FA_14776 \FA_INST_0[1].FA_INST_1[390].FA_  ( .A(A[902]), .B(n124), .CI(
        C[902]), .CO(C[903]) );
  FA_14775 \FA_INST_0[1].FA_INST_1[391].FA_  ( .A(A[903]), .B(n123), .CI(
        C[903]), .CO(C[904]) );
  FA_14774 \FA_INST_0[1].FA_INST_1[392].FA_  ( .A(A[904]), .B(n122), .CI(
        C[904]), .CO(C[905]) );
  FA_14773 \FA_INST_0[1].FA_INST_1[393].FA_  ( .A(A[905]), .B(n121), .CI(
        C[905]), .CO(C[906]) );
  FA_14772 \FA_INST_0[1].FA_INST_1[394].FA_  ( .A(A[906]), .B(n120), .CI(
        C[906]), .CO(C[907]) );
  FA_14771 \FA_INST_0[1].FA_INST_1[395].FA_  ( .A(A[907]), .B(n119), .CI(
        C[907]), .CO(C[908]) );
  FA_14770 \FA_INST_0[1].FA_INST_1[396].FA_  ( .A(A[908]), .B(n118), .CI(
        C[908]), .CO(C[909]) );
  FA_14769 \FA_INST_0[1].FA_INST_1[397].FA_  ( .A(A[909]), .B(n117), .CI(
        C[909]), .CO(C[910]) );
  FA_14768 \FA_INST_0[1].FA_INST_1[398].FA_  ( .A(A[910]), .B(n116), .CI(
        C[910]), .CO(C[911]) );
  FA_14767 \FA_INST_0[1].FA_INST_1[399].FA_  ( .A(A[911]), .B(n115), .CI(
        C[911]), .CO(C[912]) );
  FA_14766 \FA_INST_0[1].FA_INST_1[400].FA_  ( .A(A[912]), .B(n114), .CI(
        C[912]), .CO(C[913]) );
  FA_14765 \FA_INST_0[1].FA_INST_1[401].FA_  ( .A(A[913]), .B(n113), .CI(
        C[913]), .CO(C[914]) );
  FA_14764 \FA_INST_0[1].FA_INST_1[402].FA_  ( .A(A[914]), .B(n112), .CI(
        C[914]), .CO(C[915]) );
  FA_14763 \FA_INST_0[1].FA_INST_1[403].FA_  ( .A(A[915]), .B(n111), .CI(
        C[915]), .CO(C[916]) );
  FA_14762 \FA_INST_0[1].FA_INST_1[404].FA_  ( .A(A[916]), .B(n110), .CI(
        C[916]), .CO(C[917]) );
  FA_14761 \FA_INST_0[1].FA_INST_1[405].FA_  ( .A(A[917]), .B(n109), .CI(
        C[917]), .CO(C[918]) );
  FA_14760 \FA_INST_0[1].FA_INST_1[406].FA_  ( .A(A[918]), .B(n108), .CI(
        C[918]), .CO(C[919]) );
  FA_14759 \FA_INST_0[1].FA_INST_1[407].FA_  ( .A(A[919]), .B(n107), .CI(
        C[919]), .CO(C[920]) );
  FA_14758 \FA_INST_0[1].FA_INST_1[408].FA_  ( .A(A[920]), .B(n106), .CI(
        C[920]), .CO(C[921]) );
  FA_14757 \FA_INST_0[1].FA_INST_1[409].FA_  ( .A(A[921]), .B(n105), .CI(
        C[921]), .CO(C[922]) );
  FA_14756 \FA_INST_0[1].FA_INST_1[410].FA_  ( .A(A[922]), .B(n104), .CI(
        C[922]), .CO(C[923]) );
  FA_14755 \FA_INST_0[1].FA_INST_1[411].FA_  ( .A(A[923]), .B(n103), .CI(
        C[923]), .CO(C[924]) );
  FA_14754 \FA_INST_0[1].FA_INST_1[412].FA_  ( .A(A[924]), .B(n102), .CI(
        C[924]), .CO(C[925]) );
  FA_14753 \FA_INST_0[1].FA_INST_1[413].FA_  ( .A(A[925]), .B(n101), .CI(
        C[925]), .CO(C[926]) );
  FA_14752 \FA_INST_0[1].FA_INST_1[414].FA_  ( .A(A[926]), .B(n100), .CI(
        C[926]), .CO(C[927]) );
  FA_14751 \FA_INST_0[1].FA_INST_1[415].FA_  ( .A(A[927]), .B(n99), .CI(C[927]), .CO(C[928]) );
  FA_14750 \FA_INST_0[1].FA_INST_1[416].FA_  ( .A(A[928]), .B(n98), .CI(C[928]), .CO(C[929]) );
  FA_14749 \FA_INST_0[1].FA_INST_1[417].FA_  ( .A(A[929]), .B(n97), .CI(C[929]), .CO(C[930]) );
  FA_14748 \FA_INST_0[1].FA_INST_1[418].FA_  ( .A(A[930]), .B(n96), .CI(C[930]), .CO(C[931]) );
  FA_14747 \FA_INST_0[1].FA_INST_1[419].FA_  ( .A(A[931]), .B(n95), .CI(C[931]), .CO(C[932]) );
  FA_14746 \FA_INST_0[1].FA_INST_1[420].FA_  ( .A(A[932]), .B(n94), .CI(C[932]), .CO(C[933]) );
  FA_14745 \FA_INST_0[1].FA_INST_1[421].FA_  ( .A(A[933]), .B(n93), .CI(C[933]), .CO(C[934]) );
  FA_14744 \FA_INST_0[1].FA_INST_1[422].FA_  ( .A(A[934]), .B(n92), .CI(C[934]), .CO(C[935]) );
  FA_14743 \FA_INST_0[1].FA_INST_1[423].FA_  ( .A(A[935]), .B(n91), .CI(C[935]), .CO(C[936]) );
  FA_14742 \FA_INST_0[1].FA_INST_1[424].FA_  ( .A(A[936]), .B(n90), .CI(C[936]), .CO(C[937]) );
  FA_14741 \FA_INST_0[1].FA_INST_1[425].FA_  ( .A(A[937]), .B(n89), .CI(C[937]), .CO(C[938]) );
  FA_14740 \FA_INST_0[1].FA_INST_1[426].FA_  ( .A(A[938]), .B(n88), .CI(C[938]), .CO(C[939]) );
  FA_14739 \FA_INST_0[1].FA_INST_1[427].FA_  ( .A(A[939]), .B(n87), .CI(C[939]), .CO(C[940]) );
  FA_14738 \FA_INST_0[1].FA_INST_1[428].FA_  ( .A(A[940]), .B(n86), .CI(C[940]), .CO(C[941]) );
  FA_14737 \FA_INST_0[1].FA_INST_1[429].FA_  ( .A(A[941]), .B(n85), .CI(C[941]), .CO(C[942]) );
  FA_14736 \FA_INST_0[1].FA_INST_1[430].FA_  ( .A(A[942]), .B(n84), .CI(C[942]), .CO(C[943]) );
  FA_14735 \FA_INST_0[1].FA_INST_1[431].FA_  ( .A(A[943]), .B(n83), .CI(C[943]), .CO(C[944]) );
  FA_14734 \FA_INST_0[1].FA_INST_1[432].FA_  ( .A(A[944]), .B(n82), .CI(C[944]), .CO(C[945]) );
  FA_14733 \FA_INST_0[1].FA_INST_1[433].FA_  ( .A(A[945]), .B(n81), .CI(C[945]), .CO(C[946]) );
  FA_14732 \FA_INST_0[1].FA_INST_1[434].FA_  ( .A(A[946]), .B(n80), .CI(C[946]), .CO(C[947]) );
  FA_14731 \FA_INST_0[1].FA_INST_1[435].FA_  ( .A(A[947]), .B(n79), .CI(C[947]), .CO(C[948]) );
  FA_14730 \FA_INST_0[1].FA_INST_1[436].FA_  ( .A(A[948]), .B(n78), .CI(C[948]), .CO(C[949]) );
  FA_14729 \FA_INST_0[1].FA_INST_1[437].FA_  ( .A(A[949]), .B(n77), .CI(C[949]), .CO(C[950]) );
  FA_14728 \FA_INST_0[1].FA_INST_1[438].FA_  ( .A(A[950]), .B(n76), .CI(C[950]), .CO(C[951]) );
  FA_14727 \FA_INST_0[1].FA_INST_1[439].FA_  ( .A(A[951]), .B(n75), .CI(C[951]), .CO(C[952]) );
  FA_14726 \FA_INST_0[1].FA_INST_1[440].FA_  ( .A(A[952]), .B(n74), .CI(C[952]), .CO(C[953]) );
  FA_14725 \FA_INST_0[1].FA_INST_1[441].FA_  ( .A(A[953]), .B(n73), .CI(C[953]), .CO(C[954]) );
  FA_14724 \FA_INST_0[1].FA_INST_1[442].FA_  ( .A(A[954]), .B(n72), .CI(C[954]), .CO(C[955]) );
  FA_14723 \FA_INST_0[1].FA_INST_1[443].FA_  ( .A(A[955]), .B(n71), .CI(C[955]), .CO(C[956]) );
  FA_14722 \FA_INST_0[1].FA_INST_1[444].FA_  ( .A(A[956]), .B(n70), .CI(C[956]), .CO(C[957]) );
  FA_14721 \FA_INST_0[1].FA_INST_1[445].FA_  ( .A(A[957]), .B(n69), .CI(C[957]), .CO(C[958]) );
  FA_14720 \FA_INST_0[1].FA_INST_1[446].FA_  ( .A(A[958]), .B(n68), .CI(C[958]), .CO(C[959]) );
  FA_14719 \FA_INST_0[1].FA_INST_1[447].FA_  ( .A(A[959]), .B(n67), .CI(C[959]), .CO(C[960]) );
  FA_14718 \FA_INST_0[1].FA_INST_1[448].FA_  ( .A(A[960]), .B(n66), .CI(C[960]), .CO(C[961]) );
  FA_14717 \FA_INST_0[1].FA_INST_1[449].FA_  ( .A(A[961]), .B(n65), .CI(C[961]), .CO(C[962]) );
  FA_14716 \FA_INST_0[1].FA_INST_1[450].FA_  ( .A(A[962]), .B(n64), .CI(C[962]), .CO(C[963]) );
  FA_14715 \FA_INST_0[1].FA_INST_1[451].FA_  ( .A(A[963]), .B(n63), .CI(C[963]), .CO(C[964]) );
  FA_14714 \FA_INST_0[1].FA_INST_1[452].FA_  ( .A(A[964]), .B(n62), .CI(C[964]), .CO(C[965]) );
  FA_14713 \FA_INST_0[1].FA_INST_1[453].FA_  ( .A(A[965]), .B(n61), .CI(C[965]), .CO(C[966]) );
  FA_14712 \FA_INST_0[1].FA_INST_1[454].FA_  ( .A(A[966]), .B(n60), .CI(C[966]), .CO(C[967]) );
  FA_14711 \FA_INST_0[1].FA_INST_1[455].FA_  ( .A(A[967]), .B(n59), .CI(C[967]), .CO(C[968]) );
  FA_14710 \FA_INST_0[1].FA_INST_1[456].FA_  ( .A(A[968]), .B(n58), .CI(C[968]), .CO(C[969]) );
  FA_14709 \FA_INST_0[1].FA_INST_1[457].FA_  ( .A(A[969]), .B(n57), .CI(C[969]), .CO(C[970]) );
  FA_14708 \FA_INST_0[1].FA_INST_1[458].FA_  ( .A(A[970]), .B(n56), .CI(C[970]), .CO(C[971]) );
  FA_14707 \FA_INST_0[1].FA_INST_1[459].FA_  ( .A(A[971]), .B(n55), .CI(C[971]), .CO(C[972]) );
  FA_14706 \FA_INST_0[1].FA_INST_1[460].FA_  ( .A(A[972]), .B(n54), .CI(C[972]), .CO(C[973]) );
  FA_14705 \FA_INST_0[1].FA_INST_1[461].FA_  ( .A(A[973]), .B(n53), .CI(C[973]), .CO(C[974]) );
  FA_14704 \FA_INST_0[1].FA_INST_1[462].FA_  ( .A(A[974]), .B(n52), .CI(C[974]), .CO(C[975]) );
  FA_14703 \FA_INST_0[1].FA_INST_1[463].FA_  ( .A(A[975]), .B(n51), .CI(C[975]), .CO(C[976]) );
  FA_14702 \FA_INST_0[1].FA_INST_1[464].FA_  ( .A(A[976]), .B(n50), .CI(C[976]), .CO(C[977]) );
  FA_14701 \FA_INST_0[1].FA_INST_1[465].FA_  ( .A(A[977]), .B(n49), .CI(C[977]), .CO(C[978]) );
  FA_14700 \FA_INST_0[1].FA_INST_1[466].FA_  ( .A(A[978]), .B(n48), .CI(C[978]), .CO(C[979]) );
  FA_14699 \FA_INST_0[1].FA_INST_1[467].FA_  ( .A(A[979]), .B(n47), .CI(C[979]), .CO(C[980]) );
  FA_14698 \FA_INST_0[1].FA_INST_1[468].FA_  ( .A(A[980]), .B(n46), .CI(C[980]), .CO(C[981]) );
  FA_14697 \FA_INST_0[1].FA_INST_1[469].FA_  ( .A(A[981]), .B(n45), .CI(C[981]), .CO(C[982]) );
  FA_14696 \FA_INST_0[1].FA_INST_1[470].FA_  ( .A(A[982]), .B(n44), .CI(C[982]), .CO(C[983]) );
  FA_14695 \FA_INST_0[1].FA_INST_1[471].FA_  ( .A(A[983]), .B(n43), .CI(C[983]), .CO(C[984]) );
  FA_14694 \FA_INST_0[1].FA_INST_1[472].FA_  ( .A(A[984]), .B(n42), .CI(C[984]), .CO(C[985]) );
  FA_14693 \FA_INST_0[1].FA_INST_1[473].FA_  ( .A(A[985]), .B(n41), .CI(C[985]), .CO(C[986]) );
  FA_14692 \FA_INST_0[1].FA_INST_1[474].FA_  ( .A(A[986]), .B(n40), .CI(C[986]), .CO(C[987]) );
  FA_14691 \FA_INST_0[1].FA_INST_1[475].FA_  ( .A(A[987]), .B(n39), .CI(C[987]), .CO(C[988]) );
  FA_14690 \FA_INST_0[1].FA_INST_1[476].FA_  ( .A(A[988]), .B(n38), .CI(C[988]), .CO(C[989]) );
  FA_14689 \FA_INST_0[1].FA_INST_1[477].FA_  ( .A(A[989]), .B(n37), .CI(C[989]), .CO(C[990]) );
  FA_14688 \FA_INST_0[1].FA_INST_1[478].FA_  ( .A(A[990]), .B(n36), .CI(C[990]), .CO(C[991]) );
  FA_14687 \FA_INST_0[1].FA_INST_1[479].FA_  ( .A(A[991]), .B(n35), .CI(C[991]), .CO(C[992]) );
  FA_14686 \FA_INST_0[1].FA_INST_1[480].FA_  ( .A(A[992]), .B(n34), .CI(C[992]), .CO(C[993]) );
  FA_14685 \FA_INST_0[1].FA_INST_1[481].FA_  ( .A(A[993]), .B(n33), .CI(C[993]), .CO(C[994]) );
  FA_14684 \FA_INST_0[1].FA_INST_1[482].FA_  ( .A(A[994]), .B(n32), .CI(C[994]), .CO(C[995]) );
  FA_14683 \FA_INST_0[1].FA_INST_1[483].FA_  ( .A(A[995]), .B(n31), .CI(C[995]), .CO(C[996]) );
  FA_14682 \FA_INST_0[1].FA_INST_1[484].FA_  ( .A(A[996]), .B(n30), .CI(C[996]), .CO(C[997]) );
  FA_14681 \FA_INST_0[1].FA_INST_1[485].FA_  ( .A(A[997]), .B(n29), .CI(C[997]), .CO(C[998]) );
  FA_14680 \FA_INST_0[1].FA_INST_1[486].FA_  ( .A(A[998]), .B(n28), .CI(C[998]), .CO(C[999]) );
  FA_14679 \FA_INST_0[1].FA_INST_1[487].FA_  ( .A(A[999]), .B(n27), .CI(C[999]), .CO(C[1000]) );
  FA_14678 \FA_INST_0[1].FA_INST_1[488].FA_  ( .A(A[1000]), .B(n26), .CI(
        C[1000]), .CO(C[1001]) );
  FA_14677 \FA_INST_0[1].FA_INST_1[489].FA_  ( .A(A[1001]), .B(n25), .CI(
        C[1001]), .CO(C[1002]) );
  FA_14676 \FA_INST_0[1].FA_INST_1[490].FA_  ( .A(A[1002]), .B(n24), .CI(
        C[1002]), .CO(C[1003]) );
  FA_14675 \FA_INST_0[1].FA_INST_1[491].FA_  ( .A(A[1003]), .B(n23), .CI(
        C[1003]), .CO(C[1004]) );
  FA_14674 \FA_INST_0[1].FA_INST_1[492].FA_  ( .A(A[1004]), .B(n22), .CI(
        C[1004]), .CO(C[1005]) );
  FA_14673 \FA_INST_0[1].FA_INST_1[493].FA_  ( .A(A[1005]), .B(n21), .CI(
        C[1005]), .CO(C[1006]) );
  FA_14672 \FA_INST_0[1].FA_INST_1[494].FA_  ( .A(A[1006]), .B(n20), .CI(
        C[1006]), .CO(C[1007]) );
  FA_14671 \FA_INST_0[1].FA_INST_1[495].FA_  ( .A(A[1007]), .B(n19), .CI(
        C[1007]), .CO(C[1008]) );
  FA_14670 \FA_INST_0[1].FA_INST_1[496].FA_  ( .A(A[1008]), .B(n18), .CI(
        C[1008]), .CO(C[1009]) );
  FA_14669 \FA_INST_0[1].FA_INST_1[497].FA_  ( .A(A[1009]), .B(n17), .CI(
        C[1009]), .CO(C[1010]) );
  FA_14668 \FA_INST_0[1].FA_INST_1[498].FA_  ( .A(A[1010]), .B(n16), .CI(
        C[1010]), .CO(C[1011]) );
  FA_14667 \FA_INST_0[1].FA_INST_1[499].FA_  ( .A(A[1011]), .B(n15), .CI(
        C[1011]), .CO(C[1012]) );
  FA_14666 \FA_INST_0[1].FA_INST_1[500].FA_  ( .A(A[1012]), .B(n14), .CI(
        C[1012]), .CO(C[1013]) );
  FA_14665 \FA_INST_0[1].FA_INST_1[501].FA_  ( .A(A[1013]), .B(n13), .CI(
        C[1013]), .CO(C[1014]) );
  FA_14664 \FA_INST_0[1].FA_INST_1[502].FA_  ( .A(A[1014]), .B(n12), .CI(
        C[1014]), .CO(C[1015]) );
  FA_14663 \FA_INST_0[1].FA_INST_1[503].FA_  ( .A(A[1015]), .B(n11), .CI(
        C[1015]), .CO(C[1016]) );
  FA_14662 \FA_INST_0[1].FA_INST_1[504].FA_  ( .A(A[1016]), .B(n10), .CI(
        C[1016]), .CO(C[1017]) );
  FA_14661 \FA_INST_0[1].FA_INST_1[505].FA_  ( .A(A[1017]), .B(n9), .CI(
        C[1017]), .CO(C[1018]) );
  FA_14660 \FA_INST_0[1].FA_INST_1[506].FA_  ( .A(A[1018]), .B(n8), .CI(
        C[1018]), .CO(C[1019]) );
  FA_14659 \FA_INST_0[1].FA_INST_1[507].FA_  ( .A(A[1019]), .B(n7), .CI(
        C[1019]), .CO(C[1020]) );
  FA_14658 \FA_INST_0[1].FA_INST_1[508].FA_  ( .A(A[1020]), .B(n6), .CI(
        C[1020]), .CO(C[1021]) );
  FA_14657 \FA_INST_0[1].FA_INST_1[509].FA_  ( .A(A[1021]), .B(n5), .CI(
        C[1021]), .CO(C[1022]) );
  FA_14656 \FA_INST_0[1].FA_INST_1[510].FA_  ( .A(A[1022]), .B(n4), .CI(
        C[1022]), .CO(C[1023]) );
  FA_14655 \FA_INST_0[1].FA_INST_1[511].FA_  ( .A(A[1023]), .B(n3), .CI(
        C[1023]), .CO(C[1024]) );
  FA_14654 \FA_INST_1[1024].FA_  ( .A(A[1024]), .B(1'b1), .CI(C[1024]), .CO(
        C[1025]) );
  FA_14653 \FA_INST_1[1025].FA_  ( .A(A[1025]), .B(1'b1), .CI(C[1025]), .CO(O)
         );
  IV U2 ( .A(B[27]), .Z(n999) );
  IV U3 ( .A(B[28]), .Z(n998) );
  IV U4 ( .A(B[29]), .Z(n997) );
  IV U5 ( .A(B[30]), .Z(n996) );
  IV U6 ( .A(B[31]), .Z(n995) );
  IV U7 ( .A(B[32]), .Z(n994) );
  IV U8 ( .A(B[33]), .Z(n993) );
  IV U9 ( .A(B[34]), .Z(n992) );
  IV U10 ( .A(B[35]), .Z(n991) );
  IV U11 ( .A(B[36]), .Z(n990) );
  IV U12 ( .A(B[927]), .Z(n99) );
  IV U13 ( .A(B[37]), .Z(n989) );
  IV U14 ( .A(B[38]), .Z(n988) );
  IV U15 ( .A(B[39]), .Z(n987) );
  IV U16 ( .A(B[40]), .Z(n986) );
  IV U17 ( .A(B[41]), .Z(n985) );
  IV U18 ( .A(B[42]), .Z(n984) );
  IV U19 ( .A(B[43]), .Z(n983) );
  IV U20 ( .A(B[44]), .Z(n982) );
  IV U21 ( .A(B[45]), .Z(n981) );
  IV U22 ( .A(B[46]), .Z(n980) );
  IV U23 ( .A(B[928]), .Z(n98) );
  IV U24 ( .A(B[47]), .Z(n979) );
  IV U25 ( .A(B[48]), .Z(n978) );
  IV U26 ( .A(B[49]), .Z(n977) );
  IV U27 ( .A(B[50]), .Z(n976) );
  IV U28 ( .A(B[51]), .Z(n975) );
  IV U29 ( .A(B[52]), .Z(n974) );
  IV U30 ( .A(B[53]), .Z(n973) );
  IV U31 ( .A(B[54]), .Z(n972) );
  IV U32 ( .A(B[55]), .Z(n971) );
  IV U33 ( .A(B[56]), .Z(n970) );
  IV U34 ( .A(B[929]), .Z(n97) );
  IV U35 ( .A(B[57]), .Z(n969) );
  IV U36 ( .A(B[58]), .Z(n968) );
  IV U37 ( .A(B[59]), .Z(n967) );
  IV U38 ( .A(B[60]), .Z(n966) );
  IV U39 ( .A(B[61]), .Z(n965) );
  IV U40 ( .A(B[62]), .Z(n964) );
  IV U41 ( .A(B[63]), .Z(n963) );
  IV U42 ( .A(B[64]), .Z(n962) );
  IV U43 ( .A(B[65]), .Z(n961) );
  IV U44 ( .A(B[66]), .Z(n960) );
  IV U45 ( .A(B[930]), .Z(n96) );
  IV U46 ( .A(B[67]), .Z(n959) );
  IV U47 ( .A(B[68]), .Z(n958) );
  IV U48 ( .A(B[69]), .Z(n957) );
  IV U49 ( .A(B[70]), .Z(n956) );
  IV U50 ( .A(B[71]), .Z(n955) );
  IV U51 ( .A(B[72]), .Z(n954) );
  IV U52 ( .A(B[73]), .Z(n953) );
  IV U53 ( .A(B[74]), .Z(n952) );
  IV U54 ( .A(B[75]), .Z(n951) );
  IV U55 ( .A(B[76]), .Z(n950) );
  IV U56 ( .A(B[931]), .Z(n95) );
  IV U57 ( .A(B[77]), .Z(n949) );
  IV U58 ( .A(B[78]), .Z(n948) );
  IV U59 ( .A(B[79]), .Z(n947) );
  IV U60 ( .A(B[80]), .Z(n946) );
  IV U61 ( .A(B[81]), .Z(n945) );
  IV U62 ( .A(B[82]), .Z(n944) );
  IV U63 ( .A(B[83]), .Z(n943) );
  IV U64 ( .A(B[84]), .Z(n942) );
  IV U65 ( .A(B[85]), .Z(n941) );
  IV U66 ( .A(B[86]), .Z(n940) );
  IV U67 ( .A(B[932]), .Z(n94) );
  IV U68 ( .A(B[87]), .Z(n939) );
  IV U69 ( .A(B[88]), .Z(n938) );
  IV U70 ( .A(B[89]), .Z(n937) );
  IV U71 ( .A(B[90]), .Z(n936) );
  IV U72 ( .A(B[91]), .Z(n935) );
  IV U73 ( .A(B[92]), .Z(n934) );
  IV U74 ( .A(B[93]), .Z(n933) );
  IV U75 ( .A(B[94]), .Z(n932) );
  IV U76 ( .A(B[95]), .Z(n931) );
  IV U77 ( .A(B[96]), .Z(n930) );
  IV U78 ( .A(B[933]), .Z(n93) );
  IV U79 ( .A(B[97]), .Z(n929) );
  IV U80 ( .A(B[98]), .Z(n928) );
  IV U81 ( .A(B[99]), .Z(n927) );
  IV U82 ( .A(B[100]), .Z(n926) );
  IV U83 ( .A(B[101]), .Z(n925) );
  IV U84 ( .A(B[102]), .Z(n924) );
  IV U85 ( .A(B[103]), .Z(n923) );
  IV U86 ( .A(B[104]), .Z(n922) );
  IV U87 ( .A(B[105]), .Z(n921) );
  IV U88 ( .A(B[106]), .Z(n920) );
  IV U89 ( .A(B[934]), .Z(n92) );
  IV U90 ( .A(B[107]), .Z(n919) );
  IV U91 ( .A(B[108]), .Z(n918) );
  IV U92 ( .A(B[109]), .Z(n917) );
  IV U93 ( .A(B[110]), .Z(n916) );
  IV U94 ( .A(B[111]), .Z(n915) );
  IV U95 ( .A(B[112]), .Z(n914) );
  IV U96 ( .A(B[113]), .Z(n913) );
  IV U97 ( .A(B[114]), .Z(n912) );
  IV U98 ( .A(B[115]), .Z(n911) );
  IV U99 ( .A(B[116]), .Z(n910) );
  IV U100 ( .A(B[935]), .Z(n91) );
  IV U101 ( .A(B[117]), .Z(n909) );
  IV U102 ( .A(B[118]), .Z(n908) );
  IV U103 ( .A(B[119]), .Z(n907) );
  IV U104 ( .A(B[120]), .Z(n906) );
  IV U105 ( .A(B[121]), .Z(n905) );
  IV U106 ( .A(B[122]), .Z(n904) );
  IV U107 ( .A(B[123]), .Z(n903) );
  IV U108 ( .A(B[124]), .Z(n902) );
  IV U109 ( .A(B[125]), .Z(n901) );
  IV U110 ( .A(B[126]), .Z(n900) );
  IV U111 ( .A(B[936]), .Z(n90) );
  IV U112 ( .A(B[1017]), .Z(n9) );
  IV U113 ( .A(B[127]), .Z(n899) );
  IV U114 ( .A(B[128]), .Z(n898) );
  IV U115 ( .A(B[129]), .Z(n897) );
  IV U116 ( .A(B[130]), .Z(n896) );
  IV U117 ( .A(B[131]), .Z(n895) );
  IV U118 ( .A(B[132]), .Z(n894) );
  IV U119 ( .A(B[133]), .Z(n893) );
  IV U120 ( .A(B[134]), .Z(n892) );
  IV U121 ( .A(B[135]), .Z(n891) );
  IV U122 ( .A(B[136]), .Z(n890) );
  IV U123 ( .A(B[937]), .Z(n89) );
  IV U124 ( .A(B[137]), .Z(n889) );
  IV U125 ( .A(B[138]), .Z(n888) );
  IV U126 ( .A(B[139]), .Z(n887) );
  IV U127 ( .A(B[140]), .Z(n886) );
  IV U128 ( .A(B[141]), .Z(n885) );
  IV U129 ( .A(B[142]), .Z(n884) );
  IV U130 ( .A(B[143]), .Z(n883) );
  IV U131 ( .A(B[144]), .Z(n882) );
  IV U132 ( .A(B[145]), .Z(n881) );
  IV U133 ( .A(B[146]), .Z(n880) );
  IV U134 ( .A(B[938]), .Z(n88) );
  IV U135 ( .A(B[147]), .Z(n879) );
  IV U136 ( .A(B[148]), .Z(n878) );
  IV U137 ( .A(B[149]), .Z(n877) );
  IV U138 ( .A(B[150]), .Z(n876) );
  IV U139 ( .A(B[151]), .Z(n875) );
  IV U140 ( .A(B[152]), .Z(n874) );
  IV U141 ( .A(B[153]), .Z(n873) );
  IV U142 ( .A(B[154]), .Z(n872) );
  IV U143 ( .A(B[155]), .Z(n871) );
  IV U144 ( .A(B[156]), .Z(n870) );
  IV U145 ( .A(B[939]), .Z(n87) );
  IV U146 ( .A(B[157]), .Z(n869) );
  IV U147 ( .A(B[158]), .Z(n868) );
  IV U148 ( .A(B[159]), .Z(n867) );
  IV U149 ( .A(B[160]), .Z(n866) );
  IV U150 ( .A(B[161]), .Z(n865) );
  IV U151 ( .A(B[162]), .Z(n864) );
  IV U152 ( .A(B[163]), .Z(n863) );
  IV U153 ( .A(B[164]), .Z(n862) );
  IV U154 ( .A(B[165]), .Z(n861) );
  IV U155 ( .A(B[166]), .Z(n860) );
  IV U156 ( .A(B[940]), .Z(n86) );
  IV U157 ( .A(B[167]), .Z(n859) );
  IV U158 ( .A(B[168]), .Z(n858) );
  IV U159 ( .A(B[169]), .Z(n857) );
  IV U160 ( .A(B[170]), .Z(n856) );
  IV U161 ( .A(B[171]), .Z(n855) );
  IV U162 ( .A(B[172]), .Z(n854) );
  IV U163 ( .A(B[173]), .Z(n853) );
  IV U164 ( .A(B[174]), .Z(n852) );
  IV U165 ( .A(B[175]), .Z(n851) );
  IV U166 ( .A(B[176]), .Z(n850) );
  IV U167 ( .A(B[941]), .Z(n85) );
  IV U168 ( .A(B[177]), .Z(n849) );
  IV U169 ( .A(B[178]), .Z(n848) );
  IV U170 ( .A(B[179]), .Z(n847) );
  IV U171 ( .A(B[180]), .Z(n846) );
  IV U172 ( .A(B[181]), .Z(n845) );
  IV U173 ( .A(B[182]), .Z(n844) );
  IV U174 ( .A(B[183]), .Z(n843) );
  IV U175 ( .A(B[184]), .Z(n842) );
  IV U176 ( .A(B[185]), .Z(n841) );
  IV U177 ( .A(B[186]), .Z(n840) );
  IV U178 ( .A(B[942]), .Z(n84) );
  IV U179 ( .A(B[187]), .Z(n839) );
  IV U180 ( .A(B[188]), .Z(n838) );
  IV U181 ( .A(B[189]), .Z(n837) );
  IV U182 ( .A(B[190]), .Z(n836) );
  IV U183 ( .A(B[191]), .Z(n835) );
  IV U184 ( .A(B[192]), .Z(n834) );
  IV U185 ( .A(B[193]), .Z(n833) );
  IV U186 ( .A(B[194]), .Z(n832) );
  IV U187 ( .A(B[195]), .Z(n831) );
  IV U188 ( .A(B[196]), .Z(n830) );
  IV U189 ( .A(B[943]), .Z(n83) );
  IV U190 ( .A(B[197]), .Z(n829) );
  IV U191 ( .A(B[198]), .Z(n828) );
  IV U192 ( .A(B[199]), .Z(n827) );
  IV U193 ( .A(B[200]), .Z(n826) );
  IV U194 ( .A(B[201]), .Z(n825) );
  IV U195 ( .A(B[202]), .Z(n824) );
  IV U196 ( .A(B[203]), .Z(n823) );
  IV U197 ( .A(B[204]), .Z(n822) );
  IV U198 ( .A(B[205]), .Z(n821) );
  IV U199 ( .A(B[206]), .Z(n820) );
  IV U200 ( .A(B[944]), .Z(n82) );
  IV U201 ( .A(B[207]), .Z(n819) );
  IV U202 ( .A(B[208]), .Z(n818) );
  IV U203 ( .A(B[209]), .Z(n817) );
  IV U204 ( .A(B[210]), .Z(n816) );
  IV U205 ( .A(B[211]), .Z(n815) );
  IV U206 ( .A(B[212]), .Z(n814) );
  IV U207 ( .A(B[213]), .Z(n813) );
  IV U208 ( .A(B[214]), .Z(n812) );
  IV U209 ( .A(B[215]), .Z(n811) );
  IV U210 ( .A(B[216]), .Z(n810) );
  IV U211 ( .A(B[945]), .Z(n81) );
  IV U212 ( .A(B[217]), .Z(n809) );
  IV U213 ( .A(B[218]), .Z(n808) );
  IV U214 ( .A(B[219]), .Z(n807) );
  IV U215 ( .A(B[220]), .Z(n806) );
  IV U216 ( .A(B[221]), .Z(n805) );
  IV U217 ( .A(B[222]), .Z(n804) );
  IV U218 ( .A(B[223]), .Z(n803) );
  IV U219 ( .A(B[224]), .Z(n802) );
  IV U220 ( .A(B[225]), .Z(n801) );
  IV U221 ( .A(B[226]), .Z(n800) );
  IV U222 ( .A(B[946]), .Z(n80) );
  IV U223 ( .A(B[1018]), .Z(n8) );
  IV U224 ( .A(B[227]), .Z(n799) );
  IV U225 ( .A(B[228]), .Z(n798) );
  IV U226 ( .A(B[229]), .Z(n797) );
  IV U227 ( .A(B[230]), .Z(n796) );
  IV U228 ( .A(B[231]), .Z(n795) );
  IV U229 ( .A(B[232]), .Z(n794) );
  IV U230 ( .A(B[233]), .Z(n793) );
  IV U231 ( .A(B[234]), .Z(n792) );
  IV U232 ( .A(B[235]), .Z(n791) );
  IV U233 ( .A(B[236]), .Z(n790) );
  IV U234 ( .A(B[947]), .Z(n79) );
  IV U235 ( .A(B[237]), .Z(n789) );
  IV U236 ( .A(B[238]), .Z(n788) );
  IV U237 ( .A(B[239]), .Z(n787) );
  IV U238 ( .A(B[240]), .Z(n786) );
  IV U239 ( .A(B[241]), .Z(n785) );
  IV U240 ( .A(B[242]), .Z(n784) );
  IV U241 ( .A(B[243]), .Z(n783) );
  IV U242 ( .A(B[244]), .Z(n782) );
  IV U243 ( .A(B[245]), .Z(n781) );
  IV U244 ( .A(B[246]), .Z(n780) );
  IV U245 ( .A(B[948]), .Z(n78) );
  IV U246 ( .A(B[247]), .Z(n779) );
  IV U247 ( .A(B[248]), .Z(n778) );
  IV U248 ( .A(B[249]), .Z(n777) );
  IV U249 ( .A(B[250]), .Z(n776) );
  IV U250 ( .A(B[251]), .Z(n775) );
  IV U251 ( .A(B[252]), .Z(n774) );
  IV U252 ( .A(B[253]), .Z(n773) );
  IV U253 ( .A(B[254]), .Z(n772) );
  IV U254 ( .A(B[255]), .Z(n771) );
  IV U255 ( .A(B[256]), .Z(n770) );
  IV U256 ( .A(B[949]), .Z(n77) );
  IV U257 ( .A(B[257]), .Z(n769) );
  IV U258 ( .A(B[258]), .Z(n768) );
  IV U259 ( .A(B[259]), .Z(n767) );
  IV U260 ( .A(B[260]), .Z(n766) );
  IV U261 ( .A(B[261]), .Z(n765) );
  IV U262 ( .A(B[262]), .Z(n764) );
  IV U263 ( .A(B[263]), .Z(n763) );
  IV U264 ( .A(B[264]), .Z(n762) );
  IV U265 ( .A(B[265]), .Z(n761) );
  IV U266 ( .A(B[266]), .Z(n760) );
  IV U267 ( .A(B[950]), .Z(n76) );
  IV U268 ( .A(B[267]), .Z(n759) );
  IV U269 ( .A(B[268]), .Z(n758) );
  IV U270 ( .A(B[269]), .Z(n757) );
  IV U271 ( .A(B[270]), .Z(n756) );
  IV U272 ( .A(B[271]), .Z(n755) );
  IV U273 ( .A(B[272]), .Z(n754) );
  IV U274 ( .A(B[273]), .Z(n753) );
  IV U275 ( .A(B[274]), .Z(n752) );
  IV U276 ( .A(B[275]), .Z(n751) );
  IV U277 ( .A(B[276]), .Z(n750) );
  IV U278 ( .A(B[951]), .Z(n75) );
  IV U279 ( .A(B[277]), .Z(n749) );
  IV U280 ( .A(B[278]), .Z(n748) );
  IV U281 ( .A(B[279]), .Z(n747) );
  IV U282 ( .A(B[280]), .Z(n746) );
  IV U283 ( .A(B[281]), .Z(n745) );
  IV U284 ( .A(B[282]), .Z(n744) );
  IV U285 ( .A(B[283]), .Z(n743) );
  IV U286 ( .A(B[284]), .Z(n742) );
  IV U287 ( .A(B[285]), .Z(n741) );
  IV U288 ( .A(B[286]), .Z(n740) );
  IV U289 ( .A(B[952]), .Z(n74) );
  IV U290 ( .A(B[287]), .Z(n739) );
  IV U291 ( .A(B[288]), .Z(n738) );
  IV U292 ( .A(B[289]), .Z(n737) );
  IV U293 ( .A(B[290]), .Z(n736) );
  IV U294 ( .A(B[291]), .Z(n735) );
  IV U295 ( .A(B[292]), .Z(n734) );
  IV U296 ( .A(B[293]), .Z(n733) );
  IV U297 ( .A(B[294]), .Z(n732) );
  IV U298 ( .A(B[295]), .Z(n731) );
  IV U299 ( .A(B[296]), .Z(n730) );
  IV U300 ( .A(B[953]), .Z(n73) );
  IV U301 ( .A(B[297]), .Z(n729) );
  IV U302 ( .A(B[298]), .Z(n728) );
  IV U303 ( .A(B[299]), .Z(n727) );
  IV U304 ( .A(B[300]), .Z(n726) );
  IV U305 ( .A(B[301]), .Z(n725) );
  IV U306 ( .A(B[302]), .Z(n724) );
  IV U307 ( .A(B[303]), .Z(n723) );
  IV U308 ( .A(B[304]), .Z(n722) );
  IV U309 ( .A(B[305]), .Z(n721) );
  IV U310 ( .A(B[306]), .Z(n720) );
  IV U311 ( .A(B[954]), .Z(n72) );
  IV U312 ( .A(B[307]), .Z(n719) );
  IV U313 ( .A(B[308]), .Z(n718) );
  IV U314 ( .A(B[309]), .Z(n717) );
  IV U315 ( .A(B[310]), .Z(n716) );
  IV U316 ( .A(B[311]), .Z(n715) );
  IV U317 ( .A(B[312]), .Z(n714) );
  IV U318 ( .A(B[313]), .Z(n713) );
  IV U319 ( .A(B[314]), .Z(n712) );
  IV U320 ( .A(B[315]), .Z(n711) );
  IV U321 ( .A(B[316]), .Z(n710) );
  IV U322 ( .A(B[955]), .Z(n71) );
  IV U323 ( .A(B[317]), .Z(n709) );
  IV U324 ( .A(B[318]), .Z(n708) );
  IV U325 ( .A(B[319]), .Z(n707) );
  IV U326 ( .A(B[320]), .Z(n706) );
  IV U327 ( .A(B[321]), .Z(n705) );
  IV U328 ( .A(B[322]), .Z(n704) );
  IV U329 ( .A(B[323]), .Z(n703) );
  IV U330 ( .A(B[324]), .Z(n702) );
  IV U331 ( .A(B[325]), .Z(n701) );
  IV U332 ( .A(B[326]), .Z(n700) );
  IV U333 ( .A(B[956]), .Z(n70) );
  IV U334 ( .A(B[1019]), .Z(n7) );
  IV U335 ( .A(B[327]), .Z(n699) );
  IV U336 ( .A(B[328]), .Z(n698) );
  IV U337 ( .A(B[329]), .Z(n697) );
  IV U338 ( .A(B[330]), .Z(n696) );
  IV U339 ( .A(B[331]), .Z(n695) );
  IV U340 ( .A(B[332]), .Z(n694) );
  IV U341 ( .A(B[333]), .Z(n693) );
  IV U342 ( .A(B[334]), .Z(n692) );
  IV U343 ( .A(B[335]), .Z(n691) );
  IV U344 ( .A(B[336]), .Z(n690) );
  IV U345 ( .A(B[957]), .Z(n69) );
  IV U346 ( .A(B[337]), .Z(n689) );
  IV U347 ( .A(B[338]), .Z(n688) );
  IV U348 ( .A(B[339]), .Z(n687) );
  IV U349 ( .A(B[340]), .Z(n686) );
  IV U350 ( .A(B[341]), .Z(n685) );
  IV U351 ( .A(B[342]), .Z(n684) );
  IV U352 ( .A(B[343]), .Z(n683) );
  IV U353 ( .A(B[344]), .Z(n682) );
  IV U354 ( .A(B[345]), .Z(n681) );
  IV U355 ( .A(B[346]), .Z(n680) );
  IV U356 ( .A(B[958]), .Z(n68) );
  IV U357 ( .A(B[347]), .Z(n679) );
  IV U358 ( .A(B[348]), .Z(n678) );
  IV U359 ( .A(B[349]), .Z(n677) );
  IV U360 ( .A(B[350]), .Z(n676) );
  IV U361 ( .A(B[351]), .Z(n675) );
  IV U362 ( .A(B[352]), .Z(n674) );
  IV U363 ( .A(B[353]), .Z(n673) );
  IV U364 ( .A(B[354]), .Z(n672) );
  IV U365 ( .A(B[355]), .Z(n671) );
  IV U366 ( .A(B[356]), .Z(n670) );
  IV U367 ( .A(B[959]), .Z(n67) );
  IV U368 ( .A(B[357]), .Z(n669) );
  IV U369 ( .A(B[358]), .Z(n668) );
  IV U370 ( .A(B[359]), .Z(n667) );
  IV U371 ( .A(B[360]), .Z(n666) );
  IV U372 ( .A(B[361]), .Z(n665) );
  IV U373 ( .A(B[362]), .Z(n664) );
  IV U374 ( .A(B[363]), .Z(n663) );
  IV U375 ( .A(B[364]), .Z(n662) );
  IV U376 ( .A(B[365]), .Z(n661) );
  IV U377 ( .A(B[366]), .Z(n660) );
  IV U378 ( .A(B[960]), .Z(n66) );
  IV U379 ( .A(B[367]), .Z(n659) );
  IV U380 ( .A(B[368]), .Z(n658) );
  IV U381 ( .A(B[369]), .Z(n657) );
  IV U382 ( .A(B[370]), .Z(n656) );
  IV U383 ( .A(B[371]), .Z(n655) );
  IV U384 ( .A(B[372]), .Z(n654) );
  IV U385 ( .A(B[373]), .Z(n653) );
  IV U386 ( .A(B[374]), .Z(n652) );
  IV U387 ( .A(B[375]), .Z(n651) );
  IV U388 ( .A(B[376]), .Z(n650) );
  IV U389 ( .A(B[961]), .Z(n65) );
  IV U390 ( .A(B[377]), .Z(n649) );
  IV U391 ( .A(B[378]), .Z(n648) );
  IV U392 ( .A(B[379]), .Z(n647) );
  IV U393 ( .A(B[380]), .Z(n646) );
  IV U394 ( .A(B[381]), .Z(n645) );
  IV U395 ( .A(B[382]), .Z(n644) );
  IV U396 ( .A(B[383]), .Z(n643) );
  IV U397 ( .A(B[384]), .Z(n642) );
  IV U398 ( .A(B[385]), .Z(n641) );
  IV U399 ( .A(B[386]), .Z(n640) );
  IV U400 ( .A(B[962]), .Z(n64) );
  IV U401 ( .A(B[387]), .Z(n639) );
  IV U402 ( .A(B[388]), .Z(n638) );
  IV U403 ( .A(B[389]), .Z(n637) );
  IV U404 ( .A(B[390]), .Z(n636) );
  IV U405 ( .A(B[391]), .Z(n635) );
  IV U406 ( .A(B[392]), .Z(n634) );
  IV U407 ( .A(B[393]), .Z(n633) );
  IV U408 ( .A(B[394]), .Z(n632) );
  IV U409 ( .A(B[395]), .Z(n631) );
  IV U410 ( .A(B[396]), .Z(n630) );
  IV U411 ( .A(B[963]), .Z(n63) );
  IV U412 ( .A(B[397]), .Z(n629) );
  IV U413 ( .A(B[398]), .Z(n628) );
  IV U414 ( .A(B[399]), .Z(n627) );
  IV U415 ( .A(B[400]), .Z(n626) );
  IV U416 ( .A(B[401]), .Z(n625) );
  IV U417 ( .A(B[402]), .Z(n624) );
  IV U418 ( .A(B[403]), .Z(n623) );
  IV U419 ( .A(B[404]), .Z(n622) );
  IV U420 ( .A(B[405]), .Z(n621) );
  IV U421 ( .A(B[406]), .Z(n620) );
  IV U422 ( .A(B[964]), .Z(n62) );
  IV U423 ( .A(B[407]), .Z(n619) );
  IV U424 ( .A(B[408]), .Z(n618) );
  IV U425 ( .A(B[409]), .Z(n617) );
  IV U426 ( .A(B[410]), .Z(n616) );
  IV U427 ( .A(B[411]), .Z(n615) );
  IV U428 ( .A(B[412]), .Z(n614) );
  IV U429 ( .A(B[413]), .Z(n613) );
  IV U430 ( .A(B[414]), .Z(n612) );
  IV U431 ( .A(B[415]), .Z(n611) );
  IV U432 ( .A(B[416]), .Z(n610) );
  IV U433 ( .A(B[965]), .Z(n61) );
  IV U434 ( .A(B[417]), .Z(n609) );
  IV U435 ( .A(B[418]), .Z(n608) );
  IV U436 ( .A(B[419]), .Z(n607) );
  IV U437 ( .A(B[420]), .Z(n606) );
  IV U438 ( .A(B[421]), .Z(n605) );
  IV U439 ( .A(B[422]), .Z(n604) );
  IV U440 ( .A(B[423]), .Z(n603) );
  IV U441 ( .A(B[424]), .Z(n602) );
  IV U442 ( .A(B[425]), .Z(n601) );
  IV U443 ( .A(B[426]), .Z(n600) );
  IV U444 ( .A(B[966]), .Z(n60) );
  IV U445 ( .A(B[1020]), .Z(n6) );
  IV U446 ( .A(B[427]), .Z(n599) );
  IV U447 ( .A(B[428]), .Z(n598) );
  IV U448 ( .A(B[429]), .Z(n597) );
  IV U449 ( .A(B[430]), .Z(n596) );
  IV U450 ( .A(B[431]), .Z(n595) );
  IV U451 ( .A(B[432]), .Z(n594) );
  IV U452 ( .A(B[433]), .Z(n593) );
  IV U453 ( .A(B[434]), .Z(n592) );
  IV U454 ( .A(B[435]), .Z(n591) );
  IV U455 ( .A(B[436]), .Z(n590) );
  IV U456 ( .A(B[967]), .Z(n59) );
  IV U457 ( .A(B[437]), .Z(n589) );
  IV U458 ( .A(B[438]), .Z(n588) );
  IV U459 ( .A(B[439]), .Z(n587) );
  IV U460 ( .A(B[440]), .Z(n586) );
  IV U461 ( .A(B[441]), .Z(n585) );
  IV U462 ( .A(B[442]), .Z(n584) );
  IV U463 ( .A(B[443]), .Z(n583) );
  IV U464 ( .A(B[444]), .Z(n582) );
  IV U465 ( .A(B[445]), .Z(n581) );
  IV U466 ( .A(B[446]), .Z(n580) );
  IV U467 ( .A(B[968]), .Z(n58) );
  IV U468 ( .A(B[447]), .Z(n579) );
  IV U469 ( .A(B[448]), .Z(n578) );
  IV U470 ( .A(B[449]), .Z(n577) );
  IV U471 ( .A(B[450]), .Z(n576) );
  IV U472 ( .A(B[451]), .Z(n575) );
  IV U473 ( .A(B[452]), .Z(n574) );
  IV U474 ( .A(B[453]), .Z(n573) );
  IV U475 ( .A(B[454]), .Z(n572) );
  IV U476 ( .A(B[455]), .Z(n571) );
  IV U477 ( .A(B[456]), .Z(n570) );
  IV U478 ( .A(B[969]), .Z(n57) );
  IV U479 ( .A(B[457]), .Z(n569) );
  IV U480 ( .A(B[458]), .Z(n568) );
  IV U481 ( .A(B[459]), .Z(n567) );
  IV U482 ( .A(B[460]), .Z(n566) );
  IV U483 ( .A(B[461]), .Z(n565) );
  IV U484 ( .A(B[462]), .Z(n564) );
  IV U485 ( .A(B[463]), .Z(n563) );
  IV U486 ( .A(B[464]), .Z(n562) );
  IV U487 ( .A(B[465]), .Z(n561) );
  IV U488 ( .A(B[466]), .Z(n560) );
  IV U489 ( .A(B[970]), .Z(n56) );
  IV U490 ( .A(B[467]), .Z(n559) );
  IV U491 ( .A(B[468]), .Z(n558) );
  IV U492 ( .A(B[469]), .Z(n557) );
  IV U493 ( .A(B[470]), .Z(n556) );
  IV U494 ( .A(B[471]), .Z(n555) );
  IV U495 ( .A(B[472]), .Z(n554) );
  IV U496 ( .A(B[473]), .Z(n553) );
  IV U497 ( .A(B[474]), .Z(n552) );
  IV U498 ( .A(B[475]), .Z(n551) );
  IV U499 ( .A(B[476]), .Z(n550) );
  IV U500 ( .A(B[971]), .Z(n55) );
  IV U501 ( .A(B[477]), .Z(n549) );
  IV U502 ( .A(B[478]), .Z(n548) );
  IV U503 ( .A(B[479]), .Z(n547) );
  IV U504 ( .A(B[480]), .Z(n546) );
  IV U505 ( .A(B[481]), .Z(n545) );
  IV U506 ( .A(B[482]), .Z(n544) );
  IV U507 ( .A(B[483]), .Z(n543) );
  IV U508 ( .A(B[484]), .Z(n542) );
  IV U509 ( .A(B[485]), .Z(n541) );
  IV U510 ( .A(B[486]), .Z(n540) );
  IV U511 ( .A(B[972]), .Z(n54) );
  IV U512 ( .A(B[487]), .Z(n539) );
  IV U513 ( .A(B[488]), .Z(n538) );
  IV U514 ( .A(B[489]), .Z(n537) );
  IV U515 ( .A(B[490]), .Z(n536) );
  IV U516 ( .A(B[491]), .Z(n535) );
  IV U517 ( .A(B[492]), .Z(n534) );
  IV U518 ( .A(B[493]), .Z(n533) );
  IV U519 ( .A(B[494]), .Z(n532) );
  IV U520 ( .A(B[495]), .Z(n531) );
  IV U521 ( .A(B[496]), .Z(n530) );
  IV U522 ( .A(B[973]), .Z(n53) );
  IV U523 ( .A(B[497]), .Z(n529) );
  IV U524 ( .A(B[498]), .Z(n528) );
  IV U525 ( .A(B[499]), .Z(n527) );
  IV U526 ( .A(B[500]), .Z(n526) );
  IV U527 ( .A(B[501]), .Z(n525) );
  IV U528 ( .A(B[502]), .Z(n524) );
  IV U529 ( .A(B[503]), .Z(n523) );
  IV U530 ( .A(B[504]), .Z(n522) );
  IV U531 ( .A(B[505]), .Z(n521) );
  IV U532 ( .A(B[506]), .Z(n520) );
  IV U533 ( .A(B[974]), .Z(n52) );
  IV U534 ( .A(B[507]), .Z(n519) );
  IV U535 ( .A(B[508]), .Z(n518) );
  IV U536 ( .A(B[509]), .Z(n517) );
  IV U537 ( .A(B[510]), .Z(n516) );
  IV U538 ( .A(B[511]), .Z(n515) );
  IV U539 ( .A(B[512]), .Z(n514) );
  IV U540 ( .A(B[513]), .Z(n513) );
  IV U541 ( .A(B[514]), .Z(n512) );
  IV U542 ( .A(B[515]), .Z(n511) );
  IV U543 ( .A(B[516]), .Z(n510) );
  IV U544 ( .A(B[975]), .Z(n51) );
  IV U545 ( .A(B[517]), .Z(n509) );
  IV U546 ( .A(B[518]), .Z(n508) );
  IV U547 ( .A(B[519]), .Z(n507) );
  IV U548 ( .A(B[520]), .Z(n506) );
  IV U549 ( .A(B[521]), .Z(n505) );
  IV U550 ( .A(B[522]), .Z(n504) );
  IV U551 ( .A(B[523]), .Z(n503) );
  IV U552 ( .A(B[524]), .Z(n502) );
  IV U553 ( .A(B[525]), .Z(n501) );
  IV U554 ( .A(B[526]), .Z(n500) );
  IV U555 ( .A(B[976]), .Z(n50) );
  IV U556 ( .A(B[1021]), .Z(n5) );
  IV U557 ( .A(B[527]), .Z(n499) );
  IV U558 ( .A(B[528]), .Z(n498) );
  IV U559 ( .A(B[529]), .Z(n497) );
  IV U560 ( .A(B[530]), .Z(n496) );
  IV U561 ( .A(B[531]), .Z(n495) );
  IV U562 ( .A(B[532]), .Z(n494) );
  IV U563 ( .A(B[533]), .Z(n493) );
  IV U564 ( .A(B[534]), .Z(n492) );
  IV U565 ( .A(B[535]), .Z(n491) );
  IV U566 ( .A(B[536]), .Z(n490) );
  IV U567 ( .A(B[977]), .Z(n49) );
  IV U568 ( .A(B[537]), .Z(n489) );
  IV U569 ( .A(B[538]), .Z(n488) );
  IV U570 ( .A(B[539]), .Z(n487) );
  IV U571 ( .A(B[540]), .Z(n486) );
  IV U572 ( .A(B[541]), .Z(n485) );
  IV U573 ( .A(B[542]), .Z(n484) );
  IV U574 ( .A(B[543]), .Z(n483) );
  IV U575 ( .A(B[544]), .Z(n482) );
  IV U576 ( .A(B[545]), .Z(n481) );
  IV U577 ( .A(B[546]), .Z(n480) );
  IV U578 ( .A(B[978]), .Z(n48) );
  IV U579 ( .A(B[547]), .Z(n479) );
  IV U580 ( .A(B[548]), .Z(n478) );
  IV U581 ( .A(B[549]), .Z(n477) );
  IV U582 ( .A(B[550]), .Z(n476) );
  IV U583 ( .A(B[551]), .Z(n475) );
  IV U584 ( .A(B[552]), .Z(n474) );
  IV U585 ( .A(B[553]), .Z(n473) );
  IV U586 ( .A(B[554]), .Z(n472) );
  IV U587 ( .A(B[555]), .Z(n471) );
  IV U588 ( .A(B[556]), .Z(n470) );
  IV U589 ( .A(B[979]), .Z(n47) );
  IV U590 ( .A(B[557]), .Z(n469) );
  IV U591 ( .A(B[558]), .Z(n468) );
  IV U592 ( .A(B[559]), .Z(n467) );
  IV U593 ( .A(B[560]), .Z(n466) );
  IV U594 ( .A(B[561]), .Z(n465) );
  IV U595 ( .A(B[562]), .Z(n464) );
  IV U596 ( .A(B[563]), .Z(n463) );
  IV U597 ( .A(B[564]), .Z(n462) );
  IV U598 ( .A(B[565]), .Z(n461) );
  IV U599 ( .A(B[566]), .Z(n460) );
  IV U600 ( .A(B[980]), .Z(n46) );
  IV U601 ( .A(B[567]), .Z(n459) );
  IV U602 ( .A(B[568]), .Z(n458) );
  IV U603 ( .A(B[569]), .Z(n457) );
  IV U604 ( .A(B[570]), .Z(n456) );
  IV U605 ( .A(B[571]), .Z(n455) );
  IV U606 ( .A(B[572]), .Z(n454) );
  IV U607 ( .A(B[573]), .Z(n453) );
  IV U608 ( .A(B[574]), .Z(n452) );
  IV U609 ( .A(B[575]), .Z(n451) );
  IV U610 ( .A(B[576]), .Z(n450) );
  IV U611 ( .A(B[981]), .Z(n45) );
  IV U612 ( .A(B[577]), .Z(n449) );
  IV U613 ( .A(B[578]), .Z(n448) );
  IV U614 ( .A(B[579]), .Z(n447) );
  IV U615 ( .A(B[580]), .Z(n446) );
  IV U616 ( .A(B[581]), .Z(n445) );
  IV U617 ( .A(B[582]), .Z(n444) );
  IV U618 ( .A(B[583]), .Z(n443) );
  IV U619 ( .A(B[584]), .Z(n442) );
  IV U620 ( .A(B[585]), .Z(n441) );
  IV U621 ( .A(B[586]), .Z(n440) );
  IV U622 ( .A(B[982]), .Z(n44) );
  IV U623 ( .A(B[587]), .Z(n439) );
  IV U624 ( .A(B[588]), .Z(n438) );
  IV U625 ( .A(B[589]), .Z(n437) );
  IV U626 ( .A(B[590]), .Z(n436) );
  IV U627 ( .A(B[591]), .Z(n435) );
  IV U628 ( .A(B[592]), .Z(n434) );
  IV U629 ( .A(B[593]), .Z(n433) );
  IV U630 ( .A(B[594]), .Z(n432) );
  IV U631 ( .A(B[595]), .Z(n431) );
  IV U632 ( .A(B[596]), .Z(n430) );
  IV U633 ( .A(B[983]), .Z(n43) );
  IV U634 ( .A(B[597]), .Z(n429) );
  IV U635 ( .A(B[598]), .Z(n428) );
  IV U636 ( .A(B[599]), .Z(n427) );
  IV U637 ( .A(B[600]), .Z(n426) );
  IV U638 ( .A(B[601]), .Z(n425) );
  IV U639 ( .A(B[602]), .Z(n424) );
  IV U640 ( .A(B[603]), .Z(n423) );
  IV U641 ( .A(B[604]), .Z(n422) );
  IV U642 ( .A(B[605]), .Z(n421) );
  IV U643 ( .A(B[606]), .Z(n420) );
  IV U644 ( .A(B[984]), .Z(n42) );
  IV U645 ( .A(B[607]), .Z(n419) );
  IV U646 ( .A(B[608]), .Z(n418) );
  IV U647 ( .A(B[609]), .Z(n417) );
  IV U648 ( .A(B[610]), .Z(n416) );
  IV U649 ( .A(B[611]), .Z(n415) );
  IV U650 ( .A(B[612]), .Z(n414) );
  IV U651 ( .A(B[613]), .Z(n413) );
  IV U652 ( .A(B[614]), .Z(n412) );
  IV U653 ( .A(B[615]), .Z(n411) );
  IV U654 ( .A(B[616]), .Z(n410) );
  IV U655 ( .A(B[985]), .Z(n41) );
  IV U656 ( .A(B[617]), .Z(n409) );
  IV U657 ( .A(B[618]), .Z(n408) );
  IV U658 ( .A(B[619]), .Z(n407) );
  IV U659 ( .A(B[620]), .Z(n406) );
  IV U660 ( .A(B[621]), .Z(n405) );
  IV U661 ( .A(B[622]), .Z(n404) );
  IV U662 ( .A(B[623]), .Z(n403) );
  IV U663 ( .A(B[624]), .Z(n402) );
  IV U664 ( .A(B[625]), .Z(n401) );
  IV U665 ( .A(B[626]), .Z(n400) );
  IV U666 ( .A(B[986]), .Z(n40) );
  IV U667 ( .A(B[1022]), .Z(n4) );
  IV U668 ( .A(B[627]), .Z(n399) );
  IV U669 ( .A(B[628]), .Z(n398) );
  IV U670 ( .A(B[629]), .Z(n397) );
  IV U671 ( .A(B[630]), .Z(n396) );
  IV U672 ( .A(B[631]), .Z(n395) );
  IV U673 ( .A(B[632]), .Z(n394) );
  IV U674 ( .A(B[633]), .Z(n393) );
  IV U675 ( .A(B[634]), .Z(n392) );
  IV U676 ( .A(B[635]), .Z(n391) );
  IV U677 ( .A(B[636]), .Z(n390) );
  IV U678 ( .A(B[987]), .Z(n39) );
  IV U679 ( .A(B[637]), .Z(n389) );
  IV U680 ( .A(B[638]), .Z(n388) );
  IV U681 ( .A(B[639]), .Z(n387) );
  IV U682 ( .A(B[640]), .Z(n386) );
  IV U683 ( .A(B[641]), .Z(n385) );
  IV U684 ( .A(B[642]), .Z(n384) );
  IV U685 ( .A(B[643]), .Z(n383) );
  IV U686 ( .A(B[644]), .Z(n382) );
  IV U687 ( .A(B[645]), .Z(n381) );
  IV U688 ( .A(B[646]), .Z(n380) );
  IV U689 ( .A(B[988]), .Z(n38) );
  IV U690 ( .A(B[647]), .Z(n379) );
  IV U691 ( .A(B[648]), .Z(n378) );
  IV U692 ( .A(B[649]), .Z(n377) );
  IV U693 ( .A(B[650]), .Z(n376) );
  IV U694 ( .A(B[651]), .Z(n375) );
  IV U695 ( .A(B[652]), .Z(n374) );
  IV U696 ( .A(B[653]), .Z(n373) );
  IV U697 ( .A(B[654]), .Z(n372) );
  IV U698 ( .A(B[655]), .Z(n371) );
  IV U699 ( .A(B[656]), .Z(n370) );
  IV U700 ( .A(B[989]), .Z(n37) );
  IV U701 ( .A(B[657]), .Z(n369) );
  IV U702 ( .A(B[658]), .Z(n368) );
  IV U703 ( .A(B[659]), .Z(n367) );
  IV U704 ( .A(B[660]), .Z(n366) );
  IV U705 ( .A(B[661]), .Z(n365) );
  IV U706 ( .A(B[662]), .Z(n364) );
  IV U707 ( .A(B[663]), .Z(n363) );
  IV U708 ( .A(B[664]), .Z(n362) );
  IV U709 ( .A(B[665]), .Z(n361) );
  IV U710 ( .A(B[666]), .Z(n360) );
  IV U711 ( .A(B[990]), .Z(n36) );
  IV U712 ( .A(B[667]), .Z(n359) );
  IV U713 ( .A(B[668]), .Z(n358) );
  IV U714 ( .A(B[669]), .Z(n357) );
  IV U715 ( .A(B[670]), .Z(n356) );
  IV U716 ( .A(B[671]), .Z(n355) );
  IV U717 ( .A(B[672]), .Z(n354) );
  IV U718 ( .A(B[673]), .Z(n353) );
  IV U719 ( .A(B[674]), .Z(n352) );
  IV U720 ( .A(B[675]), .Z(n351) );
  IV U721 ( .A(B[676]), .Z(n350) );
  IV U722 ( .A(B[991]), .Z(n35) );
  IV U723 ( .A(B[677]), .Z(n349) );
  IV U724 ( .A(B[678]), .Z(n348) );
  IV U725 ( .A(B[679]), .Z(n347) );
  IV U726 ( .A(B[680]), .Z(n346) );
  IV U727 ( .A(B[681]), .Z(n345) );
  IV U728 ( .A(B[682]), .Z(n344) );
  IV U729 ( .A(B[683]), .Z(n343) );
  IV U730 ( .A(B[684]), .Z(n342) );
  IV U731 ( .A(B[685]), .Z(n341) );
  IV U732 ( .A(B[686]), .Z(n340) );
  IV U733 ( .A(B[992]), .Z(n34) );
  IV U734 ( .A(B[687]), .Z(n339) );
  IV U735 ( .A(B[688]), .Z(n338) );
  IV U736 ( .A(B[689]), .Z(n337) );
  IV U737 ( .A(B[690]), .Z(n336) );
  IV U738 ( .A(B[691]), .Z(n335) );
  IV U739 ( .A(B[692]), .Z(n334) );
  IV U740 ( .A(B[693]), .Z(n333) );
  IV U741 ( .A(B[694]), .Z(n332) );
  IV U742 ( .A(B[695]), .Z(n331) );
  IV U743 ( .A(B[696]), .Z(n330) );
  IV U744 ( .A(B[993]), .Z(n33) );
  IV U745 ( .A(B[697]), .Z(n329) );
  IV U746 ( .A(B[698]), .Z(n328) );
  IV U747 ( .A(B[699]), .Z(n327) );
  IV U748 ( .A(B[700]), .Z(n326) );
  IV U749 ( .A(B[701]), .Z(n325) );
  IV U750 ( .A(B[702]), .Z(n324) );
  IV U751 ( .A(B[703]), .Z(n323) );
  IV U752 ( .A(B[704]), .Z(n322) );
  IV U753 ( .A(B[705]), .Z(n321) );
  IV U754 ( .A(B[706]), .Z(n320) );
  IV U755 ( .A(B[994]), .Z(n32) );
  IV U756 ( .A(B[707]), .Z(n319) );
  IV U757 ( .A(B[708]), .Z(n318) );
  IV U758 ( .A(B[709]), .Z(n317) );
  IV U759 ( .A(B[710]), .Z(n316) );
  IV U760 ( .A(B[711]), .Z(n315) );
  IV U761 ( .A(B[712]), .Z(n314) );
  IV U762 ( .A(B[713]), .Z(n313) );
  IV U763 ( .A(B[714]), .Z(n312) );
  IV U764 ( .A(B[715]), .Z(n311) );
  IV U765 ( .A(B[716]), .Z(n310) );
  IV U766 ( .A(B[995]), .Z(n31) );
  IV U767 ( .A(B[717]), .Z(n309) );
  IV U768 ( .A(B[718]), .Z(n308) );
  IV U769 ( .A(B[719]), .Z(n307) );
  IV U770 ( .A(B[720]), .Z(n306) );
  IV U771 ( .A(B[721]), .Z(n305) );
  IV U772 ( .A(B[722]), .Z(n304) );
  IV U773 ( .A(B[723]), .Z(n303) );
  IV U774 ( .A(B[724]), .Z(n302) );
  IV U775 ( .A(B[725]), .Z(n301) );
  IV U776 ( .A(B[726]), .Z(n300) );
  IV U777 ( .A(B[996]), .Z(n30) );
  IV U778 ( .A(B[1023]), .Z(n3) );
  IV U779 ( .A(B[727]), .Z(n299) );
  IV U780 ( .A(B[728]), .Z(n298) );
  IV U781 ( .A(B[729]), .Z(n297) );
  IV U782 ( .A(B[730]), .Z(n296) );
  IV U783 ( .A(B[731]), .Z(n295) );
  IV U784 ( .A(B[732]), .Z(n294) );
  IV U785 ( .A(B[733]), .Z(n293) );
  IV U786 ( .A(B[734]), .Z(n292) );
  IV U787 ( .A(B[735]), .Z(n291) );
  IV U788 ( .A(B[736]), .Z(n290) );
  IV U789 ( .A(B[997]), .Z(n29) );
  IV U790 ( .A(B[737]), .Z(n289) );
  IV U791 ( .A(B[738]), .Z(n288) );
  IV U792 ( .A(B[739]), .Z(n287) );
  IV U793 ( .A(B[740]), .Z(n286) );
  IV U794 ( .A(B[741]), .Z(n285) );
  IV U795 ( .A(B[742]), .Z(n284) );
  IV U796 ( .A(B[743]), .Z(n283) );
  IV U797 ( .A(B[744]), .Z(n282) );
  IV U798 ( .A(B[745]), .Z(n281) );
  IV U799 ( .A(B[746]), .Z(n280) );
  IV U800 ( .A(B[998]), .Z(n28) );
  IV U801 ( .A(B[747]), .Z(n279) );
  IV U802 ( .A(B[748]), .Z(n278) );
  IV U803 ( .A(B[749]), .Z(n277) );
  IV U804 ( .A(B[750]), .Z(n276) );
  IV U805 ( .A(B[751]), .Z(n275) );
  IV U806 ( .A(B[752]), .Z(n274) );
  IV U807 ( .A(B[753]), .Z(n273) );
  IV U808 ( .A(B[754]), .Z(n272) );
  IV U809 ( .A(B[755]), .Z(n271) );
  IV U810 ( .A(B[756]), .Z(n270) );
  IV U811 ( .A(B[999]), .Z(n27) );
  IV U812 ( .A(B[757]), .Z(n269) );
  IV U813 ( .A(B[758]), .Z(n268) );
  IV U814 ( .A(B[759]), .Z(n267) );
  IV U815 ( .A(B[760]), .Z(n266) );
  IV U816 ( .A(B[761]), .Z(n265) );
  IV U817 ( .A(B[762]), .Z(n264) );
  IV U818 ( .A(B[763]), .Z(n263) );
  IV U819 ( .A(B[764]), .Z(n262) );
  IV U820 ( .A(B[765]), .Z(n261) );
  IV U821 ( .A(B[766]), .Z(n260) );
  IV U822 ( .A(B[1000]), .Z(n26) );
  IV U823 ( .A(B[767]), .Z(n259) );
  IV U824 ( .A(B[768]), .Z(n258) );
  IV U825 ( .A(B[769]), .Z(n257) );
  IV U826 ( .A(B[770]), .Z(n256) );
  IV U827 ( .A(B[771]), .Z(n255) );
  IV U828 ( .A(B[772]), .Z(n254) );
  IV U829 ( .A(B[773]), .Z(n253) );
  IV U830 ( .A(B[774]), .Z(n252) );
  IV U831 ( .A(B[775]), .Z(n251) );
  IV U832 ( .A(B[776]), .Z(n250) );
  IV U833 ( .A(B[1001]), .Z(n25) );
  IV U834 ( .A(B[777]), .Z(n249) );
  IV U835 ( .A(B[778]), .Z(n248) );
  IV U836 ( .A(B[779]), .Z(n247) );
  IV U837 ( .A(B[780]), .Z(n246) );
  IV U838 ( .A(B[781]), .Z(n245) );
  IV U839 ( .A(B[782]), .Z(n244) );
  IV U840 ( .A(B[783]), .Z(n243) );
  IV U841 ( .A(B[784]), .Z(n242) );
  IV U842 ( .A(B[785]), .Z(n241) );
  IV U843 ( .A(B[786]), .Z(n240) );
  IV U844 ( .A(B[1002]), .Z(n24) );
  IV U845 ( .A(B[787]), .Z(n239) );
  IV U846 ( .A(B[788]), .Z(n238) );
  IV U847 ( .A(B[789]), .Z(n237) );
  IV U848 ( .A(B[790]), .Z(n236) );
  IV U849 ( .A(B[791]), .Z(n235) );
  IV U850 ( .A(B[792]), .Z(n234) );
  IV U851 ( .A(B[793]), .Z(n233) );
  IV U852 ( .A(B[794]), .Z(n232) );
  IV U853 ( .A(B[795]), .Z(n231) );
  IV U854 ( .A(B[796]), .Z(n230) );
  IV U855 ( .A(B[1003]), .Z(n23) );
  IV U856 ( .A(B[797]), .Z(n229) );
  IV U857 ( .A(B[798]), .Z(n228) );
  IV U858 ( .A(B[799]), .Z(n227) );
  IV U859 ( .A(B[800]), .Z(n226) );
  IV U860 ( .A(B[801]), .Z(n225) );
  IV U861 ( .A(B[802]), .Z(n224) );
  IV U862 ( .A(B[803]), .Z(n223) );
  IV U863 ( .A(B[804]), .Z(n222) );
  IV U864 ( .A(B[805]), .Z(n221) );
  IV U865 ( .A(B[806]), .Z(n220) );
  IV U866 ( .A(B[1004]), .Z(n22) );
  IV U867 ( .A(B[807]), .Z(n219) );
  IV U868 ( .A(B[808]), .Z(n218) );
  IV U869 ( .A(B[809]), .Z(n217) );
  IV U870 ( .A(B[810]), .Z(n216) );
  IV U871 ( .A(B[811]), .Z(n215) );
  IV U872 ( .A(B[812]), .Z(n214) );
  IV U873 ( .A(B[813]), .Z(n213) );
  IV U874 ( .A(B[814]), .Z(n212) );
  IV U875 ( .A(B[815]), .Z(n211) );
  IV U876 ( .A(B[816]), .Z(n210) );
  IV U877 ( .A(B[1005]), .Z(n21) );
  IV U878 ( .A(B[817]), .Z(n209) );
  IV U879 ( .A(B[818]), .Z(n208) );
  IV U880 ( .A(B[819]), .Z(n207) );
  IV U881 ( .A(B[820]), .Z(n206) );
  IV U882 ( .A(B[821]), .Z(n205) );
  IV U883 ( .A(B[822]), .Z(n204) );
  IV U884 ( .A(B[823]), .Z(n203) );
  IV U885 ( .A(B[824]), .Z(n202) );
  IV U886 ( .A(B[825]), .Z(n201) );
  IV U887 ( .A(B[826]), .Z(n200) );
  IV U888 ( .A(B[1006]), .Z(n20) );
  IV U889 ( .A(B[827]), .Z(n199) );
  IV U890 ( .A(B[828]), .Z(n198) );
  IV U891 ( .A(B[829]), .Z(n197) );
  IV U892 ( .A(B[830]), .Z(n196) );
  IV U893 ( .A(B[831]), .Z(n195) );
  IV U894 ( .A(B[832]), .Z(n194) );
  IV U895 ( .A(B[833]), .Z(n193) );
  IV U896 ( .A(B[834]), .Z(n192) );
  IV U897 ( .A(B[835]), .Z(n191) );
  IV U898 ( .A(B[836]), .Z(n190) );
  IV U899 ( .A(B[1007]), .Z(n19) );
  IV U900 ( .A(B[837]), .Z(n189) );
  IV U901 ( .A(B[838]), .Z(n188) );
  IV U902 ( .A(B[839]), .Z(n187) );
  IV U903 ( .A(B[840]), .Z(n186) );
  IV U904 ( .A(B[841]), .Z(n185) );
  IV U905 ( .A(B[842]), .Z(n184) );
  IV U906 ( .A(B[843]), .Z(n183) );
  IV U907 ( .A(B[844]), .Z(n182) );
  IV U908 ( .A(B[845]), .Z(n181) );
  IV U909 ( .A(B[846]), .Z(n180) );
  IV U910 ( .A(B[1008]), .Z(n18) );
  IV U911 ( .A(B[847]), .Z(n179) );
  IV U912 ( .A(B[848]), .Z(n178) );
  IV U913 ( .A(B[849]), .Z(n177) );
  IV U914 ( .A(B[850]), .Z(n176) );
  IV U915 ( .A(B[851]), .Z(n175) );
  IV U916 ( .A(B[852]), .Z(n174) );
  IV U917 ( .A(B[853]), .Z(n173) );
  IV U918 ( .A(B[854]), .Z(n172) );
  IV U919 ( .A(B[855]), .Z(n171) );
  IV U920 ( .A(B[856]), .Z(n170) );
  IV U921 ( .A(B[1009]), .Z(n17) );
  IV U922 ( .A(B[857]), .Z(n169) );
  IV U923 ( .A(B[858]), .Z(n168) );
  IV U924 ( .A(B[859]), .Z(n167) );
  IV U925 ( .A(B[860]), .Z(n166) );
  IV U926 ( .A(B[861]), .Z(n165) );
  IV U927 ( .A(B[862]), .Z(n164) );
  IV U928 ( .A(B[863]), .Z(n163) );
  IV U929 ( .A(B[864]), .Z(n162) );
  IV U930 ( .A(B[865]), .Z(n161) );
  IV U931 ( .A(B[866]), .Z(n160) );
  IV U932 ( .A(B[1010]), .Z(n16) );
  IV U933 ( .A(B[867]), .Z(n159) );
  IV U934 ( .A(B[868]), .Z(n158) );
  IV U935 ( .A(B[869]), .Z(n157) );
  IV U936 ( .A(B[870]), .Z(n156) );
  IV U937 ( .A(B[871]), .Z(n155) );
  IV U938 ( .A(B[872]), .Z(n154) );
  IV U939 ( .A(B[873]), .Z(n153) );
  IV U940 ( .A(B[874]), .Z(n152) );
  IV U941 ( .A(B[875]), .Z(n151) );
  IV U942 ( .A(B[876]), .Z(n150) );
  IV U943 ( .A(B[1011]), .Z(n15) );
  IV U944 ( .A(B[877]), .Z(n149) );
  IV U945 ( .A(B[878]), .Z(n148) );
  IV U946 ( .A(B[879]), .Z(n147) );
  IV U947 ( .A(B[880]), .Z(n146) );
  IV U948 ( .A(B[881]), .Z(n145) );
  IV U949 ( .A(B[882]), .Z(n144) );
  IV U950 ( .A(B[883]), .Z(n143) );
  IV U951 ( .A(B[884]), .Z(n142) );
  IV U952 ( .A(B[885]), .Z(n141) );
  IV U953 ( .A(B[886]), .Z(n140) );
  IV U954 ( .A(B[1012]), .Z(n14) );
  IV U955 ( .A(B[887]), .Z(n139) );
  IV U956 ( .A(B[888]), .Z(n138) );
  IV U957 ( .A(B[889]), .Z(n137) );
  IV U958 ( .A(B[890]), .Z(n136) );
  IV U959 ( .A(B[891]), .Z(n135) );
  IV U960 ( .A(B[892]), .Z(n134) );
  IV U961 ( .A(B[893]), .Z(n133) );
  IV U962 ( .A(B[894]), .Z(n132) );
  IV U963 ( .A(B[895]), .Z(n131) );
  IV U964 ( .A(B[896]), .Z(n130) );
  IV U965 ( .A(B[1013]), .Z(n13) );
  IV U966 ( .A(B[897]), .Z(n129) );
  IV U967 ( .A(B[898]), .Z(n128) );
  IV U968 ( .A(B[899]), .Z(n127) );
  IV U969 ( .A(B[900]), .Z(n126) );
  IV U970 ( .A(B[901]), .Z(n125) );
  IV U971 ( .A(B[902]), .Z(n124) );
  IV U972 ( .A(B[903]), .Z(n123) );
  IV U973 ( .A(B[904]), .Z(n122) );
  IV U974 ( .A(B[905]), .Z(n121) );
  IV U975 ( .A(B[906]), .Z(n120) );
  IV U976 ( .A(B[1014]), .Z(n12) );
  IV U977 ( .A(B[907]), .Z(n119) );
  IV U978 ( .A(B[908]), .Z(n118) );
  IV U979 ( .A(B[909]), .Z(n117) );
  IV U980 ( .A(B[910]), .Z(n116) );
  IV U981 ( .A(B[911]), .Z(n115) );
  IV U982 ( .A(B[912]), .Z(n114) );
  IV U983 ( .A(B[913]), .Z(n113) );
  IV U984 ( .A(B[914]), .Z(n112) );
  IV U985 ( .A(B[915]), .Z(n111) );
  IV U986 ( .A(B[916]), .Z(n110) );
  IV U987 ( .A(B[1015]), .Z(n11) );
  IV U988 ( .A(B[917]), .Z(n109) );
  IV U989 ( .A(B[918]), .Z(n108) );
  IV U990 ( .A(B[919]), .Z(n107) );
  IV U991 ( .A(B[920]), .Z(n106) );
  IV U992 ( .A(B[921]), .Z(n105) );
  IV U993 ( .A(B[922]), .Z(n104) );
  IV U994 ( .A(B[923]), .Z(n103) );
  IV U995 ( .A(B[0]), .Z(n1026) );
  IV U996 ( .A(B[1]), .Z(n1025) );
  IV U997 ( .A(B[2]), .Z(n1024) );
  IV U998 ( .A(B[3]), .Z(n1023) );
  IV U999 ( .A(B[4]), .Z(n1022) );
  IV U1000 ( .A(B[5]), .Z(n1021) );
  IV U1001 ( .A(B[6]), .Z(n1020) );
  IV U1002 ( .A(B[924]), .Z(n102) );
  IV U1003 ( .A(B[7]), .Z(n1019) );
  IV U1004 ( .A(B[8]), .Z(n1018) );
  IV U1005 ( .A(B[9]), .Z(n1017) );
  IV U1006 ( .A(B[10]), .Z(n1016) );
  IV U1007 ( .A(B[11]), .Z(n1015) );
  IV U1008 ( .A(B[12]), .Z(n1014) );
  IV U1009 ( .A(B[13]), .Z(n1013) );
  IV U1010 ( .A(B[14]), .Z(n1012) );
  IV U1011 ( .A(B[15]), .Z(n1011) );
  IV U1012 ( .A(B[16]), .Z(n1010) );
  IV U1013 ( .A(B[925]), .Z(n101) );
  IV U1014 ( .A(B[17]), .Z(n1009) );
  IV U1015 ( .A(B[18]), .Z(n1008) );
  IV U1016 ( .A(B[19]), .Z(n1007) );
  IV U1017 ( .A(B[20]), .Z(n1006) );
  IV U1018 ( .A(B[21]), .Z(n1005) );
  IV U1019 ( .A(B[22]), .Z(n1004) );
  IV U1020 ( .A(B[23]), .Z(n1003) );
  IV U1021 ( .A(B[24]), .Z(n1002) );
  IV U1022 ( .A(B[25]), .Z(n1001) );
  IV U1023 ( .A(B[26]), .Z(n1000) );
  IV U1024 ( .A(B[926]), .Z(n100) );
  IV U1025 ( .A(B[1016]), .Z(n10) );
endmodule


module FA_13627 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XNOR U1 ( .A(CI), .B(A), .Z(S) );
endmodule


module FA_13628 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  NANDN U1 ( .A(CI), .B(S), .Z(CO) );
  XNOR U2 ( .A(A), .B(CI), .Z(S) );
endmodule


module FA_13629 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13630 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13631 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13632 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13633 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13634 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13635 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13636 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13637 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13638 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13639 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13640 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13641 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13642 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13643 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13644 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13645 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13646 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13647 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13648 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13649 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13650 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13651 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13652 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13653 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13654 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13655 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13656 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13657 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13658 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13659 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13660 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13661 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13662 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13663 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13664 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13665 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13666 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13667 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13668 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13669 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13670 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13671 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13672 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13673 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13674 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13675 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13676 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13677 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13678 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13679 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13680 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13681 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13682 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13683 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13684 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13685 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13686 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13687 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13688 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13689 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13690 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13691 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13692 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13693 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13694 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13695 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13696 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13697 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13698 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13699 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13700 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13701 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13702 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13703 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13704 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13705 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13706 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13707 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13708 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13709 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13710 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13711 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13712 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13713 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13714 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13715 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13716 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13717 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13718 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13719 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13720 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13721 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13722 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13723 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13724 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13725 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13726 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13727 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13728 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13729 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13730 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13731 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13732 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13733 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13734 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13735 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13736 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13737 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13738 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13739 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13740 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13741 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13742 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13743 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13744 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13745 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13746 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13747 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13748 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13749 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13750 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13751 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13752 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13753 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13754 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13755 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13756 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13757 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13758 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13759 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13760 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13761 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13762 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13763 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13764 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13765 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13766 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13767 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13768 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13769 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13770 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13771 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13772 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13773 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13774 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13775 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13776 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13777 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13778 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13779 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13780 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13781 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13782 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13783 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13784 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13785 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13786 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13787 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13788 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13789 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13790 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13791 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13792 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13793 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13794 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13795 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13796 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13797 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13798 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13799 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13800 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13801 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13802 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13803 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13804 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13805 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13806 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13807 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13808 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13809 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13810 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13811 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13812 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13813 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13814 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13815 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13816 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13817 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13818 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13819 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13820 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13821 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13822 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13823 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13824 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13825 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13826 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13827 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13828 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13829 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13830 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13831 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13832 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13833 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13834 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13835 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13836 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13837 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13838 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13839 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13840 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13841 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13842 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13843 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13844 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13845 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13846 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13847 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13848 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13849 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13850 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13851 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13852 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13853 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13854 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13855 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13856 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13857 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13858 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13859 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13860 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13861 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13862 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13863 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13864 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13865 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13866 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13867 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13868 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13869 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13870 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13871 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13872 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13873 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13874 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13875 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13876 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13877 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13878 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13879 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13880 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13881 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13882 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13883 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13884 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13885 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13886 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13887 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13888 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13889 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13890 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13891 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13892 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13893 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13894 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13895 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13896 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13897 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13898 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13899 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13900 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13901 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13902 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13903 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13904 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13905 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13906 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13907 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13908 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13909 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13910 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13911 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13912 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13913 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13914 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13915 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13916 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13917 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13918 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13919 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13920 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13921 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13922 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13923 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13924 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13925 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13926 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13927 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13928 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13929 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13930 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13931 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13932 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13933 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13934 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13935 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13936 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13937 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13938 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13939 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13940 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13941 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13942 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13943 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13944 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13945 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13946 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13947 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13948 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13949 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13950 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13951 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13952 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13953 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13954 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13955 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13956 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13957 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13958 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13959 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13960 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13961 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13962 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13963 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13964 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13965 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13966 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13967 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13968 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13969 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13970 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13971 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13972 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13973 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13974 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13975 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13976 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13977 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13978 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13979 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13980 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13981 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13982 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13983 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13984 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13985 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13986 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13987 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13988 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13989 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13990 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13991 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13992 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13993 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13994 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13995 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13996 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13997 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13998 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13999 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14000 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14001 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14002 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14003 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14004 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14005 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14006 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14007 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14008 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14009 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14010 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14011 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14012 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14013 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14014 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14015 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14016 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14017 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14018 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14019 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14020 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14021 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14022 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14023 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14024 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14025 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14026 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14027 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14028 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14029 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14030 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14031 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14032 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14033 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14034 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14035 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14036 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14037 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14038 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14039 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14040 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14041 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14042 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14043 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14044 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14045 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14046 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14047 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14048 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14049 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14050 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14051 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14052 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14053 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14054 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14055 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14056 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14057 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14058 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14059 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14060 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14061 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14062 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14063 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14064 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14065 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14066 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14067 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14068 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14069 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14070 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14071 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14072 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14073 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14074 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14075 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14076 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14077 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14078 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14079 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14080 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14081 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14082 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14083 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14084 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14085 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14086 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14087 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14088 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14089 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14090 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14091 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14092 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14093 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14094 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14095 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14096 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14097 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14098 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14099 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14100 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14101 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14102 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14103 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14104 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14105 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14106 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14107 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14108 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14109 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14110 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14111 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14112 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14113 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14114 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14115 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14116 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14117 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14118 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14119 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14120 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14121 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14122 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14123 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14124 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14125 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14126 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14127 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14128 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14129 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14130 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14131 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14132 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14133 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14134 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14135 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14136 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14137 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14138 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14139 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14140 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14141 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14142 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14143 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14144 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14145 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14146 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14147 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14148 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14149 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14150 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14151 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14152 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14153 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14154 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14155 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14156 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14157 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14158 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14159 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14160 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14161 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14162 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14163 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14164 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14165 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14166 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14167 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14168 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14169 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14170 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14171 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14172 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14173 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14174 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14175 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14176 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14177 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14178 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14179 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14180 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14181 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14182 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14183 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14184 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14185 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14186 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14187 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14188 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14189 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14190 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14191 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14192 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14193 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14194 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14195 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14196 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14197 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14198 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14199 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14200 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14201 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14202 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14203 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14204 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14205 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14206 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14207 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14208 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14209 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14210 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14211 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14212 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14213 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14214 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14215 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14216 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14217 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14218 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14219 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14220 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14221 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14222 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14223 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14224 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14225 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14226 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14227 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14228 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14229 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14230 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14231 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14232 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14233 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14234 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14235 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14236 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14237 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14238 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14239 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14240 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14241 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14242 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14243 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14244 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14245 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14246 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14247 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14248 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14249 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14250 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14251 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14252 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14253 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14254 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14255 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14256 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14257 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14258 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14259 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14260 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14261 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14262 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14263 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14264 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14265 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14266 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14267 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14268 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14269 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14270 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14271 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14272 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14273 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14274 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14275 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14276 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14277 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14278 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14279 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14280 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14281 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14282 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14283 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14284 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14285 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14286 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14287 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14288 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14289 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14290 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14291 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14292 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14293 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14294 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14295 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14296 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14297 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14298 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14299 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14300 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14301 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14302 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14303 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14304 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14305 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14306 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14307 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14308 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14309 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14310 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14311 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14312 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14313 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14314 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14315 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14316 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14317 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14318 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14319 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14320 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14321 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14322 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14323 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14324 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14325 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14326 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14327 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14328 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14329 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14330 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14331 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14332 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14333 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14334 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14335 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14336 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14337 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14338 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14339 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14340 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14341 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14342 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14343 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14344 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14345 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14346 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14347 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14348 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14349 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14350 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14351 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14352 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14353 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14354 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14355 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14356 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14357 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14358 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14359 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14360 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14361 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14362 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14363 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14364 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14365 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14366 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14367 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14368 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14369 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14370 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14371 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14372 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14373 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14374 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14375 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14376 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14377 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14378 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14379 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14380 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14381 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14382 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14383 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14384 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14385 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14386 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14387 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14388 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14389 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14390 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14391 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14392 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14393 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14394 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14395 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14396 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14397 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14398 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14399 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14400 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14401 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14402 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14403 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14404 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14405 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14406 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14407 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14408 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14409 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14410 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14411 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14412 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14413 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14414 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14415 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14416 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14417 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14418 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14419 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14420 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14421 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14422 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14423 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14424 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14425 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14426 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14427 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14428 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14429 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14430 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14431 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14432 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14433 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14434 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14435 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14436 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14437 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14438 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14439 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14440 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14441 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14442 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14443 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14444 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14445 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14446 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14447 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14448 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14449 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14450 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14451 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14452 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14453 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14454 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14455 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14456 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14457 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14458 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14459 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14460 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14461 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14462 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14463 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14464 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14465 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14466 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14467 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14468 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14469 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14470 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14471 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14472 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14473 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14474 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14475 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14476 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14477 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14478 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14479 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14480 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14481 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14482 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14483 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14484 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14485 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14486 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14487 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14488 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14489 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14490 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14491 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14492 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14493 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14494 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14495 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14496 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14497 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14498 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14499 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14500 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14501 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14502 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14503 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14504 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14505 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14506 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14507 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14508 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14509 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14510 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14511 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14512 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14513 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14514 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14515 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14516 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14517 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14518 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14519 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14520 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14521 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14522 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14523 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14524 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14525 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14526 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14527 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14528 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14529 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14530 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14531 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14532 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14533 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14534 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14535 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14536 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14537 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14538 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14539 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14540 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14541 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14542 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14543 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14544 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14545 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14546 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14547 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14548 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14549 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14550 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14551 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14552 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14553 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14554 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14555 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14556 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14557 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14558 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14559 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14560 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14561 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14562 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14563 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14564 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14565 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14566 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14567 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14568 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14569 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14570 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14571 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14572 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14573 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14574 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14575 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14576 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14577 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14578 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14579 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14580 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14581 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14582 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14583 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14584 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14585 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14586 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14587 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14588 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14589 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14590 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14591 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14592 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14593 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14594 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14595 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14596 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14597 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14598 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14599 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14600 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14601 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14602 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14603 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14604 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14605 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14606 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14607 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14608 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14609 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14610 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14611 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14612 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14613 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14614 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14615 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14616 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14617 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14618 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14619 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14620 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14621 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14622 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14623 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14624 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14625 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14626 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14627 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14628 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14629 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14630 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14631 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14632 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14633 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14634 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14635 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14636 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14637 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14638 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14639 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14640 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14641 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14642 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14643 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14644 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14645 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14646 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14647 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14648 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14649 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14650 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14651 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14652 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XNOR U1 ( .A(B), .B(A), .Z(S) );
  OR U2 ( .A(B), .B(A), .Z(CO) );
endmodule


module SUB_N1026_0 ( A, B, S, CO );
  input [1025:0] A;
  input [1025:0] B;
  output [1025:0] S;
  output CO;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026;
  wire   [1025:1] C;

  FA_14652 \FA_INST_0[0].FA_INST_1[0].FA_  ( .A(A[0]), .B(n1026), .CI(1'b1), 
        .S(S[0]), .CO(C[1]) );
  FA_14651 \FA_INST_0[0].FA_INST_1[1].FA_  ( .A(A[1]), .B(n1025), .CI(C[1]), 
        .S(S[1]), .CO(C[2]) );
  FA_14650 \FA_INST_0[0].FA_INST_1[2].FA_  ( .A(A[2]), .B(n1024), .CI(C[2]), 
        .S(S[2]), .CO(C[3]) );
  FA_14649 \FA_INST_0[0].FA_INST_1[3].FA_  ( .A(A[3]), .B(n1023), .CI(C[3]), 
        .S(S[3]), .CO(C[4]) );
  FA_14648 \FA_INST_0[0].FA_INST_1[4].FA_  ( .A(A[4]), .B(n1022), .CI(C[4]), 
        .S(S[4]), .CO(C[5]) );
  FA_14647 \FA_INST_0[0].FA_INST_1[5].FA_  ( .A(A[5]), .B(n1021), .CI(C[5]), 
        .S(S[5]), .CO(C[6]) );
  FA_14646 \FA_INST_0[0].FA_INST_1[6].FA_  ( .A(A[6]), .B(n1020), .CI(C[6]), 
        .S(S[6]), .CO(C[7]) );
  FA_14645 \FA_INST_0[0].FA_INST_1[7].FA_  ( .A(A[7]), .B(n1019), .CI(C[7]), 
        .S(S[7]), .CO(C[8]) );
  FA_14644 \FA_INST_0[0].FA_INST_1[8].FA_  ( .A(A[8]), .B(n1018), .CI(C[8]), 
        .S(S[8]), .CO(C[9]) );
  FA_14643 \FA_INST_0[0].FA_INST_1[9].FA_  ( .A(A[9]), .B(n1017), .CI(C[9]), 
        .S(S[9]), .CO(C[10]) );
  FA_14642 \FA_INST_0[0].FA_INST_1[10].FA_  ( .A(A[10]), .B(n1016), .CI(C[10]), 
        .S(S[10]), .CO(C[11]) );
  FA_14641 \FA_INST_0[0].FA_INST_1[11].FA_  ( .A(A[11]), .B(n1015), .CI(C[11]), 
        .S(S[11]), .CO(C[12]) );
  FA_14640 \FA_INST_0[0].FA_INST_1[12].FA_  ( .A(A[12]), .B(n1014), .CI(C[12]), 
        .S(S[12]), .CO(C[13]) );
  FA_14639 \FA_INST_0[0].FA_INST_1[13].FA_  ( .A(A[13]), .B(n1013), .CI(C[13]), 
        .S(S[13]), .CO(C[14]) );
  FA_14638 \FA_INST_0[0].FA_INST_1[14].FA_  ( .A(A[14]), .B(n1012), .CI(C[14]), 
        .S(S[14]), .CO(C[15]) );
  FA_14637 \FA_INST_0[0].FA_INST_1[15].FA_  ( .A(A[15]), .B(n1011), .CI(C[15]), 
        .S(S[15]), .CO(C[16]) );
  FA_14636 \FA_INST_0[0].FA_INST_1[16].FA_  ( .A(A[16]), .B(n1010), .CI(C[16]), 
        .S(S[16]), .CO(C[17]) );
  FA_14635 \FA_INST_0[0].FA_INST_1[17].FA_  ( .A(A[17]), .B(n1009), .CI(C[17]), 
        .S(S[17]), .CO(C[18]) );
  FA_14634 \FA_INST_0[0].FA_INST_1[18].FA_  ( .A(A[18]), .B(n1008), .CI(C[18]), 
        .S(S[18]), .CO(C[19]) );
  FA_14633 \FA_INST_0[0].FA_INST_1[19].FA_  ( .A(A[19]), .B(n1007), .CI(C[19]), 
        .S(S[19]), .CO(C[20]) );
  FA_14632 \FA_INST_0[0].FA_INST_1[20].FA_  ( .A(A[20]), .B(n1006), .CI(C[20]), 
        .S(S[20]), .CO(C[21]) );
  FA_14631 \FA_INST_0[0].FA_INST_1[21].FA_  ( .A(A[21]), .B(n1005), .CI(C[21]), 
        .S(S[21]), .CO(C[22]) );
  FA_14630 \FA_INST_0[0].FA_INST_1[22].FA_  ( .A(A[22]), .B(n1004), .CI(C[22]), 
        .S(S[22]), .CO(C[23]) );
  FA_14629 \FA_INST_0[0].FA_INST_1[23].FA_  ( .A(A[23]), .B(n1003), .CI(C[23]), 
        .S(S[23]), .CO(C[24]) );
  FA_14628 \FA_INST_0[0].FA_INST_1[24].FA_  ( .A(A[24]), .B(n1002), .CI(C[24]), 
        .S(S[24]), .CO(C[25]) );
  FA_14627 \FA_INST_0[0].FA_INST_1[25].FA_  ( .A(A[25]), .B(n1001), .CI(C[25]), 
        .S(S[25]), .CO(C[26]) );
  FA_14626 \FA_INST_0[0].FA_INST_1[26].FA_  ( .A(A[26]), .B(n1000), .CI(C[26]), 
        .S(S[26]), .CO(C[27]) );
  FA_14625 \FA_INST_0[0].FA_INST_1[27].FA_  ( .A(A[27]), .B(n999), .CI(C[27]), 
        .S(S[27]), .CO(C[28]) );
  FA_14624 \FA_INST_0[0].FA_INST_1[28].FA_  ( .A(A[28]), .B(n998), .CI(C[28]), 
        .S(S[28]), .CO(C[29]) );
  FA_14623 \FA_INST_0[0].FA_INST_1[29].FA_  ( .A(A[29]), .B(n997), .CI(C[29]), 
        .S(S[29]), .CO(C[30]) );
  FA_14622 \FA_INST_0[0].FA_INST_1[30].FA_  ( .A(A[30]), .B(n996), .CI(C[30]), 
        .S(S[30]), .CO(C[31]) );
  FA_14621 \FA_INST_0[0].FA_INST_1[31].FA_  ( .A(A[31]), .B(n995), .CI(C[31]), 
        .S(S[31]), .CO(C[32]) );
  FA_14620 \FA_INST_0[0].FA_INST_1[32].FA_  ( .A(A[32]), .B(n994), .CI(C[32]), 
        .S(S[32]), .CO(C[33]) );
  FA_14619 \FA_INST_0[0].FA_INST_1[33].FA_  ( .A(A[33]), .B(n993), .CI(C[33]), 
        .S(S[33]), .CO(C[34]) );
  FA_14618 \FA_INST_0[0].FA_INST_1[34].FA_  ( .A(A[34]), .B(n992), .CI(C[34]), 
        .S(S[34]), .CO(C[35]) );
  FA_14617 \FA_INST_0[0].FA_INST_1[35].FA_  ( .A(A[35]), .B(n991), .CI(C[35]), 
        .S(S[35]), .CO(C[36]) );
  FA_14616 \FA_INST_0[0].FA_INST_1[36].FA_  ( .A(A[36]), .B(n990), .CI(C[36]), 
        .S(S[36]), .CO(C[37]) );
  FA_14615 \FA_INST_0[0].FA_INST_1[37].FA_  ( .A(A[37]), .B(n989), .CI(C[37]), 
        .S(S[37]), .CO(C[38]) );
  FA_14614 \FA_INST_0[0].FA_INST_1[38].FA_  ( .A(A[38]), .B(n988), .CI(C[38]), 
        .S(S[38]), .CO(C[39]) );
  FA_14613 \FA_INST_0[0].FA_INST_1[39].FA_  ( .A(A[39]), .B(n987), .CI(C[39]), 
        .S(S[39]), .CO(C[40]) );
  FA_14612 \FA_INST_0[0].FA_INST_1[40].FA_  ( .A(A[40]), .B(n986), .CI(C[40]), 
        .S(S[40]), .CO(C[41]) );
  FA_14611 \FA_INST_0[0].FA_INST_1[41].FA_  ( .A(A[41]), .B(n985), .CI(C[41]), 
        .S(S[41]), .CO(C[42]) );
  FA_14610 \FA_INST_0[0].FA_INST_1[42].FA_  ( .A(A[42]), .B(n984), .CI(C[42]), 
        .S(S[42]), .CO(C[43]) );
  FA_14609 \FA_INST_0[0].FA_INST_1[43].FA_  ( .A(A[43]), .B(n983), .CI(C[43]), 
        .S(S[43]), .CO(C[44]) );
  FA_14608 \FA_INST_0[0].FA_INST_1[44].FA_  ( .A(A[44]), .B(n982), .CI(C[44]), 
        .S(S[44]), .CO(C[45]) );
  FA_14607 \FA_INST_0[0].FA_INST_1[45].FA_  ( .A(A[45]), .B(n981), .CI(C[45]), 
        .S(S[45]), .CO(C[46]) );
  FA_14606 \FA_INST_0[0].FA_INST_1[46].FA_  ( .A(A[46]), .B(n980), .CI(C[46]), 
        .S(S[46]), .CO(C[47]) );
  FA_14605 \FA_INST_0[0].FA_INST_1[47].FA_  ( .A(A[47]), .B(n979), .CI(C[47]), 
        .S(S[47]), .CO(C[48]) );
  FA_14604 \FA_INST_0[0].FA_INST_1[48].FA_  ( .A(A[48]), .B(n978), .CI(C[48]), 
        .S(S[48]), .CO(C[49]) );
  FA_14603 \FA_INST_0[0].FA_INST_1[49].FA_  ( .A(A[49]), .B(n977), .CI(C[49]), 
        .S(S[49]), .CO(C[50]) );
  FA_14602 \FA_INST_0[0].FA_INST_1[50].FA_  ( .A(A[50]), .B(n976), .CI(C[50]), 
        .S(S[50]), .CO(C[51]) );
  FA_14601 \FA_INST_0[0].FA_INST_1[51].FA_  ( .A(A[51]), .B(n975), .CI(C[51]), 
        .S(S[51]), .CO(C[52]) );
  FA_14600 \FA_INST_0[0].FA_INST_1[52].FA_  ( .A(A[52]), .B(n974), .CI(C[52]), 
        .S(S[52]), .CO(C[53]) );
  FA_14599 \FA_INST_0[0].FA_INST_1[53].FA_  ( .A(A[53]), .B(n973), .CI(C[53]), 
        .S(S[53]), .CO(C[54]) );
  FA_14598 \FA_INST_0[0].FA_INST_1[54].FA_  ( .A(A[54]), .B(n972), .CI(C[54]), 
        .S(S[54]), .CO(C[55]) );
  FA_14597 \FA_INST_0[0].FA_INST_1[55].FA_  ( .A(A[55]), .B(n971), .CI(C[55]), 
        .S(S[55]), .CO(C[56]) );
  FA_14596 \FA_INST_0[0].FA_INST_1[56].FA_  ( .A(A[56]), .B(n970), .CI(C[56]), 
        .S(S[56]), .CO(C[57]) );
  FA_14595 \FA_INST_0[0].FA_INST_1[57].FA_  ( .A(A[57]), .B(n969), .CI(C[57]), 
        .S(S[57]), .CO(C[58]) );
  FA_14594 \FA_INST_0[0].FA_INST_1[58].FA_  ( .A(A[58]), .B(n968), .CI(C[58]), 
        .S(S[58]), .CO(C[59]) );
  FA_14593 \FA_INST_0[0].FA_INST_1[59].FA_  ( .A(A[59]), .B(n967), .CI(C[59]), 
        .S(S[59]), .CO(C[60]) );
  FA_14592 \FA_INST_0[0].FA_INST_1[60].FA_  ( .A(A[60]), .B(n966), .CI(C[60]), 
        .S(S[60]), .CO(C[61]) );
  FA_14591 \FA_INST_0[0].FA_INST_1[61].FA_  ( .A(A[61]), .B(n965), .CI(C[61]), 
        .S(S[61]), .CO(C[62]) );
  FA_14590 \FA_INST_0[0].FA_INST_1[62].FA_  ( .A(A[62]), .B(n964), .CI(C[62]), 
        .S(S[62]), .CO(C[63]) );
  FA_14589 \FA_INST_0[0].FA_INST_1[63].FA_  ( .A(A[63]), .B(n963), .CI(C[63]), 
        .S(S[63]), .CO(C[64]) );
  FA_14588 \FA_INST_0[0].FA_INST_1[64].FA_  ( .A(A[64]), .B(n962), .CI(C[64]), 
        .S(S[64]), .CO(C[65]) );
  FA_14587 \FA_INST_0[0].FA_INST_1[65].FA_  ( .A(A[65]), .B(n961), .CI(C[65]), 
        .S(S[65]), .CO(C[66]) );
  FA_14586 \FA_INST_0[0].FA_INST_1[66].FA_  ( .A(A[66]), .B(n960), .CI(C[66]), 
        .S(S[66]), .CO(C[67]) );
  FA_14585 \FA_INST_0[0].FA_INST_1[67].FA_  ( .A(A[67]), .B(n959), .CI(C[67]), 
        .S(S[67]), .CO(C[68]) );
  FA_14584 \FA_INST_0[0].FA_INST_1[68].FA_  ( .A(A[68]), .B(n958), .CI(C[68]), 
        .S(S[68]), .CO(C[69]) );
  FA_14583 \FA_INST_0[0].FA_INST_1[69].FA_  ( .A(A[69]), .B(n957), .CI(C[69]), 
        .S(S[69]), .CO(C[70]) );
  FA_14582 \FA_INST_0[0].FA_INST_1[70].FA_  ( .A(A[70]), .B(n956), .CI(C[70]), 
        .S(S[70]), .CO(C[71]) );
  FA_14581 \FA_INST_0[0].FA_INST_1[71].FA_  ( .A(A[71]), .B(n955), .CI(C[71]), 
        .S(S[71]), .CO(C[72]) );
  FA_14580 \FA_INST_0[0].FA_INST_1[72].FA_  ( .A(A[72]), .B(n954), .CI(C[72]), 
        .S(S[72]), .CO(C[73]) );
  FA_14579 \FA_INST_0[0].FA_INST_1[73].FA_  ( .A(A[73]), .B(n953), .CI(C[73]), 
        .S(S[73]), .CO(C[74]) );
  FA_14578 \FA_INST_0[0].FA_INST_1[74].FA_  ( .A(A[74]), .B(n952), .CI(C[74]), 
        .S(S[74]), .CO(C[75]) );
  FA_14577 \FA_INST_0[0].FA_INST_1[75].FA_  ( .A(A[75]), .B(n951), .CI(C[75]), 
        .S(S[75]), .CO(C[76]) );
  FA_14576 \FA_INST_0[0].FA_INST_1[76].FA_  ( .A(A[76]), .B(n950), .CI(C[76]), 
        .S(S[76]), .CO(C[77]) );
  FA_14575 \FA_INST_0[0].FA_INST_1[77].FA_  ( .A(A[77]), .B(n949), .CI(C[77]), 
        .S(S[77]), .CO(C[78]) );
  FA_14574 \FA_INST_0[0].FA_INST_1[78].FA_  ( .A(A[78]), .B(n948), .CI(C[78]), 
        .S(S[78]), .CO(C[79]) );
  FA_14573 \FA_INST_0[0].FA_INST_1[79].FA_  ( .A(A[79]), .B(n947), .CI(C[79]), 
        .S(S[79]), .CO(C[80]) );
  FA_14572 \FA_INST_0[0].FA_INST_1[80].FA_  ( .A(A[80]), .B(n946), .CI(C[80]), 
        .S(S[80]), .CO(C[81]) );
  FA_14571 \FA_INST_0[0].FA_INST_1[81].FA_  ( .A(A[81]), .B(n945), .CI(C[81]), 
        .S(S[81]), .CO(C[82]) );
  FA_14570 \FA_INST_0[0].FA_INST_1[82].FA_  ( .A(A[82]), .B(n944), .CI(C[82]), 
        .S(S[82]), .CO(C[83]) );
  FA_14569 \FA_INST_0[0].FA_INST_1[83].FA_  ( .A(A[83]), .B(n943), .CI(C[83]), 
        .S(S[83]), .CO(C[84]) );
  FA_14568 \FA_INST_0[0].FA_INST_1[84].FA_  ( .A(A[84]), .B(n942), .CI(C[84]), 
        .S(S[84]), .CO(C[85]) );
  FA_14567 \FA_INST_0[0].FA_INST_1[85].FA_  ( .A(A[85]), .B(n941), .CI(C[85]), 
        .S(S[85]), .CO(C[86]) );
  FA_14566 \FA_INST_0[0].FA_INST_1[86].FA_  ( .A(A[86]), .B(n940), .CI(C[86]), 
        .S(S[86]), .CO(C[87]) );
  FA_14565 \FA_INST_0[0].FA_INST_1[87].FA_  ( .A(A[87]), .B(n939), .CI(C[87]), 
        .S(S[87]), .CO(C[88]) );
  FA_14564 \FA_INST_0[0].FA_INST_1[88].FA_  ( .A(A[88]), .B(n938), .CI(C[88]), 
        .S(S[88]), .CO(C[89]) );
  FA_14563 \FA_INST_0[0].FA_INST_1[89].FA_  ( .A(A[89]), .B(n937), .CI(C[89]), 
        .S(S[89]), .CO(C[90]) );
  FA_14562 \FA_INST_0[0].FA_INST_1[90].FA_  ( .A(A[90]), .B(n936), .CI(C[90]), 
        .S(S[90]), .CO(C[91]) );
  FA_14561 \FA_INST_0[0].FA_INST_1[91].FA_  ( .A(A[91]), .B(n935), .CI(C[91]), 
        .S(S[91]), .CO(C[92]) );
  FA_14560 \FA_INST_0[0].FA_INST_1[92].FA_  ( .A(A[92]), .B(n934), .CI(C[92]), 
        .S(S[92]), .CO(C[93]) );
  FA_14559 \FA_INST_0[0].FA_INST_1[93].FA_  ( .A(A[93]), .B(n933), .CI(C[93]), 
        .S(S[93]), .CO(C[94]) );
  FA_14558 \FA_INST_0[0].FA_INST_1[94].FA_  ( .A(A[94]), .B(n932), .CI(C[94]), 
        .S(S[94]), .CO(C[95]) );
  FA_14557 \FA_INST_0[0].FA_INST_1[95].FA_  ( .A(A[95]), .B(n931), .CI(C[95]), 
        .S(S[95]), .CO(C[96]) );
  FA_14556 \FA_INST_0[0].FA_INST_1[96].FA_  ( .A(A[96]), .B(n930), .CI(C[96]), 
        .S(S[96]), .CO(C[97]) );
  FA_14555 \FA_INST_0[0].FA_INST_1[97].FA_  ( .A(A[97]), .B(n929), .CI(C[97]), 
        .S(S[97]), .CO(C[98]) );
  FA_14554 \FA_INST_0[0].FA_INST_1[98].FA_  ( .A(A[98]), .B(n928), .CI(C[98]), 
        .S(S[98]), .CO(C[99]) );
  FA_14553 \FA_INST_0[0].FA_INST_1[99].FA_  ( .A(A[99]), .B(n927), .CI(C[99]), 
        .S(S[99]), .CO(C[100]) );
  FA_14552 \FA_INST_0[0].FA_INST_1[100].FA_  ( .A(A[100]), .B(n926), .CI(
        C[100]), .S(S[100]), .CO(C[101]) );
  FA_14551 \FA_INST_0[0].FA_INST_1[101].FA_  ( .A(A[101]), .B(n925), .CI(
        C[101]), .S(S[101]), .CO(C[102]) );
  FA_14550 \FA_INST_0[0].FA_INST_1[102].FA_  ( .A(A[102]), .B(n924), .CI(
        C[102]), .S(S[102]), .CO(C[103]) );
  FA_14549 \FA_INST_0[0].FA_INST_1[103].FA_  ( .A(A[103]), .B(n923), .CI(
        C[103]), .S(S[103]), .CO(C[104]) );
  FA_14548 \FA_INST_0[0].FA_INST_1[104].FA_  ( .A(A[104]), .B(n922), .CI(
        C[104]), .S(S[104]), .CO(C[105]) );
  FA_14547 \FA_INST_0[0].FA_INST_1[105].FA_  ( .A(A[105]), .B(n921), .CI(
        C[105]), .S(S[105]), .CO(C[106]) );
  FA_14546 \FA_INST_0[0].FA_INST_1[106].FA_  ( .A(A[106]), .B(n920), .CI(
        C[106]), .S(S[106]), .CO(C[107]) );
  FA_14545 \FA_INST_0[0].FA_INST_1[107].FA_  ( .A(A[107]), .B(n919), .CI(
        C[107]), .S(S[107]), .CO(C[108]) );
  FA_14544 \FA_INST_0[0].FA_INST_1[108].FA_  ( .A(A[108]), .B(n918), .CI(
        C[108]), .S(S[108]), .CO(C[109]) );
  FA_14543 \FA_INST_0[0].FA_INST_1[109].FA_  ( .A(A[109]), .B(n917), .CI(
        C[109]), .S(S[109]), .CO(C[110]) );
  FA_14542 \FA_INST_0[0].FA_INST_1[110].FA_  ( .A(A[110]), .B(n916), .CI(
        C[110]), .S(S[110]), .CO(C[111]) );
  FA_14541 \FA_INST_0[0].FA_INST_1[111].FA_  ( .A(A[111]), .B(n915), .CI(
        C[111]), .S(S[111]), .CO(C[112]) );
  FA_14540 \FA_INST_0[0].FA_INST_1[112].FA_  ( .A(A[112]), .B(n914), .CI(
        C[112]), .S(S[112]), .CO(C[113]) );
  FA_14539 \FA_INST_0[0].FA_INST_1[113].FA_  ( .A(A[113]), .B(n913), .CI(
        C[113]), .S(S[113]), .CO(C[114]) );
  FA_14538 \FA_INST_0[0].FA_INST_1[114].FA_  ( .A(A[114]), .B(n912), .CI(
        C[114]), .S(S[114]), .CO(C[115]) );
  FA_14537 \FA_INST_0[0].FA_INST_1[115].FA_  ( .A(A[115]), .B(n911), .CI(
        C[115]), .S(S[115]), .CO(C[116]) );
  FA_14536 \FA_INST_0[0].FA_INST_1[116].FA_  ( .A(A[116]), .B(n910), .CI(
        C[116]), .S(S[116]), .CO(C[117]) );
  FA_14535 \FA_INST_0[0].FA_INST_1[117].FA_  ( .A(A[117]), .B(n909), .CI(
        C[117]), .S(S[117]), .CO(C[118]) );
  FA_14534 \FA_INST_0[0].FA_INST_1[118].FA_  ( .A(A[118]), .B(n908), .CI(
        C[118]), .S(S[118]), .CO(C[119]) );
  FA_14533 \FA_INST_0[0].FA_INST_1[119].FA_  ( .A(A[119]), .B(n907), .CI(
        C[119]), .S(S[119]), .CO(C[120]) );
  FA_14532 \FA_INST_0[0].FA_INST_1[120].FA_  ( .A(A[120]), .B(n906), .CI(
        C[120]), .S(S[120]), .CO(C[121]) );
  FA_14531 \FA_INST_0[0].FA_INST_1[121].FA_  ( .A(A[121]), .B(n905), .CI(
        C[121]), .S(S[121]), .CO(C[122]) );
  FA_14530 \FA_INST_0[0].FA_INST_1[122].FA_  ( .A(A[122]), .B(n904), .CI(
        C[122]), .S(S[122]), .CO(C[123]) );
  FA_14529 \FA_INST_0[0].FA_INST_1[123].FA_  ( .A(A[123]), .B(n903), .CI(
        C[123]), .S(S[123]), .CO(C[124]) );
  FA_14528 \FA_INST_0[0].FA_INST_1[124].FA_  ( .A(A[124]), .B(n902), .CI(
        C[124]), .S(S[124]), .CO(C[125]) );
  FA_14527 \FA_INST_0[0].FA_INST_1[125].FA_  ( .A(A[125]), .B(n901), .CI(
        C[125]), .S(S[125]), .CO(C[126]) );
  FA_14526 \FA_INST_0[0].FA_INST_1[126].FA_  ( .A(A[126]), .B(n900), .CI(
        C[126]), .S(S[126]), .CO(C[127]) );
  FA_14525 \FA_INST_0[0].FA_INST_1[127].FA_  ( .A(A[127]), .B(n899), .CI(
        C[127]), .S(S[127]), .CO(C[128]) );
  FA_14524 \FA_INST_0[0].FA_INST_1[128].FA_  ( .A(A[128]), .B(n898), .CI(
        C[128]), .S(S[128]), .CO(C[129]) );
  FA_14523 \FA_INST_0[0].FA_INST_1[129].FA_  ( .A(A[129]), .B(n897), .CI(
        C[129]), .S(S[129]), .CO(C[130]) );
  FA_14522 \FA_INST_0[0].FA_INST_1[130].FA_  ( .A(A[130]), .B(n896), .CI(
        C[130]), .S(S[130]), .CO(C[131]) );
  FA_14521 \FA_INST_0[0].FA_INST_1[131].FA_  ( .A(A[131]), .B(n895), .CI(
        C[131]), .S(S[131]), .CO(C[132]) );
  FA_14520 \FA_INST_0[0].FA_INST_1[132].FA_  ( .A(A[132]), .B(n894), .CI(
        C[132]), .S(S[132]), .CO(C[133]) );
  FA_14519 \FA_INST_0[0].FA_INST_1[133].FA_  ( .A(A[133]), .B(n893), .CI(
        C[133]), .S(S[133]), .CO(C[134]) );
  FA_14518 \FA_INST_0[0].FA_INST_1[134].FA_  ( .A(A[134]), .B(n892), .CI(
        C[134]), .S(S[134]), .CO(C[135]) );
  FA_14517 \FA_INST_0[0].FA_INST_1[135].FA_  ( .A(A[135]), .B(n891), .CI(
        C[135]), .S(S[135]), .CO(C[136]) );
  FA_14516 \FA_INST_0[0].FA_INST_1[136].FA_  ( .A(A[136]), .B(n890), .CI(
        C[136]), .S(S[136]), .CO(C[137]) );
  FA_14515 \FA_INST_0[0].FA_INST_1[137].FA_  ( .A(A[137]), .B(n889), .CI(
        C[137]), .S(S[137]), .CO(C[138]) );
  FA_14514 \FA_INST_0[0].FA_INST_1[138].FA_  ( .A(A[138]), .B(n888), .CI(
        C[138]), .S(S[138]), .CO(C[139]) );
  FA_14513 \FA_INST_0[0].FA_INST_1[139].FA_  ( .A(A[139]), .B(n887), .CI(
        C[139]), .S(S[139]), .CO(C[140]) );
  FA_14512 \FA_INST_0[0].FA_INST_1[140].FA_  ( .A(A[140]), .B(n886), .CI(
        C[140]), .S(S[140]), .CO(C[141]) );
  FA_14511 \FA_INST_0[0].FA_INST_1[141].FA_  ( .A(A[141]), .B(n885), .CI(
        C[141]), .S(S[141]), .CO(C[142]) );
  FA_14510 \FA_INST_0[0].FA_INST_1[142].FA_  ( .A(A[142]), .B(n884), .CI(
        C[142]), .S(S[142]), .CO(C[143]) );
  FA_14509 \FA_INST_0[0].FA_INST_1[143].FA_  ( .A(A[143]), .B(n883), .CI(
        C[143]), .S(S[143]), .CO(C[144]) );
  FA_14508 \FA_INST_0[0].FA_INST_1[144].FA_  ( .A(A[144]), .B(n882), .CI(
        C[144]), .S(S[144]), .CO(C[145]) );
  FA_14507 \FA_INST_0[0].FA_INST_1[145].FA_  ( .A(A[145]), .B(n881), .CI(
        C[145]), .S(S[145]), .CO(C[146]) );
  FA_14506 \FA_INST_0[0].FA_INST_1[146].FA_  ( .A(A[146]), .B(n880), .CI(
        C[146]), .S(S[146]), .CO(C[147]) );
  FA_14505 \FA_INST_0[0].FA_INST_1[147].FA_  ( .A(A[147]), .B(n879), .CI(
        C[147]), .S(S[147]), .CO(C[148]) );
  FA_14504 \FA_INST_0[0].FA_INST_1[148].FA_  ( .A(A[148]), .B(n878), .CI(
        C[148]), .S(S[148]), .CO(C[149]) );
  FA_14503 \FA_INST_0[0].FA_INST_1[149].FA_  ( .A(A[149]), .B(n877), .CI(
        C[149]), .S(S[149]), .CO(C[150]) );
  FA_14502 \FA_INST_0[0].FA_INST_1[150].FA_  ( .A(A[150]), .B(n876), .CI(
        C[150]), .S(S[150]), .CO(C[151]) );
  FA_14501 \FA_INST_0[0].FA_INST_1[151].FA_  ( .A(A[151]), .B(n875), .CI(
        C[151]), .S(S[151]), .CO(C[152]) );
  FA_14500 \FA_INST_0[0].FA_INST_1[152].FA_  ( .A(A[152]), .B(n874), .CI(
        C[152]), .S(S[152]), .CO(C[153]) );
  FA_14499 \FA_INST_0[0].FA_INST_1[153].FA_  ( .A(A[153]), .B(n873), .CI(
        C[153]), .S(S[153]), .CO(C[154]) );
  FA_14498 \FA_INST_0[0].FA_INST_1[154].FA_  ( .A(A[154]), .B(n872), .CI(
        C[154]), .S(S[154]), .CO(C[155]) );
  FA_14497 \FA_INST_0[0].FA_INST_1[155].FA_  ( .A(A[155]), .B(n871), .CI(
        C[155]), .S(S[155]), .CO(C[156]) );
  FA_14496 \FA_INST_0[0].FA_INST_1[156].FA_  ( .A(A[156]), .B(n870), .CI(
        C[156]), .S(S[156]), .CO(C[157]) );
  FA_14495 \FA_INST_0[0].FA_INST_1[157].FA_  ( .A(A[157]), .B(n869), .CI(
        C[157]), .S(S[157]), .CO(C[158]) );
  FA_14494 \FA_INST_0[0].FA_INST_1[158].FA_  ( .A(A[158]), .B(n868), .CI(
        C[158]), .S(S[158]), .CO(C[159]) );
  FA_14493 \FA_INST_0[0].FA_INST_1[159].FA_  ( .A(A[159]), .B(n867), .CI(
        C[159]), .S(S[159]), .CO(C[160]) );
  FA_14492 \FA_INST_0[0].FA_INST_1[160].FA_  ( .A(A[160]), .B(n866), .CI(
        C[160]), .S(S[160]), .CO(C[161]) );
  FA_14491 \FA_INST_0[0].FA_INST_1[161].FA_  ( .A(A[161]), .B(n865), .CI(
        C[161]), .S(S[161]), .CO(C[162]) );
  FA_14490 \FA_INST_0[0].FA_INST_1[162].FA_  ( .A(A[162]), .B(n864), .CI(
        C[162]), .S(S[162]), .CO(C[163]) );
  FA_14489 \FA_INST_0[0].FA_INST_1[163].FA_  ( .A(A[163]), .B(n863), .CI(
        C[163]), .S(S[163]), .CO(C[164]) );
  FA_14488 \FA_INST_0[0].FA_INST_1[164].FA_  ( .A(A[164]), .B(n862), .CI(
        C[164]), .S(S[164]), .CO(C[165]) );
  FA_14487 \FA_INST_0[0].FA_INST_1[165].FA_  ( .A(A[165]), .B(n861), .CI(
        C[165]), .S(S[165]), .CO(C[166]) );
  FA_14486 \FA_INST_0[0].FA_INST_1[166].FA_  ( .A(A[166]), .B(n860), .CI(
        C[166]), .S(S[166]), .CO(C[167]) );
  FA_14485 \FA_INST_0[0].FA_INST_1[167].FA_  ( .A(A[167]), .B(n859), .CI(
        C[167]), .S(S[167]), .CO(C[168]) );
  FA_14484 \FA_INST_0[0].FA_INST_1[168].FA_  ( .A(A[168]), .B(n858), .CI(
        C[168]), .S(S[168]), .CO(C[169]) );
  FA_14483 \FA_INST_0[0].FA_INST_1[169].FA_  ( .A(A[169]), .B(n857), .CI(
        C[169]), .S(S[169]), .CO(C[170]) );
  FA_14482 \FA_INST_0[0].FA_INST_1[170].FA_  ( .A(A[170]), .B(n856), .CI(
        C[170]), .S(S[170]), .CO(C[171]) );
  FA_14481 \FA_INST_0[0].FA_INST_1[171].FA_  ( .A(A[171]), .B(n855), .CI(
        C[171]), .S(S[171]), .CO(C[172]) );
  FA_14480 \FA_INST_0[0].FA_INST_1[172].FA_  ( .A(A[172]), .B(n854), .CI(
        C[172]), .S(S[172]), .CO(C[173]) );
  FA_14479 \FA_INST_0[0].FA_INST_1[173].FA_  ( .A(A[173]), .B(n853), .CI(
        C[173]), .S(S[173]), .CO(C[174]) );
  FA_14478 \FA_INST_0[0].FA_INST_1[174].FA_  ( .A(A[174]), .B(n852), .CI(
        C[174]), .S(S[174]), .CO(C[175]) );
  FA_14477 \FA_INST_0[0].FA_INST_1[175].FA_  ( .A(A[175]), .B(n851), .CI(
        C[175]), .S(S[175]), .CO(C[176]) );
  FA_14476 \FA_INST_0[0].FA_INST_1[176].FA_  ( .A(A[176]), .B(n850), .CI(
        C[176]), .S(S[176]), .CO(C[177]) );
  FA_14475 \FA_INST_0[0].FA_INST_1[177].FA_  ( .A(A[177]), .B(n849), .CI(
        C[177]), .S(S[177]), .CO(C[178]) );
  FA_14474 \FA_INST_0[0].FA_INST_1[178].FA_  ( .A(A[178]), .B(n848), .CI(
        C[178]), .S(S[178]), .CO(C[179]) );
  FA_14473 \FA_INST_0[0].FA_INST_1[179].FA_  ( .A(A[179]), .B(n847), .CI(
        C[179]), .S(S[179]), .CO(C[180]) );
  FA_14472 \FA_INST_0[0].FA_INST_1[180].FA_  ( .A(A[180]), .B(n846), .CI(
        C[180]), .S(S[180]), .CO(C[181]) );
  FA_14471 \FA_INST_0[0].FA_INST_1[181].FA_  ( .A(A[181]), .B(n845), .CI(
        C[181]), .S(S[181]), .CO(C[182]) );
  FA_14470 \FA_INST_0[0].FA_INST_1[182].FA_  ( .A(A[182]), .B(n844), .CI(
        C[182]), .S(S[182]), .CO(C[183]) );
  FA_14469 \FA_INST_0[0].FA_INST_1[183].FA_  ( .A(A[183]), .B(n843), .CI(
        C[183]), .S(S[183]), .CO(C[184]) );
  FA_14468 \FA_INST_0[0].FA_INST_1[184].FA_  ( .A(A[184]), .B(n842), .CI(
        C[184]), .S(S[184]), .CO(C[185]) );
  FA_14467 \FA_INST_0[0].FA_INST_1[185].FA_  ( .A(A[185]), .B(n841), .CI(
        C[185]), .S(S[185]), .CO(C[186]) );
  FA_14466 \FA_INST_0[0].FA_INST_1[186].FA_  ( .A(A[186]), .B(n840), .CI(
        C[186]), .S(S[186]), .CO(C[187]) );
  FA_14465 \FA_INST_0[0].FA_INST_1[187].FA_  ( .A(A[187]), .B(n839), .CI(
        C[187]), .S(S[187]), .CO(C[188]) );
  FA_14464 \FA_INST_0[0].FA_INST_1[188].FA_  ( .A(A[188]), .B(n838), .CI(
        C[188]), .S(S[188]), .CO(C[189]) );
  FA_14463 \FA_INST_0[0].FA_INST_1[189].FA_  ( .A(A[189]), .B(n837), .CI(
        C[189]), .S(S[189]), .CO(C[190]) );
  FA_14462 \FA_INST_0[0].FA_INST_1[190].FA_  ( .A(A[190]), .B(n836), .CI(
        C[190]), .S(S[190]), .CO(C[191]) );
  FA_14461 \FA_INST_0[0].FA_INST_1[191].FA_  ( .A(A[191]), .B(n835), .CI(
        C[191]), .S(S[191]), .CO(C[192]) );
  FA_14460 \FA_INST_0[0].FA_INST_1[192].FA_  ( .A(A[192]), .B(n834), .CI(
        C[192]), .S(S[192]), .CO(C[193]) );
  FA_14459 \FA_INST_0[0].FA_INST_1[193].FA_  ( .A(A[193]), .B(n833), .CI(
        C[193]), .S(S[193]), .CO(C[194]) );
  FA_14458 \FA_INST_0[0].FA_INST_1[194].FA_  ( .A(A[194]), .B(n832), .CI(
        C[194]), .S(S[194]), .CO(C[195]) );
  FA_14457 \FA_INST_0[0].FA_INST_1[195].FA_  ( .A(A[195]), .B(n831), .CI(
        C[195]), .S(S[195]), .CO(C[196]) );
  FA_14456 \FA_INST_0[0].FA_INST_1[196].FA_  ( .A(A[196]), .B(n830), .CI(
        C[196]), .S(S[196]), .CO(C[197]) );
  FA_14455 \FA_INST_0[0].FA_INST_1[197].FA_  ( .A(A[197]), .B(n829), .CI(
        C[197]), .S(S[197]), .CO(C[198]) );
  FA_14454 \FA_INST_0[0].FA_INST_1[198].FA_  ( .A(A[198]), .B(n828), .CI(
        C[198]), .S(S[198]), .CO(C[199]) );
  FA_14453 \FA_INST_0[0].FA_INST_1[199].FA_  ( .A(A[199]), .B(n827), .CI(
        C[199]), .S(S[199]), .CO(C[200]) );
  FA_14452 \FA_INST_0[0].FA_INST_1[200].FA_  ( .A(A[200]), .B(n826), .CI(
        C[200]), .S(S[200]), .CO(C[201]) );
  FA_14451 \FA_INST_0[0].FA_INST_1[201].FA_  ( .A(A[201]), .B(n825), .CI(
        C[201]), .S(S[201]), .CO(C[202]) );
  FA_14450 \FA_INST_0[0].FA_INST_1[202].FA_  ( .A(A[202]), .B(n824), .CI(
        C[202]), .S(S[202]), .CO(C[203]) );
  FA_14449 \FA_INST_0[0].FA_INST_1[203].FA_  ( .A(A[203]), .B(n823), .CI(
        C[203]), .S(S[203]), .CO(C[204]) );
  FA_14448 \FA_INST_0[0].FA_INST_1[204].FA_  ( .A(A[204]), .B(n822), .CI(
        C[204]), .S(S[204]), .CO(C[205]) );
  FA_14447 \FA_INST_0[0].FA_INST_1[205].FA_  ( .A(A[205]), .B(n821), .CI(
        C[205]), .S(S[205]), .CO(C[206]) );
  FA_14446 \FA_INST_0[0].FA_INST_1[206].FA_  ( .A(A[206]), .B(n820), .CI(
        C[206]), .S(S[206]), .CO(C[207]) );
  FA_14445 \FA_INST_0[0].FA_INST_1[207].FA_  ( .A(A[207]), .B(n819), .CI(
        C[207]), .S(S[207]), .CO(C[208]) );
  FA_14444 \FA_INST_0[0].FA_INST_1[208].FA_  ( .A(A[208]), .B(n818), .CI(
        C[208]), .S(S[208]), .CO(C[209]) );
  FA_14443 \FA_INST_0[0].FA_INST_1[209].FA_  ( .A(A[209]), .B(n817), .CI(
        C[209]), .S(S[209]), .CO(C[210]) );
  FA_14442 \FA_INST_0[0].FA_INST_1[210].FA_  ( .A(A[210]), .B(n816), .CI(
        C[210]), .S(S[210]), .CO(C[211]) );
  FA_14441 \FA_INST_0[0].FA_INST_1[211].FA_  ( .A(A[211]), .B(n815), .CI(
        C[211]), .S(S[211]), .CO(C[212]) );
  FA_14440 \FA_INST_0[0].FA_INST_1[212].FA_  ( .A(A[212]), .B(n814), .CI(
        C[212]), .S(S[212]), .CO(C[213]) );
  FA_14439 \FA_INST_0[0].FA_INST_1[213].FA_  ( .A(A[213]), .B(n813), .CI(
        C[213]), .S(S[213]), .CO(C[214]) );
  FA_14438 \FA_INST_0[0].FA_INST_1[214].FA_  ( .A(A[214]), .B(n812), .CI(
        C[214]), .S(S[214]), .CO(C[215]) );
  FA_14437 \FA_INST_0[0].FA_INST_1[215].FA_  ( .A(A[215]), .B(n811), .CI(
        C[215]), .S(S[215]), .CO(C[216]) );
  FA_14436 \FA_INST_0[0].FA_INST_1[216].FA_  ( .A(A[216]), .B(n810), .CI(
        C[216]), .S(S[216]), .CO(C[217]) );
  FA_14435 \FA_INST_0[0].FA_INST_1[217].FA_  ( .A(A[217]), .B(n809), .CI(
        C[217]), .S(S[217]), .CO(C[218]) );
  FA_14434 \FA_INST_0[0].FA_INST_1[218].FA_  ( .A(A[218]), .B(n808), .CI(
        C[218]), .S(S[218]), .CO(C[219]) );
  FA_14433 \FA_INST_0[0].FA_INST_1[219].FA_  ( .A(A[219]), .B(n807), .CI(
        C[219]), .S(S[219]), .CO(C[220]) );
  FA_14432 \FA_INST_0[0].FA_INST_1[220].FA_  ( .A(A[220]), .B(n806), .CI(
        C[220]), .S(S[220]), .CO(C[221]) );
  FA_14431 \FA_INST_0[0].FA_INST_1[221].FA_  ( .A(A[221]), .B(n805), .CI(
        C[221]), .S(S[221]), .CO(C[222]) );
  FA_14430 \FA_INST_0[0].FA_INST_1[222].FA_  ( .A(A[222]), .B(n804), .CI(
        C[222]), .S(S[222]), .CO(C[223]) );
  FA_14429 \FA_INST_0[0].FA_INST_1[223].FA_  ( .A(A[223]), .B(n803), .CI(
        C[223]), .S(S[223]), .CO(C[224]) );
  FA_14428 \FA_INST_0[0].FA_INST_1[224].FA_  ( .A(A[224]), .B(n802), .CI(
        C[224]), .S(S[224]), .CO(C[225]) );
  FA_14427 \FA_INST_0[0].FA_INST_1[225].FA_  ( .A(A[225]), .B(n801), .CI(
        C[225]), .S(S[225]), .CO(C[226]) );
  FA_14426 \FA_INST_0[0].FA_INST_1[226].FA_  ( .A(A[226]), .B(n800), .CI(
        C[226]), .S(S[226]), .CO(C[227]) );
  FA_14425 \FA_INST_0[0].FA_INST_1[227].FA_  ( .A(A[227]), .B(n799), .CI(
        C[227]), .S(S[227]), .CO(C[228]) );
  FA_14424 \FA_INST_0[0].FA_INST_1[228].FA_  ( .A(A[228]), .B(n798), .CI(
        C[228]), .S(S[228]), .CO(C[229]) );
  FA_14423 \FA_INST_0[0].FA_INST_1[229].FA_  ( .A(A[229]), .B(n797), .CI(
        C[229]), .S(S[229]), .CO(C[230]) );
  FA_14422 \FA_INST_0[0].FA_INST_1[230].FA_  ( .A(A[230]), .B(n796), .CI(
        C[230]), .S(S[230]), .CO(C[231]) );
  FA_14421 \FA_INST_0[0].FA_INST_1[231].FA_  ( .A(A[231]), .B(n795), .CI(
        C[231]), .S(S[231]), .CO(C[232]) );
  FA_14420 \FA_INST_0[0].FA_INST_1[232].FA_  ( .A(A[232]), .B(n794), .CI(
        C[232]), .S(S[232]), .CO(C[233]) );
  FA_14419 \FA_INST_0[0].FA_INST_1[233].FA_  ( .A(A[233]), .B(n793), .CI(
        C[233]), .S(S[233]), .CO(C[234]) );
  FA_14418 \FA_INST_0[0].FA_INST_1[234].FA_  ( .A(A[234]), .B(n792), .CI(
        C[234]), .S(S[234]), .CO(C[235]) );
  FA_14417 \FA_INST_0[0].FA_INST_1[235].FA_  ( .A(A[235]), .B(n791), .CI(
        C[235]), .S(S[235]), .CO(C[236]) );
  FA_14416 \FA_INST_0[0].FA_INST_1[236].FA_  ( .A(A[236]), .B(n790), .CI(
        C[236]), .S(S[236]), .CO(C[237]) );
  FA_14415 \FA_INST_0[0].FA_INST_1[237].FA_  ( .A(A[237]), .B(n789), .CI(
        C[237]), .S(S[237]), .CO(C[238]) );
  FA_14414 \FA_INST_0[0].FA_INST_1[238].FA_  ( .A(A[238]), .B(n788), .CI(
        C[238]), .S(S[238]), .CO(C[239]) );
  FA_14413 \FA_INST_0[0].FA_INST_1[239].FA_  ( .A(A[239]), .B(n787), .CI(
        C[239]), .S(S[239]), .CO(C[240]) );
  FA_14412 \FA_INST_0[0].FA_INST_1[240].FA_  ( .A(A[240]), .B(n786), .CI(
        C[240]), .S(S[240]), .CO(C[241]) );
  FA_14411 \FA_INST_0[0].FA_INST_1[241].FA_  ( .A(A[241]), .B(n785), .CI(
        C[241]), .S(S[241]), .CO(C[242]) );
  FA_14410 \FA_INST_0[0].FA_INST_1[242].FA_  ( .A(A[242]), .B(n784), .CI(
        C[242]), .S(S[242]), .CO(C[243]) );
  FA_14409 \FA_INST_0[0].FA_INST_1[243].FA_  ( .A(A[243]), .B(n783), .CI(
        C[243]), .S(S[243]), .CO(C[244]) );
  FA_14408 \FA_INST_0[0].FA_INST_1[244].FA_  ( .A(A[244]), .B(n782), .CI(
        C[244]), .S(S[244]), .CO(C[245]) );
  FA_14407 \FA_INST_0[0].FA_INST_1[245].FA_  ( .A(A[245]), .B(n781), .CI(
        C[245]), .S(S[245]), .CO(C[246]) );
  FA_14406 \FA_INST_0[0].FA_INST_1[246].FA_  ( .A(A[246]), .B(n780), .CI(
        C[246]), .S(S[246]), .CO(C[247]) );
  FA_14405 \FA_INST_0[0].FA_INST_1[247].FA_  ( .A(A[247]), .B(n779), .CI(
        C[247]), .S(S[247]), .CO(C[248]) );
  FA_14404 \FA_INST_0[0].FA_INST_1[248].FA_  ( .A(A[248]), .B(n778), .CI(
        C[248]), .S(S[248]), .CO(C[249]) );
  FA_14403 \FA_INST_0[0].FA_INST_1[249].FA_  ( .A(A[249]), .B(n777), .CI(
        C[249]), .S(S[249]), .CO(C[250]) );
  FA_14402 \FA_INST_0[0].FA_INST_1[250].FA_  ( .A(A[250]), .B(n776), .CI(
        C[250]), .S(S[250]), .CO(C[251]) );
  FA_14401 \FA_INST_0[0].FA_INST_1[251].FA_  ( .A(A[251]), .B(n775), .CI(
        C[251]), .S(S[251]), .CO(C[252]) );
  FA_14400 \FA_INST_0[0].FA_INST_1[252].FA_  ( .A(A[252]), .B(n774), .CI(
        C[252]), .S(S[252]), .CO(C[253]) );
  FA_14399 \FA_INST_0[0].FA_INST_1[253].FA_  ( .A(A[253]), .B(n773), .CI(
        C[253]), .S(S[253]), .CO(C[254]) );
  FA_14398 \FA_INST_0[0].FA_INST_1[254].FA_  ( .A(A[254]), .B(n772), .CI(
        C[254]), .S(S[254]), .CO(C[255]) );
  FA_14397 \FA_INST_0[0].FA_INST_1[255].FA_  ( .A(A[255]), .B(n771), .CI(
        C[255]), .S(S[255]), .CO(C[256]) );
  FA_14396 \FA_INST_0[0].FA_INST_1[256].FA_  ( .A(A[256]), .B(n770), .CI(
        C[256]), .S(S[256]), .CO(C[257]) );
  FA_14395 \FA_INST_0[0].FA_INST_1[257].FA_  ( .A(A[257]), .B(n769), .CI(
        C[257]), .S(S[257]), .CO(C[258]) );
  FA_14394 \FA_INST_0[0].FA_INST_1[258].FA_  ( .A(A[258]), .B(n768), .CI(
        C[258]), .S(S[258]), .CO(C[259]) );
  FA_14393 \FA_INST_0[0].FA_INST_1[259].FA_  ( .A(A[259]), .B(n767), .CI(
        C[259]), .S(S[259]), .CO(C[260]) );
  FA_14392 \FA_INST_0[0].FA_INST_1[260].FA_  ( .A(A[260]), .B(n766), .CI(
        C[260]), .S(S[260]), .CO(C[261]) );
  FA_14391 \FA_INST_0[0].FA_INST_1[261].FA_  ( .A(A[261]), .B(n765), .CI(
        C[261]), .S(S[261]), .CO(C[262]) );
  FA_14390 \FA_INST_0[0].FA_INST_1[262].FA_  ( .A(A[262]), .B(n764), .CI(
        C[262]), .S(S[262]), .CO(C[263]) );
  FA_14389 \FA_INST_0[0].FA_INST_1[263].FA_  ( .A(A[263]), .B(n763), .CI(
        C[263]), .S(S[263]), .CO(C[264]) );
  FA_14388 \FA_INST_0[0].FA_INST_1[264].FA_  ( .A(A[264]), .B(n762), .CI(
        C[264]), .S(S[264]), .CO(C[265]) );
  FA_14387 \FA_INST_0[0].FA_INST_1[265].FA_  ( .A(A[265]), .B(n761), .CI(
        C[265]), .S(S[265]), .CO(C[266]) );
  FA_14386 \FA_INST_0[0].FA_INST_1[266].FA_  ( .A(A[266]), .B(n760), .CI(
        C[266]), .S(S[266]), .CO(C[267]) );
  FA_14385 \FA_INST_0[0].FA_INST_1[267].FA_  ( .A(A[267]), .B(n759), .CI(
        C[267]), .S(S[267]), .CO(C[268]) );
  FA_14384 \FA_INST_0[0].FA_INST_1[268].FA_  ( .A(A[268]), .B(n758), .CI(
        C[268]), .S(S[268]), .CO(C[269]) );
  FA_14383 \FA_INST_0[0].FA_INST_1[269].FA_  ( .A(A[269]), .B(n757), .CI(
        C[269]), .S(S[269]), .CO(C[270]) );
  FA_14382 \FA_INST_0[0].FA_INST_1[270].FA_  ( .A(A[270]), .B(n756), .CI(
        C[270]), .S(S[270]), .CO(C[271]) );
  FA_14381 \FA_INST_0[0].FA_INST_1[271].FA_  ( .A(A[271]), .B(n755), .CI(
        C[271]), .S(S[271]), .CO(C[272]) );
  FA_14380 \FA_INST_0[0].FA_INST_1[272].FA_  ( .A(A[272]), .B(n754), .CI(
        C[272]), .S(S[272]), .CO(C[273]) );
  FA_14379 \FA_INST_0[0].FA_INST_1[273].FA_  ( .A(A[273]), .B(n753), .CI(
        C[273]), .S(S[273]), .CO(C[274]) );
  FA_14378 \FA_INST_0[0].FA_INST_1[274].FA_  ( .A(A[274]), .B(n752), .CI(
        C[274]), .S(S[274]), .CO(C[275]) );
  FA_14377 \FA_INST_0[0].FA_INST_1[275].FA_  ( .A(A[275]), .B(n751), .CI(
        C[275]), .S(S[275]), .CO(C[276]) );
  FA_14376 \FA_INST_0[0].FA_INST_1[276].FA_  ( .A(A[276]), .B(n750), .CI(
        C[276]), .S(S[276]), .CO(C[277]) );
  FA_14375 \FA_INST_0[0].FA_INST_1[277].FA_  ( .A(A[277]), .B(n749), .CI(
        C[277]), .S(S[277]), .CO(C[278]) );
  FA_14374 \FA_INST_0[0].FA_INST_1[278].FA_  ( .A(A[278]), .B(n748), .CI(
        C[278]), .S(S[278]), .CO(C[279]) );
  FA_14373 \FA_INST_0[0].FA_INST_1[279].FA_  ( .A(A[279]), .B(n747), .CI(
        C[279]), .S(S[279]), .CO(C[280]) );
  FA_14372 \FA_INST_0[0].FA_INST_1[280].FA_  ( .A(A[280]), .B(n746), .CI(
        C[280]), .S(S[280]), .CO(C[281]) );
  FA_14371 \FA_INST_0[0].FA_INST_1[281].FA_  ( .A(A[281]), .B(n745), .CI(
        C[281]), .S(S[281]), .CO(C[282]) );
  FA_14370 \FA_INST_0[0].FA_INST_1[282].FA_  ( .A(A[282]), .B(n744), .CI(
        C[282]), .S(S[282]), .CO(C[283]) );
  FA_14369 \FA_INST_0[0].FA_INST_1[283].FA_  ( .A(A[283]), .B(n743), .CI(
        C[283]), .S(S[283]), .CO(C[284]) );
  FA_14368 \FA_INST_0[0].FA_INST_1[284].FA_  ( .A(A[284]), .B(n742), .CI(
        C[284]), .S(S[284]), .CO(C[285]) );
  FA_14367 \FA_INST_0[0].FA_INST_1[285].FA_  ( .A(A[285]), .B(n741), .CI(
        C[285]), .S(S[285]), .CO(C[286]) );
  FA_14366 \FA_INST_0[0].FA_INST_1[286].FA_  ( .A(A[286]), .B(n740), .CI(
        C[286]), .S(S[286]), .CO(C[287]) );
  FA_14365 \FA_INST_0[0].FA_INST_1[287].FA_  ( .A(A[287]), .B(n739), .CI(
        C[287]), .S(S[287]), .CO(C[288]) );
  FA_14364 \FA_INST_0[0].FA_INST_1[288].FA_  ( .A(A[288]), .B(n738), .CI(
        C[288]), .S(S[288]), .CO(C[289]) );
  FA_14363 \FA_INST_0[0].FA_INST_1[289].FA_  ( .A(A[289]), .B(n737), .CI(
        C[289]), .S(S[289]), .CO(C[290]) );
  FA_14362 \FA_INST_0[0].FA_INST_1[290].FA_  ( .A(A[290]), .B(n736), .CI(
        C[290]), .S(S[290]), .CO(C[291]) );
  FA_14361 \FA_INST_0[0].FA_INST_1[291].FA_  ( .A(A[291]), .B(n735), .CI(
        C[291]), .S(S[291]), .CO(C[292]) );
  FA_14360 \FA_INST_0[0].FA_INST_1[292].FA_  ( .A(A[292]), .B(n734), .CI(
        C[292]), .S(S[292]), .CO(C[293]) );
  FA_14359 \FA_INST_0[0].FA_INST_1[293].FA_  ( .A(A[293]), .B(n733), .CI(
        C[293]), .S(S[293]), .CO(C[294]) );
  FA_14358 \FA_INST_0[0].FA_INST_1[294].FA_  ( .A(A[294]), .B(n732), .CI(
        C[294]), .S(S[294]), .CO(C[295]) );
  FA_14357 \FA_INST_0[0].FA_INST_1[295].FA_  ( .A(A[295]), .B(n731), .CI(
        C[295]), .S(S[295]), .CO(C[296]) );
  FA_14356 \FA_INST_0[0].FA_INST_1[296].FA_  ( .A(A[296]), .B(n730), .CI(
        C[296]), .S(S[296]), .CO(C[297]) );
  FA_14355 \FA_INST_0[0].FA_INST_1[297].FA_  ( .A(A[297]), .B(n729), .CI(
        C[297]), .S(S[297]), .CO(C[298]) );
  FA_14354 \FA_INST_0[0].FA_INST_1[298].FA_  ( .A(A[298]), .B(n728), .CI(
        C[298]), .S(S[298]), .CO(C[299]) );
  FA_14353 \FA_INST_0[0].FA_INST_1[299].FA_  ( .A(A[299]), .B(n727), .CI(
        C[299]), .S(S[299]), .CO(C[300]) );
  FA_14352 \FA_INST_0[0].FA_INST_1[300].FA_  ( .A(A[300]), .B(n726), .CI(
        C[300]), .S(S[300]), .CO(C[301]) );
  FA_14351 \FA_INST_0[0].FA_INST_1[301].FA_  ( .A(A[301]), .B(n725), .CI(
        C[301]), .S(S[301]), .CO(C[302]) );
  FA_14350 \FA_INST_0[0].FA_INST_1[302].FA_  ( .A(A[302]), .B(n724), .CI(
        C[302]), .S(S[302]), .CO(C[303]) );
  FA_14349 \FA_INST_0[0].FA_INST_1[303].FA_  ( .A(A[303]), .B(n723), .CI(
        C[303]), .S(S[303]), .CO(C[304]) );
  FA_14348 \FA_INST_0[0].FA_INST_1[304].FA_  ( .A(A[304]), .B(n722), .CI(
        C[304]), .S(S[304]), .CO(C[305]) );
  FA_14347 \FA_INST_0[0].FA_INST_1[305].FA_  ( .A(A[305]), .B(n721), .CI(
        C[305]), .S(S[305]), .CO(C[306]) );
  FA_14346 \FA_INST_0[0].FA_INST_1[306].FA_  ( .A(A[306]), .B(n720), .CI(
        C[306]), .S(S[306]), .CO(C[307]) );
  FA_14345 \FA_INST_0[0].FA_INST_1[307].FA_  ( .A(A[307]), .B(n719), .CI(
        C[307]), .S(S[307]), .CO(C[308]) );
  FA_14344 \FA_INST_0[0].FA_INST_1[308].FA_  ( .A(A[308]), .B(n718), .CI(
        C[308]), .S(S[308]), .CO(C[309]) );
  FA_14343 \FA_INST_0[0].FA_INST_1[309].FA_  ( .A(A[309]), .B(n717), .CI(
        C[309]), .S(S[309]), .CO(C[310]) );
  FA_14342 \FA_INST_0[0].FA_INST_1[310].FA_  ( .A(A[310]), .B(n716), .CI(
        C[310]), .S(S[310]), .CO(C[311]) );
  FA_14341 \FA_INST_0[0].FA_INST_1[311].FA_  ( .A(A[311]), .B(n715), .CI(
        C[311]), .S(S[311]), .CO(C[312]) );
  FA_14340 \FA_INST_0[0].FA_INST_1[312].FA_  ( .A(A[312]), .B(n714), .CI(
        C[312]), .S(S[312]), .CO(C[313]) );
  FA_14339 \FA_INST_0[0].FA_INST_1[313].FA_  ( .A(A[313]), .B(n713), .CI(
        C[313]), .S(S[313]), .CO(C[314]) );
  FA_14338 \FA_INST_0[0].FA_INST_1[314].FA_  ( .A(A[314]), .B(n712), .CI(
        C[314]), .S(S[314]), .CO(C[315]) );
  FA_14337 \FA_INST_0[0].FA_INST_1[315].FA_  ( .A(A[315]), .B(n711), .CI(
        C[315]), .S(S[315]), .CO(C[316]) );
  FA_14336 \FA_INST_0[0].FA_INST_1[316].FA_  ( .A(A[316]), .B(n710), .CI(
        C[316]), .S(S[316]), .CO(C[317]) );
  FA_14335 \FA_INST_0[0].FA_INST_1[317].FA_  ( .A(A[317]), .B(n709), .CI(
        C[317]), .S(S[317]), .CO(C[318]) );
  FA_14334 \FA_INST_0[0].FA_INST_1[318].FA_  ( .A(A[318]), .B(n708), .CI(
        C[318]), .S(S[318]), .CO(C[319]) );
  FA_14333 \FA_INST_0[0].FA_INST_1[319].FA_  ( .A(A[319]), .B(n707), .CI(
        C[319]), .S(S[319]), .CO(C[320]) );
  FA_14332 \FA_INST_0[0].FA_INST_1[320].FA_  ( .A(A[320]), .B(n706), .CI(
        C[320]), .S(S[320]), .CO(C[321]) );
  FA_14331 \FA_INST_0[0].FA_INST_1[321].FA_  ( .A(A[321]), .B(n705), .CI(
        C[321]), .S(S[321]), .CO(C[322]) );
  FA_14330 \FA_INST_0[0].FA_INST_1[322].FA_  ( .A(A[322]), .B(n704), .CI(
        C[322]), .S(S[322]), .CO(C[323]) );
  FA_14329 \FA_INST_0[0].FA_INST_1[323].FA_  ( .A(A[323]), .B(n703), .CI(
        C[323]), .S(S[323]), .CO(C[324]) );
  FA_14328 \FA_INST_0[0].FA_INST_1[324].FA_  ( .A(A[324]), .B(n702), .CI(
        C[324]), .S(S[324]), .CO(C[325]) );
  FA_14327 \FA_INST_0[0].FA_INST_1[325].FA_  ( .A(A[325]), .B(n701), .CI(
        C[325]), .S(S[325]), .CO(C[326]) );
  FA_14326 \FA_INST_0[0].FA_INST_1[326].FA_  ( .A(A[326]), .B(n700), .CI(
        C[326]), .S(S[326]), .CO(C[327]) );
  FA_14325 \FA_INST_0[0].FA_INST_1[327].FA_  ( .A(A[327]), .B(n699), .CI(
        C[327]), .S(S[327]), .CO(C[328]) );
  FA_14324 \FA_INST_0[0].FA_INST_1[328].FA_  ( .A(A[328]), .B(n698), .CI(
        C[328]), .S(S[328]), .CO(C[329]) );
  FA_14323 \FA_INST_0[0].FA_INST_1[329].FA_  ( .A(A[329]), .B(n697), .CI(
        C[329]), .S(S[329]), .CO(C[330]) );
  FA_14322 \FA_INST_0[0].FA_INST_1[330].FA_  ( .A(A[330]), .B(n696), .CI(
        C[330]), .S(S[330]), .CO(C[331]) );
  FA_14321 \FA_INST_0[0].FA_INST_1[331].FA_  ( .A(A[331]), .B(n695), .CI(
        C[331]), .S(S[331]), .CO(C[332]) );
  FA_14320 \FA_INST_0[0].FA_INST_1[332].FA_  ( .A(A[332]), .B(n694), .CI(
        C[332]), .S(S[332]), .CO(C[333]) );
  FA_14319 \FA_INST_0[0].FA_INST_1[333].FA_  ( .A(A[333]), .B(n693), .CI(
        C[333]), .S(S[333]), .CO(C[334]) );
  FA_14318 \FA_INST_0[0].FA_INST_1[334].FA_  ( .A(A[334]), .B(n692), .CI(
        C[334]), .S(S[334]), .CO(C[335]) );
  FA_14317 \FA_INST_0[0].FA_INST_1[335].FA_  ( .A(A[335]), .B(n691), .CI(
        C[335]), .S(S[335]), .CO(C[336]) );
  FA_14316 \FA_INST_0[0].FA_INST_1[336].FA_  ( .A(A[336]), .B(n690), .CI(
        C[336]), .S(S[336]), .CO(C[337]) );
  FA_14315 \FA_INST_0[0].FA_INST_1[337].FA_  ( .A(A[337]), .B(n689), .CI(
        C[337]), .S(S[337]), .CO(C[338]) );
  FA_14314 \FA_INST_0[0].FA_INST_1[338].FA_  ( .A(A[338]), .B(n688), .CI(
        C[338]), .S(S[338]), .CO(C[339]) );
  FA_14313 \FA_INST_0[0].FA_INST_1[339].FA_  ( .A(A[339]), .B(n687), .CI(
        C[339]), .S(S[339]), .CO(C[340]) );
  FA_14312 \FA_INST_0[0].FA_INST_1[340].FA_  ( .A(A[340]), .B(n686), .CI(
        C[340]), .S(S[340]), .CO(C[341]) );
  FA_14311 \FA_INST_0[0].FA_INST_1[341].FA_  ( .A(A[341]), .B(n685), .CI(
        C[341]), .S(S[341]), .CO(C[342]) );
  FA_14310 \FA_INST_0[0].FA_INST_1[342].FA_  ( .A(A[342]), .B(n684), .CI(
        C[342]), .S(S[342]), .CO(C[343]) );
  FA_14309 \FA_INST_0[0].FA_INST_1[343].FA_  ( .A(A[343]), .B(n683), .CI(
        C[343]), .S(S[343]), .CO(C[344]) );
  FA_14308 \FA_INST_0[0].FA_INST_1[344].FA_  ( .A(A[344]), .B(n682), .CI(
        C[344]), .S(S[344]), .CO(C[345]) );
  FA_14307 \FA_INST_0[0].FA_INST_1[345].FA_  ( .A(A[345]), .B(n681), .CI(
        C[345]), .S(S[345]), .CO(C[346]) );
  FA_14306 \FA_INST_0[0].FA_INST_1[346].FA_  ( .A(A[346]), .B(n680), .CI(
        C[346]), .S(S[346]), .CO(C[347]) );
  FA_14305 \FA_INST_0[0].FA_INST_1[347].FA_  ( .A(A[347]), .B(n679), .CI(
        C[347]), .S(S[347]), .CO(C[348]) );
  FA_14304 \FA_INST_0[0].FA_INST_1[348].FA_  ( .A(A[348]), .B(n678), .CI(
        C[348]), .S(S[348]), .CO(C[349]) );
  FA_14303 \FA_INST_0[0].FA_INST_1[349].FA_  ( .A(A[349]), .B(n677), .CI(
        C[349]), .S(S[349]), .CO(C[350]) );
  FA_14302 \FA_INST_0[0].FA_INST_1[350].FA_  ( .A(A[350]), .B(n676), .CI(
        C[350]), .S(S[350]), .CO(C[351]) );
  FA_14301 \FA_INST_0[0].FA_INST_1[351].FA_  ( .A(A[351]), .B(n675), .CI(
        C[351]), .S(S[351]), .CO(C[352]) );
  FA_14300 \FA_INST_0[0].FA_INST_1[352].FA_  ( .A(A[352]), .B(n674), .CI(
        C[352]), .S(S[352]), .CO(C[353]) );
  FA_14299 \FA_INST_0[0].FA_INST_1[353].FA_  ( .A(A[353]), .B(n673), .CI(
        C[353]), .S(S[353]), .CO(C[354]) );
  FA_14298 \FA_INST_0[0].FA_INST_1[354].FA_  ( .A(A[354]), .B(n672), .CI(
        C[354]), .S(S[354]), .CO(C[355]) );
  FA_14297 \FA_INST_0[0].FA_INST_1[355].FA_  ( .A(A[355]), .B(n671), .CI(
        C[355]), .S(S[355]), .CO(C[356]) );
  FA_14296 \FA_INST_0[0].FA_INST_1[356].FA_  ( .A(A[356]), .B(n670), .CI(
        C[356]), .S(S[356]), .CO(C[357]) );
  FA_14295 \FA_INST_0[0].FA_INST_1[357].FA_  ( .A(A[357]), .B(n669), .CI(
        C[357]), .S(S[357]), .CO(C[358]) );
  FA_14294 \FA_INST_0[0].FA_INST_1[358].FA_  ( .A(A[358]), .B(n668), .CI(
        C[358]), .S(S[358]), .CO(C[359]) );
  FA_14293 \FA_INST_0[0].FA_INST_1[359].FA_  ( .A(A[359]), .B(n667), .CI(
        C[359]), .S(S[359]), .CO(C[360]) );
  FA_14292 \FA_INST_0[0].FA_INST_1[360].FA_  ( .A(A[360]), .B(n666), .CI(
        C[360]), .S(S[360]), .CO(C[361]) );
  FA_14291 \FA_INST_0[0].FA_INST_1[361].FA_  ( .A(A[361]), .B(n665), .CI(
        C[361]), .S(S[361]), .CO(C[362]) );
  FA_14290 \FA_INST_0[0].FA_INST_1[362].FA_  ( .A(A[362]), .B(n664), .CI(
        C[362]), .S(S[362]), .CO(C[363]) );
  FA_14289 \FA_INST_0[0].FA_INST_1[363].FA_  ( .A(A[363]), .B(n663), .CI(
        C[363]), .S(S[363]), .CO(C[364]) );
  FA_14288 \FA_INST_0[0].FA_INST_1[364].FA_  ( .A(A[364]), .B(n662), .CI(
        C[364]), .S(S[364]), .CO(C[365]) );
  FA_14287 \FA_INST_0[0].FA_INST_1[365].FA_  ( .A(A[365]), .B(n661), .CI(
        C[365]), .S(S[365]), .CO(C[366]) );
  FA_14286 \FA_INST_0[0].FA_INST_1[366].FA_  ( .A(A[366]), .B(n660), .CI(
        C[366]), .S(S[366]), .CO(C[367]) );
  FA_14285 \FA_INST_0[0].FA_INST_1[367].FA_  ( .A(A[367]), .B(n659), .CI(
        C[367]), .S(S[367]), .CO(C[368]) );
  FA_14284 \FA_INST_0[0].FA_INST_1[368].FA_  ( .A(A[368]), .B(n658), .CI(
        C[368]), .S(S[368]), .CO(C[369]) );
  FA_14283 \FA_INST_0[0].FA_INST_1[369].FA_  ( .A(A[369]), .B(n657), .CI(
        C[369]), .S(S[369]), .CO(C[370]) );
  FA_14282 \FA_INST_0[0].FA_INST_1[370].FA_  ( .A(A[370]), .B(n656), .CI(
        C[370]), .S(S[370]), .CO(C[371]) );
  FA_14281 \FA_INST_0[0].FA_INST_1[371].FA_  ( .A(A[371]), .B(n655), .CI(
        C[371]), .S(S[371]), .CO(C[372]) );
  FA_14280 \FA_INST_0[0].FA_INST_1[372].FA_  ( .A(A[372]), .B(n654), .CI(
        C[372]), .S(S[372]), .CO(C[373]) );
  FA_14279 \FA_INST_0[0].FA_INST_1[373].FA_  ( .A(A[373]), .B(n653), .CI(
        C[373]), .S(S[373]), .CO(C[374]) );
  FA_14278 \FA_INST_0[0].FA_INST_1[374].FA_  ( .A(A[374]), .B(n652), .CI(
        C[374]), .S(S[374]), .CO(C[375]) );
  FA_14277 \FA_INST_0[0].FA_INST_1[375].FA_  ( .A(A[375]), .B(n651), .CI(
        C[375]), .S(S[375]), .CO(C[376]) );
  FA_14276 \FA_INST_0[0].FA_INST_1[376].FA_  ( .A(A[376]), .B(n650), .CI(
        C[376]), .S(S[376]), .CO(C[377]) );
  FA_14275 \FA_INST_0[0].FA_INST_1[377].FA_  ( .A(A[377]), .B(n649), .CI(
        C[377]), .S(S[377]), .CO(C[378]) );
  FA_14274 \FA_INST_0[0].FA_INST_1[378].FA_  ( .A(A[378]), .B(n648), .CI(
        C[378]), .S(S[378]), .CO(C[379]) );
  FA_14273 \FA_INST_0[0].FA_INST_1[379].FA_  ( .A(A[379]), .B(n647), .CI(
        C[379]), .S(S[379]), .CO(C[380]) );
  FA_14272 \FA_INST_0[0].FA_INST_1[380].FA_  ( .A(A[380]), .B(n646), .CI(
        C[380]), .S(S[380]), .CO(C[381]) );
  FA_14271 \FA_INST_0[0].FA_INST_1[381].FA_  ( .A(A[381]), .B(n645), .CI(
        C[381]), .S(S[381]), .CO(C[382]) );
  FA_14270 \FA_INST_0[0].FA_INST_1[382].FA_  ( .A(A[382]), .B(n644), .CI(
        C[382]), .S(S[382]), .CO(C[383]) );
  FA_14269 \FA_INST_0[0].FA_INST_1[383].FA_  ( .A(A[383]), .B(n643), .CI(
        C[383]), .S(S[383]), .CO(C[384]) );
  FA_14268 \FA_INST_0[0].FA_INST_1[384].FA_  ( .A(A[384]), .B(n642), .CI(
        C[384]), .S(S[384]), .CO(C[385]) );
  FA_14267 \FA_INST_0[0].FA_INST_1[385].FA_  ( .A(A[385]), .B(n641), .CI(
        C[385]), .S(S[385]), .CO(C[386]) );
  FA_14266 \FA_INST_0[0].FA_INST_1[386].FA_  ( .A(A[386]), .B(n640), .CI(
        C[386]), .S(S[386]), .CO(C[387]) );
  FA_14265 \FA_INST_0[0].FA_INST_1[387].FA_  ( .A(A[387]), .B(n639), .CI(
        C[387]), .S(S[387]), .CO(C[388]) );
  FA_14264 \FA_INST_0[0].FA_INST_1[388].FA_  ( .A(A[388]), .B(n638), .CI(
        C[388]), .S(S[388]), .CO(C[389]) );
  FA_14263 \FA_INST_0[0].FA_INST_1[389].FA_  ( .A(A[389]), .B(n637), .CI(
        C[389]), .S(S[389]), .CO(C[390]) );
  FA_14262 \FA_INST_0[0].FA_INST_1[390].FA_  ( .A(A[390]), .B(n636), .CI(
        C[390]), .S(S[390]), .CO(C[391]) );
  FA_14261 \FA_INST_0[0].FA_INST_1[391].FA_  ( .A(A[391]), .B(n635), .CI(
        C[391]), .S(S[391]), .CO(C[392]) );
  FA_14260 \FA_INST_0[0].FA_INST_1[392].FA_  ( .A(A[392]), .B(n634), .CI(
        C[392]), .S(S[392]), .CO(C[393]) );
  FA_14259 \FA_INST_0[0].FA_INST_1[393].FA_  ( .A(A[393]), .B(n633), .CI(
        C[393]), .S(S[393]), .CO(C[394]) );
  FA_14258 \FA_INST_0[0].FA_INST_1[394].FA_  ( .A(A[394]), .B(n632), .CI(
        C[394]), .S(S[394]), .CO(C[395]) );
  FA_14257 \FA_INST_0[0].FA_INST_1[395].FA_  ( .A(A[395]), .B(n631), .CI(
        C[395]), .S(S[395]), .CO(C[396]) );
  FA_14256 \FA_INST_0[0].FA_INST_1[396].FA_  ( .A(A[396]), .B(n630), .CI(
        C[396]), .S(S[396]), .CO(C[397]) );
  FA_14255 \FA_INST_0[0].FA_INST_1[397].FA_  ( .A(A[397]), .B(n629), .CI(
        C[397]), .S(S[397]), .CO(C[398]) );
  FA_14254 \FA_INST_0[0].FA_INST_1[398].FA_  ( .A(A[398]), .B(n628), .CI(
        C[398]), .S(S[398]), .CO(C[399]) );
  FA_14253 \FA_INST_0[0].FA_INST_1[399].FA_  ( .A(A[399]), .B(n627), .CI(
        C[399]), .S(S[399]), .CO(C[400]) );
  FA_14252 \FA_INST_0[0].FA_INST_1[400].FA_  ( .A(A[400]), .B(n626), .CI(
        C[400]), .S(S[400]), .CO(C[401]) );
  FA_14251 \FA_INST_0[0].FA_INST_1[401].FA_  ( .A(A[401]), .B(n625), .CI(
        C[401]), .S(S[401]), .CO(C[402]) );
  FA_14250 \FA_INST_0[0].FA_INST_1[402].FA_  ( .A(A[402]), .B(n624), .CI(
        C[402]), .S(S[402]), .CO(C[403]) );
  FA_14249 \FA_INST_0[0].FA_INST_1[403].FA_  ( .A(A[403]), .B(n623), .CI(
        C[403]), .S(S[403]), .CO(C[404]) );
  FA_14248 \FA_INST_0[0].FA_INST_1[404].FA_  ( .A(A[404]), .B(n622), .CI(
        C[404]), .S(S[404]), .CO(C[405]) );
  FA_14247 \FA_INST_0[0].FA_INST_1[405].FA_  ( .A(A[405]), .B(n621), .CI(
        C[405]), .S(S[405]), .CO(C[406]) );
  FA_14246 \FA_INST_0[0].FA_INST_1[406].FA_  ( .A(A[406]), .B(n620), .CI(
        C[406]), .S(S[406]), .CO(C[407]) );
  FA_14245 \FA_INST_0[0].FA_INST_1[407].FA_  ( .A(A[407]), .B(n619), .CI(
        C[407]), .S(S[407]), .CO(C[408]) );
  FA_14244 \FA_INST_0[0].FA_INST_1[408].FA_  ( .A(A[408]), .B(n618), .CI(
        C[408]), .S(S[408]), .CO(C[409]) );
  FA_14243 \FA_INST_0[0].FA_INST_1[409].FA_  ( .A(A[409]), .B(n617), .CI(
        C[409]), .S(S[409]), .CO(C[410]) );
  FA_14242 \FA_INST_0[0].FA_INST_1[410].FA_  ( .A(A[410]), .B(n616), .CI(
        C[410]), .S(S[410]), .CO(C[411]) );
  FA_14241 \FA_INST_0[0].FA_INST_1[411].FA_  ( .A(A[411]), .B(n615), .CI(
        C[411]), .S(S[411]), .CO(C[412]) );
  FA_14240 \FA_INST_0[0].FA_INST_1[412].FA_  ( .A(A[412]), .B(n614), .CI(
        C[412]), .S(S[412]), .CO(C[413]) );
  FA_14239 \FA_INST_0[0].FA_INST_1[413].FA_  ( .A(A[413]), .B(n613), .CI(
        C[413]), .S(S[413]), .CO(C[414]) );
  FA_14238 \FA_INST_0[0].FA_INST_1[414].FA_  ( .A(A[414]), .B(n612), .CI(
        C[414]), .S(S[414]), .CO(C[415]) );
  FA_14237 \FA_INST_0[0].FA_INST_1[415].FA_  ( .A(A[415]), .B(n611), .CI(
        C[415]), .S(S[415]), .CO(C[416]) );
  FA_14236 \FA_INST_0[0].FA_INST_1[416].FA_  ( .A(A[416]), .B(n610), .CI(
        C[416]), .S(S[416]), .CO(C[417]) );
  FA_14235 \FA_INST_0[0].FA_INST_1[417].FA_  ( .A(A[417]), .B(n609), .CI(
        C[417]), .S(S[417]), .CO(C[418]) );
  FA_14234 \FA_INST_0[0].FA_INST_1[418].FA_  ( .A(A[418]), .B(n608), .CI(
        C[418]), .S(S[418]), .CO(C[419]) );
  FA_14233 \FA_INST_0[0].FA_INST_1[419].FA_  ( .A(A[419]), .B(n607), .CI(
        C[419]), .S(S[419]), .CO(C[420]) );
  FA_14232 \FA_INST_0[0].FA_INST_1[420].FA_  ( .A(A[420]), .B(n606), .CI(
        C[420]), .S(S[420]), .CO(C[421]) );
  FA_14231 \FA_INST_0[0].FA_INST_1[421].FA_  ( .A(A[421]), .B(n605), .CI(
        C[421]), .S(S[421]), .CO(C[422]) );
  FA_14230 \FA_INST_0[0].FA_INST_1[422].FA_  ( .A(A[422]), .B(n604), .CI(
        C[422]), .S(S[422]), .CO(C[423]) );
  FA_14229 \FA_INST_0[0].FA_INST_1[423].FA_  ( .A(A[423]), .B(n603), .CI(
        C[423]), .S(S[423]), .CO(C[424]) );
  FA_14228 \FA_INST_0[0].FA_INST_1[424].FA_  ( .A(A[424]), .B(n602), .CI(
        C[424]), .S(S[424]), .CO(C[425]) );
  FA_14227 \FA_INST_0[0].FA_INST_1[425].FA_  ( .A(A[425]), .B(n601), .CI(
        C[425]), .S(S[425]), .CO(C[426]) );
  FA_14226 \FA_INST_0[0].FA_INST_1[426].FA_  ( .A(A[426]), .B(n600), .CI(
        C[426]), .S(S[426]), .CO(C[427]) );
  FA_14225 \FA_INST_0[0].FA_INST_1[427].FA_  ( .A(A[427]), .B(n599), .CI(
        C[427]), .S(S[427]), .CO(C[428]) );
  FA_14224 \FA_INST_0[0].FA_INST_1[428].FA_  ( .A(A[428]), .B(n598), .CI(
        C[428]), .S(S[428]), .CO(C[429]) );
  FA_14223 \FA_INST_0[0].FA_INST_1[429].FA_  ( .A(A[429]), .B(n597), .CI(
        C[429]), .S(S[429]), .CO(C[430]) );
  FA_14222 \FA_INST_0[0].FA_INST_1[430].FA_  ( .A(A[430]), .B(n596), .CI(
        C[430]), .S(S[430]), .CO(C[431]) );
  FA_14221 \FA_INST_0[0].FA_INST_1[431].FA_  ( .A(A[431]), .B(n595), .CI(
        C[431]), .S(S[431]), .CO(C[432]) );
  FA_14220 \FA_INST_0[0].FA_INST_1[432].FA_  ( .A(A[432]), .B(n594), .CI(
        C[432]), .S(S[432]), .CO(C[433]) );
  FA_14219 \FA_INST_0[0].FA_INST_1[433].FA_  ( .A(A[433]), .B(n593), .CI(
        C[433]), .S(S[433]), .CO(C[434]) );
  FA_14218 \FA_INST_0[0].FA_INST_1[434].FA_  ( .A(A[434]), .B(n592), .CI(
        C[434]), .S(S[434]), .CO(C[435]) );
  FA_14217 \FA_INST_0[0].FA_INST_1[435].FA_  ( .A(A[435]), .B(n591), .CI(
        C[435]), .S(S[435]), .CO(C[436]) );
  FA_14216 \FA_INST_0[0].FA_INST_1[436].FA_  ( .A(A[436]), .B(n590), .CI(
        C[436]), .S(S[436]), .CO(C[437]) );
  FA_14215 \FA_INST_0[0].FA_INST_1[437].FA_  ( .A(A[437]), .B(n589), .CI(
        C[437]), .S(S[437]), .CO(C[438]) );
  FA_14214 \FA_INST_0[0].FA_INST_1[438].FA_  ( .A(A[438]), .B(n588), .CI(
        C[438]), .S(S[438]), .CO(C[439]) );
  FA_14213 \FA_INST_0[0].FA_INST_1[439].FA_  ( .A(A[439]), .B(n587), .CI(
        C[439]), .S(S[439]), .CO(C[440]) );
  FA_14212 \FA_INST_0[0].FA_INST_1[440].FA_  ( .A(A[440]), .B(n586), .CI(
        C[440]), .S(S[440]), .CO(C[441]) );
  FA_14211 \FA_INST_0[0].FA_INST_1[441].FA_  ( .A(A[441]), .B(n585), .CI(
        C[441]), .S(S[441]), .CO(C[442]) );
  FA_14210 \FA_INST_0[0].FA_INST_1[442].FA_  ( .A(A[442]), .B(n584), .CI(
        C[442]), .S(S[442]), .CO(C[443]) );
  FA_14209 \FA_INST_0[0].FA_INST_1[443].FA_  ( .A(A[443]), .B(n583), .CI(
        C[443]), .S(S[443]), .CO(C[444]) );
  FA_14208 \FA_INST_0[0].FA_INST_1[444].FA_  ( .A(A[444]), .B(n582), .CI(
        C[444]), .S(S[444]), .CO(C[445]) );
  FA_14207 \FA_INST_0[0].FA_INST_1[445].FA_  ( .A(A[445]), .B(n581), .CI(
        C[445]), .S(S[445]), .CO(C[446]) );
  FA_14206 \FA_INST_0[0].FA_INST_1[446].FA_  ( .A(A[446]), .B(n580), .CI(
        C[446]), .S(S[446]), .CO(C[447]) );
  FA_14205 \FA_INST_0[0].FA_INST_1[447].FA_  ( .A(A[447]), .B(n579), .CI(
        C[447]), .S(S[447]), .CO(C[448]) );
  FA_14204 \FA_INST_0[0].FA_INST_1[448].FA_  ( .A(A[448]), .B(n578), .CI(
        C[448]), .S(S[448]), .CO(C[449]) );
  FA_14203 \FA_INST_0[0].FA_INST_1[449].FA_  ( .A(A[449]), .B(n577), .CI(
        C[449]), .S(S[449]), .CO(C[450]) );
  FA_14202 \FA_INST_0[0].FA_INST_1[450].FA_  ( .A(A[450]), .B(n576), .CI(
        C[450]), .S(S[450]), .CO(C[451]) );
  FA_14201 \FA_INST_0[0].FA_INST_1[451].FA_  ( .A(A[451]), .B(n575), .CI(
        C[451]), .S(S[451]), .CO(C[452]) );
  FA_14200 \FA_INST_0[0].FA_INST_1[452].FA_  ( .A(A[452]), .B(n574), .CI(
        C[452]), .S(S[452]), .CO(C[453]) );
  FA_14199 \FA_INST_0[0].FA_INST_1[453].FA_  ( .A(A[453]), .B(n573), .CI(
        C[453]), .S(S[453]), .CO(C[454]) );
  FA_14198 \FA_INST_0[0].FA_INST_1[454].FA_  ( .A(A[454]), .B(n572), .CI(
        C[454]), .S(S[454]), .CO(C[455]) );
  FA_14197 \FA_INST_0[0].FA_INST_1[455].FA_  ( .A(A[455]), .B(n571), .CI(
        C[455]), .S(S[455]), .CO(C[456]) );
  FA_14196 \FA_INST_0[0].FA_INST_1[456].FA_  ( .A(A[456]), .B(n570), .CI(
        C[456]), .S(S[456]), .CO(C[457]) );
  FA_14195 \FA_INST_0[0].FA_INST_1[457].FA_  ( .A(A[457]), .B(n569), .CI(
        C[457]), .S(S[457]), .CO(C[458]) );
  FA_14194 \FA_INST_0[0].FA_INST_1[458].FA_  ( .A(A[458]), .B(n568), .CI(
        C[458]), .S(S[458]), .CO(C[459]) );
  FA_14193 \FA_INST_0[0].FA_INST_1[459].FA_  ( .A(A[459]), .B(n567), .CI(
        C[459]), .S(S[459]), .CO(C[460]) );
  FA_14192 \FA_INST_0[0].FA_INST_1[460].FA_  ( .A(A[460]), .B(n566), .CI(
        C[460]), .S(S[460]), .CO(C[461]) );
  FA_14191 \FA_INST_0[0].FA_INST_1[461].FA_  ( .A(A[461]), .B(n565), .CI(
        C[461]), .S(S[461]), .CO(C[462]) );
  FA_14190 \FA_INST_0[0].FA_INST_1[462].FA_  ( .A(A[462]), .B(n564), .CI(
        C[462]), .S(S[462]), .CO(C[463]) );
  FA_14189 \FA_INST_0[0].FA_INST_1[463].FA_  ( .A(A[463]), .B(n563), .CI(
        C[463]), .S(S[463]), .CO(C[464]) );
  FA_14188 \FA_INST_0[0].FA_INST_1[464].FA_  ( .A(A[464]), .B(n562), .CI(
        C[464]), .S(S[464]), .CO(C[465]) );
  FA_14187 \FA_INST_0[0].FA_INST_1[465].FA_  ( .A(A[465]), .B(n561), .CI(
        C[465]), .S(S[465]), .CO(C[466]) );
  FA_14186 \FA_INST_0[0].FA_INST_1[466].FA_  ( .A(A[466]), .B(n560), .CI(
        C[466]), .S(S[466]), .CO(C[467]) );
  FA_14185 \FA_INST_0[0].FA_INST_1[467].FA_  ( .A(A[467]), .B(n559), .CI(
        C[467]), .S(S[467]), .CO(C[468]) );
  FA_14184 \FA_INST_0[0].FA_INST_1[468].FA_  ( .A(A[468]), .B(n558), .CI(
        C[468]), .S(S[468]), .CO(C[469]) );
  FA_14183 \FA_INST_0[0].FA_INST_1[469].FA_  ( .A(A[469]), .B(n557), .CI(
        C[469]), .S(S[469]), .CO(C[470]) );
  FA_14182 \FA_INST_0[0].FA_INST_1[470].FA_  ( .A(A[470]), .B(n556), .CI(
        C[470]), .S(S[470]), .CO(C[471]) );
  FA_14181 \FA_INST_0[0].FA_INST_1[471].FA_  ( .A(A[471]), .B(n555), .CI(
        C[471]), .S(S[471]), .CO(C[472]) );
  FA_14180 \FA_INST_0[0].FA_INST_1[472].FA_  ( .A(A[472]), .B(n554), .CI(
        C[472]), .S(S[472]), .CO(C[473]) );
  FA_14179 \FA_INST_0[0].FA_INST_1[473].FA_  ( .A(A[473]), .B(n553), .CI(
        C[473]), .S(S[473]), .CO(C[474]) );
  FA_14178 \FA_INST_0[0].FA_INST_1[474].FA_  ( .A(A[474]), .B(n552), .CI(
        C[474]), .S(S[474]), .CO(C[475]) );
  FA_14177 \FA_INST_0[0].FA_INST_1[475].FA_  ( .A(A[475]), .B(n551), .CI(
        C[475]), .S(S[475]), .CO(C[476]) );
  FA_14176 \FA_INST_0[0].FA_INST_1[476].FA_  ( .A(A[476]), .B(n550), .CI(
        C[476]), .S(S[476]), .CO(C[477]) );
  FA_14175 \FA_INST_0[0].FA_INST_1[477].FA_  ( .A(A[477]), .B(n549), .CI(
        C[477]), .S(S[477]), .CO(C[478]) );
  FA_14174 \FA_INST_0[0].FA_INST_1[478].FA_  ( .A(A[478]), .B(n548), .CI(
        C[478]), .S(S[478]), .CO(C[479]) );
  FA_14173 \FA_INST_0[0].FA_INST_1[479].FA_  ( .A(A[479]), .B(n547), .CI(
        C[479]), .S(S[479]), .CO(C[480]) );
  FA_14172 \FA_INST_0[0].FA_INST_1[480].FA_  ( .A(A[480]), .B(n546), .CI(
        C[480]), .S(S[480]), .CO(C[481]) );
  FA_14171 \FA_INST_0[0].FA_INST_1[481].FA_  ( .A(A[481]), .B(n545), .CI(
        C[481]), .S(S[481]), .CO(C[482]) );
  FA_14170 \FA_INST_0[0].FA_INST_1[482].FA_  ( .A(A[482]), .B(n544), .CI(
        C[482]), .S(S[482]), .CO(C[483]) );
  FA_14169 \FA_INST_0[0].FA_INST_1[483].FA_  ( .A(A[483]), .B(n543), .CI(
        C[483]), .S(S[483]), .CO(C[484]) );
  FA_14168 \FA_INST_0[0].FA_INST_1[484].FA_  ( .A(A[484]), .B(n542), .CI(
        C[484]), .S(S[484]), .CO(C[485]) );
  FA_14167 \FA_INST_0[0].FA_INST_1[485].FA_  ( .A(A[485]), .B(n541), .CI(
        C[485]), .S(S[485]), .CO(C[486]) );
  FA_14166 \FA_INST_0[0].FA_INST_1[486].FA_  ( .A(A[486]), .B(n540), .CI(
        C[486]), .S(S[486]), .CO(C[487]) );
  FA_14165 \FA_INST_0[0].FA_INST_1[487].FA_  ( .A(A[487]), .B(n539), .CI(
        C[487]), .S(S[487]), .CO(C[488]) );
  FA_14164 \FA_INST_0[0].FA_INST_1[488].FA_  ( .A(A[488]), .B(n538), .CI(
        C[488]), .S(S[488]), .CO(C[489]) );
  FA_14163 \FA_INST_0[0].FA_INST_1[489].FA_  ( .A(A[489]), .B(n537), .CI(
        C[489]), .S(S[489]), .CO(C[490]) );
  FA_14162 \FA_INST_0[0].FA_INST_1[490].FA_  ( .A(A[490]), .B(n536), .CI(
        C[490]), .S(S[490]), .CO(C[491]) );
  FA_14161 \FA_INST_0[0].FA_INST_1[491].FA_  ( .A(A[491]), .B(n535), .CI(
        C[491]), .S(S[491]), .CO(C[492]) );
  FA_14160 \FA_INST_0[0].FA_INST_1[492].FA_  ( .A(A[492]), .B(n534), .CI(
        C[492]), .S(S[492]), .CO(C[493]) );
  FA_14159 \FA_INST_0[0].FA_INST_1[493].FA_  ( .A(A[493]), .B(n533), .CI(
        C[493]), .S(S[493]), .CO(C[494]) );
  FA_14158 \FA_INST_0[0].FA_INST_1[494].FA_  ( .A(A[494]), .B(n532), .CI(
        C[494]), .S(S[494]), .CO(C[495]) );
  FA_14157 \FA_INST_0[0].FA_INST_1[495].FA_  ( .A(A[495]), .B(n531), .CI(
        C[495]), .S(S[495]), .CO(C[496]) );
  FA_14156 \FA_INST_0[0].FA_INST_1[496].FA_  ( .A(A[496]), .B(n530), .CI(
        C[496]), .S(S[496]), .CO(C[497]) );
  FA_14155 \FA_INST_0[0].FA_INST_1[497].FA_  ( .A(A[497]), .B(n529), .CI(
        C[497]), .S(S[497]), .CO(C[498]) );
  FA_14154 \FA_INST_0[0].FA_INST_1[498].FA_  ( .A(A[498]), .B(n528), .CI(
        C[498]), .S(S[498]), .CO(C[499]) );
  FA_14153 \FA_INST_0[0].FA_INST_1[499].FA_  ( .A(A[499]), .B(n527), .CI(
        C[499]), .S(S[499]), .CO(C[500]) );
  FA_14152 \FA_INST_0[0].FA_INST_1[500].FA_  ( .A(A[500]), .B(n526), .CI(
        C[500]), .S(S[500]), .CO(C[501]) );
  FA_14151 \FA_INST_0[0].FA_INST_1[501].FA_  ( .A(A[501]), .B(n525), .CI(
        C[501]), .S(S[501]), .CO(C[502]) );
  FA_14150 \FA_INST_0[0].FA_INST_1[502].FA_  ( .A(A[502]), .B(n524), .CI(
        C[502]), .S(S[502]), .CO(C[503]) );
  FA_14149 \FA_INST_0[0].FA_INST_1[503].FA_  ( .A(A[503]), .B(n523), .CI(
        C[503]), .S(S[503]), .CO(C[504]) );
  FA_14148 \FA_INST_0[0].FA_INST_1[504].FA_  ( .A(A[504]), .B(n522), .CI(
        C[504]), .S(S[504]), .CO(C[505]) );
  FA_14147 \FA_INST_0[0].FA_INST_1[505].FA_  ( .A(A[505]), .B(n521), .CI(
        C[505]), .S(S[505]), .CO(C[506]) );
  FA_14146 \FA_INST_0[0].FA_INST_1[506].FA_  ( .A(A[506]), .B(n520), .CI(
        C[506]), .S(S[506]), .CO(C[507]) );
  FA_14145 \FA_INST_0[0].FA_INST_1[507].FA_  ( .A(A[507]), .B(n519), .CI(
        C[507]), .S(S[507]), .CO(C[508]) );
  FA_14144 \FA_INST_0[0].FA_INST_1[508].FA_  ( .A(A[508]), .B(n518), .CI(
        C[508]), .S(S[508]), .CO(C[509]) );
  FA_14143 \FA_INST_0[0].FA_INST_1[509].FA_  ( .A(A[509]), .B(n517), .CI(
        C[509]), .S(S[509]), .CO(C[510]) );
  FA_14142 \FA_INST_0[0].FA_INST_1[510].FA_  ( .A(A[510]), .B(n516), .CI(
        C[510]), .S(S[510]), .CO(C[511]) );
  FA_14141 \FA_INST_0[0].FA_INST_1[511].FA_  ( .A(A[511]), .B(n515), .CI(
        C[511]), .S(S[511]), .CO(C[512]) );
  FA_14140 \FA_INST_0[1].FA_INST_1[0].FA_  ( .A(A[512]), .B(n514), .CI(C[512]), 
        .S(S[512]), .CO(C[513]) );
  FA_14139 \FA_INST_0[1].FA_INST_1[1].FA_  ( .A(A[513]), .B(n513), .CI(C[513]), 
        .S(S[513]), .CO(C[514]) );
  FA_14138 \FA_INST_0[1].FA_INST_1[2].FA_  ( .A(A[514]), .B(n512), .CI(C[514]), 
        .S(S[514]), .CO(C[515]) );
  FA_14137 \FA_INST_0[1].FA_INST_1[3].FA_  ( .A(A[515]), .B(n511), .CI(C[515]), 
        .S(S[515]), .CO(C[516]) );
  FA_14136 \FA_INST_0[1].FA_INST_1[4].FA_  ( .A(A[516]), .B(n510), .CI(C[516]), 
        .S(S[516]), .CO(C[517]) );
  FA_14135 \FA_INST_0[1].FA_INST_1[5].FA_  ( .A(A[517]), .B(n509), .CI(C[517]), 
        .S(S[517]), .CO(C[518]) );
  FA_14134 \FA_INST_0[1].FA_INST_1[6].FA_  ( .A(A[518]), .B(n508), .CI(C[518]), 
        .S(S[518]), .CO(C[519]) );
  FA_14133 \FA_INST_0[1].FA_INST_1[7].FA_  ( .A(A[519]), .B(n507), .CI(C[519]), 
        .S(S[519]), .CO(C[520]) );
  FA_14132 \FA_INST_0[1].FA_INST_1[8].FA_  ( .A(A[520]), .B(n506), .CI(C[520]), 
        .S(S[520]), .CO(C[521]) );
  FA_14131 \FA_INST_0[1].FA_INST_1[9].FA_  ( .A(A[521]), .B(n505), .CI(C[521]), 
        .S(S[521]), .CO(C[522]) );
  FA_14130 \FA_INST_0[1].FA_INST_1[10].FA_  ( .A(A[522]), .B(n504), .CI(C[522]), .S(S[522]), .CO(C[523]) );
  FA_14129 \FA_INST_0[1].FA_INST_1[11].FA_  ( .A(A[523]), .B(n503), .CI(C[523]), .S(S[523]), .CO(C[524]) );
  FA_14128 \FA_INST_0[1].FA_INST_1[12].FA_  ( .A(A[524]), .B(n502), .CI(C[524]), .S(S[524]), .CO(C[525]) );
  FA_14127 \FA_INST_0[1].FA_INST_1[13].FA_  ( .A(A[525]), .B(n501), .CI(C[525]), .S(S[525]), .CO(C[526]) );
  FA_14126 \FA_INST_0[1].FA_INST_1[14].FA_  ( .A(A[526]), .B(n500), .CI(C[526]), .S(S[526]), .CO(C[527]) );
  FA_14125 \FA_INST_0[1].FA_INST_1[15].FA_  ( .A(A[527]), .B(n499), .CI(C[527]), .S(S[527]), .CO(C[528]) );
  FA_14124 \FA_INST_0[1].FA_INST_1[16].FA_  ( .A(A[528]), .B(n498), .CI(C[528]), .S(S[528]), .CO(C[529]) );
  FA_14123 \FA_INST_0[1].FA_INST_1[17].FA_  ( .A(A[529]), .B(n497), .CI(C[529]), .S(S[529]), .CO(C[530]) );
  FA_14122 \FA_INST_0[1].FA_INST_1[18].FA_  ( .A(A[530]), .B(n496), .CI(C[530]), .S(S[530]), .CO(C[531]) );
  FA_14121 \FA_INST_0[1].FA_INST_1[19].FA_  ( .A(A[531]), .B(n495), .CI(C[531]), .S(S[531]), .CO(C[532]) );
  FA_14120 \FA_INST_0[1].FA_INST_1[20].FA_  ( .A(A[532]), .B(n494), .CI(C[532]), .S(S[532]), .CO(C[533]) );
  FA_14119 \FA_INST_0[1].FA_INST_1[21].FA_  ( .A(A[533]), .B(n493), .CI(C[533]), .S(S[533]), .CO(C[534]) );
  FA_14118 \FA_INST_0[1].FA_INST_1[22].FA_  ( .A(A[534]), .B(n492), .CI(C[534]), .S(S[534]), .CO(C[535]) );
  FA_14117 \FA_INST_0[1].FA_INST_1[23].FA_  ( .A(A[535]), .B(n491), .CI(C[535]), .S(S[535]), .CO(C[536]) );
  FA_14116 \FA_INST_0[1].FA_INST_1[24].FA_  ( .A(A[536]), .B(n490), .CI(C[536]), .S(S[536]), .CO(C[537]) );
  FA_14115 \FA_INST_0[1].FA_INST_1[25].FA_  ( .A(A[537]), .B(n489), .CI(C[537]), .S(S[537]), .CO(C[538]) );
  FA_14114 \FA_INST_0[1].FA_INST_1[26].FA_  ( .A(A[538]), .B(n488), .CI(C[538]), .S(S[538]), .CO(C[539]) );
  FA_14113 \FA_INST_0[1].FA_INST_1[27].FA_  ( .A(A[539]), .B(n487), .CI(C[539]), .S(S[539]), .CO(C[540]) );
  FA_14112 \FA_INST_0[1].FA_INST_1[28].FA_  ( .A(A[540]), .B(n486), .CI(C[540]), .S(S[540]), .CO(C[541]) );
  FA_14111 \FA_INST_0[1].FA_INST_1[29].FA_  ( .A(A[541]), .B(n485), .CI(C[541]), .S(S[541]), .CO(C[542]) );
  FA_14110 \FA_INST_0[1].FA_INST_1[30].FA_  ( .A(A[542]), .B(n484), .CI(C[542]), .S(S[542]), .CO(C[543]) );
  FA_14109 \FA_INST_0[1].FA_INST_1[31].FA_  ( .A(A[543]), .B(n483), .CI(C[543]), .S(S[543]), .CO(C[544]) );
  FA_14108 \FA_INST_0[1].FA_INST_1[32].FA_  ( .A(A[544]), .B(n482), .CI(C[544]), .S(S[544]), .CO(C[545]) );
  FA_14107 \FA_INST_0[1].FA_INST_1[33].FA_  ( .A(A[545]), .B(n481), .CI(C[545]), .S(S[545]), .CO(C[546]) );
  FA_14106 \FA_INST_0[1].FA_INST_1[34].FA_  ( .A(A[546]), .B(n480), .CI(C[546]), .S(S[546]), .CO(C[547]) );
  FA_14105 \FA_INST_0[1].FA_INST_1[35].FA_  ( .A(A[547]), .B(n479), .CI(C[547]), .S(S[547]), .CO(C[548]) );
  FA_14104 \FA_INST_0[1].FA_INST_1[36].FA_  ( .A(A[548]), .B(n478), .CI(C[548]), .S(S[548]), .CO(C[549]) );
  FA_14103 \FA_INST_0[1].FA_INST_1[37].FA_  ( .A(A[549]), .B(n477), .CI(C[549]), .S(S[549]), .CO(C[550]) );
  FA_14102 \FA_INST_0[1].FA_INST_1[38].FA_  ( .A(A[550]), .B(n476), .CI(C[550]), .S(S[550]), .CO(C[551]) );
  FA_14101 \FA_INST_0[1].FA_INST_1[39].FA_  ( .A(A[551]), .B(n475), .CI(C[551]), .S(S[551]), .CO(C[552]) );
  FA_14100 \FA_INST_0[1].FA_INST_1[40].FA_  ( .A(A[552]), .B(n474), .CI(C[552]), .S(S[552]), .CO(C[553]) );
  FA_14099 \FA_INST_0[1].FA_INST_1[41].FA_  ( .A(A[553]), .B(n473), .CI(C[553]), .S(S[553]), .CO(C[554]) );
  FA_14098 \FA_INST_0[1].FA_INST_1[42].FA_  ( .A(A[554]), .B(n472), .CI(C[554]), .S(S[554]), .CO(C[555]) );
  FA_14097 \FA_INST_0[1].FA_INST_1[43].FA_  ( .A(A[555]), .B(n471), .CI(C[555]), .S(S[555]), .CO(C[556]) );
  FA_14096 \FA_INST_0[1].FA_INST_1[44].FA_  ( .A(A[556]), .B(n470), .CI(C[556]), .S(S[556]), .CO(C[557]) );
  FA_14095 \FA_INST_0[1].FA_INST_1[45].FA_  ( .A(A[557]), .B(n469), .CI(C[557]), .S(S[557]), .CO(C[558]) );
  FA_14094 \FA_INST_0[1].FA_INST_1[46].FA_  ( .A(A[558]), .B(n468), .CI(C[558]), .S(S[558]), .CO(C[559]) );
  FA_14093 \FA_INST_0[1].FA_INST_1[47].FA_  ( .A(A[559]), .B(n467), .CI(C[559]), .S(S[559]), .CO(C[560]) );
  FA_14092 \FA_INST_0[1].FA_INST_1[48].FA_  ( .A(A[560]), .B(n466), .CI(C[560]), .S(S[560]), .CO(C[561]) );
  FA_14091 \FA_INST_0[1].FA_INST_1[49].FA_  ( .A(A[561]), .B(n465), .CI(C[561]), .S(S[561]), .CO(C[562]) );
  FA_14090 \FA_INST_0[1].FA_INST_1[50].FA_  ( .A(A[562]), .B(n464), .CI(C[562]), .S(S[562]), .CO(C[563]) );
  FA_14089 \FA_INST_0[1].FA_INST_1[51].FA_  ( .A(A[563]), .B(n463), .CI(C[563]), .S(S[563]), .CO(C[564]) );
  FA_14088 \FA_INST_0[1].FA_INST_1[52].FA_  ( .A(A[564]), .B(n462), .CI(C[564]), .S(S[564]), .CO(C[565]) );
  FA_14087 \FA_INST_0[1].FA_INST_1[53].FA_  ( .A(A[565]), .B(n461), .CI(C[565]), .S(S[565]), .CO(C[566]) );
  FA_14086 \FA_INST_0[1].FA_INST_1[54].FA_  ( .A(A[566]), .B(n460), .CI(C[566]), .S(S[566]), .CO(C[567]) );
  FA_14085 \FA_INST_0[1].FA_INST_1[55].FA_  ( .A(A[567]), .B(n459), .CI(C[567]), .S(S[567]), .CO(C[568]) );
  FA_14084 \FA_INST_0[1].FA_INST_1[56].FA_  ( .A(A[568]), .B(n458), .CI(C[568]), .S(S[568]), .CO(C[569]) );
  FA_14083 \FA_INST_0[1].FA_INST_1[57].FA_  ( .A(A[569]), .B(n457), .CI(C[569]), .S(S[569]), .CO(C[570]) );
  FA_14082 \FA_INST_0[1].FA_INST_1[58].FA_  ( .A(A[570]), .B(n456), .CI(C[570]), .S(S[570]), .CO(C[571]) );
  FA_14081 \FA_INST_0[1].FA_INST_1[59].FA_  ( .A(A[571]), .B(n455), .CI(C[571]), .S(S[571]), .CO(C[572]) );
  FA_14080 \FA_INST_0[1].FA_INST_1[60].FA_  ( .A(A[572]), .B(n454), .CI(C[572]), .S(S[572]), .CO(C[573]) );
  FA_14079 \FA_INST_0[1].FA_INST_1[61].FA_  ( .A(A[573]), .B(n453), .CI(C[573]), .S(S[573]), .CO(C[574]) );
  FA_14078 \FA_INST_0[1].FA_INST_1[62].FA_  ( .A(A[574]), .B(n452), .CI(C[574]), .S(S[574]), .CO(C[575]) );
  FA_14077 \FA_INST_0[1].FA_INST_1[63].FA_  ( .A(A[575]), .B(n451), .CI(C[575]), .S(S[575]), .CO(C[576]) );
  FA_14076 \FA_INST_0[1].FA_INST_1[64].FA_  ( .A(A[576]), .B(n450), .CI(C[576]), .S(S[576]), .CO(C[577]) );
  FA_14075 \FA_INST_0[1].FA_INST_1[65].FA_  ( .A(A[577]), .B(n449), .CI(C[577]), .S(S[577]), .CO(C[578]) );
  FA_14074 \FA_INST_0[1].FA_INST_1[66].FA_  ( .A(A[578]), .B(n448), .CI(C[578]), .S(S[578]), .CO(C[579]) );
  FA_14073 \FA_INST_0[1].FA_INST_1[67].FA_  ( .A(A[579]), .B(n447), .CI(C[579]), .S(S[579]), .CO(C[580]) );
  FA_14072 \FA_INST_0[1].FA_INST_1[68].FA_  ( .A(A[580]), .B(n446), .CI(C[580]), .S(S[580]), .CO(C[581]) );
  FA_14071 \FA_INST_0[1].FA_INST_1[69].FA_  ( .A(A[581]), .B(n445), .CI(C[581]), .S(S[581]), .CO(C[582]) );
  FA_14070 \FA_INST_0[1].FA_INST_1[70].FA_  ( .A(A[582]), .B(n444), .CI(C[582]), .S(S[582]), .CO(C[583]) );
  FA_14069 \FA_INST_0[1].FA_INST_1[71].FA_  ( .A(A[583]), .B(n443), .CI(C[583]), .S(S[583]), .CO(C[584]) );
  FA_14068 \FA_INST_0[1].FA_INST_1[72].FA_  ( .A(A[584]), .B(n442), .CI(C[584]), .S(S[584]), .CO(C[585]) );
  FA_14067 \FA_INST_0[1].FA_INST_1[73].FA_  ( .A(A[585]), .B(n441), .CI(C[585]), .S(S[585]), .CO(C[586]) );
  FA_14066 \FA_INST_0[1].FA_INST_1[74].FA_  ( .A(A[586]), .B(n440), .CI(C[586]), .S(S[586]), .CO(C[587]) );
  FA_14065 \FA_INST_0[1].FA_INST_1[75].FA_  ( .A(A[587]), .B(n439), .CI(C[587]), .S(S[587]), .CO(C[588]) );
  FA_14064 \FA_INST_0[1].FA_INST_1[76].FA_  ( .A(A[588]), .B(n438), .CI(C[588]), .S(S[588]), .CO(C[589]) );
  FA_14063 \FA_INST_0[1].FA_INST_1[77].FA_  ( .A(A[589]), .B(n437), .CI(C[589]), .S(S[589]), .CO(C[590]) );
  FA_14062 \FA_INST_0[1].FA_INST_1[78].FA_  ( .A(A[590]), .B(n436), .CI(C[590]), .S(S[590]), .CO(C[591]) );
  FA_14061 \FA_INST_0[1].FA_INST_1[79].FA_  ( .A(A[591]), .B(n435), .CI(C[591]), .S(S[591]), .CO(C[592]) );
  FA_14060 \FA_INST_0[1].FA_INST_1[80].FA_  ( .A(A[592]), .B(n434), .CI(C[592]), .S(S[592]), .CO(C[593]) );
  FA_14059 \FA_INST_0[1].FA_INST_1[81].FA_  ( .A(A[593]), .B(n433), .CI(C[593]), .S(S[593]), .CO(C[594]) );
  FA_14058 \FA_INST_0[1].FA_INST_1[82].FA_  ( .A(A[594]), .B(n432), .CI(C[594]), .S(S[594]), .CO(C[595]) );
  FA_14057 \FA_INST_0[1].FA_INST_1[83].FA_  ( .A(A[595]), .B(n431), .CI(C[595]), .S(S[595]), .CO(C[596]) );
  FA_14056 \FA_INST_0[1].FA_INST_1[84].FA_  ( .A(A[596]), .B(n430), .CI(C[596]), .S(S[596]), .CO(C[597]) );
  FA_14055 \FA_INST_0[1].FA_INST_1[85].FA_  ( .A(A[597]), .B(n429), .CI(C[597]), .S(S[597]), .CO(C[598]) );
  FA_14054 \FA_INST_0[1].FA_INST_1[86].FA_  ( .A(A[598]), .B(n428), .CI(C[598]), .S(S[598]), .CO(C[599]) );
  FA_14053 \FA_INST_0[1].FA_INST_1[87].FA_  ( .A(A[599]), .B(n427), .CI(C[599]), .S(S[599]), .CO(C[600]) );
  FA_14052 \FA_INST_0[1].FA_INST_1[88].FA_  ( .A(A[600]), .B(n426), .CI(C[600]), .S(S[600]), .CO(C[601]) );
  FA_14051 \FA_INST_0[1].FA_INST_1[89].FA_  ( .A(A[601]), .B(n425), .CI(C[601]), .S(S[601]), .CO(C[602]) );
  FA_14050 \FA_INST_0[1].FA_INST_1[90].FA_  ( .A(A[602]), .B(n424), .CI(C[602]), .S(S[602]), .CO(C[603]) );
  FA_14049 \FA_INST_0[1].FA_INST_1[91].FA_  ( .A(A[603]), .B(n423), .CI(C[603]), .S(S[603]), .CO(C[604]) );
  FA_14048 \FA_INST_0[1].FA_INST_1[92].FA_  ( .A(A[604]), .B(n422), .CI(C[604]), .S(S[604]), .CO(C[605]) );
  FA_14047 \FA_INST_0[1].FA_INST_1[93].FA_  ( .A(A[605]), .B(n421), .CI(C[605]), .S(S[605]), .CO(C[606]) );
  FA_14046 \FA_INST_0[1].FA_INST_1[94].FA_  ( .A(A[606]), .B(n420), .CI(C[606]), .S(S[606]), .CO(C[607]) );
  FA_14045 \FA_INST_0[1].FA_INST_1[95].FA_  ( .A(A[607]), .B(n419), .CI(C[607]), .S(S[607]), .CO(C[608]) );
  FA_14044 \FA_INST_0[1].FA_INST_1[96].FA_  ( .A(A[608]), .B(n418), .CI(C[608]), .S(S[608]), .CO(C[609]) );
  FA_14043 \FA_INST_0[1].FA_INST_1[97].FA_  ( .A(A[609]), .B(n417), .CI(C[609]), .S(S[609]), .CO(C[610]) );
  FA_14042 \FA_INST_0[1].FA_INST_1[98].FA_  ( .A(A[610]), .B(n416), .CI(C[610]), .S(S[610]), .CO(C[611]) );
  FA_14041 \FA_INST_0[1].FA_INST_1[99].FA_  ( .A(A[611]), .B(n415), .CI(C[611]), .S(S[611]), .CO(C[612]) );
  FA_14040 \FA_INST_0[1].FA_INST_1[100].FA_  ( .A(A[612]), .B(n414), .CI(
        C[612]), .S(S[612]), .CO(C[613]) );
  FA_14039 \FA_INST_0[1].FA_INST_1[101].FA_  ( .A(A[613]), .B(n413), .CI(
        C[613]), .S(S[613]), .CO(C[614]) );
  FA_14038 \FA_INST_0[1].FA_INST_1[102].FA_  ( .A(A[614]), .B(n412), .CI(
        C[614]), .S(S[614]), .CO(C[615]) );
  FA_14037 \FA_INST_0[1].FA_INST_1[103].FA_  ( .A(A[615]), .B(n411), .CI(
        C[615]), .S(S[615]), .CO(C[616]) );
  FA_14036 \FA_INST_0[1].FA_INST_1[104].FA_  ( .A(A[616]), .B(n410), .CI(
        C[616]), .S(S[616]), .CO(C[617]) );
  FA_14035 \FA_INST_0[1].FA_INST_1[105].FA_  ( .A(A[617]), .B(n409), .CI(
        C[617]), .S(S[617]), .CO(C[618]) );
  FA_14034 \FA_INST_0[1].FA_INST_1[106].FA_  ( .A(A[618]), .B(n408), .CI(
        C[618]), .S(S[618]), .CO(C[619]) );
  FA_14033 \FA_INST_0[1].FA_INST_1[107].FA_  ( .A(A[619]), .B(n407), .CI(
        C[619]), .S(S[619]), .CO(C[620]) );
  FA_14032 \FA_INST_0[1].FA_INST_1[108].FA_  ( .A(A[620]), .B(n406), .CI(
        C[620]), .S(S[620]), .CO(C[621]) );
  FA_14031 \FA_INST_0[1].FA_INST_1[109].FA_  ( .A(A[621]), .B(n405), .CI(
        C[621]), .S(S[621]), .CO(C[622]) );
  FA_14030 \FA_INST_0[1].FA_INST_1[110].FA_  ( .A(A[622]), .B(n404), .CI(
        C[622]), .S(S[622]), .CO(C[623]) );
  FA_14029 \FA_INST_0[1].FA_INST_1[111].FA_  ( .A(A[623]), .B(n403), .CI(
        C[623]), .S(S[623]), .CO(C[624]) );
  FA_14028 \FA_INST_0[1].FA_INST_1[112].FA_  ( .A(A[624]), .B(n402), .CI(
        C[624]), .S(S[624]), .CO(C[625]) );
  FA_14027 \FA_INST_0[1].FA_INST_1[113].FA_  ( .A(A[625]), .B(n401), .CI(
        C[625]), .S(S[625]), .CO(C[626]) );
  FA_14026 \FA_INST_0[1].FA_INST_1[114].FA_  ( .A(A[626]), .B(n400), .CI(
        C[626]), .S(S[626]), .CO(C[627]) );
  FA_14025 \FA_INST_0[1].FA_INST_1[115].FA_  ( .A(A[627]), .B(n399), .CI(
        C[627]), .S(S[627]), .CO(C[628]) );
  FA_14024 \FA_INST_0[1].FA_INST_1[116].FA_  ( .A(A[628]), .B(n398), .CI(
        C[628]), .S(S[628]), .CO(C[629]) );
  FA_14023 \FA_INST_0[1].FA_INST_1[117].FA_  ( .A(A[629]), .B(n397), .CI(
        C[629]), .S(S[629]), .CO(C[630]) );
  FA_14022 \FA_INST_0[1].FA_INST_1[118].FA_  ( .A(A[630]), .B(n396), .CI(
        C[630]), .S(S[630]), .CO(C[631]) );
  FA_14021 \FA_INST_0[1].FA_INST_1[119].FA_  ( .A(A[631]), .B(n395), .CI(
        C[631]), .S(S[631]), .CO(C[632]) );
  FA_14020 \FA_INST_0[1].FA_INST_1[120].FA_  ( .A(A[632]), .B(n394), .CI(
        C[632]), .S(S[632]), .CO(C[633]) );
  FA_14019 \FA_INST_0[1].FA_INST_1[121].FA_  ( .A(A[633]), .B(n393), .CI(
        C[633]), .S(S[633]), .CO(C[634]) );
  FA_14018 \FA_INST_0[1].FA_INST_1[122].FA_  ( .A(A[634]), .B(n392), .CI(
        C[634]), .S(S[634]), .CO(C[635]) );
  FA_14017 \FA_INST_0[1].FA_INST_1[123].FA_  ( .A(A[635]), .B(n391), .CI(
        C[635]), .S(S[635]), .CO(C[636]) );
  FA_14016 \FA_INST_0[1].FA_INST_1[124].FA_  ( .A(A[636]), .B(n390), .CI(
        C[636]), .S(S[636]), .CO(C[637]) );
  FA_14015 \FA_INST_0[1].FA_INST_1[125].FA_  ( .A(A[637]), .B(n389), .CI(
        C[637]), .S(S[637]), .CO(C[638]) );
  FA_14014 \FA_INST_0[1].FA_INST_1[126].FA_  ( .A(A[638]), .B(n388), .CI(
        C[638]), .S(S[638]), .CO(C[639]) );
  FA_14013 \FA_INST_0[1].FA_INST_1[127].FA_  ( .A(A[639]), .B(n387), .CI(
        C[639]), .S(S[639]), .CO(C[640]) );
  FA_14012 \FA_INST_0[1].FA_INST_1[128].FA_  ( .A(A[640]), .B(n386), .CI(
        C[640]), .S(S[640]), .CO(C[641]) );
  FA_14011 \FA_INST_0[1].FA_INST_1[129].FA_  ( .A(A[641]), .B(n385), .CI(
        C[641]), .S(S[641]), .CO(C[642]) );
  FA_14010 \FA_INST_0[1].FA_INST_1[130].FA_  ( .A(A[642]), .B(n384), .CI(
        C[642]), .S(S[642]), .CO(C[643]) );
  FA_14009 \FA_INST_0[1].FA_INST_1[131].FA_  ( .A(A[643]), .B(n383), .CI(
        C[643]), .S(S[643]), .CO(C[644]) );
  FA_14008 \FA_INST_0[1].FA_INST_1[132].FA_  ( .A(A[644]), .B(n382), .CI(
        C[644]), .S(S[644]), .CO(C[645]) );
  FA_14007 \FA_INST_0[1].FA_INST_1[133].FA_  ( .A(A[645]), .B(n381), .CI(
        C[645]), .S(S[645]), .CO(C[646]) );
  FA_14006 \FA_INST_0[1].FA_INST_1[134].FA_  ( .A(A[646]), .B(n380), .CI(
        C[646]), .S(S[646]), .CO(C[647]) );
  FA_14005 \FA_INST_0[1].FA_INST_1[135].FA_  ( .A(A[647]), .B(n379), .CI(
        C[647]), .S(S[647]), .CO(C[648]) );
  FA_14004 \FA_INST_0[1].FA_INST_1[136].FA_  ( .A(A[648]), .B(n378), .CI(
        C[648]), .S(S[648]), .CO(C[649]) );
  FA_14003 \FA_INST_0[1].FA_INST_1[137].FA_  ( .A(A[649]), .B(n377), .CI(
        C[649]), .S(S[649]), .CO(C[650]) );
  FA_14002 \FA_INST_0[1].FA_INST_1[138].FA_  ( .A(A[650]), .B(n376), .CI(
        C[650]), .S(S[650]), .CO(C[651]) );
  FA_14001 \FA_INST_0[1].FA_INST_1[139].FA_  ( .A(A[651]), .B(n375), .CI(
        C[651]), .S(S[651]), .CO(C[652]) );
  FA_14000 \FA_INST_0[1].FA_INST_1[140].FA_  ( .A(A[652]), .B(n374), .CI(
        C[652]), .S(S[652]), .CO(C[653]) );
  FA_13999 \FA_INST_0[1].FA_INST_1[141].FA_  ( .A(A[653]), .B(n373), .CI(
        C[653]), .S(S[653]), .CO(C[654]) );
  FA_13998 \FA_INST_0[1].FA_INST_1[142].FA_  ( .A(A[654]), .B(n372), .CI(
        C[654]), .S(S[654]), .CO(C[655]) );
  FA_13997 \FA_INST_0[1].FA_INST_1[143].FA_  ( .A(A[655]), .B(n371), .CI(
        C[655]), .S(S[655]), .CO(C[656]) );
  FA_13996 \FA_INST_0[1].FA_INST_1[144].FA_  ( .A(A[656]), .B(n370), .CI(
        C[656]), .S(S[656]), .CO(C[657]) );
  FA_13995 \FA_INST_0[1].FA_INST_1[145].FA_  ( .A(A[657]), .B(n369), .CI(
        C[657]), .S(S[657]), .CO(C[658]) );
  FA_13994 \FA_INST_0[1].FA_INST_1[146].FA_  ( .A(A[658]), .B(n368), .CI(
        C[658]), .S(S[658]), .CO(C[659]) );
  FA_13993 \FA_INST_0[1].FA_INST_1[147].FA_  ( .A(A[659]), .B(n367), .CI(
        C[659]), .S(S[659]), .CO(C[660]) );
  FA_13992 \FA_INST_0[1].FA_INST_1[148].FA_  ( .A(A[660]), .B(n366), .CI(
        C[660]), .S(S[660]), .CO(C[661]) );
  FA_13991 \FA_INST_0[1].FA_INST_1[149].FA_  ( .A(A[661]), .B(n365), .CI(
        C[661]), .S(S[661]), .CO(C[662]) );
  FA_13990 \FA_INST_0[1].FA_INST_1[150].FA_  ( .A(A[662]), .B(n364), .CI(
        C[662]), .S(S[662]), .CO(C[663]) );
  FA_13989 \FA_INST_0[1].FA_INST_1[151].FA_  ( .A(A[663]), .B(n363), .CI(
        C[663]), .S(S[663]), .CO(C[664]) );
  FA_13988 \FA_INST_0[1].FA_INST_1[152].FA_  ( .A(A[664]), .B(n362), .CI(
        C[664]), .S(S[664]), .CO(C[665]) );
  FA_13987 \FA_INST_0[1].FA_INST_1[153].FA_  ( .A(A[665]), .B(n361), .CI(
        C[665]), .S(S[665]), .CO(C[666]) );
  FA_13986 \FA_INST_0[1].FA_INST_1[154].FA_  ( .A(A[666]), .B(n360), .CI(
        C[666]), .S(S[666]), .CO(C[667]) );
  FA_13985 \FA_INST_0[1].FA_INST_1[155].FA_  ( .A(A[667]), .B(n359), .CI(
        C[667]), .S(S[667]), .CO(C[668]) );
  FA_13984 \FA_INST_0[1].FA_INST_1[156].FA_  ( .A(A[668]), .B(n358), .CI(
        C[668]), .S(S[668]), .CO(C[669]) );
  FA_13983 \FA_INST_0[1].FA_INST_1[157].FA_  ( .A(A[669]), .B(n357), .CI(
        C[669]), .S(S[669]), .CO(C[670]) );
  FA_13982 \FA_INST_0[1].FA_INST_1[158].FA_  ( .A(A[670]), .B(n356), .CI(
        C[670]), .S(S[670]), .CO(C[671]) );
  FA_13981 \FA_INST_0[1].FA_INST_1[159].FA_  ( .A(A[671]), .B(n355), .CI(
        C[671]), .S(S[671]), .CO(C[672]) );
  FA_13980 \FA_INST_0[1].FA_INST_1[160].FA_  ( .A(A[672]), .B(n354), .CI(
        C[672]), .S(S[672]), .CO(C[673]) );
  FA_13979 \FA_INST_0[1].FA_INST_1[161].FA_  ( .A(A[673]), .B(n353), .CI(
        C[673]), .S(S[673]), .CO(C[674]) );
  FA_13978 \FA_INST_0[1].FA_INST_1[162].FA_  ( .A(A[674]), .B(n352), .CI(
        C[674]), .S(S[674]), .CO(C[675]) );
  FA_13977 \FA_INST_0[1].FA_INST_1[163].FA_  ( .A(A[675]), .B(n351), .CI(
        C[675]), .S(S[675]), .CO(C[676]) );
  FA_13976 \FA_INST_0[1].FA_INST_1[164].FA_  ( .A(A[676]), .B(n350), .CI(
        C[676]), .S(S[676]), .CO(C[677]) );
  FA_13975 \FA_INST_0[1].FA_INST_1[165].FA_  ( .A(A[677]), .B(n349), .CI(
        C[677]), .S(S[677]), .CO(C[678]) );
  FA_13974 \FA_INST_0[1].FA_INST_1[166].FA_  ( .A(A[678]), .B(n348), .CI(
        C[678]), .S(S[678]), .CO(C[679]) );
  FA_13973 \FA_INST_0[1].FA_INST_1[167].FA_  ( .A(A[679]), .B(n347), .CI(
        C[679]), .S(S[679]), .CO(C[680]) );
  FA_13972 \FA_INST_0[1].FA_INST_1[168].FA_  ( .A(A[680]), .B(n346), .CI(
        C[680]), .S(S[680]), .CO(C[681]) );
  FA_13971 \FA_INST_0[1].FA_INST_1[169].FA_  ( .A(A[681]), .B(n345), .CI(
        C[681]), .S(S[681]), .CO(C[682]) );
  FA_13970 \FA_INST_0[1].FA_INST_1[170].FA_  ( .A(A[682]), .B(n344), .CI(
        C[682]), .S(S[682]), .CO(C[683]) );
  FA_13969 \FA_INST_0[1].FA_INST_1[171].FA_  ( .A(A[683]), .B(n343), .CI(
        C[683]), .S(S[683]), .CO(C[684]) );
  FA_13968 \FA_INST_0[1].FA_INST_1[172].FA_  ( .A(A[684]), .B(n342), .CI(
        C[684]), .S(S[684]), .CO(C[685]) );
  FA_13967 \FA_INST_0[1].FA_INST_1[173].FA_  ( .A(A[685]), .B(n341), .CI(
        C[685]), .S(S[685]), .CO(C[686]) );
  FA_13966 \FA_INST_0[1].FA_INST_1[174].FA_  ( .A(A[686]), .B(n340), .CI(
        C[686]), .S(S[686]), .CO(C[687]) );
  FA_13965 \FA_INST_0[1].FA_INST_1[175].FA_  ( .A(A[687]), .B(n339), .CI(
        C[687]), .S(S[687]), .CO(C[688]) );
  FA_13964 \FA_INST_0[1].FA_INST_1[176].FA_  ( .A(A[688]), .B(n338), .CI(
        C[688]), .S(S[688]), .CO(C[689]) );
  FA_13963 \FA_INST_0[1].FA_INST_1[177].FA_  ( .A(A[689]), .B(n337), .CI(
        C[689]), .S(S[689]), .CO(C[690]) );
  FA_13962 \FA_INST_0[1].FA_INST_1[178].FA_  ( .A(A[690]), .B(n336), .CI(
        C[690]), .S(S[690]), .CO(C[691]) );
  FA_13961 \FA_INST_0[1].FA_INST_1[179].FA_  ( .A(A[691]), .B(n335), .CI(
        C[691]), .S(S[691]), .CO(C[692]) );
  FA_13960 \FA_INST_0[1].FA_INST_1[180].FA_  ( .A(A[692]), .B(n334), .CI(
        C[692]), .S(S[692]), .CO(C[693]) );
  FA_13959 \FA_INST_0[1].FA_INST_1[181].FA_  ( .A(A[693]), .B(n333), .CI(
        C[693]), .S(S[693]), .CO(C[694]) );
  FA_13958 \FA_INST_0[1].FA_INST_1[182].FA_  ( .A(A[694]), .B(n332), .CI(
        C[694]), .S(S[694]), .CO(C[695]) );
  FA_13957 \FA_INST_0[1].FA_INST_1[183].FA_  ( .A(A[695]), .B(n331), .CI(
        C[695]), .S(S[695]), .CO(C[696]) );
  FA_13956 \FA_INST_0[1].FA_INST_1[184].FA_  ( .A(A[696]), .B(n330), .CI(
        C[696]), .S(S[696]), .CO(C[697]) );
  FA_13955 \FA_INST_0[1].FA_INST_1[185].FA_  ( .A(A[697]), .B(n329), .CI(
        C[697]), .S(S[697]), .CO(C[698]) );
  FA_13954 \FA_INST_0[1].FA_INST_1[186].FA_  ( .A(A[698]), .B(n328), .CI(
        C[698]), .S(S[698]), .CO(C[699]) );
  FA_13953 \FA_INST_0[1].FA_INST_1[187].FA_  ( .A(A[699]), .B(n327), .CI(
        C[699]), .S(S[699]), .CO(C[700]) );
  FA_13952 \FA_INST_0[1].FA_INST_1[188].FA_  ( .A(A[700]), .B(n326), .CI(
        C[700]), .S(S[700]), .CO(C[701]) );
  FA_13951 \FA_INST_0[1].FA_INST_1[189].FA_  ( .A(A[701]), .B(n325), .CI(
        C[701]), .S(S[701]), .CO(C[702]) );
  FA_13950 \FA_INST_0[1].FA_INST_1[190].FA_  ( .A(A[702]), .B(n324), .CI(
        C[702]), .S(S[702]), .CO(C[703]) );
  FA_13949 \FA_INST_0[1].FA_INST_1[191].FA_  ( .A(A[703]), .B(n323), .CI(
        C[703]), .S(S[703]), .CO(C[704]) );
  FA_13948 \FA_INST_0[1].FA_INST_1[192].FA_  ( .A(A[704]), .B(n322), .CI(
        C[704]), .S(S[704]), .CO(C[705]) );
  FA_13947 \FA_INST_0[1].FA_INST_1[193].FA_  ( .A(A[705]), .B(n321), .CI(
        C[705]), .S(S[705]), .CO(C[706]) );
  FA_13946 \FA_INST_0[1].FA_INST_1[194].FA_  ( .A(A[706]), .B(n320), .CI(
        C[706]), .S(S[706]), .CO(C[707]) );
  FA_13945 \FA_INST_0[1].FA_INST_1[195].FA_  ( .A(A[707]), .B(n319), .CI(
        C[707]), .S(S[707]), .CO(C[708]) );
  FA_13944 \FA_INST_0[1].FA_INST_1[196].FA_  ( .A(A[708]), .B(n318), .CI(
        C[708]), .S(S[708]), .CO(C[709]) );
  FA_13943 \FA_INST_0[1].FA_INST_1[197].FA_  ( .A(A[709]), .B(n317), .CI(
        C[709]), .S(S[709]), .CO(C[710]) );
  FA_13942 \FA_INST_0[1].FA_INST_1[198].FA_  ( .A(A[710]), .B(n316), .CI(
        C[710]), .S(S[710]), .CO(C[711]) );
  FA_13941 \FA_INST_0[1].FA_INST_1[199].FA_  ( .A(A[711]), .B(n315), .CI(
        C[711]), .S(S[711]), .CO(C[712]) );
  FA_13940 \FA_INST_0[1].FA_INST_1[200].FA_  ( .A(A[712]), .B(n314), .CI(
        C[712]), .S(S[712]), .CO(C[713]) );
  FA_13939 \FA_INST_0[1].FA_INST_1[201].FA_  ( .A(A[713]), .B(n313), .CI(
        C[713]), .S(S[713]), .CO(C[714]) );
  FA_13938 \FA_INST_0[1].FA_INST_1[202].FA_  ( .A(A[714]), .B(n312), .CI(
        C[714]), .S(S[714]), .CO(C[715]) );
  FA_13937 \FA_INST_0[1].FA_INST_1[203].FA_  ( .A(A[715]), .B(n311), .CI(
        C[715]), .S(S[715]), .CO(C[716]) );
  FA_13936 \FA_INST_0[1].FA_INST_1[204].FA_  ( .A(A[716]), .B(n310), .CI(
        C[716]), .S(S[716]), .CO(C[717]) );
  FA_13935 \FA_INST_0[1].FA_INST_1[205].FA_  ( .A(A[717]), .B(n309), .CI(
        C[717]), .S(S[717]), .CO(C[718]) );
  FA_13934 \FA_INST_0[1].FA_INST_1[206].FA_  ( .A(A[718]), .B(n308), .CI(
        C[718]), .S(S[718]), .CO(C[719]) );
  FA_13933 \FA_INST_0[1].FA_INST_1[207].FA_  ( .A(A[719]), .B(n307), .CI(
        C[719]), .S(S[719]), .CO(C[720]) );
  FA_13932 \FA_INST_0[1].FA_INST_1[208].FA_  ( .A(A[720]), .B(n306), .CI(
        C[720]), .S(S[720]), .CO(C[721]) );
  FA_13931 \FA_INST_0[1].FA_INST_1[209].FA_  ( .A(A[721]), .B(n305), .CI(
        C[721]), .S(S[721]), .CO(C[722]) );
  FA_13930 \FA_INST_0[1].FA_INST_1[210].FA_  ( .A(A[722]), .B(n304), .CI(
        C[722]), .S(S[722]), .CO(C[723]) );
  FA_13929 \FA_INST_0[1].FA_INST_1[211].FA_  ( .A(A[723]), .B(n303), .CI(
        C[723]), .S(S[723]), .CO(C[724]) );
  FA_13928 \FA_INST_0[1].FA_INST_1[212].FA_  ( .A(A[724]), .B(n302), .CI(
        C[724]), .S(S[724]), .CO(C[725]) );
  FA_13927 \FA_INST_0[1].FA_INST_1[213].FA_  ( .A(A[725]), .B(n301), .CI(
        C[725]), .S(S[725]), .CO(C[726]) );
  FA_13926 \FA_INST_0[1].FA_INST_1[214].FA_  ( .A(A[726]), .B(n300), .CI(
        C[726]), .S(S[726]), .CO(C[727]) );
  FA_13925 \FA_INST_0[1].FA_INST_1[215].FA_  ( .A(A[727]), .B(n299), .CI(
        C[727]), .S(S[727]), .CO(C[728]) );
  FA_13924 \FA_INST_0[1].FA_INST_1[216].FA_  ( .A(A[728]), .B(n298), .CI(
        C[728]), .S(S[728]), .CO(C[729]) );
  FA_13923 \FA_INST_0[1].FA_INST_1[217].FA_  ( .A(A[729]), .B(n297), .CI(
        C[729]), .S(S[729]), .CO(C[730]) );
  FA_13922 \FA_INST_0[1].FA_INST_1[218].FA_  ( .A(A[730]), .B(n296), .CI(
        C[730]), .S(S[730]), .CO(C[731]) );
  FA_13921 \FA_INST_0[1].FA_INST_1[219].FA_  ( .A(A[731]), .B(n295), .CI(
        C[731]), .S(S[731]), .CO(C[732]) );
  FA_13920 \FA_INST_0[1].FA_INST_1[220].FA_  ( .A(A[732]), .B(n294), .CI(
        C[732]), .S(S[732]), .CO(C[733]) );
  FA_13919 \FA_INST_0[1].FA_INST_1[221].FA_  ( .A(A[733]), .B(n293), .CI(
        C[733]), .S(S[733]), .CO(C[734]) );
  FA_13918 \FA_INST_0[1].FA_INST_1[222].FA_  ( .A(A[734]), .B(n292), .CI(
        C[734]), .S(S[734]), .CO(C[735]) );
  FA_13917 \FA_INST_0[1].FA_INST_1[223].FA_  ( .A(A[735]), .B(n291), .CI(
        C[735]), .S(S[735]), .CO(C[736]) );
  FA_13916 \FA_INST_0[1].FA_INST_1[224].FA_  ( .A(A[736]), .B(n290), .CI(
        C[736]), .S(S[736]), .CO(C[737]) );
  FA_13915 \FA_INST_0[1].FA_INST_1[225].FA_  ( .A(A[737]), .B(n289), .CI(
        C[737]), .S(S[737]), .CO(C[738]) );
  FA_13914 \FA_INST_0[1].FA_INST_1[226].FA_  ( .A(A[738]), .B(n288), .CI(
        C[738]), .S(S[738]), .CO(C[739]) );
  FA_13913 \FA_INST_0[1].FA_INST_1[227].FA_  ( .A(A[739]), .B(n287), .CI(
        C[739]), .S(S[739]), .CO(C[740]) );
  FA_13912 \FA_INST_0[1].FA_INST_1[228].FA_  ( .A(A[740]), .B(n286), .CI(
        C[740]), .S(S[740]), .CO(C[741]) );
  FA_13911 \FA_INST_0[1].FA_INST_1[229].FA_  ( .A(A[741]), .B(n285), .CI(
        C[741]), .S(S[741]), .CO(C[742]) );
  FA_13910 \FA_INST_0[1].FA_INST_1[230].FA_  ( .A(A[742]), .B(n284), .CI(
        C[742]), .S(S[742]), .CO(C[743]) );
  FA_13909 \FA_INST_0[1].FA_INST_1[231].FA_  ( .A(A[743]), .B(n283), .CI(
        C[743]), .S(S[743]), .CO(C[744]) );
  FA_13908 \FA_INST_0[1].FA_INST_1[232].FA_  ( .A(A[744]), .B(n282), .CI(
        C[744]), .S(S[744]), .CO(C[745]) );
  FA_13907 \FA_INST_0[1].FA_INST_1[233].FA_  ( .A(A[745]), .B(n281), .CI(
        C[745]), .S(S[745]), .CO(C[746]) );
  FA_13906 \FA_INST_0[1].FA_INST_1[234].FA_  ( .A(A[746]), .B(n280), .CI(
        C[746]), .S(S[746]), .CO(C[747]) );
  FA_13905 \FA_INST_0[1].FA_INST_1[235].FA_  ( .A(A[747]), .B(n279), .CI(
        C[747]), .S(S[747]), .CO(C[748]) );
  FA_13904 \FA_INST_0[1].FA_INST_1[236].FA_  ( .A(A[748]), .B(n278), .CI(
        C[748]), .S(S[748]), .CO(C[749]) );
  FA_13903 \FA_INST_0[1].FA_INST_1[237].FA_  ( .A(A[749]), .B(n277), .CI(
        C[749]), .S(S[749]), .CO(C[750]) );
  FA_13902 \FA_INST_0[1].FA_INST_1[238].FA_  ( .A(A[750]), .B(n276), .CI(
        C[750]), .S(S[750]), .CO(C[751]) );
  FA_13901 \FA_INST_0[1].FA_INST_1[239].FA_  ( .A(A[751]), .B(n275), .CI(
        C[751]), .S(S[751]), .CO(C[752]) );
  FA_13900 \FA_INST_0[1].FA_INST_1[240].FA_  ( .A(A[752]), .B(n274), .CI(
        C[752]), .S(S[752]), .CO(C[753]) );
  FA_13899 \FA_INST_0[1].FA_INST_1[241].FA_  ( .A(A[753]), .B(n273), .CI(
        C[753]), .S(S[753]), .CO(C[754]) );
  FA_13898 \FA_INST_0[1].FA_INST_1[242].FA_  ( .A(A[754]), .B(n272), .CI(
        C[754]), .S(S[754]), .CO(C[755]) );
  FA_13897 \FA_INST_0[1].FA_INST_1[243].FA_  ( .A(A[755]), .B(n271), .CI(
        C[755]), .S(S[755]), .CO(C[756]) );
  FA_13896 \FA_INST_0[1].FA_INST_1[244].FA_  ( .A(A[756]), .B(n270), .CI(
        C[756]), .S(S[756]), .CO(C[757]) );
  FA_13895 \FA_INST_0[1].FA_INST_1[245].FA_  ( .A(A[757]), .B(n269), .CI(
        C[757]), .S(S[757]), .CO(C[758]) );
  FA_13894 \FA_INST_0[1].FA_INST_1[246].FA_  ( .A(A[758]), .B(n268), .CI(
        C[758]), .S(S[758]), .CO(C[759]) );
  FA_13893 \FA_INST_0[1].FA_INST_1[247].FA_  ( .A(A[759]), .B(n267), .CI(
        C[759]), .S(S[759]), .CO(C[760]) );
  FA_13892 \FA_INST_0[1].FA_INST_1[248].FA_  ( .A(A[760]), .B(n266), .CI(
        C[760]), .S(S[760]), .CO(C[761]) );
  FA_13891 \FA_INST_0[1].FA_INST_1[249].FA_  ( .A(A[761]), .B(n265), .CI(
        C[761]), .S(S[761]), .CO(C[762]) );
  FA_13890 \FA_INST_0[1].FA_INST_1[250].FA_  ( .A(A[762]), .B(n264), .CI(
        C[762]), .S(S[762]), .CO(C[763]) );
  FA_13889 \FA_INST_0[1].FA_INST_1[251].FA_  ( .A(A[763]), .B(n263), .CI(
        C[763]), .S(S[763]), .CO(C[764]) );
  FA_13888 \FA_INST_0[1].FA_INST_1[252].FA_  ( .A(A[764]), .B(n262), .CI(
        C[764]), .S(S[764]), .CO(C[765]) );
  FA_13887 \FA_INST_0[1].FA_INST_1[253].FA_  ( .A(A[765]), .B(n261), .CI(
        C[765]), .S(S[765]), .CO(C[766]) );
  FA_13886 \FA_INST_0[1].FA_INST_1[254].FA_  ( .A(A[766]), .B(n260), .CI(
        C[766]), .S(S[766]), .CO(C[767]) );
  FA_13885 \FA_INST_0[1].FA_INST_1[255].FA_  ( .A(A[767]), .B(n259), .CI(
        C[767]), .S(S[767]), .CO(C[768]) );
  FA_13884 \FA_INST_0[1].FA_INST_1[256].FA_  ( .A(A[768]), .B(n258), .CI(
        C[768]), .S(S[768]), .CO(C[769]) );
  FA_13883 \FA_INST_0[1].FA_INST_1[257].FA_  ( .A(A[769]), .B(n257), .CI(
        C[769]), .S(S[769]), .CO(C[770]) );
  FA_13882 \FA_INST_0[1].FA_INST_1[258].FA_  ( .A(A[770]), .B(n256), .CI(
        C[770]), .S(S[770]), .CO(C[771]) );
  FA_13881 \FA_INST_0[1].FA_INST_1[259].FA_  ( .A(A[771]), .B(n255), .CI(
        C[771]), .S(S[771]), .CO(C[772]) );
  FA_13880 \FA_INST_0[1].FA_INST_1[260].FA_  ( .A(A[772]), .B(n254), .CI(
        C[772]), .S(S[772]), .CO(C[773]) );
  FA_13879 \FA_INST_0[1].FA_INST_1[261].FA_  ( .A(A[773]), .B(n253), .CI(
        C[773]), .S(S[773]), .CO(C[774]) );
  FA_13878 \FA_INST_0[1].FA_INST_1[262].FA_  ( .A(A[774]), .B(n252), .CI(
        C[774]), .S(S[774]), .CO(C[775]) );
  FA_13877 \FA_INST_0[1].FA_INST_1[263].FA_  ( .A(A[775]), .B(n251), .CI(
        C[775]), .S(S[775]), .CO(C[776]) );
  FA_13876 \FA_INST_0[1].FA_INST_1[264].FA_  ( .A(A[776]), .B(n250), .CI(
        C[776]), .S(S[776]), .CO(C[777]) );
  FA_13875 \FA_INST_0[1].FA_INST_1[265].FA_  ( .A(A[777]), .B(n249), .CI(
        C[777]), .S(S[777]), .CO(C[778]) );
  FA_13874 \FA_INST_0[1].FA_INST_1[266].FA_  ( .A(A[778]), .B(n248), .CI(
        C[778]), .S(S[778]), .CO(C[779]) );
  FA_13873 \FA_INST_0[1].FA_INST_1[267].FA_  ( .A(A[779]), .B(n247), .CI(
        C[779]), .S(S[779]), .CO(C[780]) );
  FA_13872 \FA_INST_0[1].FA_INST_1[268].FA_  ( .A(A[780]), .B(n246), .CI(
        C[780]), .S(S[780]), .CO(C[781]) );
  FA_13871 \FA_INST_0[1].FA_INST_1[269].FA_  ( .A(A[781]), .B(n245), .CI(
        C[781]), .S(S[781]), .CO(C[782]) );
  FA_13870 \FA_INST_0[1].FA_INST_1[270].FA_  ( .A(A[782]), .B(n244), .CI(
        C[782]), .S(S[782]), .CO(C[783]) );
  FA_13869 \FA_INST_0[1].FA_INST_1[271].FA_  ( .A(A[783]), .B(n243), .CI(
        C[783]), .S(S[783]), .CO(C[784]) );
  FA_13868 \FA_INST_0[1].FA_INST_1[272].FA_  ( .A(A[784]), .B(n242), .CI(
        C[784]), .S(S[784]), .CO(C[785]) );
  FA_13867 \FA_INST_0[1].FA_INST_1[273].FA_  ( .A(A[785]), .B(n241), .CI(
        C[785]), .S(S[785]), .CO(C[786]) );
  FA_13866 \FA_INST_0[1].FA_INST_1[274].FA_  ( .A(A[786]), .B(n240), .CI(
        C[786]), .S(S[786]), .CO(C[787]) );
  FA_13865 \FA_INST_0[1].FA_INST_1[275].FA_  ( .A(A[787]), .B(n239), .CI(
        C[787]), .S(S[787]), .CO(C[788]) );
  FA_13864 \FA_INST_0[1].FA_INST_1[276].FA_  ( .A(A[788]), .B(n238), .CI(
        C[788]), .S(S[788]), .CO(C[789]) );
  FA_13863 \FA_INST_0[1].FA_INST_1[277].FA_  ( .A(A[789]), .B(n237), .CI(
        C[789]), .S(S[789]), .CO(C[790]) );
  FA_13862 \FA_INST_0[1].FA_INST_1[278].FA_  ( .A(A[790]), .B(n236), .CI(
        C[790]), .S(S[790]), .CO(C[791]) );
  FA_13861 \FA_INST_0[1].FA_INST_1[279].FA_  ( .A(A[791]), .B(n235), .CI(
        C[791]), .S(S[791]), .CO(C[792]) );
  FA_13860 \FA_INST_0[1].FA_INST_1[280].FA_  ( .A(A[792]), .B(n234), .CI(
        C[792]), .S(S[792]), .CO(C[793]) );
  FA_13859 \FA_INST_0[1].FA_INST_1[281].FA_  ( .A(A[793]), .B(n233), .CI(
        C[793]), .S(S[793]), .CO(C[794]) );
  FA_13858 \FA_INST_0[1].FA_INST_1[282].FA_  ( .A(A[794]), .B(n232), .CI(
        C[794]), .S(S[794]), .CO(C[795]) );
  FA_13857 \FA_INST_0[1].FA_INST_1[283].FA_  ( .A(A[795]), .B(n231), .CI(
        C[795]), .S(S[795]), .CO(C[796]) );
  FA_13856 \FA_INST_0[1].FA_INST_1[284].FA_  ( .A(A[796]), .B(n230), .CI(
        C[796]), .S(S[796]), .CO(C[797]) );
  FA_13855 \FA_INST_0[1].FA_INST_1[285].FA_  ( .A(A[797]), .B(n229), .CI(
        C[797]), .S(S[797]), .CO(C[798]) );
  FA_13854 \FA_INST_0[1].FA_INST_1[286].FA_  ( .A(A[798]), .B(n228), .CI(
        C[798]), .S(S[798]), .CO(C[799]) );
  FA_13853 \FA_INST_0[1].FA_INST_1[287].FA_  ( .A(A[799]), .B(n227), .CI(
        C[799]), .S(S[799]), .CO(C[800]) );
  FA_13852 \FA_INST_0[1].FA_INST_1[288].FA_  ( .A(A[800]), .B(n226), .CI(
        C[800]), .S(S[800]), .CO(C[801]) );
  FA_13851 \FA_INST_0[1].FA_INST_1[289].FA_  ( .A(A[801]), .B(n225), .CI(
        C[801]), .S(S[801]), .CO(C[802]) );
  FA_13850 \FA_INST_0[1].FA_INST_1[290].FA_  ( .A(A[802]), .B(n224), .CI(
        C[802]), .S(S[802]), .CO(C[803]) );
  FA_13849 \FA_INST_0[1].FA_INST_1[291].FA_  ( .A(A[803]), .B(n223), .CI(
        C[803]), .S(S[803]), .CO(C[804]) );
  FA_13848 \FA_INST_0[1].FA_INST_1[292].FA_  ( .A(A[804]), .B(n222), .CI(
        C[804]), .S(S[804]), .CO(C[805]) );
  FA_13847 \FA_INST_0[1].FA_INST_1[293].FA_  ( .A(A[805]), .B(n221), .CI(
        C[805]), .S(S[805]), .CO(C[806]) );
  FA_13846 \FA_INST_0[1].FA_INST_1[294].FA_  ( .A(A[806]), .B(n220), .CI(
        C[806]), .S(S[806]), .CO(C[807]) );
  FA_13845 \FA_INST_0[1].FA_INST_1[295].FA_  ( .A(A[807]), .B(n219), .CI(
        C[807]), .S(S[807]), .CO(C[808]) );
  FA_13844 \FA_INST_0[1].FA_INST_1[296].FA_  ( .A(A[808]), .B(n218), .CI(
        C[808]), .S(S[808]), .CO(C[809]) );
  FA_13843 \FA_INST_0[1].FA_INST_1[297].FA_  ( .A(A[809]), .B(n217), .CI(
        C[809]), .S(S[809]), .CO(C[810]) );
  FA_13842 \FA_INST_0[1].FA_INST_1[298].FA_  ( .A(A[810]), .B(n216), .CI(
        C[810]), .S(S[810]), .CO(C[811]) );
  FA_13841 \FA_INST_0[1].FA_INST_1[299].FA_  ( .A(A[811]), .B(n215), .CI(
        C[811]), .S(S[811]), .CO(C[812]) );
  FA_13840 \FA_INST_0[1].FA_INST_1[300].FA_  ( .A(A[812]), .B(n214), .CI(
        C[812]), .S(S[812]), .CO(C[813]) );
  FA_13839 \FA_INST_0[1].FA_INST_1[301].FA_  ( .A(A[813]), .B(n213), .CI(
        C[813]), .S(S[813]), .CO(C[814]) );
  FA_13838 \FA_INST_0[1].FA_INST_1[302].FA_  ( .A(A[814]), .B(n212), .CI(
        C[814]), .S(S[814]), .CO(C[815]) );
  FA_13837 \FA_INST_0[1].FA_INST_1[303].FA_  ( .A(A[815]), .B(n211), .CI(
        C[815]), .S(S[815]), .CO(C[816]) );
  FA_13836 \FA_INST_0[1].FA_INST_1[304].FA_  ( .A(A[816]), .B(n210), .CI(
        C[816]), .S(S[816]), .CO(C[817]) );
  FA_13835 \FA_INST_0[1].FA_INST_1[305].FA_  ( .A(A[817]), .B(n209), .CI(
        C[817]), .S(S[817]), .CO(C[818]) );
  FA_13834 \FA_INST_0[1].FA_INST_1[306].FA_  ( .A(A[818]), .B(n208), .CI(
        C[818]), .S(S[818]), .CO(C[819]) );
  FA_13833 \FA_INST_0[1].FA_INST_1[307].FA_  ( .A(A[819]), .B(n207), .CI(
        C[819]), .S(S[819]), .CO(C[820]) );
  FA_13832 \FA_INST_0[1].FA_INST_1[308].FA_  ( .A(A[820]), .B(n206), .CI(
        C[820]), .S(S[820]), .CO(C[821]) );
  FA_13831 \FA_INST_0[1].FA_INST_1[309].FA_  ( .A(A[821]), .B(n205), .CI(
        C[821]), .S(S[821]), .CO(C[822]) );
  FA_13830 \FA_INST_0[1].FA_INST_1[310].FA_  ( .A(A[822]), .B(n204), .CI(
        C[822]), .S(S[822]), .CO(C[823]) );
  FA_13829 \FA_INST_0[1].FA_INST_1[311].FA_  ( .A(A[823]), .B(n203), .CI(
        C[823]), .S(S[823]), .CO(C[824]) );
  FA_13828 \FA_INST_0[1].FA_INST_1[312].FA_  ( .A(A[824]), .B(n202), .CI(
        C[824]), .S(S[824]), .CO(C[825]) );
  FA_13827 \FA_INST_0[1].FA_INST_1[313].FA_  ( .A(A[825]), .B(n201), .CI(
        C[825]), .S(S[825]), .CO(C[826]) );
  FA_13826 \FA_INST_0[1].FA_INST_1[314].FA_  ( .A(A[826]), .B(n200), .CI(
        C[826]), .S(S[826]), .CO(C[827]) );
  FA_13825 \FA_INST_0[1].FA_INST_1[315].FA_  ( .A(A[827]), .B(n199), .CI(
        C[827]), .S(S[827]), .CO(C[828]) );
  FA_13824 \FA_INST_0[1].FA_INST_1[316].FA_  ( .A(A[828]), .B(n198), .CI(
        C[828]), .S(S[828]), .CO(C[829]) );
  FA_13823 \FA_INST_0[1].FA_INST_1[317].FA_  ( .A(A[829]), .B(n197), .CI(
        C[829]), .S(S[829]), .CO(C[830]) );
  FA_13822 \FA_INST_0[1].FA_INST_1[318].FA_  ( .A(A[830]), .B(n196), .CI(
        C[830]), .S(S[830]), .CO(C[831]) );
  FA_13821 \FA_INST_0[1].FA_INST_1[319].FA_  ( .A(A[831]), .B(n195), .CI(
        C[831]), .S(S[831]), .CO(C[832]) );
  FA_13820 \FA_INST_0[1].FA_INST_1[320].FA_  ( .A(A[832]), .B(n194), .CI(
        C[832]), .S(S[832]), .CO(C[833]) );
  FA_13819 \FA_INST_0[1].FA_INST_1[321].FA_  ( .A(A[833]), .B(n193), .CI(
        C[833]), .S(S[833]), .CO(C[834]) );
  FA_13818 \FA_INST_0[1].FA_INST_1[322].FA_  ( .A(A[834]), .B(n192), .CI(
        C[834]), .S(S[834]), .CO(C[835]) );
  FA_13817 \FA_INST_0[1].FA_INST_1[323].FA_  ( .A(A[835]), .B(n191), .CI(
        C[835]), .S(S[835]), .CO(C[836]) );
  FA_13816 \FA_INST_0[1].FA_INST_1[324].FA_  ( .A(A[836]), .B(n190), .CI(
        C[836]), .S(S[836]), .CO(C[837]) );
  FA_13815 \FA_INST_0[1].FA_INST_1[325].FA_  ( .A(A[837]), .B(n189), .CI(
        C[837]), .S(S[837]), .CO(C[838]) );
  FA_13814 \FA_INST_0[1].FA_INST_1[326].FA_  ( .A(A[838]), .B(n188), .CI(
        C[838]), .S(S[838]), .CO(C[839]) );
  FA_13813 \FA_INST_0[1].FA_INST_1[327].FA_  ( .A(A[839]), .B(n187), .CI(
        C[839]), .S(S[839]), .CO(C[840]) );
  FA_13812 \FA_INST_0[1].FA_INST_1[328].FA_  ( .A(A[840]), .B(n186), .CI(
        C[840]), .S(S[840]), .CO(C[841]) );
  FA_13811 \FA_INST_0[1].FA_INST_1[329].FA_  ( .A(A[841]), .B(n185), .CI(
        C[841]), .S(S[841]), .CO(C[842]) );
  FA_13810 \FA_INST_0[1].FA_INST_1[330].FA_  ( .A(A[842]), .B(n184), .CI(
        C[842]), .S(S[842]), .CO(C[843]) );
  FA_13809 \FA_INST_0[1].FA_INST_1[331].FA_  ( .A(A[843]), .B(n183), .CI(
        C[843]), .S(S[843]), .CO(C[844]) );
  FA_13808 \FA_INST_0[1].FA_INST_1[332].FA_  ( .A(A[844]), .B(n182), .CI(
        C[844]), .S(S[844]), .CO(C[845]) );
  FA_13807 \FA_INST_0[1].FA_INST_1[333].FA_  ( .A(A[845]), .B(n181), .CI(
        C[845]), .S(S[845]), .CO(C[846]) );
  FA_13806 \FA_INST_0[1].FA_INST_1[334].FA_  ( .A(A[846]), .B(n180), .CI(
        C[846]), .S(S[846]), .CO(C[847]) );
  FA_13805 \FA_INST_0[1].FA_INST_1[335].FA_  ( .A(A[847]), .B(n179), .CI(
        C[847]), .S(S[847]), .CO(C[848]) );
  FA_13804 \FA_INST_0[1].FA_INST_1[336].FA_  ( .A(A[848]), .B(n178), .CI(
        C[848]), .S(S[848]), .CO(C[849]) );
  FA_13803 \FA_INST_0[1].FA_INST_1[337].FA_  ( .A(A[849]), .B(n177), .CI(
        C[849]), .S(S[849]), .CO(C[850]) );
  FA_13802 \FA_INST_0[1].FA_INST_1[338].FA_  ( .A(A[850]), .B(n176), .CI(
        C[850]), .S(S[850]), .CO(C[851]) );
  FA_13801 \FA_INST_0[1].FA_INST_1[339].FA_  ( .A(A[851]), .B(n175), .CI(
        C[851]), .S(S[851]), .CO(C[852]) );
  FA_13800 \FA_INST_0[1].FA_INST_1[340].FA_  ( .A(A[852]), .B(n174), .CI(
        C[852]), .S(S[852]), .CO(C[853]) );
  FA_13799 \FA_INST_0[1].FA_INST_1[341].FA_  ( .A(A[853]), .B(n173), .CI(
        C[853]), .S(S[853]), .CO(C[854]) );
  FA_13798 \FA_INST_0[1].FA_INST_1[342].FA_  ( .A(A[854]), .B(n172), .CI(
        C[854]), .S(S[854]), .CO(C[855]) );
  FA_13797 \FA_INST_0[1].FA_INST_1[343].FA_  ( .A(A[855]), .B(n171), .CI(
        C[855]), .S(S[855]), .CO(C[856]) );
  FA_13796 \FA_INST_0[1].FA_INST_1[344].FA_  ( .A(A[856]), .B(n170), .CI(
        C[856]), .S(S[856]), .CO(C[857]) );
  FA_13795 \FA_INST_0[1].FA_INST_1[345].FA_  ( .A(A[857]), .B(n169), .CI(
        C[857]), .S(S[857]), .CO(C[858]) );
  FA_13794 \FA_INST_0[1].FA_INST_1[346].FA_  ( .A(A[858]), .B(n168), .CI(
        C[858]), .S(S[858]), .CO(C[859]) );
  FA_13793 \FA_INST_0[1].FA_INST_1[347].FA_  ( .A(A[859]), .B(n167), .CI(
        C[859]), .S(S[859]), .CO(C[860]) );
  FA_13792 \FA_INST_0[1].FA_INST_1[348].FA_  ( .A(A[860]), .B(n166), .CI(
        C[860]), .S(S[860]), .CO(C[861]) );
  FA_13791 \FA_INST_0[1].FA_INST_1[349].FA_  ( .A(A[861]), .B(n165), .CI(
        C[861]), .S(S[861]), .CO(C[862]) );
  FA_13790 \FA_INST_0[1].FA_INST_1[350].FA_  ( .A(A[862]), .B(n164), .CI(
        C[862]), .S(S[862]), .CO(C[863]) );
  FA_13789 \FA_INST_0[1].FA_INST_1[351].FA_  ( .A(A[863]), .B(n163), .CI(
        C[863]), .S(S[863]), .CO(C[864]) );
  FA_13788 \FA_INST_0[1].FA_INST_1[352].FA_  ( .A(A[864]), .B(n162), .CI(
        C[864]), .S(S[864]), .CO(C[865]) );
  FA_13787 \FA_INST_0[1].FA_INST_1[353].FA_  ( .A(A[865]), .B(n161), .CI(
        C[865]), .S(S[865]), .CO(C[866]) );
  FA_13786 \FA_INST_0[1].FA_INST_1[354].FA_  ( .A(A[866]), .B(n160), .CI(
        C[866]), .S(S[866]), .CO(C[867]) );
  FA_13785 \FA_INST_0[1].FA_INST_1[355].FA_  ( .A(A[867]), .B(n159), .CI(
        C[867]), .S(S[867]), .CO(C[868]) );
  FA_13784 \FA_INST_0[1].FA_INST_1[356].FA_  ( .A(A[868]), .B(n158), .CI(
        C[868]), .S(S[868]), .CO(C[869]) );
  FA_13783 \FA_INST_0[1].FA_INST_1[357].FA_  ( .A(A[869]), .B(n157), .CI(
        C[869]), .S(S[869]), .CO(C[870]) );
  FA_13782 \FA_INST_0[1].FA_INST_1[358].FA_  ( .A(A[870]), .B(n156), .CI(
        C[870]), .S(S[870]), .CO(C[871]) );
  FA_13781 \FA_INST_0[1].FA_INST_1[359].FA_  ( .A(A[871]), .B(n155), .CI(
        C[871]), .S(S[871]), .CO(C[872]) );
  FA_13780 \FA_INST_0[1].FA_INST_1[360].FA_  ( .A(A[872]), .B(n154), .CI(
        C[872]), .S(S[872]), .CO(C[873]) );
  FA_13779 \FA_INST_0[1].FA_INST_1[361].FA_  ( .A(A[873]), .B(n153), .CI(
        C[873]), .S(S[873]), .CO(C[874]) );
  FA_13778 \FA_INST_0[1].FA_INST_1[362].FA_  ( .A(A[874]), .B(n152), .CI(
        C[874]), .S(S[874]), .CO(C[875]) );
  FA_13777 \FA_INST_0[1].FA_INST_1[363].FA_  ( .A(A[875]), .B(n151), .CI(
        C[875]), .S(S[875]), .CO(C[876]) );
  FA_13776 \FA_INST_0[1].FA_INST_1[364].FA_  ( .A(A[876]), .B(n150), .CI(
        C[876]), .S(S[876]), .CO(C[877]) );
  FA_13775 \FA_INST_0[1].FA_INST_1[365].FA_  ( .A(A[877]), .B(n149), .CI(
        C[877]), .S(S[877]), .CO(C[878]) );
  FA_13774 \FA_INST_0[1].FA_INST_1[366].FA_  ( .A(A[878]), .B(n148), .CI(
        C[878]), .S(S[878]), .CO(C[879]) );
  FA_13773 \FA_INST_0[1].FA_INST_1[367].FA_  ( .A(A[879]), .B(n147), .CI(
        C[879]), .S(S[879]), .CO(C[880]) );
  FA_13772 \FA_INST_0[1].FA_INST_1[368].FA_  ( .A(A[880]), .B(n146), .CI(
        C[880]), .S(S[880]), .CO(C[881]) );
  FA_13771 \FA_INST_0[1].FA_INST_1[369].FA_  ( .A(A[881]), .B(n145), .CI(
        C[881]), .S(S[881]), .CO(C[882]) );
  FA_13770 \FA_INST_0[1].FA_INST_1[370].FA_  ( .A(A[882]), .B(n144), .CI(
        C[882]), .S(S[882]), .CO(C[883]) );
  FA_13769 \FA_INST_0[1].FA_INST_1[371].FA_  ( .A(A[883]), .B(n143), .CI(
        C[883]), .S(S[883]), .CO(C[884]) );
  FA_13768 \FA_INST_0[1].FA_INST_1[372].FA_  ( .A(A[884]), .B(n142), .CI(
        C[884]), .S(S[884]), .CO(C[885]) );
  FA_13767 \FA_INST_0[1].FA_INST_1[373].FA_  ( .A(A[885]), .B(n141), .CI(
        C[885]), .S(S[885]), .CO(C[886]) );
  FA_13766 \FA_INST_0[1].FA_INST_1[374].FA_  ( .A(A[886]), .B(n140), .CI(
        C[886]), .S(S[886]), .CO(C[887]) );
  FA_13765 \FA_INST_0[1].FA_INST_1[375].FA_  ( .A(A[887]), .B(n139), .CI(
        C[887]), .S(S[887]), .CO(C[888]) );
  FA_13764 \FA_INST_0[1].FA_INST_1[376].FA_  ( .A(A[888]), .B(n138), .CI(
        C[888]), .S(S[888]), .CO(C[889]) );
  FA_13763 \FA_INST_0[1].FA_INST_1[377].FA_  ( .A(A[889]), .B(n137), .CI(
        C[889]), .S(S[889]), .CO(C[890]) );
  FA_13762 \FA_INST_0[1].FA_INST_1[378].FA_  ( .A(A[890]), .B(n136), .CI(
        C[890]), .S(S[890]), .CO(C[891]) );
  FA_13761 \FA_INST_0[1].FA_INST_1[379].FA_  ( .A(A[891]), .B(n135), .CI(
        C[891]), .S(S[891]), .CO(C[892]) );
  FA_13760 \FA_INST_0[1].FA_INST_1[380].FA_  ( .A(A[892]), .B(n134), .CI(
        C[892]), .S(S[892]), .CO(C[893]) );
  FA_13759 \FA_INST_0[1].FA_INST_1[381].FA_  ( .A(A[893]), .B(n133), .CI(
        C[893]), .S(S[893]), .CO(C[894]) );
  FA_13758 \FA_INST_0[1].FA_INST_1[382].FA_  ( .A(A[894]), .B(n132), .CI(
        C[894]), .S(S[894]), .CO(C[895]) );
  FA_13757 \FA_INST_0[1].FA_INST_1[383].FA_  ( .A(A[895]), .B(n131), .CI(
        C[895]), .S(S[895]), .CO(C[896]) );
  FA_13756 \FA_INST_0[1].FA_INST_1[384].FA_  ( .A(A[896]), .B(n130), .CI(
        C[896]), .S(S[896]), .CO(C[897]) );
  FA_13755 \FA_INST_0[1].FA_INST_1[385].FA_  ( .A(A[897]), .B(n129), .CI(
        C[897]), .S(S[897]), .CO(C[898]) );
  FA_13754 \FA_INST_0[1].FA_INST_1[386].FA_  ( .A(A[898]), .B(n128), .CI(
        C[898]), .S(S[898]), .CO(C[899]) );
  FA_13753 \FA_INST_0[1].FA_INST_1[387].FA_  ( .A(A[899]), .B(n127), .CI(
        C[899]), .S(S[899]), .CO(C[900]) );
  FA_13752 \FA_INST_0[1].FA_INST_1[388].FA_  ( .A(A[900]), .B(n126), .CI(
        C[900]), .S(S[900]), .CO(C[901]) );
  FA_13751 \FA_INST_0[1].FA_INST_1[389].FA_  ( .A(A[901]), .B(n125), .CI(
        C[901]), .S(S[901]), .CO(C[902]) );
  FA_13750 \FA_INST_0[1].FA_INST_1[390].FA_  ( .A(A[902]), .B(n124), .CI(
        C[902]), .S(S[902]), .CO(C[903]) );
  FA_13749 \FA_INST_0[1].FA_INST_1[391].FA_  ( .A(A[903]), .B(n123), .CI(
        C[903]), .S(S[903]), .CO(C[904]) );
  FA_13748 \FA_INST_0[1].FA_INST_1[392].FA_  ( .A(A[904]), .B(n122), .CI(
        C[904]), .S(S[904]), .CO(C[905]) );
  FA_13747 \FA_INST_0[1].FA_INST_1[393].FA_  ( .A(A[905]), .B(n121), .CI(
        C[905]), .S(S[905]), .CO(C[906]) );
  FA_13746 \FA_INST_0[1].FA_INST_1[394].FA_  ( .A(A[906]), .B(n120), .CI(
        C[906]), .S(S[906]), .CO(C[907]) );
  FA_13745 \FA_INST_0[1].FA_INST_1[395].FA_  ( .A(A[907]), .B(n119), .CI(
        C[907]), .S(S[907]), .CO(C[908]) );
  FA_13744 \FA_INST_0[1].FA_INST_1[396].FA_  ( .A(A[908]), .B(n118), .CI(
        C[908]), .S(S[908]), .CO(C[909]) );
  FA_13743 \FA_INST_0[1].FA_INST_1[397].FA_  ( .A(A[909]), .B(n117), .CI(
        C[909]), .S(S[909]), .CO(C[910]) );
  FA_13742 \FA_INST_0[1].FA_INST_1[398].FA_  ( .A(A[910]), .B(n116), .CI(
        C[910]), .S(S[910]), .CO(C[911]) );
  FA_13741 \FA_INST_0[1].FA_INST_1[399].FA_  ( .A(A[911]), .B(n115), .CI(
        C[911]), .S(S[911]), .CO(C[912]) );
  FA_13740 \FA_INST_0[1].FA_INST_1[400].FA_  ( .A(A[912]), .B(n114), .CI(
        C[912]), .S(S[912]), .CO(C[913]) );
  FA_13739 \FA_INST_0[1].FA_INST_1[401].FA_  ( .A(A[913]), .B(n113), .CI(
        C[913]), .S(S[913]), .CO(C[914]) );
  FA_13738 \FA_INST_0[1].FA_INST_1[402].FA_  ( .A(A[914]), .B(n112), .CI(
        C[914]), .S(S[914]), .CO(C[915]) );
  FA_13737 \FA_INST_0[1].FA_INST_1[403].FA_  ( .A(A[915]), .B(n111), .CI(
        C[915]), .S(S[915]), .CO(C[916]) );
  FA_13736 \FA_INST_0[1].FA_INST_1[404].FA_  ( .A(A[916]), .B(n110), .CI(
        C[916]), .S(S[916]), .CO(C[917]) );
  FA_13735 \FA_INST_0[1].FA_INST_1[405].FA_  ( .A(A[917]), .B(n109), .CI(
        C[917]), .S(S[917]), .CO(C[918]) );
  FA_13734 \FA_INST_0[1].FA_INST_1[406].FA_  ( .A(A[918]), .B(n108), .CI(
        C[918]), .S(S[918]), .CO(C[919]) );
  FA_13733 \FA_INST_0[1].FA_INST_1[407].FA_  ( .A(A[919]), .B(n107), .CI(
        C[919]), .S(S[919]), .CO(C[920]) );
  FA_13732 \FA_INST_0[1].FA_INST_1[408].FA_  ( .A(A[920]), .B(n106), .CI(
        C[920]), .S(S[920]), .CO(C[921]) );
  FA_13731 \FA_INST_0[1].FA_INST_1[409].FA_  ( .A(A[921]), .B(n105), .CI(
        C[921]), .S(S[921]), .CO(C[922]) );
  FA_13730 \FA_INST_0[1].FA_INST_1[410].FA_  ( .A(A[922]), .B(n104), .CI(
        C[922]), .S(S[922]), .CO(C[923]) );
  FA_13729 \FA_INST_0[1].FA_INST_1[411].FA_  ( .A(A[923]), .B(n103), .CI(
        C[923]), .S(S[923]), .CO(C[924]) );
  FA_13728 \FA_INST_0[1].FA_INST_1[412].FA_  ( .A(A[924]), .B(n102), .CI(
        C[924]), .S(S[924]), .CO(C[925]) );
  FA_13727 \FA_INST_0[1].FA_INST_1[413].FA_  ( .A(A[925]), .B(n101), .CI(
        C[925]), .S(S[925]), .CO(C[926]) );
  FA_13726 \FA_INST_0[1].FA_INST_1[414].FA_  ( .A(A[926]), .B(n100), .CI(
        C[926]), .S(S[926]), .CO(C[927]) );
  FA_13725 \FA_INST_0[1].FA_INST_1[415].FA_  ( .A(A[927]), .B(n99), .CI(C[927]), .S(S[927]), .CO(C[928]) );
  FA_13724 \FA_INST_0[1].FA_INST_1[416].FA_  ( .A(A[928]), .B(n98), .CI(C[928]), .S(S[928]), .CO(C[929]) );
  FA_13723 \FA_INST_0[1].FA_INST_1[417].FA_  ( .A(A[929]), .B(n97), .CI(C[929]), .S(S[929]), .CO(C[930]) );
  FA_13722 \FA_INST_0[1].FA_INST_1[418].FA_  ( .A(A[930]), .B(n96), .CI(C[930]), .S(S[930]), .CO(C[931]) );
  FA_13721 \FA_INST_0[1].FA_INST_1[419].FA_  ( .A(A[931]), .B(n95), .CI(C[931]), .S(S[931]), .CO(C[932]) );
  FA_13720 \FA_INST_0[1].FA_INST_1[420].FA_  ( .A(A[932]), .B(n94), .CI(C[932]), .S(S[932]), .CO(C[933]) );
  FA_13719 \FA_INST_0[1].FA_INST_1[421].FA_  ( .A(A[933]), .B(n93), .CI(C[933]), .S(S[933]), .CO(C[934]) );
  FA_13718 \FA_INST_0[1].FA_INST_1[422].FA_  ( .A(A[934]), .B(n92), .CI(C[934]), .S(S[934]), .CO(C[935]) );
  FA_13717 \FA_INST_0[1].FA_INST_1[423].FA_  ( .A(A[935]), .B(n91), .CI(C[935]), .S(S[935]), .CO(C[936]) );
  FA_13716 \FA_INST_0[1].FA_INST_1[424].FA_  ( .A(A[936]), .B(n90), .CI(C[936]), .S(S[936]), .CO(C[937]) );
  FA_13715 \FA_INST_0[1].FA_INST_1[425].FA_  ( .A(A[937]), .B(n89), .CI(C[937]), .S(S[937]), .CO(C[938]) );
  FA_13714 \FA_INST_0[1].FA_INST_1[426].FA_  ( .A(A[938]), .B(n88), .CI(C[938]), .S(S[938]), .CO(C[939]) );
  FA_13713 \FA_INST_0[1].FA_INST_1[427].FA_  ( .A(A[939]), .B(n87), .CI(C[939]), .S(S[939]), .CO(C[940]) );
  FA_13712 \FA_INST_0[1].FA_INST_1[428].FA_  ( .A(A[940]), .B(n86), .CI(C[940]), .S(S[940]), .CO(C[941]) );
  FA_13711 \FA_INST_0[1].FA_INST_1[429].FA_  ( .A(A[941]), .B(n85), .CI(C[941]), .S(S[941]), .CO(C[942]) );
  FA_13710 \FA_INST_0[1].FA_INST_1[430].FA_  ( .A(A[942]), .B(n84), .CI(C[942]), .S(S[942]), .CO(C[943]) );
  FA_13709 \FA_INST_0[1].FA_INST_1[431].FA_  ( .A(A[943]), .B(n83), .CI(C[943]), .S(S[943]), .CO(C[944]) );
  FA_13708 \FA_INST_0[1].FA_INST_1[432].FA_  ( .A(A[944]), .B(n82), .CI(C[944]), .S(S[944]), .CO(C[945]) );
  FA_13707 \FA_INST_0[1].FA_INST_1[433].FA_  ( .A(A[945]), .B(n81), .CI(C[945]), .S(S[945]), .CO(C[946]) );
  FA_13706 \FA_INST_0[1].FA_INST_1[434].FA_  ( .A(A[946]), .B(n80), .CI(C[946]), .S(S[946]), .CO(C[947]) );
  FA_13705 \FA_INST_0[1].FA_INST_1[435].FA_  ( .A(A[947]), .B(n79), .CI(C[947]), .S(S[947]), .CO(C[948]) );
  FA_13704 \FA_INST_0[1].FA_INST_1[436].FA_  ( .A(A[948]), .B(n78), .CI(C[948]), .S(S[948]), .CO(C[949]) );
  FA_13703 \FA_INST_0[1].FA_INST_1[437].FA_  ( .A(A[949]), .B(n77), .CI(C[949]), .S(S[949]), .CO(C[950]) );
  FA_13702 \FA_INST_0[1].FA_INST_1[438].FA_  ( .A(A[950]), .B(n76), .CI(C[950]), .S(S[950]), .CO(C[951]) );
  FA_13701 \FA_INST_0[1].FA_INST_1[439].FA_  ( .A(A[951]), .B(n75), .CI(C[951]), .S(S[951]), .CO(C[952]) );
  FA_13700 \FA_INST_0[1].FA_INST_1[440].FA_  ( .A(A[952]), .B(n74), .CI(C[952]), .S(S[952]), .CO(C[953]) );
  FA_13699 \FA_INST_0[1].FA_INST_1[441].FA_  ( .A(A[953]), .B(n73), .CI(C[953]), .S(S[953]), .CO(C[954]) );
  FA_13698 \FA_INST_0[1].FA_INST_1[442].FA_  ( .A(A[954]), .B(n72), .CI(C[954]), .S(S[954]), .CO(C[955]) );
  FA_13697 \FA_INST_0[1].FA_INST_1[443].FA_  ( .A(A[955]), .B(n71), .CI(C[955]), .S(S[955]), .CO(C[956]) );
  FA_13696 \FA_INST_0[1].FA_INST_1[444].FA_  ( .A(A[956]), .B(n70), .CI(C[956]), .S(S[956]), .CO(C[957]) );
  FA_13695 \FA_INST_0[1].FA_INST_1[445].FA_  ( .A(A[957]), .B(n69), .CI(C[957]), .S(S[957]), .CO(C[958]) );
  FA_13694 \FA_INST_0[1].FA_INST_1[446].FA_  ( .A(A[958]), .B(n68), .CI(C[958]), .S(S[958]), .CO(C[959]) );
  FA_13693 \FA_INST_0[1].FA_INST_1[447].FA_  ( .A(A[959]), .B(n67), .CI(C[959]), .S(S[959]), .CO(C[960]) );
  FA_13692 \FA_INST_0[1].FA_INST_1[448].FA_  ( .A(A[960]), .B(n66), .CI(C[960]), .S(S[960]), .CO(C[961]) );
  FA_13691 \FA_INST_0[1].FA_INST_1[449].FA_  ( .A(A[961]), .B(n65), .CI(C[961]), .S(S[961]), .CO(C[962]) );
  FA_13690 \FA_INST_0[1].FA_INST_1[450].FA_  ( .A(A[962]), .B(n64), .CI(C[962]), .S(S[962]), .CO(C[963]) );
  FA_13689 \FA_INST_0[1].FA_INST_1[451].FA_  ( .A(A[963]), .B(n63), .CI(C[963]), .S(S[963]), .CO(C[964]) );
  FA_13688 \FA_INST_0[1].FA_INST_1[452].FA_  ( .A(A[964]), .B(n62), .CI(C[964]), .S(S[964]), .CO(C[965]) );
  FA_13687 \FA_INST_0[1].FA_INST_1[453].FA_  ( .A(A[965]), .B(n61), .CI(C[965]), .S(S[965]), .CO(C[966]) );
  FA_13686 \FA_INST_0[1].FA_INST_1[454].FA_  ( .A(A[966]), .B(n60), .CI(C[966]), .S(S[966]), .CO(C[967]) );
  FA_13685 \FA_INST_0[1].FA_INST_1[455].FA_  ( .A(A[967]), .B(n59), .CI(C[967]), .S(S[967]), .CO(C[968]) );
  FA_13684 \FA_INST_0[1].FA_INST_1[456].FA_  ( .A(A[968]), .B(n58), .CI(C[968]), .S(S[968]), .CO(C[969]) );
  FA_13683 \FA_INST_0[1].FA_INST_1[457].FA_  ( .A(A[969]), .B(n57), .CI(C[969]), .S(S[969]), .CO(C[970]) );
  FA_13682 \FA_INST_0[1].FA_INST_1[458].FA_  ( .A(A[970]), .B(n56), .CI(C[970]), .S(S[970]), .CO(C[971]) );
  FA_13681 \FA_INST_0[1].FA_INST_1[459].FA_  ( .A(A[971]), .B(n55), .CI(C[971]), .S(S[971]), .CO(C[972]) );
  FA_13680 \FA_INST_0[1].FA_INST_1[460].FA_  ( .A(A[972]), .B(n54), .CI(C[972]), .S(S[972]), .CO(C[973]) );
  FA_13679 \FA_INST_0[1].FA_INST_1[461].FA_  ( .A(A[973]), .B(n53), .CI(C[973]), .S(S[973]), .CO(C[974]) );
  FA_13678 \FA_INST_0[1].FA_INST_1[462].FA_  ( .A(A[974]), .B(n52), .CI(C[974]), .S(S[974]), .CO(C[975]) );
  FA_13677 \FA_INST_0[1].FA_INST_1[463].FA_  ( .A(A[975]), .B(n51), .CI(C[975]), .S(S[975]), .CO(C[976]) );
  FA_13676 \FA_INST_0[1].FA_INST_1[464].FA_  ( .A(A[976]), .B(n50), .CI(C[976]), .S(S[976]), .CO(C[977]) );
  FA_13675 \FA_INST_0[1].FA_INST_1[465].FA_  ( .A(A[977]), .B(n49), .CI(C[977]), .S(S[977]), .CO(C[978]) );
  FA_13674 \FA_INST_0[1].FA_INST_1[466].FA_  ( .A(A[978]), .B(n48), .CI(C[978]), .S(S[978]), .CO(C[979]) );
  FA_13673 \FA_INST_0[1].FA_INST_1[467].FA_  ( .A(A[979]), .B(n47), .CI(C[979]), .S(S[979]), .CO(C[980]) );
  FA_13672 \FA_INST_0[1].FA_INST_1[468].FA_  ( .A(A[980]), .B(n46), .CI(C[980]), .S(S[980]), .CO(C[981]) );
  FA_13671 \FA_INST_0[1].FA_INST_1[469].FA_  ( .A(A[981]), .B(n45), .CI(C[981]), .S(S[981]), .CO(C[982]) );
  FA_13670 \FA_INST_0[1].FA_INST_1[470].FA_  ( .A(A[982]), .B(n44), .CI(C[982]), .S(S[982]), .CO(C[983]) );
  FA_13669 \FA_INST_0[1].FA_INST_1[471].FA_  ( .A(A[983]), .B(n43), .CI(C[983]), .S(S[983]), .CO(C[984]) );
  FA_13668 \FA_INST_0[1].FA_INST_1[472].FA_  ( .A(A[984]), .B(n42), .CI(C[984]), .S(S[984]), .CO(C[985]) );
  FA_13667 \FA_INST_0[1].FA_INST_1[473].FA_  ( .A(A[985]), .B(n41), .CI(C[985]), .S(S[985]), .CO(C[986]) );
  FA_13666 \FA_INST_0[1].FA_INST_1[474].FA_  ( .A(A[986]), .B(n40), .CI(C[986]), .S(S[986]), .CO(C[987]) );
  FA_13665 \FA_INST_0[1].FA_INST_1[475].FA_  ( .A(A[987]), .B(n39), .CI(C[987]), .S(S[987]), .CO(C[988]) );
  FA_13664 \FA_INST_0[1].FA_INST_1[476].FA_  ( .A(A[988]), .B(n38), .CI(C[988]), .S(S[988]), .CO(C[989]) );
  FA_13663 \FA_INST_0[1].FA_INST_1[477].FA_  ( .A(A[989]), .B(n37), .CI(C[989]), .S(S[989]), .CO(C[990]) );
  FA_13662 \FA_INST_0[1].FA_INST_1[478].FA_  ( .A(A[990]), .B(n36), .CI(C[990]), .S(S[990]), .CO(C[991]) );
  FA_13661 \FA_INST_0[1].FA_INST_1[479].FA_  ( .A(A[991]), .B(n35), .CI(C[991]), .S(S[991]), .CO(C[992]) );
  FA_13660 \FA_INST_0[1].FA_INST_1[480].FA_  ( .A(A[992]), .B(n34), .CI(C[992]), .S(S[992]), .CO(C[993]) );
  FA_13659 \FA_INST_0[1].FA_INST_1[481].FA_  ( .A(A[993]), .B(n33), .CI(C[993]), .S(S[993]), .CO(C[994]) );
  FA_13658 \FA_INST_0[1].FA_INST_1[482].FA_  ( .A(A[994]), .B(n32), .CI(C[994]), .S(S[994]), .CO(C[995]) );
  FA_13657 \FA_INST_0[1].FA_INST_1[483].FA_  ( .A(A[995]), .B(n31), .CI(C[995]), .S(S[995]), .CO(C[996]) );
  FA_13656 \FA_INST_0[1].FA_INST_1[484].FA_  ( .A(A[996]), .B(n30), .CI(C[996]), .S(S[996]), .CO(C[997]) );
  FA_13655 \FA_INST_0[1].FA_INST_1[485].FA_  ( .A(A[997]), .B(n29), .CI(C[997]), .S(S[997]), .CO(C[998]) );
  FA_13654 \FA_INST_0[1].FA_INST_1[486].FA_  ( .A(A[998]), .B(n28), .CI(C[998]), .S(S[998]), .CO(C[999]) );
  FA_13653 \FA_INST_0[1].FA_INST_1[487].FA_  ( .A(A[999]), .B(n27), .CI(C[999]), .S(S[999]), .CO(C[1000]) );
  FA_13652 \FA_INST_0[1].FA_INST_1[488].FA_  ( .A(A[1000]), .B(n26), .CI(
        C[1000]), .S(S[1000]), .CO(C[1001]) );
  FA_13651 \FA_INST_0[1].FA_INST_1[489].FA_  ( .A(A[1001]), .B(n25), .CI(
        C[1001]), .S(S[1001]), .CO(C[1002]) );
  FA_13650 \FA_INST_0[1].FA_INST_1[490].FA_  ( .A(A[1002]), .B(n24), .CI(
        C[1002]), .S(S[1002]), .CO(C[1003]) );
  FA_13649 \FA_INST_0[1].FA_INST_1[491].FA_  ( .A(A[1003]), .B(n23), .CI(
        C[1003]), .S(S[1003]), .CO(C[1004]) );
  FA_13648 \FA_INST_0[1].FA_INST_1[492].FA_  ( .A(A[1004]), .B(n22), .CI(
        C[1004]), .S(S[1004]), .CO(C[1005]) );
  FA_13647 \FA_INST_0[1].FA_INST_1[493].FA_  ( .A(A[1005]), .B(n21), .CI(
        C[1005]), .S(S[1005]), .CO(C[1006]) );
  FA_13646 \FA_INST_0[1].FA_INST_1[494].FA_  ( .A(A[1006]), .B(n20), .CI(
        C[1006]), .S(S[1006]), .CO(C[1007]) );
  FA_13645 \FA_INST_0[1].FA_INST_1[495].FA_  ( .A(A[1007]), .B(n19), .CI(
        C[1007]), .S(S[1007]), .CO(C[1008]) );
  FA_13644 \FA_INST_0[1].FA_INST_1[496].FA_  ( .A(A[1008]), .B(n18), .CI(
        C[1008]), .S(S[1008]), .CO(C[1009]) );
  FA_13643 \FA_INST_0[1].FA_INST_1[497].FA_  ( .A(A[1009]), .B(n17), .CI(
        C[1009]), .S(S[1009]), .CO(C[1010]) );
  FA_13642 \FA_INST_0[1].FA_INST_1[498].FA_  ( .A(A[1010]), .B(n16), .CI(
        C[1010]), .S(S[1010]), .CO(C[1011]) );
  FA_13641 \FA_INST_0[1].FA_INST_1[499].FA_  ( .A(A[1011]), .B(n15), .CI(
        C[1011]), .S(S[1011]), .CO(C[1012]) );
  FA_13640 \FA_INST_0[1].FA_INST_1[500].FA_  ( .A(A[1012]), .B(n14), .CI(
        C[1012]), .S(S[1012]), .CO(C[1013]) );
  FA_13639 \FA_INST_0[1].FA_INST_1[501].FA_  ( .A(A[1013]), .B(n13), .CI(
        C[1013]), .S(S[1013]), .CO(C[1014]) );
  FA_13638 \FA_INST_0[1].FA_INST_1[502].FA_  ( .A(A[1014]), .B(n12), .CI(
        C[1014]), .S(S[1014]), .CO(C[1015]) );
  FA_13637 \FA_INST_0[1].FA_INST_1[503].FA_  ( .A(A[1015]), .B(n11), .CI(
        C[1015]), .S(S[1015]), .CO(C[1016]) );
  FA_13636 \FA_INST_0[1].FA_INST_1[504].FA_  ( .A(A[1016]), .B(n10), .CI(
        C[1016]), .S(S[1016]), .CO(C[1017]) );
  FA_13635 \FA_INST_0[1].FA_INST_1[505].FA_  ( .A(A[1017]), .B(n9), .CI(
        C[1017]), .S(S[1017]), .CO(C[1018]) );
  FA_13634 \FA_INST_0[1].FA_INST_1[506].FA_  ( .A(A[1018]), .B(n8), .CI(
        C[1018]), .S(S[1018]), .CO(C[1019]) );
  FA_13633 \FA_INST_0[1].FA_INST_1[507].FA_  ( .A(A[1019]), .B(n7), .CI(
        C[1019]), .S(S[1019]), .CO(C[1020]) );
  FA_13632 \FA_INST_0[1].FA_INST_1[508].FA_  ( .A(A[1020]), .B(n6), .CI(
        C[1020]), .S(S[1020]), .CO(C[1021]) );
  FA_13631 \FA_INST_0[1].FA_INST_1[509].FA_  ( .A(A[1021]), .B(n5), .CI(
        C[1021]), .S(S[1021]), .CO(C[1022]) );
  FA_13630 \FA_INST_0[1].FA_INST_1[510].FA_  ( .A(A[1022]), .B(n4), .CI(
        C[1022]), .S(S[1022]), .CO(C[1023]) );
  FA_13629 \FA_INST_0[1].FA_INST_1[511].FA_  ( .A(A[1023]), .B(n3), .CI(
        C[1023]), .S(S[1023]), .CO(C[1024]) );
  FA_13628 \FA_INST_1[1024].FA_  ( .A(A[1024]), .B(1'b1), .CI(C[1024]), .S(
        S[1024]), .CO(C[1025]) );
  FA_13627 \FA_INST_1[1025].FA_  ( .A(A[1025]), .B(1'b1), .CI(C[1025]), .S(
        S[1025]) );
  IV U2 ( .A(B[27]), .Z(n999) );
  IV U3 ( .A(B[28]), .Z(n998) );
  IV U4 ( .A(B[29]), .Z(n997) );
  IV U5 ( .A(B[30]), .Z(n996) );
  IV U6 ( .A(B[31]), .Z(n995) );
  IV U7 ( .A(B[32]), .Z(n994) );
  IV U8 ( .A(B[33]), .Z(n993) );
  IV U9 ( .A(B[34]), .Z(n992) );
  IV U10 ( .A(B[35]), .Z(n991) );
  IV U11 ( .A(B[36]), .Z(n990) );
  IV U12 ( .A(B[927]), .Z(n99) );
  IV U13 ( .A(B[37]), .Z(n989) );
  IV U14 ( .A(B[38]), .Z(n988) );
  IV U15 ( .A(B[39]), .Z(n987) );
  IV U16 ( .A(B[40]), .Z(n986) );
  IV U17 ( .A(B[41]), .Z(n985) );
  IV U18 ( .A(B[42]), .Z(n984) );
  IV U19 ( .A(B[43]), .Z(n983) );
  IV U20 ( .A(B[44]), .Z(n982) );
  IV U21 ( .A(B[45]), .Z(n981) );
  IV U22 ( .A(B[46]), .Z(n980) );
  IV U23 ( .A(B[928]), .Z(n98) );
  IV U24 ( .A(B[47]), .Z(n979) );
  IV U25 ( .A(B[48]), .Z(n978) );
  IV U26 ( .A(B[49]), .Z(n977) );
  IV U27 ( .A(B[50]), .Z(n976) );
  IV U28 ( .A(B[51]), .Z(n975) );
  IV U29 ( .A(B[52]), .Z(n974) );
  IV U30 ( .A(B[53]), .Z(n973) );
  IV U31 ( .A(B[54]), .Z(n972) );
  IV U32 ( .A(B[55]), .Z(n971) );
  IV U33 ( .A(B[56]), .Z(n970) );
  IV U34 ( .A(B[929]), .Z(n97) );
  IV U35 ( .A(B[57]), .Z(n969) );
  IV U36 ( .A(B[58]), .Z(n968) );
  IV U37 ( .A(B[59]), .Z(n967) );
  IV U38 ( .A(B[60]), .Z(n966) );
  IV U39 ( .A(B[61]), .Z(n965) );
  IV U40 ( .A(B[62]), .Z(n964) );
  IV U41 ( .A(B[63]), .Z(n963) );
  IV U42 ( .A(B[64]), .Z(n962) );
  IV U43 ( .A(B[65]), .Z(n961) );
  IV U44 ( .A(B[66]), .Z(n960) );
  IV U45 ( .A(B[930]), .Z(n96) );
  IV U46 ( .A(B[67]), .Z(n959) );
  IV U47 ( .A(B[68]), .Z(n958) );
  IV U48 ( .A(B[69]), .Z(n957) );
  IV U49 ( .A(B[70]), .Z(n956) );
  IV U50 ( .A(B[71]), .Z(n955) );
  IV U51 ( .A(B[72]), .Z(n954) );
  IV U52 ( .A(B[73]), .Z(n953) );
  IV U53 ( .A(B[74]), .Z(n952) );
  IV U54 ( .A(B[75]), .Z(n951) );
  IV U55 ( .A(B[76]), .Z(n950) );
  IV U56 ( .A(B[931]), .Z(n95) );
  IV U57 ( .A(B[77]), .Z(n949) );
  IV U58 ( .A(B[78]), .Z(n948) );
  IV U59 ( .A(B[79]), .Z(n947) );
  IV U60 ( .A(B[80]), .Z(n946) );
  IV U61 ( .A(B[81]), .Z(n945) );
  IV U62 ( .A(B[82]), .Z(n944) );
  IV U63 ( .A(B[83]), .Z(n943) );
  IV U64 ( .A(B[84]), .Z(n942) );
  IV U65 ( .A(B[85]), .Z(n941) );
  IV U66 ( .A(B[86]), .Z(n940) );
  IV U67 ( .A(B[932]), .Z(n94) );
  IV U68 ( .A(B[87]), .Z(n939) );
  IV U69 ( .A(B[88]), .Z(n938) );
  IV U70 ( .A(B[89]), .Z(n937) );
  IV U71 ( .A(B[90]), .Z(n936) );
  IV U72 ( .A(B[91]), .Z(n935) );
  IV U73 ( .A(B[92]), .Z(n934) );
  IV U74 ( .A(B[93]), .Z(n933) );
  IV U75 ( .A(B[94]), .Z(n932) );
  IV U76 ( .A(B[95]), .Z(n931) );
  IV U77 ( .A(B[96]), .Z(n930) );
  IV U78 ( .A(B[933]), .Z(n93) );
  IV U79 ( .A(B[97]), .Z(n929) );
  IV U80 ( .A(B[98]), .Z(n928) );
  IV U81 ( .A(B[99]), .Z(n927) );
  IV U82 ( .A(B[100]), .Z(n926) );
  IV U83 ( .A(B[101]), .Z(n925) );
  IV U84 ( .A(B[102]), .Z(n924) );
  IV U85 ( .A(B[103]), .Z(n923) );
  IV U86 ( .A(B[104]), .Z(n922) );
  IV U87 ( .A(B[105]), .Z(n921) );
  IV U88 ( .A(B[106]), .Z(n920) );
  IV U89 ( .A(B[934]), .Z(n92) );
  IV U90 ( .A(B[107]), .Z(n919) );
  IV U91 ( .A(B[108]), .Z(n918) );
  IV U92 ( .A(B[109]), .Z(n917) );
  IV U93 ( .A(B[110]), .Z(n916) );
  IV U94 ( .A(B[111]), .Z(n915) );
  IV U95 ( .A(B[112]), .Z(n914) );
  IV U96 ( .A(B[113]), .Z(n913) );
  IV U97 ( .A(B[114]), .Z(n912) );
  IV U98 ( .A(B[115]), .Z(n911) );
  IV U99 ( .A(B[116]), .Z(n910) );
  IV U100 ( .A(B[935]), .Z(n91) );
  IV U101 ( .A(B[117]), .Z(n909) );
  IV U102 ( .A(B[118]), .Z(n908) );
  IV U103 ( .A(B[119]), .Z(n907) );
  IV U104 ( .A(B[120]), .Z(n906) );
  IV U105 ( .A(B[121]), .Z(n905) );
  IV U106 ( .A(B[122]), .Z(n904) );
  IV U107 ( .A(B[123]), .Z(n903) );
  IV U108 ( .A(B[124]), .Z(n902) );
  IV U109 ( .A(B[125]), .Z(n901) );
  IV U110 ( .A(B[126]), .Z(n900) );
  IV U111 ( .A(B[936]), .Z(n90) );
  IV U112 ( .A(B[1017]), .Z(n9) );
  IV U113 ( .A(B[127]), .Z(n899) );
  IV U114 ( .A(B[128]), .Z(n898) );
  IV U115 ( .A(B[129]), .Z(n897) );
  IV U116 ( .A(B[130]), .Z(n896) );
  IV U117 ( .A(B[131]), .Z(n895) );
  IV U118 ( .A(B[132]), .Z(n894) );
  IV U119 ( .A(B[133]), .Z(n893) );
  IV U120 ( .A(B[134]), .Z(n892) );
  IV U121 ( .A(B[135]), .Z(n891) );
  IV U122 ( .A(B[136]), .Z(n890) );
  IV U123 ( .A(B[937]), .Z(n89) );
  IV U124 ( .A(B[137]), .Z(n889) );
  IV U125 ( .A(B[138]), .Z(n888) );
  IV U126 ( .A(B[139]), .Z(n887) );
  IV U127 ( .A(B[140]), .Z(n886) );
  IV U128 ( .A(B[141]), .Z(n885) );
  IV U129 ( .A(B[142]), .Z(n884) );
  IV U130 ( .A(B[143]), .Z(n883) );
  IV U131 ( .A(B[144]), .Z(n882) );
  IV U132 ( .A(B[145]), .Z(n881) );
  IV U133 ( .A(B[146]), .Z(n880) );
  IV U134 ( .A(B[938]), .Z(n88) );
  IV U135 ( .A(B[147]), .Z(n879) );
  IV U136 ( .A(B[148]), .Z(n878) );
  IV U137 ( .A(B[149]), .Z(n877) );
  IV U138 ( .A(B[150]), .Z(n876) );
  IV U139 ( .A(B[151]), .Z(n875) );
  IV U140 ( .A(B[152]), .Z(n874) );
  IV U141 ( .A(B[153]), .Z(n873) );
  IV U142 ( .A(B[154]), .Z(n872) );
  IV U143 ( .A(B[155]), .Z(n871) );
  IV U144 ( .A(B[156]), .Z(n870) );
  IV U145 ( .A(B[939]), .Z(n87) );
  IV U146 ( .A(B[157]), .Z(n869) );
  IV U147 ( .A(B[158]), .Z(n868) );
  IV U148 ( .A(B[159]), .Z(n867) );
  IV U149 ( .A(B[160]), .Z(n866) );
  IV U150 ( .A(B[161]), .Z(n865) );
  IV U151 ( .A(B[162]), .Z(n864) );
  IV U152 ( .A(B[163]), .Z(n863) );
  IV U153 ( .A(B[164]), .Z(n862) );
  IV U154 ( .A(B[165]), .Z(n861) );
  IV U155 ( .A(B[166]), .Z(n860) );
  IV U156 ( .A(B[940]), .Z(n86) );
  IV U157 ( .A(B[167]), .Z(n859) );
  IV U158 ( .A(B[168]), .Z(n858) );
  IV U159 ( .A(B[169]), .Z(n857) );
  IV U160 ( .A(B[170]), .Z(n856) );
  IV U161 ( .A(B[171]), .Z(n855) );
  IV U162 ( .A(B[172]), .Z(n854) );
  IV U163 ( .A(B[173]), .Z(n853) );
  IV U164 ( .A(B[174]), .Z(n852) );
  IV U165 ( .A(B[175]), .Z(n851) );
  IV U166 ( .A(B[176]), .Z(n850) );
  IV U167 ( .A(B[941]), .Z(n85) );
  IV U168 ( .A(B[177]), .Z(n849) );
  IV U169 ( .A(B[178]), .Z(n848) );
  IV U170 ( .A(B[179]), .Z(n847) );
  IV U171 ( .A(B[180]), .Z(n846) );
  IV U172 ( .A(B[181]), .Z(n845) );
  IV U173 ( .A(B[182]), .Z(n844) );
  IV U174 ( .A(B[183]), .Z(n843) );
  IV U175 ( .A(B[184]), .Z(n842) );
  IV U176 ( .A(B[185]), .Z(n841) );
  IV U177 ( .A(B[186]), .Z(n840) );
  IV U178 ( .A(B[942]), .Z(n84) );
  IV U179 ( .A(B[187]), .Z(n839) );
  IV U180 ( .A(B[188]), .Z(n838) );
  IV U181 ( .A(B[189]), .Z(n837) );
  IV U182 ( .A(B[190]), .Z(n836) );
  IV U183 ( .A(B[191]), .Z(n835) );
  IV U184 ( .A(B[192]), .Z(n834) );
  IV U185 ( .A(B[193]), .Z(n833) );
  IV U186 ( .A(B[194]), .Z(n832) );
  IV U187 ( .A(B[195]), .Z(n831) );
  IV U188 ( .A(B[196]), .Z(n830) );
  IV U189 ( .A(B[943]), .Z(n83) );
  IV U190 ( .A(B[197]), .Z(n829) );
  IV U191 ( .A(B[198]), .Z(n828) );
  IV U192 ( .A(B[199]), .Z(n827) );
  IV U193 ( .A(B[200]), .Z(n826) );
  IV U194 ( .A(B[201]), .Z(n825) );
  IV U195 ( .A(B[202]), .Z(n824) );
  IV U196 ( .A(B[203]), .Z(n823) );
  IV U197 ( .A(B[204]), .Z(n822) );
  IV U198 ( .A(B[205]), .Z(n821) );
  IV U199 ( .A(B[206]), .Z(n820) );
  IV U200 ( .A(B[944]), .Z(n82) );
  IV U201 ( .A(B[207]), .Z(n819) );
  IV U202 ( .A(B[208]), .Z(n818) );
  IV U203 ( .A(B[209]), .Z(n817) );
  IV U204 ( .A(B[210]), .Z(n816) );
  IV U205 ( .A(B[211]), .Z(n815) );
  IV U206 ( .A(B[212]), .Z(n814) );
  IV U207 ( .A(B[213]), .Z(n813) );
  IV U208 ( .A(B[214]), .Z(n812) );
  IV U209 ( .A(B[215]), .Z(n811) );
  IV U210 ( .A(B[216]), .Z(n810) );
  IV U211 ( .A(B[945]), .Z(n81) );
  IV U212 ( .A(B[217]), .Z(n809) );
  IV U213 ( .A(B[218]), .Z(n808) );
  IV U214 ( .A(B[219]), .Z(n807) );
  IV U215 ( .A(B[220]), .Z(n806) );
  IV U216 ( .A(B[221]), .Z(n805) );
  IV U217 ( .A(B[222]), .Z(n804) );
  IV U218 ( .A(B[223]), .Z(n803) );
  IV U219 ( .A(B[224]), .Z(n802) );
  IV U220 ( .A(B[225]), .Z(n801) );
  IV U221 ( .A(B[226]), .Z(n800) );
  IV U222 ( .A(B[946]), .Z(n80) );
  IV U223 ( .A(B[1018]), .Z(n8) );
  IV U224 ( .A(B[227]), .Z(n799) );
  IV U225 ( .A(B[228]), .Z(n798) );
  IV U226 ( .A(B[229]), .Z(n797) );
  IV U227 ( .A(B[230]), .Z(n796) );
  IV U228 ( .A(B[231]), .Z(n795) );
  IV U229 ( .A(B[232]), .Z(n794) );
  IV U230 ( .A(B[233]), .Z(n793) );
  IV U231 ( .A(B[234]), .Z(n792) );
  IV U232 ( .A(B[235]), .Z(n791) );
  IV U233 ( .A(B[236]), .Z(n790) );
  IV U234 ( .A(B[947]), .Z(n79) );
  IV U235 ( .A(B[237]), .Z(n789) );
  IV U236 ( .A(B[238]), .Z(n788) );
  IV U237 ( .A(B[239]), .Z(n787) );
  IV U238 ( .A(B[240]), .Z(n786) );
  IV U239 ( .A(B[241]), .Z(n785) );
  IV U240 ( .A(B[242]), .Z(n784) );
  IV U241 ( .A(B[243]), .Z(n783) );
  IV U242 ( .A(B[244]), .Z(n782) );
  IV U243 ( .A(B[245]), .Z(n781) );
  IV U244 ( .A(B[246]), .Z(n780) );
  IV U245 ( .A(B[948]), .Z(n78) );
  IV U246 ( .A(B[247]), .Z(n779) );
  IV U247 ( .A(B[248]), .Z(n778) );
  IV U248 ( .A(B[249]), .Z(n777) );
  IV U249 ( .A(B[250]), .Z(n776) );
  IV U250 ( .A(B[251]), .Z(n775) );
  IV U251 ( .A(B[252]), .Z(n774) );
  IV U252 ( .A(B[253]), .Z(n773) );
  IV U253 ( .A(B[254]), .Z(n772) );
  IV U254 ( .A(B[255]), .Z(n771) );
  IV U255 ( .A(B[256]), .Z(n770) );
  IV U256 ( .A(B[949]), .Z(n77) );
  IV U257 ( .A(B[257]), .Z(n769) );
  IV U258 ( .A(B[258]), .Z(n768) );
  IV U259 ( .A(B[259]), .Z(n767) );
  IV U260 ( .A(B[260]), .Z(n766) );
  IV U261 ( .A(B[261]), .Z(n765) );
  IV U262 ( .A(B[262]), .Z(n764) );
  IV U263 ( .A(B[263]), .Z(n763) );
  IV U264 ( .A(B[264]), .Z(n762) );
  IV U265 ( .A(B[265]), .Z(n761) );
  IV U266 ( .A(B[266]), .Z(n760) );
  IV U267 ( .A(B[950]), .Z(n76) );
  IV U268 ( .A(B[267]), .Z(n759) );
  IV U269 ( .A(B[268]), .Z(n758) );
  IV U270 ( .A(B[269]), .Z(n757) );
  IV U271 ( .A(B[270]), .Z(n756) );
  IV U272 ( .A(B[271]), .Z(n755) );
  IV U273 ( .A(B[272]), .Z(n754) );
  IV U274 ( .A(B[273]), .Z(n753) );
  IV U275 ( .A(B[274]), .Z(n752) );
  IV U276 ( .A(B[275]), .Z(n751) );
  IV U277 ( .A(B[276]), .Z(n750) );
  IV U278 ( .A(B[951]), .Z(n75) );
  IV U279 ( .A(B[277]), .Z(n749) );
  IV U280 ( .A(B[278]), .Z(n748) );
  IV U281 ( .A(B[279]), .Z(n747) );
  IV U282 ( .A(B[280]), .Z(n746) );
  IV U283 ( .A(B[281]), .Z(n745) );
  IV U284 ( .A(B[282]), .Z(n744) );
  IV U285 ( .A(B[283]), .Z(n743) );
  IV U286 ( .A(B[284]), .Z(n742) );
  IV U287 ( .A(B[285]), .Z(n741) );
  IV U288 ( .A(B[286]), .Z(n740) );
  IV U289 ( .A(B[952]), .Z(n74) );
  IV U290 ( .A(B[287]), .Z(n739) );
  IV U291 ( .A(B[288]), .Z(n738) );
  IV U292 ( .A(B[289]), .Z(n737) );
  IV U293 ( .A(B[290]), .Z(n736) );
  IV U294 ( .A(B[291]), .Z(n735) );
  IV U295 ( .A(B[292]), .Z(n734) );
  IV U296 ( .A(B[293]), .Z(n733) );
  IV U297 ( .A(B[294]), .Z(n732) );
  IV U298 ( .A(B[295]), .Z(n731) );
  IV U299 ( .A(B[296]), .Z(n730) );
  IV U300 ( .A(B[953]), .Z(n73) );
  IV U301 ( .A(B[297]), .Z(n729) );
  IV U302 ( .A(B[298]), .Z(n728) );
  IV U303 ( .A(B[299]), .Z(n727) );
  IV U304 ( .A(B[300]), .Z(n726) );
  IV U305 ( .A(B[301]), .Z(n725) );
  IV U306 ( .A(B[302]), .Z(n724) );
  IV U307 ( .A(B[303]), .Z(n723) );
  IV U308 ( .A(B[304]), .Z(n722) );
  IV U309 ( .A(B[305]), .Z(n721) );
  IV U310 ( .A(B[306]), .Z(n720) );
  IV U311 ( .A(B[954]), .Z(n72) );
  IV U312 ( .A(B[307]), .Z(n719) );
  IV U313 ( .A(B[308]), .Z(n718) );
  IV U314 ( .A(B[309]), .Z(n717) );
  IV U315 ( .A(B[310]), .Z(n716) );
  IV U316 ( .A(B[311]), .Z(n715) );
  IV U317 ( .A(B[312]), .Z(n714) );
  IV U318 ( .A(B[313]), .Z(n713) );
  IV U319 ( .A(B[314]), .Z(n712) );
  IV U320 ( .A(B[315]), .Z(n711) );
  IV U321 ( .A(B[316]), .Z(n710) );
  IV U322 ( .A(B[955]), .Z(n71) );
  IV U323 ( .A(B[317]), .Z(n709) );
  IV U324 ( .A(B[318]), .Z(n708) );
  IV U325 ( .A(B[319]), .Z(n707) );
  IV U326 ( .A(B[320]), .Z(n706) );
  IV U327 ( .A(B[321]), .Z(n705) );
  IV U328 ( .A(B[322]), .Z(n704) );
  IV U329 ( .A(B[323]), .Z(n703) );
  IV U330 ( .A(B[324]), .Z(n702) );
  IV U331 ( .A(B[325]), .Z(n701) );
  IV U332 ( .A(B[326]), .Z(n700) );
  IV U333 ( .A(B[956]), .Z(n70) );
  IV U334 ( .A(B[1019]), .Z(n7) );
  IV U335 ( .A(B[327]), .Z(n699) );
  IV U336 ( .A(B[328]), .Z(n698) );
  IV U337 ( .A(B[329]), .Z(n697) );
  IV U338 ( .A(B[330]), .Z(n696) );
  IV U339 ( .A(B[331]), .Z(n695) );
  IV U340 ( .A(B[332]), .Z(n694) );
  IV U341 ( .A(B[333]), .Z(n693) );
  IV U342 ( .A(B[334]), .Z(n692) );
  IV U343 ( .A(B[335]), .Z(n691) );
  IV U344 ( .A(B[336]), .Z(n690) );
  IV U345 ( .A(B[957]), .Z(n69) );
  IV U346 ( .A(B[337]), .Z(n689) );
  IV U347 ( .A(B[338]), .Z(n688) );
  IV U348 ( .A(B[339]), .Z(n687) );
  IV U349 ( .A(B[340]), .Z(n686) );
  IV U350 ( .A(B[341]), .Z(n685) );
  IV U351 ( .A(B[342]), .Z(n684) );
  IV U352 ( .A(B[343]), .Z(n683) );
  IV U353 ( .A(B[344]), .Z(n682) );
  IV U354 ( .A(B[345]), .Z(n681) );
  IV U355 ( .A(B[346]), .Z(n680) );
  IV U356 ( .A(B[958]), .Z(n68) );
  IV U357 ( .A(B[347]), .Z(n679) );
  IV U358 ( .A(B[348]), .Z(n678) );
  IV U359 ( .A(B[349]), .Z(n677) );
  IV U360 ( .A(B[350]), .Z(n676) );
  IV U361 ( .A(B[351]), .Z(n675) );
  IV U362 ( .A(B[352]), .Z(n674) );
  IV U363 ( .A(B[353]), .Z(n673) );
  IV U364 ( .A(B[354]), .Z(n672) );
  IV U365 ( .A(B[355]), .Z(n671) );
  IV U366 ( .A(B[356]), .Z(n670) );
  IV U367 ( .A(B[959]), .Z(n67) );
  IV U368 ( .A(B[357]), .Z(n669) );
  IV U369 ( .A(B[358]), .Z(n668) );
  IV U370 ( .A(B[359]), .Z(n667) );
  IV U371 ( .A(B[360]), .Z(n666) );
  IV U372 ( .A(B[361]), .Z(n665) );
  IV U373 ( .A(B[362]), .Z(n664) );
  IV U374 ( .A(B[363]), .Z(n663) );
  IV U375 ( .A(B[364]), .Z(n662) );
  IV U376 ( .A(B[365]), .Z(n661) );
  IV U377 ( .A(B[366]), .Z(n660) );
  IV U378 ( .A(B[960]), .Z(n66) );
  IV U379 ( .A(B[367]), .Z(n659) );
  IV U380 ( .A(B[368]), .Z(n658) );
  IV U381 ( .A(B[369]), .Z(n657) );
  IV U382 ( .A(B[370]), .Z(n656) );
  IV U383 ( .A(B[371]), .Z(n655) );
  IV U384 ( .A(B[372]), .Z(n654) );
  IV U385 ( .A(B[373]), .Z(n653) );
  IV U386 ( .A(B[374]), .Z(n652) );
  IV U387 ( .A(B[375]), .Z(n651) );
  IV U388 ( .A(B[376]), .Z(n650) );
  IV U389 ( .A(B[961]), .Z(n65) );
  IV U390 ( .A(B[377]), .Z(n649) );
  IV U391 ( .A(B[378]), .Z(n648) );
  IV U392 ( .A(B[379]), .Z(n647) );
  IV U393 ( .A(B[380]), .Z(n646) );
  IV U394 ( .A(B[381]), .Z(n645) );
  IV U395 ( .A(B[382]), .Z(n644) );
  IV U396 ( .A(B[383]), .Z(n643) );
  IV U397 ( .A(B[384]), .Z(n642) );
  IV U398 ( .A(B[385]), .Z(n641) );
  IV U399 ( .A(B[386]), .Z(n640) );
  IV U400 ( .A(B[962]), .Z(n64) );
  IV U401 ( .A(B[387]), .Z(n639) );
  IV U402 ( .A(B[388]), .Z(n638) );
  IV U403 ( .A(B[389]), .Z(n637) );
  IV U404 ( .A(B[390]), .Z(n636) );
  IV U405 ( .A(B[391]), .Z(n635) );
  IV U406 ( .A(B[392]), .Z(n634) );
  IV U407 ( .A(B[393]), .Z(n633) );
  IV U408 ( .A(B[394]), .Z(n632) );
  IV U409 ( .A(B[395]), .Z(n631) );
  IV U410 ( .A(B[396]), .Z(n630) );
  IV U411 ( .A(B[963]), .Z(n63) );
  IV U412 ( .A(B[397]), .Z(n629) );
  IV U413 ( .A(B[398]), .Z(n628) );
  IV U414 ( .A(B[399]), .Z(n627) );
  IV U415 ( .A(B[400]), .Z(n626) );
  IV U416 ( .A(B[401]), .Z(n625) );
  IV U417 ( .A(B[402]), .Z(n624) );
  IV U418 ( .A(B[403]), .Z(n623) );
  IV U419 ( .A(B[404]), .Z(n622) );
  IV U420 ( .A(B[405]), .Z(n621) );
  IV U421 ( .A(B[406]), .Z(n620) );
  IV U422 ( .A(B[964]), .Z(n62) );
  IV U423 ( .A(B[407]), .Z(n619) );
  IV U424 ( .A(B[408]), .Z(n618) );
  IV U425 ( .A(B[409]), .Z(n617) );
  IV U426 ( .A(B[410]), .Z(n616) );
  IV U427 ( .A(B[411]), .Z(n615) );
  IV U428 ( .A(B[412]), .Z(n614) );
  IV U429 ( .A(B[413]), .Z(n613) );
  IV U430 ( .A(B[414]), .Z(n612) );
  IV U431 ( .A(B[415]), .Z(n611) );
  IV U432 ( .A(B[416]), .Z(n610) );
  IV U433 ( .A(B[965]), .Z(n61) );
  IV U434 ( .A(B[417]), .Z(n609) );
  IV U435 ( .A(B[418]), .Z(n608) );
  IV U436 ( .A(B[419]), .Z(n607) );
  IV U437 ( .A(B[420]), .Z(n606) );
  IV U438 ( .A(B[421]), .Z(n605) );
  IV U439 ( .A(B[422]), .Z(n604) );
  IV U440 ( .A(B[423]), .Z(n603) );
  IV U441 ( .A(B[424]), .Z(n602) );
  IV U442 ( .A(B[425]), .Z(n601) );
  IV U443 ( .A(B[426]), .Z(n600) );
  IV U444 ( .A(B[966]), .Z(n60) );
  IV U445 ( .A(B[1020]), .Z(n6) );
  IV U446 ( .A(B[427]), .Z(n599) );
  IV U447 ( .A(B[428]), .Z(n598) );
  IV U448 ( .A(B[429]), .Z(n597) );
  IV U449 ( .A(B[430]), .Z(n596) );
  IV U450 ( .A(B[431]), .Z(n595) );
  IV U451 ( .A(B[432]), .Z(n594) );
  IV U452 ( .A(B[433]), .Z(n593) );
  IV U453 ( .A(B[434]), .Z(n592) );
  IV U454 ( .A(B[435]), .Z(n591) );
  IV U455 ( .A(B[436]), .Z(n590) );
  IV U456 ( .A(B[967]), .Z(n59) );
  IV U457 ( .A(B[437]), .Z(n589) );
  IV U458 ( .A(B[438]), .Z(n588) );
  IV U459 ( .A(B[439]), .Z(n587) );
  IV U460 ( .A(B[440]), .Z(n586) );
  IV U461 ( .A(B[441]), .Z(n585) );
  IV U462 ( .A(B[442]), .Z(n584) );
  IV U463 ( .A(B[443]), .Z(n583) );
  IV U464 ( .A(B[444]), .Z(n582) );
  IV U465 ( .A(B[445]), .Z(n581) );
  IV U466 ( .A(B[446]), .Z(n580) );
  IV U467 ( .A(B[968]), .Z(n58) );
  IV U468 ( .A(B[447]), .Z(n579) );
  IV U469 ( .A(B[448]), .Z(n578) );
  IV U470 ( .A(B[449]), .Z(n577) );
  IV U471 ( .A(B[450]), .Z(n576) );
  IV U472 ( .A(B[451]), .Z(n575) );
  IV U473 ( .A(B[452]), .Z(n574) );
  IV U474 ( .A(B[453]), .Z(n573) );
  IV U475 ( .A(B[454]), .Z(n572) );
  IV U476 ( .A(B[455]), .Z(n571) );
  IV U477 ( .A(B[456]), .Z(n570) );
  IV U478 ( .A(B[969]), .Z(n57) );
  IV U479 ( .A(B[457]), .Z(n569) );
  IV U480 ( .A(B[458]), .Z(n568) );
  IV U481 ( .A(B[459]), .Z(n567) );
  IV U482 ( .A(B[460]), .Z(n566) );
  IV U483 ( .A(B[461]), .Z(n565) );
  IV U484 ( .A(B[462]), .Z(n564) );
  IV U485 ( .A(B[463]), .Z(n563) );
  IV U486 ( .A(B[464]), .Z(n562) );
  IV U487 ( .A(B[465]), .Z(n561) );
  IV U488 ( .A(B[466]), .Z(n560) );
  IV U489 ( .A(B[970]), .Z(n56) );
  IV U490 ( .A(B[467]), .Z(n559) );
  IV U491 ( .A(B[468]), .Z(n558) );
  IV U492 ( .A(B[469]), .Z(n557) );
  IV U493 ( .A(B[470]), .Z(n556) );
  IV U494 ( .A(B[471]), .Z(n555) );
  IV U495 ( .A(B[472]), .Z(n554) );
  IV U496 ( .A(B[473]), .Z(n553) );
  IV U497 ( .A(B[474]), .Z(n552) );
  IV U498 ( .A(B[475]), .Z(n551) );
  IV U499 ( .A(B[476]), .Z(n550) );
  IV U500 ( .A(B[971]), .Z(n55) );
  IV U501 ( .A(B[477]), .Z(n549) );
  IV U502 ( .A(B[478]), .Z(n548) );
  IV U503 ( .A(B[479]), .Z(n547) );
  IV U504 ( .A(B[480]), .Z(n546) );
  IV U505 ( .A(B[481]), .Z(n545) );
  IV U506 ( .A(B[482]), .Z(n544) );
  IV U507 ( .A(B[483]), .Z(n543) );
  IV U508 ( .A(B[484]), .Z(n542) );
  IV U509 ( .A(B[485]), .Z(n541) );
  IV U510 ( .A(B[486]), .Z(n540) );
  IV U511 ( .A(B[972]), .Z(n54) );
  IV U512 ( .A(B[487]), .Z(n539) );
  IV U513 ( .A(B[488]), .Z(n538) );
  IV U514 ( .A(B[489]), .Z(n537) );
  IV U515 ( .A(B[490]), .Z(n536) );
  IV U516 ( .A(B[491]), .Z(n535) );
  IV U517 ( .A(B[492]), .Z(n534) );
  IV U518 ( .A(B[493]), .Z(n533) );
  IV U519 ( .A(B[494]), .Z(n532) );
  IV U520 ( .A(B[495]), .Z(n531) );
  IV U521 ( .A(B[496]), .Z(n530) );
  IV U522 ( .A(B[973]), .Z(n53) );
  IV U523 ( .A(B[497]), .Z(n529) );
  IV U524 ( .A(B[498]), .Z(n528) );
  IV U525 ( .A(B[499]), .Z(n527) );
  IV U526 ( .A(B[500]), .Z(n526) );
  IV U527 ( .A(B[501]), .Z(n525) );
  IV U528 ( .A(B[502]), .Z(n524) );
  IV U529 ( .A(B[503]), .Z(n523) );
  IV U530 ( .A(B[504]), .Z(n522) );
  IV U531 ( .A(B[505]), .Z(n521) );
  IV U532 ( .A(B[506]), .Z(n520) );
  IV U533 ( .A(B[974]), .Z(n52) );
  IV U534 ( .A(B[507]), .Z(n519) );
  IV U535 ( .A(B[508]), .Z(n518) );
  IV U536 ( .A(B[509]), .Z(n517) );
  IV U537 ( .A(B[510]), .Z(n516) );
  IV U538 ( .A(B[511]), .Z(n515) );
  IV U539 ( .A(B[512]), .Z(n514) );
  IV U540 ( .A(B[513]), .Z(n513) );
  IV U541 ( .A(B[514]), .Z(n512) );
  IV U542 ( .A(B[515]), .Z(n511) );
  IV U543 ( .A(B[516]), .Z(n510) );
  IV U544 ( .A(B[975]), .Z(n51) );
  IV U545 ( .A(B[517]), .Z(n509) );
  IV U546 ( .A(B[518]), .Z(n508) );
  IV U547 ( .A(B[519]), .Z(n507) );
  IV U548 ( .A(B[520]), .Z(n506) );
  IV U549 ( .A(B[521]), .Z(n505) );
  IV U550 ( .A(B[522]), .Z(n504) );
  IV U551 ( .A(B[523]), .Z(n503) );
  IV U552 ( .A(B[524]), .Z(n502) );
  IV U553 ( .A(B[525]), .Z(n501) );
  IV U554 ( .A(B[526]), .Z(n500) );
  IV U555 ( .A(B[976]), .Z(n50) );
  IV U556 ( .A(B[1021]), .Z(n5) );
  IV U557 ( .A(B[527]), .Z(n499) );
  IV U558 ( .A(B[528]), .Z(n498) );
  IV U559 ( .A(B[529]), .Z(n497) );
  IV U560 ( .A(B[530]), .Z(n496) );
  IV U561 ( .A(B[531]), .Z(n495) );
  IV U562 ( .A(B[532]), .Z(n494) );
  IV U563 ( .A(B[533]), .Z(n493) );
  IV U564 ( .A(B[534]), .Z(n492) );
  IV U565 ( .A(B[535]), .Z(n491) );
  IV U566 ( .A(B[536]), .Z(n490) );
  IV U567 ( .A(B[977]), .Z(n49) );
  IV U568 ( .A(B[537]), .Z(n489) );
  IV U569 ( .A(B[538]), .Z(n488) );
  IV U570 ( .A(B[539]), .Z(n487) );
  IV U571 ( .A(B[540]), .Z(n486) );
  IV U572 ( .A(B[541]), .Z(n485) );
  IV U573 ( .A(B[542]), .Z(n484) );
  IV U574 ( .A(B[543]), .Z(n483) );
  IV U575 ( .A(B[544]), .Z(n482) );
  IV U576 ( .A(B[545]), .Z(n481) );
  IV U577 ( .A(B[546]), .Z(n480) );
  IV U578 ( .A(B[978]), .Z(n48) );
  IV U579 ( .A(B[547]), .Z(n479) );
  IV U580 ( .A(B[548]), .Z(n478) );
  IV U581 ( .A(B[549]), .Z(n477) );
  IV U582 ( .A(B[550]), .Z(n476) );
  IV U583 ( .A(B[551]), .Z(n475) );
  IV U584 ( .A(B[552]), .Z(n474) );
  IV U585 ( .A(B[553]), .Z(n473) );
  IV U586 ( .A(B[554]), .Z(n472) );
  IV U587 ( .A(B[555]), .Z(n471) );
  IV U588 ( .A(B[556]), .Z(n470) );
  IV U589 ( .A(B[979]), .Z(n47) );
  IV U590 ( .A(B[557]), .Z(n469) );
  IV U591 ( .A(B[558]), .Z(n468) );
  IV U592 ( .A(B[559]), .Z(n467) );
  IV U593 ( .A(B[560]), .Z(n466) );
  IV U594 ( .A(B[561]), .Z(n465) );
  IV U595 ( .A(B[562]), .Z(n464) );
  IV U596 ( .A(B[563]), .Z(n463) );
  IV U597 ( .A(B[564]), .Z(n462) );
  IV U598 ( .A(B[565]), .Z(n461) );
  IV U599 ( .A(B[566]), .Z(n460) );
  IV U600 ( .A(B[980]), .Z(n46) );
  IV U601 ( .A(B[567]), .Z(n459) );
  IV U602 ( .A(B[568]), .Z(n458) );
  IV U603 ( .A(B[569]), .Z(n457) );
  IV U604 ( .A(B[570]), .Z(n456) );
  IV U605 ( .A(B[571]), .Z(n455) );
  IV U606 ( .A(B[572]), .Z(n454) );
  IV U607 ( .A(B[573]), .Z(n453) );
  IV U608 ( .A(B[574]), .Z(n452) );
  IV U609 ( .A(B[575]), .Z(n451) );
  IV U610 ( .A(B[576]), .Z(n450) );
  IV U611 ( .A(B[981]), .Z(n45) );
  IV U612 ( .A(B[577]), .Z(n449) );
  IV U613 ( .A(B[578]), .Z(n448) );
  IV U614 ( .A(B[579]), .Z(n447) );
  IV U615 ( .A(B[580]), .Z(n446) );
  IV U616 ( .A(B[581]), .Z(n445) );
  IV U617 ( .A(B[582]), .Z(n444) );
  IV U618 ( .A(B[583]), .Z(n443) );
  IV U619 ( .A(B[584]), .Z(n442) );
  IV U620 ( .A(B[585]), .Z(n441) );
  IV U621 ( .A(B[586]), .Z(n440) );
  IV U622 ( .A(B[982]), .Z(n44) );
  IV U623 ( .A(B[587]), .Z(n439) );
  IV U624 ( .A(B[588]), .Z(n438) );
  IV U625 ( .A(B[589]), .Z(n437) );
  IV U626 ( .A(B[590]), .Z(n436) );
  IV U627 ( .A(B[591]), .Z(n435) );
  IV U628 ( .A(B[592]), .Z(n434) );
  IV U629 ( .A(B[593]), .Z(n433) );
  IV U630 ( .A(B[594]), .Z(n432) );
  IV U631 ( .A(B[595]), .Z(n431) );
  IV U632 ( .A(B[596]), .Z(n430) );
  IV U633 ( .A(B[983]), .Z(n43) );
  IV U634 ( .A(B[597]), .Z(n429) );
  IV U635 ( .A(B[598]), .Z(n428) );
  IV U636 ( .A(B[599]), .Z(n427) );
  IV U637 ( .A(B[600]), .Z(n426) );
  IV U638 ( .A(B[601]), .Z(n425) );
  IV U639 ( .A(B[602]), .Z(n424) );
  IV U640 ( .A(B[603]), .Z(n423) );
  IV U641 ( .A(B[604]), .Z(n422) );
  IV U642 ( .A(B[605]), .Z(n421) );
  IV U643 ( .A(B[606]), .Z(n420) );
  IV U644 ( .A(B[984]), .Z(n42) );
  IV U645 ( .A(B[607]), .Z(n419) );
  IV U646 ( .A(B[608]), .Z(n418) );
  IV U647 ( .A(B[609]), .Z(n417) );
  IV U648 ( .A(B[610]), .Z(n416) );
  IV U649 ( .A(B[611]), .Z(n415) );
  IV U650 ( .A(B[612]), .Z(n414) );
  IV U651 ( .A(B[613]), .Z(n413) );
  IV U652 ( .A(B[614]), .Z(n412) );
  IV U653 ( .A(B[615]), .Z(n411) );
  IV U654 ( .A(B[616]), .Z(n410) );
  IV U655 ( .A(B[985]), .Z(n41) );
  IV U656 ( .A(B[617]), .Z(n409) );
  IV U657 ( .A(B[618]), .Z(n408) );
  IV U658 ( .A(B[619]), .Z(n407) );
  IV U659 ( .A(B[620]), .Z(n406) );
  IV U660 ( .A(B[621]), .Z(n405) );
  IV U661 ( .A(B[622]), .Z(n404) );
  IV U662 ( .A(B[623]), .Z(n403) );
  IV U663 ( .A(B[624]), .Z(n402) );
  IV U664 ( .A(B[625]), .Z(n401) );
  IV U665 ( .A(B[626]), .Z(n400) );
  IV U666 ( .A(B[986]), .Z(n40) );
  IV U667 ( .A(B[1022]), .Z(n4) );
  IV U668 ( .A(B[627]), .Z(n399) );
  IV U669 ( .A(B[628]), .Z(n398) );
  IV U670 ( .A(B[629]), .Z(n397) );
  IV U671 ( .A(B[630]), .Z(n396) );
  IV U672 ( .A(B[631]), .Z(n395) );
  IV U673 ( .A(B[632]), .Z(n394) );
  IV U674 ( .A(B[633]), .Z(n393) );
  IV U675 ( .A(B[634]), .Z(n392) );
  IV U676 ( .A(B[635]), .Z(n391) );
  IV U677 ( .A(B[636]), .Z(n390) );
  IV U678 ( .A(B[987]), .Z(n39) );
  IV U679 ( .A(B[637]), .Z(n389) );
  IV U680 ( .A(B[638]), .Z(n388) );
  IV U681 ( .A(B[639]), .Z(n387) );
  IV U682 ( .A(B[640]), .Z(n386) );
  IV U683 ( .A(B[641]), .Z(n385) );
  IV U684 ( .A(B[642]), .Z(n384) );
  IV U685 ( .A(B[643]), .Z(n383) );
  IV U686 ( .A(B[644]), .Z(n382) );
  IV U687 ( .A(B[645]), .Z(n381) );
  IV U688 ( .A(B[646]), .Z(n380) );
  IV U689 ( .A(B[988]), .Z(n38) );
  IV U690 ( .A(B[647]), .Z(n379) );
  IV U691 ( .A(B[648]), .Z(n378) );
  IV U692 ( .A(B[649]), .Z(n377) );
  IV U693 ( .A(B[650]), .Z(n376) );
  IV U694 ( .A(B[651]), .Z(n375) );
  IV U695 ( .A(B[652]), .Z(n374) );
  IV U696 ( .A(B[653]), .Z(n373) );
  IV U697 ( .A(B[654]), .Z(n372) );
  IV U698 ( .A(B[655]), .Z(n371) );
  IV U699 ( .A(B[656]), .Z(n370) );
  IV U700 ( .A(B[989]), .Z(n37) );
  IV U701 ( .A(B[657]), .Z(n369) );
  IV U702 ( .A(B[658]), .Z(n368) );
  IV U703 ( .A(B[659]), .Z(n367) );
  IV U704 ( .A(B[660]), .Z(n366) );
  IV U705 ( .A(B[661]), .Z(n365) );
  IV U706 ( .A(B[662]), .Z(n364) );
  IV U707 ( .A(B[663]), .Z(n363) );
  IV U708 ( .A(B[664]), .Z(n362) );
  IV U709 ( .A(B[665]), .Z(n361) );
  IV U710 ( .A(B[666]), .Z(n360) );
  IV U711 ( .A(B[990]), .Z(n36) );
  IV U712 ( .A(B[667]), .Z(n359) );
  IV U713 ( .A(B[668]), .Z(n358) );
  IV U714 ( .A(B[669]), .Z(n357) );
  IV U715 ( .A(B[670]), .Z(n356) );
  IV U716 ( .A(B[671]), .Z(n355) );
  IV U717 ( .A(B[672]), .Z(n354) );
  IV U718 ( .A(B[673]), .Z(n353) );
  IV U719 ( .A(B[674]), .Z(n352) );
  IV U720 ( .A(B[675]), .Z(n351) );
  IV U721 ( .A(B[676]), .Z(n350) );
  IV U722 ( .A(B[991]), .Z(n35) );
  IV U723 ( .A(B[677]), .Z(n349) );
  IV U724 ( .A(B[678]), .Z(n348) );
  IV U725 ( .A(B[679]), .Z(n347) );
  IV U726 ( .A(B[680]), .Z(n346) );
  IV U727 ( .A(B[681]), .Z(n345) );
  IV U728 ( .A(B[682]), .Z(n344) );
  IV U729 ( .A(B[683]), .Z(n343) );
  IV U730 ( .A(B[684]), .Z(n342) );
  IV U731 ( .A(B[685]), .Z(n341) );
  IV U732 ( .A(B[686]), .Z(n340) );
  IV U733 ( .A(B[992]), .Z(n34) );
  IV U734 ( .A(B[687]), .Z(n339) );
  IV U735 ( .A(B[688]), .Z(n338) );
  IV U736 ( .A(B[689]), .Z(n337) );
  IV U737 ( .A(B[690]), .Z(n336) );
  IV U738 ( .A(B[691]), .Z(n335) );
  IV U739 ( .A(B[692]), .Z(n334) );
  IV U740 ( .A(B[693]), .Z(n333) );
  IV U741 ( .A(B[694]), .Z(n332) );
  IV U742 ( .A(B[695]), .Z(n331) );
  IV U743 ( .A(B[696]), .Z(n330) );
  IV U744 ( .A(B[993]), .Z(n33) );
  IV U745 ( .A(B[697]), .Z(n329) );
  IV U746 ( .A(B[698]), .Z(n328) );
  IV U747 ( .A(B[699]), .Z(n327) );
  IV U748 ( .A(B[700]), .Z(n326) );
  IV U749 ( .A(B[701]), .Z(n325) );
  IV U750 ( .A(B[702]), .Z(n324) );
  IV U751 ( .A(B[703]), .Z(n323) );
  IV U752 ( .A(B[704]), .Z(n322) );
  IV U753 ( .A(B[705]), .Z(n321) );
  IV U754 ( .A(B[706]), .Z(n320) );
  IV U755 ( .A(B[994]), .Z(n32) );
  IV U756 ( .A(B[707]), .Z(n319) );
  IV U757 ( .A(B[708]), .Z(n318) );
  IV U758 ( .A(B[709]), .Z(n317) );
  IV U759 ( .A(B[710]), .Z(n316) );
  IV U760 ( .A(B[711]), .Z(n315) );
  IV U761 ( .A(B[712]), .Z(n314) );
  IV U762 ( .A(B[713]), .Z(n313) );
  IV U763 ( .A(B[714]), .Z(n312) );
  IV U764 ( .A(B[715]), .Z(n311) );
  IV U765 ( .A(B[716]), .Z(n310) );
  IV U766 ( .A(B[995]), .Z(n31) );
  IV U767 ( .A(B[717]), .Z(n309) );
  IV U768 ( .A(B[718]), .Z(n308) );
  IV U769 ( .A(B[719]), .Z(n307) );
  IV U770 ( .A(B[720]), .Z(n306) );
  IV U771 ( .A(B[721]), .Z(n305) );
  IV U772 ( .A(B[722]), .Z(n304) );
  IV U773 ( .A(B[723]), .Z(n303) );
  IV U774 ( .A(B[724]), .Z(n302) );
  IV U775 ( .A(B[725]), .Z(n301) );
  IV U776 ( .A(B[726]), .Z(n300) );
  IV U777 ( .A(B[996]), .Z(n30) );
  IV U778 ( .A(B[1023]), .Z(n3) );
  IV U779 ( .A(B[727]), .Z(n299) );
  IV U780 ( .A(B[728]), .Z(n298) );
  IV U781 ( .A(B[729]), .Z(n297) );
  IV U782 ( .A(B[730]), .Z(n296) );
  IV U783 ( .A(B[731]), .Z(n295) );
  IV U784 ( .A(B[732]), .Z(n294) );
  IV U785 ( .A(B[733]), .Z(n293) );
  IV U786 ( .A(B[734]), .Z(n292) );
  IV U787 ( .A(B[735]), .Z(n291) );
  IV U788 ( .A(B[736]), .Z(n290) );
  IV U789 ( .A(B[997]), .Z(n29) );
  IV U790 ( .A(B[737]), .Z(n289) );
  IV U791 ( .A(B[738]), .Z(n288) );
  IV U792 ( .A(B[739]), .Z(n287) );
  IV U793 ( .A(B[740]), .Z(n286) );
  IV U794 ( .A(B[741]), .Z(n285) );
  IV U795 ( .A(B[742]), .Z(n284) );
  IV U796 ( .A(B[743]), .Z(n283) );
  IV U797 ( .A(B[744]), .Z(n282) );
  IV U798 ( .A(B[745]), .Z(n281) );
  IV U799 ( .A(B[746]), .Z(n280) );
  IV U800 ( .A(B[998]), .Z(n28) );
  IV U801 ( .A(B[747]), .Z(n279) );
  IV U802 ( .A(B[748]), .Z(n278) );
  IV U803 ( .A(B[749]), .Z(n277) );
  IV U804 ( .A(B[750]), .Z(n276) );
  IV U805 ( .A(B[751]), .Z(n275) );
  IV U806 ( .A(B[752]), .Z(n274) );
  IV U807 ( .A(B[753]), .Z(n273) );
  IV U808 ( .A(B[754]), .Z(n272) );
  IV U809 ( .A(B[755]), .Z(n271) );
  IV U810 ( .A(B[756]), .Z(n270) );
  IV U811 ( .A(B[999]), .Z(n27) );
  IV U812 ( .A(B[757]), .Z(n269) );
  IV U813 ( .A(B[758]), .Z(n268) );
  IV U814 ( .A(B[759]), .Z(n267) );
  IV U815 ( .A(B[760]), .Z(n266) );
  IV U816 ( .A(B[761]), .Z(n265) );
  IV U817 ( .A(B[762]), .Z(n264) );
  IV U818 ( .A(B[763]), .Z(n263) );
  IV U819 ( .A(B[764]), .Z(n262) );
  IV U820 ( .A(B[765]), .Z(n261) );
  IV U821 ( .A(B[766]), .Z(n260) );
  IV U822 ( .A(B[1000]), .Z(n26) );
  IV U823 ( .A(B[767]), .Z(n259) );
  IV U824 ( .A(B[768]), .Z(n258) );
  IV U825 ( .A(B[769]), .Z(n257) );
  IV U826 ( .A(B[770]), .Z(n256) );
  IV U827 ( .A(B[771]), .Z(n255) );
  IV U828 ( .A(B[772]), .Z(n254) );
  IV U829 ( .A(B[773]), .Z(n253) );
  IV U830 ( .A(B[774]), .Z(n252) );
  IV U831 ( .A(B[775]), .Z(n251) );
  IV U832 ( .A(B[776]), .Z(n250) );
  IV U833 ( .A(B[1001]), .Z(n25) );
  IV U834 ( .A(B[777]), .Z(n249) );
  IV U835 ( .A(B[778]), .Z(n248) );
  IV U836 ( .A(B[779]), .Z(n247) );
  IV U837 ( .A(B[780]), .Z(n246) );
  IV U838 ( .A(B[781]), .Z(n245) );
  IV U839 ( .A(B[782]), .Z(n244) );
  IV U840 ( .A(B[783]), .Z(n243) );
  IV U841 ( .A(B[784]), .Z(n242) );
  IV U842 ( .A(B[785]), .Z(n241) );
  IV U843 ( .A(B[786]), .Z(n240) );
  IV U844 ( .A(B[1002]), .Z(n24) );
  IV U845 ( .A(B[787]), .Z(n239) );
  IV U846 ( .A(B[788]), .Z(n238) );
  IV U847 ( .A(B[789]), .Z(n237) );
  IV U848 ( .A(B[790]), .Z(n236) );
  IV U849 ( .A(B[791]), .Z(n235) );
  IV U850 ( .A(B[792]), .Z(n234) );
  IV U851 ( .A(B[793]), .Z(n233) );
  IV U852 ( .A(B[794]), .Z(n232) );
  IV U853 ( .A(B[795]), .Z(n231) );
  IV U854 ( .A(B[796]), .Z(n230) );
  IV U855 ( .A(B[1003]), .Z(n23) );
  IV U856 ( .A(B[797]), .Z(n229) );
  IV U857 ( .A(B[798]), .Z(n228) );
  IV U858 ( .A(B[799]), .Z(n227) );
  IV U859 ( .A(B[800]), .Z(n226) );
  IV U860 ( .A(B[801]), .Z(n225) );
  IV U861 ( .A(B[802]), .Z(n224) );
  IV U862 ( .A(B[803]), .Z(n223) );
  IV U863 ( .A(B[804]), .Z(n222) );
  IV U864 ( .A(B[805]), .Z(n221) );
  IV U865 ( .A(B[806]), .Z(n220) );
  IV U866 ( .A(B[1004]), .Z(n22) );
  IV U867 ( .A(B[807]), .Z(n219) );
  IV U868 ( .A(B[808]), .Z(n218) );
  IV U869 ( .A(B[809]), .Z(n217) );
  IV U870 ( .A(B[810]), .Z(n216) );
  IV U871 ( .A(B[811]), .Z(n215) );
  IV U872 ( .A(B[812]), .Z(n214) );
  IV U873 ( .A(B[813]), .Z(n213) );
  IV U874 ( .A(B[814]), .Z(n212) );
  IV U875 ( .A(B[815]), .Z(n211) );
  IV U876 ( .A(B[816]), .Z(n210) );
  IV U877 ( .A(B[1005]), .Z(n21) );
  IV U878 ( .A(B[817]), .Z(n209) );
  IV U879 ( .A(B[818]), .Z(n208) );
  IV U880 ( .A(B[819]), .Z(n207) );
  IV U881 ( .A(B[820]), .Z(n206) );
  IV U882 ( .A(B[821]), .Z(n205) );
  IV U883 ( .A(B[822]), .Z(n204) );
  IV U884 ( .A(B[823]), .Z(n203) );
  IV U885 ( .A(B[824]), .Z(n202) );
  IV U886 ( .A(B[825]), .Z(n201) );
  IV U887 ( .A(B[826]), .Z(n200) );
  IV U888 ( .A(B[1006]), .Z(n20) );
  IV U889 ( .A(B[827]), .Z(n199) );
  IV U890 ( .A(B[828]), .Z(n198) );
  IV U891 ( .A(B[829]), .Z(n197) );
  IV U892 ( .A(B[830]), .Z(n196) );
  IV U893 ( .A(B[831]), .Z(n195) );
  IV U894 ( .A(B[832]), .Z(n194) );
  IV U895 ( .A(B[833]), .Z(n193) );
  IV U896 ( .A(B[834]), .Z(n192) );
  IV U897 ( .A(B[835]), .Z(n191) );
  IV U898 ( .A(B[836]), .Z(n190) );
  IV U899 ( .A(B[1007]), .Z(n19) );
  IV U900 ( .A(B[837]), .Z(n189) );
  IV U901 ( .A(B[838]), .Z(n188) );
  IV U902 ( .A(B[839]), .Z(n187) );
  IV U903 ( .A(B[840]), .Z(n186) );
  IV U904 ( .A(B[841]), .Z(n185) );
  IV U905 ( .A(B[842]), .Z(n184) );
  IV U906 ( .A(B[843]), .Z(n183) );
  IV U907 ( .A(B[844]), .Z(n182) );
  IV U908 ( .A(B[845]), .Z(n181) );
  IV U909 ( .A(B[846]), .Z(n180) );
  IV U910 ( .A(B[1008]), .Z(n18) );
  IV U911 ( .A(B[847]), .Z(n179) );
  IV U912 ( .A(B[848]), .Z(n178) );
  IV U913 ( .A(B[849]), .Z(n177) );
  IV U914 ( .A(B[850]), .Z(n176) );
  IV U915 ( .A(B[851]), .Z(n175) );
  IV U916 ( .A(B[852]), .Z(n174) );
  IV U917 ( .A(B[853]), .Z(n173) );
  IV U918 ( .A(B[854]), .Z(n172) );
  IV U919 ( .A(B[855]), .Z(n171) );
  IV U920 ( .A(B[856]), .Z(n170) );
  IV U921 ( .A(B[1009]), .Z(n17) );
  IV U922 ( .A(B[857]), .Z(n169) );
  IV U923 ( .A(B[858]), .Z(n168) );
  IV U924 ( .A(B[859]), .Z(n167) );
  IV U925 ( .A(B[860]), .Z(n166) );
  IV U926 ( .A(B[861]), .Z(n165) );
  IV U927 ( .A(B[862]), .Z(n164) );
  IV U928 ( .A(B[863]), .Z(n163) );
  IV U929 ( .A(B[864]), .Z(n162) );
  IV U930 ( .A(B[865]), .Z(n161) );
  IV U931 ( .A(B[866]), .Z(n160) );
  IV U932 ( .A(B[1010]), .Z(n16) );
  IV U933 ( .A(B[867]), .Z(n159) );
  IV U934 ( .A(B[868]), .Z(n158) );
  IV U935 ( .A(B[869]), .Z(n157) );
  IV U936 ( .A(B[870]), .Z(n156) );
  IV U937 ( .A(B[871]), .Z(n155) );
  IV U938 ( .A(B[872]), .Z(n154) );
  IV U939 ( .A(B[873]), .Z(n153) );
  IV U940 ( .A(B[874]), .Z(n152) );
  IV U941 ( .A(B[875]), .Z(n151) );
  IV U942 ( .A(B[876]), .Z(n150) );
  IV U943 ( .A(B[1011]), .Z(n15) );
  IV U944 ( .A(B[877]), .Z(n149) );
  IV U945 ( .A(B[878]), .Z(n148) );
  IV U946 ( .A(B[879]), .Z(n147) );
  IV U947 ( .A(B[880]), .Z(n146) );
  IV U948 ( .A(B[881]), .Z(n145) );
  IV U949 ( .A(B[882]), .Z(n144) );
  IV U950 ( .A(B[883]), .Z(n143) );
  IV U951 ( .A(B[884]), .Z(n142) );
  IV U952 ( .A(B[885]), .Z(n141) );
  IV U953 ( .A(B[886]), .Z(n140) );
  IV U954 ( .A(B[1012]), .Z(n14) );
  IV U955 ( .A(B[887]), .Z(n139) );
  IV U956 ( .A(B[888]), .Z(n138) );
  IV U957 ( .A(B[889]), .Z(n137) );
  IV U958 ( .A(B[890]), .Z(n136) );
  IV U959 ( .A(B[891]), .Z(n135) );
  IV U960 ( .A(B[892]), .Z(n134) );
  IV U961 ( .A(B[893]), .Z(n133) );
  IV U962 ( .A(B[894]), .Z(n132) );
  IV U963 ( .A(B[895]), .Z(n131) );
  IV U964 ( .A(B[896]), .Z(n130) );
  IV U965 ( .A(B[1013]), .Z(n13) );
  IV U966 ( .A(B[897]), .Z(n129) );
  IV U967 ( .A(B[898]), .Z(n128) );
  IV U968 ( .A(B[899]), .Z(n127) );
  IV U969 ( .A(B[900]), .Z(n126) );
  IV U970 ( .A(B[901]), .Z(n125) );
  IV U971 ( .A(B[902]), .Z(n124) );
  IV U972 ( .A(B[903]), .Z(n123) );
  IV U973 ( .A(B[904]), .Z(n122) );
  IV U974 ( .A(B[905]), .Z(n121) );
  IV U975 ( .A(B[906]), .Z(n120) );
  IV U976 ( .A(B[1014]), .Z(n12) );
  IV U977 ( .A(B[907]), .Z(n119) );
  IV U978 ( .A(B[908]), .Z(n118) );
  IV U979 ( .A(B[909]), .Z(n117) );
  IV U980 ( .A(B[910]), .Z(n116) );
  IV U981 ( .A(B[911]), .Z(n115) );
  IV U982 ( .A(B[912]), .Z(n114) );
  IV U983 ( .A(B[913]), .Z(n113) );
  IV U984 ( .A(B[914]), .Z(n112) );
  IV U985 ( .A(B[915]), .Z(n111) );
  IV U986 ( .A(B[916]), .Z(n110) );
  IV U987 ( .A(B[1015]), .Z(n11) );
  IV U988 ( .A(B[917]), .Z(n109) );
  IV U989 ( .A(B[918]), .Z(n108) );
  IV U990 ( .A(B[919]), .Z(n107) );
  IV U991 ( .A(B[920]), .Z(n106) );
  IV U992 ( .A(B[921]), .Z(n105) );
  IV U993 ( .A(B[922]), .Z(n104) );
  IV U994 ( .A(B[923]), .Z(n103) );
  IV U995 ( .A(B[0]), .Z(n1026) );
  IV U996 ( .A(B[1]), .Z(n1025) );
  IV U997 ( .A(B[2]), .Z(n1024) );
  IV U998 ( .A(B[3]), .Z(n1023) );
  IV U999 ( .A(B[4]), .Z(n1022) );
  IV U1000 ( .A(B[5]), .Z(n1021) );
  IV U1001 ( .A(B[6]), .Z(n1020) );
  IV U1002 ( .A(B[924]), .Z(n102) );
  IV U1003 ( .A(B[7]), .Z(n1019) );
  IV U1004 ( .A(B[8]), .Z(n1018) );
  IV U1005 ( .A(B[9]), .Z(n1017) );
  IV U1006 ( .A(B[10]), .Z(n1016) );
  IV U1007 ( .A(B[11]), .Z(n1015) );
  IV U1008 ( .A(B[12]), .Z(n1014) );
  IV U1009 ( .A(B[13]), .Z(n1013) );
  IV U1010 ( .A(B[14]), .Z(n1012) );
  IV U1011 ( .A(B[15]), .Z(n1011) );
  IV U1012 ( .A(B[16]), .Z(n1010) );
  IV U1013 ( .A(B[925]), .Z(n101) );
  IV U1014 ( .A(B[17]), .Z(n1009) );
  IV U1015 ( .A(B[18]), .Z(n1008) );
  IV U1016 ( .A(B[19]), .Z(n1007) );
  IV U1017 ( .A(B[20]), .Z(n1006) );
  IV U1018 ( .A(B[21]), .Z(n1005) );
  IV U1019 ( .A(B[22]), .Z(n1004) );
  IV U1020 ( .A(B[23]), .Z(n1003) );
  IV U1021 ( .A(B[24]), .Z(n1002) );
  IV U1022 ( .A(B[25]), .Z(n1001) );
  IV U1023 ( .A(B[26]), .Z(n1000) );
  IV U1024 ( .A(B[926]), .Z(n100) );
  IV U1025 ( .A(B[1016]), .Z(n10) );
endmodule


module MUX_N1026_1 ( A, B, S, O );
  input [1025:0] A;
  input [1025:0] B;
  output [1025:0] O;
  input S;


  ANDN U1 ( .B(A[9]), .A(S), .Z(O[9]) );
  ANDN U2 ( .B(A[99]), .A(S), .Z(O[99]) );
  ANDN U3 ( .B(A[999]), .A(S), .Z(O[999]) );
  ANDN U4 ( .B(A[998]), .A(S), .Z(O[998]) );
  ANDN U5 ( .B(A[997]), .A(S), .Z(O[997]) );
  ANDN U6 ( .B(A[996]), .A(S), .Z(O[996]) );
  ANDN U7 ( .B(A[995]), .A(S), .Z(O[995]) );
  ANDN U8 ( .B(A[994]), .A(S), .Z(O[994]) );
  ANDN U9 ( .B(A[993]), .A(S), .Z(O[993]) );
  ANDN U10 ( .B(A[992]), .A(S), .Z(O[992]) );
  ANDN U11 ( .B(A[991]), .A(S), .Z(O[991]) );
  ANDN U12 ( .B(A[990]), .A(S), .Z(O[990]) );
  ANDN U13 ( .B(A[98]), .A(S), .Z(O[98]) );
  ANDN U14 ( .B(A[989]), .A(S), .Z(O[989]) );
  ANDN U15 ( .B(A[988]), .A(S), .Z(O[988]) );
  ANDN U16 ( .B(A[987]), .A(S), .Z(O[987]) );
  ANDN U17 ( .B(A[986]), .A(S), .Z(O[986]) );
  ANDN U18 ( .B(A[985]), .A(S), .Z(O[985]) );
  ANDN U19 ( .B(A[984]), .A(S), .Z(O[984]) );
  ANDN U20 ( .B(A[983]), .A(S), .Z(O[983]) );
  ANDN U21 ( .B(A[982]), .A(S), .Z(O[982]) );
  ANDN U22 ( .B(A[981]), .A(S), .Z(O[981]) );
  ANDN U23 ( .B(A[980]), .A(S), .Z(O[980]) );
  ANDN U24 ( .B(A[97]), .A(S), .Z(O[97]) );
  ANDN U25 ( .B(A[979]), .A(S), .Z(O[979]) );
  ANDN U26 ( .B(A[978]), .A(S), .Z(O[978]) );
  ANDN U27 ( .B(A[977]), .A(S), .Z(O[977]) );
  ANDN U28 ( .B(A[976]), .A(S), .Z(O[976]) );
  ANDN U29 ( .B(A[975]), .A(S), .Z(O[975]) );
  ANDN U30 ( .B(A[974]), .A(S), .Z(O[974]) );
  ANDN U31 ( .B(A[973]), .A(S), .Z(O[973]) );
  ANDN U32 ( .B(A[972]), .A(S), .Z(O[972]) );
  ANDN U33 ( .B(A[971]), .A(S), .Z(O[971]) );
  ANDN U34 ( .B(A[970]), .A(S), .Z(O[970]) );
  ANDN U35 ( .B(A[96]), .A(S), .Z(O[96]) );
  ANDN U36 ( .B(A[969]), .A(S), .Z(O[969]) );
  ANDN U37 ( .B(A[968]), .A(S), .Z(O[968]) );
  ANDN U38 ( .B(A[967]), .A(S), .Z(O[967]) );
  ANDN U39 ( .B(A[966]), .A(S), .Z(O[966]) );
  ANDN U40 ( .B(A[965]), .A(S), .Z(O[965]) );
  ANDN U41 ( .B(A[964]), .A(S), .Z(O[964]) );
  ANDN U42 ( .B(A[963]), .A(S), .Z(O[963]) );
  ANDN U43 ( .B(A[962]), .A(S), .Z(O[962]) );
  ANDN U44 ( .B(A[961]), .A(S), .Z(O[961]) );
  ANDN U45 ( .B(A[960]), .A(S), .Z(O[960]) );
  ANDN U46 ( .B(A[95]), .A(S), .Z(O[95]) );
  ANDN U47 ( .B(A[959]), .A(S), .Z(O[959]) );
  ANDN U48 ( .B(A[958]), .A(S), .Z(O[958]) );
  ANDN U49 ( .B(A[957]), .A(S), .Z(O[957]) );
  ANDN U50 ( .B(A[956]), .A(S), .Z(O[956]) );
  ANDN U51 ( .B(A[955]), .A(S), .Z(O[955]) );
  ANDN U52 ( .B(A[954]), .A(S), .Z(O[954]) );
  ANDN U53 ( .B(A[953]), .A(S), .Z(O[953]) );
  ANDN U54 ( .B(A[952]), .A(S), .Z(O[952]) );
  ANDN U55 ( .B(A[951]), .A(S), .Z(O[951]) );
  ANDN U56 ( .B(A[950]), .A(S), .Z(O[950]) );
  ANDN U57 ( .B(A[94]), .A(S), .Z(O[94]) );
  ANDN U58 ( .B(A[949]), .A(S), .Z(O[949]) );
  ANDN U59 ( .B(A[948]), .A(S), .Z(O[948]) );
  ANDN U60 ( .B(A[947]), .A(S), .Z(O[947]) );
  ANDN U61 ( .B(A[946]), .A(S), .Z(O[946]) );
  ANDN U62 ( .B(A[945]), .A(S), .Z(O[945]) );
  ANDN U63 ( .B(A[944]), .A(S), .Z(O[944]) );
  ANDN U64 ( .B(A[943]), .A(S), .Z(O[943]) );
  ANDN U65 ( .B(A[942]), .A(S), .Z(O[942]) );
  ANDN U66 ( .B(A[941]), .A(S), .Z(O[941]) );
  ANDN U67 ( .B(A[940]), .A(S), .Z(O[940]) );
  ANDN U68 ( .B(A[93]), .A(S), .Z(O[93]) );
  ANDN U69 ( .B(A[939]), .A(S), .Z(O[939]) );
  ANDN U70 ( .B(A[938]), .A(S), .Z(O[938]) );
  ANDN U71 ( .B(A[937]), .A(S), .Z(O[937]) );
  ANDN U72 ( .B(A[936]), .A(S), .Z(O[936]) );
  ANDN U73 ( .B(A[935]), .A(S), .Z(O[935]) );
  ANDN U74 ( .B(A[934]), .A(S), .Z(O[934]) );
  ANDN U75 ( .B(A[933]), .A(S), .Z(O[933]) );
  ANDN U76 ( .B(A[932]), .A(S), .Z(O[932]) );
  ANDN U77 ( .B(A[931]), .A(S), .Z(O[931]) );
  ANDN U78 ( .B(A[930]), .A(S), .Z(O[930]) );
  ANDN U79 ( .B(A[92]), .A(S), .Z(O[92]) );
  ANDN U80 ( .B(A[929]), .A(S), .Z(O[929]) );
  ANDN U81 ( .B(A[928]), .A(S), .Z(O[928]) );
  ANDN U82 ( .B(A[927]), .A(S), .Z(O[927]) );
  ANDN U83 ( .B(A[926]), .A(S), .Z(O[926]) );
  ANDN U84 ( .B(A[925]), .A(S), .Z(O[925]) );
  ANDN U85 ( .B(A[924]), .A(S), .Z(O[924]) );
  ANDN U86 ( .B(A[923]), .A(S), .Z(O[923]) );
  ANDN U87 ( .B(A[922]), .A(S), .Z(O[922]) );
  ANDN U88 ( .B(A[921]), .A(S), .Z(O[921]) );
  ANDN U89 ( .B(A[920]), .A(S), .Z(O[920]) );
  ANDN U90 ( .B(A[91]), .A(S), .Z(O[91]) );
  ANDN U91 ( .B(A[919]), .A(S), .Z(O[919]) );
  ANDN U92 ( .B(A[918]), .A(S), .Z(O[918]) );
  ANDN U93 ( .B(A[917]), .A(S), .Z(O[917]) );
  ANDN U94 ( .B(A[916]), .A(S), .Z(O[916]) );
  ANDN U95 ( .B(A[915]), .A(S), .Z(O[915]) );
  ANDN U96 ( .B(A[914]), .A(S), .Z(O[914]) );
  ANDN U97 ( .B(A[913]), .A(S), .Z(O[913]) );
  ANDN U98 ( .B(A[912]), .A(S), .Z(O[912]) );
  ANDN U99 ( .B(A[911]), .A(S), .Z(O[911]) );
  ANDN U100 ( .B(A[910]), .A(S), .Z(O[910]) );
  ANDN U101 ( .B(A[90]), .A(S), .Z(O[90]) );
  ANDN U102 ( .B(A[909]), .A(S), .Z(O[909]) );
  ANDN U103 ( .B(A[908]), .A(S), .Z(O[908]) );
  ANDN U104 ( .B(A[907]), .A(S), .Z(O[907]) );
  ANDN U105 ( .B(A[906]), .A(S), .Z(O[906]) );
  ANDN U106 ( .B(A[905]), .A(S), .Z(O[905]) );
  ANDN U107 ( .B(A[904]), .A(S), .Z(O[904]) );
  ANDN U108 ( .B(A[903]), .A(S), .Z(O[903]) );
  ANDN U109 ( .B(A[902]), .A(S), .Z(O[902]) );
  ANDN U110 ( .B(A[901]), .A(S), .Z(O[901]) );
  ANDN U111 ( .B(A[900]), .A(S), .Z(O[900]) );
  ANDN U112 ( .B(A[8]), .A(S), .Z(O[8]) );
  ANDN U113 ( .B(A[89]), .A(S), .Z(O[89]) );
  ANDN U114 ( .B(A[899]), .A(S), .Z(O[899]) );
  ANDN U115 ( .B(A[898]), .A(S), .Z(O[898]) );
  ANDN U116 ( .B(A[897]), .A(S), .Z(O[897]) );
  ANDN U117 ( .B(A[896]), .A(S), .Z(O[896]) );
  ANDN U118 ( .B(A[895]), .A(S), .Z(O[895]) );
  ANDN U119 ( .B(A[894]), .A(S), .Z(O[894]) );
  ANDN U120 ( .B(A[893]), .A(S), .Z(O[893]) );
  ANDN U121 ( .B(A[892]), .A(S), .Z(O[892]) );
  ANDN U122 ( .B(A[891]), .A(S), .Z(O[891]) );
  ANDN U123 ( .B(A[890]), .A(S), .Z(O[890]) );
  ANDN U124 ( .B(A[88]), .A(S), .Z(O[88]) );
  ANDN U125 ( .B(A[889]), .A(S), .Z(O[889]) );
  ANDN U126 ( .B(A[888]), .A(S), .Z(O[888]) );
  ANDN U127 ( .B(A[887]), .A(S), .Z(O[887]) );
  ANDN U128 ( .B(A[886]), .A(S), .Z(O[886]) );
  ANDN U129 ( .B(A[885]), .A(S), .Z(O[885]) );
  ANDN U130 ( .B(A[884]), .A(S), .Z(O[884]) );
  ANDN U131 ( .B(A[883]), .A(S), .Z(O[883]) );
  ANDN U132 ( .B(A[882]), .A(S), .Z(O[882]) );
  ANDN U133 ( .B(A[881]), .A(S), .Z(O[881]) );
  ANDN U134 ( .B(A[880]), .A(S), .Z(O[880]) );
  ANDN U135 ( .B(A[87]), .A(S), .Z(O[87]) );
  ANDN U136 ( .B(A[879]), .A(S), .Z(O[879]) );
  ANDN U137 ( .B(A[878]), .A(S), .Z(O[878]) );
  ANDN U138 ( .B(A[877]), .A(S), .Z(O[877]) );
  ANDN U139 ( .B(A[876]), .A(S), .Z(O[876]) );
  ANDN U140 ( .B(A[875]), .A(S), .Z(O[875]) );
  ANDN U141 ( .B(A[874]), .A(S), .Z(O[874]) );
  ANDN U142 ( .B(A[873]), .A(S), .Z(O[873]) );
  ANDN U143 ( .B(A[872]), .A(S), .Z(O[872]) );
  ANDN U144 ( .B(A[871]), .A(S), .Z(O[871]) );
  ANDN U145 ( .B(A[870]), .A(S), .Z(O[870]) );
  ANDN U146 ( .B(A[86]), .A(S), .Z(O[86]) );
  ANDN U147 ( .B(A[869]), .A(S), .Z(O[869]) );
  ANDN U148 ( .B(A[868]), .A(S), .Z(O[868]) );
  ANDN U149 ( .B(A[867]), .A(S), .Z(O[867]) );
  ANDN U150 ( .B(A[866]), .A(S), .Z(O[866]) );
  ANDN U151 ( .B(A[865]), .A(S), .Z(O[865]) );
  ANDN U152 ( .B(A[864]), .A(S), .Z(O[864]) );
  ANDN U153 ( .B(A[863]), .A(S), .Z(O[863]) );
  ANDN U154 ( .B(A[862]), .A(S), .Z(O[862]) );
  ANDN U155 ( .B(A[861]), .A(S), .Z(O[861]) );
  ANDN U156 ( .B(A[860]), .A(S), .Z(O[860]) );
  ANDN U157 ( .B(A[85]), .A(S), .Z(O[85]) );
  ANDN U158 ( .B(A[859]), .A(S), .Z(O[859]) );
  ANDN U159 ( .B(A[858]), .A(S), .Z(O[858]) );
  ANDN U160 ( .B(A[857]), .A(S), .Z(O[857]) );
  ANDN U161 ( .B(A[856]), .A(S), .Z(O[856]) );
  ANDN U162 ( .B(A[855]), .A(S), .Z(O[855]) );
  ANDN U163 ( .B(A[854]), .A(S), .Z(O[854]) );
  ANDN U164 ( .B(A[853]), .A(S), .Z(O[853]) );
  ANDN U165 ( .B(A[852]), .A(S), .Z(O[852]) );
  ANDN U166 ( .B(A[851]), .A(S), .Z(O[851]) );
  ANDN U167 ( .B(A[850]), .A(S), .Z(O[850]) );
  ANDN U168 ( .B(A[84]), .A(S), .Z(O[84]) );
  ANDN U169 ( .B(A[849]), .A(S), .Z(O[849]) );
  ANDN U170 ( .B(A[848]), .A(S), .Z(O[848]) );
  ANDN U171 ( .B(A[847]), .A(S), .Z(O[847]) );
  ANDN U172 ( .B(A[846]), .A(S), .Z(O[846]) );
  ANDN U173 ( .B(A[845]), .A(S), .Z(O[845]) );
  ANDN U174 ( .B(A[844]), .A(S), .Z(O[844]) );
  ANDN U175 ( .B(A[843]), .A(S), .Z(O[843]) );
  ANDN U176 ( .B(A[842]), .A(S), .Z(O[842]) );
  ANDN U177 ( .B(A[841]), .A(S), .Z(O[841]) );
  ANDN U178 ( .B(A[840]), .A(S), .Z(O[840]) );
  ANDN U179 ( .B(A[83]), .A(S), .Z(O[83]) );
  ANDN U180 ( .B(A[839]), .A(S), .Z(O[839]) );
  ANDN U181 ( .B(A[838]), .A(S), .Z(O[838]) );
  ANDN U182 ( .B(A[837]), .A(S), .Z(O[837]) );
  ANDN U183 ( .B(A[836]), .A(S), .Z(O[836]) );
  ANDN U184 ( .B(A[835]), .A(S), .Z(O[835]) );
  ANDN U185 ( .B(A[834]), .A(S), .Z(O[834]) );
  ANDN U186 ( .B(A[833]), .A(S), .Z(O[833]) );
  ANDN U187 ( .B(A[832]), .A(S), .Z(O[832]) );
  ANDN U188 ( .B(A[831]), .A(S), .Z(O[831]) );
  ANDN U189 ( .B(A[830]), .A(S), .Z(O[830]) );
  ANDN U190 ( .B(A[82]), .A(S), .Z(O[82]) );
  ANDN U191 ( .B(A[829]), .A(S), .Z(O[829]) );
  ANDN U192 ( .B(A[828]), .A(S), .Z(O[828]) );
  ANDN U193 ( .B(A[827]), .A(S), .Z(O[827]) );
  ANDN U194 ( .B(A[826]), .A(S), .Z(O[826]) );
  ANDN U195 ( .B(A[825]), .A(S), .Z(O[825]) );
  ANDN U196 ( .B(A[824]), .A(S), .Z(O[824]) );
  ANDN U197 ( .B(A[823]), .A(S), .Z(O[823]) );
  ANDN U198 ( .B(A[822]), .A(S), .Z(O[822]) );
  ANDN U199 ( .B(A[821]), .A(S), .Z(O[821]) );
  ANDN U200 ( .B(A[820]), .A(S), .Z(O[820]) );
  ANDN U201 ( .B(A[81]), .A(S), .Z(O[81]) );
  ANDN U202 ( .B(A[819]), .A(S), .Z(O[819]) );
  ANDN U203 ( .B(A[818]), .A(S), .Z(O[818]) );
  ANDN U204 ( .B(A[817]), .A(S), .Z(O[817]) );
  ANDN U205 ( .B(A[816]), .A(S), .Z(O[816]) );
  ANDN U206 ( .B(A[815]), .A(S), .Z(O[815]) );
  ANDN U207 ( .B(A[814]), .A(S), .Z(O[814]) );
  ANDN U208 ( .B(A[813]), .A(S), .Z(O[813]) );
  ANDN U209 ( .B(A[812]), .A(S), .Z(O[812]) );
  ANDN U210 ( .B(A[811]), .A(S), .Z(O[811]) );
  ANDN U211 ( .B(A[810]), .A(S), .Z(O[810]) );
  ANDN U212 ( .B(A[80]), .A(S), .Z(O[80]) );
  ANDN U213 ( .B(A[809]), .A(S), .Z(O[809]) );
  ANDN U214 ( .B(A[808]), .A(S), .Z(O[808]) );
  ANDN U215 ( .B(A[807]), .A(S), .Z(O[807]) );
  ANDN U216 ( .B(A[806]), .A(S), .Z(O[806]) );
  ANDN U217 ( .B(A[805]), .A(S), .Z(O[805]) );
  ANDN U218 ( .B(A[804]), .A(S), .Z(O[804]) );
  ANDN U219 ( .B(A[803]), .A(S), .Z(O[803]) );
  ANDN U220 ( .B(A[802]), .A(S), .Z(O[802]) );
  ANDN U221 ( .B(A[801]), .A(S), .Z(O[801]) );
  ANDN U222 ( .B(A[800]), .A(S), .Z(O[800]) );
  ANDN U223 ( .B(A[7]), .A(S), .Z(O[7]) );
  ANDN U224 ( .B(A[79]), .A(S), .Z(O[79]) );
  ANDN U225 ( .B(A[799]), .A(S), .Z(O[799]) );
  ANDN U226 ( .B(A[798]), .A(S), .Z(O[798]) );
  ANDN U227 ( .B(A[797]), .A(S), .Z(O[797]) );
  ANDN U228 ( .B(A[796]), .A(S), .Z(O[796]) );
  ANDN U229 ( .B(A[795]), .A(S), .Z(O[795]) );
  ANDN U230 ( .B(A[794]), .A(S), .Z(O[794]) );
  ANDN U231 ( .B(A[793]), .A(S), .Z(O[793]) );
  ANDN U232 ( .B(A[792]), .A(S), .Z(O[792]) );
  ANDN U233 ( .B(A[791]), .A(S), .Z(O[791]) );
  ANDN U234 ( .B(A[790]), .A(S), .Z(O[790]) );
  ANDN U235 ( .B(A[78]), .A(S), .Z(O[78]) );
  ANDN U236 ( .B(A[789]), .A(S), .Z(O[789]) );
  ANDN U237 ( .B(A[788]), .A(S), .Z(O[788]) );
  ANDN U238 ( .B(A[787]), .A(S), .Z(O[787]) );
  ANDN U239 ( .B(A[786]), .A(S), .Z(O[786]) );
  ANDN U240 ( .B(A[785]), .A(S), .Z(O[785]) );
  ANDN U241 ( .B(A[784]), .A(S), .Z(O[784]) );
  ANDN U242 ( .B(A[783]), .A(S), .Z(O[783]) );
  ANDN U243 ( .B(A[782]), .A(S), .Z(O[782]) );
  ANDN U244 ( .B(A[781]), .A(S), .Z(O[781]) );
  ANDN U245 ( .B(A[780]), .A(S), .Z(O[780]) );
  ANDN U246 ( .B(A[77]), .A(S), .Z(O[77]) );
  ANDN U247 ( .B(A[779]), .A(S), .Z(O[779]) );
  ANDN U248 ( .B(A[778]), .A(S), .Z(O[778]) );
  ANDN U249 ( .B(A[777]), .A(S), .Z(O[777]) );
  ANDN U250 ( .B(A[776]), .A(S), .Z(O[776]) );
  ANDN U251 ( .B(A[775]), .A(S), .Z(O[775]) );
  ANDN U252 ( .B(A[774]), .A(S), .Z(O[774]) );
  ANDN U253 ( .B(A[773]), .A(S), .Z(O[773]) );
  ANDN U254 ( .B(A[772]), .A(S), .Z(O[772]) );
  ANDN U255 ( .B(A[771]), .A(S), .Z(O[771]) );
  ANDN U256 ( .B(A[770]), .A(S), .Z(O[770]) );
  ANDN U257 ( .B(A[76]), .A(S), .Z(O[76]) );
  ANDN U258 ( .B(A[769]), .A(S), .Z(O[769]) );
  ANDN U259 ( .B(A[768]), .A(S), .Z(O[768]) );
  ANDN U260 ( .B(A[767]), .A(S), .Z(O[767]) );
  ANDN U261 ( .B(A[766]), .A(S), .Z(O[766]) );
  ANDN U262 ( .B(A[765]), .A(S), .Z(O[765]) );
  ANDN U263 ( .B(A[764]), .A(S), .Z(O[764]) );
  ANDN U264 ( .B(A[763]), .A(S), .Z(O[763]) );
  ANDN U265 ( .B(A[762]), .A(S), .Z(O[762]) );
  ANDN U266 ( .B(A[761]), .A(S), .Z(O[761]) );
  ANDN U267 ( .B(A[760]), .A(S), .Z(O[760]) );
  ANDN U268 ( .B(A[75]), .A(S), .Z(O[75]) );
  ANDN U269 ( .B(A[759]), .A(S), .Z(O[759]) );
  ANDN U270 ( .B(A[758]), .A(S), .Z(O[758]) );
  ANDN U271 ( .B(A[757]), .A(S), .Z(O[757]) );
  ANDN U272 ( .B(A[756]), .A(S), .Z(O[756]) );
  ANDN U273 ( .B(A[755]), .A(S), .Z(O[755]) );
  ANDN U274 ( .B(A[754]), .A(S), .Z(O[754]) );
  ANDN U275 ( .B(A[753]), .A(S), .Z(O[753]) );
  ANDN U276 ( .B(A[752]), .A(S), .Z(O[752]) );
  ANDN U277 ( .B(A[751]), .A(S), .Z(O[751]) );
  ANDN U278 ( .B(A[750]), .A(S), .Z(O[750]) );
  ANDN U279 ( .B(A[74]), .A(S), .Z(O[74]) );
  ANDN U280 ( .B(A[749]), .A(S), .Z(O[749]) );
  ANDN U281 ( .B(A[748]), .A(S), .Z(O[748]) );
  ANDN U282 ( .B(A[747]), .A(S), .Z(O[747]) );
  ANDN U283 ( .B(A[746]), .A(S), .Z(O[746]) );
  ANDN U284 ( .B(A[745]), .A(S), .Z(O[745]) );
  ANDN U285 ( .B(A[744]), .A(S), .Z(O[744]) );
  ANDN U286 ( .B(A[743]), .A(S), .Z(O[743]) );
  ANDN U287 ( .B(A[742]), .A(S), .Z(O[742]) );
  ANDN U288 ( .B(A[741]), .A(S), .Z(O[741]) );
  ANDN U289 ( .B(A[740]), .A(S), .Z(O[740]) );
  ANDN U290 ( .B(A[73]), .A(S), .Z(O[73]) );
  ANDN U291 ( .B(A[739]), .A(S), .Z(O[739]) );
  ANDN U292 ( .B(A[738]), .A(S), .Z(O[738]) );
  ANDN U293 ( .B(A[737]), .A(S), .Z(O[737]) );
  ANDN U294 ( .B(A[736]), .A(S), .Z(O[736]) );
  ANDN U295 ( .B(A[735]), .A(S), .Z(O[735]) );
  ANDN U296 ( .B(A[734]), .A(S), .Z(O[734]) );
  ANDN U297 ( .B(A[733]), .A(S), .Z(O[733]) );
  ANDN U298 ( .B(A[732]), .A(S), .Z(O[732]) );
  ANDN U299 ( .B(A[731]), .A(S), .Z(O[731]) );
  ANDN U300 ( .B(A[730]), .A(S), .Z(O[730]) );
  ANDN U301 ( .B(A[72]), .A(S), .Z(O[72]) );
  ANDN U302 ( .B(A[729]), .A(S), .Z(O[729]) );
  ANDN U303 ( .B(A[728]), .A(S), .Z(O[728]) );
  ANDN U304 ( .B(A[727]), .A(S), .Z(O[727]) );
  ANDN U305 ( .B(A[726]), .A(S), .Z(O[726]) );
  ANDN U306 ( .B(A[725]), .A(S), .Z(O[725]) );
  ANDN U307 ( .B(A[724]), .A(S), .Z(O[724]) );
  ANDN U308 ( .B(A[723]), .A(S), .Z(O[723]) );
  ANDN U309 ( .B(A[722]), .A(S), .Z(O[722]) );
  ANDN U310 ( .B(A[721]), .A(S), .Z(O[721]) );
  ANDN U311 ( .B(A[720]), .A(S), .Z(O[720]) );
  ANDN U312 ( .B(A[71]), .A(S), .Z(O[71]) );
  ANDN U313 ( .B(A[719]), .A(S), .Z(O[719]) );
  ANDN U314 ( .B(A[718]), .A(S), .Z(O[718]) );
  ANDN U315 ( .B(A[717]), .A(S), .Z(O[717]) );
  ANDN U316 ( .B(A[716]), .A(S), .Z(O[716]) );
  ANDN U317 ( .B(A[715]), .A(S), .Z(O[715]) );
  ANDN U318 ( .B(A[714]), .A(S), .Z(O[714]) );
  ANDN U319 ( .B(A[713]), .A(S), .Z(O[713]) );
  ANDN U320 ( .B(A[712]), .A(S), .Z(O[712]) );
  ANDN U321 ( .B(A[711]), .A(S), .Z(O[711]) );
  ANDN U322 ( .B(A[710]), .A(S), .Z(O[710]) );
  ANDN U323 ( .B(A[70]), .A(S), .Z(O[70]) );
  ANDN U324 ( .B(A[709]), .A(S), .Z(O[709]) );
  ANDN U325 ( .B(A[708]), .A(S), .Z(O[708]) );
  ANDN U326 ( .B(A[707]), .A(S), .Z(O[707]) );
  ANDN U327 ( .B(A[706]), .A(S), .Z(O[706]) );
  ANDN U328 ( .B(A[705]), .A(S), .Z(O[705]) );
  ANDN U329 ( .B(A[704]), .A(S), .Z(O[704]) );
  ANDN U330 ( .B(A[703]), .A(S), .Z(O[703]) );
  ANDN U331 ( .B(A[702]), .A(S), .Z(O[702]) );
  ANDN U332 ( .B(A[701]), .A(S), .Z(O[701]) );
  ANDN U333 ( .B(A[700]), .A(S), .Z(O[700]) );
  ANDN U334 ( .B(A[6]), .A(S), .Z(O[6]) );
  ANDN U335 ( .B(A[69]), .A(S), .Z(O[69]) );
  ANDN U336 ( .B(A[699]), .A(S), .Z(O[699]) );
  ANDN U337 ( .B(A[698]), .A(S), .Z(O[698]) );
  ANDN U338 ( .B(A[697]), .A(S), .Z(O[697]) );
  ANDN U339 ( .B(A[696]), .A(S), .Z(O[696]) );
  ANDN U340 ( .B(A[695]), .A(S), .Z(O[695]) );
  ANDN U341 ( .B(A[694]), .A(S), .Z(O[694]) );
  ANDN U342 ( .B(A[693]), .A(S), .Z(O[693]) );
  ANDN U343 ( .B(A[692]), .A(S), .Z(O[692]) );
  ANDN U344 ( .B(A[691]), .A(S), .Z(O[691]) );
  ANDN U345 ( .B(A[690]), .A(S), .Z(O[690]) );
  ANDN U346 ( .B(A[68]), .A(S), .Z(O[68]) );
  ANDN U347 ( .B(A[689]), .A(S), .Z(O[689]) );
  ANDN U348 ( .B(A[688]), .A(S), .Z(O[688]) );
  ANDN U349 ( .B(A[687]), .A(S), .Z(O[687]) );
  ANDN U350 ( .B(A[686]), .A(S), .Z(O[686]) );
  ANDN U351 ( .B(A[685]), .A(S), .Z(O[685]) );
  ANDN U352 ( .B(A[684]), .A(S), .Z(O[684]) );
  ANDN U353 ( .B(A[683]), .A(S), .Z(O[683]) );
  ANDN U354 ( .B(A[682]), .A(S), .Z(O[682]) );
  ANDN U355 ( .B(A[681]), .A(S), .Z(O[681]) );
  ANDN U356 ( .B(A[680]), .A(S), .Z(O[680]) );
  ANDN U357 ( .B(A[67]), .A(S), .Z(O[67]) );
  ANDN U358 ( .B(A[679]), .A(S), .Z(O[679]) );
  ANDN U359 ( .B(A[678]), .A(S), .Z(O[678]) );
  ANDN U360 ( .B(A[677]), .A(S), .Z(O[677]) );
  ANDN U361 ( .B(A[676]), .A(S), .Z(O[676]) );
  ANDN U362 ( .B(A[675]), .A(S), .Z(O[675]) );
  ANDN U363 ( .B(A[674]), .A(S), .Z(O[674]) );
  ANDN U364 ( .B(A[673]), .A(S), .Z(O[673]) );
  ANDN U365 ( .B(A[672]), .A(S), .Z(O[672]) );
  ANDN U366 ( .B(A[671]), .A(S), .Z(O[671]) );
  ANDN U367 ( .B(A[670]), .A(S), .Z(O[670]) );
  ANDN U368 ( .B(A[66]), .A(S), .Z(O[66]) );
  ANDN U369 ( .B(A[669]), .A(S), .Z(O[669]) );
  ANDN U370 ( .B(A[668]), .A(S), .Z(O[668]) );
  ANDN U371 ( .B(A[667]), .A(S), .Z(O[667]) );
  ANDN U372 ( .B(A[666]), .A(S), .Z(O[666]) );
  ANDN U373 ( .B(A[665]), .A(S), .Z(O[665]) );
  ANDN U374 ( .B(A[664]), .A(S), .Z(O[664]) );
  ANDN U375 ( .B(A[663]), .A(S), .Z(O[663]) );
  ANDN U376 ( .B(A[662]), .A(S), .Z(O[662]) );
  ANDN U377 ( .B(A[661]), .A(S), .Z(O[661]) );
  ANDN U378 ( .B(A[660]), .A(S), .Z(O[660]) );
  ANDN U379 ( .B(A[65]), .A(S), .Z(O[65]) );
  ANDN U380 ( .B(A[659]), .A(S), .Z(O[659]) );
  ANDN U381 ( .B(A[658]), .A(S), .Z(O[658]) );
  ANDN U382 ( .B(A[657]), .A(S), .Z(O[657]) );
  ANDN U383 ( .B(A[656]), .A(S), .Z(O[656]) );
  ANDN U384 ( .B(A[655]), .A(S), .Z(O[655]) );
  ANDN U385 ( .B(A[654]), .A(S), .Z(O[654]) );
  ANDN U386 ( .B(A[653]), .A(S), .Z(O[653]) );
  ANDN U387 ( .B(A[652]), .A(S), .Z(O[652]) );
  ANDN U388 ( .B(A[651]), .A(S), .Z(O[651]) );
  ANDN U389 ( .B(A[650]), .A(S), .Z(O[650]) );
  ANDN U390 ( .B(A[64]), .A(S), .Z(O[64]) );
  ANDN U391 ( .B(A[649]), .A(S), .Z(O[649]) );
  ANDN U392 ( .B(A[648]), .A(S), .Z(O[648]) );
  ANDN U393 ( .B(A[647]), .A(S), .Z(O[647]) );
  ANDN U394 ( .B(A[646]), .A(S), .Z(O[646]) );
  ANDN U395 ( .B(A[645]), .A(S), .Z(O[645]) );
  ANDN U396 ( .B(A[644]), .A(S), .Z(O[644]) );
  ANDN U397 ( .B(A[643]), .A(S), .Z(O[643]) );
  ANDN U398 ( .B(A[642]), .A(S), .Z(O[642]) );
  ANDN U399 ( .B(A[641]), .A(S), .Z(O[641]) );
  ANDN U400 ( .B(A[640]), .A(S), .Z(O[640]) );
  ANDN U401 ( .B(A[63]), .A(S), .Z(O[63]) );
  ANDN U402 ( .B(A[639]), .A(S), .Z(O[639]) );
  ANDN U403 ( .B(A[638]), .A(S), .Z(O[638]) );
  ANDN U404 ( .B(A[637]), .A(S), .Z(O[637]) );
  ANDN U405 ( .B(A[636]), .A(S), .Z(O[636]) );
  ANDN U406 ( .B(A[635]), .A(S), .Z(O[635]) );
  ANDN U407 ( .B(A[634]), .A(S), .Z(O[634]) );
  ANDN U408 ( .B(A[633]), .A(S), .Z(O[633]) );
  ANDN U409 ( .B(A[632]), .A(S), .Z(O[632]) );
  ANDN U410 ( .B(A[631]), .A(S), .Z(O[631]) );
  ANDN U411 ( .B(A[630]), .A(S), .Z(O[630]) );
  ANDN U412 ( .B(A[62]), .A(S), .Z(O[62]) );
  ANDN U413 ( .B(A[629]), .A(S), .Z(O[629]) );
  ANDN U414 ( .B(A[628]), .A(S), .Z(O[628]) );
  ANDN U415 ( .B(A[627]), .A(S), .Z(O[627]) );
  ANDN U416 ( .B(A[626]), .A(S), .Z(O[626]) );
  ANDN U417 ( .B(A[625]), .A(S), .Z(O[625]) );
  ANDN U418 ( .B(A[624]), .A(S), .Z(O[624]) );
  ANDN U419 ( .B(A[623]), .A(S), .Z(O[623]) );
  ANDN U420 ( .B(A[622]), .A(S), .Z(O[622]) );
  ANDN U421 ( .B(A[621]), .A(S), .Z(O[621]) );
  ANDN U422 ( .B(A[620]), .A(S), .Z(O[620]) );
  ANDN U423 ( .B(A[61]), .A(S), .Z(O[61]) );
  ANDN U424 ( .B(A[619]), .A(S), .Z(O[619]) );
  ANDN U425 ( .B(A[618]), .A(S), .Z(O[618]) );
  ANDN U426 ( .B(A[617]), .A(S), .Z(O[617]) );
  ANDN U427 ( .B(A[616]), .A(S), .Z(O[616]) );
  ANDN U428 ( .B(A[615]), .A(S), .Z(O[615]) );
  ANDN U429 ( .B(A[614]), .A(S), .Z(O[614]) );
  ANDN U430 ( .B(A[613]), .A(S), .Z(O[613]) );
  ANDN U431 ( .B(A[612]), .A(S), .Z(O[612]) );
  ANDN U432 ( .B(A[611]), .A(S), .Z(O[611]) );
  ANDN U433 ( .B(A[610]), .A(S), .Z(O[610]) );
  ANDN U434 ( .B(A[60]), .A(S), .Z(O[60]) );
  ANDN U435 ( .B(A[609]), .A(S), .Z(O[609]) );
  ANDN U436 ( .B(A[608]), .A(S), .Z(O[608]) );
  ANDN U437 ( .B(A[607]), .A(S), .Z(O[607]) );
  ANDN U438 ( .B(A[606]), .A(S), .Z(O[606]) );
  ANDN U439 ( .B(A[605]), .A(S), .Z(O[605]) );
  ANDN U440 ( .B(A[604]), .A(S), .Z(O[604]) );
  ANDN U441 ( .B(A[603]), .A(S), .Z(O[603]) );
  ANDN U442 ( .B(A[602]), .A(S), .Z(O[602]) );
  ANDN U443 ( .B(A[601]), .A(S), .Z(O[601]) );
  ANDN U444 ( .B(A[600]), .A(S), .Z(O[600]) );
  ANDN U445 ( .B(A[5]), .A(S), .Z(O[5]) );
  ANDN U446 ( .B(A[59]), .A(S), .Z(O[59]) );
  ANDN U447 ( .B(A[599]), .A(S), .Z(O[599]) );
  ANDN U448 ( .B(A[598]), .A(S), .Z(O[598]) );
  ANDN U449 ( .B(A[597]), .A(S), .Z(O[597]) );
  ANDN U450 ( .B(A[596]), .A(S), .Z(O[596]) );
  ANDN U451 ( .B(A[595]), .A(S), .Z(O[595]) );
  ANDN U452 ( .B(A[594]), .A(S), .Z(O[594]) );
  ANDN U453 ( .B(A[593]), .A(S), .Z(O[593]) );
  ANDN U454 ( .B(A[592]), .A(S), .Z(O[592]) );
  ANDN U455 ( .B(A[591]), .A(S), .Z(O[591]) );
  ANDN U456 ( .B(A[590]), .A(S), .Z(O[590]) );
  ANDN U457 ( .B(A[58]), .A(S), .Z(O[58]) );
  ANDN U458 ( .B(A[589]), .A(S), .Z(O[589]) );
  ANDN U459 ( .B(A[588]), .A(S), .Z(O[588]) );
  ANDN U460 ( .B(A[587]), .A(S), .Z(O[587]) );
  ANDN U461 ( .B(A[586]), .A(S), .Z(O[586]) );
  ANDN U462 ( .B(A[585]), .A(S), .Z(O[585]) );
  ANDN U463 ( .B(A[584]), .A(S), .Z(O[584]) );
  ANDN U464 ( .B(A[583]), .A(S), .Z(O[583]) );
  ANDN U465 ( .B(A[582]), .A(S), .Z(O[582]) );
  ANDN U466 ( .B(A[581]), .A(S), .Z(O[581]) );
  ANDN U467 ( .B(A[580]), .A(S), .Z(O[580]) );
  ANDN U468 ( .B(A[57]), .A(S), .Z(O[57]) );
  ANDN U469 ( .B(A[579]), .A(S), .Z(O[579]) );
  ANDN U470 ( .B(A[578]), .A(S), .Z(O[578]) );
  ANDN U471 ( .B(A[577]), .A(S), .Z(O[577]) );
  ANDN U472 ( .B(A[576]), .A(S), .Z(O[576]) );
  ANDN U473 ( .B(A[575]), .A(S), .Z(O[575]) );
  ANDN U474 ( .B(A[574]), .A(S), .Z(O[574]) );
  ANDN U475 ( .B(A[573]), .A(S), .Z(O[573]) );
  ANDN U476 ( .B(A[572]), .A(S), .Z(O[572]) );
  ANDN U477 ( .B(A[571]), .A(S), .Z(O[571]) );
  ANDN U478 ( .B(A[570]), .A(S), .Z(O[570]) );
  ANDN U479 ( .B(A[56]), .A(S), .Z(O[56]) );
  ANDN U480 ( .B(A[569]), .A(S), .Z(O[569]) );
  ANDN U481 ( .B(A[568]), .A(S), .Z(O[568]) );
  ANDN U482 ( .B(A[567]), .A(S), .Z(O[567]) );
  ANDN U483 ( .B(A[566]), .A(S), .Z(O[566]) );
  ANDN U484 ( .B(A[565]), .A(S), .Z(O[565]) );
  ANDN U485 ( .B(A[564]), .A(S), .Z(O[564]) );
  ANDN U486 ( .B(A[563]), .A(S), .Z(O[563]) );
  ANDN U487 ( .B(A[562]), .A(S), .Z(O[562]) );
  ANDN U488 ( .B(A[561]), .A(S), .Z(O[561]) );
  ANDN U489 ( .B(A[560]), .A(S), .Z(O[560]) );
  ANDN U490 ( .B(A[55]), .A(S), .Z(O[55]) );
  ANDN U491 ( .B(A[559]), .A(S), .Z(O[559]) );
  ANDN U492 ( .B(A[558]), .A(S), .Z(O[558]) );
  ANDN U493 ( .B(A[557]), .A(S), .Z(O[557]) );
  ANDN U494 ( .B(A[556]), .A(S), .Z(O[556]) );
  ANDN U495 ( .B(A[555]), .A(S), .Z(O[555]) );
  ANDN U496 ( .B(A[554]), .A(S), .Z(O[554]) );
  ANDN U497 ( .B(A[553]), .A(S), .Z(O[553]) );
  ANDN U498 ( .B(A[552]), .A(S), .Z(O[552]) );
  ANDN U499 ( .B(A[551]), .A(S), .Z(O[551]) );
  ANDN U500 ( .B(A[550]), .A(S), .Z(O[550]) );
  ANDN U501 ( .B(A[54]), .A(S), .Z(O[54]) );
  ANDN U502 ( .B(A[549]), .A(S), .Z(O[549]) );
  ANDN U503 ( .B(A[548]), .A(S), .Z(O[548]) );
  ANDN U504 ( .B(A[547]), .A(S), .Z(O[547]) );
  ANDN U505 ( .B(A[546]), .A(S), .Z(O[546]) );
  ANDN U506 ( .B(A[545]), .A(S), .Z(O[545]) );
  ANDN U507 ( .B(A[544]), .A(S), .Z(O[544]) );
  ANDN U508 ( .B(A[543]), .A(S), .Z(O[543]) );
  ANDN U509 ( .B(A[542]), .A(S), .Z(O[542]) );
  ANDN U510 ( .B(A[541]), .A(S), .Z(O[541]) );
  ANDN U511 ( .B(A[540]), .A(S), .Z(O[540]) );
  ANDN U512 ( .B(A[53]), .A(S), .Z(O[53]) );
  ANDN U513 ( .B(A[539]), .A(S), .Z(O[539]) );
  ANDN U514 ( .B(A[538]), .A(S), .Z(O[538]) );
  ANDN U515 ( .B(A[537]), .A(S), .Z(O[537]) );
  ANDN U516 ( .B(A[536]), .A(S), .Z(O[536]) );
  ANDN U517 ( .B(A[535]), .A(S), .Z(O[535]) );
  ANDN U518 ( .B(A[534]), .A(S), .Z(O[534]) );
  ANDN U519 ( .B(A[533]), .A(S), .Z(O[533]) );
  ANDN U520 ( .B(A[532]), .A(S), .Z(O[532]) );
  ANDN U521 ( .B(A[531]), .A(S), .Z(O[531]) );
  ANDN U522 ( .B(A[530]), .A(S), .Z(O[530]) );
  ANDN U523 ( .B(A[52]), .A(S), .Z(O[52]) );
  ANDN U524 ( .B(A[529]), .A(S), .Z(O[529]) );
  ANDN U525 ( .B(A[528]), .A(S), .Z(O[528]) );
  ANDN U526 ( .B(A[527]), .A(S), .Z(O[527]) );
  ANDN U527 ( .B(A[526]), .A(S), .Z(O[526]) );
  ANDN U528 ( .B(A[525]), .A(S), .Z(O[525]) );
  ANDN U529 ( .B(A[524]), .A(S), .Z(O[524]) );
  ANDN U530 ( .B(A[523]), .A(S), .Z(O[523]) );
  ANDN U531 ( .B(A[522]), .A(S), .Z(O[522]) );
  ANDN U532 ( .B(A[521]), .A(S), .Z(O[521]) );
  ANDN U533 ( .B(A[520]), .A(S), .Z(O[520]) );
  ANDN U534 ( .B(A[51]), .A(S), .Z(O[51]) );
  ANDN U535 ( .B(A[519]), .A(S), .Z(O[519]) );
  ANDN U536 ( .B(A[518]), .A(S), .Z(O[518]) );
  ANDN U537 ( .B(A[517]), .A(S), .Z(O[517]) );
  ANDN U538 ( .B(A[516]), .A(S), .Z(O[516]) );
  ANDN U539 ( .B(A[515]), .A(S), .Z(O[515]) );
  ANDN U540 ( .B(A[514]), .A(S), .Z(O[514]) );
  ANDN U541 ( .B(A[513]), .A(S), .Z(O[513]) );
  ANDN U542 ( .B(A[512]), .A(S), .Z(O[512]) );
  ANDN U543 ( .B(A[511]), .A(S), .Z(O[511]) );
  ANDN U544 ( .B(A[510]), .A(S), .Z(O[510]) );
  ANDN U545 ( .B(A[50]), .A(S), .Z(O[50]) );
  ANDN U546 ( .B(A[509]), .A(S), .Z(O[509]) );
  ANDN U547 ( .B(A[508]), .A(S), .Z(O[508]) );
  ANDN U548 ( .B(A[507]), .A(S), .Z(O[507]) );
  ANDN U549 ( .B(A[506]), .A(S), .Z(O[506]) );
  ANDN U550 ( .B(A[505]), .A(S), .Z(O[505]) );
  ANDN U551 ( .B(A[504]), .A(S), .Z(O[504]) );
  ANDN U552 ( .B(A[503]), .A(S), .Z(O[503]) );
  ANDN U553 ( .B(A[502]), .A(S), .Z(O[502]) );
  ANDN U554 ( .B(A[501]), .A(S), .Z(O[501]) );
  ANDN U555 ( .B(A[500]), .A(S), .Z(O[500]) );
  ANDN U556 ( .B(A[4]), .A(S), .Z(O[4]) );
  ANDN U557 ( .B(A[49]), .A(S), .Z(O[49]) );
  ANDN U558 ( .B(A[499]), .A(S), .Z(O[499]) );
  ANDN U559 ( .B(A[498]), .A(S), .Z(O[498]) );
  ANDN U560 ( .B(A[497]), .A(S), .Z(O[497]) );
  ANDN U561 ( .B(A[496]), .A(S), .Z(O[496]) );
  ANDN U562 ( .B(A[495]), .A(S), .Z(O[495]) );
  ANDN U563 ( .B(A[494]), .A(S), .Z(O[494]) );
  ANDN U564 ( .B(A[493]), .A(S), .Z(O[493]) );
  ANDN U565 ( .B(A[492]), .A(S), .Z(O[492]) );
  ANDN U566 ( .B(A[491]), .A(S), .Z(O[491]) );
  ANDN U567 ( .B(A[490]), .A(S), .Z(O[490]) );
  ANDN U568 ( .B(A[48]), .A(S), .Z(O[48]) );
  ANDN U569 ( .B(A[489]), .A(S), .Z(O[489]) );
  ANDN U570 ( .B(A[488]), .A(S), .Z(O[488]) );
  ANDN U571 ( .B(A[487]), .A(S), .Z(O[487]) );
  ANDN U572 ( .B(A[486]), .A(S), .Z(O[486]) );
  ANDN U573 ( .B(A[485]), .A(S), .Z(O[485]) );
  ANDN U574 ( .B(A[484]), .A(S), .Z(O[484]) );
  ANDN U575 ( .B(A[483]), .A(S), .Z(O[483]) );
  ANDN U576 ( .B(A[482]), .A(S), .Z(O[482]) );
  ANDN U577 ( .B(A[481]), .A(S), .Z(O[481]) );
  ANDN U578 ( .B(A[480]), .A(S), .Z(O[480]) );
  ANDN U579 ( .B(A[47]), .A(S), .Z(O[47]) );
  ANDN U580 ( .B(A[479]), .A(S), .Z(O[479]) );
  ANDN U581 ( .B(A[478]), .A(S), .Z(O[478]) );
  ANDN U582 ( .B(A[477]), .A(S), .Z(O[477]) );
  ANDN U583 ( .B(A[476]), .A(S), .Z(O[476]) );
  ANDN U584 ( .B(A[475]), .A(S), .Z(O[475]) );
  ANDN U585 ( .B(A[474]), .A(S), .Z(O[474]) );
  ANDN U586 ( .B(A[473]), .A(S), .Z(O[473]) );
  ANDN U587 ( .B(A[472]), .A(S), .Z(O[472]) );
  ANDN U588 ( .B(A[471]), .A(S), .Z(O[471]) );
  ANDN U589 ( .B(A[470]), .A(S), .Z(O[470]) );
  ANDN U590 ( .B(A[46]), .A(S), .Z(O[46]) );
  ANDN U591 ( .B(A[469]), .A(S), .Z(O[469]) );
  ANDN U592 ( .B(A[468]), .A(S), .Z(O[468]) );
  ANDN U593 ( .B(A[467]), .A(S), .Z(O[467]) );
  ANDN U594 ( .B(A[466]), .A(S), .Z(O[466]) );
  ANDN U595 ( .B(A[465]), .A(S), .Z(O[465]) );
  ANDN U596 ( .B(A[464]), .A(S), .Z(O[464]) );
  ANDN U597 ( .B(A[463]), .A(S), .Z(O[463]) );
  ANDN U598 ( .B(A[462]), .A(S), .Z(O[462]) );
  ANDN U599 ( .B(A[461]), .A(S), .Z(O[461]) );
  ANDN U600 ( .B(A[460]), .A(S), .Z(O[460]) );
  ANDN U601 ( .B(A[45]), .A(S), .Z(O[45]) );
  ANDN U602 ( .B(A[459]), .A(S), .Z(O[459]) );
  ANDN U603 ( .B(A[458]), .A(S), .Z(O[458]) );
  ANDN U604 ( .B(A[457]), .A(S), .Z(O[457]) );
  ANDN U605 ( .B(A[456]), .A(S), .Z(O[456]) );
  ANDN U606 ( .B(A[455]), .A(S), .Z(O[455]) );
  ANDN U607 ( .B(A[454]), .A(S), .Z(O[454]) );
  ANDN U608 ( .B(A[453]), .A(S), .Z(O[453]) );
  ANDN U609 ( .B(A[452]), .A(S), .Z(O[452]) );
  ANDN U610 ( .B(A[451]), .A(S), .Z(O[451]) );
  ANDN U611 ( .B(A[450]), .A(S), .Z(O[450]) );
  ANDN U612 ( .B(A[44]), .A(S), .Z(O[44]) );
  ANDN U613 ( .B(A[449]), .A(S), .Z(O[449]) );
  ANDN U614 ( .B(A[448]), .A(S), .Z(O[448]) );
  ANDN U615 ( .B(A[447]), .A(S), .Z(O[447]) );
  ANDN U616 ( .B(A[446]), .A(S), .Z(O[446]) );
  ANDN U617 ( .B(A[445]), .A(S), .Z(O[445]) );
  ANDN U618 ( .B(A[444]), .A(S), .Z(O[444]) );
  ANDN U619 ( .B(A[443]), .A(S), .Z(O[443]) );
  ANDN U620 ( .B(A[442]), .A(S), .Z(O[442]) );
  ANDN U621 ( .B(A[441]), .A(S), .Z(O[441]) );
  ANDN U622 ( .B(A[440]), .A(S), .Z(O[440]) );
  ANDN U623 ( .B(A[43]), .A(S), .Z(O[43]) );
  ANDN U624 ( .B(A[439]), .A(S), .Z(O[439]) );
  ANDN U625 ( .B(A[438]), .A(S), .Z(O[438]) );
  ANDN U626 ( .B(A[437]), .A(S), .Z(O[437]) );
  ANDN U627 ( .B(A[436]), .A(S), .Z(O[436]) );
  ANDN U628 ( .B(A[435]), .A(S), .Z(O[435]) );
  ANDN U629 ( .B(A[434]), .A(S), .Z(O[434]) );
  ANDN U630 ( .B(A[433]), .A(S), .Z(O[433]) );
  ANDN U631 ( .B(A[432]), .A(S), .Z(O[432]) );
  ANDN U632 ( .B(A[431]), .A(S), .Z(O[431]) );
  ANDN U633 ( .B(A[430]), .A(S), .Z(O[430]) );
  ANDN U634 ( .B(A[42]), .A(S), .Z(O[42]) );
  ANDN U635 ( .B(A[429]), .A(S), .Z(O[429]) );
  ANDN U636 ( .B(A[428]), .A(S), .Z(O[428]) );
  ANDN U637 ( .B(A[427]), .A(S), .Z(O[427]) );
  ANDN U638 ( .B(A[426]), .A(S), .Z(O[426]) );
  ANDN U639 ( .B(A[425]), .A(S), .Z(O[425]) );
  ANDN U640 ( .B(A[424]), .A(S), .Z(O[424]) );
  ANDN U641 ( .B(A[423]), .A(S), .Z(O[423]) );
  ANDN U642 ( .B(A[422]), .A(S), .Z(O[422]) );
  ANDN U643 ( .B(A[421]), .A(S), .Z(O[421]) );
  ANDN U644 ( .B(A[420]), .A(S), .Z(O[420]) );
  ANDN U645 ( .B(A[41]), .A(S), .Z(O[41]) );
  ANDN U646 ( .B(A[419]), .A(S), .Z(O[419]) );
  ANDN U647 ( .B(A[418]), .A(S), .Z(O[418]) );
  ANDN U648 ( .B(A[417]), .A(S), .Z(O[417]) );
  ANDN U649 ( .B(A[416]), .A(S), .Z(O[416]) );
  ANDN U650 ( .B(A[415]), .A(S), .Z(O[415]) );
  ANDN U651 ( .B(A[414]), .A(S), .Z(O[414]) );
  ANDN U652 ( .B(A[413]), .A(S), .Z(O[413]) );
  ANDN U653 ( .B(A[412]), .A(S), .Z(O[412]) );
  ANDN U654 ( .B(A[411]), .A(S), .Z(O[411]) );
  ANDN U655 ( .B(A[410]), .A(S), .Z(O[410]) );
  ANDN U656 ( .B(A[40]), .A(S), .Z(O[40]) );
  ANDN U657 ( .B(A[409]), .A(S), .Z(O[409]) );
  ANDN U658 ( .B(A[408]), .A(S), .Z(O[408]) );
  ANDN U659 ( .B(A[407]), .A(S), .Z(O[407]) );
  ANDN U660 ( .B(A[406]), .A(S), .Z(O[406]) );
  ANDN U661 ( .B(A[405]), .A(S), .Z(O[405]) );
  ANDN U662 ( .B(A[404]), .A(S), .Z(O[404]) );
  ANDN U663 ( .B(A[403]), .A(S), .Z(O[403]) );
  ANDN U664 ( .B(A[402]), .A(S), .Z(O[402]) );
  ANDN U665 ( .B(A[401]), .A(S), .Z(O[401]) );
  ANDN U666 ( .B(A[400]), .A(S), .Z(O[400]) );
  ANDN U667 ( .B(A[3]), .A(S), .Z(O[3]) );
  ANDN U668 ( .B(A[39]), .A(S), .Z(O[39]) );
  ANDN U669 ( .B(A[399]), .A(S), .Z(O[399]) );
  ANDN U670 ( .B(A[398]), .A(S), .Z(O[398]) );
  ANDN U671 ( .B(A[397]), .A(S), .Z(O[397]) );
  ANDN U672 ( .B(A[396]), .A(S), .Z(O[396]) );
  ANDN U673 ( .B(A[395]), .A(S), .Z(O[395]) );
  ANDN U674 ( .B(A[394]), .A(S), .Z(O[394]) );
  ANDN U675 ( .B(A[393]), .A(S), .Z(O[393]) );
  ANDN U676 ( .B(A[392]), .A(S), .Z(O[392]) );
  ANDN U677 ( .B(A[391]), .A(S), .Z(O[391]) );
  ANDN U678 ( .B(A[390]), .A(S), .Z(O[390]) );
  ANDN U679 ( .B(A[38]), .A(S), .Z(O[38]) );
  ANDN U680 ( .B(A[389]), .A(S), .Z(O[389]) );
  ANDN U681 ( .B(A[388]), .A(S), .Z(O[388]) );
  ANDN U682 ( .B(A[387]), .A(S), .Z(O[387]) );
  ANDN U683 ( .B(A[386]), .A(S), .Z(O[386]) );
  ANDN U684 ( .B(A[385]), .A(S), .Z(O[385]) );
  ANDN U685 ( .B(A[384]), .A(S), .Z(O[384]) );
  ANDN U686 ( .B(A[383]), .A(S), .Z(O[383]) );
  ANDN U687 ( .B(A[382]), .A(S), .Z(O[382]) );
  ANDN U688 ( .B(A[381]), .A(S), .Z(O[381]) );
  ANDN U689 ( .B(A[380]), .A(S), .Z(O[380]) );
  ANDN U690 ( .B(A[37]), .A(S), .Z(O[37]) );
  ANDN U691 ( .B(A[379]), .A(S), .Z(O[379]) );
  ANDN U692 ( .B(A[378]), .A(S), .Z(O[378]) );
  ANDN U693 ( .B(A[377]), .A(S), .Z(O[377]) );
  ANDN U694 ( .B(A[376]), .A(S), .Z(O[376]) );
  ANDN U695 ( .B(A[375]), .A(S), .Z(O[375]) );
  ANDN U696 ( .B(A[374]), .A(S), .Z(O[374]) );
  ANDN U697 ( .B(A[373]), .A(S), .Z(O[373]) );
  ANDN U698 ( .B(A[372]), .A(S), .Z(O[372]) );
  ANDN U699 ( .B(A[371]), .A(S), .Z(O[371]) );
  ANDN U700 ( .B(A[370]), .A(S), .Z(O[370]) );
  ANDN U701 ( .B(A[36]), .A(S), .Z(O[36]) );
  ANDN U702 ( .B(A[369]), .A(S), .Z(O[369]) );
  ANDN U703 ( .B(A[368]), .A(S), .Z(O[368]) );
  ANDN U704 ( .B(A[367]), .A(S), .Z(O[367]) );
  ANDN U705 ( .B(A[366]), .A(S), .Z(O[366]) );
  ANDN U706 ( .B(A[365]), .A(S), .Z(O[365]) );
  ANDN U707 ( .B(A[364]), .A(S), .Z(O[364]) );
  ANDN U708 ( .B(A[363]), .A(S), .Z(O[363]) );
  ANDN U709 ( .B(A[362]), .A(S), .Z(O[362]) );
  ANDN U710 ( .B(A[361]), .A(S), .Z(O[361]) );
  ANDN U711 ( .B(A[360]), .A(S), .Z(O[360]) );
  ANDN U712 ( .B(A[35]), .A(S), .Z(O[35]) );
  ANDN U713 ( .B(A[359]), .A(S), .Z(O[359]) );
  ANDN U714 ( .B(A[358]), .A(S), .Z(O[358]) );
  ANDN U715 ( .B(A[357]), .A(S), .Z(O[357]) );
  ANDN U716 ( .B(A[356]), .A(S), .Z(O[356]) );
  ANDN U717 ( .B(A[355]), .A(S), .Z(O[355]) );
  ANDN U718 ( .B(A[354]), .A(S), .Z(O[354]) );
  ANDN U719 ( .B(A[353]), .A(S), .Z(O[353]) );
  ANDN U720 ( .B(A[352]), .A(S), .Z(O[352]) );
  ANDN U721 ( .B(A[351]), .A(S), .Z(O[351]) );
  ANDN U722 ( .B(A[350]), .A(S), .Z(O[350]) );
  ANDN U723 ( .B(A[34]), .A(S), .Z(O[34]) );
  ANDN U724 ( .B(A[349]), .A(S), .Z(O[349]) );
  ANDN U725 ( .B(A[348]), .A(S), .Z(O[348]) );
  ANDN U726 ( .B(A[347]), .A(S), .Z(O[347]) );
  ANDN U727 ( .B(A[346]), .A(S), .Z(O[346]) );
  ANDN U728 ( .B(A[345]), .A(S), .Z(O[345]) );
  ANDN U729 ( .B(A[344]), .A(S), .Z(O[344]) );
  ANDN U730 ( .B(A[343]), .A(S), .Z(O[343]) );
  ANDN U731 ( .B(A[342]), .A(S), .Z(O[342]) );
  ANDN U732 ( .B(A[341]), .A(S), .Z(O[341]) );
  ANDN U733 ( .B(A[340]), .A(S), .Z(O[340]) );
  ANDN U734 ( .B(A[33]), .A(S), .Z(O[33]) );
  ANDN U735 ( .B(A[339]), .A(S), .Z(O[339]) );
  ANDN U736 ( .B(A[338]), .A(S), .Z(O[338]) );
  ANDN U737 ( .B(A[337]), .A(S), .Z(O[337]) );
  ANDN U738 ( .B(A[336]), .A(S), .Z(O[336]) );
  ANDN U739 ( .B(A[335]), .A(S), .Z(O[335]) );
  ANDN U740 ( .B(A[334]), .A(S), .Z(O[334]) );
  ANDN U741 ( .B(A[333]), .A(S), .Z(O[333]) );
  ANDN U742 ( .B(A[332]), .A(S), .Z(O[332]) );
  ANDN U743 ( .B(A[331]), .A(S), .Z(O[331]) );
  ANDN U744 ( .B(A[330]), .A(S), .Z(O[330]) );
  ANDN U745 ( .B(A[32]), .A(S), .Z(O[32]) );
  ANDN U746 ( .B(A[329]), .A(S), .Z(O[329]) );
  ANDN U747 ( .B(A[328]), .A(S), .Z(O[328]) );
  ANDN U748 ( .B(A[327]), .A(S), .Z(O[327]) );
  ANDN U749 ( .B(A[326]), .A(S), .Z(O[326]) );
  ANDN U750 ( .B(A[325]), .A(S), .Z(O[325]) );
  ANDN U751 ( .B(A[324]), .A(S), .Z(O[324]) );
  ANDN U752 ( .B(A[323]), .A(S), .Z(O[323]) );
  ANDN U753 ( .B(A[322]), .A(S), .Z(O[322]) );
  ANDN U754 ( .B(A[321]), .A(S), .Z(O[321]) );
  ANDN U755 ( .B(A[320]), .A(S), .Z(O[320]) );
  ANDN U756 ( .B(A[31]), .A(S), .Z(O[31]) );
  ANDN U757 ( .B(A[319]), .A(S), .Z(O[319]) );
  ANDN U758 ( .B(A[318]), .A(S), .Z(O[318]) );
  ANDN U759 ( .B(A[317]), .A(S), .Z(O[317]) );
  ANDN U760 ( .B(A[316]), .A(S), .Z(O[316]) );
  ANDN U761 ( .B(A[315]), .A(S), .Z(O[315]) );
  ANDN U762 ( .B(A[314]), .A(S), .Z(O[314]) );
  ANDN U763 ( .B(A[313]), .A(S), .Z(O[313]) );
  ANDN U764 ( .B(A[312]), .A(S), .Z(O[312]) );
  ANDN U765 ( .B(A[311]), .A(S), .Z(O[311]) );
  ANDN U766 ( .B(A[310]), .A(S), .Z(O[310]) );
  ANDN U767 ( .B(A[30]), .A(S), .Z(O[30]) );
  ANDN U768 ( .B(A[309]), .A(S), .Z(O[309]) );
  ANDN U769 ( .B(A[308]), .A(S), .Z(O[308]) );
  ANDN U770 ( .B(A[307]), .A(S), .Z(O[307]) );
  ANDN U771 ( .B(A[306]), .A(S), .Z(O[306]) );
  ANDN U772 ( .B(A[305]), .A(S), .Z(O[305]) );
  ANDN U773 ( .B(A[304]), .A(S), .Z(O[304]) );
  ANDN U774 ( .B(A[303]), .A(S), .Z(O[303]) );
  ANDN U775 ( .B(A[302]), .A(S), .Z(O[302]) );
  ANDN U776 ( .B(A[301]), .A(S), .Z(O[301]) );
  ANDN U777 ( .B(A[300]), .A(S), .Z(O[300]) );
  ANDN U778 ( .B(A[2]), .A(S), .Z(O[2]) );
  ANDN U779 ( .B(A[29]), .A(S), .Z(O[29]) );
  ANDN U780 ( .B(A[299]), .A(S), .Z(O[299]) );
  ANDN U781 ( .B(A[298]), .A(S), .Z(O[298]) );
  ANDN U782 ( .B(A[297]), .A(S), .Z(O[297]) );
  ANDN U783 ( .B(A[296]), .A(S), .Z(O[296]) );
  ANDN U784 ( .B(A[295]), .A(S), .Z(O[295]) );
  ANDN U785 ( .B(A[294]), .A(S), .Z(O[294]) );
  ANDN U786 ( .B(A[293]), .A(S), .Z(O[293]) );
  ANDN U787 ( .B(A[292]), .A(S), .Z(O[292]) );
  ANDN U788 ( .B(A[291]), .A(S), .Z(O[291]) );
  ANDN U789 ( .B(A[290]), .A(S), .Z(O[290]) );
  ANDN U790 ( .B(A[28]), .A(S), .Z(O[28]) );
  ANDN U791 ( .B(A[289]), .A(S), .Z(O[289]) );
  ANDN U792 ( .B(A[288]), .A(S), .Z(O[288]) );
  ANDN U793 ( .B(A[287]), .A(S), .Z(O[287]) );
  ANDN U794 ( .B(A[286]), .A(S), .Z(O[286]) );
  ANDN U795 ( .B(A[285]), .A(S), .Z(O[285]) );
  ANDN U796 ( .B(A[284]), .A(S), .Z(O[284]) );
  ANDN U797 ( .B(A[283]), .A(S), .Z(O[283]) );
  ANDN U798 ( .B(A[282]), .A(S), .Z(O[282]) );
  ANDN U799 ( .B(A[281]), .A(S), .Z(O[281]) );
  ANDN U800 ( .B(A[280]), .A(S), .Z(O[280]) );
  ANDN U801 ( .B(A[27]), .A(S), .Z(O[27]) );
  ANDN U802 ( .B(A[279]), .A(S), .Z(O[279]) );
  ANDN U803 ( .B(A[278]), .A(S), .Z(O[278]) );
  ANDN U804 ( .B(A[277]), .A(S), .Z(O[277]) );
  ANDN U805 ( .B(A[276]), .A(S), .Z(O[276]) );
  ANDN U806 ( .B(A[275]), .A(S), .Z(O[275]) );
  ANDN U807 ( .B(A[274]), .A(S), .Z(O[274]) );
  ANDN U808 ( .B(A[273]), .A(S), .Z(O[273]) );
  ANDN U809 ( .B(A[272]), .A(S), .Z(O[272]) );
  ANDN U810 ( .B(A[271]), .A(S), .Z(O[271]) );
  ANDN U811 ( .B(A[270]), .A(S), .Z(O[270]) );
  ANDN U812 ( .B(A[26]), .A(S), .Z(O[26]) );
  ANDN U813 ( .B(A[269]), .A(S), .Z(O[269]) );
  ANDN U814 ( .B(A[268]), .A(S), .Z(O[268]) );
  ANDN U815 ( .B(A[267]), .A(S), .Z(O[267]) );
  ANDN U816 ( .B(A[266]), .A(S), .Z(O[266]) );
  ANDN U817 ( .B(A[265]), .A(S), .Z(O[265]) );
  ANDN U818 ( .B(A[264]), .A(S), .Z(O[264]) );
  ANDN U819 ( .B(A[263]), .A(S), .Z(O[263]) );
  ANDN U820 ( .B(A[262]), .A(S), .Z(O[262]) );
  ANDN U821 ( .B(A[261]), .A(S), .Z(O[261]) );
  ANDN U822 ( .B(A[260]), .A(S), .Z(O[260]) );
  ANDN U823 ( .B(A[25]), .A(S), .Z(O[25]) );
  ANDN U824 ( .B(A[259]), .A(S), .Z(O[259]) );
  ANDN U825 ( .B(A[258]), .A(S), .Z(O[258]) );
  ANDN U826 ( .B(A[257]), .A(S), .Z(O[257]) );
  ANDN U827 ( .B(A[256]), .A(S), .Z(O[256]) );
  ANDN U828 ( .B(A[255]), .A(S), .Z(O[255]) );
  ANDN U829 ( .B(A[254]), .A(S), .Z(O[254]) );
  ANDN U830 ( .B(A[253]), .A(S), .Z(O[253]) );
  ANDN U831 ( .B(A[252]), .A(S), .Z(O[252]) );
  ANDN U832 ( .B(A[251]), .A(S), .Z(O[251]) );
  ANDN U833 ( .B(A[250]), .A(S), .Z(O[250]) );
  ANDN U834 ( .B(A[24]), .A(S), .Z(O[24]) );
  ANDN U835 ( .B(A[249]), .A(S), .Z(O[249]) );
  ANDN U836 ( .B(A[248]), .A(S), .Z(O[248]) );
  ANDN U837 ( .B(A[247]), .A(S), .Z(O[247]) );
  ANDN U838 ( .B(A[246]), .A(S), .Z(O[246]) );
  ANDN U839 ( .B(A[245]), .A(S), .Z(O[245]) );
  ANDN U840 ( .B(A[244]), .A(S), .Z(O[244]) );
  ANDN U841 ( .B(A[243]), .A(S), .Z(O[243]) );
  ANDN U842 ( .B(A[242]), .A(S), .Z(O[242]) );
  ANDN U843 ( .B(A[241]), .A(S), .Z(O[241]) );
  ANDN U844 ( .B(A[240]), .A(S), .Z(O[240]) );
  ANDN U845 ( .B(A[23]), .A(S), .Z(O[23]) );
  ANDN U846 ( .B(A[239]), .A(S), .Z(O[239]) );
  ANDN U847 ( .B(A[238]), .A(S), .Z(O[238]) );
  ANDN U848 ( .B(A[237]), .A(S), .Z(O[237]) );
  ANDN U849 ( .B(A[236]), .A(S), .Z(O[236]) );
  ANDN U850 ( .B(A[235]), .A(S), .Z(O[235]) );
  ANDN U851 ( .B(A[234]), .A(S), .Z(O[234]) );
  ANDN U852 ( .B(A[233]), .A(S), .Z(O[233]) );
  ANDN U853 ( .B(A[232]), .A(S), .Z(O[232]) );
  ANDN U854 ( .B(A[231]), .A(S), .Z(O[231]) );
  ANDN U855 ( .B(A[230]), .A(S), .Z(O[230]) );
  ANDN U856 ( .B(A[22]), .A(S), .Z(O[22]) );
  ANDN U857 ( .B(A[229]), .A(S), .Z(O[229]) );
  ANDN U858 ( .B(A[228]), .A(S), .Z(O[228]) );
  ANDN U859 ( .B(A[227]), .A(S), .Z(O[227]) );
  ANDN U860 ( .B(A[226]), .A(S), .Z(O[226]) );
  ANDN U861 ( .B(A[225]), .A(S), .Z(O[225]) );
  ANDN U862 ( .B(A[224]), .A(S), .Z(O[224]) );
  ANDN U863 ( .B(A[223]), .A(S), .Z(O[223]) );
  ANDN U864 ( .B(A[222]), .A(S), .Z(O[222]) );
  ANDN U865 ( .B(A[221]), .A(S), .Z(O[221]) );
  ANDN U866 ( .B(A[220]), .A(S), .Z(O[220]) );
  ANDN U867 ( .B(A[21]), .A(S), .Z(O[21]) );
  ANDN U868 ( .B(A[219]), .A(S), .Z(O[219]) );
  ANDN U869 ( .B(A[218]), .A(S), .Z(O[218]) );
  ANDN U870 ( .B(A[217]), .A(S), .Z(O[217]) );
  ANDN U871 ( .B(A[216]), .A(S), .Z(O[216]) );
  ANDN U872 ( .B(A[215]), .A(S), .Z(O[215]) );
  ANDN U873 ( .B(A[214]), .A(S), .Z(O[214]) );
  ANDN U874 ( .B(A[213]), .A(S), .Z(O[213]) );
  ANDN U875 ( .B(A[212]), .A(S), .Z(O[212]) );
  ANDN U876 ( .B(A[211]), .A(S), .Z(O[211]) );
  ANDN U877 ( .B(A[210]), .A(S), .Z(O[210]) );
  ANDN U878 ( .B(A[20]), .A(S), .Z(O[20]) );
  ANDN U879 ( .B(A[209]), .A(S), .Z(O[209]) );
  ANDN U880 ( .B(A[208]), .A(S), .Z(O[208]) );
  ANDN U881 ( .B(A[207]), .A(S), .Z(O[207]) );
  ANDN U882 ( .B(A[206]), .A(S), .Z(O[206]) );
  ANDN U883 ( .B(A[205]), .A(S), .Z(O[205]) );
  ANDN U884 ( .B(A[204]), .A(S), .Z(O[204]) );
  ANDN U885 ( .B(A[203]), .A(S), .Z(O[203]) );
  ANDN U886 ( .B(A[202]), .A(S), .Z(O[202]) );
  ANDN U887 ( .B(A[201]), .A(S), .Z(O[201]) );
  ANDN U888 ( .B(A[200]), .A(S), .Z(O[200]) );
  ANDN U889 ( .B(A[1]), .A(S), .Z(O[1]) );
  ANDN U890 ( .B(A[19]), .A(S), .Z(O[19]) );
  ANDN U891 ( .B(A[199]), .A(S), .Z(O[199]) );
  ANDN U892 ( .B(A[198]), .A(S), .Z(O[198]) );
  ANDN U893 ( .B(A[197]), .A(S), .Z(O[197]) );
  ANDN U894 ( .B(A[196]), .A(S), .Z(O[196]) );
  ANDN U895 ( .B(A[195]), .A(S), .Z(O[195]) );
  ANDN U896 ( .B(A[194]), .A(S), .Z(O[194]) );
  ANDN U897 ( .B(A[193]), .A(S), .Z(O[193]) );
  ANDN U898 ( .B(A[192]), .A(S), .Z(O[192]) );
  ANDN U899 ( .B(A[191]), .A(S), .Z(O[191]) );
  ANDN U900 ( .B(A[190]), .A(S), .Z(O[190]) );
  ANDN U901 ( .B(A[18]), .A(S), .Z(O[18]) );
  ANDN U902 ( .B(A[189]), .A(S), .Z(O[189]) );
  ANDN U903 ( .B(A[188]), .A(S), .Z(O[188]) );
  ANDN U904 ( .B(A[187]), .A(S), .Z(O[187]) );
  ANDN U905 ( .B(A[186]), .A(S), .Z(O[186]) );
  ANDN U906 ( .B(A[185]), .A(S), .Z(O[185]) );
  ANDN U907 ( .B(A[184]), .A(S), .Z(O[184]) );
  ANDN U908 ( .B(A[183]), .A(S), .Z(O[183]) );
  ANDN U909 ( .B(A[182]), .A(S), .Z(O[182]) );
  ANDN U910 ( .B(A[181]), .A(S), .Z(O[181]) );
  ANDN U911 ( .B(A[180]), .A(S), .Z(O[180]) );
  ANDN U912 ( .B(A[17]), .A(S), .Z(O[17]) );
  ANDN U913 ( .B(A[179]), .A(S), .Z(O[179]) );
  ANDN U914 ( .B(A[178]), .A(S), .Z(O[178]) );
  ANDN U915 ( .B(A[177]), .A(S), .Z(O[177]) );
  ANDN U916 ( .B(A[176]), .A(S), .Z(O[176]) );
  ANDN U917 ( .B(A[175]), .A(S), .Z(O[175]) );
  ANDN U918 ( .B(A[174]), .A(S), .Z(O[174]) );
  ANDN U919 ( .B(A[173]), .A(S), .Z(O[173]) );
  ANDN U920 ( .B(A[172]), .A(S), .Z(O[172]) );
  ANDN U921 ( .B(A[171]), .A(S), .Z(O[171]) );
  ANDN U922 ( .B(A[170]), .A(S), .Z(O[170]) );
  ANDN U923 ( .B(A[16]), .A(S), .Z(O[16]) );
  ANDN U924 ( .B(A[169]), .A(S), .Z(O[169]) );
  ANDN U925 ( .B(A[168]), .A(S), .Z(O[168]) );
  ANDN U926 ( .B(A[167]), .A(S), .Z(O[167]) );
  ANDN U927 ( .B(A[166]), .A(S), .Z(O[166]) );
  ANDN U928 ( .B(A[165]), .A(S), .Z(O[165]) );
  ANDN U929 ( .B(A[164]), .A(S), .Z(O[164]) );
  ANDN U930 ( .B(A[163]), .A(S), .Z(O[163]) );
  ANDN U931 ( .B(A[162]), .A(S), .Z(O[162]) );
  ANDN U932 ( .B(A[161]), .A(S), .Z(O[161]) );
  ANDN U933 ( .B(A[160]), .A(S), .Z(O[160]) );
  ANDN U934 ( .B(A[15]), .A(S), .Z(O[15]) );
  ANDN U935 ( .B(A[159]), .A(S), .Z(O[159]) );
  ANDN U936 ( .B(A[158]), .A(S), .Z(O[158]) );
  ANDN U937 ( .B(A[157]), .A(S), .Z(O[157]) );
  ANDN U938 ( .B(A[156]), .A(S), .Z(O[156]) );
  ANDN U939 ( .B(A[155]), .A(S), .Z(O[155]) );
  ANDN U940 ( .B(A[154]), .A(S), .Z(O[154]) );
  ANDN U941 ( .B(A[153]), .A(S), .Z(O[153]) );
  ANDN U942 ( .B(A[152]), .A(S), .Z(O[152]) );
  ANDN U943 ( .B(A[151]), .A(S), .Z(O[151]) );
  ANDN U944 ( .B(A[150]), .A(S), .Z(O[150]) );
  ANDN U945 ( .B(A[14]), .A(S), .Z(O[14]) );
  ANDN U946 ( .B(A[149]), .A(S), .Z(O[149]) );
  ANDN U947 ( .B(A[148]), .A(S), .Z(O[148]) );
  ANDN U948 ( .B(A[147]), .A(S), .Z(O[147]) );
  ANDN U949 ( .B(A[146]), .A(S), .Z(O[146]) );
  ANDN U950 ( .B(A[145]), .A(S), .Z(O[145]) );
  ANDN U951 ( .B(A[144]), .A(S), .Z(O[144]) );
  ANDN U952 ( .B(A[143]), .A(S), .Z(O[143]) );
  ANDN U953 ( .B(A[142]), .A(S), .Z(O[142]) );
  ANDN U954 ( .B(A[141]), .A(S), .Z(O[141]) );
  ANDN U955 ( .B(A[140]), .A(S), .Z(O[140]) );
  ANDN U956 ( .B(A[13]), .A(S), .Z(O[13]) );
  ANDN U957 ( .B(A[139]), .A(S), .Z(O[139]) );
  ANDN U958 ( .B(A[138]), .A(S), .Z(O[138]) );
  ANDN U959 ( .B(A[137]), .A(S), .Z(O[137]) );
  ANDN U960 ( .B(A[136]), .A(S), .Z(O[136]) );
  ANDN U961 ( .B(A[135]), .A(S), .Z(O[135]) );
  ANDN U962 ( .B(A[134]), .A(S), .Z(O[134]) );
  ANDN U963 ( .B(A[133]), .A(S), .Z(O[133]) );
  ANDN U964 ( .B(A[132]), .A(S), .Z(O[132]) );
  ANDN U965 ( .B(A[131]), .A(S), .Z(O[131]) );
  ANDN U966 ( .B(A[130]), .A(S), .Z(O[130]) );
  ANDN U967 ( .B(A[12]), .A(S), .Z(O[12]) );
  ANDN U968 ( .B(A[129]), .A(S), .Z(O[129]) );
  ANDN U969 ( .B(A[128]), .A(S), .Z(O[128]) );
  ANDN U970 ( .B(A[127]), .A(S), .Z(O[127]) );
  ANDN U971 ( .B(A[126]), .A(S), .Z(O[126]) );
  ANDN U972 ( .B(A[125]), .A(S), .Z(O[125]) );
  ANDN U973 ( .B(A[124]), .A(S), .Z(O[124]) );
  ANDN U974 ( .B(A[123]), .A(S), .Z(O[123]) );
  ANDN U975 ( .B(A[122]), .A(S), .Z(O[122]) );
  ANDN U976 ( .B(A[121]), .A(S), .Z(O[121]) );
  ANDN U977 ( .B(A[120]), .A(S), .Z(O[120]) );
  ANDN U978 ( .B(A[11]), .A(S), .Z(O[11]) );
  ANDN U979 ( .B(A[119]), .A(S), .Z(O[119]) );
  ANDN U980 ( .B(A[118]), .A(S), .Z(O[118]) );
  ANDN U981 ( .B(A[117]), .A(S), .Z(O[117]) );
  ANDN U982 ( .B(A[116]), .A(S), .Z(O[116]) );
  ANDN U983 ( .B(A[115]), .A(S), .Z(O[115]) );
  ANDN U984 ( .B(A[114]), .A(S), .Z(O[114]) );
  ANDN U985 ( .B(A[113]), .A(S), .Z(O[113]) );
  ANDN U986 ( .B(A[112]), .A(S), .Z(O[112]) );
  ANDN U987 ( .B(A[111]), .A(S), .Z(O[111]) );
  ANDN U988 ( .B(A[110]), .A(S), .Z(O[110]) );
  ANDN U989 ( .B(A[10]), .A(S), .Z(O[10]) );
  ANDN U990 ( .B(A[109]), .A(S), .Z(O[109]) );
  ANDN U991 ( .B(A[108]), .A(S), .Z(O[108]) );
  ANDN U992 ( .B(A[107]), .A(S), .Z(O[107]) );
  ANDN U993 ( .B(A[106]), .A(S), .Z(O[106]) );
  ANDN U994 ( .B(A[105]), .A(S), .Z(O[105]) );
  ANDN U995 ( .B(A[104]), .A(S), .Z(O[104]) );
  ANDN U996 ( .B(A[103]), .A(S), .Z(O[103]) );
  ANDN U997 ( .B(A[102]), .A(S), .Z(O[102]) );
  ANDN U998 ( .B(A[1023]), .A(S), .Z(O[1023]) );
  ANDN U999 ( .B(A[1022]), .A(S), .Z(O[1022]) );
  ANDN U1000 ( .B(A[1021]), .A(S), .Z(O[1021]) );
  ANDN U1001 ( .B(A[1020]), .A(S), .Z(O[1020]) );
  ANDN U1002 ( .B(A[101]), .A(S), .Z(O[101]) );
  ANDN U1003 ( .B(A[1019]), .A(S), .Z(O[1019]) );
  ANDN U1004 ( .B(A[1018]), .A(S), .Z(O[1018]) );
  ANDN U1005 ( .B(A[1017]), .A(S), .Z(O[1017]) );
  ANDN U1006 ( .B(A[1016]), .A(S), .Z(O[1016]) );
  ANDN U1007 ( .B(A[1015]), .A(S), .Z(O[1015]) );
  ANDN U1008 ( .B(A[1014]), .A(S), .Z(O[1014]) );
  ANDN U1009 ( .B(A[1013]), .A(S), .Z(O[1013]) );
  ANDN U1010 ( .B(A[1012]), .A(S), .Z(O[1012]) );
  ANDN U1011 ( .B(A[1011]), .A(S), .Z(O[1011]) );
  ANDN U1012 ( .B(A[1010]), .A(S), .Z(O[1010]) );
  ANDN U1013 ( .B(A[100]), .A(S), .Z(O[100]) );
  ANDN U1014 ( .B(A[1009]), .A(S), .Z(O[1009]) );
  ANDN U1015 ( .B(A[1008]), .A(S), .Z(O[1008]) );
  ANDN U1016 ( .B(A[1007]), .A(S), .Z(O[1007]) );
  ANDN U1017 ( .B(A[1006]), .A(S), .Z(O[1006]) );
  ANDN U1018 ( .B(A[1005]), .A(S), .Z(O[1005]) );
  ANDN U1019 ( .B(A[1004]), .A(S), .Z(O[1004]) );
  ANDN U1020 ( .B(A[1003]), .A(S), .Z(O[1003]) );
  ANDN U1021 ( .B(A[1002]), .A(S), .Z(O[1002]) );
  ANDN U1022 ( .B(A[1001]), .A(S), .Z(O[1001]) );
  ANDN U1023 ( .B(A[1000]), .A(S), .Z(O[1000]) );
  ANDN U1024 ( .B(A[0]), .A(S), .Z(O[0]) );
endmodule


module MUX_N1026_2 ( A, B, S, O );
  input [1025:0] A;
  input [1025:0] B;
  output [1025:0] O;
  input S;


  ANDN U1 ( .B(A[9]), .A(S), .Z(O[9]) );
  ANDN U2 ( .B(A[99]), .A(S), .Z(O[99]) );
  ANDN U3 ( .B(A[999]), .A(S), .Z(O[999]) );
  ANDN U4 ( .B(A[998]), .A(S), .Z(O[998]) );
  ANDN U5 ( .B(A[997]), .A(S), .Z(O[997]) );
  ANDN U6 ( .B(A[996]), .A(S), .Z(O[996]) );
  ANDN U7 ( .B(A[995]), .A(S), .Z(O[995]) );
  ANDN U8 ( .B(A[994]), .A(S), .Z(O[994]) );
  ANDN U9 ( .B(A[993]), .A(S), .Z(O[993]) );
  ANDN U10 ( .B(A[992]), .A(S), .Z(O[992]) );
  ANDN U11 ( .B(A[991]), .A(S), .Z(O[991]) );
  ANDN U12 ( .B(A[990]), .A(S), .Z(O[990]) );
  ANDN U13 ( .B(A[98]), .A(S), .Z(O[98]) );
  ANDN U14 ( .B(A[989]), .A(S), .Z(O[989]) );
  ANDN U15 ( .B(A[988]), .A(S), .Z(O[988]) );
  ANDN U16 ( .B(A[987]), .A(S), .Z(O[987]) );
  ANDN U17 ( .B(A[986]), .A(S), .Z(O[986]) );
  ANDN U18 ( .B(A[985]), .A(S), .Z(O[985]) );
  ANDN U19 ( .B(A[984]), .A(S), .Z(O[984]) );
  ANDN U20 ( .B(A[983]), .A(S), .Z(O[983]) );
  ANDN U21 ( .B(A[982]), .A(S), .Z(O[982]) );
  ANDN U22 ( .B(A[981]), .A(S), .Z(O[981]) );
  ANDN U23 ( .B(A[980]), .A(S), .Z(O[980]) );
  ANDN U24 ( .B(A[97]), .A(S), .Z(O[97]) );
  ANDN U25 ( .B(A[979]), .A(S), .Z(O[979]) );
  ANDN U26 ( .B(A[978]), .A(S), .Z(O[978]) );
  ANDN U27 ( .B(A[977]), .A(S), .Z(O[977]) );
  ANDN U28 ( .B(A[976]), .A(S), .Z(O[976]) );
  ANDN U29 ( .B(A[975]), .A(S), .Z(O[975]) );
  ANDN U30 ( .B(A[974]), .A(S), .Z(O[974]) );
  ANDN U31 ( .B(A[973]), .A(S), .Z(O[973]) );
  ANDN U32 ( .B(A[972]), .A(S), .Z(O[972]) );
  ANDN U33 ( .B(A[971]), .A(S), .Z(O[971]) );
  ANDN U34 ( .B(A[970]), .A(S), .Z(O[970]) );
  ANDN U35 ( .B(A[96]), .A(S), .Z(O[96]) );
  ANDN U36 ( .B(A[969]), .A(S), .Z(O[969]) );
  ANDN U37 ( .B(A[968]), .A(S), .Z(O[968]) );
  ANDN U38 ( .B(A[967]), .A(S), .Z(O[967]) );
  ANDN U39 ( .B(A[966]), .A(S), .Z(O[966]) );
  ANDN U40 ( .B(A[965]), .A(S), .Z(O[965]) );
  ANDN U41 ( .B(A[964]), .A(S), .Z(O[964]) );
  ANDN U42 ( .B(A[963]), .A(S), .Z(O[963]) );
  ANDN U43 ( .B(A[962]), .A(S), .Z(O[962]) );
  ANDN U44 ( .B(A[961]), .A(S), .Z(O[961]) );
  ANDN U45 ( .B(A[960]), .A(S), .Z(O[960]) );
  ANDN U46 ( .B(A[95]), .A(S), .Z(O[95]) );
  ANDN U47 ( .B(A[959]), .A(S), .Z(O[959]) );
  ANDN U48 ( .B(A[958]), .A(S), .Z(O[958]) );
  ANDN U49 ( .B(A[957]), .A(S), .Z(O[957]) );
  ANDN U50 ( .B(A[956]), .A(S), .Z(O[956]) );
  ANDN U51 ( .B(A[955]), .A(S), .Z(O[955]) );
  ANDN U52 ( .B(A[954]), .A(S), .Z(O[954]) );
  ANDN U53 ( .B(A[953]), .A(S), .Z(O[953]) );
  ANDN U54 ( .B(A[952]), .A(S), .Z(O[952]) );
  ANDN U55 ( .B(A[951]), .A(S), .Z(O[951]) );
  ANDN U56 ( .B(A[950]), .A(S), .Z(O[950]) );
  ANDN U57 ( .B(A[94]), .A(S), .Z(O[94]) );
  ANDN U58 ( .B(A[949]), .A(S), .Z(O[949]) );
  ANDN U59 ( .B(A[948]), .A(S), .Z(O[948]) );
  ANDN U60 ( .B(A[947]), .A(S), .Z(O[947]) );
  ANDN U61 ( .B(A[946]), .A(S), .Z(O[946]) );
  ANDN U62 ( .B(A[945]), .A(S), .Z(O[945]) );
  ANDN U63 ( .B(A[944]), .A(S), .Z(O[944]) );
  ANDN U64 ( .B(A[943]), .A(S), .Z(O[943]) );
  ANDN U65 ( .B(A[942]), .A(S), .Z(O[942]) );
  ANDN U66 ( .B(A[941]), .A(S), .Z(O[941]) );
  ANDN U67 ( .B(A[940]), .A(S), .Z(O[940]) );
  ANDN U68 ( .B(A[93]), .A(S), .Z(O[93]) );
  ANDN U69 ( .B(A[939]), .A(S), .Z(O[939]) );
  ANDN U70 ( .B(A[938]), .A(S), .Z(O[938]) );
  ANDN U71 ( .B(A[937]), .A(S), .Z(O[937]) );
  ANDN U72 ( .B(A[936]), .A(S), .Z(O[936]) );
  ANDN U73 ( .B(A[935]), .A(S), .Z(O[935]) );
  ANDN U74 ( .B(A[934]), .A(S), .Z(O[934]) );
  ANDN U75 ( .B(A[933]), .A(S), .Z(O[933]) );
  ANDN U76 ( .B(A[932]), .A(S), .Z(O[932]) );
  ANDN U77 ( .B(A[931]), .A(S), .Z(O[931]) );
  ANDN U78 ( .B(A[930]), .A(S), .Z(O[930]) );
  ANDN U79 ( .B(A[92]), .A(S), .Z(O[92]) );
  ANDN U80 ( .B(A[929]), .A(S), .Z(O[929]) );
  ANDN U81 ( .B(A[928]), .A(S), .Z(O[928]) );
  ANDN U82 ( .B(A[927]), .A(S), .Z(O[927]) );
  ANDN U83 ( .B(A[926]), .A(S), .Z(O[926]) );
  ANDN U84 ( .B(A[925]), .A(S), .Z(O[925]) );
  ANDN U85 ( .B(A[924]), .A(S), .Z(O[924]) );
  ANDN U86 ( .B(A[923]), .A(S), .Z(O[923]) );
  ANDN U87 ( .B(A[922]), .A(S), .Z(O[922]) );
  ANDN U88 ( .B(A[921]), .A(S), .Z(O[921]) );
  ANDN U89 ( .B(A[920]), .A(S), .Z(O[920]) );
  ANDN U90 ( .B(A[91]), .A(S), .Z(O[91]) );
  ANDN U91 ( .B(A[919]), .A(S), .Z(O[919]) );
  ANDN U92 ( .B(A[918]), .A(S), .Z(O[918]) );
  ANDN U93 ( .B(A[917]), .A(S), .Z(O[917]) );
  ANDN U94 ( .B(A[916]), .A(S), .Z(O[916]) );
  ANDN U95 ( .B(A[915]), .A(S), .Z(O[915]) );
  ANDN U96 ( .B(A[914]), .A(S), .Z(O[914]) );
  ANDN U97 ( .B(A[913]), .A(S), .Z(O[913]) );
  ANDN U98 ( .B(A[912]), .A(S), .Z(O[912]) );
  ANDN U99 ( .B(A[911]), .A(S), .Z(O[911]) );
  ANDN U100 ( .B(A[910]), .A(S), .Z(O[910]) );
  ANDN U101 ( .B(A[90]), .A(S), .Z(O[90]) );
  ANDN U102 ( .B(A[909]), .A(S), .Z(O[909]) );
  ANDN U103 ( .B(A[908]), .A(S), .Z(O[908]) );
  ANDN U104 ( .B(A[907]), .A(S), .Z(O[907]) );
  ANDN U105 ( .B(A[906]), .A(S), .Z(O[906]) );
  ANDN U106 ( .B(A[905]), .A(S), .Z(O[905]) );
  ANDN U107 ( .B(A[904]), .A(S), .Z(O[904]) );
  ANDN U108 ( .B(A[903]), .A(S), .Z(O[903]) );
  ANDN U109 ( .B(A[902]), .A(S), .Z(O[902]) );
  ANDN U110 ( .B(A[901]), .A(S), .Z(O[901]) );
  ANDN U111 ( .B(A[900]), .A(S), .Z(O[900]) );
  ANDN U112 ( .B(A[8]), .A(S), .Z(O[8]) );
  ANDN U113 ( .B(A[89]), .A(S), .Z(O[89]) );
  ANDN U114 ( .B(A[899]), .A(S), .Z(O[899]) );
  ANDN U115 ( .B(A[898]), .A(S), .Z(O[898]) );
  ANDN U116 ( .B(A[897]), .A(S), .Z(O[897]) );
  ANDN U117 ( .B(A[896]), .A(S), .Z(O[896]) );
  ANDN U118 ( .B(A[895]), .A(S), .Z(O[895]) );
  ANDN U119 ( .B(A[894]), .A(S), .Z(O[894]) );
  ANDN U120 ( .B(A[893]), .A(S), .Z(O[893]) );
  ANDN U121 ( .B(A[892]), .A(S), .Z(O[892]) );
  ANDN U122 ( .B(A[891]), .A(S), .Z(O[891]) );
  ANDN U123 ( .B(A[890]), .A(S), .Z(O[890]) );
  ANDN U124 ( .B(A[88]), .A(S), .Z(O[88]) );
  ANDN U125 ( .B(A[889]), .A(S), .Z(O[889]) );
  ANDN U126 ( .B(A[888]), .A(S), .Z(O[888]) );
  ANDN U127 ( .B(A[887]), .A(S), .Z(O[887]) );
  ANDN U128 ( .B(A[886]), .A(S), .Z(O[886]) );
  ANDN U129 ( .B(A[885]), .A(S), .Z(O[885]) );
  ANDN U130 ( .B(A[884]), .A(S), .Z(O[884]) );
  ANDN U131 ( .B(A[883]), .A(S), .Z(O[883]) );
  ANDN U132 ( .B(A[882]), .A(S), .Z(O[882]) );
  ANDN U133 ( .B(A[881]), .A(S), .Z(O[881]) );
  ANDN U134 ( .B(A[880]), .A(S), .Z(O[880]) );
  ANDN U135 ( .B(A[87]), .A(S), .Z(O[87]) );
  ANDN U136 ( .B(A[879]), .A(S), .Z(O[879]) );
  ANDN U137 ( .B(A[878]), .A(S), .Z(O[878]) );
  ANDN U138 ( .B(A[877]), .A(S), .Z(O[877]) );
  ANDN U139 ( .B(A[876]), .A(S), .Z(O[876]) );
  ANDN U140 ( .B(A[875]), .A(S), .Z(O[875]) );
  ANDN U141 ( .B(A[874]), .A(S), .Z(O[874]) );
  ANDN U142 ( .B(A[873]), .A(S), .Z(O[873]) );
  ANDN U143 ( .B(A[872]), .A(S), .Z(O[872]) );
  ANDN U144 ( .B(A[871]), .A(S), .Z(O[871]) );
  ANDN U145 ( .B(A[870]), .A(S), .Z(O[870]) );
  ANDN U146 ( .B(A[86]), .A(S), .Z(O[86]) );
  ANDN U147 ( .B(A[869]), .A(S), .Z(O[869]) );
  ANDN U148 ( .B(A[868]), .A(S), .Z(O[868]) );
  ANDN U149 ( .B(A[867]), .A(S), .Z(O[867]) );
  ANDN U150 ( .B(A[866]), .A(S), .Z(O[866]) );
  ANDN U151 ( .B(A[865]), .A(S), .Z(O[865]) );
  ANDN U152 ( .B(A[864]), .A(S), .Z(O[864]) );
  ANDN U153 ( .B(A[863]), .A(S), .Z(O[863]) );
  ANDN U154 ( .B(A[862]), .A(S), .Z(O[862]) );
  ANDN U155 ( .B(A[861]), .A(S), .Z(O[861]) );
  ANDN U156 ( .B(A[860]), .A(S), .Z(O[860]) );
  ANDN U157 ( .B(A[85]), .A(S), .Z(O[85]) );
  ANDN U158 ( .B(A[859]), .A(S), .Z(O[859]) );
  ANDN U159 ( .B(A[858]), .A(S), .Z(O[858]) );
  ANDN U160 ( .B(A[857]), .A(S), .Z(O[857]) );
  ANDN U161 ( .B(A[856]), .A(S), .Z(O[856]) );
  ANDN U162 ( .B(A[855]), .A(S), .Z(O[855]) );
  ANDN U163 ( .B(A[854]), .A(S), .Z(O[854]) );
  ANDN U164 ( .B(A[853]), .A(S), .Z(O[853]) );
  ANDN U165 ( .B(A[852]), .A(S), .Z(O[852]) );
  ANDN U166 ( .B(A[851]), .A(S), .Z(O[851]) );
  ANDN U167 ( .B(A[850]), .A(S), .Z(O[850]) );
  ANDN U168 ( .B(A[84]), .A(S), .Z(O[84]) );
  ANDN U169 ( .B(A[849]), .A(S), .Z(O[849]) );
  ANDN U170 ( .B(A[848]), .A(S), .Z(O[848]) );
  ANDN U171 ( .B(A[847]), .A(S), .Z(O[847]) );
  ANDN U172 ( .B(A[846]), .A(S), .Z(O[846]) );
  ANDN U173 ( .B(A[845]), .A(S), .Z(O[845]) );
  ANDN U174 ( .B(A[844]), .A(S), .Z(O[844]) );
  ANDN U175 ( .B(A[843]), .A(S), .Z(O[843]) );
  ANDN U176 ( .B(A[842]), .A(S), .Z(O[842]) );
  ANDN U177 ( .B(A[841]), .A(S), .Z(O[841]) );
  ANDN U178 ( .B(A[840]), .A(S), .Z(O[840]) );
  ANDN U179 ( .B(A[83]), .A(S), .Z(O[83]) );
  ANDN U180 ( .B(A[839]), .A(S), .Z(O[839]) );
  ANDN U181 ( .B(A[838]), .A(S), .Z(O[838]) );
  ANDN U182 ( .B(A[837]), .A(S), .Z(O[837]) );
  ANDN U183 ( .B(A[836]), .A(S), .Z(O[836]) );
  ANDN U184 ( .B(A[835]), .A(S), .Z(O[835]) );
  ANDN U185 ( .B(A[834]), .A(S), .Z(O[834]) );
  ANDN U186 ( .B(A[833]), .A(S), .Z(O[833]) );
  ANDN U187 ( .B(A[832]), .A(S), .Z(O[832]) );
  ANDN U188 ( .B(A[831]), .A(S), .Z(O[831]) );
  ANDN U189 ( .B(A[830]), .A(S), .Z(O[830]) );
  ANDN U190 ( .B(A[82]), .A(S), .Z(O[82]) );
  ANDN U191 ( .B(A[829]), .A(S), .Z(O[829]) );
  ANDN U192 ( .B(A[828]), .A(S), .Z(O[828]) );
  ANDN U193 ( .B(A[827]), .A(S), .Z(O[827]) );
  ANDN U194 ( .B(A[826]), .A(S), .Z(O[826]) );
  ANDN U195 ( .B(A[825]), .A(S), .Z(O[825]) );
  ANDN U196 ( .B(A[824]), .A(S), .Z(O[824]) );
  ANDN U197 ( .B(A[823]), .A(S), .Z(O[823]) );
  ANDN U198 ( .B(A[822]), .A(S), .Z(O[822]) );
  ANDN U199 ( .B(A[821]), .A(S), .Z(O[821]) );
  ANDN U200 ( .B(A[820]), .A(S), .Z(O[820]) );
  ANDN U201 ( .B(A[81]), .A(S), .Z(O[81]) );
  ANDN U202 ( .B(A[819]), .A(S), .Z(O[819]) );
  ANDN U203 ( .B(A[818]), .A(S), .Z(O[818]) );
  ANDN U204 ( .B(A[817]), .A(S), .Z(O[817]) );
  ANDN U205 ( .B(A[816]), .A(S), .Z(O[816]) );
  ANDN U206 ( .B(A[815]), .A(S), .Z(O[815]) );
  ANDN U207 ( .B(A[814]), .A(S), .Z(O[814]) );
  ANDN U208 ( .B(A[813]), .A(S), .Z(O[813]) );
  ANDN U209 ( .B(A[812]), .A(S), .Z(O[812]) );
  ANDN U210 ( .B(A[811]), .A(S), .Z(O[811]) );
  ANDN U211 ( .B(A[810]), .A(S), .Z(O[810]) );
  ANDN U212 ( .B(A[80]), .A(S), .Z(O[80]) );
  ANDN U213 ( .B(A[809]), .A(S), .Z(O[809]) );
  ANDN U214 ( .B(A[808]), .A(S), .Z(O[808]) );
  ANDN U215 ( .B(A[807]), .A(S), .Z(O[807]) );
  ANDN U216 ( .B(A[806]), .A(S), .Z(O[806]) );
  ANDN U217 ( .B(A[805]), .A(S), .Z(O[805]) );
  ANDN U218 ( .B(A[804]), .A(S), .Z(O[804]) );
  ANDN U219 ( .B(A[803]), .A(S), .Z(O[803]) );
  ANDN U220 ( .B(A[802]), .A(S), .Z(O[802]) );
  ANDN U221 ( .B(A[801]), .A(S), .Z(O[801]) );
  ANDN U222 ( .B(A[800]), .A(S), .Z(O[800]) );
  ANDN U223 ( .B(A[7]), .A(S), .Z(O[7]) );
  ANDN U224 ( .B(A[79]), .A(S), .Z(O[79]) );
  ANDN U225 ( .B(A[799]), .A(S), .Z(O[799]) );
  ANDN U226 ( .B(A[798]), .A(S), .Z(O[798]) );
  ANDN U227 ( .B(A[797]), .A(S), .Z(O[797]) );
  ANDN U228 ( .B(A[796]), .A(S), .Z(O[796]) );
  ANDN U229 ( .B(A[795]), .A(S), .Z(O[795]) );
  ANDN U230 ( .B(A[794]), .A(S), .Z(O[794]) );
  ANDN U231 ( .B(A[793]), .A(S), .Z(O[793]) );
  ANDN U232 ( .B(A[792]), .A(S), .Z(O[792]) );
  ANDN U233 ( .B(A[791]), .A(S), .Z(O[791]) );
  ANDN U234 ( .B(A[790]), .A(S), .Z(O[790]) );
  ANDN U235 ( .B(A[78]), .A(S), .Z(O[78]) );
  ANDN U236 ( .B(A[789]), .A(S), .Z(O[789]) );
  ANDN U237 ( .B(A[788]), .A(S), .Z(O[788]) );
  ANDN U238 ( .B(A[787]), .A(S), .Z(O[787]) );
  ANDN U239 ( .B(A[786]), .A(S), .Z(O[786]) );
  ANDN U240 ( .B(A[785]), .A(S), .Z(O[785]) );
  ANDN U241 ( .B(A[784]), .A(S), .Z(O[784]) );
  ANDN U242 ( .B(A[783]), .A(S), .Z(O[783]) );
  ANDN U243 ( .B(A[782]), .A(S), .Z(O[782]) );
  ANDN U244 ( .B(A[781]), .A(S), .Z(O[781]) );
  ANDN U245 ( .B(A[780]), .A(S), .Z(O[780]) );
  ANDN U246 ( .B(A[77]), .A(S), .Z(O[77]) );
  ANDN U247 ( .B(A[779]), .A(S), .Z(O[779]) );
  ANDN U248 ( .B(A[778]), .A(S), .Z(O[778]) );
  ANDN U249 ( .B(A[777]), .A(S), .Z(O[777]) );
  ANDN U250 ( .B(A[776]), .A(S), .Z(O[776]) );
  ANDN U251 ( .B(A[775]), .A(S), .Z(O[775]) );
  ANDN U252 ( .B(A[774]), .A(S), .Z(O[774]) );
  ANDN U253 ( .B(A[773]), .A(S), .Z(O[773]) );
  ANDN U254 ( .B(A[772]), .A(S), .Z(O[772]) );
  ANDN U255 ( .B(A[771]), .A(S), .Z(O[771]) );
  ANDN U256 ( .B(A[770]), .A(S), .Z(O[770]) );
  ANDN U257 ( .B(A[76]), .A(S), .Z(O[76]) );
  ANDN U258 ( .B(A[769]), .A(S), .Z(O[769]) );
  ANDN U259 ( .B(A[768]), .A(S), .Z(O[768]) );
  ANDN U260 ( .B(A[767]), .A(S), .Z(O[767]) );
  ANDN U261 ( .B(A[766]), .A(S), .Z(O[766]) );
  ANDN U262 ( .B(A[765]), .A(S), .Z(O[765]) );
  ANDN U263 ( .B(A[764]), .A(S), .Z(O[764]) );
  ANDN U264 ( .B(A[763]), .A(S), .Z(O[763]) );
  ANDN U265 ( .B(A[762]), .A(S), .Z(O[762]) );
  ANDN U266 ( .B(A[761]), .A(S), .Z(O[761]) );
  ANDN U267 ( .B(A[760]), .A(S), .Z(O[760]) );
  ANDN U268 ( .B(A[75]), .A(S), .Z(O[75]) );
  ANDN U269 ( .B(A[759]), .A(S), .Z(O[759]) );
  ANDN U270 ( .B(A[758]), .A(S), .Z(O[758]) );
  ANDN U271 ( .B(A[757]), .A(S), .Z(O[757]) );
  ANDN U272 ( .B(A[756]), .A(S), .Z(O[756]) );
  ANDN U273 ( .B(A[755]), .A(S), .Z(O[755]) );
  ANDN U274 ( .B(A[754]), .A(S), .Z(O[754]) );
  ANDN U275 ( .B(A[753]), .A(S), .Z(O[753]) );
  ANDN U276 ( .B(A[752]), .A(S), .Z(O[752]) );
  ANDN U277 ( .B(A[751]), .A(S), .Z(O[751]) );
  ANDN U278 ( .B(A[750]), .A(S), .Z(O[750]) );
  ANDN U279 ( .B(A[74]), .A(S), .Z(O[74]) );
  ANDN U280 ( .B(A[749]), .A(S), .Z(O[749]) );
  ANDN U281 ( .B(A[748]), .A(S), .Z(O[748]) );
  ANDN U282 ( .B(A[747]), .A(S), .Z(O[747]) );
  ANDN U283 ( .B(A[746]), .A(S), .Z(O[746]) );
  ANDN U284 ( .B(A[745]), .A(S), .Z(O[745]) );
  ANDN U285 ( .B(A[744]), .A(S), .Z(O[744]) );
  ANDN U286 ( .B(A[743]), .A(S), .Z(O[743]) );
  ANDN U287 ( .B(A[742]), .A(S), .Z(O[742]) );
  ANDN U288 ( .B(A[741]), .A(S), .Z(O[741]) );
  ANDN U289 ( .B(A[740]), .A(S), .Z(O[740]) );
  ANDN U290 ( .B(A[73]), .A(S), .Z(O[73]) );
  ANDN U291 ( .B(A[739]), .A(S), .Z(O[739]) );
  ANDN U292 ( .B(A[738]), .A(S), .Z(O[738]) );
  ANDN U293 ( .B(A[737]), .A(S), .Z(O[737]) );
  ANDN U294 ( .B(A[736]), .A(S), .Z(O[736]) );
  ANDN U295 ( .B(A[735]), .A(S), .Z(O[735]) );
  ANDN U296 ( .B(A[734]), .A(S), .Z(O[734]) );
  ANDN U297 ( .B(A[733]), .A(S), .Z(O[733]) );
  ANDN U298 ( .B(A[732]), .A(S), .Z(O[732]) );
  ANDN U299 ( .B(A[731]), .A(S), .Z(O[731]) );
  ANDN U300 ( .B(A[730]), .A(S), .Z(O[730]) );
  ANDN U301 ( .B(A[72]), .A(S), .Z(O[72]) );
  ANDN U302 ( .B(A[729]), .A(S), .Z(O[729]) );
  ANDN U303 ( .B(A[728]), .A(S), .Z(O[728]) );
  ANDN U304 ( .B(A[727]), .A(S), .Z(O[727]) );
  ANDN U305 ( .B(A[726]), .A(S), .Z(O[726]) );
  ANDN U306 ( .B(A[725]), .A(S), .Z(O[725]) );
  ANDN U307 ( .B(A[724]), .A(S), .Z(O[724]) );
  ANDN U308 ( .B(A[723]), .A(S), .Z(O[723]) );
  ANDN U309 ( .B(A[722]), .A(S), .Z(O[722]) );
  ANDN U310 ( .B(A[721]), .A(S), .Z(O[721]) );
  ANDN U311 ( .B(A[720]), .A(S), .Z(O[720]) );
  ANDN U312 ( .B(A[71]), .A(S), .Z(O[71]) );
  ANDN U313 ( .B(A[719]), .A(S), .Z(O[719]) );
  ANDN U314 ( .B(A[718]), .A(S), .Z(O[718]) );
  ANDN U315 ( .B(A[717]), .A(S), .Z(O[717]) );
  ANDN U316 ( .B(A[716]), .A(S), .Z(O[716]) );
  ANDN U317 ( .B(A[715]), .A(S), .Z(O[715]) );
  ANDN U318 ( .B(A[714]), .A(S), .Z(O[714]) );
  ANDN U319 ( .B(A[713]), .A(S), .Z(O[713]) );
  ANDN U320 ( .B(A[712]), .A(S), .Z(O[712]) );
  ANDN U321 ( .B(A[711]), .A(S), .Z(O[711]) );
  ANDN U322 ( .B(A[710]), .A(S), .Z(O[710]) );
  ANDN U323 ( .B(A[70]), .A(S), .Z(O[70]) );
  ANDN U324 ( .B(A[709]), .A(S), .Z(O[709]) );
  ANDN U325 ( .B(A[708]), .A(S), .Z(O[708]) );
  ANDN U326 ( .B(A[707]), .A(S), .Z(O[707]) );
  ANDN U327 ( .B(A[706]), .A(S), .Z(O[706]) );
  ANDN U328 ( .B(A[705]), .A(S), .Z(O[705]) );
  ANDN U329 ( .B(A[704]), .A(S), .Z(O[704]) );
  ANDN U330 ( .B(A[703]), .A(S), .Z(O[703]) );
  ANDN U331 ( .B(A[702]), .A(S), .Z(O[702]) );
  ANDN U332 ( .B(A[701]), .A(S), .Z(O[701]) );
  ANDN U333 ( .B(A[700]), .A(S), .Z(O[700]) );
  ANDN U334 ( .B(A[6]), .A(S), .Z(O[6]) );
  ANDN U335 ( .B(A[69]), .A(S), .Z(O[69]) );
  ANDN U336 ( .B(A[699]), .A(S), .Z(O[699]) );
  ANDN U337 ( .B(A[698]), .A(S), .Z(O[698]) );
  ANDN U338 ( .B(A[697]), .A(S), .Z(O[697]) );
  ANDN U339 ( .B(A[696]), .A(S), .Z(O[696]) );
  ANDN U340 ( .B(A[695]), .A(S), .Z(O[695]) );
  ANDN U341 ( .B(A[694]), .A(S), .Z(O[694]) );
  ANDN U342 ( .B(A[693]), .A(S), .Z(O[693]) );
  ANDN U343 ( .B(A[692]), .A(S), .Z(O[692]) );
  ANDN U344 ( .B(A[691]), .A(S), .Z(O[691]) );
  ANDN U345 ( .B(A[690]), .A(S), .Z(O[690]) );
  ANDN U346 ( .B(A[68]), .A(S), .Z(O[68]) );
  ANDN U347 ( .B(A[689]), .A(S), .Z(O[689]) );
  ANDN U348 ( .B(A[688]), .A(S), .Z(O[688]) );
  ANDN U349 ( .B(A[687]), .A(S), .Z(O[687]) );
  ANDN U350 ( .B(A[686]), .A(S), .Z(O[686]) );
  ANDN U351 ( .B(A[685]), .A(S), .Z(O[685]) );
  ANDN U352 ( .B(A[684]), .A(S), .Z(O[684]) );
  ANDN U353 ( .B(A[683]), .A(S), .Z(O[683]) );
  ANDN U354 ( .B(A[682]), .A(S), .Z(O[682]) );
  ANDN U355 ( .B(A[681]), .A(S), .Z(O[681]) );
  ANDN U356 ( .B(A[680]), .A(S), .Z(O[680]) );
  ANDN U357 ( .B(A[67]), .A(S), .Z(O[67]) );
  ANDN U358 ( .B(A[679]), .A(S), .Z(O[679]) );
  ANDN U359 ( .B(A[678]), .A(S), .Z(O[678]) );
  ANDN U360 ( .B(A[677]), .A(S), .Z(O[677]) );
  ANDN U361 ( .B(A[676]), .A(S), .Z(O[676]) );
  ANDN U362 ( .B(A[675]), .A(S), .Z(O[675]) );
  ANDN U363 ( .B(A[674]), .A(S), .Z(O[674]) );
  ANDN U364 ( .B(A[673]), .A(S), .Z(O[673]) );
  ANDN U365 ( .B(A[672]), .A(S), .Z(O[672]) );
  ANDN U366 ( .B(A[671]), .A(S), .Z(O[671]) );
  ANDN U367 ( .B(A[670]), .A(S), .Z(O[670]) );
  ANDN U368 ( .B(A[66]), .A(S), .Z(O[66]) );
  ANDN U369 ( .B(A[669]), .A(S), .Z(O[669]) );
  ANDN U370 ( .B(A[668]), .A(S), .Z(O[668]) );
  ANDN U371 ( .B(A[667]), .A(S), .Z(O[667]) );
  ANDN U372 ( .B(A[666]), .A(S), .Z(O[666]) );
  ANDN U373 ( .B(A[665]), .A(S), .Z(O[665]) );
  ANDN U374 ( .B(A[664]), .A(S), .Z(O[664]) );
  ANDN U375 ( .B(A[663]), .A(S), .Z(O[663]) );
  ANDN U376 ( .B(A[662]), .A(S), .Z(O[662]) );
  ANDN U377 ( .B(A[661]), .A(S), .Z(O[661]) );
  ANDN U378 ( .B(A[660]), .A(S), .Z(O[660]) );
  ANDN U379 ( .B(A[65]), .A(S), .Z(O[65]) );
  ANDN U380 ( .B(A[659]), .A(S), .Z(O[659]) );
  ANDN U381 ( .B(A[658]), .A(S), .Z(O[658]) );
  ANDN U382 ( .B(A[657]), .A(S), .Z(O[657]) );
  ANDN U383 ( .B(A[656]), .A(S), .Z(O[656]) );
  ANDN U384 ( .B(A[655]), .A(S), .Z(O[655]) );
  ANDN U385 ( .B(A[654]), .A(S), .Z(O[654]) );
  ANDN U386 ( .B(A[653]), .A(S), .Z(O[653]) );
  ANDN U387 ( .B(A[652]), .A(S), .Z(O[652]) );
  ANDN U388 ( .B(A[651]), .A(S), .Z(O[651]) );
  ANDN U389 ( .B(A[650]), .A(S), .Z(O[650]) );
  ANDN U390 ( .B(A[64]), .A(S), .Z(O[64]) );
  ANDN U391 ( .B(A[649]), .A(S), .Z(O[649]) );
  ANDN U392 ( .B(A[648]), .A(S), .Z(O[648]) );
  ANDN U393 ( .B(A[647]), .A(S), .Z(O[647]) );
  ANDN U394 ( .B(A[646]), .A(S), .Z(O[646]) );
  ANDN U395 ( .B(A[645]), .A(S), .Z(O[645]) );
  ANDN U396 ( .B(A[644]), .A(S), .Z(O[644]) );
  ANDN U397 ( .B(A[643]), .A(S), .Z(O[643]) );
  ANDN U398 ( .B(A[642]), .A(S), .Z(O[642]) );
  ANDN U399 ( .B(A[641]), .A(S), .Z(O[641]) );
  ANDN U400 ( .B(A[640]), .A(S), .Z(O[640]) );
  ANDN U401 ( .B(A[63]), .A(S), .Z(O[63]) );
  ANDN U402 ( .B(A[639]), .A(S), .Z(O[639]) );
  ANDN U403 ( .B(A[638]), .A(S), .Z(O[638]) );
  ANDN U404 ( .B(A[637]), .A(S), .Z(O[637]) );
  ANDN U405 ( .B(A[636]), .A(S), .Z(O[636]) );
  ANDN U406 ( .B(A[635]), .A(S), .Z(O[635]) );
  ANDN U407 ( .B(A[634]), .A(S), .Z(O[634]) );
  ANDN U408 ( .B(A[633]), .A(S), .Z(O[633]) );
  ANDN U409 ( .B(A[632]), .A(S), .Z(O[632]) );
  ANDN U410 ( .B(A[631]), .A(S), .Z(O[631]) );
  ANDN U411 ( .B(A[630]), .A(S), .Z(O[630]) );
  ANDN U412 ( .B(A[62]), .A(S), .Z(O[62]) );
  ANDN U413 ( .B(A[629]), .A(S), .Z(O[629]) );
  ANDN U414 ( .B(A[628]), .A(S), .Z(O[628]) );
  ANDN U415 ( .B(A[627]), .A(S), .Z(O[627]) );
  ANDN U416 ( .B(A[626]), .A(S), .Z(O[626]) );
  ANDN U417 ( .B(A[625]), .A(S), .Z(O[625]) );
  ANDN U418 ( .B(A[624]), .A(S), .Z(O[624]) );
  ANDN U419 ( .B(A[623]), .A(S), .Z(O[623]) );
  ANDN U420 ( .B(A[622]), .A(S), .Z(O[622]) );
  ANDN U421 ( .B(A[621]), .A(S), .Z(O[621]) );
  ANDN U422 ( .B(A[620]), .A(S), .Z(O[620]) );
  ANDN U423 ( .B(A[61]), .A(S), .Z(O[61]) );
  ANDN U424 ( .B(A[619]), .A(S), .Z(O[619]) );
  ANDN U425 ( .B(A[618]), .A(S), .Z(O[618]) );
  ANDN U426 ( .B(A[617]), .A(S), .Z(O[617]) );
  ANDN U427 ( .B(A[616]), .A(S), .Z(O[616]) );
  ANDN U428 ( .B(A[615]), .A(S), .Z(O[615]) );
  ANDN U429 ( .B(A[614]), .A(S), .Z(O[614]) );
  ANDN U430 ( .B(A[613]), .A(S), .Z(O[613]) );
  ANDN U431 ( .B(A[612]), .A(S), .Z(O[612]) );
  ANDN U432 ( .B(A[611]), .A(S), .Z(O[611]) );
  ANDN U433 ( .B(A[610]), .A(S), .Z(O[610]) );
  ANDN U434 ( .B(A[60]), .A(S), .Z(O[60]) );
  ANDN U435 ( .B(A[609]), .A(S), .Z(O[609]) );
  ANDN U436 ( .B(A[608]), .A(S), .Z(O[608]) );
  ANDN U437 ( .B(A[607]), .A(S), .Z(O[607]) );
  ANDN U438 ( .B(A[606]), .A(S), .Z(O[606]) );
  ANDN U439 ( .B(A[605]), .A(S), .Z(O[605]) );
  ANDN U440 ( .B(A[604]), .A(S), .Z(O[604]) );
  ANDN U441 ( .B(A[603]), .A(S), .Z(O[603]) );
  ANDN U442 ( .B(A[602]), .A(S), .Z(O[602]) );
  ANDN U443 ( .B(A[601]), .A(S), .Z(O[601]) );
  ANDN U444 ( .B(A[600]), .A(S), .Z(O[600]) );
  ANDN U445 ( .B(A[5]), .A(S), .Z(O[5]) );
  ANDN U446 ( .B(A[59]), .A(S), .Z(O[59]) );
  ANDN U447 ( .B(A[599]), .A(S), .Z(O[599]) );
  ANDN U448 ( .B(A[598]), .A(S), .Z(O[598]) );
  ANDN U449 ( .B(A[597]), .A(S), .Z(O[597]) );
  ANDN U450 ( .B(A[596]), .A(S), .Z(O[596]) );
  ANDN U451 ( .B(A[595]), .A(S), .Z(O[595]) );
  ANDN U452 ( .B(A[594]), .A(S), .Z(O[594]) );
  ANDN U453 ( .B(A[593]), .A(S), .Z(O[593]) );
  ANDN U454 ( .B(A[592]), .A(S), .Z(O[592]) );
  ANDN U455 ( .B(A[591]), .A(S), .Z(O[591]) );
  ANDN U456 ( .B(A[590]), .A(S), .Z(O[590]) );
  ANDN U457 ( .B(A[58]), .A(S), .Z(O[58]) );
  ANDN U458 ( .B(A[589]), .A(S), .Z(O[589]) );
  ANDN U459 ( .B(A[588]), .A(S), .Z(O[588]) );
  ANDN U460 ( .B(A[587]), .A(S), .Z(O[587]) );
  ANDN U461 ( .B(A[586]), .A(S), .Z(O[586]) );
  ANDN U462 ( .B(A[585]), .A(S), .Z(O[585]) );
  ANDN U463 ( .B(A[584]), .A(S), .Z(O[584]) );
  ANDN U464 ( .B(A[583]), .A(S), .Z(O[583]) );
  ANDN U465 ( .B(A[582]), .A(S), .Z(O[582]) );
  ANDN U466 ( .B(A[581]), .A(S), .Z(O[581]) );
  ANDN U467 ( .B(A[580]), .A(S), .Z(O[580]) );
  ANDN U468 ( .B(A[57]), .A(S), .Z(O[57]) );
  ANDN U469 ( .B(A[579]), .A(S), .Z(O[579]) );
  ANDN U470 ( .B(A[578]), .A(S), .Z(O[578]) );
  ANDN U471 ( .B(A[577]), .A(S), .Z(O[577]) );
  ANDN U472 ( .B(A[576]), .A(S), .Z(O[576]) );
  ANDN U473 ( .B(A[575]), .A(S), .Z(O[575]) );
  ANDN U474 ( .B(A[574]), .A(S), .Z(O[574]) );
  ANDN U475 ( .B(A[573]), .A(S), .Z(O[573]) );
  ANDN U476 ( .B(A[572]), .A(S), .Z(O[572]) );
  ANDN U477 ( .B(A[571]), .A(S), .Z(O[571]) );
  ANDN U478 ( .B(A[570]), .A(S), .Z(O[570]) );
  ANDN U479 ( .B(A[56]), .A(S), .Z(O[56]) );
  ANDN U480 ( .B(A[569]), .A(S), .Z(O[569]) );
  ANDN U481 ( .B(A[568]), .A(S), .Z(O[568]) );
  ANDN U482 ( .B(A[567]), .A(S), .Z(O[567]) );
  ANDN U483 ( .B(A[566]), .A(S), .Z(O[566]) );
  ANDN U484 ( .B(A[565]), .A(S), .Z(O[565]) );
  ANDN U485 ( .B(A[564]), .A(S), .Z(O[564]) );
  ANDN U486 ( .B(A[563]), .A(S), .Z(O[563]) );
  ANDN U487 ( .B(A[562]), .A(S), .Z(O[562]) );
  ANDN U488 ( .B(A[561]), .A(S), .Z(O[561]) );
  ANDN U489 ( .B(A[560]), .A(S), .Z(O[560]) );
  ANDN U490 ( .B(A[55]), .A(S), .Z(O[55]) );
  ANDN U491 ( .B(A[559]), .A(S), .Z(O[559]) );
  ANDN U492 ( .B(A[558]), .A(S), .Z(O[558]) );
  ANDN U493 ( .B(A[557]), .A(S), .Z(O[557]) );
  ANDN U494 ( .B(A[556]), .A(S), .Z(O[556]) );
  ANDN U495 ( .B(A[555]), .A(S), .Z(O[555]) );
  ANDN U496 ( .B(A[554]), .A(S), .Z(O[554]) );
  ANDN U497 ( .B(A[553]), .A(S), .Z(O[553]) );
  ANDN U498 ( .B(A[552]), .A(S), .Z(O[552]) );
  ANDN U499 ( .B(A[551]), .A(S), .Z(O[551]) );
  ANDN U500 ( .B(A[550]), .A(S), .Z(O[550]) );
  ANDN U501 ( .B(A[54]), .A(S), .Z(O[54]) );
  ANDN U502 ( .B(A[549]), .A(S), .Z(O[549]) );
  ANDN U503 ( .B(A[548]), .A(S), .Z(O[548]) );
  ANDN U504 ( .B(A[547]), .A(S), .Z(O[547]) );
  ANDN U505 ( .B(A[546]), .A(S), .Z(O[546]) );
  ANDN U506 ( .B(A[545]), .A(S), .Z(O[545]) );
  ANDN U507 ( .B(A[544]), .A(S), .Z(O[544]) );
  ANDN U508 ( .B(A[543]), .A(S), .Z(O[543]) );
  ANDN U509 ( .B(A[542]), .A(S), .Z(O[542]) );
  ANDN U510 ( .B(A[541]), .A(S), .Z(O[541]) );
  ANDN U511 ( .B(A[540]), .A(S), .Z(O[540]) );
  ANDN U512 ( .B(A[53]), .A(S), .Z(O[53]) );
  ANDN U513 ( .B(A[539]), .A(S), .Z(O[539]) );
  ANDN U514 ( .B(A[538]), .A(S), .Z(O[538]) );
  ANDN U515 ( .B(A[537]), .A(S), .Z(O[537]) );
  ANDN U516 ( .B(A[536]), .A(S), .Z(O[536]) );
  ANDN U517 ( .B(A[535]), .A(S), .Z(O[535]) );
  ANDN U518 ( .B(A[534]), .A(S), .Z(O[534]) );
  ANDN U519 ( .B(A[533]), .A(S), .Z(O[533]) );
  ANDN U520 ( .B(A[532]), .A(S), .Z(O[532]) );
  ANDN U521 ( .B(A[531]), .A(S), .Z(O[531]) );
  ANDN U522 ( .B(A[530]), .A(S), .Z(O[530]) );
  ANDN U523 ( .B(A[52]), .A(S), .Z(O[52]) );
  ANDN U524 ( .B(A[529]), .A(S), .Z(O[529]) );
  ANDN U525 ( .B(A[528]), .A(S), .Z(O[528]) );
  ANDN U526 ( .B(A[527]), .A(S), .Z(O[527]) );
  ANDN U527 ( .B(A[526]), .A(S), .Z(O[526]) );
  ANDN U528 ( .B(A[525]), .A(S), .Z(O[525]) );
  ANDN U529 ( .B(A[524]), .A(S), .Z(O[524]) );
  ANDN U530 ( .B(A[523]), .A(S), .Z(O[523]) );
  ANDN U531 ( .B(A[522]), .A(S), .Z(O[522]) );
  ANDN U532 ( .B(A[521]), .A(S), .Z(O[521]) );
  ANDN U533 ( .B(A[520]), .A(S), .Z(O[520]) );
  ANDN U534 ( .B(A[51]), .A(S), .Z(O[51]) );
  ANDN U535 ( .B(A[519]), .A(S), .Z(O[519]) );
  ANDN U536 ( .B(A[518]), .A(S), .Z(O[518]) );
  ANDN U537 ( .B(A[517]), .A(S), .Z(O[517]) );
  ANDN U538 ( .B(A[516]), .A(S), .Z(O[516]) );
  ANDN U539 ( .B(A[515]), .A(S), .Z(O[515]) );
  ANDN U540 ( .B(A[514]), .A(S), .Z(O[514]) );
  ANDN U541 ( .B(A[513]), .A(S), .Z(O[513]) );
  ANDN U542 ( .B(A[512]), .A(S), .Z(O[512]) );
  ANDN U543 ( .B(A[511]), .A(S), .Z(O[511]) );
  ANDN U544 ( .B(A[510]), .A(S), .Z(O[510]) );
  ANDN U545 ( .B(A[50]), .A(S), .Z(O[50]) );
  ANDN U546 ( .B(A[509]), .A(S), .Z(O[509]) );
  ANDN U547 ( .B(A[508]), .A(S), .Z(O[508]) );
  ANDN U548 ( .B(A[507]), .A(S), .Z(O[507]) );
  ANDN U549 ( .B(A[506]), .A(S), .Z(O[506]) );
  ANDN U550 ( .B(A[505]), .A(S), .Z(O[505]) );
  ANDN U551 ( .B(A[504]), .A(S), .Z(O[504]) );
  ANDN U552 ( .B(A[503]), .A(S), .Z(O[503]) );
  ANDN U553 ( .B(A[502]), .A(S), .Z(O[502]) );
  ANDN U554 ( .B(A[501]), .A(S), .Z(O[501]) );
  ANDN U555 ( .B(A[500]), .A(S), .Z(O[500]) );
  ANDN U556 ( .B(A[4]), .A(S), .Z(O[4]) );
  ANDN U557 ( .B(A[49]), .A(S), .Z(O[49]) );
  ANDN U558 ( .B(A[499]), .A(S), .Z(O[499]) );
  ANDN U559 ( .B(A[498]), .A(S), .Z(O[498]) );
  ANDN U560 ( .B(A[497]), .A(S), .Z(O[497]) );
  ANDN U561 ( .B(A[496]), .A(S), .Z(O[496]) );
  ANDN U562 ( .B(A[495]), .A(S), .Z(O[495]) );
  ANDN U563 ( .B(A[494]), .A(S), .Z(O[494]) );
  ANDN U564 ( .B(A[493]), .A(S), .Z(O[493]) );
  ANDN U565 ( .B(A[492]), .A(S), .Z(O[492]) );
  ANDN U566 ( .B(A[491]), .A(S), .Z(O[491]) );
  ANDN U567 ( .B(A[490]), .A(S), .Z(O[490]) );
  ANDN U568 ( .B(A[48]), .A(S), .Z(O[48]) );
  ANDN U569 ( .B(A[489]), .A(S), .Z(O[489]) );
  ANDN U570 ( .B(A[488]), .A(S), .Z(O[488]) );
  ANDN U571 ( .B(A[487]), .A(S), .Z(O[487]) );
  ANDN U572 ( .B(A[486]), .A(S), .Z(O[486]) );
  ANDN U573 ( .B(A[485]), .A(S), .Z(O[485]) );
  ANDN U574 ( .B(A[484]), .A(S), .Z(O[484]) );
  ANDN U575 ( .B(A[483]), .A(S), .Z(O[483]) );
  ANDN U576 ( .B(A[482]), .A(S), .Z(O[482]) );
  ANDN U577 ( .B(A[481]), .A(S), .Z(O[481]) );
  ANDN U578 ( .B(A[480]), .A(S), .Z(O[480]) );
  ANDN U579 ( .B(A[47]), .A(S), .Z(O[47]) );
  ANDN U580 ( .B(A[479]), .A(S), .Z(O[479]) );
  ANDN U581 ( .B(A[478]), .A(S), .Z(O[478]) );
  ANDN U582 ( .B(A[477]), .A(S), .Z(O[477]) );
  ANDN U583 ( .B(A[476]), .A(S), .Z(O[476]) );
  ANDN U584 ( .B(A[475]), .A(S), .Z(O[475]) );
  ANDN U585 ( .B(A[474]), .A(S), .Z(O[474]) );
  ANDN U586 ( .B(A[473]), .A(S), .Z(O[473]) );
  ANDN U587 ( .B(A[472]), .A(S), .Z(O[472]) );
  ANDN U588 ( .B(A[471]), .A(S), .Z(O[471]) );
  ANDN U589 ( .B(A[470]), .A(S), .Z(O[470]) );
  ANDN U590 ( .B(A[46]), .A(S), .Z(O[46]) );
  ANDN U591 ( .B(A[469]), .A(S), .Z(O[469]) );
  ANDN U592 ( .B(A[468]), .A(S), .Z(O[468]) );
  ANDN U593 ( .B(A[467]), .A(S), .Z(O[467]) );
  ANDN U594 ( .B(A[466]), .A(S), .Z(O[466]) );
  ANDN U595 ( .B(A[465]), .A(S), .Z(O[465]) );
  ANDN U596 ( .B(A[464]), .A(S), .Z(O[464]) );
  ANDN U597 ( .B(A[463]), .A(S), .Z(O[463]) );
  ANDN U598 ( .B(A[462]), .A(S), .Z(O[462]) );
  ANDN U599 ( .B(A[461]), .A(S), .Z(O[461]) );
  ANDN U600 ( .B(A[460]), .A(S), .Z(O[460]) );
  ANDN U601 ( .B(A[45]), .A(S), .Z(O[45]) );
  ANDN U602 ( .B(A[459]), .A(S), .Z(O[459]) );
  ANDN U603 ( .B(A[458]), .A(S), .Z(O[458]) );
  ANDN U604 ( .B(A[457]), .A(S), .Z(O[457]) );
  ANDN U605 ( .B(A[456]), .A(S), .Z(O[456]) );
  ANDN U606 ( .B(A[455]), .A(S), .Z(O[455]) );
  ANDN U607 ( .B(A[454]), .A(S), .Z(O[454]) );
  ANDN U608 ( .B(A[453]), .A(S), .Z(O[453]) );
  ANDN U609 ( .B(A[452]), .A(S), .Z(O[452]) );
  ANDN U610 ( .B(A[451]), .A(S), .Z(O[451]) );
  ANDN U611 ( .B(A[450]), .A(S), .Z(O[450]) );
  ANDN U612 ( .B(A[44]), .A(S), .Z(O[44]) );
  ANDN U613 ( .B(A[449]), .A(S), .Z(O[449]) );
  ANDN U614 ( .B(A[448]), .A(S), .Z(O[448]) );
  ANDN U615 ( .B(A[447]), .A(S), .Z(O[447]) );
  ANDN U616 ( .B(A[446]), .A(S), .Z(O[446]) );
  ANDN U617 ( .B(A[445]), .A(S), .Z(O[445]) );
  ANDN U618 ( .B(A[444]), .A(S), .Z(O[444]) );
  ANDN U619 ( .B(A[443]), .A(S), .Z(O[443]) );
  ANDN U620 ( .B(A[442]), .A(S), .Z(O[442]) );
  ANDN U621 ( .B(A[441]), .A(S), .Z(O[441]) );
  ANDN U622 ( .B(A[440]), .A(S), .Z(O[440]) );
  ANDN U623 ( .B(A[43]), .A(S), .Z(O[43]) );
  ANDN U624 ( .B(A[439]), .A(S), .Z(O[439]) );
  ANDN U625 ( .B(A[438]), .A(S), .Z(O[438]) );
  ANDN U626 ( .B(A[437]), .A(S), .Z(O[437]) );
  ANDN U627 ( .B(A[436]), .A(S), .Z(O[436]) );
  ANDN U628 ( .B(A[435]), .A(S), .Z(O[435]) );
  ANDN U629 ( .B(A[434]), .A(S), .Z(O[434]) );
  ANDN U630 ( .B(A[433]), .A(S), .Z(O[433]) );
  ANDN U631 ( .B(A[432]), .A(S), .Z(O[432]) );
  ANDN U632 ( .B(A[431]), .A(S), .Z(O[431]) );
  ANDN U633 ( .B(A[430]), .A(S), .Z(O[430]) );
  ANDN U634 ( .B(A[42]), .A(S), .Z(O[42]) );
  ANDN U635 ( .B(A[429]), .A(S), .Z(O[429]) );
  ANDN U636 ( .B(A[428]), .A(S), .Z(O[428]) );
  ANDN U637 ( .B(A[427]), .A(S), .Z(O[427]) );
  ANDN U638 ( .B(A[426]), .A(S), .Z(O[426]) );
  ANDN U639 ( .B(A[425]), .A(S), .Z(O[425]) );
  ANDN U640 ( .B(A[424]), .A(S), .Z(O[424]) );
  ANDN U641 ( .B(A[423]), .A(S), .Z(O[423]) );
  ANDN U642 ( .B(A[422]), .A(S), .Z(O[422]) );
  ANDN U643 ( .B(A[421]), .A(S), .Z(O[421]) );
  ANDN U644 ( .B(A[420]), .A(S), .Z(O[420]) );
  ANDN U645 ( .B(A[41]), .A(S), .Z(O[41]) );
  ANDN U646 ( .B(A[419]), .A(S), .Z(O[419]) );
  ANDN U647 ( .B(A[418]), .A(S), .Z(O[418]) );
  ANDN U648 ( .B(A[417]), .A(S), .Z(O[417]) );
  ANDN U649 ( .B(A[416]), .A(S), .Z(O[416]) );
  ANDN U650 ( .B(A[415]), .A(S), .Z(O[415]) );
  ANDN U651 ( .B(A[414]), .A(S), .Z(O[414]) );
  ANDN U652 ( .B(A[413]), .A(S), .Z(O[413]) );
  ANDN U653 ( .B(A[412]), .A(S), .Z(O[412]) );
  ANDN U654 ( .B(A[411]), .A(S), .Z(O[411]) );
  ANDN U655 ( .B(A[410]), .A(S), .Z(O[410]) );
  ANDN U656 ( .B(A[40]), .A(S), .Z(O[40]) );
  ANDN U657 ( .B(A[409]), .A(S), .Z(O[409]) );
  ANDN U658 ( .B(A[408]), .A(S), .Z(O[408]) );
  ANDN U659 ( .B(A[407]), .A(S), .Z(O[407]) );
  ANDN U660 ( .B(A[406]), .A(S), .Z(O[406]) );
  ANDN U661 ( .B(A[405]), .A(S), .Z(O[405]) );
  ANDN U662 ( .B(A[404]), .A(S), .Z(O[404]) );
  ANDN U663 ( .B(A[403]), .A(S), .Z(O[403]) );
  ANDN U664 ( .B(A[402]), .A(S), .Z(O[402]) );
  ANDN U665 ( .B(A[401]), .A(S), .Z(O[401]) );
  ANDN U666 ( .B(A[400]), .A(S), .Z(O[400]) );
  ANDN U667 ( .B(A[3]), .A(S), .Z(O[3]) );
  ANDN U668 ( .B(A[39]), .A(S), .Z(O[39]) );
  ANDN U669 ( .B(A[399]), .A(S), .Z(O[399]) );
  ANDN U670 ( .B(A[398]), .A(S), .Z(O[398]) );
  ANDN U671 ( .B(A[397]), .A(S), .Z(O[397]) );
  ANDN U672 ( .B(A[396]), .A(S), .Z(O[396]) );
  ANDN U673 ( .B(A[395]), .A(S), .Z(O[395]) );
  ANDN U674 ( .B(A[394]), .A(S), .Z(O[394]) );
  ANDN U675 ( .B(A[393]), .A(S), .Z(O[393]) );
  ANDN U676 ( .B(A[392]), .A(S), .Z(O[392]) );
  ANDN U677 ( .B(A[391]), .A(S), .Z(O[391]) );
  ANDN U678 ( .B(A[390]), .A(S), .Z(O[390]) );
  ANDN U679 ( .B(A[38]), .A(S), .Z(O[38]) );
  ANDN U680 ( .B(A[389]), .A(S), .Z(O[389]) );
  ANDN U681 ( .B(A[388]), .A(S), .Z(O[388]) );
  ANDN U682 ( .B(A[387]), .A(S), .Z(O[387]) );
  ANDN U683 ( .B(A[386]), .A(S), .Z(O[386]) );
  ANDN U684 ( .B(A[385]), .A(S), .Z(O[385]) );
  ANDN U685 ( .B(A[384]), .A(S), .Z(O[384]) );
  ANDN U686 ( .B(A[383]), .A(S), .Z(O[383]) );
  ANDN U687 ( .B(A[382]), .A(S), .Z(O[382]) );
  ANDN U688 ( .B(A[381]), .A(S), .Z(O[381]) );
  ANDN U689 ( .B(A[380]), .A(S), .Z(O[380]) );
  ANDN U690 ( .B(A[37]), .A(S), .Z(O[37]) );
  ANDN U691 ( .B(A[379]), .A(S), .Z(O[379]) );
  ANDN U692 ( .B(A[378]), .A(S), .Z(O[378]) );
  ANDN U693 ( .B(A[377]), .A(S), .Z(O[377]) );
  ANDN U694 ( .B(A[376]), .A(S), .Z(O[376]) );
  ANDN U695 ( .B(A[375]), .A(S), .Z(O[375]) );
  ANDN U696 ( .B(A[374]), .A(S), .Z(O[374]) );
  ANDN U697 ( .B(A[373]), .A(S), .Z(O[373]) );
  ANDN U698 ( .B(A[372]), .A(S), .Z(O[372]) );
  ANDN U699 ( .B(A[371]), .A(S), .Z(O[371]) );
  ANDN U700 ( .B(A[370]), .A(S), .Z(O[370]) );
  ANDN U701 ( .B(A[36]), .A(S), .Z(O[36]) );
  ANDN U702 ( .B(A[369]), .A(S), .Z(O[369]) );
  ANDN U703 ( .B(A[368]), .A(S), .Z(O[368]) );
  ANDN U704 ( .B(A[367]), .A(S), .Z(O[367]) );
  ANDN U705 ( .B(A[366]), .A(S), .Z(O[366]) );
  ANDN U706 ( .B(A[365]), .A(S), .Z(O[365]) );
  ANDN U707 ( .B(A[364]), .A(S), .Z(O[364]) );
  ANDN U708 ( .B(A[363]), .A(S), .Z(O[363]) );
  ANDN U709 ( .B(A[362]), .A(S), .Z(O[362]) );
  ANDN U710 ( .B(A[361]), .A(S), .Z(O[361]) );
  ANDN U711 ( .B(A[360]), .A(S), .Z(O[360]) );
  ANDN U712 ( .B(A[35]), .A(S), .Z(O[35]) );
  ANDN U713 ( .B(A[359]), .A(S), .Z(O[359]) );
  ANDN U714 ( .B(A[358]), .A(S), .Z(O[358]) );
  ANDN U715 ( .B(A[357]), .A(S), .Z(O[357]) );
  ANDN U716 ( .B(A[356]), .A(S), .Z(O[356]) );
  ANDN U717 ( .B(A[355]), .A(S), .Z(O[355]) );
  ANDN U718 ( .B(A[354]), .A(S), .Z(O[354]) );
  ANDN U719 ( .B(A[353]), .A(S), .Z(O[353]) );
  ANDN U720 ( .B(A[352]), .A(S), .Z(O[352]) );
  ANDN U721 ( .B(A[351]), .A(S), .Z(O[351]) );
  ANDN U722 ( .B(A[350]), .A(S), .Z(O[350]) );
  ANDN U723 ( .B(A[34]), .A(S), .Z(O[34]) );
  ANDN U724 ( .B(A[349]), .A(S), .Z(O[349]) );
  ANDN U725 ( .B(A[348]), .A(S), .Z(O[348]) );
  ANDN U726 ( .B(A[347]), .A(S), .Z(O[347]) );
  ANDN U727 ( .B(A[346]), .A(S), .Z(O[346]) );
  ANDN U728 ( .B(A[345]), .A(S), .Z(O[345]) );
  ANDN U729 ( .B(A[344]), .A(S), .Z(O[344]) );
  ANDN U730 ( .B(A[343]), .A(S), .Z(O[343]) );
  ANDN U731 ( .B(A[342]), .A(S), .Z(O[342]) );
  ANDN U732 ( .B(A[341]), .A(S), .Z(O[341]) );
  ANDN U733 ( .B(A[340]), .A(S), .Z(O[340]) );
  ANDN U734 ( .B(A[33]), .A(S), .Z(O[33]) );
  ANDN U735 ( .B(A[339]), .A(S), .Z(O[339]) );
  ANDN U736 ( .B(A[338]), .A(S), .Z(O[338]) );
  ANDN U737 ( .B(A[337]), .A(S), .Z(O[337]) );
  ANDN U738 ( .B(A[336]), .A(S), .Z(O[336]) );
  ANDN U739 ( .B(A[335]), .A(S), .Z(O[335]) );
  ANDN U740 ( .B(A[334]), .A(S), .Z(O[334]) );
  ANDN U741 ( .B(A[333]), .A(S), .Z(O[333]) );
  ANDN U742 ( .B(A[332]), .A(S), .Z(O[332]) );
  ANDN U743 ( .B(A[331]), .A(S), .Z(O[331]) );
  ANDN U744 ( .B(A[330]), .A(S), .Z(O[330]) );
  ANDN U745 ( .B(A[32]), .A(S), .Z(O[32]) );
  ANDN U746 ( .B(A[329]), .A(S), .Z(O[329]) );
  ANDN U747 ( .B(A[328]), .A(S), .Z(O[328]) );
  ANDN U748 ( .B(A[327]), .A(S), .Z(O[327]) );
  ANDN U749 ( .B(A[326]), .A(S), .Z(O[326]) );
  ANDN U750 ( .B(A[325]), .A(S), .Z(O[325]) );
  ANDN U751 ( .B(A[324]), .A(S), .Z(O[324]) );
  ANDN U752 ( .B(A[323]), .A(S), .Z(O[323]) );
  ANDN U753 ( .B(A[322]), .A(S), .Z(O[322]) );
  ANDN U754 ( .B(A[321]), .A(S), .Z(O[321]) );
  ANDN U755 ( .B(A[320]), .A(S), .Z(O[320]) );
  ANDN U756 ( .B(A[31]), .A(S), .Z(O[31]) );
  ANDN U757 ( .B(A[319]), .A(S), .Z(O[319]) );
  ANDN U758 ( .B(A[318]), .A(S), .Z(O[318]) );
  ANDN U759 ( .B(A[317]), .A(S), .Z(O[317]) );
  ANDN U760 ( .B(A[316]), .A(S), .Z(O[316]) );
  ANDN U761 ( .B(A[315]), .A(S), .Z(O[315]) );
  ANDN U762 ( .B(A[314]), .A(S), .Z(O[314]) );
  ANDN U763 ( .B(A[313]), .A(S), .Z(O[313]) );
  ANDN U764 ( .B(A[312]), .A(S), .Z(O[312]) );
  ANDN U765 ( .B(A[311]), .A(S), .Z(O[311]) );
  ANDN U766 ( .B(A[310]), .A(S), .Z(O[310]) );
  ANDN U767 ( .B(A[30]), .A(S), .Z(O[30]) );
  ANDN U768 ( .B(A[309]), .A(S), .Z(O[309]) );
  ANDN U769 ( .B(A[308]), .A(S), .Z(O[308]) );
  ANDN U770 ( .B(A[307]), .A(S), .Z(O[307]) );
  ANDN U771 ( .B(A[306]), .A(S), .Z(O[306]) );
  ANDN U772 ( .B(A[305]), .A(S), .Z(O[305]) );
  ANDN U773 ( .B(A[304]), .A(S), .Z(O[304]) );
  ANDN U774 ( .B(A[303]), .A(S), .Z(O[303]) );
  ANDN U775 ( .B(A[302]), .A(S), .Z(O[302]) );
  ANDN U776 ( .B(A[301]), .A(S), .Z(O[301]) );
  ANDN U777 ( .B(A[300]), .A(S), .Z(O[300]) );
  ANDN U778 ( .B(A[2]), .A(S), .Z(O[2]) );
  ANDN U779 ( .B(A[29]), .A(S), .Z(O[29]) );
  ANDN U780 ( .B(A[299]), .A(S), .Z(O[299]) );
  ANDN U781 ( .B(A[298]), .A(S), .Z(O[298]) );
  ANDN U782 ( .B(A[297]), .A(S), .Z(O[297]) );
  ANDN U783 ( .B(A[296]), .A(S), .Z(O[296]) );
  ANDN U784 ( .B(A[295]), .A(S), .Z(O[295]) );
  ANDN U785 ( .B(A[294]), .A(S), .Z(O[294]) );
  ANDN U786 ( .B(A[293]), .A(S), .Z(O[293]) );
  ANDN U787 ( .B(A[292]), .A(S), .Z(O[292]) );
  ANDN U788 ( .B(A[291]), .A(S), .Z(O[291]) );
  ANDN U789 ( .B(A[290]), .A(S), .Z(O[290]) );
  ANDN U790 ( .B(A[28]), .A(S), .Z(O[28]) );
  ANDN U791 ( .B(A[289]), .A(S), .Z(O[289]) );
  ANDN U792 ( .B(A[288]), .A(S), .Z(O[288]) );
  ANDN U793 ( .B(A[287]), .A(S), .Z(O[287]) );
  ANDN U794 ( .B(A[286]), .A(S), .Z(O[286]) );
  ANDN U795 ( .B(A[285]), .A(S), .Z(O[285]) );
  ANDN U796 ( .B(A[284]), .A(S), .Z(O[284]) );
  ANDN U797 ( .B(A[283]), .A(S), .Z(O[283]) );
  ANDN U798 ( .B(A[282]), .A(S), .Z(O[282]) );
  ANDN U799 ( .B(A[281]), .A(S), .Z(O[281]) );
  ANDN U800 ( .B(A[280]), .A(S), .Z(O[280]) );
  ANDN U801 ( .B(A[27]), .A(S), .Z(O[27]) );
  ANDN U802 ( .B(A[279]), .A(S), .Z(O[279]) );
  ANDN U803 ( .B(A[278]), .A(S), .Z(O[278]) );
  ANDN U804 ( .B(A[277]), .A(S), .Z(O[277]) );
  ANDN U805 ( .B(A[276]), .A(S), .Z(O[276]) );
  ANDN U806 ( .B(A[275]), .A(S), .Z(O[275]) );
  ANDN U807 ( .B(A[274]), .A(S), .Z(O[274]) );
  ANDN U808 ( .B(A[273]), .A(S), .Z(O[273]) );
  ANDN U809 ( .B(A[272]), .A(S), .Z(O[272]) );
  ANDN U810 ( .B(A[271]), .A(S), .Z(O[271]) );
  ANDN U811 ( .B(A[270]), .A(S), .Z(O[270]) );
  ANDN U812 ( .B(A[26]), .A(S), .Z(O[26]) );
  ANDN U813 ( .B(A[269]), .A(S), .Z(O[269]) );
  ANDN U814 ( .B(A[268]), .A(S), .Z(O[268]) );
  ANDN U815 ( .B(A[267]), .A(S), .Z(O[267]) );
  ANDN U816 ( .B(A[266]), .A(S), .Z(O[266]) );
  ANDN U817 ( .B(A[265]), .A(S), .Z(O[265]) );
  ANDN U818 ( .B(A[264]), .A(S), .Z(O[264]) );
  ANDN U819 ( .B(A[263]), .A(S), .Z(O[263]) );
  ANDN U820 ( .B(A[262]), .A(S), .Z(O[262]) );
  ANDN U821 ( .B(A[261]), .A(S), .Z(O[261]) );
  ANDN U822 ( .B(A[260]), .A(S), .Z(O[260]) );
  ANDN U823 ( .B(A[25]), .A(S), .Z(O[25]) );
  ANDN U824 ( .B(A[259]), .A(S), .Z(O[259]) );
  ANDN U825 ( .B(A[258]), .A(S), .Z(O[258]) );
  ANDN U826 ( .B(A[257]), .A(S), .Z(O[257]) );
  ANDN U827 ( .B(A[256]), .A(S), .Z(O[256]) );
  ANDN U828 ( .B(A[255]), .A(S), .Z(O[255]) );
  ANDN U829 ( .B(A[254]), .A(S), .Z(O[254]) );
  ANDN U830 ( .B(A[253]), .A(S), .Z(O[253]) );
  ANDN U831 ( .B(A[252]), .A(S), .Z(O[252]) );
  ANDN U832 ( .B(A[251]), .A(S), .Z(O[251]) );
  ANDN U833 ( .B(A[250]), .A(S), .Z(O[250]) );
  ANDN U834 ( .B(A[24]), .A(S), .Z(O[24]) );
  ANDN U835 ( .B(A[249]), .A(S), .Z(O[249]) );
  ANDN U836 ( .B(A[248]), .A(S), .Z(O[248]) );
  ANDN U837 ( .B(A[247]), .A(S), .Z(O[247]) );
  ANDN U838 ( .B(A[246]), .A(S), .Z(O[246]) );
  ANDN U839 ( .B(A[245]), .A(S), .Z(O[245]) );
  ANDN U840 ( .B(A[244]), .A(S), .Z(O[244]) );
  ANDN U841 ( .B(A[243]), .A(S), .Z(O[243]) );
  ANDN U842 ( .B(A[242]), .A(S), .Z(O[242]) );
  ANDN U843 ( .B(A[241]), .A(S), .Z(O[241]) );
  ANDN U844 ( .B(A[240]), .A(S), .Z(O[240]) );
  ANDN U845 ( .B(A[23]), .A(S), .Z(O[23]) );
  ANDN U846 ( .B(A[239]), .A(S), .Z(O[239]) );
  ANDN U847 ( .B(A[238]), .A(S), .Z(O[238]) );
  ANDN U848 ( .B(A[237]), .A(S), .Z(O[237]) );
  ANDN U849 ( .B(A[236]), .A(S), .Z(O[236]) );
  ANDN U850 ( .B(A[235]), .A(S), .Z(O[235]) );
  ANDN U851 ( .B(A[234]), .A(S), .Z(O[234]) );
  ANDN U852 ( .B(A[233]), .A(S), .Z(O[233]) );
  ANDN U853 ( .B(A[232]), .A(S), .Z(O[232]) );
  ANDN U854 ( .B(A[231]), .A(S), .Z(O[231]) );
  ANDN U855 ( .B(A[230]), .A(S), .Z(O[230]) );
  ANDN U856 ( .B(A[22]), .A(S), .Z(O[22]) );
  ANDN U857 ( .B(A[229]), .A(S), .Z(O[229]) );
  ANDN U858 ( .B(A[228]), .A(S), .Z(O[228]) );
  ANDN U859 ( .B(A[227]), .A(S), .Z(O[227]) );
  ANDN U860 ( .B(A[226]), .A(S), .Z(O[226]) );
  ANDN U861 ( .B(A[225]), .A(S), .Z(O[225]) );
  ANDN U862 ( .B(A[224]), .A(S), .Z(O[224]) );
  ANDN U863 ( .B(A[223]), .A(S), .Z(O[223]) );
  ANDN U864 ( .B(A[222]), .A(S), .Z(O[222]) );
  ANDN U865 ( .B(A[221]), .A(S), .Z(O[221]) );
  ANDN U866 ( .B(A[220]), .A(S), .Z(O[220]) );
  ANDN U867 ( .B(A[21]), .A(S), .Z(O[21]) );
  ANDN U868 ( .B(A[219]), .A(S), .Z(O[219]) );
  ANDN U869 ( .B(A[218]), .A(S), .Z(O[218]) );
  ANDN U870 ( .B(A[217]), .A(S), .Z(O[217]) );
  ANDN U871 ( .B(A[216]), .A(S), .Z(O[216]) );
  ANDN U872 ( .B(A[215]), .A(S), .Z(O[215]) );
  ANDN U873 ( .B(A[214]), .A(S), .Z(O[214]) );
  ANDN U874 ( .B(A[213]), .A(S), .Z(O[213]) );
  ANDN U875 ( .B(A[212]), .A(S), .Z(O[212]) );
  ANDN U876 ( .B(A[211]), .A(S), .Z(O[211]) );
  ANDN U877 ( .B(A[210]), .A(S), .Z(O[210]) );
  ANDN U878 ( .B(A[20]), .A(S), .Z(O[20]) );
  ANDN U879 ( .B(A[209]), .A(S), .Z(O[209]) );
  ANDN U880 ( .B(A[208]), .A(S), .Z(O[208]) );
  ANDN U881 ( .B(A[207]), .A(S), .Z(O[207]) );
  ANDN U882 ( .B(A[206]), .A(S), .Z(O[206]) );
  ANDN U883 ( .B(A[205]), .A(S), .Z(O[205]) );
  ANDN U884 ( .B(A[204]), .A(S), .Z(O[204]) );
  ANDN U885 ( .B(A[203]), .A(S), .Z(O[203]) );
  ANDN U886 ( .B(A[202]), .A(S), .Z(O[202]) );
  ANDN U887 ( .B(A[201]), .A(S), .Z(O[201]) );
  ANDN U888 ( .B(A[200]), .A(S), .Z(O[200]) );
  ANDN U889 ( .B(A[1]), .A(S), .Z(O[1]) );
  ANDN U890 ( .B(A[19]), .A(S), .Z(O[19]) );
  ANDN U891 ( .B(A[199]), .A(S), .Z(O[199]) );
  ANDN U892 ( .B(A[198]), .A(S), .Z(O[198]) );
  ANDN U893 ( .B(A[197]), .A(S), .Z(O[197]) );
  ANDN U894 ( .B(A[196]), .A(S), .Z(O[196]) );
  ANDN U895 ( .B(A[195]), .A(S), .Z(O[195]) );
  ANDN U896 ( .B(A[194]), .A(S), .Z(O[194]) );
  ANDN U897 ( .B(A[193]), .A(S), .Z(O[193]) );
  ANDN U898 ( .B(A[192]), .A(S), .Z(O[192]) );
  ANDN U899 ( .B(A[191]), .A(S), .Z(O[191]) );
  ANDN U900 ( .B(A[190]), .A(S), .Z(O[190]) );
  ANDN U901 ( .B(A[18]), .A(S), .Z(O[18]) );
  ANDN U902 ( .B(A[189]), .A(S), .Z(O[189]) );
  ANDN U903 ( .B(A[188]), .A(S), .Z(O[188]) );
  ANDN U904 ( .B(A[187]), .A(S), .Z(O[187]) );
  ANDN U905 ( .B(A[186]), .A(S), .Z(O[186]) );
  ANDN U906 ( .B(A[185]), .A(S), .Z(O[185]) );
  ANDN U907 ( .B(A[184]), .A(S), .Z(O[184]) );
  ANDN U908 ( .B(A[183]), .A(S), .Z(O[183]) );
  ANDN U909 ( .B(A[182]), .A(S), .Z(O[182]) );
  ANDN U910 ( .B(A[181]), .A(S), .Z(O[181]) );
  ANDN U911 ( .B(A[180]), .A(S), .Z(O[180]) );
  ANDN U912 ( .B(A[17]), .A(S), .Z(O[17]) );
  ANDN U913 ( .B(A[179]), .A(S), .Z(O[179]) );
  ANDN U914 ( .B(A[178]), .A(S), .Z(O[178]) );
  ANDN U915 ( .B(A[177]), .A(S), .Z(O[177]) );
  ANDN U916 ( .B(A[176]), .A(S), .Z(O[176]) );
  ANDN U917 ( .B(A[175]), .A(S), .Z(O[175]) );
  ANDN U918 ( .B(A[174]), .A(S), .Z(O[174]) );
  ANDN U919 ( .B(A[173]), .A(S), .Z(O[173]) );
  ANDN U920 ( .B(A[172]), .A(S), .Z(O[172]) );
  ANDN U921 ( .B(A[171]), .A(S), .Z(O[171]) );
  ANDN U922 ( .B(A[170]), .A(S), .Z(O[170]) );
  ANDN U923 ( .B(A[16]), .A(S), .Z(O[16]) );
  ANDN U924 ( .B(A[169]), .A(S), .Z(O[169]) );
  ANDN U925 ( .B(A[168]), .A(S), .Z(O[168]) );
  ANDN U926 ( .B(A[167]), .A(S), .Z(O[167]) );
  ANDN U927 ( .B(A[166]), .A(S), .Z(O[166]) );
  ANDN U928 ( .B(A[165]), .A(S), .Z(O[165]) );
  ANDN U929 ( .B(A[164]), .A(S), .Z(O[164]) );
  ANDN U930 ( .B(A[163]), .A(S), .Z(O[163]) );
  ANDN U931 ( .B(A[162]), .A(S), .Z(O[162]) );
  ANDN U932 ( .B(A[161]), .A(S), .Z(O[161]) );
  ANDN U933 ( .B(A[160]), .A(S), .Z(O[160]) );
  ANDN U934 ( .B(A[15]), .A(S), .Z(O[15]) );
  ANDN U935 ( .B(A[159]), .A(S), .Z(O[159]) );
  ANDN U936 ( .B(A[158]), .A(S), .Z(O[158]) );
  ANDN U937 ( .B(A[157]), .A(S), .Z(O[157]) );
  ANDN U938 ( .B(A[156]), .A(S), .Z(O[156]) );
  ANDN U939 ( .B(A[155]), .A(S), .Z(O[155]) );
  ANDN U940 ( .B(A[154]), .A(S), .Z(O[154]) );
  ANDN U941 ( .B(A[153]), .A(S), .Z(O[153]) );
  ANDN U942 ( .B(A[152]), .A(S), .Z(O[152]) );
  ANDN U943 ( .B(A[151]), .A(S), .Z(O[151]) );
  ANDN U944 ( .B(A[150]), .A(S), .Z(O[150]) );
  ANDN U945 ( .B(A[14]), .A(S), .Z(O[14]) );
  ANDN U946 ( .B(A[149]), .A(S), .Z(O[149]) );
  ANDN U947 ( .B(A[148]), .A(S), .Z(O[148]) );
  ANDN U948 ( .B(A[147]), .A(S), .Z(O[147]) );
  ANDN U949 ( .B(A[146]), .A(S), .Z(O[146]) );
  ANDN U950 ( .B(A[145]), .A(S), .Z(O[145]) );
  ANDN U951 ( .B(A[144]), .A(S), .Z(O[144]) );
  ANDN U952 ( .B(A[143]), .A(S), .Z(O[143]) );
  ANDN U953 ( .B(A[142]), .A(S), .Z(O[142]) );
  ANDN U954 ( .B(A[141]), .A(S), .Z(O[141]) );
  ANDN U955 ( .B(A[140]), .A(S), .Z(O[140]) );
  ANDN U956 ( .B(A[13]), .A(S), .Z(O[13]) );
  ANDN U957 ( .B(A[139]), .A(S), .Z(O[139]) );
  ANDN U958 ( .B(A[138]), .A(S), .Z(O[138]) );
  ANDN U959 ( .B(A[137]), .A(S), .Z(O[137]) );
  ANDN U960 ( .B(A[136]), .A(S), .Z(O[136]) );
  ANDN U961 ( .B(A[135]), .A(S), .Z(O[135]) );
  ANDN U962 ( .B(A[134]), .A(S), .Z(O[134]) );
  ANDN U963 ( .B(A[133]), .A(S), .Z(O[133]) );
  ANDN U964 ( .B(A[132]), .A(S), .Z(O[132]) );
  ANDN U965 ( .B(A[131]), .A(S), .Z(O[131]) );
  ANDN U966 ( .B(A[130]), .A(S), .Z(O[130]) );
  ANDN U967 ( .B(A[12]), .A(S), .Z(O[12]) );
  ANDN U968 ( .B(A[129]), .A(S), .Z(O[129]) );
  ANDN U969 ( .B(A[128]), .A(S), .Z(O[128]) );
  ANDN U970 ( .B(A[127]), .A(S), .Z(O[127]) );
  ANDN U971 ( .B(A[126]), .A(S), .Z(O[126]) );
  ANDN U972 ( .B(A[125]), .A(S), .Z(O[125]) );
  ANDN U973 ( .B(A[124]), .A(S), .Z(O[124]) );
  ANDN U974 ( .B(A[123]), .A(S), .Z(O[123]) );
  ANDN U975 ( .B(A[122]), .A(S), .Z(O[122]) );
  ANDN U976 ( .B(A[121]), .A(S), .Z(O[121]) );
  ANDN U977 ( .B(A[120]), .A(S), .Z(O[120]) );
  ANDN U978 ( .B(A[11]), .A(S), .Z(O[11]) );
  ANDN U979 ( .B(A[119]), .A(S), .Z(O[119]) );
  ANDN U980 ( .B(A[118]), .A(S), .Z(O[118]) );
  ANDN U981 ( .B(A[117]), .A(S), .Z(O[117]) );
  ANDN U982 ( .B(A[116]), .A(S), .Z(O[116]) );
  ANDN U983 ( .B(A[115]), .A(S), .Z(O[115]) );
  ANDN U984 ( .B(A[114]), .A(S), .Z(O[114]) );
  ANDN U985 ( .B(A[113]), .A(S), .Z(O[113]) );
  ANDN U986 ( .B(A[112]), .A(S), .Z(O[112]) );
  ANDN U987 ( .B(A[111]), .A(S), .Z(O[111]) );
  ANDN U988 ( .B(A[110]), .A(S), .Z(O[110]) );
  ANDN U989 ( .B(A[10]), .A(S), .Z(O[10]) );
  ANDN U990 ( .B(A[109]), .A(S), .Z(O[109]) );
  ANDN U991 ( .B(A[108]), .A(S), .Z(O[108]) );
  ANDN U992 ( .B(A[107]), .A(S), .Z(O[107]) );
  ANDN U993 ( .B(A[106]), .A(S), .Z(O[106]) );
  ANDN U994 ( .B(A[105]), .A(S), .Z(O[105]) );
  ANDN U995 ( .B(A[104]), .A(S), .Z(O[104]) );
  ANDN U996 ( .B(A[103]), .A(S), .Z(O[103]) );
  ANDN U997 ( .B(A[102]), .A(S), .Z(O[102]) );
  ANDN U998 ( .B(A[1023]), .A(S), .Z(O[1023]) );
  ANDN U999 ( .B(A[1022]), .A(S), .Z(O[1022]) );
  ANDN U1000 ( .B(A[1021]), .A(S), .Z(O[1021]) );
  ANDN U1001 ( .B(A[1020]), .A(S), .Z(O[1020]) );
  ANDN U1002 ( .B(A[101]), .A(S), .Z(O[101]) );
  ANDN U1003 ( .B(A[1019]), .A(S), .Z(O[1019]) );
  ANDN U1004 ( .B(A[1018]), .A(S), .Z(O[1018]) );
  ANDN U1005 ( .B(A[1017]), .A(S), .Z(O[1017]) );
  ANDN U1006 ( .B(A[1016]), .A(S), .Z(O[1016]) );
  ANDN U1007 ( .B(A[1015]), .A(S), .Z(O[1015]) );
  ANDN U1008 ( .B(A[1014]), .A(S), .Z(O[1014]) );
  ANDN U1009 ( .B(A[1013]), .A(S), .Z(O[1013]) );
  ANDN U1010 ( .B(A[1012]), .A(S), .Z(O[1012]) );
  ANDN U1011 ( .B(A[1011]), .A(S), .Z(O[1011]) );
  ANDN U1012 ( .B(A[1010]), .A(S), .Z(O[1010]) );
  ANDN U1013 ( .B(A[100]), .A(S), .Z(O[100]) );
  ANDN U1014 ( .B(A[1009]), .A(S), .Z(O[1009]) );
  ANDN U1015 ( .B(A[1008]), .A(S), .Z(O[1008]) );
  ANDN U1016 ( .B(A[1007]), .A(S), .Z(O[1007]) );
  ANDN U1017 ( .B(A[1006]), .A(S), .Z(O[1006]) );
  ANDN U1018 ( .B(A[1005]), .A(S), .Z(O[1005]) );
  ANDN U1019 ( .B(A[1004]), .A(S), .Z(O[1004]) );
  ANDN U1020 ( .B(A[1003]), .A(S), .Z(O[1003]) );
  ANDN U1021 ( .B(A[1002]), .A(S), .Z(O[1002]) );
  ANDN U1022 ( .B(A[1001]), .A(S), .Z(O[1001]) );
  ANDN U1023 ( .B(A[1000]), .A(S), .Z(O[1000]) );
  ANDN U1024 ( .B(A[0]), .A(S), .Z(O[0]) );
endmodule


module FA_12601 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  AND U1 ( .A(CI), .B(B), .Z(CO) );
endmodule


module FA_12602 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  AND U1 ( .A(CI), .B(B), .Z(CO) );
endmodule


module FA_12603 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12604 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12605 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12606 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12607 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12608 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12609 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12610 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12611 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12612 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12613 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12614 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12615 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12616 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12617 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12618 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12619 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12620 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12621 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12622 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12623 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12624 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12625 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12626 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12627 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12628 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12629 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12630 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12631 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12632 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12633 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12634 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12635 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12636 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12637 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12638 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12639 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12640 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12641 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12642 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12643 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12644 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12645 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12646 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12647 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12648 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12649 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12650 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12651 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12652 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12653 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12654 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12655 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12656 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12657 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12658 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12659 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12660 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12661 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12662 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12663 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12664 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12665 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12666 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12667 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12668 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12669 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12670 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12671 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12672 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12673 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12674 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12675 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12676 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12677 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12678 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12679 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12680 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12681 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12682 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12683 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12684 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12685 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12686 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12687 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12688 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12689 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12690 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12691 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12692 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12693 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12694 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12695 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12696 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12697 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12698 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12699 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12700 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12701 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12702 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12703 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12704 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12705 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12706 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12707 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12708 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12709 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12710 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12711 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12712 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12713 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12714 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12715 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12716 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12717 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12718 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12719 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12720 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12721 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12722 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12723 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12724 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12725 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12726 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12727 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12728 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12729 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12730 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12731 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12732 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12733 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12734 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12735 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12736 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12737 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12738 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12739 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12740 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12741 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12742 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12743 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12744 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12745 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12746 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12747 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12748 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12749 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12750 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12751 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12752 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12753 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12754 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12755 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12756 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12757 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12758 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12759 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12760 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12761 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12762 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12763 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12764 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12765 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12766 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12767 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12768 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12769 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12770 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12771 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12772 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12773 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12774 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12775 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12776 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12777 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12778 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12779 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12780 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12781 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12782 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12783 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12784 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12785 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12786 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12787 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12788 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12789 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12790 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12791 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12792 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12793 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12794 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12795 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12796 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12797 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12798 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12799 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12800 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12801 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12802 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12803 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12804 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12805 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12806 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12807 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12808 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12809 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12810 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12811 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12812 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12813 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12814 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12815 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12816 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12817 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12818 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12819 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12820 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12821 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12822 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12823 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12824 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12825 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12826 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12827 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12828 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12829 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12830 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12831 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12832 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12833 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12834 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12835 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12836 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12837 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12838 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12839 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12840 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12841 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12842 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12843 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12844 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12845 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12846 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12847 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12848 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12849 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12850 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12851 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12852 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12853 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12854 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12855 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12856 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12857 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12858 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12859 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12860 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12861 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12862 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12863 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12864 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12865 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12866 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12867 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12868 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12869 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12870 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12871 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12872 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12873 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12874 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12875 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12876 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12877 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12878 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12879 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12880 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12881 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12882 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12883 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12884 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12885 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12886 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12887 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12888 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12889 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12890 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12891 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12892 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12893 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12894 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12895 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12896 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12897 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12898 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12899 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12900 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12901 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12902 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12903 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12904 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12905 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12906 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12907 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12908 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12909 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12910 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12911 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12912 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12913 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12914 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12915 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12916 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12917 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12918 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12919 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12920 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12921 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12922 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12923 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12924 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12925 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12926 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12927 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12928 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12929 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12930 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12931 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12932 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12933 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12934 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12935 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12936 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12937 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12938 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12939 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12940 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12941 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12942 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12943 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12944 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12945 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12946 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12947 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12948 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12949 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12950 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12951 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12952 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12953 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12954 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12955 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12956 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12957 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12958 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12959 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12960 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12961 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12962 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12963 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12964 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12965 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12966 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12967 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12968 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12969 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12970 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12971 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12972 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12973 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12974 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12975 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12976 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12977 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12978 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12979 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12980 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12981 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12982 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12983 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12984 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12985 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12986 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12987 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12988 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12989 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12990 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12991 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12992 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12993 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12994 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12995 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12996 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12997 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12998 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_12999 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13000 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13001 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13002 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13003 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13004 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13005 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13006 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13007 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13008 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13009 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13010 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13011 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13012 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13013 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13014 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13015 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13016 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13017 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13018 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13019 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13020 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13021 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13022 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13023 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13024 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13025 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13026 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13027 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13028 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13029 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13030 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13031 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13032 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13033 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13034 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13035 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13036 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13037 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13038 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13039 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13040 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13041 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13042 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13043 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13044 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13045 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13046 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13047 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13048 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13049 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13050 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13051 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13052 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13053 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13054 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13055 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13056 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13057 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13058 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13059 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13060 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13061 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13062 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13063 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13064 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13065 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13066 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13067 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13068 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13069 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13070 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13071 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13072 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13073 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13074 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13075 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13076 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13077 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13078 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13079 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13080 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13081 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13082 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13083 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13084 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13085 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13086 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13087 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13088 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13089 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13090 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13091 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13092 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13093 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13094 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13095 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13096 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13097 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13098 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13099 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13100 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13101 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13102 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13103 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13104 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13105 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13106 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13107 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13108 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13109 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13110 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13111 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13112 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13113 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13114 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13115 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13116 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13117 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13118 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13119 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13120 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13121 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13122 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13123 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13124 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13125 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13126 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13127 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13128 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13129 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13130 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13131 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13132 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13133 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13134 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13135 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13136 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13137 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13138 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13139 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13140 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13141 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13142 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13143 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13144 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13145 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13146 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13147 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13148 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13149 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13150 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13151 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13152 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13153 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13154 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13155 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13156 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13157 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13158 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13159 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13160 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13161 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13162 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13163 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13164 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13165 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13166 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13167 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13168 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13169 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13170 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13171 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13172 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13173 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13174 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13175 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13176 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13177 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13178 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13179 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13180 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13181 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13182 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13183 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13184 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13185 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13186 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13187 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13188 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13189 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13190 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13191 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13192 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13193 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13194 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13195 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13196 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13197 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13198 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13199 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13200 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13201 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13202 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13203 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13204 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13205 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13206 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13207 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13208 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13209 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13210 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13211 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13212 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13213 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13214 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13215 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13216 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13217 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13218 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13219 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13220 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13221 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13222 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13223 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13224 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13225 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13226 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13227 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13228 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13229 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13230 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13231 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13232 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13233 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13234 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13235 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13236 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13237 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13238 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13239 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13240 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13241 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13242 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13243 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13244 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13245 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13246 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13247 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13248 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13249 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13250 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13251 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13252 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13253 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13254 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13255 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13256 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13257 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13258 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13259 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13260 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13261 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13262 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13263 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13264 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13265 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13266 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13267 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13268 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13269 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13270 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13271 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13272 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13273 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13274 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13275 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13276 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13277 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13278 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13279 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13280 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13281 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13282 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13283 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13284 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13285 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13286 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13287 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13288 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13289 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13290 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13291 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13292 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13293 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13294 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13295 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13296 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13297 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13298 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13299 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13300 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13301 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13302 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13303 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13304 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13305 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13306 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13307 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13308 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13309 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13310 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13311 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13312 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13313 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13314 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13315 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13316 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13317 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13318 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13319 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13320 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13321 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13322 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13323 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13324 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13325 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13326 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13327 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13328 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13329 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13330 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13331 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13332 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13333 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13334 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13335 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13336 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13337 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13338 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13339 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13340 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13341 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13342 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13343 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13344 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13345 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13346 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13347 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13348 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13349 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13350 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13351 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13352 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13353 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13354 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13355 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13356 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13357 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13358 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13359 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13360 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13361 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13362 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13363 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13364 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13365 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13366 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13367 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13368 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13369 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13370 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13371 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13372 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13373 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13374 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13375 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13376 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13377 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13378 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13379 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13380 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13381 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13382 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13383 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13384 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13385 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13386 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13387 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13388 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13389 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13390 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13391 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13392 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13393 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13394 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13395 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13396 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13397 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13398 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13399 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13400 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13401 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13402 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13403 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13404 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13405 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13406 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13407 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13408 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13409 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13410 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13411 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13412 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13413 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13414 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13415 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13416 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13417 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13418 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13419 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13420 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13421 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13422 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13423 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13424 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13425 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13426 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13427 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13428 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13429 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13430 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13431 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13432 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13433 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13434 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13435 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13436 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13437 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13438 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13439 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13440 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13441 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13442 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13443 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13444 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13445 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13446 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13447 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13448 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13449 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13450 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13451 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13452 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13453 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13454 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13455 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13456 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13457 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13458 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13459 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13460 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13461 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13462 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13463 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13464 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13465 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13466 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13467 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13468 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13469 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13470 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13471 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13472 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13473 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13474 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13475 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13476 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13477 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13478 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13479 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13480 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13481 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13482 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13483 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13484 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13485 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13486 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13487 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13488 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13489 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13490 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13491 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13492 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13493 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13494 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13495 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13496 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13497 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13498 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13499 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13500 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13501 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13502 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13503 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13504 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13505 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13506 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13507 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13508 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13509 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13510 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13511 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13512 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13513 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13514 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13515 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13516 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13517 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13518 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13519 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13520 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13521 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13522 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13523 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13524 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13525 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13526 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13527 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13528 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13529 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13530 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13531 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13532 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13533 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13534 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13535 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13536 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13537 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13538 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13539 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13540 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13541 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13542 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13543 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13544 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13545 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13546 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13547 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13548 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13549 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13550 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13551 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13552 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13553 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13554 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13555 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13556 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13557 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13558 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13559 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13560 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13561 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13562 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13563 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13564 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13565 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13566 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13567 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13568 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13569 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13570 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13571 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13572 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13573 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13574 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13575 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13576 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13577 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13578 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13579 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13580 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13581 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13582 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13583 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13584 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13585 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13586 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13587 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13588 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13589 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13590 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13591 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13592 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13593 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13594 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13595 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13596 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13597 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13598 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13599 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13600 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13601 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13602 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13603 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13604 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13605 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13606 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13607 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13608 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13609 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13610 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13611 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13612 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13613 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13614 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13615 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13616 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13617 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13618 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13619 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13620 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13621 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13622 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13623 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13624 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13625 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_13626 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  OR U1 ( .A(B), .B(A), .Z(CO) );
endmodule


module COMP_N1026_1 ( A, B, O );
  input [1025:0] A;
  input [1025:0] B;
  output O;
  wire   n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
         n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
         n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
         n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
         n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
         n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
         n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
         n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
         n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
         n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
         n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
         n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
         n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
         n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
         n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
         n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
         n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
         n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
         n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
         n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
         n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
         n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
         n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
         n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
         n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
         n2048, n2049, n2050, n2051, n2052, n2053;
  wire   [1025:1] C;

  FA_13626 \FA_INST_0[0].FA_INST_1[0].FA_  ( .A(A[0]), .B(n1028), .CI(1'b1), 
        .CO(C[1]) );
  FA_13625 \FA_INST_0[0].FA_INST_1[1].FA_  ( .A(A[1]), .B(n1029), .CI(C[1]), 
        .CO(C[2]) );
  FA_13624 \FA_INST_0[0].FA_INST_1[2].FA_  ( .A(A[2]), .B(n1030), .CI(C[2]), 
        .CO(C[3]) );
  FA_13623 \FA_INST_0[0].FA_INST_1[3].FA_  ( .A(A[3]), .B(n1031), .CI(C[3]), 
        .CO(C[4]) );
  FA_13622 \FA_INST_0[0].FA_INST_1[4].FA_  ( .A(A[4]), .B(n1032), .CI(C[4]), 
        .CO(C[5]) );
  FA_13621 \FA_INST_0[0].FA_INST_1[5].FA_  ( .A(A[5]), .B(n1033), .CI(C[5]), 
        .CO(C[6]) );
  FA_13620 \FA_INST_0[0].FA_INST_1[6].FA_  ( .A(A[6]), .B(n1034), .CI(C[6]), 
        .CO(C[7]) );
  FA_13619 \FA_INST_0[0].FA_INST_1[7].FA_  ( .A(A[7]), .B(n1035), .CI(C[7]), 
        .CO(C[8]) );
  FA_13618 \FA_INST_0[0].FA_INST_1[8].FA_  ( .A(A[8]), .B(n1036), .CI(C[8]), 
        .CO(C[9]) );
  FA_13617 \FA_INST_0[0].FA_INST_1[9].FA_  ( .A(A[9]), .B(n1037), .CI(C[9]), 
        .CO(C[10]) );
  FA_13616 \FA_INST_0[0].FA_INST_1[10].FA_  ( .A(A[10]), .B(n1038), .CI(C[10]), 
        .CO(C[11]) );
  FA_13615 \FA_INST_0[0].FA_INST_1[11].FA_  ( .A(A[11]), .B(n1039), .CI(C[11]), 
        .CO(C[12]) );
  FA_13614 \FA_INST_0[0].FA_INST_1[12].FA_  ( .A(A[12]), .B(n1040), .CI(C[12]), 
        .CO(C[13]) );
  FA_13613 \FA_INST_0[0].FA_INST_1[13].FA_  ( .A(A[13]), .B(n1041), .CI(C[13]), 
        .CO(C[14]) );
  FA_13612 \FA_INST_0[0].FA_INST_1[14].FA_  ( .A(A[14]), .B(n1042), .CI(C[14]), 
        .CO(C[15]) );
  FA_13611 \FA_INST_0[0].FA_INST_1[15].FA_  ( .A(A[15]), .B(n1043), .CI(C[15]), 
        .CO(C[16]) );
  FA_13610 \FA_INST_0[0].FA_INST_1[16].FA_  ( .A(A[16]), .B(n1044), .CI(C[16]), 
        .CO(C[17]) );
  FA_13609 \FA_INST_0[0].FA_INST_1[17].FA_  ( .A(A[17]), .B(n1045), .CI(C[17]), 
        .CO(C[18]) );
  FA_13608 \FA_INST_0[0].FA_INST_1[18].FA_  ( .A(A[18]), .B(n1046), .CI(C[18]), 
        .CO(C[19]) );
  FA_13607 \FA_INST_0[0].FA_INST_1[19].FA_  ( .A(A[19]), .B(n1047), .CI(C[19]), 
        .CO(C[20]) );
  FA_13606 \FA_INST_0[0].FA_INST_1[20].FA_  ( .A(A[20]), .B(n1048), .CI(C[20]), 
        .CO(C[21]) );
  FA_13605 \FA_INST_0[0].FA_INST_1[21].FA_  ( .A(A[21]), .B(n1049), .CI(C[21]), 
        .CO(C[22]) );
  FA_13604 \FA_INST_0[0].FA_INST_1[22].FA_  ( .A(A[22]), .B(n1050), .CI(C[22]), 
        .CO(C[23]) );
  FA_13603 \FA_INST_0[0].FA_INST_1[23].FA_  ( .A(A[23]), .B(n1051), .CI(C[23]), 
        .CO(C[24]) );
  FA_13602 \FA_INST_0[0].FA_INST_1[24].FA_  ( .A(A[24]), .B(n1052), .CI(C[24]), 
        .CO(C[25]) );
  FA_13601 \FA_INST_0[0].FA_INST_1[25].FA_  ( .A(A[25]), .B(n1053), .CI(C[25]), 
        .CO(C[26]) );
  FA_13600 \FA_INST_0[0].FA_INST_1[26].FA_  ( .A(A[26]), .B(n1054), .CI(C[26]), 
        .CO(C[27]) );
  FA_13599 \FA_INST_0[0].FA_INST_1[27].FA_  ( .A(A[27]), .B(n1055), .CI(C[27]), 
        .CO(C[28]) );
  FA_13598 \FA_INST_0[0].FA_INST_1[28].FA_  ( .A(A[28]), .B(n1056), .CI(C[28]), 
        .CO(C[29]) );
  FA_13597 \FA_INST_0[0].FA_INST_1[29].FA_  ( .A(A[29]), .B(n1057), .CI(C[29]), 
        .CO(C[30]) );
  FA_13596 \FA_INST_0[0].FA_INST_1[30].FA_  ( .A(A[30]), .B(n1058), .CI(C[30]), 
        .CO(C[31]) );
  FA_13595 \FA_INST_0[0].FA_INST_1[31].FA_  ( .A(A[31]), .B(n1059), .CI(C[31]), 
        .CO(C[32]) );
  FA_13594 \FA_INST_0[0].FA_INST_1[32].FA_  ( .A(A[32]), .B(n1060), .CI(C[32]), 
        .CO(C[33]) );
  FA_13593 \FA_INST_0[0].FA_INST_1[33].FA_  ( .A(A[33]), .B(n1061), .CI(C[33]), 
        .CO(C[34]) );
  FA_13592 \FA_INST_0[0].FA_INST_1[34].FA_  ( .A(A[34]), .B(n1062), .CI(C[34]), 
        .CO(C[35]) );
  FA_13591 \FA_INST_0[0].FA_INST_1[35].FA_  ( .A(A[35]), .B(n1063), .CI(C[35]), 
        .CO(C[36]) );
  FA_13590 \FA_INST_0[0].FA_INST_1[36].FA_  ( .A(A[36]), .B(n1064), .CI(C[36]), 
        .CO(C[37]) );
  FA_13589 \FA_INST_0[0].FA_INST_1[37].FA_  ( .A(A[37]), .B(n1065), .CI(C[37]), 
        .CO(C[38]) );
  FA_13588 \FA_INST_0[0].FA_INST_1[38].FA_  ( .A(A[38]), .B(n1066), .CI(C[38]), 
        .CO(C[39]) );
  FA_13587 \FA_INST_0[0].FA_INST_1[39].FA_  ( .A(A[39]), .B(n1067), .CI(C[39]), 
        .CO(C[40]) );
  FA_13586 \FA_INST_0[0].FA_INST_1[40].FA_  ( .A(A[40]), .B(n1068), .CI(C[40]), 
        .CO(C[41]) );
  FA_13585 \FA_INST_0[0].FA_INST_1[41].FA_  ( .A(A[41]), .B(n1069), .CI(C[41]), 
        .CO(C[42]) );
  FA_13584 \FA_INST_0[0].FA_INST_1[42].FA_  ( .A(A[42]), .B(n1070), .CI(C[42]), 
        .CO(C[43]) );
  FA_13583 \FA_INST_0[0].FA_INST_1[43].FA_  ( .A(A[43]), .B(n1071), .CI(C[43]), 
        .CO(C[44]) );
  FA_13582 \FA_INST_0[0].FA_INST_1[44].FA_  ( .A(A[44]), .B(n1072), .CI(C[44]), 
        .CO(C[45]) );
  FA_13581 \FA_INST_0[0].FA_INST_1[45].FA_  ( .A(A[45]), .B(n1073), .CI(C[45]), 
        .CO(C[46]) );
  FA_13580 \FA_INST_0[0].FA_INST_1[46].FA_  ( .A(A[46]), .B(n1074), .CI(C[46]), 
        .CO(C[47]) );
  FA_13579 \FA_INST_0[0].FA_INST_1[47].FA_  ( .A(A[47]), .B(n1075), .CI(C[47]), 
        .CO(C[48]) );
  FA_13578 \FA_INST_0[0].FA_INST_1[48].FA_  ( .A(A[48]), .B(n1076), .CI(C[48]), 
        .CO(C[49]) );
  FA_13577 \FA_INST_0[0].FA_INST_1[49].FA_  ( .A(A[49]), .B(n1077), .CI(C[49]), 
        .CO(C[50]) );
  FA_13576 \FA_INST_0[0].FA_INST_1[50].FA_  ( .A(A[50]), .B(n1078), .CI(C[50]), 
        .CO(C[51]) );
  FA_13575 \FA_INST_0[0].FA_INST_1[51].FA_  ( .A(A[51]), .B(n1079), .CI(C[51]), 
        .CO(C[52]) );
  FA_13574 \FA_INST_0[0].FA_INST_1[52].FA_  ( .A(A[52]), .B(n1080), .CI(C[52]), 
        .CO(C[53]) );
  FA_13573 \FA_INST_0[0].FA_INST_1[53].FA_  ( .A(A[53]), .B(n1081), .CI(C[53]), 
        .CO(C[54]) );
  FA_13572 \FA_INST_0[0].FA_INST_1[54].FA_  ( .A(A[54]), .B(n1082), .CI(C[54]), 
        .CO(C[55]) );
  FA_13571 \FA_INST_0[0].FA_INST_1[55].FA_  ( .A(A[55]), .B(n1083), .CI(C[55]), 
        .CO(C[56]) );
  FA_13570 \FA_INST_0[0].FA_INST_1[56].FA_  ( .A(A[56]), .B(n1084), .CI(C[56]), 
        .CO(C[57]) );
  FA_13569 \FA_INST_0[0].FA_INST_1[57].FA_  ( .A(A[57]), .B(n1085), .CI(C[57]), 
        .CO(C[58]) );
  FA_13568 \FA_INST_0[0].FA_INST_1[58].FA_  ( .A(A[58]), .B(n1086), .CI(C[58]), 
        .CO(C[59]) );
  FA_13567 \FA_INST_0[0].FA_INST_1[59].FA_  ( .A(A[59]), .B(n1087), .CI(C[59]), 
        .CO(C[60]) );
  FA_13566 \FA_INST_0[0].FA_INST_1[60].FA_  ( .A(A[60]), .B(n1088), .CI(C[60]), 
        .CO(C[61]) );
  FA_13565 \FA_INST_0[0].FA_INST_1[61].FA_  ( .A(A[61]), .B(n1089), .CI(C[61]), 
        .CO(C[62]) );
  FA_13564 \FA_INST_0[0].FA_INST_1[62].FA_  ( .A(A[62]), .B(n1090), .CI(C[62]), 
        .CO(C[63]) );
  FA_13563 \FA_INST_0[0].FA_INST_1[63].FA_  ( .A(A[63]), .B(n1091), .CI(C[63]), 
        .CO(C[64]) );
  FA_13562 \FA_INST_0[0].FA_INST_1[64].FA_  ( .A(A[64]), .B(n1092), .CI(C[64]), 
        .CO(C[65]) );
  FA_13561 \FA_INST_0[0].FA_INST_1[65].FA_  ( .A(A[65]), .B(n1093), .CI(C[65]), 
        .CO(C[66]) );
  FA_13560 \FA_INST_0[0].FA_INST_1[66].FA_  ( .A(A[66]), .B(n1094), .CI(C[66]), 
        .CO(C[67]) );
  FA_13559 \FA_INST_0[0].FA_INST_1[67].FA_  ( .A(A[67]), .B(n1095), .CI(C[67]), 
        .CO(C[68]) );
  FA_13558 \FA_INST_0[0].FA_INST_1[68].FA_  ( .A(A[68]), .B(n1096), .CI(C[68]), 
        .CO(C[69]) );
  FA_13557 \FA_INST_0[0].FA_INST_1[69].FA_  ( .A(A[69]), .B(n1097), .CI(C[69]), 
        .CO(C[70]) );
  FA_13556 \FA_INST_0[0].FA_INST_1[70].FA_  ( .A(A[70]), .B(n1098), .CI(C[70]), 
        .CO(C[71]) );
  FA_13555 \FA_INST_0[0].FA_INST_1[71].FA_  ( .A(A[71]), .B(n1099), .CI(C[71]), 
        .CO(C[72]) );
  FA_13554 \FA_INST_0[0].FA_INST_1[72].FA_  ( .A(A[72]), .B(n1100), .CI(C[72]), 
        .CO(C[73]) );
  FA_13553 \FA_INST_0[0].FA_INST_1[73].FA_  ( .A(A[73]), .B(n1101), .CI(C[73]), 
        .CO(C[74]) );
  FA_13552 \FA_INST_0[0].FA_INST_1[74].FA_  ( .A(A[74]), .B(n1102), .CI(C[74]), 
        .CO(C[75]) );
  FA_13551 \FA_INST_0[0].FA_INST_1[75].FA_  ( .A(A[75]), .B(n1103), .CI(C[75]), 
        .CO(C[76]) );
  FA_13550 \FA_INST_0[0].FA_INST_1[76].FA_  ( .A(A[76]), .B(n1104), .CI(C[76]), 
        .CO(C[77]) );
  FA_13549 \FA_INST_0[0].FA_INST_1[77].FA_  ( .A(A[77]), .B(n1105), .CI(C[77]), 
        .CO(C[78]) );
  FA_13548 \FA_INST_0[0].FA_INST_1[78].FA_  ( .A(A[78]), .B(n1106), .CI(C[78]), 
        .CO(C[79]) );
  FA_13547 \FA_INST_0[0].FA_INST_1[79].FA_  ( .A(A[79]), .B(n1107), .CI(C[79]), 
        .CO(C[80]) );
  FA_13546 \FA_INST_0[0].FA_INST_1[80].FA_  ( .A(A[80]), .B(n1108), .CI(C[80]), 
        .CO(C[81]) );
  FA_13545 \FA_INST_0[0].FA_INST_1[81].FA_  ( .A(A[81]), .B(n1109), .CI(C[81]), 
        .CO(C[82]) );
  FA_13544 \FA_INST_0[0].FA_INST_1[82].FA_  ( .A(A[82]), .B(n1110), .CI(C[82]), 
        .CO(C[83]) );
  FA_13543 \FA_INST_0[0].FA_INST_1[83].FA_  ( .A(A[83]), .B(n1111), .CI(C[83]), 
        .CO(C[84]) );
  FA_13542 \FA_INST_0[0].FA_INST_1[84].FA_  ( .A(A[84]), .B(n1112), .CI(C[84]), 
        .CO(C[85]) );
  FA_13541 \FA_INST_0[0].FA_INST_1[85].FA_  ( .A(A[85]), .B(n1113), .CI(C[85]), 
        .CO(C[86]) );
  FA_13540 \FA_INST_0[0].FA_INST_1[86].FA_  ( .A(A[86]), .B(n1114), .CI(C[86]), 
        .CO(C[87]) );
  FA_13539 \FA_INST_0[0].FA_INST_1[87].FA_  ( .A(A[87]), .B(n1115), .CI(C[87]), 
        .CO(C[88]) );
  FA_13538 \FA_INST_0[0].FA_INST_1[88].FA_  ( .A(A[88]), .B(n1116), .CI(C[88]), 
        .CO(C[89]) );
  FA_13537 \FA_INST_0[0].FA_INST_1[89].FA_  ( .A(A[89]), .B(n1117), .CI(C[89]), 
        .CO(C[90]) );
  FA_13536 \FA_INST_0[0].FA_INST_1[90].FA_  ( .A(A[90]), .B(n1118), .CI(C[90]), 
        .CO(C[91]) );
  FA_13535 \FA_INST_0[0].FA_INST_1[91].FA_  ( .A(A[91]), .B(n1119), .CI(C[91]), 
        .CO(C[92]) );
  FA_13534 \FA_INST_0[0].FA_INST_1[92].FA_  ( .A(A[92]), .B(n1120), .CI(C[92]), 
        .CO(C[93]) );
  FA_13533 \FA_INST_0[0].FA_INST_1[93].FA_  ( .A(A[93]), .B(n1121), .CI(C[93]), 
        .CO(C[94]) );
  FA_13532 \FA_INST_0[0].FA_INST_1[94].FA_  ( .A(A[94]), .B(n1122), .CI(C[94]), 
        .CO(C[95]) );
  FA_13531 \FA_INST_0[0].FA_INST_1[95].FA_  ( .A(A[95]), .B(n1123), .CI(C[95]), 
        .CO(C[96]) );
  FA_13530 \FA_INST_0[0].FA_INST_1[96].FA_  ( .A(A[96]), .B(n1124), .CI(C[96]), 
        .CO(C[97]) );
  FA_13529 \FA_INST_0[0].FA_INST_1[97].FA_  ( .A(A[97]), .B(n1125), .CI(C[97]), 
        .CO(C[98]) );
  FA_13528 \FA_INST_0[0].FA_INST_1[98].FA_  ( .A(A[98]), .B(n1126), .CI(C[98]), 
        .CO(C[99]) );
  FA_13527 \FA_INST_0[0].FA_INST_1[99].FA_  ( .A(A[99]), .B(n1127), .CI(C[99]), 
        .CO(C[100]) );
  FA_13526 \FA_INST_0[0].FA_INST_1[100].FA_  ( .A(A[100]), .B(n1128), .CI(
        C[100]), .CO(C[101]) );
  FA_13525 \FA_INST_0[0].FA_INST_1[101].FA_  ( .A(A[101]), .B(n1129), .CI(
        C[101]), .CO(C[102]) );
  FA_13524 \FA_INST_0[0].FA_INST_1[102].FA_  ( .A(A[102]), .B(n1130), .CI(
        C[102]), .CO(C[103]) );
  FA_13523 \FA_INST_0[0].FA_INST_1[103].FA_  ( .A(A[103]), .B(n1131), .CI(
        C[103]), .CO(C[104]) );
  FA_13522 \FA_INST_0[0].FA_INST_1[104].FA_  ( .A(A[104]), .B(n1132), .CI(
        C[104]), .CO(C[105]) );
  FA_13521 \FA_INST_0[0].FA_INST_1[105].FA_  ( .A(A[105]), .B(n1133), .CI(
        C[105]), .CO(C[106]) );
  FA_13520 \FA_INST_0[0].FA_INST_1[106].FA_  ( .A(A[106]), .B(n1134), .CI(
        C[106]), .CO(C[107]) );
  FA_13519 \FA_INST_0[0].FA_INST_1[107].FA_  ( .A(A[107]), .B(n1135), .CI(
        C[107]), .CO(C[108]) );
  FA_13518 \FA_INST_0[0].FA_INST_1[108].FA_  ( .A(A[108]), .B(n1136), .CI(
        C[108]), .CO(C[109]) );
  FA_13517 \FA_INST_0[0].FA_INST_1[109].FA_  ( .A(A[109]), .B(n1137), .CI(
        C[109]), .CO(C[110]) );
  FA_13516 \FA_INST_0[0].FA_INST_1[110].FA_  ( .A(A[110]), .B(n1138), .CI(
        C[110]), .CO(C[111]) );
  FA_13515 \FA_INST_0[0].FA_INST_1[111].FA_  ( .A(A[111]), .B(n1139), .CI(
        C[111]), .CO(C[112]) );
  FA_13514 \FA_INST_0[0].FA_INST_1[112].FA_  ( .A(A[112]), .B(n1140), .CI(
        C[112]), .CO(C[113]) );
  FA_13513 \FA_INST_0[0].FA_INST_1[113].FA_  ( .A(A[113]), .B(n1141), .CI(
        C[113]), .CO(C[114]) );
  FA_13512 \FA_INST_0[0].FA_INST_1[114].FA_  ( .A(A[114]), .B(n1142), .CI(
        C[114]), .CO(C[115]) );
  FA_13511 \FA_INST_0[0].FA_INST_1[115].FA_  ( .A(A[115]), .B(n1143), .CI(
        C[115]), .CO(C[116]) );
  FA_13510 \FA_INST_0[0].FA_INST_1[116].FA_  ( .A(A[116]), .B(n1144), .CI(
        C[116]), .CO(C[117]) );
  FA_13509 \FA_INST_0[0].FA_INST_1[117].FA_  ( .A(A[117]), .B(n1145), .CI(
        C[117]), .CO(C[118]) );
  FA_13508 \FA_INST_0[0].FA_INST_1[118].FA_  ( .A(A[118]), .B(n1146), .CI(
        C[118]), .CO(C[119]) );
  FA_13507 \FA_INST_0[0].FA_INST_1[119].FA_  ( .A(A[119]), .B(n1147), .CI(
        C[119]), .CO(C[120]) );
  FA_13506 \FA_INST_0[0].FA_INST_1[120].FA_  ( .A(A[120]), .B(n1148), .CI(
        C[120]), .CO(C[121]) );
  FA_13505 \FA_INST_0[0].FA_INST_1[121].FA_  ( .A(A[121]), .B(n1149), .CI(
        C[121]), .CO(C[122]) );
  FA_13504 \FA_INST_0[0].FA_INST_1[122].FA_  ( .A(A[122]), .B(n1150), .CI(
        C[122]), .CO(C[123]) );
  FA_13503 \FA_INST_0[0].FA_INST_1[123].FA_  ( .A(A[123]), .B(n1151), .CI(
        C[123]), .CO(C[124]) );
  FA_13502 \FA_INST_0[0].FA_INST_1[124].FA_  ( .A(A[124]), .B(n1152), .CI(
        C[124]), .CO(C[125]) );
  FA_13501 \FA_INST_0[0].FA_INST_1[125].FA_  ( .A(A[125]), .B(n1153), .CI(
        C[125]), .CO(C[126]) );
  FA_13500 \FA_INST_0[0].FA_INST_1[126].FA_  ( .A(A[126]), .B(n1154), .CI(
        C[126]), .CO(C[127]) );
  FA_13499 \FA_INST_0[0].FA_INST_1[127].FA_  ( .A(A[127]), .B(n1155), .CI(
        C[127]), .CO(C[128]) );
  FA_13498 \FA_INST_0[0].FA_INST_1[128].FA_  ( .A(A[128]), .B(n1156), .CI(
        C[128]), .CO(C[129]) );
  FA_13497 \FA_INST_0[0].FA_INST_1[129].FA_  ( .A(A[129]), .B(n1157), .CI(
        C[129]), .CO(C[130]) );
  FA_13496 \FA_INST_0[0].FA_INST_1[130].FA_  ( .A(A[130]), .B(n1158), .CI(
        C[130]), .CO(C[131]) );
  FA_13495 \FA_INST_0[0].FA_INST_1[131].FA_  ( .A(A[131]), .B(n1159), .CI(
        C[131]), .CO(C[132]) );
  FA_13494 \FA_INST_0[0].FA_INST_1[132].FA_  ( .A(A[132]), .B(n1160), .CI(
        C[132]), .CO(C[133]) );
  FA_13493 \FA_INST_0[0].FA_INST_1[133].FA_  ( .A(A[133]), .B(n1161), .CI(
        C[133]), .CO(C[134]) );
  FA_13492 \FA_INST_0[0].FA_INST_1[134].FA_  ( .A(A[134]), .B(n1162), .CI(
        C[134]), .CO(C[135]) );
  FA_13491 \FA_INST_0[0].FA_INST_1[135].FA_  ( .A(A[135]), .B(n1163), .CI(
        C[135]), .CO(C[136]) );
  FA_13490 \FA_INST_0[0].FA_INST_1[136].FA_  ( .A(A[136]), .B(n1164), .CI(
        C[136]), .CO(C[137]) );
  FA_13489 \FA_INST_0[0].FA_INST_1[137].FA_  ( .A(A[137]), .B(n1165), .CI(
        C[137]), .CO(C[138]) );
  FA_13488 \FA_INST_0[0].FA_INST_1[138].FA_  ( .A(A[138]), .B(n1166), .CI(
        C[138]), .CO(C[139]) );
  FA_13487 \FA_INST_0[0].FA_INST_1[139].FA_  ( .A(A[139]), .B(n1167), .CI(
        C[139]), .CO(C[140]) );
  FA_13486 \FA_INST_0[0].FA_INST_1[140].FA_  ( .A(A[140]), .B(n1168), .CI(
        C[140]), .CO(C[141]) );
  FA_13485 \FA_INST_0[0].FA_INST_1[141].FA_  ( .A(A[141]), .B(n1169), .CI(
        C[141]), .CO(C[142]) );
  FA_13484 \FA_INST_0[0].FA_INST_1[142].FA_  ( .A(A[142]), .B(n1170), .CI(
        C[142]), .CO(C[143]) );
  FA_13483 \FA_INST_0[0].FA_INST_1[143].FA_  ( .A(A[143]), .B(n1171), .CI(
        C[143]), .CO(C[144]) );
  FA_13482 \FA_INST_0[0].FA_INST_1[144].FA_  ( .A(A[144]), .B(n1172), .CI(
        C[144]), .CO(C[145]) );
  FA_13481 \FA_INST_0[0].FA_INST_1[145].FA_  ( .A(A[145]), .B(n1173), .CI(
        C[145]), .CO(C[146]) );
  FA_13480 \FA_INST_0[0].FA_INST_1[146].FA_  ( .A(A[146]), .B(n1174), .CI(
        C[146]), .CO(C[147]) );
  FA_13479 \FA_INST_0[0].FA_INST_1[147].FA_  ( .A(A[147]), .B(n1175), .CI(
        C[147]), .CO(C[148]) );
  FA_13478 \FA_INST_0[0].FA_INST_1[148].FA_  ( .A(A[148]), .B(n1176), .CI(
        C[148]), .CO(C[149]) );
  FA_13477 \FA_INST_0[0].FA_INST_1[149].FA_  ( .A(A[149]), .B(n1177), .CI(
        C[149]), .CO(C[150]) );
  FA_13476 \FA_INST_0[0].FA_INST_1[150].FA_  ( .A(A[150]), .B(n1178), .CI(
        C[150]), .CO(C[151]) );
  FA_13475 \FA_INST_0[0].FA_INST_1[151].FA_  ( .A(A[151]), .B(n1179), .CI(
        C[151]), .CO(C[152]) );
  FA_13474 \FA_INST_0[0].FA_INST_1[152].FA_  ( .A(A[152]), .B(n1180), .CI(
        C[152]), .CO(C[153]) );
  FA_13473 \FA_INST_0[0].FA_INST_1[153].FA_  ( .A(A[153]), .B(n1181), .CI(
        C[153]), .CO(C[154]) );
  FA_13472 \FA_INST_0[0].FA_INST_1[154].FA_  ( .A(A[154]), .B(n1182), .CI(
        C[154]), .CO(C[155]) );
  FA_13471 \FA_INST_0[0].FA_INST_1[155].FA_  ( .A(A[155]), .B(n1183), .CI(
        C[155]), .CO(C[156]) );
  FA_13470 \FA_INST_0[0].FA_INST_1[156].FA_  ( .A(A[156]), .B(n1184), .CI(
        C[156]), .CO(C[157]) );
  FA_13469 \FA_INST_0[0].FA_INST_1[157].FA_  ( .A(A[157]), .B(n1185), .CI(
        C[157]), .CO(C[158]) );
  FA_13468 \FA_INST_0[0].FA_INST_1[158].FA_  ( .A(A[158]), .B(n1186), .CI(
        C[158]), .CO(C[159]) );
  FA_13467 \FA_INST_0[0].FA_INST_1[159].FA_  ( .A(A[159]), .B(n1187), .CI(
        C[159]), .CO(C[160]) );
  FA_13466 \FA_INST_0[0].FA_INST_1[160].FA_  ( .A(A[160]), .B(n1188), .CI(
        C[160]), .CO(C[161]) );
  FA_13465 \FA_INST_0[0].FA_INST_1[161].FA_  ( .A(A[161]), .B(n1189), .CI(
        C[161]), .CO(C[162]) );
  FA_13464 \FA_INST_0[0].FA_INST_1[162].FA_  ( .A(A[162]), .B(n1190), .CI(
        C[162]), .CO(C[163]) );
  FA_13463 \FA_INST_0[0].FA_INST_1[163].FA_  ( .A(A[163]), .B(n1191), .CI(
        C[163]), .CO(C[164]) );
  FA_13462 \FA_INST_0[0].FA_INST_1[164].FA_  ( .A(A[164]), .B(n1192), .CI(
        C[164]), .CO(C[165]) );
  FA_13461 \FA_INST_0[0].FA_INST_1[165].FA_  ( .A(A[165]), .B(n1193), .CI(
        C[165]), .CO(C[166]) );
  FA_13460 \FA_INST_0[0].FA_INST_1[166].FA_  ( .A(A[166]), .B(n1194), .CI(
        C[166]), .CO(C[167]) );
  FA_13459 \FA_INST_0[0].FA_INST_1[167].FA_  ( .A(A[167]), .B(n1195), .CI(
        C[167]), .CO(C[168]) );
  FA_13458 \FA_INST_0[0].FA_INST_1[168].FA_  ( .A(A[168]), .B(n1196), .CI(
        C[168]), .CO(C[169]) );
  FA_13457 \FA_INST_0[0].FA_INST_1[169].FA_  ( .A(A[169]), .B(n1197), .CI(
        C[169]), .CO(C[170]) );
  FA_13456 \FA_INST_0[0].FA_INST_1[170].FA_  ( .A(A[170]), .B(n1198), .CI(
        C[170]), .CO(C[171]) );
  FA_13455 \FA_INST_0[0].FA_INST_1[171].FA_  ( .A(A[171]), .B(n1199), .CI(
        C[171]), .CO(C[172]) );
  FA_13454 \FA_INST_0[0].FA_INST_1[172].FA_  ( .A(A[172]), .B(n1200), .CI(
        C[172]), .CO(C[173]) );
  FA_13453 \FA_INST_0[0].FA_INST_1[173].FA_  ( .A(A[173]), .B(n1201), .CI(
        C[173]), .CO(C[174]) );
  FA_13452 \FA_INST_0[0].FA_INST_1[174].FA_  ( .A(A[174]), .B(n1202), .CI(
        C[174]), .CO(C[175]) );
  FA_13451 \FA_INST_0[0].FA_INST_1[175].FA_  ( .A(A[175]), .B(n1203), .CI(
        C[175]), .CO(C[176]) );
  FA_13450 \FA_INST_0[0].FA_INST_1[176].FA_  ( .A(A[176]), .B(n1204), .CI(
        C[176]), .CO(C[177]) );
  FA_13449 \FA_INST_0[0].FA_INST_1[177].FA_  ( .A(A[177]), .B(n1205), .CI(
        C[177]), .CO(C[178]) );
  FA_13448 \FA_INST_0[0].FA_INST_1[178].FA_  ( .A(A[178]), .B(n1206), .CI(
        C[178]), .CO(C[179]) );
  FA_13447 \FA_INST_0[0].FA_INST_1[179].FA_  ( .A(A[179]), .B(n1207), .CI(
        C[179]), .CO(C[180]) );
  FA_13446 \FA_INST_0[0].FA_INST_1[180].FA_  ( .A(A[180]), .B(n1208), .CI(
        C[180]), .CO(C[181]) );
  FA_13445 \FA_INST_0[0].FA_INST_1[181].FA_  ( .A(A[181]), .B(n1209), .CI(
        C[181]), .CO(C[182]) );
  FA_13444 \FA_INST_0[0].FA_INST_1[182].FA_  ( .A(A[182]), .B(n1210), .CI(
        C[182]), .CO(C[183]) );
  FA_13443 \FA_INST_0[0].FA_INST_1[183].FA_  ( .A(A[183]), .B(n1211), .CI(
        C[183]), .CO(C[184]) );
  FA_13442 \FA_INST_0[0].FA_INST_1[184].FA_  ( .A(A[184]), .B(n1212), .CI(
        C[184]), .CO(C[185]) );
  FA_13441 \FA_INST_0[0].FA_INST_1[185].FA_  ( .A(A[185]), .B(n1213), .CI(
        C[185]), .CO(C[186]) );
  FA_13440 \FA_INST_0[0].FA_INST_1[186].FA_  ( .A(A[186]), .B(n1214), .CI(
        C[186]), .CO(C[187]) );
  FA_13439 \FA_INST_0[0].FA_INST_1[187].FA_  ( .A(A[187]), .B(n1215), .CI(
        C[187]), .CO(C[188]) );
  FA_13438 \FA_INST_0[0].FA_INST_1[188].FA_  ( .A(A[188]), .B(n1216), .CI(
        C[188]), .CO(C[189]) );
  FA_13437 \FA_INST_0[0].FA_INST_1[189].FA_  ( .A(A[189]), .B(n1217), .CI(
        C[189]), .CO(C[190]) );
  FA_13436 \FA_INST_0[0].FA_INST_1[190].FA_  ( .A(A[190]), .B(n1218), .CI(
        C[190]), .CO(C[191]) );
  FA_13435 \FA_INST_0[0].FA_INST_1[191].FA_  ( .A(A[191]), .B(n1219), .CI(
        C[191]), .CO(C[192]) );
  FA_13434 \FA_INST_0[0].FA_INST_1[192].FA_  ( .A(A[192]), .B(n1220), .CI(
        C[192]), .CO(C[193]) );
  FA_13433 \FA_INST_0[0].FA_INST_1[193].FA_  ( .A(A[193]), .B(n1221), .CI(
        C[193]), .CO(C[194]) );
  FA_13432 \FA_INST_0[0].FA_INST_1[194].FA_  ( .A(A[194]), .B(n1222), .CI(
        C[194]), .CO(C[195]) );
  FA_13431 \FA_INST_0[0].FA_INST_1[195].FA_  ( .A(A[195]), .B(n1223), .CI(
        C[195]), .CO(C[196]) );
  FA_13430 \FA_INST_0[0].FA_INST_1[196].FA_  ( .A(A[196]), .B(n1224), .CI(
        C[196]), .CO(C[197]) );
  FA_13429 \FA_INST_0[0].FA_INST_1[197].FA_  ( .A(A[197]), .B(n1225), .CI(
        C[197]), .CO(C[198]) );
  FA_13428 \FA_INST_0[0].FA_INST_1[198].FA_  ( .A(A[198]), .B(n1226), .CI(
        C[198]), .CO(C[199]) );
  FA_13427 \FA_INST_0[0].FA_INST_1[199].FA_  ( .A(A[199]), .B(n1227), .CI(
        C[199]), .CO(C[200]) );
  FA_13426 \FA_INST_0[0].FA_INST_1[200].FA_  ( .A(A[200]), .B(n1228), .CI(
        C[200]), .CO(C[201]) );
  FA_13425 \FA_INST_0[0].FA_INST_1[201].FA_  ( .A(A[201]), .B(n1229), .CI(
        C[201]), .CO(C[202]) );
  FA_13424 \FA_INST_0[0].FA_INST_1[202].FA_  ( .A(A[202]), .B(n1230), .CI(
        C[202]), .CO(C[203]) );
  FA_13423 \FA_INST_0[0].FA_INST_1[203].FA_  ( .A(A[203]), .B(n1231), .CI(
        C[203]), .CO(C[204]) );
  FA_13422 \FA_INST_0[0].FA_INST_1[204].FA_  ( .A(A[204]), .B(n1232), .CI(
        C[204]), .CO(C[205]) );
  FA_13421 \FA_INST_0[0].FA_INST_1[205].FA_  ( .A(A[205]), .B(n1233), .CI(
        C[205]), .CO(C[206]) );
  FA_13420 \FA_INST_0[0].FA_INST_1[206].FA_  ( .A(A[206]), .B(n1234), .CI(
        C[206]), .CO(C[207]) );
  FA_13419 \FA_INST_0[0].FA_INST_1[207].FA_  ( .A(A[207]), .B(n1235), .CI(
        C[207]), .CO(C[208]) );
  FA_13418 \FA_INST_0[0].FA_INST_1[208].FA_  ( .A(A[208]), .B(n1236), .CI(
        C[208]), .CO(C[209]) );
  FA_13417 \FA_INST_0[0].FA_INST_1[209].FA_  ( .A(A[209]), .B(n1237), .CI(
        C[209]), .CO(C[210]) );
  FA_13416 \FA_INST_0[0].FA_INST_1[210].FA_  ( .A(A[210]), .B(n1238), .CI(
        C[210]), .CO(C[211]) );
  FA_13415 \FA_INST_0[0].FA_INST_1[211].FA_  ( .A(A[211]), .B(n1239), .CI(
        C[211]), .CO(C[212]) );
  FA_13414 \FA_INST_0[0].FA_INST_1[212].FA_  ( .A(A[212]), .B(n1240), .CI(
        C[212]), .CO(C[213]) );
  FA_13413 \FA_INST_0[0].FA_INST_1[213].FA_  ( .A(A[213]), .B(n1241), .CI(
        C[213]), .CO(C[214]) );
  FA_13412 \FA_INST_0[0].FA_INST_1[214].FA_  ( .A(A[214]), .B(n1242), .CI(
        C[214]), .CO(C[215]) );
  FA_13411 \FA_INST_0[0].FA_INST_1[215].FA_  ( .A(A[215]), .B(n1243), .CI(
        C[215]), .CO(C[216]) );
  FA_13410 \FA_INST_0[0].FA_INST_1[216].FA_  ( .A(A[216]), .B(n1244), .CI(
        C[216]), .CO(C[217]) );
  FA_13409 \FA_INST_0[0].FA_INST_1[217].FA_  ( .A(A[217]), .B(n1245), .CI(
        C[217]), .CO(C[218]) );
  FA_13408 \FA_INST_0[0].FA_INST_1[218].FA_  ( .A(A[218]), .B(n1246), .CI(
        C[218]), .CO(C[219]) );
  FA_13407 \FA_INST_0[0].FA_INST_1[219].FA_  ( .A(A[219]), .B(n1247), .CI(
        C[219]), .CO(C[220]) );
  FA_13406 \FA_INST_0[0].FA_INST_1[220].FA_  ( .A(A[220]), .B(n1248), .CI(
        C[220]), .CO(C[221]) );
  FA_13405 \FA_INST_0[0].FA_INST_1[221].FA_  ( .A(A[221]), .B(n1249), .CI(
        C[221]), .CO(C[222]) );
  FA_13404 \FA_INST_0[0].FA_INST_1[222].FA_  ( .A(A[222]), .B(n1250), .CI(
        C[222]), .CO(C[223]) );
  FA_13403 \FA_INST_0[0].FA_INST_1[223].FA_  ( .A(A[223]), .B(n1251), .CI(
        C[223]), .CO(C[224]) );
  FA_13402 \FA_INST_0[0].FA_INST_1[224].FA_  ( .A(A[224]), .B(n1252), .CI(
        C[224]), .CO(C[225]) );
  FA_13401 \FA_INST_0[0].FA_INST_1[225].FA_  ( .A(A[225]), .B(n1253), .CI(
        C[225]), .CO(C[226]) );
  FA_13400 \FA_INST_0[0].FA_INST_1[226].FA_  ( .A(A[226]), .B(n1254), .CI(
        C[226]), .CO(C[227]) );
  FA_13399 \FA_INST_0[0].FA_INST_1[227].FA_  ( .A(A[227]), .B(n1255), .CI(
        C[227]), .CO(C[228]) );
  FA_13398 \FA_INST_0[0].FA_INST_1[228].FA_  ( .A(A[228]), .B(n1256), .CI(
        C[228]), .CO(C[229]) );
  FA_13397 \FA_INST_0[0].FA_INST_1[229].FA_  ( .A(A[229]), .B(n1257), .CI(
        C[229]), .CO(C[230]) );
  FA_13396 \FA_INST_0[0].FA_INST_1[230].FA_  ( .A(A[230]), .B(n1258), .CI(
        C[230]), .CO(C[231]) );
  FA_13395 \FA_INST_0[0].FA_INST_1[231].FA_  ( .A(A[231]), .B(n1259), .CI(
        C[231]), .CO(C[232]) );
  FA_13394 \FA_INST_0[0].FA_INST_1[232].FA_  ( .A(A[232]), .B(n1260), .CI(
        C[232]), .CO(C[233]) );
  FA_13393 \FA_INST_0[0].FA_INST_1[233].FA_  ( .A(A[233]), .B(n1261), .CI(
        C[233]), .CO(C[234]) );
  FA_13392 \FA_INST_0[0].FA_INST_1[234].FA_  ( .A(A[234]), .B(n1262), .CI(
        C[234]), .CO(C[235]) );
  FA_13391 \FA_INST_0[0].FA_INST_1[235].FA_  ( .A(A[235]), .B(n1263), .CI(
        C[235]), .CO(C[236]) );
  FA_13390 \FA_INST_0[0].FA_INST_1[236].FA_  ( .A(A[236]), .B(n1264), .CI(
        C[236]), .CO(C[237]) );
  FA_13389 \FA_INST_0[0].FA_INST_1[237].FA_  ( .A(A[237]), .B(n1265), .CI(
        C[237]), .CO(C[238]) );
  FA_13388 \FA_INST_0[0].FA_INST_1[238].FA_  ( .A(A[238]), .B(n1266), .CI(
        C[238]), .CO(C[239]) );
  FA_13387 \FA_INST_0[0].FA_INST_1[239].FA_  ( .A(A[239]), .B(n1267), .CI(
        C[239]), .CO(C[240]) );
  FA_13386 \FA_INST_0[0].FA_INST_1[240].FA_  ( .A(A[240]), .B(n1268), .CI(
        C[240]), .CO(C[241]) );
  FA_13385 \FA_INST_0[0].FA_INST_1[241].FA_  ( .A(A[241]), .B(n1269), .CI(
        C[241]), .CO(C[242]) );
  FA_13384 \FA_INST_0[0].FA_INST_1[242].FA_  ( .A(A[242]), .B(n1270), .CI(
        C[242]), .CO(C[243]) );
  FA_13383 \FA_INST_0[0].FA_INST_1[243].FA_  ( .A(A[243]), .B(n1271), .CI(
        C[243]), .CO(C[244]) );
  FA_13382 \FA_INST_0[0].FA_INST_1[244].FA_  ( .A(A[244]), .B(n1272), .CI(
        C[244]), .CO(C[245]) );
  FA_13381 \FA_INST_0[0].FA_INST_1[245].FA_  ( .A(A[245]), .B(n1273), .CI(
        C[245]), .CO(C[246]) );
  FA_13380 \FA_INST_0[0].FA_INST_1[246].FA_  ( .A(A[246]), .B(n1274), .CI(
        C[246]), .CO(C[247]) );
  FA_13379 \FA_INST_0[0].FA_INST_1[247].FA_  ( .A(A[247]), .B(n1275), .CI(
        C[247]), .CO(C[248]) );
  FA_13378 \FA_INST_0[0].FA_INST_1[248].FA_  ( .A(A[248]), .B(n1276), .CI(
        C[248]), .CO(C[249]) );
  FA_13377 \FA_INST_0[0].FA_INST_1[249].FA_  ( .A(A[249]), .B(n1277), .CI(
        C[249]), .CO(C[250]) );
  FA_13376 \FA_INST_0[0].FA_INST_1[250].FA_  ( .A(A[250]), .B(n1278), .CI(
        C[250]), .CO(C[251]) );
  FA_13375 \FA_INST_0[0].FA_INST_1[251].FA_  ( .A(A[251]), .B(n1279), .CI(
        C[251]), .CO(C[252]) );
  FA_13374 \FA_INST_0[0].FA_INST_1[252].FA_  ( .A(A[252]), .B(n1280), .CI(
        C[252]), .CO(C[253]) );
  FA_13373 \FA_INST_0[0].FA_INST_1[253].FA_  ( .A(A[253]), .B(n1281), .CI(
        C[253]), .CO(C[254]) );
  FA_13372 \FA_INST_0[0].FA_INST_1[254].FA_  ( .A(A[254]), .B(n1282), .CI(
        C[254]), .CO(C[255]) );
  FA_13371 \FA_INST_0[0].FA_INST_1[255].FA_  ( .A(A[255]), .B(n1283), .CI(
        C[255]), .CO(C[256]) );
  FA_13370 \FA_INST_0[0].FA_INST_1[256].FA_  ( .A(A[256]), .B(n1284), .CI(
        C[256]), .CO(C[257]) );
  FA_13369 \FA_INST_0[0].FA_INST_1[257].FA_  ( .A(A[257]), .B(n1285), .CI(
        C[257]), .CO(C[258]) );
  FA_13368 \FA_INST_0[0].FA_INST_1[258].FA_  ( .A(A[258]), .B(n1286), .CI(
        C[258]), .CO(C[259]) );
  FA_13367 \FA_INST_0[0].FA_INST_1[259].FA_  ( .A(A[259]), .B(n1287), .CI(
        C[259]), .CO(C[260]) );
  FA_13366 \FA_INST_0[0].FA_INST_1[260].FA_  ( .A(A[260]), .B(n1288), .CI(
        C[260]), .CO(C[261]) );
  FA_13365 \FA_INST_0[0].FA_INST_1[261].FA_  ( .A(A[261]), .B(n1289), .CI(
        C[261]), .CO(C[262]) );
  FA_13364 \FA_INST_0[0].FA_INST_1[262].FA_  ( .A(A[262]), .B(n1290), .CI(
        C[262]), .CO(C[263]) );
  FA_13363 \FA_INST_0[0].FA_INST_1[263].FA_  ( .A(A[263]), .B(n1291), .CI(
        C[263]), .CO(C[264]) );
  FA_13362 \FA_INST_0[0].FA_INST_1[264].FA_  ( .A(A[264]), .B(n1292), .CI(
        C[264]), .CO(C[265]) );
  FA_13361 \FA_INST_0[0].FA_INST_1[265].FA_  ( .A(A[265]), .B(n1293), .CI(
        C[265]), .CO(C[266]) );
  FA_13360 \FA_INST_0[0].FA_INST_1[266].FA_  ( .A(A[266]), .B(n1294), .CI(
        C[266]), .CO(C[267]) );
  FA_13359 \FA_INST_0[0].FA_INST_1[267].FA_  ( .A(A[267]), .B(n1295), .CI(
        C[267]), .CO(C[268]) );
  FA_13358 \FA_INST_0[0].FA_INST_1[268].FA_  ( .A(A[268]), .B(n1296), .CI(
        C[268]), .CO(C[269]) );
  FA_13357 \FA_INST_0[0].FA_INST_1[269].FA_  ( .A(A[269]), .B(n1297), .CI(
        C[269]), .CO(C[270]) );
  FA_13356 \FA_INST_0[0].FA_INST_1[270].FA_  ( .A(A[270]), .B(n1298), .CI(
        C[270]), .CO(C[271]) );
  FA_13355 \FA_INST_0[0].FA_INST_1[271].FA_  ( .A(A[271]), .B(n1299), .CI(
        C[271]), .CO(C[272]) );
  FA_13354 \FA_INST_0[0].FA_INST_1[272].FA_  ( .A(A[272]), .B(n1300), .CI(
        C[272]), .CO(C[273]) );
  FA_13353 \FA_INST_0[0].FA_INST_1[273].FA_  ( .A(A[273]), .B(n1301), .CI(
        C[273]), .CO(C[274]) );
  FA_13352 \FA_INST_0[0].FA_INST_1[274].FA_  ( .A(A[274]), .B(n1302), .CI(
        C[274]), .CO(C[275]) );
  FA_13351 \FA_INST_0[0].FA_INST_1[275].FA_  ( .A(A[275]), .B(n1303), .CI(
        C[275]), .CO(C[276]) );
  FA_13350 \FA_INST_0[0].FA_INST_1[276].FA_  ( .A(A[276]), .B(n1304), .CI(
        C[276]), .CO(C[277]) );
  FA_13349 \FA_INST_0[0].FA_INST_1[277].FA_  ( .A(A[277]), .B(n1305), .CI(
        C[277]), .CO(C[278]) );
  FA_13348 \FA_INST_0[0].FA_INST_1[278].FA_  ( .A(A[278]), .B(n1306), .CI(
        C[278]), .CO(C[279]) );
  FA_13347 \FA_INST_0[0].FA_INST_1[279].FA_  ( .A(A[279]), .B(n1307), .CI(
        C[279]), .CO(C[280]) );
  FA_13346 \FA_INST_0[0].FA_INST_1[280].FA_  ( .A(A[280]), .B(n1308), .CI(
        C[280]), .CO(C[281]) );
  FA_13345 \FA_INST_0[0].FA_INST_1[281].FA_  ( .A(A[281]), .B(n1309), .CI(
        C[281]), .CO(C[282]) );
  FA_13344 \FA_INST_0[0].FA_INST_1[282].FA_  ( .A(A[282]), .B(n1310), .CI(
        C[282]), .CO(C[283]) );
  FA_13343 \FA_INST_0[0].FA_INST_1[283].FA_  ( .A(A[283]), .B(n1311), .CI(
        C[283]), .CO(C[284]) );
  FA_13342 \FA_INST_0[0].FA_INST_1[284].FA_  ( .A(A[284]), .B(n1312), .CI(
        C[284]), .CO(C[285]) );
  FA_13341 \FA_INST_0[0].FA_INST_1[285].FA_  ( .A(A[285]), .B(n1313), .CI(
        C[285]), .CO(C[286]) );
  FA_13340 \FA_INST_0[0].FA_INST_1[286].FA_  ( .A(A[286]), .B(n1314), .CI(
        C[286]), .CO(C[287]) );
  FA_13339 \FA_INST_0[0].FA_INST_1[287].FA_  ( .A(A[287]), .B(n1315), .CI(
        C[287]), .CO(C[288]) );
  FA_13338 \FA_INST_0[0].FA_INST_1[288].FA_  ( .A(A[288]), .B(n1316), .CI(
        C[288]), .CO(C[289]) );
  FA_13337 \FA_INST_0[0].FA_INST_1[289].FA_  ( .A(A[289]), .B(n1317), .CI(
        C[289]), .CO(C[290]) );
  FA_13336 \FA_INST_0[0].FA_INST_1[290].FA_  ( .A(A[290]), .B(n1318), .CI(
        C[290]), .CO(C[291]) );
  FA_13335 \FA_INST_0[0].FA_INST_1[291].FA_  ( .A(A[291]), .B(n1319), .CI(
        C[291]), .CO(C[292]) );
  FA_13334 \FA_INST_0[0].FA_INST_1[292].FA_  ( .A(A[292]), .B(n1320), .CI(
        C[292]), .CO(C[293]) );
  FA_13333 \FA_INST_0[0].FA_INST_1[293].FA_  ( .A(A[293]), .B(n1321), .CI(
        C[293]), .CO(C[294]) );
  FA_13332 \FA_INST_0[0].FA_INST_1[294].FA_  ( .A(A[294]), .B(n1322), .CI(
        C[294]), .CO(C[295]) );
  FA_13331 \FA_INST_0[0].FA_INST_1[295].FA_  ( .A(A[295]), .B(n1323), .CI(
        C[295]), .CO(C[296]) );
  FA_13330 \FA_INST_0[0].FA_INST_1[296].FA_  ( .A(A[296]), .B(n1324), .CI(
        C[296]), .CO(C[297]) );
  FA_13329 \FA_INST_0[0].FA_INST_1[297].FA_  ( .A(A[297]), .B(n1325), .CI(
        C[297]), .CO(C[298]) );
  FA_13328 \FA_INST_0[0].FA_INST_1[298].FA_  ( .A(A[298]), .B(n1326), .CI(
        C[298]), .CO(C[299]) );
  FA_13327 \FA_INST_0[0].FA_INST_1[299].FA_  ( .A(A[299]), .B(n1327), .CI(
        C[299]), .CO(C[300]) );
  FA_13326 \FA_INST_0[0].FA_INST_1[300].FA_  ( .A(A[300]), .B(n1328), .CI(
        C[300]), .CO(C[301]) );
  FA_13325 \FA_INST_0[0].FA_INST_1[301].FA_  ( .A(A[301]), .B(n1329), .CI(
        C[301]), .CO(C[302]) );
  FA_13324 \FA_INST_0[0].FA_INST_1[302].FA_  ( .A(A[302]), .B(n1330), .CI(
        C[302]), .CO(C[303]) );
  FA_13323 \FA_INST_0[0].FA_INST_1[303].FA_  ( .A(A[303]), .B(n1331), .CI(
        C[303]), .CO(C[304]) );
  FA_13322 \FA_INST_0[0].FA_INST_1[304].FA_  ( .A(A[304]), .B(n1332), .CI(
        C[304]), .CO(C[305]) );
  FA_13321 \FA_INST_0[0].FA_INST_1[305].FA_  ( .A(A[305]), .B(n1333), .CI(
        C[305]), .CO(C[306]) );
  FA_13320 \FA_INST_0[0].FA_INST_1[306].FA_  ( .A(A[306]), .B(n1334), .CI(
        C[306]), .CO(C[307]) );
  FA_13319 \FA_INST_0[0].FA_INST_1[307].FA_  ( .A(A[307]), .B(n1335), .CI(
        C[307]), .CO(C[308]) );
  FA_13318 \FA_INST_0[0].FA_INST_1[308].FA_  ( .A(A[308]), .B(n1336), .CI(
        C[308]), .CO(C[309]) );
  FA_13317 \FA_INST_0[0].FA_INST_1[309].FA_  ( .A(A[309]), .B(n1337), .CI(
        C[309]), .CO(C[310]) );
  FA_13316 \FA_INST_0[0].FA_INST_1[310].FA_  ( .A(A[310]), .B(n1338), .CI(
        C[310]), .CO(C[311]) );
  FA_13315 \FA_INST_0[0].FA_INST_1[311].FA_  ( .A(A[311]), .B(n1339), .CI(
        C[311]), .CO(C[312]) );
  FA_13314 \FA_INST_0[0].FA_INST_1[312].FA_  ( .A(A[312]), .B(n1340), .CI(
        C[312]), .CO(C[313]) );
  FA_13313 \FA_INST_0[0].FA_INST_1[313].FA_  ( .A(A[313]), .B(n1341), .CI(
        C[313]), .CO(C[314]) );
  FA_13312 \FA_INST_0[0].FA_INST_1[314].FA_  ( .A(A[314]), .B(n1342), .CI(
        C[314]), .CO(C[315]) );
  FA_13311 \FA_INST_0[0].FA_INST_1[315].FA_  ( .A(A[315]), .B(n1343), .CI(
        C[315]), .CO(C[316]) );
  FA_13310 \FA_INST_0[0].FA_INST_1[316].FA_  ( .A(A[316]), .B(n1344), .CI(
        C[316]), .CO(C[317]) );
  FA_13309 \FA_INST_0[0].FA_INST_1[317].FA_  ( .A(A[317]), .B(n1345), .CI(
        C[317]), .CO(C[318]) );
  FA_13308 \FA_INST_0[0].FA_INST_1[318].FA_  ( .A(A[318]), .B(n1346), .CI(
        C[318]), .CO(C[319]) );
  FA_13307 \FA_INST_0[0].FA_INST_1[319].FA_  ( .A(A[319]), .B(n1347), .CI(
        C[319]), .CO(C[320]) );
  FA_13306 \FA_INST_0[0].FA_INST_1[320].FA_  ( .A(A[320]), .B(n1348), .CI(
        C[320]), .CO(C[321]) );
  FA_13305 \FA_INST_0[0].FA_INST_1[321].FA_  ( .A(A[321]), .B(n1349), .CI(
        C[321]), .CO(C[322]) );
  FA_13304 \FA_INST_0[0].FA_INST_1[322].FA_  ( .A(A[322]), .B(n1350), .CI(
        C[322]), .CO(C[323]) );
  FA_13303 \FA_INST_0[0].FA_INST_1[323].FA_  ( .A(A[323]), .B(n1351), .CI(
        C[323]), .CO(C[324]) );
  FA_13302 \FA_INST_0[0].FA_INST_1[324].FA_  ( .A(A[324]), .B(n1352), .CI(
        C[324]), .CO(C[325]) );
  FA_13301 \FA_INST_0[0].FA_INST_1[325].FA_  ( .A(A[325]), .B(n1353), .CI(
        C[325]), .CO(C[326]) );
  FA_13300 \FA_INST_0[0].FA_INST_1[326].FA_  ( .A(A[326]), .B(n1354), .CI(
        C[326]), .CO(C[327]) );
  FA_13299 \FA_INST_0[0].FA_INST_1[327].FA_  ( .A(A[327]), .B(n1355), .CI(
        C[327]), .CO(C[328]) );
  FA_13298 \FA_INST_0[0].FA_INST_1[328].FA_  ( .A(A[328]), .B(n1356), .CI(
        C[328]), .CO(C[329]) );
  FA_13297 \FA_INST_0[0].FA_INST_1[329].FA_  ( .A(A[329]), .B(n1357), .CI(
        C[329]), .CO(C[330]) );
  FA_13296 \FA_INST_0[0].FA_INST_1[330].FA_  ( .A(A[330]), .B(n1358), .CI(
        C[330]), .CO(C[331]) );
  FA_13295 \FA_INST_0[0].FA_INST_1[331].FA_  ( .A(A[331]), .B(n1359), .CI(
        C[331]), .CO(C[332]) );
  FA_13294 \FA_INST_0[0].FA_INST_1[332].FA_  ( .A(A[332]), .B(n1360), .CI(
        C[332]), .CO(C[333]) );
  FA_13293 \FA_INST_0[0].FA_INST_1[333].FA_  ( .A(A[333]), .B(n1361), .CI(
        C[333]), .CO(C[334]) );
  FA_13292 \FA_INST_0[0].FA_INST_1[334].FA_  ( .A(A[334]), .B(n1362), .CI(
        C[334]), .CO(C[335]) );
  FA_13291 \FA_INST_0[0].FA_INST_1[335].FA_  ( .A(A[335]), .B(n1363), .CI(
        C[335]), .CO(C[336]) );
  FA_13290 \FA_INST_0[0].FA_INST_1[336].FA_  ( .A(A[336]), .B(n1364), .CI(
        C[336]), .CO(C[337]) );
  FA_13289 \FA_INST_0[0].FA_INST_1[337].FA_  ( .A(A[337]), .B(n1365), .CI(
        C[337]), .CO(C[338]) );
  FA_13288 \FA_INST_0[0].FA_INST_1[338].FA_  ( .A(A[338]), .B(n1366), .CI(
        C[338]), .CO(C[339]) );
  FA_13287 \FA_INST_0[0].FA_INST_1[339].FA_  ( .A(A[339]), .B(n1367), .CI(
        C[339]), .CO(C[340]) );
  FA_13286 \FA_INST_0[0].FA_INST_1[340].FA_  ( .A(A[340]), .B(n1368), .CI(
        C[340]), .CO(C[341]) );
  FA_13285 \FA_INST_0[0].FA_INST_1[341].FA_  ( .A(A[341]), .B(n1369), .CI(
        C[341]), .CO(C[342]) );
  FA_13284 \FA_INST_0[0].FA_INST_1[342].FA_  ( .A(A[342]), .B(n1370), .CI(
        C[342]), .CO(C[343]) );
  FA_13283 \FA_INST_0[0].FA_INST_1[343].FA_  ( .A(A[343]), .B(n1371), .CI(
        C[343]), .CO(C[344]) );
  FA_13282 \FA_INST_0[0].FA_INST_1[344].FA_  ( .A(A[344]), .B(n1372), .CI(
        C[344]), .CO(C[345]) );
  FA_13281 \FA_INST_0[0].FA_INST_1[345].FA_  ( .A(A[345]), .B(n1373), .CI(
        C[345]), .CO(C[346]) );
  FA_13280 \FA_INST_0[0].FA_INST_1[346].FA_  ( .A(A[346]), .B(n1374), .CI(
        C[346]), .CO(C[347]) );
  FA_13279 \FA_INST_0[0].FA_INST_1[347].FA_  ( .A(A[347]), .B(n1375), .CI(
        C[347]), .CO(C[348]) );
  FA_13278 \FA_INST_0[0].FA_INST_1[348].FA_  ( .A(A[348]), .B(n1376), .CI(
        C[348]), .CO(C[349]) );
  FA_13277 \FA_INST_0[0].FA_INST_1[349].FA_  ( .A(A[349]), .B(n1377), .CI(
        C[349]), .CO(C[350]) );
  FA_13276 \FA_INST_0[0].FA_INST_1[350].FA_  ( .A(A[350]), .B(n1378), .CI(
        C[350]), .CO(C[351]) );
  FA_13275 \FA_INST_0[0].FA_INST_1[351].FA_  ( .A(A[351]), .B(n1379), .CI(
        C[351]), .CO(C[352]) );
  FA_13274 \FA_INST_0[0].FA_INST_1[352].FA_  ( .A(A[352]), .B(n1380), .CI(
        C[352]), .CO(C[353]) );
  FA_13273 \FA_INST_0[0].FA_INST_1[353].FA_  ( .A(A[353]), .B(n1381), .CI(
        C[353]), .CO(C[354]) );
  FA_13272 \FA_INST_0[0].FA_INST_1[354].FA_  ( .A(A[354]), .B(n1382), .CI(
        C[354]), .CO(C[355]) );
  FA_13271 \FA_INST_0[0].FA_INST_1[355].FA_  ( .A(A[355]), .B(n1383), .CI(
        C[355]), .CO(C[356]) );
  FA_13270 \FA_INST_0[0].FA_INST_1[356].FA_  ( .A(A[356]), .B(n1384), .CI(
        C[356]), .CO(C[357]) );
  FA_13269 \FA_INST_0[0].FA_INST_1[357].FA_  ( .A(A[357]), .B(n1385), .CI(
        C[357]), .CO(C[358]) );
  FA_13268 \FA_INST_0[0].FA_INST_1[358].FA_  ( .A(A[358]), .B(n1386), .CI(
        C[358]), .CO(C[359]) );
  FA_13267 \FA_INST_0[0].FA_INST_1[359].FA_  ( .A(A[359]), .B(n1387), .CI(
        C[359]), .CO(C[360]) );
  FA_13266 \FA_INST_0[0].FA_INST_1[360].FA_  ( .A(A[360]), .B(n1388), .CI(
        C[360]), .CO(C[361]) );
  FA_13265 \FA_INST_0[0].FA_INST_1[361].FA_  ( .A(A[361]), .B(n1389), .CI(
        C[361]), .CO(C[362]) );
  FA_13264 \FA_INST_0[0].FA_INST_1[362].FA_  ( .A(A[362]), .B(n1390), .CI(
        C[362]), .CO(C[363]) );
  FA_13263 \FA_INST_0[0].FA_INST_1[363].FA_  ( .A(A[363]), .B(n1391), .CI(
        C[363]), .CO(C[364]) );
  FA_13262 \FA_INST_0[0].FA_INST_1[364].FA_  ( .A(A[364]), .B(n1392), .CI(
        C[364]), .CO(C[365]) );
  FA_13261 \FA_INST_0[0].FA_INST_1[365].FA_  ( .A(A[365]), .B(n1393), .CI(
        C[365]), .CO(C[366]) );
  FA_13260 \FA_INST_0[0].FA_INST_1[366].FA_  ( .A(A[366]), .B(n1394), .CI(
        C[366]), .CO(C[367]) );
  FA_13259 \FA_INST_0[0].FA_INST_1[367].FA_  ( .A(A[367]), .B(n1395), .CI(
        C[367]), .CO(C[368]) );
  FA_13258 \FA_INST_0[0].FA_INST_1[368].FA_  ( .A(A[368]), .B(n1396), .CI(
        C[368]), .CO(C[369]) );
  FA_13257 \FA_INST_0[0].FA_INST_1[369].FA_  ( .A(A[369]), .B(n1397), .CI(
        C[369]), .CO(C[370]) );
  FA_13256 \FA_INST_0[0].FA_INST_1[370].FA_  ( .A(A[370]), .B(n1398), .CI(
        C[370]), .CO(C[371]) );
  FA_13255 \FA_INST_0[0].FA_INST_1[371].FA_  ( .A(A[371]), .B(n1399), .CI(
        C[371]), .CO(C[372]) );
  FA_13254 \FA_INST_0[0].FA_INST_1[372].FA_  ( .A(A[372]), .B(n1400), .CI(
        C[372]), .CO(C[373]) );
  FA_13253 \FA_INST_0[0].FA_INST_1[373].FA_  ( .A(A[373]), .B(n1401), .CI(
        C[373]), .CO(C[374]) );
  FA_13252 \FA_INST_0[0].FA_INST_1[374].FA_  ( .A(A[374]), .B(n1402), .CI(
        C[374]), .CO(C[375]) );
  FA_13251 \FA_INST_0[0].FA_INST_1[375].FA_  ( .A(A[375]), .B(n1403), .CI(
        C[375]), .CO(C[376]) );
  FA_13250 \FA_INST_0[0].FA_INST_1[376].FA_  ( .A(A[376]), .B(n1404), .CI(
        C[376]), .CO(C[377]) );
  FA_13249 \FA_INST_0[0].FA_INST_1[377].FA_  ( .A(A[377]), .B(n1405), .CI(
        C[377]), .CO(C[378]) );
  FA_13248 \FA_INST_0[0].FA_INST_1[378].FA_  ( .A(A[378]), .B(n1406), .CI(
        C[378]), .CO(C[379]) );
  FA_13247 \FA_INST_0[0].FA_INST_1[379].FA_  ( .A(A[379]), .B(n1407), .CI(
        C[379]), .CO(C[380]) );
  FA_13246 \FA_INST_0[0].FA_INST_1[380].FA_  ( .A(A[380]), .B(n1408), .CI(
        C[380]), .CO(C[381]) );
  FA_13245 \FA_INST_0[0].FA_INST_1[381].FA_  ( .A(A[381]), .B(n1409), .CI(
        C[381]), .CO(C[382]) );
  FA_13244 \FA_INST_0[0].FA_INST_1[382].FA_  ( .A(A[382]), .B(n1410), .CI(
        C[382]), .CO(C[383]) );
  FA_13243 \FA_INST_0[0].FA_INST_1[383].FA_  ( .A(A[383]), .B(n1411), .CI(
        C[383]), .CO(C[384]) );
  FA_13242 \FA_INST_0[0].FA_INST_1[384].FA_  ( .A(A[384]), .B(n1412), .CI(
        C[384]), .CO(C[385]) );
  FA_13241 \FA_INST_0[0].FA_INST_1[385].FA_  ( .A(A[385]), .B(n1413), .CI(
        C[385]), .CO(C[386]) );
  FA_13240 \FA_INST_0[0].FA_INST_1[386].FA_  ( .A(A[386]), .B(n1414), .CI(
        C[386]), .CO(C[387]) );
  FA_13239 \FA_INST_0[0].FA_INST_1[387].FA_  ( .A(A[387]), .B(n1415), .CI(
        C[387]), .CO(C[388]) );
  FA_13238 \FA_INST_0[0].FA_INST_1[388].FA_  ( .A(A[388]), .B(n1416), .CI(
        C[388]), .CO(C[389]) );
  FA_13237 \FA_INST_0[0].FA_INST_1[389].FA_  ( .A(A[389]), .B(n1417), .CI(
        C[389]), .CO(C[390]) );
  FA_13236 \FA_INST_0[0].FA_INST_1[390].FA_  ( .A(A[390]), .B(n1418), .CI(
        C[390]), .CO(C[391]) );
  FA_13235 \FA_INST_0[0].FA_INST_1[391].FA_  ( .A(A[391]), .B(n1419), .CI(
        C[391]), .CO(C[392]) );
  FA_13234 \FA_INST_0[0].FA_INST_1[392].FA_  ( .A(A[392]), .B(n1420), .CI(
        C[392]), .CO(C[393]) );
  FA_13233 \FA_INST_0[0].FA_INST_1[393].FA_  ( .A(A[393]), .B(n1421), .CI(
        C[393]), .CO(C[394]) );
  FA_13232 \FA_INST_0[0].FA_INST_1[394].FA_  ( .A(A[394]), .B(n1422), .CI(
        C[394]), .CO(C[395]) );
  FA_13231 \FA_INST_0[0].FA_INST_1[395].FA_  ( .A(A[395]), .B(n1423), .CI(
        C[395]), .CO(C[396]) );
  FA_13230 \FA_INST_0[0].FA_INST_1[396].FA_  ( .A(A[396]), .B(n1424), .CI(
        C[396]), .CO(C[397]) );
  FA_13229 \FA_INST_0[0].FA_INST_1[397].FA_  ( .A(A[397]), .B(n1425), .CI(
        C[397]), .CO(C[398]) );
  FA_13228 \FA_INST_0[0].FA_INST_1[398].FA_  ( .A(A[398]), .B(n1426), .CI(
        C[398]), .CO(C[399]) );
  FA_13227 \FA_INST_0[0].FA_INST_1[399].FA_  ( .A(A[399]), .B(n1427), .CI(
        C[399]), .CO(C[400]) );
  FA_13226 \FA_INST_0[0].FA_INST_1[400].FA_  ( .A(A[400]), .B(n1428), .CI(
        C[400]), .CO(C[401]) );
  FA_13225 \FA_INST_0[0].FA_INST_1[401].FA_  ( .A(A[401]), .B(n1429), .CI(
        C[401]), .CO(C[402]) );
  FA_13224 \FA_INST_0[0].FA_INST_1[402].FA_  ( .A(A[402]), .B(n1430), .CI(
        C[402]), .CO(C[403]) );
  FA_13223 \FA_INST_0[0].FA_INST_1[403].FA_  ( .A(A[403]), .B(n1431), .CI(
        C[403]), .CO(C[404]) );
  FA_13222 \FA_INST_0[0].FA_INST_1[404].FA_  ( .A(A[404]), .B(n1432), .CI(
        C[404]), .CO(C[405]) );
  FA_13221 \FA_INST_0[0].FA_INST_1[405].FA_  ( .A(A[405]), .B(n1433), .CI(
        C[405]), .CO(C[406]) );
  FA_13220 \FA_INST_0[0].FA_INST_1[406].FA_  ( .A(A[406]), .B(n1434), .CI(
        C[406]), .CO(C[407]) );
  FA_13219 \FA_INST_0[0].FA_INST_1[407].FA_  ( .A(A[407]), .B(n1435), .CI(
        C[407]), .CO(C[408]) );
  FA_13218 \FA_INST_0[0].FA_INST_1[408].FA_  ( .A(A[408]), .B(n1436), .CI(
        C[408]), .CO(C[409]) );
  FA_13217 \FA_INST_0[0].FA_INST_1[409].FA_  ( .A(A[409]), .B(n1437), .CI(
        C[409]), .CO(C[410]) );
  FA_13216 \FA_INST_0[0].FA_INST_1[410].FA_  ( .A(A[410]), .B(n1438), .CI(
        C[410]), .CO(C[411]) );
  FA_13215 \FA_INST_0[0].FA_INST_1[411].FA_  ( .A(A[411]), .B(n1439), .CI(
        C[411]), .CO(C[412]) );
  FA_13214 \FA_INST_0[0].FA_INST_1[412].FA_  ( .A(A[412]), .B(n1440), .CI(
        C[412]), .CO(C[413]) );
  FA_13213 \FA_INST_0[0].FA_INST_1[413].FA_  ( .A(A[413]), .B(n1441), .CI(
        C[413]), .CO(C[414]) );
  FA_13212 \FA_INST_0[0].FA_INST_1[414].FA_  ( .A(A[414]), .B(n1442), .CI(
        C[414]), .CO(C[415]) );
  FA_13211 \FA_INST_0[0].FA_INST_1[415].FA_  ( .A(A[415]), .B(n1443), .CI(
        C[415]), .CO(C[416]) );
  FA_13210 \FA_INST_0[0].FA_INST_1[416].FA_  ( .A(A[416]), .B(n1444), .CI(
        C[416]), .CO(C[417]) );
  FA_13209 \FA_INST_0[0].FA_INST_1[417].FA_  ( .A(A[417]), .B(n1445), .CI(
        C[417]), .CO(C[418]) );
  FA_13208 \FA_INST_0[0].FA_INST_1[418].FA_  ( .A(A[418]), .B(n1446), .CI(
        C[418]), .CO(C[419]) );
  FA_13207 \FA_INST_0[0].FA_INST_1[419].FA_  ( .A(A[419]), .B(n1447), .CI(
        C[419]), .CO(C[420]) );
  FA_13206 \FA_INST_0[0].FA_INST_1[420].FA_  ( .A(A[420]), .B(n1448), .CI(
        C[420]), .CO(C[421]) );
  FA_13205 \FA_INST_0[0].FA_INST_1[421].FA_  ( .A(A[421]), .B(n1449), .CI(
        C[421]), .CO(C[422]) );
  FA_13204 \FA_INST_0[0].FA_INST_1[422].FA_  ( .A(A[422]), .B(n1450), .CI(
        C[422]), .CO(C[423]) );
  FA_13203 \FA_INST_0[0].FA_INST_1[423].FA_  ( .A(A[423]), .B(n1451), .CI(
        C[423]), .CO(C[424]) );
  FA_13202 \FA_INST_0[0].FA_INST_1[424].FA_  ( .A(A[424]), .B(n1452), .CI(
        C[424]), .CO(C[425]) );
  FA_13201 \FA_INST_0[0].FA_INST_1[425].FA_  ( .A(A[425]), .B(n1453), .CI(
        C[425]), .CO(C[426]) );
  FA_13200 \FA_INST_0[0].FA_INST_1[426].FA_  ( .A(A[426]), .B(n1454), .CI(
        C[426]), .CO(C[427]) );
  FA_13199 \FA_INST_0[0].FA_INST_1[427].FA_  ( .A(A[427]), .B(n1455), .CI(
        C[427]), .CO(C[428]) );
  FA_13198 \FA_INST_0[0].FA_INST_1[428].FA_  ( .A(A[428]), .B(n1456), .CI(
        C[428]), .CO(C[429]) );
  FA_13197 \FA_INST_0[0].FA_INST_1[429].FA_  ( .A(A[429]), .B(n1457), .CI(
        C[429]), .CO(C[430]) );
  FA_13196 \FA_INST_0[0].FA_INST_1[430].FA_  ( .A(A[430]), .B(n1458), .CI(
        C[430]), .CO(C[431]) );
  FA_13195 \FA_INST_0[0].FA_INST_1[431].FA_  ( .A(A[431]), .B(n1459), .CI(
        C[431]), .CO(C[432]) );
  FA_13194 \FA_INST_0[0].FA_INST_1[432].FA_  ( .A(A[432]), .B(n1460), .CI(
        C[432]), .CO(C[433]) );
  FA_13193 \FA_INST_0[0].FA_INST_1[433].FA_  ( .A(A[433]), .B(n1461), .CI(
        C[433]), .CO(C[434]) );
  FA_13192 \FA_INST_0[0].FA_INST_1[434].FA_  ( .A(A[434]), .B(n1462), .CI(
        C[434]), .CO(C[435]) );
  FA_13191 \FA_INST_0[0].FA_INST_1[435].FA_  ( .A(A[435]), .B(n1463), .CI(
        C[435]), .CO(C[436]) );
  FA_13190 \FA_INST_0[0].FA_INST_1[436].FA_  ( .A(A[436]), .B(n1464), .CI(
        C[436]), .CO(C[437]) );
  FA_13189 \FA_INST_0[0].FA_INST_1[437].FA_  ( .A(A[437]), .B(n1465), .CI(
        C[437]), .CO(C[438]) );
  FA_13188 \FA_INST_0[0].FA_INST_1[438].FA_  ( .A(A[438]), .B(n1466), .CI(
        C[438]), .CO(C[439]) );
  FA_13187 \FA_INST_0[0].FA_INST_1[439].FA_  ( .A(A[439]), .B(n1467), .CI(
        C[439]), .CO(C[440]) );
  FA_13186 \FA_INST_0[0].FA_INST_1[440].FA_  ( .A(A[440]), .B(n1468), .CI(
        C[440]), .CO(C[441]) );
  FA_13185 \FA_INST_0[0].FA_INST_1[441].FA_  ( .A(A[441]), .B(n1469), .CI(
        C[441]), .CO(C[442]) );
  FA_13184 \FA_INST_0[0].FA_INST_1[442].FA_  ( .A(A[442]), .B(n1470), .CI(
        C[442]), .CO(C[443]) );
  FA_13183 \FA_INST_0[0].FA_INST_1[443].FA_  ( .A(A[443]), .B(n1471), .CI(
        C[443]), .CO(C[444]) );
  FA_13182 \FA_INST_0[0].FA_INST_1[444].FA_  ( .A(A[444]), .B(n1472), .CI(
        C[444]), .CO(C[445]) );
  FA_13181 \FA_INST_0[0].FA_INST_1[445].FA_  ( .A(A[445]), .B(n1473), .CI(
        C[445]), .CO(C[446]) );
  FA_13180 \FA_INST_0[0].FA_INST_1[446].FA_  ( .A(A[446]), .B(n1474), .CI(
        C[446]), .CO(C[447]) );
  FA_13179 \FA_INST_0[0].FA_INST_1[447].FA_  ( .A(A[447]), .B(n1475), .CI(
        C[447]), .CO(C[448]) );
  FA_13178 \FA_INST_0[0].FA_INST_1[448].FA_  ( .A(A[448]), .B(n1476), .CI(
        C[448]), .CO(C[449]) );
  FA_13177 \FA_INST_0[0].FA_INST_1[449].FA_  ( .A(A[449]), .B(n1477), .CI(
        C[449]), .CO(C[450]) );
  FA_13176 \FA_INST_0[0].FA_INST_1[450].FA_  ( .A(A[450]), .B(n1478), .CI(
        C[450]), .CO(C[451]) );
  FA_13175 \FA_INST_0[0].FA_INST_1[451].FA_  ( .A(A[451]), .B(n1479), .CI(
        C[451]), .CO(C[452]) );
  FA_13174 \FA_INST_0[0].FA_INST_1[452].FA_  ( .A(A[452]), .B(n1480), .CI(
        C[452]), .CO(C[453]) );
  FA_13173 \FA_INST_0[0].FA_INST_1[453].FA_  ( .A(A[453]), .B(n1481), .CI(
        C[453]), .CO(C[454]) );
  FA_13172 \FA_INST_0[0].FA_INST_1[454].FA_  ( .A(A[454]), .B(n1482), .CI(
        C[454]), .CO(C[455]) );
  FA_13171 \FA_INST_0[0].FA_INST_1[455].FA_  ( .A(A[455]), .B(n1483), .CI(
        C[455]), .CO(C[456]) );
  FA_13170 \FA_INST_0[0].FA_INST_1[456].FA_  ( .A(A[456]), .B(n1484), .CI(
        C[456]), .CO(C[457]) );
  FA_13169 \FA_INST_0[0].FA_INST_1[457].FA_  ( .A(A[457]), .B(n1485), .CI(
        C[457]), .CO(C[458]) );
  FA_13168 \FA_INST_0[0].FA_INST_1[458].FA_  ( .A(A[458]), .B(n1486), .CI(
        C[458]), .CO(C[459]) );
  FA_13167 \FA_INST_0[0].FA_INST_1[459].FA_  ( .A(A[459]), .B(n1487), .CI(
        C[459]), .CO(C[460]) );
  FA_13166 \FA_INST_0[0].FA_INST_1[460].FA_  ( .A(A[460]), .B(n1488), .CI(
        C[460]), .CO(C[461]) );
  FA_13165 \FA_INST_0[0].FA_INST_1[461].FA_  ( .A(A[461]), .B(n1489), .CI(
        C[461]), .CO(C[462]) );
  FA_13164 \FA_INST_0[0].FA_INST_1[462].FA_  ( .A(A[462]), .B(n1490), .CI(
        C[462]), .CO(C[463]) );
  FA_13163 \FA_INST_0[0].FA_INST_1[463].FA_  ( .A(A[463]), .B(n1491), .CI(
        C[463]), .CO(C[464]) );
  FA_13162 \FA_INST_0[0].FA_INST_1[464].FA_  ( .A(A[464]), .B(n1492), .CI(
        C[464]), .CO(C[465]) );
  FA_13161 \FA_INST_0[0].FA_INST_1[465].FA_  ( .A(A[465]), .B(n1493), .CI(
        C[465]), .CO(C[466]) );
  FA_13160 \FA_INST_0[0].FA_INST_1[466].FA_  ( .A(A[466]), .B(n1494), .CI(
        C[466]), .CO(C[467]) );
  FA_13159 \FA_INST_0[0].FA_INST_1[467].FA_  ( .A(A[467]), .B(n1495), .CI(
        C[467]), .CO(C[468]) );
  FA_13158 \FA_INST_0[0].FA_INST_1[468].FA_  ( .A(A[468]), .B(n1496), .CI(
        C[468]), .CO(C[469]) );
  FA_13157 \FA_INST_0[0].FA_INST_1[469].FA_  ( .A(A[469]), .B(n1497), .CI(
        C[469]), .CO(C[470]) );
  FA_13156 \FA_INST_0[0].FA_INST_1[470].FA_  ( .A(A[470]), .B(n1498), .CI(
        C[470]), .CO(C[471]) );
  FA_13155 \FA_INST_0[0].FA_INST_1[471].FA_  ( .A(A[471]), .B(n1499), .CI(
        C[471]), .CO(C[472]) );
  FA_13154 \FA_INST_0[0].FA_INST_1[472].FA_  ( .A(A[472]), .B(n1500), .CI(
        C[472]), .CO(C[473]) );
  FA_13153 \FA_INST_0[0].FA_INST_1[473].FA_  ( .A(A[473]), .B(n1501), .CI(
        C[473]), .CO(C[474]) );
  FA_13152 \FA_INST_0[0].FA_INST_1[474].FA_  ( .A(A[474]), .B(n1502), .CI(
        C[474]), .CO(C[475]) );
  FA_13151 \FA_INST_0[0].FA_INST_1[475].FA_  ( .A(A[475]), .B(n1503), .CI(
        C[475]), .CO(C[476]) );
  FA_13150 \FA_INST_0[0].FA_INST_1[476].FA_  ( .A(A[476]), .B(n1504), .CI(
        C[476]), .CO(C[477]) );
  FA_13149 \FA_INST_0[0].FA_INST_1[477].FA_  ( .A(A[477]), .B(n1505), .CI(
        C[477]), .CO(C[478]) );
  FA_13148 \FA_INST_0[0].FA_INST_1[478].FA_  ( .A(A[478]), .B(n1506), .CI(
        C[478]), .CO(C[479]) );
  FA_13147 \FA_INST_0[0].FA_INST_1[479].FA_  ( .A(A[479]), .B(n1507), .CI(
        C[479]), .CO(C[480]) );
  FA_13146 \FA_INST_0[0].FA_INST_1[480].FA_  ( .A(A[480]), .B(n1508), .CI(
        C[480]), .CO(C[481]) );
  FA_13145 \FA_INST_0[0].FA_INST_1[481].FA_  ( .A(A[481]), .B(n1509), .CI(
        C[481]), .CO(C[482]) );
  FA_13144 \FA_INST_0[0].FA_INST_1[482].FA_  ( .A(A[482]), .B(n1510), .CI(
        C[482]), .CO(C[483]) );
  FA_13143 \FA_INST_0[0].FA_INST_1[483].FA_  ( .A(A[483]), .B(n1511), .CI(
        C[483]), .CO(C[484]) );
  FA_13142 \FA_INST_0[0].FA_INST_1[484].FA_  ( .A(A[484]), .B(n1512), .CI(
        C[484]), .CO(C[485]) );
  FA_13141 \FA_INST_0[0].FA_INST_1[485].FA_  ( .A(A[485]), .B(n1513), .CI(
        C[485]), .CO(C[486]) );
  FA_13140 \FA_INST_0[0].FA_INST_1[486].FA_  ( .A(A[486]), .B(n1514), .CI(
        C[486]), .CO(C[487]) );
  FA_13139 \FA_INST_0[0].FA_INST_1[487].FA_  ( .A(A[487]), .B(n1515), .CI(
        C[487]), .CO(C[488]) );
  FA_13138 \FA_INST_0[0].FA_INST_1[488].FA_  ( .A(A[488]), .B(n1516), .CI(
        C[488]), .CO(C[489]) );
  FA_13137 \FA_INST_0[0].FA_INST_1[489].FA_  ( .A(A[489]), .B(n1517), .CI(
        C[489]), .CO(C[490]) );
  FA_13136 \FA_INST_0[0].FA_INST_1[490].FA_  ( .A(A[490]), .B(n1518), .CI(
        C[490]), .CO(C[491]) );
  FA_13135 \FA_INST_0[0].FA_INST_1[491].FA_  ( .A(A[491]), .B(n1519), .CI(
        C[491]), .CO(C[492]) );
  FA_13134 \FA_INST_0[0].FA_INST_1[492].FA_  ( .A(A[492]), .B(n1520), .CI(
        C[492]), .CO(C[493]) );
  FA_13133 \FA_INST_0[0].FA_INST_1[493].FA_  ( .A(A[493]), .B(n1521), .CI(
        C[493]), .CO(C[494]) );
  FA_13132 \FA_INST_0[0].FA_INST_1[494].FA_  ( .A(A[494]), .B(n1522), .CI(
        C[494]), .CO(C[495]) );
  FA_13131 \FA_INST_0[0].FA_INST_1[495].FA_  ( .A(A[495]), .B(n1523), .CI(
        C[495]), .CO(C[496]) );
  FA_13130 \FA_INST_0[0].FA_INST_1[496].FA_  ( .A(A[496]), .B(n1524), .CI(
        C[496]), .CO(C[497]) );
  FA_13129 \FA_INST_0[0].FA_INST_1[497].FA_  ( .A(A[497]), .B(n1525), .CI(
        C[497]), .CO(C[498]) );
  FA_13128 \FA_INST_0[0].FA_INST_1[498].FA_  ( .A(A[498]), .B(n1526), .CI(
        C[498]), .CO(C[499]) );
  FA_13127 \FA_INST_0[0].FA_INST_1[499].FA_  ( .A(A[499]), .B(n1527), .CI(
        C[499]), .CO(C[500]) );
  FA_13126 \FA_INST_0[0].FA_INST_1[500].FA_  ( .A(A[500]), .B(n1528), .CI(
        C[500]), .CO(C[501]) );
  FA_13125 \FA_INST_0[0].FA_INST_1[501].FA_  ( .A(A[501]), .B(n1529), .CI(
        C[501]), .CO(C[502]) );
  FA_13124 \FA_INST_0[0].FA_INST_1[502].FA_  ( .A(A[502]), .B(n1530), .CI(
        C[502]), .CO(C[503]) );
  FA_13123 \FA_INST_0[0].FA_INST_1[503].FA_  ( .A(A[503]), .B(n1531), .CI(
        C[503]), .CO(C[504]) );
  FA_13122 \FA_INST_0[0].FA_INST_1[504].FA_  ( .A(A[504]), .B(n1532), .CI(
        C[504]), .CO(C[505]) );
  FA_13121 \FA_INST_0[0].FA_INST_1[505].FA_  ( .A(A[505]), .B(n1533), .CI(
        C[505]), .CO(C[506]) );
  FA_13120 \FA_INST_0[0].FA_INST_1[506].FA_  ( .A(A[506]), .B(n1534), .CI(
        C[506]), .CO(C[507]) );
  FA_13119 \FA_INST_0[0].FA_INST_1[507].FA_  ( .A(A[507]), .B(n1535), .CI(
        C[507]), .CO(C[508]) );
  FA_13118 \FA_INST_0[0].FA_INST_1[508].FA_  ( .A(A[508]), .B(n1536), .CI(
        C[508]), .CO(C[509]) );
  FA_13117 \FA_INST_0[0].FA_INST_1[509].FA_  ( .A(A[509]), .B(n1537), .CI(
        C[509]), .CO(C[510]) );
  FA_13116 \FA_INST_0[0].FA_INST_1[510].FA_  ( .A(A[510]), .B(n1538), .CI(
        C[510]), .CO(C[511]) );
  FA_13115 \FA_INST_0[0].FA_INST_1[511].FA_  ( .A(A[511]), .B(n1539), .CI(
        C[511]), .CO(C[512]) );
  FA_13114 \FA_INST_0[1].FA_INST_1[0].FA_  ( .A(A[512]), .B(n1540), .CI(C[512]), .CO(C[513]) );
  FA_13113 \FA_INST_0[1].FA_INST_1[1].FA_  ( .A(A[513]), .B(n1541), .CI(C[513]), .CO(C[514]) );
  FA_13112 \FA_INST_0[1].FA_INST_1[2].FA_  ( .A(A[514]), .B(n1542), .CI(C[514]), .CO(C[515]) );
  FA_13111 \FA_INST_0[1].FA_INST_1[3].FA_  ( .A(A[515]), .B(n1543), .CI(C[515]), .CO(C[516]) );
  FA_13110 \FA_INST_0[1].FA_INST_1[4].FA_  ( .A(A[516]), .B(n1544), .CI(C[516]), .CO(C[517]) );
  FA_13109 \FA_INST_0[1].FA_INST_1[5].FA_  ( .A(A[517]), .B(n1545), .CI(C[517]), .CO(C[518]) );
  FA_13108 \FA_INST_0[1].FA_INST_1[6].FA_  ( .A(A[518]), .B(n1546), .CI(C[518]), .CO(C[519]) );
  FA_13107 \FA_INST_0[1].FA_INST_1[7].FA_  ( .A(A[519]), .B(n1547), .CI(C[519]), .CO(C[520]) );
  FA_13106 \FA_INST_0[1].FA_INST_1[8].FA_  ( .A(A[520]), .B(n1548), .CI(C[520]), .CO(C[521]) );
  FA_13105 \FA_INST_0[1].FA_INST_1[9].FA_  ( .A(A[521]), .B(n1549), .CI(C[521]), .CO(C[522]) );
  FA_13104 \FA_INST_0[1].FA_INST_1[10].FA_  ( .A(A[522]), .B(n1550), .CI(
        C[522]), .CO(C[523]) );
  FA_13103 \FA_INST_0[1].FA_INST_1[11].FA_  ( .A(A[523]), .B(n1551), .CI(
        C[523]), .CO(C[524]) );
  FA_13102 \FA_INST_0[1].FA_INST_1[12].FA_  ( .A(A[524]), .B(n1552), .CI(
        C[524]), .CO(C[525]) );
  FA_13101 \FA_INST_0[1].FA_INST_1[13].FA_  ( .A(A[525]), .B(n1553), .CI(
        C[525]), .CO(C[526]) );
  FA_13100 \FA_INST_0[1].FA_INST_1[14].FA_  ( .A(A[526]), .B(n1554), .CI(
        C[526]), .CO(C[527]) );
  FA_13099 \FA_INST_0[1].FA_INST_1[15].FA_  ( .A(A[527]), .B(n1555), .CI(
        C[527]), .CO(C[528]) );
  FA_13098 \FA_INST_0[1].FA_INST_1[16].FA_  ( .A(A[528]), .B(n1556), .CI(
        C[528]), .CO(C[529]) );
  FA_13097 \FA_INST_0[1].FA_INST_1[17].FA_  ( .A(A[529]), .B(n1557), .CI(
        C[529]), .CO(C[530]) );
  FA_13096 \FA_INST_0[1].FA_INST_1[18].FA_  ( .A(A[530]), .B(n1558), .CI(
        C[530]), .CO(C[531]) );
  FA_13095 \FA_INST_0[1].FA_INST_1[19].FA_  ( .A(A[531]), .B(n1559), .CI(
        C[531]), .CO(C[532]) );
  FA_13094 \FA_INST_0[1].FA_INST_1[20].FA_  ( .A(A[532]), .B(n1560), .CI(
        C[532]), .CO(C[533]) );
  FA_13093 \FA_INST_0[1].FA_INST_1[21].FA_  ( .A(A[533]), .B(n1561), .CI(
        C[533]), .CO(C[534]) );
  FA_13092 \FA_INST_0[1].FA_INST_1[22].FA_  ( .A(A[534]), .B(n1562), .CI(
        C[534]), .CO(C[535]) );
  FA_13091 \FA_INST_0[1].FA_INST_1[23].FA_  ( .A(A[535]), .B(n1563), .CI(
        C[535]), .CO(C[536]) );
  FA_13090 \FA_INST_0[1].FA_INST_1[24].FA_  ( .A(A[536]), .B(n1564), .CI(
        C[536]), .CO(C[537]) );
  FA_13089 \FA_INST_0[1].FA_INST_1[25].FA_  ( .A(A[537]), .B(n1565), .CI(
        C[537]), .CO(C[538]) );
  FA_13088 \FA_INST_0[1].FA_INST_1[26].FA_  ( .A(A[538]), .B(n1566), .CI(
        C[538]), .CO(C[539]) );
  FA_13087 \FA_INST_0[1].FA_INST_1[27].FA_  ( .A(A[539]), .B(n1567), .CI(
        C[539]), .CO(C[540]) );
  FA_13086 \FA_INST_0[1].FA_INST_1[28].FA_  ( .A(A[540]), .B(n1568), .CI(
        C[540]), .CO(C[541]) );
  FA_13085 \FA_INST_0[1].FA_INST_1[29].FA_  ( .A(A[541]), .B(n1569), .CI(
        C[541]), .CO(C[542]) );
  FA_13084 \FA_INST_0[1].FA_INST_1[30].FA_  ( .A(A[542]), .B(n1570), .CI(
        C[542]), .CO(C[543]) );
  FA_13083 \FA_INST_0[1].FA_INST_1[31].FA_  ( .A(A[543]), .B(n1571), .CI(
        C[543]), .CO(C[544]) );
  FA_13082 \FA_INST_0[1].FA_INST_1[32].FA_  ( .A(A[544]), .B(n1572), .CI(
        C[544]), .CO(C[545]) );
  FA_13081 \FA_INST_0[1].FA_INST_1[33].FA_  ( .A(A[545]), .B(n1573), .CI(
        C[545]), .CO(C[546]) );
  FA_13080 \FA_INST_0[1].FA_INST_1[34].FA_  ( .A(A[546]), .B(n1574), .CI(
        C[546]), .CO(C[547]) );
  FA_13079 \FA_INST_0[1].FA_INST_1[35].FA_  ( .A(A[547]), .B(n1575), .CI(
        C[547]), .CO(C[548]) );
  FA_13078 \FA_INST_0[1].FA_INST_1[36].FA_  ( .A(A[548]), .B(n1576), .CI(
        C[548]), .CO(C[549]) );
  FA_13077 \FA_INST_0[1].FA_INST_1[37].FA_  ( .A(A[549]), .B(n1577), .CI(
        C[549]), .CO(C[550]) );
  FA_13076 \FA_INST_0[1].FA_INST_1[38].FA_  ( .A(A[550]), .B(n1578), .CI(
        C[550]), .CO(C[551]) );
  FA_13075 \FA_INST_0[1].FA_INST_1[39].FA_  ( .A(A[551]), .B(n1579), .CI(
        C[551]), .CO(C[552]) );
  FA_13074 \FA_INST_0[1].FA_INST_1[40].FA_  ( .A(A[552]), .B(n1580), .CI(
        C[552]), .CO(C[553]) );
  FA_13073 \FA_INST_0[1].FA_INST_1[41].FA_  ( .A(A[553]), .B(n1581), .CI(
        C[553]), .CO(C[554]) );
  FA_13072 \FA_INST_0[1].FA_INST_1[42].FA_  ( .A(A[554]), .B(n1582), .CI(
        C[554]), .CO(C[555]) );
  FA_13071 \FA_INST_0[1].FA_INST_1[43].FA_  ( .A(A[555]), .B(n1583), .CI(
        C[555]), .CO(C[556]) );
  FA_13070 \FA_INST_0[1].FA_INST_1[44].FA_  ( .A(A[556]), .B(n1584), .CI(
        C[556]), .CO(C[557]) );
  FA_13069 \FA_INST_0[1].FA_INST_1[45].FA_  ( .A(A[557]), .B(n1585), .CI(
        C[557]), .CO(C[558]) );
  FA_13068 \FA_INST_0[1].FA_INST_1[46].FA_  ( .A(A[558]), .B(n1586), .CI(
        C[558]), .CO(C[559]) );
  FA_13067 \FA_INST_0[1].FA_INST_1[47].FA_  ( .A(A[559]), .B(n1587), .CI(
        C[559]), .CO(C[560]) );
  FA_13066 \FA_INST_0[1].FA_INST_1[48].FA_  ( .A(A[560]), .B(n1588), .CI(
        C[560]), .CO(C[561]) );
  FA_13065 \FA_INST_0[1].FA_INST_1[49].FA_  ( .A(A[561]), .B(n1589), .CI(
        C[561]), .CO(C[562]) );
  FA_13064 \FA_INST_0[1].FA_INST_1[50].FA_  ( .A(A[562]), .B(n1590), .CI(
        C[562]), .CO(C[563]) );
  FA_13063 \FA_INST_0[1].FA_INST_1[51].FA_  ( .A(A[563]), .B(n1591), .CI(
        C[563]), .CO(C[564]) );
  FA_13062 \FA_INST_0[1].FA_INST_1[52].FA_  ( .A(A[564]), .B(n1592), .CI(
        C[564]), .CO(C[565]) );
  FA_13061 \FA_INST_0[1].FA_INST_1[53].FA_  ( .A(A[565]), .B(n1593), .CI(
        C[565]), .CO(C[566]) );
  FA_13060 \FA_INST_0[1].FA_INST_1[54].FA_  ( .A(A[566]), .B(n1594), .CI(
        C[566]), .CO(C[567]) );
  FA_13059 \FA_INST_0[1].FA_INST_1[55].FA_  ( .A(A[567]), .B(n1595), .CI(
        C[567]), .CO(C[568]) );
  FA_13058 \FA_INST_0[1].FA_INST_1[56].FA_  ( .A(A[568]), .B(n1596), .CI(
        C[568]), .CO(C[569]) );
  FA_13057 \FA_INST_0[1].FA_INST_1[57].FA_  ( .A(A[569]), .B(n1597), .CI(
        C[569]), .CO(C[570]) );
  FA_13056 \FA_INST_0[1].FA_INST_1[58].FA_  ( .A(A[570]), .B(n1598), .CI(
        C[570]), .CO(C[571]) );
  FA_13055 \FA_INST_0[1].FA_INST_1[59].FA_  ( .A(A[571]), .B(n1599), .CI(
        C[571]), .CO(C[572]) );
  FA_13054 \FA_INST_0[1].FA_INST_1[60].FA_  ( .A(A[572]), .B(n1600), .CI(
        C[572]), .CO(C[573]) );
  FA_13053 \FA_INST_0[1].FA_INST_1[61].FA_  ( .A(A[573]), .B(n1601), .CI(
        C[573]), .CO(C[574]) );
  FA_13052 \FA_INST_0[1].FA_INST_1[62].FA_  ( .A(A[574]), .B(n1602), .CI(
        C[574]), .CO(C[575]) );
  FA_13051 \FA_INST_0[1].FA_INST_1[63].FA_  ( .A(A[575]), .B(n1603), .CI(
        C[575]), .CO(C[576]) );
  FA_13050 \FA_INST_0[1].FA_INST_1[64].FA_  ( .A(A[576]), .B(n1604), .CI(
        C[576]), .CO(C[577]) );
  FA_13049 \FA_INST_0[1].FA_INST_1[65].FA_  ( .A(A[577]), .B(n1605), .CI(
        C[577]), .CO(C[578]) );
  FA_13048 \FA_INST_0[1].FA_INST_1[66].FA_  ( .A(A[578]), .B(n1606), .CI(
        C[578]), .CO(C[579]) );
  FA_13047 \FA_INST_0[1].FA_INST_1[67].FA_  ( .A(A[579]), .B(n1607), .CI(
        C[579]), .CO(C[580]) );
  FA_13046 \FA_INST_0[1].FA_INST_1[68].FA_  ( .A(A[580]), .B(n1608), .CI(
        C[580]), .CO(C[581]) );
  FA_13045 \FA_INST_0[1].FA_INST_1[69].FA_  ( .A(A[581]), .B(n1609), .CI(
        C[581]), .CO(C[582]) );
  FA_13044 \FA_INST_0[1].FA_INST_1[70].FA_  ( .A(A[582]), .B(n1610), .CI(
        C[582]), .CO(C[583]) );
  FA_13043 \FA_INST_0[1].FA_INST_1[71].FA_  ( .A(A[583]), .B(n1611), .CI(
        C[583]), .CO(C[584]) );
  FA_13042 \FA_INST_0[1].FA_INST_1[72].FA_  ( .A(A[584]), .B(n1612), .CI(
        C[584]), .CO(C[585]) );
  FA_13041 \FA_INST_0[1].FA_INST_1[73].FA_  ( .A(A[585]), .B(n1613), .CI(
        C[585]), .CO(C[586]) );
  FA_13040 \FA_INST_0[1].FA_INST_1[74].FA_  ( .A(A[586]), .B(n1614), .CI(
        C[586]), .CO(C[587]) );
  FA_13039 \FA_INST_0[1].FA_INST_1[75].FA_  ( .A(A[587]), .B(n1615), .CI(
        C[587]), .CO(C[588]) );
  FA_13038 \FA_INST_0[1].FA_INST_1[76].FA_  ( .A(A[588]), .B(n1616), .CI(
        C[588]), .CO(C[589]) );
  FA_13037 \FA_INST_0[1].FA_INST_1[77].FA_  ( .A(A[589]), .B(n1617), .CI(
        C[589]), .CO(C[590]) );
  FA_13036 \FA_INST_0[1].FA_INST_1[78].FA_  ( .A(A[590]), .B(n1618), .CI(
        C[590]), .CO(C[591]) );
  FA_13035 \FA_INST_0[1].FA_INST_1[79].FA_  ( .A(A[591]), .B(n1619), .CI(
        C[591]), .CO(C[592]) );
  FA_13034 \FA_INST_0[1].FA_INST_1[80].FA_  ( .A(A[592]), .B(n1620), .CI(
        C[592]), .CO(C[593]) );
  FA_13033 \FA_INST_0[1].FA_INST_1[81].FA_  ( .A(A[593]), .B(n1621), .CI(
        C[593]), .CO(C[594]) );
  FA_13032 \FA_INST_0[1].FA_INST_1[82].FA_  ( .A(A[594]), .B(n1622), .CI(
        C[594]), .CO(C[595]) );
  FA_13031 \FA_INST_0[1].FA_INST_1[83].FA_  ( .A(A[595]), .B(n1623), .CI(
        C[595]), .CO(C[596]) );
  FA_13030 \FA_INST_0[1].FA_INST_1[84].FA_  ( .A(A[596]), .B(n1624), .CI(
        C[596]), .CO(C[597]) );
  FA_13029 \FA_INST_0[1].FA_INST_1[85].FA_  ( .A(A[597]), .B(n1625), .CI(
        C[597]), .CO(C[598]) );
  FA_13028 \FA_INST_0[1].FA_INST_1[86].FA_  ( .A(A[598]), .B(n1626), .CI(
        C[598]), .CO(C[599]) );
  FA_13027 \FA_INST_0[1].FA_INST_1[87].FA_  ( .A(A[599]), .B(n1627), .CI(
        C[599]), .CO(C[600]) );
  FA_13026 \FA_INST_0[1].FA_INST_1[88].FA_  ( .A(A[600]), .B(n1628), .CI(
        C[600]), .CO(C[601]) );
  FA_13025 \FA_INST_0[1].FA_INST_1[89].FA_  ( .A(A[601]), .B(n1629), .CI(
        C[601]), .CO(C[602]) );
  FA_13024 \FA_INST_0[1].FA_INST_1[90].FA_  ( .A(A[602]), .B(n1630), .CI(
        C[602]), .CO(C[603]) );
  FA_13023 \FA_INST_0[1].FA_INST_1[91].FA_  ( .A(A[603]), .B(n1631), .CI(
        C[603]), .CO(C[604]) );
  FA_13022 \FA_INST_0[1].FA_INST_1[92].FA_  ( .A(A[604]), .B(n1632), .CI(
        C[604]), .CO(C[605]) );
  FA_13021 \FA_INST_0[1].FA_INST_1[93].FA_  ( .A(A[605]), .B(n1633), .CI(
        C[605]), .CO(C[606]) );
  FA_13020 \FA_INST_0[1].FA_INST_1[94].FA_  ( .A(A[606]), .B(n1634), .CI(
        C[606]), .CO(C[607]) );
  FA_13019 \FA_INST_0[1].FA_INST_1[95].FA_  ( .A(A[607]), .B(n1635), .CI(
        C[607]), .CO(C[608]) );
  FA_13018 \FA_INST_0[1].FA_INST_1[96].FA_  ( .A(A[608]), .B(n1636), .CI(
        C[608]), .CO(C[609]) );
  FA_13017 \FA_INST_0[1].FA_INST_1[97].FA_  ( .A(A[609]), .B(n1637), .CI(
        C[609]), .CO(C[610]) );
  FA_13016 \FA_INST_0[1].FA_INST_1[98].FA_  ( .A(A[610]), .B(n1638), .CI(
        C[610]), .CO(C[611]) );
  FA_13015 \FA_INST_0[1].FA_INST_1[99].FA_  ( .A(A[611]), .B(n1639), .CI(
        C[611]), .CO(C[612]) );
  FA_13014 \FA_INST_0[1].FA_INST_1[100].FA_  ( .A(A[612]), .B(n1640), .CI(
        C[612]), .CO(C[613]) );
  FA_13013 \FA_INST_0[1].FA_INST_1[101].FA_  ( .A(A[613]), .B(n1641), .CI(
        C[613]), .CO(C[614]) );
  FA_13012 \FA_INST_0[1].FA_INST_1[102].FA_  ( .A(A[614]), .B(n1642), .CI(
        C[614]), .CO(C[615]) );
  FA_13011 \FA_INST_0[1].FA_INST_1[103].FA_  ( .A(A[615]), .B(n1643), .CI(
        C[615]), .CO(C[616]) );
  FA_13010 \FA_INST_0[1].FA_INST_1[104].FA_  ( .A(A[616]), .B(n1644), .CI(
        C[616]), .CO(C[617]) );
  FA_13009 \FA_INST_0[1].FA_INST_1[105].FA_  ( .A(A[617]), .B(n1645), .CI(
        C[617]), .CO(C[618]) );
  FA_13008 \FA_INST_0[1].FA_INST_1[106].FA_  ( .A(A[618]), .B(n1646), .CI(
        C[618]), .CO(C[619]) );
  FA_13007 \FA_INST_0[1].FA_INST_1[107].FA_  ( .A(A[619]), .B(n1647), .CI(
        C[619]), .CO(C[620]) );
  FA_13006 \FA_INST_0[1].FA_INST_1[108].FA_  ( .A(A[620]), .B(n1648), .CI(
        C[620]), .CO(C[621]) );
  FA_13005 \FA_INST_0[1].FA_INST_1[109].FA_  ( .A(A[621]), .B(n1649), .CI(
        C[621]), .CO(C[622]) );
  FA_13004 \FA_INST_0[1].FA_INST_1[110].FA_  ( .A(A[622]), .B(n1650), .CI(
        C[622]), .CO(C[623]) );
  FA_13003 \FA_INST_0[1].FA_INST_1[111].FA_  ( .A(A[623]), .B(n1651), .CI(
        C[623]), .CO(C[624]) );
  FA_13002 \FA_INST_0[1].FA_INST_1[112].FA_  ( .A(A[624]), .B(n1652), .CI(
        C[624]), .CO(C[625]) );
  FA_13001 \FA_INST_0[1].FA_INST_1[113].FA_  ( .A(A[625]), .B(n1653), .CI(
        C[625]), .CO(C[626]) );
  FA_13000 \FA_INST_0[1].FA_INST_1[114].FA_  ( .A(A[626]), .B(n1654), .CI(
        C[626]), .CO(C[627]) );
  FA_12999 \FA_INST_0[1].FA_INST_1[115].FA_  ( .A(A[627]), .B(n1655), .CI(
        C[627]), .CO(C[628]) );
  FA_12998 \FA_INST_0[1].FA_INST_1[116].FA_  ( .A(A[628]), .B(n1656), .CI(
        C[628]), .CO(C[629]) );
  FA_12997 \FA_INST_0[1].FA_INST_1[117].FA_  ( .A(A[629]), .B(n1657), .CI(
        C[629]), .CO(C[630]) );
  FA_12996 \FA_INST_0[1].FA_INST_1[118].FA_  ( .A(A[630]), .B(n1658), .CI(
        C[630]), .CO(C[631]) );
  FA_12995 \FA_INST_0[1].FA_INST_1[119].FA_  ( .A(A[631]), .B(n1659), .CI(
        C[631]), .CO(C[632]) );
  FA_12994 \FA_INST_0[1].FA_INST_1[120].FA_  ( .A(A[632]), .B(n1660), .CI(
        C[632]), .CO(C[633]) );
  FA_12993 \FA_INST_0[1].FA_INST_1[121].FA_  ( .A(A[633]), .B(n1661), .CI(
        C[633]), .CO(C[634]) );
  FA_12992 \FA_INST_0[1].FA_INST_1[122].FA_  ( .A(A[634]), .B(n1662), .CI(
        C[634]), .CO(C[635]) );
  FA_12991 \FA_INST_0[1].FA_INST_1[123].FA_  ( .A(A[635]), .B(n1663), .CI(
        C[635]), .CO(C[636]) );
  FA_12990 \FA_INST_0[1].FA_INST_1[124].FA_  ( .A(A[636]), .B(n1664), .CI(
        C[636]), .CO(C[637]) );
  FA_12989 \FA_INST_0[1].FA_INST_1[125].FA_  ( .A(A[637]), .B(n1665), .CI(
        C[637]), .CO(C[638]) );
  FA_12988 \FA_INST_0[1].FA_INST_1[126].FA_  ( .A(A[638]), .B(n1666), .CI(
        C[638]), .CO(C[639]) );
  FA_12987 \FA_INST_0[1].FA_INST_1[127].FA_  ( .A(A[639]), .B(n1667), .CI(
        C[639]), .CO(C[640]) );
  FA_12986 \FA_INST_0[1].FA_INST_1[128].FA_  ( .A(A[640]), .B(n1668), .CI(
        C[640]), .CO(C[641]) );
  FA_12985 \FA_INST_0[1].FA_INST_1[129].FA_  ( .A(A[641]), .B(n1669), .CI(
        C[641]), .CO(C[642]) );
  FA_12984 \FA_INST_0[1].FA_INST_1[130].FA_  ( .A(A[642]), .B(n1670), .CI(
        C[642]), .CO(C[643]) );
  FA_12983 \FA_INST_0[1].FA_INST_1[131].FA_  ( .A(A[643]), .B(n1671), .CI(
        C[643]), .CO(C[644]) );
  FA_12982 \FA_INST_0[1].FA_INST_1[132].FA_  ( .A(A[644]), .B(n1672), .CI(
        C[644]), .CO(C[645]) );
  FA_12981 \FA_INST_0[1].FA_INST_1[133].FA_  ( .A(A[645]), .B(n1673), .CI(
        C[645]), .CO(C[646]) );
  FA_12980 \FA_INST_0[1].FA_INST_1[134].FA_  ( .A(A[646]), .B(n1674), .CI(
        C[646]), .CO(C[647]) );
  FA_12979 \FA_INST_0[1].FA_INST_1[135].FA_  ( .A(A[647]), .B(n1675), .CI(
        C[647]), .CO(C[648]) );
  FA_12978 \FA_INST_0[1].FA_INST_1[136].FA_  ( .A(A[648]), .B(n1676), .CI(
        C[648]), .CO(C[649]) );
  FA_12977 \FA_INST_0[1].FA_INST_1[137].FA_  ( .A(A[649]), .B(n1677), .CI(
        C[649]), .CO(C[650]) );
  FA_12976 \FA_INST_0[1].FA_INST_1[138].FA_  ( .A(A[650]), .B(n1678), .CI(
        C[650]), .CO(C[651]) );
  FA_12975 \FA_INST_0[1].FA_INST_1[139].FA_  ( .A(A[651]), .B(n1679), .CI(
        C[651]), .CO(C[652]) );
  FA_12974 \FA_INST_0[1].FA_INST_1[140].FA_  ( .A(A[652]), .B(n1680), .CI(
        C[652]), .CO(C[653]) );
  FA_12973 \FA_INST_0[1].FA_INST_1[141].FA_  ( .A(A[653]), .B(n1681), .CI(
        C[653]), .CO(C[654]) );
  FA_12972 \FA_INST_0[1].FA_INST_1[142].FA_  ( .A(A[654]), .B(n1682), .CI(
        C[654]), .CO(C[655]) );
  FA_12971 \FA_INST_0[1].FA_INST_1[143].FA_  ( .A(A[655]), .B(n1683), .CI(
        C[655]), .CO(C[656]) );
  FA_12970 \FA_INST_0[1].FA_INST_1[144].FA_  ( .A(A[656]), .B(n1684), .CI(
        C[656]), .CO(C[657]) );
  FA_12969 \FA_INST_0[1].FA_INST_1[145].FA_  ( .A(A[657]), .B(n1685), .CI(
        C[657]), .CO(C[658]) );
  FA_12968 \FA_INST_0[1].FA_INST_1[146].FA_  ( .A(A[658]), .B(n1686), .CI(
        C[658]), .CO(C[659]) );
  FA_12967 \FA_INST_0[1].FA_INST_1[147].FA_  ( .A(A[659]), .B(n1687), .CI(
        C[659]), .CO(C[660]) );
  FA_12966 \FA_INST_0[1].FA_INST_1[148].FA_  ( .A(A[660]), .B(n1688), .CI(
        C[660]), .CO(C[661]) );
  FA_12965 \FA_INST_0[1].FA_INST_1[149].FA_  ( .A(A[661]), .B(n1689), .CI(
        C[661]), .CO(C[662]) );
  FA_12964 \FA_INST_0[1].FA_INST_1[150].FA_  ( .A(A[662]), .B(n1690), .CI(
        C[662]), .CO(C[663]) );
  FA_12963 \FA_INST_0[1].FA_INST_1[151].FA_  ( .A(A[663]), .B(n1691), .CI(
        C[663]), .CO(C[664]) );
  FA_12962 \FA_INST_0[1].FA_INST_1[152].FA_  ( .A(A[664]), .B(n1692), .CI(
        C[664]), .CO(C[665]) );
  FA_12961 \FA_INST_0[1].FA_INST_1[153].FA_  ( .A(A[665]), .B(n1693), .CI(
        C[665]), .CO(C[666]) );
  FA_12960 \FA_INST_0[1].FA_INST_1[154].FA_  ( .A(A[666]), .B(n1694), .CI(
        C[666]), .CO(C[667]) );
  FA_12959 \FA_INST_0[1].FA_INST_1[155].FA_  ( .A(A[667]), .B(n1695), .CI(
        C[667]), .CO(C[668]) );
  FA_12958 \FA_INST_0[1].FA_INST_1[156].FA_  ( .A(A[668]), .B(n1696), .CI(
        C[668]), .CO(C[669]) );
  FA_12957 \FA_INST_0[1].FA_INST_1[157].FA_  ( .A(A[669]), .B(n1697), .CI(
        C[669]), .CO(C[670]) );
  FA_12956 \FA_INST_0[1].FA_INST_1[158].FA_  ( .A(A[670]), .B(n1698), .CI(
        C[670]), .CO(C[671]) );
  FA_12955 \FA_INST_0[1].FA_INST_1[159].FA_  ( .A(A[671]), .B(n1699), .CI(
        C[671]), .CO(C[672]) );
  FA_12954 \FA_INST_0[1].FA_INST_1[160].FA_  ( .A(A[672]), .B(n1700), .CI(
        C[672]), .CO(C[673]) );
  FA_12953 \FA_INST_0[1].FA_INST_1[161].FA_  ( .A(A[673]), .B(n1701), .CI(
        C[673]), .CO(C[674]) );
  FA_12952 \FA_INST_0[1].FA_INST_1[162].FA_  ( .A(A[674]), .B(n1702), .CI(
        C[674]), .CO(C[675]) );
  FA_12951 \FA_INST_0[1].FA_INST_1[163].FA_  ( .A(A[675]), .B(n1703), .CI(
        C[675]), .CO(C[676]) );
  FA_12950 \FA_INST_0[1].FA_INST_1[164].FA_  ( .A(A[676]), .B(n1704), .CI(
        C[676]), .CO(C[677]) );
  FA_12949 \FA_INST_0[1].FA_INST_1[165].FA_  ( .A(A[677]), .B(n1705), .CI(
        C[677]), .CO(C[678]) );
  FA_12948 \FA_INST_0[1].FA_INST_1[166].FA_  ( .A(A[678]), .B(n1706), .CI(
        C[678]), .CO(C[679]) );
  FA_12947 \FA_INST_0[1].FA_INST_1[167].FA_  ( .A(A[679]), .B(n1707), .CI(
        C[679]), .CO(C[680]) );
  FA_12946 \FA_INST_0[1].FA_INST_1[168].FA_  ( .A(A[680]), .B(n1708), .CI(
        C[680]), .CO(C[681]) );
  FA_12945 \FA_INST_0[1].FA_INST_1[169].FA_  ( .A(A[681]), .B(n1709), .CI(
        C[681]), .CO(C[682]) );
  FA_12944 \FA_INST_0[1].FA_INST_1[170].FA_  ( .A(A[682]), .B(n1710), .CI(
        C[682]), .CO(C[683]) );
  FA_12943 \FA_INST_0[1].FA_INST_1[171].FA_  ( .A(A[683]), .B(n1711), .CI(
        C[683]), .CO(C[684]) );
  FA_12942 \FA_INST_0[1].FA_INST_1[172].FA_  ( .A(A[684]), .B(n1712), .CI(
        C[684]), .CO(C[685]) );
  FA_12941 \FA_INST_0[1].FA_INST_1[173].FA_  ( .A(A[685]), .B(n1713), .CI(
        C[685]), .CO(C[686]) );
  FA_12940 \FA_INST_0[1].FA_INST_1[174].FA_  ( .A(A[686]), .B(n1714), .CI(
        C[686]), .CO(C[687]) );
  FA_12939 \FA_INST_0[1].FA_INST_1[175].FA_  ( .A(A[687]), .B(n1715), .CI(
        C[687]), .CO(C[688]) );
  FA_12938 \FA_INST_0[1].FA_INST_1[176].FA_  ( .A(A[688]), .B(n1716), .CI(
        C[688]), .CO(C[689]) );
  FA_12937 \FA_INST_0[1].FA_INST_1[177].FA_  ( .A(A[689]), .B(n1717), .CI(
        C[689]), .CO(C[690]) );
  FA_12936 \FA_INST_0[1].FA_INST_1[178].FA_  ( .A(A[690]), .B(n1718), .CI(
        C[690]), .CO(C[691]) );
  FA_12935 \FA_INST_0[1].FA_INST_1[179].FA_  ( .A(A[691]), .B(n1719), .CI(
        C[691]), .CO(C[692]) );
  FA_12934 \FA_INST_0[1].FA_INST_1[180].FA_  ( .A(A[692]), .B(n1720), .CI(
        C[692]), .CO(C[693]) );
  FA_12933 \FA_INST_0[1].FA_INST_1[181].FA_  ( .A(A[693]), .B(n1721), .CI(
        C[693]), .CO(C[694]) );
  FA_12932 \FA_INST_0[1].FA_INST_1[182].FA_  ( .A(A[694]), .B(n1722), .CI(
        C[694]), .CO(C[695]) );
  FA_12931 \FA_INST_0[1].FA_INST_1[183].FA_  ( .A(A[695]), .B(n1723), .CI(
        C[695]), .CO(C[696]) );
  FA_12930 \FA_INST_0[1].FA_INST_1[184].FA_  ( .A(A[696]), .B(n1724), .CI(
        C[696]), .CO(C[697]) );
  FA_12929 \FA_INST_0[1].FA_INST_1[185].FA_  ( .A(A[697]), .B(n1725), .CI(
        C[697]), .CO(C[698]) );
  FA_12928 \FA_INST_0[1].FA_INST_1[186].FA_  ( .A(A[698]), .B(n1726), .CI(
        C[698]), .CO(C[699]) );
  FA_12927 \FA_INST_0[1].FA_INST_1[187].FA_  ( .A(A[699]), .B(n1727), .CI(
        C[699]), .CO(C[700]) );
  FA_12926 \FA_INST_0[1].FA_INST_1[188].FA_  ( .A(A[700]), .B(n1728), .CI(
        C[700]), .CO(C[701]) );
  FA_12925 \FA_INST_0[1].FA_INST_1[189].FA_  ( .A(A[701]), .B(n1729), .CI(
        C[701]), .CO(C[702]) );
  FA_12924 \FA_INST_0[1].FA_INST_1[190].FA_  ( .A(A[702]), .B(n1730), .CI(
        C[702]), .CO(C[703]) );
  FA_12923 \FA_INST_0[1].FA_INST_1[191].FA_  ( .A(A[703]), .B(n1731), .CI(
        C[703]), .CO(C[704]) );
  FA_12922 \FA_INST_0[1].FA_INST_1[192].FA_  ( .A(A[704]), .B(n1732), .CI(
        C[704]), .CO(C[705]) );
  FA_12921 \FA_INST_0[1].FA_INST_1[193].FA_  ( .A(A[705]), .B(n1733), .CI(
        C[705]), .CO(C[706]) );
  FA_12920 \FA_INST_0[1].FA_INST_1[194].FA_  ( .A(A[706]), .B(n1734), .CI(
        C[706]), .CO(C[707]) );
  FA_12919 \FA_INST_0[1].FA_INST_1[195].FA_  ( .A(A[707]), .B(n1735), .CI(
        C[707]), .CO(C[708]) );
  FA_12918 \FA_INST_0[1].FA_INST_1[196].FA_  ( .A(A[708]), .B(n1736), .CI(
        C[708]), .CO(C[709]) );
  FA_12917 \FA_INST_0[1].FA_INST_1[197].FA_  ( .A(A[709]), .B(n1737), .CI(
        C[709]), .CO(C[710]) );
  FA_12916 \FA_INST_0[1].FA_INST_1[198].FA_  ( .A(A[710]), .B(n1738), .CI(
        C[710]), .CO(C[711]) );
  FA_12915 \FA_INST_0[1].FA_INST_1[199].FA_  ( .A(A[711]), .B(n1739), .CI(
        C[711]), .CO(C[712]) );
  FA_12914 \FA_INST_0[1].FA_INST_1[200].FA_  ( .A(A[712]), .B(n1740), .CI(
        C[712]), .CO(C[713]) );
  FA_12913 \FA_INST_0[1].FA_INST_1[201].FA_  ( .A(A[713]), .B(n1741), .CI(
        C[713]), .CO(C[714]) );
  FA_12912 \FA_INST_0[1].FA_INST_1[202].FA_  ( .A(A[714]), .B(n1742), .CI(
        C[714]), .CO(C[715]) );
  FA_12911 \FA_INST_0[1].FA_INST_1[203].FA_  ( .A(A[715]), .B(n1743), .CI(
        C[715]), .CO(C[716]) );
  FA_12910 \FA_INST_0[1].FA_INST_1[204].FA_  ( .A(A[716]), .B(n1744), .CI(
        C[716]), .CO(C[717]) );
  FA_12909 \FA_INST_0[1].FA_INST_1[205].FA_  ( .A(A[717]), .B(n1745), .CI(
        C[717]), .CO(C[718]) );
  FA_12908 \FA_INST_0[1].FA_INST_1[206].FA_  ( .A(A[718]), .B(n1746), .CI(
        C[718]), .CO(C[719]) );
  FA_12907 \FA_INST_0[1].FA_INST_1[207].FA_  ( .A(A[719]), .B(n1747), .CI(
        C[719]), .CO(C[720]) );
  FA_12906 \FA_INST_0[1].FA_INST_1[208].FA_  ( .A(A[720]), .B(n1748), .CI(
        C[720]), .CO(C[721]) );
  FA_12905 \FA_INST_0[1].FA_INST_1[209].FA_  ( .A(A[721]), .B(n1749), .CI(
        C[721]), .CO(C[722]) );
  FA_12904 \FA_INST_0[1].FA_INST_1[210].FA_  ( .A(A[722]), .B(n1750), .CI(
        C[722]), .CO(C[723]) );
  FA_12903 \FA_INST_0[1].FA_INST_1[211].FA_  ( .A(A[723]), .B(n1751), .CI(
        C[723]), .CO(C[724]) );
  FA_12902 \FA_INST_0[1].FA_INST_1[212].FA_  ( .A(A[724]), .B(n1752), .CI(
        C[724]), .CO(C[725]) );
  FA_12901 \FA_INST_0[1].FA_INST_1[213].FA_  ( .A(A[725]), .B(n1753), .CI(
        C[725]), .CO(C[726]) );
  FA_12900 \FA_INST_0[1].FA_INST_1[214].FA_  ( .A(A[726]), .B(n1754), .CI(
        C[726]), .CO(C[727]) );
  FA_12899 \FA_INST_0[1].FA_INST_1[215].FA_  ( .A(A[727]), .B(n1755), .CI(
        C[727]), .CO(C[728]) );
  FA_12898 \FA_INST_0[1].FA_INST_1[216].FA_  ( .A(A[728]), .B(n1756), .CI(
        C[728]), .CO(C[729]) );
  FA_12897 \FA_INST_0[1].FA_INST_1[217].FA_  ( .A(A[729]), .B(n1757), .CI(
        C[729]), .CO(C[730]) );
  FA_12896 \FA_INST_0[1].FA_INST_1[218].FA_  ( .A(A[730]), .B(n1758), .CI(
        C[730]), .CO(C[731]) );
  FA_12895 \FA_INST_0[1].FA_INST_1[219].FA_  ( .A(A[731]), .B(n1759), .CI(
        C[731]), .CO(C[732]) );
  FA_12894 \FA_INST_0[1].FA_INST_1[220].FA_  ( .A(A[732]), .B(n1760), .CI(
        C[732]), .CO(C[733]) );
  FA_12893 \FA_INST_0[1].FA_INST_1[221].FA_  ( .A(A[733]), .B(n1761), .CI(
        C[733]), .CO(C[734]) );
  FA_12892 \FA_INST_0[1].FA_INST_1[222].FA_  ( .A(A[734]), .B(n1762), .CI(
        C[734]), .CO(C[735]) );
  FA_12891 \FA_INST_0[1].FA_INST_1[223].FA_  ( .A(A[735]), .B(n1763), .CI(
        C[735]), .CO(C[736]) );
  FA_12890 \FA_INST_0[1].FA_INST_1[224].FA_  ( .A(A[736]), .B(n1764), .CI(
        C[736]), .CO(C[737]) );
  FA_12889 \FA_INST_0[1].FA_INST_1[225].FA_  ( .A(A[737]), .B(n1765), .CI(
        C[737]), .CO(C[738]) );
  FA_12888 \FA_INST_0[1].FA_INST_1[226].FA_  ( .A(A[738]), .B(n1766), .CI(
        C[738]), .CO(C[739]) );
  FA_12887 \FA_INST_0[1].FA_INST_1[227].FA_  ( .A(A[739]), .B(n1767), .CI(
        C[739]), .CO(C[740]) );
  FA_12886 \FA_INST_0[1].FA_INST_1[228].FA_  ( .A(A[740]), .B(n1768), .CI(
        C[740]), .CO(C[741]) );
  FA_12885 \FA_INST_0[1].FA_INST_1[229].FA_  ( .A(A[741]), .B(n1769), .CI(
        C[741]), .CO(C[742]) );
  FA_12884 \FA_INST_0[1].FA_INST_1[230].FA_  ( .A(A[742]), .B(n1770), .CI(
        C[742]), .CO(C[743]) );
  FA_12883 \FA_INST_0[1].FA_INST_1[231].FA_  ( .A(A[743]), .B(n1771), .CI(
        C[743]), .CO(C[744]) );
  FA_12882 \FA_INST_0[1].FA_INST_1[232].FA_  ( .A(A[744]), .B(n1772), .CI(
        C[744]), .CO(C[745]) );
  FA_12881 \FA_INST_0[1].FA_INST_1[233].FA_  ( .A(A[745]), .B(n1773), .CI(
        C[745]), .CO(C[746]) );
  FA_12880 \FA_INST_0[1].FA_INST_1[234].FA_  ( .A(A[746]), .B(n1774), .CI(
        C[746]), .CO(C[747]) );
  FA_12879 \FA_INST_0[1].FA_INST_1[235].FA_  ( .A(A[747]), .B(n1775), .CI(
        C[747]), .CO(C[748]) );
  FA_12878 \FA_INST_0[1].FA_INST_1[236].FA_  ( .A(A[748]), .B(n1776), .CI(
        C[748]), .CO(C[749]) );
  FA_12877 \FA_INST_0[1].FA_INST_1[237].FA_  ( .A(A[749]), .B(n1777), .CI(
        C[749]), .CO(C[750]) );
  FA_12876 \FA_INST_0[1].FA_INST_1[238].FA_  ( .A(A[750]), .B(n1778), .CI(
        C[750]), .CO(C[751]) );
  FA_12875 \FA_INST_0[1].FA_INST_1[239].FA_  ( .A(A[751]), .B(n1779), .CI(
        C[751]), .CO(C[752]) );
  FA_12874 \FA_INST_0[1].FA_INST_1[240].FA_  ( .A(A[752]), .B(n1780), .CI(
        C[752]), .CO(C[753]) );
  FA_12873 \FA_INST_0[1].FA_INST_1[241].FA_  ( .A(A[753]), .B(n1781), .CI(
        C[753]), .CO(C[754]) );
  FA_12872 \FA_INST_0[1].FA_INST_1[242].FA_  ( .A(A[754]), .B(n1782), .CI(
        C[754]), .CO(C[755]) );
  FA_12871 \FA_INST_0[1].FA_INST_1[243].FA_  ( .A(A[755]), .B(n1783), .CI(
        C[755]), .CO(C[756]) );
  FA_12870 \FA_INST_0[1].FA_INST_1[244].FA_  ( .A(A[756]), .B(n1784), .CI(
        C[756]), .CO(C[757]) );
  FA_12869 \FA_INST_0[1].FA_INST_1[245].FA_  ( .A(A[757]), .B(n1785), .CI(
        C[757]), .CO(C[758]) );
  FA_12868 \FA_INST_0[1].FA_INST_1[246].FA_  ( .A(A[758]), .B(n1786), .CI(
        C[758]), .CO(C[759]) );
  FA_12867 \FA_INST_0[1].FA_INST_1[247].FA_  ( .A(A[759]), .B(n1787), .CI(
        C[759]), .CO(C[760]) );
  FA_12866 \FA_INST_0[1].FA_INST_1[248].FA_  ( .A(A[760]), .B(n1788), .CI(
        C[760]), .CO(C[761]) );
  FA_12865 \FA_INST_0[1].FA_INST_1[249].FA_  ( .A(A[761]), .B(n1789), .CI(
        C[761]), .CO(C[762]) );
  FA_12864 \FA_INST_0[1].FA_INST_1[250].FA_  ( .A(A[762]), .B(n1790), .CI(
        C[762]), .CO(C[763]) );
  FA_12863 \FA_INST_0[1].FA_INST_1[251].FA_  ( .A(A[763]), .B(n1791), .CI(
        C[763]), .CO(C[764]) );
  FA_12862 \FA_INST_0[1].FA_INST_1[252].FA_  ( .A(A[764]), .B(n1792), .CI(
        C[764]), .CO(C[765]) );
  FA_12861 \FA_INST_0[1].FA_INST_1[253].FA_  ( .A(A[765]), .B(n1793), .CI(
        C[765]), .CO(C[766]) );
  FA_12860 \FA_INST_0[1].FA_INST_1[254].FA_  ( .A(A[766]), .B(n1794), .CI(
        C[766]), .CO(C[767]) );
  FA_12859 \FA_INST_0[1].FA_INST_1[255].FA_  ( .A(A[767]), .B(n1795), .CI(
        C[767]), .CO(C[768]) );
  FA_12858 \FA_INST_0[1].FA_INST_1[256].FA_  ( .A(A[768]), .B(n1796), .CI(
        C[768]), .CO(C[769]) );
  FA_12857 \FA_INST_0[1].FA_INST_1[257].FA_  ( .A(A[769]), .B(n1797), .CI(
        C[769]), .CO(C[770]) );
  FA_12856 \FA_INST_0[1].FA_INST_1[258].FA_  ( .A(A[770]), .B(n1798), .CI(
        C[770]), .CO(C[771]) );
  FA_12855 \FA_INST_0[1].FA_INST_1[259].FA_  ( .A(A[771]), .B(n1799), .CI(
        C[771]), .CO(C[772]) );
  FA_12854 \FA_INST_0[1].FA_INST_1[260].FA_  ( .A(A[772]), .B(n1800), .CI(
        C[772]), .CO(C[773]) );
  FA_12853 \FA_INST_0[1].FA_INST_1[261].FA_  ( .A(A[773]), .B(n1801), .CI(
        C[773]), .CO(C[774]) );
  FA_12852 \FA_INST_0[1].FA_INST_1[262].FA_  ( .A(A[774]), .B(n1802), .CI(
        C[774]), .CO(C[775]) );
  FA_12851 \FA_INST_0[1].FA_INST_1[263].FA_  ( .A(A[775]), .B(n1803), .CI(
        C[775]), .CO(C[776]) );
  FA_12850 \FA_INST_0[1].FA_INST_1[264].FA_  ( .A(A[776]), .B(n1804), .CI(
        C[776]), .CO(C[777]) );
  FA_12849 \FA_INST_0[1].FA_INST_1[265].FA_  ( .A(A[777]), .B(n1805), .CI(
        C[777]), .CO(C[778]) );
  FA_12848 \FA_INST_0[1].FA_INST_1[266].FA_  ( .A(A[778]), .B(n1806), .CI(
        C[778]), .CO(C[779]) );
  FA_12847 \FA_INST_0[1].FA_INST_1[267].FA_  ( .A(A[779]), .B(n1807), .CI(
        C[779]), .CO(C[780]) );
  FA_12846 \FA_INST_0[1].FA_INST_1[268].FA_  ( .A(A[780]), .B(n1808), .CI(
        C[780]), .CO(C[781]) );
  FA_12845 \FA_INST_0[1].FA_INST_1[269].FA_  ( .A(A[781]), .B(n1809), .CI(
        C[781]), .CO(C[782]) );
  FA_12844 \FA_INST_0[1].FA_INST_1[270].FA_  ( .A(A[782]), .B(n1810), .CI(
        C[782]), .CO(C[783]) );
  FA_12843 \FA_INST_0[1].FA_INST_1[271].FA_  ( .A(A[783]), .B(n1811), .CI(
        C[783]), .CO(C[784]) );
  FA_12842 \FA_INST_0[1].FA_INST_1[272].FA_  ( .A(A[784]), .B(n1812), .CI(
        C[784]), .CO(C[785]) );
  FA_12841 \FA_INST_0[1].FA_INST_1[273].FA_  ( .A(A[785]), .B(n1813), .CI(
        C[785]), .CO(C[786]) );
  FA_12840 \FA_INST_0[1].FA_INST_1[274].FA_  ( .A(A[786]), .B(n1814), .CI(
        C[786]), .CO(C[787]) );
  FA_12839 \FA_INST_0[1].FA_INST_1[275].FA_  ( .A(A[787]), .B(n1815), .CI(
        C[787]), .CO(C[788]) );
  FA_12838 \FA_INST_0[1].FA_INST_1[276].FA_  ( .A(A[788]), .B(n1816), .CI(
        C[788]), .CO(C[789]) );
  FA_12837 \FA_INST_0[1].FA_INST_1[277].FA_  ( .A(A[789]), .B(n1817), .CI(
        C[789]), .CO(C[790]) );
  FA_12836 \FA_INST_0[1].FA_INST_1[278].FA_  ( .A(A[790]), .B(n1818), .CI(
        C[790]), .CO(C[791]) );
  FA_12835 \FA_INST_0[1].FA_INST_1[279].FA_  ( .A(A[791]), .B(n1819), .CI(
        C[791]), .CO(C[792]) );
  FA_12834 \FA_INST_0[1].FA_INST_1[280].FA_  ( .A(A[792]), .B(n1820), .CI(
        C[792]), .CO(C[793]) );
  FA_12833 \FA_INST_0[1].FA_INST_1[281].FA_  ( .A(A[793]), .B(n1821), .CI(
        C[793]), .CO(C[794]) );
  FA_12832 \FA_INST_0[1].FA_INST_1[282].FA_  ( .A(A[794]), .B(n1822), .CI(
        C[794]), .CO(C[795]) );
  FA_12831 \FA_INST_0[1].FA_INST_1[283].FA_  ( .A(A[795]), .B(n1823), .CI(
        C[795]), .CO(C[796]) );
  FA_12830 \FA_INST_0[1].FA_INST_1[284].FA_  ( .A(A[796]), .B(n1824), .CI(
        C[796]), .CO(C[797]) );
  FA_12829 \FA_INST_0[1].FA_INST_1[285].FA_  ( .A(A[797]), .B(n1825), .CI(
        C[797]), .CO(C[798]) );
  FA_12828 \FA_INST_0[1].FA_INST_1[286].FA_  ( .A(A[798]), .B(n1826), .CI(
        C[798]), .CO(C[799]) );
  FA_12827 \FA_INST_0[1].FA_INST_1[287].FA_  ( .A(A[799]), .B(n1827), .CI(
        C[799]), .CO(C[800]) );
  FA_12826 \FA_INST_0[1].FA_INST_1[288].FA_  ( .A(A[800]), .B(n1828), .CI(
        C[800]), .CO(C[801]) );
  FA_12825 \FA_INST_0[1].FA_INST_1[289].FA_  ( .A(A[801]), .B(n1829), .CI(
        C[801]), .CO(C[802]) );
  FA_12824 \FA_INST_0[1].FA_INST_1[290].FA_  ( .A(A[802]), .B(n1830), .CI(
        C[802]), .CO(C[803]) );
  FA_12823 \FA_INST_0[1].FA_INST_1[291].FA_  ( .A(A[803]), .B(n1831), .CI(
        C[803]), .CO(C[804]) );
  FA_12822 \FA_INST_0[1].FA_INST_1[292].FA_  ( .A(A[804]), .B(n1832), .CI(
        C[804]), .CO(C[805]) );
  FA_12821 \FA_INST_0[1].FA_INST_1[293].FA_  ( .A(A[805]), .B(n1833), .CI(
        C[805]), .CO(C[806]) );
  FA_12820 \FA_INST_0[1].FA_INST_1[294].FA_  ( .A(A[806]), .B(n1834), .CI(
        C[806]), .CO(C[807]) );
  FA_12819 \FA_INST_0[1].FA_INST_1[295].FA_  ( .A(A[807]), .B(n1835), .CI(
        C[807]), .CO(C[808]) );
  FA_12818 \FA_INST_0[1].FA_INST_1[296].FA_  ( .A(A[808]), .B(n1836), .CI(
        C[808]), .CO(C[809]) );
  FA_12817 \FA_INST_0[1].FA_INST_1[297].FA_  ( .A(A[809]), .B(n1837), .CI(
        C[809]), .CO(C[810]) );
  FA_12816 \FA_INST_0[1].FA_INST_1[298].FA_  ( .A(A[810]), .B(n1838), .CI(
        C[810]), .CO(C[811]) );
  FA_12815 \FA_INST_0[1].FA_INST_1[299].FA_  ( .A(A[811]), .B(n1839), .CI(
        C[811]), .CO(C[812]) );
  FA_12814 \FA_INST_0[1].FA_INST_1[300].FA_  ( .A(A[812]), .B(n1840), .CI(
        C[812]), .CO(C[813]) );
  FA_12813 \FA_INST_0[1].FA_INST_1[301].FA_  ( .A(A[813]), .B(n1841), .CI(
        C[813]), .CO(C[814]) );
  FA_12812 \FA_INST_0[1].FA_INST_1[302].FA_  ( .A(A[814]), .B(n1842), .CI(
        C[814]), .CO(C[815]) );
  FA_12811 \FA_INST_0[1].FA_INST_1[303].FA_  ( .A(A[815]), .B(n1843), .CI(
        C[815]), .CO(C[816]) );
  FA_12810 \FA_INST_0[1].FA_INST_1[304].FA_  ( .A(A[816]), .B(n1844), .CI(
        C[816]), .CO(C[817]) );
  FA_12809 \FA_INST_0[1].FA_INST_1[305].FA_  ( .A(A[817]), .B(n1845), .CI(
        C[817]), .CO(C[818]) );
  FA_12808 \FA_INST_0[1].FA_INST_1[306].FA_  ( .A(A[818]), .B(n1846), .CI(
        C[818]), .CO(C[819]) );
  FA_12807 \FA_INST_0[1].FA_INST_1[307].FA_  ( .A(A[819]), .B(n1847), .CI(
        C[819]), .CO(C[820]) );
  FA_12806 \FA_INST_0[1].FA_INST_1[308].FA_  ( .A(A[820]), .B(n1848), .CI(
        C[820]), .CO(C[821]) );
  FA_12805 \FA_INST_0[1].FA_INST_1[309].FA_  ( .A(A[821]), .B(n1849), .CI(
        C[821]), .CO(C[822]) );
  FA_12804 \FA_INST_0[1].FA_INST_1[310].FA_  ( .A(A[822]), .B(n1850), .CI(
        C[822]), .CO(C[823]) );
  FA_12803 \FA_INST_0[1].FA_INST_1[311].FA_  ( .A(A[823]), .B(n1851), .CI(
        C[823]), .CO(C[824]) );
  FA_12802 \FA_INST_0[1].FA_INST_1[312].FA_  ( .A(A[824]), .B(n1852), .CI(
        C[824]), .CO(C[825]) );
  FA_12801 \FA_INST_0[1].FA_INST_1[313].FA_  ( .A(A[825]), .B(n1853), .CI(
        C[825]), .CO(C[826]) );
  FA_12800 \FA_INST_0[1].FA_INST_1[314].FA_  ( .A(A[826]), .B(n1854), .CI(
        C[826]), .CO(C[827]) );
  FA_12799 \FA_INST_0[1].FA_INST_1[315].FA_  ( .A(A[827]), .B(n1855), .CI(
        C[827]), .CO(C[828]) );
  FA_12798 \FA_INST_0[1].FA_INST_1[316].FA_  ( .A(A[828]), .B(n1856), .CI(
        C[828]), .CO(C[829]) );
  FA_12797 \FA_INST_0[1].FA_INST_1[317].FA_  ( .A(A[829]), .B(n1857), .CI(
        C[829]), .CO(C[830]) );
  FA_12796 \FA_INST_0[1].FA_INST_1[318].FA_  ( .A(A[830]), .B(n1858), .CI(
        C[830]), .CO(C[831]) );
  FA_12795 \FA_INST_0[1].FA_INST_1[319].FA_  ( .A(A[831]), .B(n1859), .CI(
        C[831]), .CO(C[832]) );
  FA_12794 \FA_INST_0[1].FA_INST_1[320].FA_  ( .A(A[832]), .B(n1860), .CI(
        C[832]), .CO(C[833]) );
  FA_12793 \FA_INST_0[1].FA_INST_1[321].FA_  ( .A(A[833]), .B(n1861), .CI(
        C[833]), .CO(C[834]) );
  FA_12792 \FA_INST_0[1].FA_INST_1[322].FA_  ( .A(A[834]), .B(n1862), .CI(
        C[834]), .CO(C[835]) );
  FA_12791 \FA_INST_0[1].FA_INST_1[323].FA_  ( .A(A[835]), .B(n1863), .CI(
        C[835]), .CO(C[836]) );
  FA_12790 \FA_INST_0[1].FA_INST_1[324].FA_  ( .A(A[836]), .B(n1864), .CI(
        C[836]), .CO(C[837]) );
  FA_12789 \FA_INST_0[1].FA_INST_1[325].FA_  ( .A(A[837]), .B(n1865), .CI(
        C[837]), .CO(C[838]) );
  FA_12788 \FA_INST_0[1].FA_INST_1[326].FA_  ( .A(A[838]), .B(n1866), .CI(
        C[838]), .CO(C[839]) );
  FA_12787 \FA_INST_0[1].FA_INST_1[327].FA_  ( .A(A[839]), .B(n1867), .CI(
        C[839]), .CO(C[840]) );
  FA_12786 \FA_INST_0[1].FA_INST_1[328].FA_  ( .A(A[840]), .B(n1868), .CI(
        C[840]), .CO(C[841]) );
  FA_12785 \FA_INST_0[1].FA_INST_1[329].FA_  ( .A(A[841]), .B(n1869), .CI(
        C[841]), .CO(C[842]) );
  FA_12784 \FA_INST_0[1].FA_INST_1[330].FA_  ( .A(A[842]), .B(n1870), .CI(
        C[842]), .CO(C[843]) );
  FA_12783 \FA_INST_0[1].FA_INST_1[331].FA_  ( .A(A[843]), .B(n1871), .CI(
        C[843]), .CO(C[844]) );
  FA_12782 \FA_INST_0[1].FA_INST_1[332].FA_  ( .A(A[844]), .B(n1872), .CI(
        C[844]), .CO(C[845]) );
  FA_12781 \FA_INST_0[1].FA_INST_1[333].FA_  ( .A(A[845]), .B(n1873), .CI(
        C[845]), .CO(C[846]) );
  FA_12780 \FA_INST_0[1].FA_INST_1[334].FA_  ( .A(A[846]), .B(n1874), .CI(
        C[846]), .CO(C[847]) );
  FA_12779 \FA_INST_0[1].FA_INST_1[335].FA_  ( .A(A[847]), .B(n1875), .CI(
        C[847]), .CO(C[848]) );
  FA_12778 \FA_INST_0[1].FA_INST_1[336].FA_  ( .A(A[848]), .B(n1876), .CI(
        C[848]), .CO(C[849]) );
  FA_12777 \FA_INST_0[1].FA_INST_1[337].FA_  ( .A(A[849]), .B(n1877), .CI(
        C[849]), .CO(C[850]) );
  FA_12776 \FA_INST_0[1].FA_INST_1[338].FA_  ( .A(A[850]), .B(n1878), .CI(
        C[850]), .CO(C[851]) );
  FA_12775 \FA_INST_0[1].FA_INST_1[339].FA_  ( .A(A[851]), .B(n1879), .CI(
        C[851]), .CO(C[852]) );
  FA_12774 \FA_INST_0[1].FA_INST_1[340].FA_  ( .A(A[852]), .B(n1880), .CI(
        C[852]), .CO(C[853]) );
  FA_12773 \FA_INST_0[1].FA_INST_1[341].FA_  ( .A(A[853]), .B(n1881), .CI(
        C[853]), .CO(C[854]) );
  FA_12772 \FA_INST_0[1].FA_INST_1[342].FA_  ( .A(A[854]), .B(n1882), .CI(
        C[854]), .CO(C[855]) );
  FA_12771 \FA_INST_0[1].FA_INST_1[343].FA_  ( .A(A[855]), .B(n1883), .CI(
        C[855]), .CO(C[856]) );
  FA_12770 \FA_INST_0[1].FA_INST_1[344].FA_  ( .A(A[856]), .B(n1884), .CI(
        C[856]), .CO(C[857]) );
  FA_12769 \FA_INST_0[1].FA_INST_1[345].FA_  ( .A(A[857]), .B(n1885), .CI(
        C[857]), .CO(C[858]) );
  FA_12768 \FA_INST_0[1].FA_INST_1[346].FA_  ( .A(A[858]), .B(n1886), .CI(
        C[858]), .CO(C[859]) );
  FA_12767 \FA_INST_0[1].FA_INST_1[347].FA_  ( .A(A[859]), .B(n1887), .CI(
        C[859]), .CO(C[860]) );
  FA_12766 \FA_INST_0[1].FA_INST_1[348].FA_  ( .A(A[860]), .B(n1888), .CI(
        C[860]), .CO(C[861]) );
  FA_12765 \FA_INST_0[1].FA_INST_1[349].FA_  ( .A(A[861]), .B(n1889), .CI(
        C[861]), .CO(C[862]) );
  FA_12764 \FA_INST_0[1].FA_INST_1[350].FA_  ( .A(A[862]), .B(n1890), .CI(
        C[862]), .CO(C[863]) );
  FA_12763 \FA_INST_0[1].FA_INST_1[351].FA_  ( .A(A[863]), .B(n1891), .CI(
        C[863]), .CO(C[864]) );
  FA_12762 \FA_INST_0[1].FA_INST_1[352].FA_  ( .A(A[864]), .B(n1892), .CI(
        C[864]), .CO(C[865]) );
  FA_12761 \FA_INST_0[1].FA_INST_1[353].FA_  ( .A(A[865]), .B(n1893), .CI(
        C[865]), .CO(C[866]) );
  FA_12760 \FA_INST_0[1].FA_INST_1[354].FA_  ( .A(A[866]), .B(n1894), .CI(
        C[866]), .CO(C[867]) );
  FA_12759 \FA_INST_0[1].FA_INST_1[355].FA_  ( .A(A[867]), .B(n1895), .CI(
        C[867]), .CO(C[868]) );
  FA_12758 \FA_INST_0[1].FA_INST_1[356].FA_  ( .A(A[868]), .B(n1896), .CI(
        C[868]), .CO(C[869]) );
  FA_12757 \FA_INST_0[1].FA_INST_1[357].FA_  ( .A(A[869]), .B(n1897), .CI(
        C[869]), .CO(C[870]) );
  FA_12756 \FA_INST_0[1].FA_INST_1[358].FA_  ( .A(A[870]), .B(n1898), .CI(
        C[870]), .CO(C[871]) );
  FA_12755 \FA_INST_0[1].FA_INST_1[359].FA_  ( .A(A[871]), .B(n1899), .CI(
        C[871]), .CO(C[872]) );
  FA_12754 \FA_INST_0[1].FA_INST_1[360].FA_  ( .A(A[872]), .B(n1900), .CI(
        C[872]), .CO(C[873]) );
  FA_12753 \FA_INST_0[1].FA_INST_1[361].FA_  ( .A(A[873]), .B(n1901), .CI(
        C[873]), .CO(C[874]) );
  FA_12752 \FA_INST_0[1].FA_INST_1[362].FA_  ( .A(A[874]), .B(n1902), .CI(
        C[874]), .CO(C[875]) );
  FA_12751 \FA_INST_0[1].FA_INST_1[363].FA_  ( .A(A[875]), .B(n1903), .CI(
        C[875]), .CO(C[876]) );
  FA_12750 \FA_INST_0[1].FA_INST_1[364].FA_  ( .A(A[876]), .B(n1904), .CI(
        C[876]), .CO(C[877]) );
  FA_12749 \FA_INST_0[1].FA_INST_1[365].FA_  ( .A(A[877]), .B(n1905), .CI(
        C[877]), .CO(C[878]) );
  FA_12748 \FA_INST_0[1].FA_INST_1[366].FA_  ( .A(A[878]), .B(n1906), .CI(
        C[878]), .CO(C[879]) );
  FA_12747 \FA_INST_0[1].FA_INST_1[367].FA_  ( .A(A[879]), .B(n1907), .CI(
        C[879]), .CO(C[880]) );
  FA_12746 \FA_INST_0[1].FA_INST_1[368].FA_  ( .A(A[880]), .B(n1908), .CI(
        C[880]), .CO(C[881]) );
  FA_12745 \FA_INST_0[1].FA_INST_1[369].FA_  ( .A(A[881]), .B(n1909), .CI(
        C[881]), .CO(C[882]) );
  FA_12744 \FA_INST_0[1].FA_INST_1[370].FA_  ( .A(A[882]), .B(n1910), .CI(
        C[882]), .CO(C[883]) );
  FA_12743 \FA_INST_0[1].FA_INST_1[371].FA_  ( .A(A[883]), .B(n1911), .CI(
        C[883]), .CO(C[884]) );
  FA_12742 \FA_INST_0[1].FA_INST_1[372].FA_  ( .A(A[884]), .B(n1912), .CI(
        C[884]), .CO(C[885]) );
  FA_12741 \FA_INST_0[1].FA_INST_1[373].FA_  ( .A(A[885]), .B(n1913), .CI(
        C[885]), .CO(C[886]) );
  FA_12740 \FA_INST_0[1].FA_INST_1[374].FA_  ( .A(A[886]), .B(n1914), .CI(
        C[886]), .CO(C[887]) );
  FA_12739 \FA_INST_0[1].FA_INST_1[375].FA_  ( .A(A[887]), .B(n1915), .CI(
        C[887]), .CO(C[888]) );
  FA_12738 \FA_INST_0[1].FA_INST_1[376].FA_  ( .A(A[888]), .B(n1916), .CI(
        C[888]), .CO(C[889]) );
  FA_12737 \FA_INST_0[1].FA_INST_1[377].FA_  ( .A(A[889]), .B(n1917), .CI(
        C[889]), .CO(C[890]) );
  FA_12736 \FA_INST_0[1].FA_INST_1[378].FA_  ( .A(A[890]), .B(n1918), .CI(
        C[890]), .CO(C[891]) );
  FA_12735 \FA_INST_0[1].FA_INST_1[379].FA_  ( .A(A[891]), .B(n1919), .CI(
        C[891]), .CO(C[892]) );
  FA_12734 \FA_INST_0[1].FA_INST_1[380].FA_  ( .A(A[892]), .B(n1920), .CI(
        C[892]), .CO(C[893]) );
  FA_12733 \FA_INST_0[1].FA_INST_1[381].FA_  ( .A(A[893]), .B(n1921), .CI(
        C[893]), .CO(C[894]) );
  FA_12732 \FA_INST_0[1].FA_INST_1[382].FA_  ( .A(A[894]), .B(n1922), .CI(
        C[894]), .CO(C[895]) );
  FA_12731 \FA_INST_0[1].FA_INST_1[383].FA_  ( .A(A[895]), .B(n1923), .CI(
        C[895]), .CO(C[896]) );
  FA_12730 \FA_INST_0[1].FA_INST_1[384].FA_  ( .A(A[896]), .B(n1924), .CI(
        C[896]), .CO(C[897]) );
  FA_12729 \FA_INST_0[1].FA_INST_1[385].FA_  ( .A(A[897]), .B(n1925), .CI(
        C[897]), .CO(C[898]) );
  FA_12728 \FA_INST_0[1].FA_INST_1[386].FA_  ( .A(A[898]), .B(n1926), .CI(
        C[898]), .CO(C[899]) );
  FA_12727 \FA_INST_0[1].FA_INST_1[387].FA_  ( .A(A[899]), .B(n1927), .CI(
        C[899]), .CO(C[900]) );
  FA_12726 \FA_INST_0[1].FA_INST_1[388].FA_  ( .A(A[900]), .B(n1928), .CI(
        C[900]), .CO(C[901]) );
  FA_12725 \FA_INST_0[1].FA_INST_1[389].FA_  ( .A(A[901]), .B(n1929), .CI(
        C[901]), .CO(C[902]) );
  FA_12724 \FA_INST_0[1].FA_INST_1[390].FA_  ( .A(A[902]), .B(n1930), .CI(
        C[902]), .CO(C[903]) );
  FA_12723 \FA_INST_0[1].FA_INST_1[391].FA_  ( .A(A[903]), .B(n1931), .CI(
        C[903]), .CO(C[904]) );
  FA_12722 \FA_INST_0[1].FA_INST_1[392].FA_  ( .A(A[904]), .B(n1932), .CI(
        C[904]), .CO(C[905]) );
  FA_12721 \FA_INST_0[1].FA_INST_1[393].FA_  ( .A(A[905]), .B(n1933), .CI(
        C[905]), .CO(C[906]) );
  FA_12720 \FA_INST_0[1].FA_INST_1[394].FA_  ( .A(A[906]), .B(n1934), .CI(
        C[906]), .CO(C[907]) );
  FA_12719 \FA_INST_0[1].FA_INST_1[395].FA_  ( .A(A[907]), .B(n1935), .CI(
        C[907]), .CO(C[908]) );
  FA_12718 \FA_INST_0[1].FA_INST_1[396].FA_  ( .A(A[908]), .B(n1936), .CI(
        C[908]), .CO(C[909]) );
  FA_12717 \FA_INST_0[1].FA_INST_1[397].FA_  ( .A(A[909]), .B(n1937), .CI(
        C[909]), .CO(C[910]) );
  FA_12716 \FA_INST_0[1].FA_INST_1[398].FA_  ( .A(A[910]), .B(n1938), .CI(
        C[910]), .CO(C[911]) );
  FA_12715 \FA_INST_0[1].FA_INST_1[399].FA_  ( .A(A[911]), .B(n1939), .CI(
        C[911]), .CO(C[912]) );
  FA_12714 \FA_INST_0[1].FA_INST_1[400].FA_  ( .A(A[912]), .B(n1940), .CI(
        C[912]), .CO(C[913]) );
  FA_12713 \FA_INST_0[1].FA_INST_1[401].FA_  ( .A(A[913]), .B(n1941), .CI(
        C[913]), .CO(C[914]) );
  FA_12712 \FA_INST_0[1].FA_INST_1[402].FA_  ( .A(A[914]), .B(n1942), .CI(
        C[914]), .CO(C[915]) );
  FA_12711 \FA_INST_0[1].FA_INST_1[403].FA_  ( .A(A[915]), .B(n1943), .CI(
        C[915]), .CO(C[916]) );
  FA_12710 \FA_INST_0[1].FA_INST_1[404].FA_  ( .A(A[916]), .B(n1944), .CI(
        C[916]), .CO(C[917]) );
  FA_12709 \FA_INST_0[1].FA_INST_1[405].FA_  ( .A(A[917]), .B(n1945), .CI(
        C[917]), .CO(C[918]) );
  FA_12708 \FA_INST_0[1].FA_INST_1[406].FA_  ( .A(A[918]), .B(n1946), .CI(
        C[918]), .CO(C[919]) );
  FA_12707 \FA_INST_0[1].FA_INST_1[407].FA_  ( .A(A[919]), .B(n1947), .CI(
        C[919]), .CO(C[920]) );
  FA_12706 \FA_INST_0[1].FA_INST_1[408].FA_  ( .A(A[920]), .B(n1948), .CI(
        C[920]), .CO(C[921]) );
  FA_12705 \FA_INST_0[1].FA_INST_1[409].FA_  ( .A(A[921]), .B(n1949), .CI(
        C[921]), .CO(C[922]) );
  FA_12704 \FA_INST_0[1].FA_INST_1[410].FA_  ( .A(A[922]), .B(n1950), .CI(
        C[922]), .CO(C[923]) );
  FA_12703 \FA_INST_0[1].FA_INST_1[411].FA_  ( .A(A[923]), .B(n1951), .CI(
        C[923]), .CO(C[924]) );
  FA_12702 \FA_INST_0[1].FA_INST_1[412].FA_  ( .A(A[924]), .B(n1952), .CI(
        C[924]), .CO(C[925]) );
  FA_12701 \FA_INST_0[1].FA_INST_1[413].FA_  ( .A(A[925]), .B(n1953), .CI(
        C[925]), .CO(C[926]) );
  FA_12700 \FA_INST_0[1].FA_INST_1[414].FA_  ( .A(A[926]), .B(n1954), .CI(
        C[926]), .CO(C[927]) );
  FA_12699 \FA_INST_0[1].FA_INST_1[415].FA_  ( .A(A[927]), .B(n1955), .CI(
        C[927]), .CO(C[928]) );
  FA_12698 \FA_INST_0[1].FA_INST_1[416].FA_  ( .A(A[928]), .B(n1956), .CI(
        C[928]), .CO(C[929]) );
  FA_12697 \FA_INST_0[1].FA_INST_1[417].FA_  ( .A(A[929]), .B(n1957), .CI(
        C[929]), .CO(C[930]) );
  FA_12696 \FA_INST_0[1].FA_INST_1[418].FA_  ( .A(A[930]), .B(n1958), .CI(
        C[930]), .CO(C[931]) );
  FA_12695 \FA_INST_0[1].FA_INST_1[419].FA_  ( .A(A[931]), .B(n1959), .CI(
        C[931]), .CO(C[932]) );
  FA_12694 \FA_INST_0[1].FA_INST_1[420].FA_  ( .A(A[932]), .B(n1960), .CI(
        C[932]), .CO(C[933]) );
  FA_12693 \FA_INST_0[1].FA_INST_1[421].FA_  ( .A(A[933]), .B(n1961), .CI(
        C[933]), .CO(C[934]) );
  FA_12692 \FA_INST_0[1].FA_INST_1[422].FA_  ( .A(A[934]), .B(n1962), .CI(
        C[934]), .CO(C[935]) );
  FA_12691 \FA_INST_0[1].FA_INST_1[423].FA_  ( .A(A[935]), .B(n1963), .CI(
        C[935]), .CO(C[936]) );
  FA_12690 \FA_INST_0[1].FA_INST_1[424].FA_  ( .A(A[936]), .B(n1964), .CI(
        C[936]), .CO(C[937]) );
  FA_12689 \FA_INST_0[1].FA_INST_1[425].FA_  ( .A(A[937]), .B(n1965), .CI(
        C[937]), .CO(C[938]) );
  FA_12688 \FA_INST_0[1].FA_INST_1[426].FA_  ( .A(A[938]), .B(n1966), .CI(
        C[938]), .CO(C[939]) );
  FA_12687 \FA_INST_0[1].FA_INST_1[427].FA_  ( .A(A[939]), .B(n1967), .CI(
        C[939]), .CO(C[940]) );
  FA_12686 \FA_INST_0[1].FA_INST_1[428].FA_  ( .A(A[940]), .B(n1968), .CI(
        C[940]), .CO(C[941]) );
  FA_12685 \FA_INST_0[1].FA_INST_1[429].FA_  ( .A(A[941]), .B(n1969), .CI(
        C[941]), .CO(C[942]) );
  FA_12684 \FA_INST_0[1].FA_INST_1[430].FA_  ( .A(A[942]), .B(n1970), .CI(
        C[942]), .CO(C[943]) );
  FA_12683 \FA_INST_0[1].FA_INST_1[431].FA_  ( .A(A[943]), .B(n1971), .CI(
        C[943]), .CO(C[944]) );
  FA_12682 \FA_INST_0[1].FA_INST_1[432].FA_  ( .A(A[944]), .B(n1972), .CI(
        C[944]), .CO(C[945]) );
  FA_12681 \FA_INST_0[1].FA_INST_1[433].FA_  ( .A(A[945]), .B(n1973), .CI(
        C[945]), .CO(C[946]) );
  FA_12680 \FA_INST_0[1].FA_INST_1[434].FA_  ( .A(A[946]), .B(n1974), .CI(
        C[946]), .CO(C[947]) );
  FA_12679 \FA_INST_0[1].FA_INST_1[435].FA_  ( .A(A[947]), .B(n1975), .CI(
        C[947]), .CO(C[948]) );
  FA_12678 \FA_INST_0[1].FA_INST_1[436].FA_  ( .A(A[948]), .B(n1976), .CI(
        C[948]), .CO(C[949]) );
  FA_12677 \FA_INST_0[1].FA_INST_1[437].FA_  ( .A(A[949]), .B(n1977), .CI(
        C[949]), .CO(C[950]) );
  FA_12676 \FA_INST_0[1].FA_INST_1[438].FA_  ( .A(A[950]), .B(n1978), .CI(
        C[950]), .CO(C[951]) );
  FA_12675 \FA_INST_0[1].FA_INST_1[439].FA_  ( .A(A[951]), .B(n1979), .CI(
        C[951]), .CO(C[952]) );
  FA_12674 \FA_INST_0[1].FA_INST_1[440].FA_  ( .A(A[952]), .B(n1980), .CI(
        C[952]), .CO(C[953]) );
  FA_12673 \FA_INST_0[1].FA_INST_1[441].FA_  ( .A(A[953]), .B(n1981), .CI(
        C[953]), .CO(C[954]) );
  FA_12672 \FA_INST_0[1].FA_INST_1[442].FA_  ( .A(A[954]), .B(n1982), .CI(
        C[954]), .CO(C[955]) );
  FA_12671 \FA_INST_0[1].FA_INST_1[443].FA_  ( .A(A[955]), .B(n1983), .CI(
        C[955]), .CO(C[956]) );
  FA_12670 \FA_INST_0[1].FA_INST_1[444].FA_  ( .A(A[956]), .B(n1984), .CI(
        C[956]), .CO(C[957]) );
  FA_12669 \FA_INST_0[1].FA_INST_1[445].FA_  ( .A(A[957]), .B(n1985), .CI(
        C[957]), .CO(C[958]) );
  FA_12668 \FA_INST_0[1].FA_INST_1[446].FA_  ( .A(A[958]), .B(n1986), .CI(
        C[958]), .CO(C[959]) );
  FA_12667 \FA_INST_0[1].FA_INST_1[447].FA_  ( .A(A[959]), .B(n1987), .CI(
        C[959]), .CO(C[960]) );
  FA_12666 \FA_INST_0[1].FA_INST_1[448].FA_  ( .A(A[960]), .B(n1988), .CI(
        C[960]), .CO(C[961]) );
  FA_12665 \FA_INST_0[1].FA_INST_1[449].FA_  ( .A(A[961]), .B(n1989), .CI(
        C[961]), .CO(C[962]) );
  FA_12664 \FA_INST_0[1].FA_INST_1[450].FA_  ( .A(A[962]), .B(n1990), .CI(
        C[962]), .CO(C[963]) );
  FA_12663 \FA_INST_0[1].FA_INST_1[451].FA_  ( .A(A[963]), .B(n1991), .CI(
        C[963]), .CO(C[964]) );
  FA_12662 \FA_INST_0[1].FA_INST_1[452].FA_  ( .A(A[964]), .B(n1992), .CI(
        C[964]), .CO(C[965]) );
  FA_12661 \FA_INST_0[1].FA_INST_1[453].FA_  ( .A(A[965]), .B(n1993), .CI(
        C[965]), .CO(C[966]) );
  FA_12660 \FA_INST_0[1].FA_INST_1[454].FA_  ( .A(A[966]), .B(n1994), .CI(
        C[966]), .CO(C[967]) );
  FA_12659 \FA_INST_0[1].FA_INST_1[455].FA_  ( .A(A[967]), .B(n1995), .CI(
        C[967]), .CO(C[968]) );
  FA_12658 \FA_INST_0[1].FA_INST_1[456].FA_  ( .A(A[968]), .B(n1996), .CI(
        C[968]), .CO(C[969]) );
  FA_12657 \FA_INST_0[1].FA_INST_1[457].FA_  ( .A(A[969]), .B(n1997), .CI(
        C[969]), .CO(C[970]) );
  FA_12656 \FA_INST_0[1].FA_INST_1[458].FA_  ( .A(A[970]), .B(n1998), .CI(
        C[970]), .CO(C[971]) );
  FA_12655 \FA_INST_0[1].FA_INST_1[459].FA_  ( .A(A[971]), .B(n1999), .CI(
        C[971]), .CO(C[972]) );
  FA_12654 \FA_INST_0[1].FA_INST_1[460].FA_  ( .A(A[972]), .B(n2000), .CI(
        C[972]), .CO(C[973]) );
  FA_12653 \FA_INST_0[1].FA_INST_1[461].FA_  ( .A(A[973]), .B(n2001), .CI(
        C[973]), .CO(C[974]) );
  FA_12652 \FA_INST_0[1].FA_INST_1[462].FA_  ( .A(A[974]), .B(n2002), .CI(
        C[974]), .CO(C[975]) );
  FA_12651 \FA_INST_0[1].FA_INST_1[463].FA_  ( .A(A[975]), .B(n2003), .CI(
        C[975]), .CO(C[976]) );
  FA_12650 \FA_INST_0[1].FA_INST_1[464].FA_  ( .A(A[976]), .B(n2004), .CI(
        C[976]), .CO(C[977]) );
  FA_12649 \FA_INST_0[1].FA_INST_1[465].FA_  ( .A(A[977]), .B(n2005), .CI(
        C[977]), .CO(C[978]) );
  FA_12648 \FA_INST_0[1].FA_INST_1[466].FA_  ( .A(A[978]), .B(n2006), .CI(
        C[978]), .CO(C[979]) );
  FA_12647 \FA_INST_0[1].FA_INST_1[467].FA_  ( .A(A[979]), .B(n2007), .CI(
        C[979]), .CO(C[980]) );
  FA_12646 \FA_INST_0[1].FA_INST_1[468].FA_  ( .A(A[980]), .B(n2008), .CI(
        C[980]), .CO(C[981]) );
  FA_12645 \FA_INST_0[1].FA_INST_1[469].FA_  ( .A(A[981]), .B(n2009), .CI(
        C[981]), .CO(C[982]) );
  FA_12644 \FA_INST_0[1].FA_INST_1[470].FA_  ( .A(A[982]), .B(n2010), .CI(
        C[982]), .CO(C[983]) );
  FA_12643 \FA_INST_0[1].FA_INST_1[471].FA_  ( .A(A[983]), .B(n2011), .CI(
        C[983]), .CO(C[984]) );
  FA_12642 \FA_INST_0[1].FA_INST_1[472].FA_  ( .A(A[984]), .B(n2012), .CI(
        C[984]), .CO(C[985]) );
  FA_12641 \FA_INST_0[1].FA_INST_1[473].FA_  ( .A(A[985]), .B(n2013), .CI(
        C[985]), .CO(C[986]) );
  FA_12640 \FA_INST_0[1].FA_INST_1[474].FA_  ( .A(A[986]), .B(n2014), .CI(
        C[986]), .CO(C[987]) );
  FA_12639 \FA_INST_0[1].FA_INST_1[475].FA_  ( .A(A[987]), .B(n2015), .CI(
        C[987]), .CO(C[988]) );
  FA_12638 \FA_INST_0[1].FA_INST_1[476].FA_  ( .A(A[988]), .B(n2016), .CI(
        C[988]), .CO(C[989]) );
  FA_12637 \FA_INST_0[1].FA_INST_1[477].FA_  ( .A(A[989]), .B(n2017), .CI(
        C[989]), .CO(C[990]) );
  FA_12636 \FA_INST_0[1].FA_INST_1[478].FA_  ( .A(A[990]), .B(n2018), .CI(
        C[990]), .CO(C[991]) );
  FA_12635 \FA_INST_0[1].FA_INST_1[479].FA_  ( .A(A[991]), .B(n2019), .CI(
        C[991]), .CO(C[992]) );
  FA_12634 \FA_INST_0[1].FA_INST_1[480].FA_  ( .A(A[992]), .B(n2020), .CI(
        C[992]), .CO(C[993]) );
  FA_12633 \FA_INST_0[1].FA_INST_1[481].FA_  ( .A(A[993]), .B(n2021), .CI(
        C[993]), .CO(C[994]) );
  FA_12632 \FA_INST_0[1].FA_INST_1[482].FA_  ( .A(A[994]), .B(n2022), .CI(
        C[994]), .CO(C[995]) );
  FA_12631 \FA_INST_0[1].FA_INST_1[483].FA_  ( .A(A[995]), .B(n2023), .CI(
        C[995]), .CO(C[996]) );
  FA_12630 \FA_INST_0[1].FA_INST_1[484].FA_  ( .A(A[996]), .B(n2024), .CI(
        C[996]), .CO(C[997]) );
  FA_12629 \FA_INST_0[1].FA_INST_1[485].FA_  ( .A(A[997]), .B(n2025), .CI(
        C[997]), .CO(C[998]) );
  FA_12628 \FA_INST_0[1].FA_INST_1[486].FA_  ( .A(A[998]), .B(n2026), .CI(
        C[998]), .CO(C[999]) );
  FA_12627 \FA_INST_0[1].FA_INST_1[487].FA_  ( .A(A[999]), .B(n2027), .CI(
        C[999]), .CO(C[1000]) );
  FA_12626 \FA_INST_0[1].FA_INST_1[488].FA_  ( .A(A[1000]), .B(n2028), .CI(
        C[1000]), .CO(C[1001]) );
  FA_12625 \FA_INST_0[1].FA_INST_1[489].FA_  ( .A(A[1001]), .B(n2029), .CI(
        C[1001]), .CO(C[1002]) );
  FA_12624 \FA_INST_0[1].FA_INST_1[490].FA_  ( .A(A[1002]), .B(n2030), .CI(
        C[1002]), .CO(C[1003]) );
  FA_12623 \FA_INST_0[1].FA_INST_1[491].FA_  ( .A(A[1003]), .B(n2031), .CI(
        C[1003]), .CO(C[1004]) );
  FA_12622 \FA_INST_0[1].FA_INST_1[492].FA_  ( .A(A[1004]), .B(n2032), .CI(
        C[1004]), .CO(C[1005]) );
  FA_12621 \FA_INST_0[1].FA_INST_1[493].FA_  ( .A(A[1005]), .B(n2033), .CI(
        C[1005]), .CO(C[1006]) );
  FA_12620 \FA_INST_0[1].FA_INST_1[494].FA_  ( .A(A[1006]), .B(n2034), .CI(
        C[1006]), .CO(C[1007]) );
  FA_12619 \FA_INST_0[1].FA_INST_1[495].FA_  ( .A(A[1007]), .B(n2035), .CI(
        C[1007]), .CO(C[1008]) );
  FA_12618 \FA_INST_0[1].FA_INST_1[496].FA_  ( .A(A[1008]), .B(n2036), .CI(
        C[1008]), .CO(C[1009]) );
  FA_12617 \FA_INST_0[1].FA_INST_1[497].FA_  ( .A(A[1009]), .B(n2037), .CI(
        C[1009]), .CO(C[1010]) );
  FA_12616 \FA_INST_0[1].FA_INST_1[498].FA_  ( .A(A[1010]), .B(n2038), .CI(
        C[1010]), .CO(C[1011]) );
  FA_12615 \FA_INST_0[1].FA_INST_1[499].FA_  ( .A(A[1011]), .B(n2039), .CI(
        C[1011]), .CO(C[1012]) );
  FA_12614 \FA_INST_0[1].FA_INST_1[500].FA_  ( .A(A[1012]), .B(n2040), .CI(
        C[1012]), .CO(C[1013]) );
  FA_12613 \FA_INST_0[1].FA_INST_1[501].FA_  ( .A(A[1013]), .B(n2041), .CI(
        C[1013]), .CO(C[1014]) );
  FA_12612 \FA_INST_0[1].FA_INST_1[502].FA_  ( .A(A[1014]), .B(n2042), .CI(
        C[1014]), .CO(C[1015]) );
  FA_12611 \FA_INST_0[1].FA_INST_1[503].FA_  ( .A(A[1015]), .B(n2043), .CI(
        C[1015]), .CO(C[1016]) );
  FA_12610 \FA_INST_0[1].FA_INST_1[504].FA_  ( .A(A[1016]), .B(n2044), .CI(
        C[1016]), .CO(C[1017]) );
  FA_12609 \FA_INST_0[1].FA_INST_1[505].FA_  ( .A(A[1017]), .B(n2045), .CI(
        C[1017]), .CO(C[1018]) );
  FA_12608 \FA_INST_0[1].FA_INST_1[506].FA_  ( .A(A[1018]), .B(n2046), .CI(
        C[1018]), .CO(C[1019]) );
  FA_12607 \FA_INST_0[1].FA_INST_1[507].FA_  ( .A(A[1019]), .B(n2047), .CI(
        C[1019]), .CO(C[1020]) );
  FA_12606 \FA_INST_0[1].FA_INST_1[508].FA_  ( .A(A[1020]), .B(n2048), .CI(
        C[1020]), .CO(C[1021]) );
  FA_12605 \FA_INST_0[1].FA_INST_1[509].FA_  ( .A(A[1021]), .B(n2049), .CI(
        C[1021]), .CO(C[1022]) );
  FA_12604 \FA_INST_0[1].FA_INST_1[510].FA_  ( .A(A[1022]), .B(n2050), .CI(
        C[1022]), .CO(C[1023]) );
  FA_12603 \FA_INST_0[1].FA_INST_1[511].FA_  ( .A(A[1023]), .B(n2051), .CI(
        C[1023]), .CO(C[1024]) );
  FA_12602 \FA_INST_1[1024].FA_  ( .A(1'b0), .B(n2052), .CI(C[1024]), .CO(
        C[1025]) );
  FA_12601 \FA_INST_1[1025].FA_  ( .A(1'b0), .B(n2053), .CI(C[1025]), .CO(O)
         );
  IV U2 ( .A(B[27]), .Z(n1055) );
  IV U3 ( .A(B[28]), .Z(n1056) );
  IV U4 ( .A(B[29]), .Z(n1057) );
  IV U5 ( .A(B[30]), .Z(n1058) );
  IV U6 ( .A(B[31]), .Z(n1059) );
  IV U7 ( .A(B[32]), .Z(n1060) );
  IV U8 ( .A(B[33]), .Z(n1061) );
  IV U9 ( .A(B[34]), .Z(n1062) );
  IV U10 ( .A(B[35]), .Z(n1063) );
  IV U11 ( .A(B[36]), .Z(n1064) );
  IV U12 ( .A(B[927]), .Z(n1955) );
  IV U13 ( .A(B[37]), .Z(n1065) );
  IV U14 ( .A(B[38]), .Z(n1066) );
  IV U15 ( .A(B[39]), .Z(n1067) );
  IV U16 ( .A(B[40]), .Z(n1068) );
  IV U17 ( .A(B[41]), .Z(n1069) );
  IV U18 ( .A(B[42]), .Z(n1070) );
  IV U19 ( .A(B[43]), .Z(n1071) );
  IV U20 ( .A(B[44]), .Z(n1072) );
  IV U21 ( .A(B[45]), .Z(n1073) );
  IV U22 ( .A(B[46]), .Z(n1074) );
  IV U23 ( .A(B[928]), .Z(n1956) );
  IV U24 ( .A(B[47]), .Z(n1075) );
  IV U25 ( .A(B[48]), .Z(n1076) );
  IV U26 ( .A(B[49]), .Z(n1077) );
  IV U27 ( .A(B[50]), .Z(n1078) );
  IV U28 ( .A(B[51]), .Z(n1079) );
  IV U29 ( .A(B[52]), .Z(n1080) );
  IV U30 ( .A(B[53]), .Z(n1081) );
  IV U31 ( .A(B[54]), .Z(n1082) );
  IV U32 ( .A(B[55]), .Z(n1083) );
  IV U33 ( .A(B[56]), .Z(n1084) );
  IV U34 ( .A(B[929]), .Z(n1957) );
  IV U35 ( .A(B[57]), .Z(n1085) );
  IV U36 ( .A(B[58]), .Z(n1086) );
  IV U37 ( .A(B[59]), .Z(n1087) );
  IV U38 ( .A(B[60]), .Z(n1088) );
  IV U39 ( .A(B[61]), .Z(n1089) );
  IV U40 ( .A(B[62]), .Z(n1090) );
  IV U41 ( .A(B[63]), .Z(n1091) );
  IV U42 ( .A(B[64]), .Z(n1092) );
  IV U43 ( .A(B[65]), .Z(n1093) );
  IV U44 ( .A(B[66]), .Z(n1094) );
  IV U45 ( .A(B[930]), .Z(n1958) );
  IV U46 ( .A(B[67]), .Z(n1095) );
  IV U47 ( .A(B[68]), .Z(n1096) );
  IV U48 ( .A(B[69]), .Z(n1097) );
  IV U49 ( .A(B[70]), .Z(n1098) );
  IV U50 ( .A(B[71]), .Z(n1099) );
  IV U51 ( .A(B[72]), .Z(n1100) );
  IV U52 ( .A(B[73]), .Z(n1101) );
  IV U53 ( .A(B[74]), .Z(n1102) );
  IV U54 ( .A(B[75]), .Z(n1103) );
  IV U55 ( .A(B[76]), .Z(n1104) );
  IV U56 ( .A(B[931]), .Z(n1959) );
  IV U57 ( .A(B[77]), .Z(n1105) );
  IV U58 ( .A(B[78]), .Z(n1106) );
  IV U59 ( .A(B[79]), .Z(n1107) );
  IV U60 ( .A(B[80]), .Z(n1108) );
  IV U61 ( .A(B[81]), .Z(n1109) );
  IV U62 ( .A(B[82]), .Z(n1110) );
  IV U63 ( .A(B[83]), .Z(n1111) );
  IV U64 ( .A(B[84]), .Z(n1112) );
  IV U65 ( .A(B[85]), .Z(n1113) );
  IV U66 ( .A(B[86]), .Z(n1114) );
  IV U67 ( .A(B[932]), .Z(n1960) );
  IV U68 ( .A(B[87]), .Z(n1115) );
  IV U69 ( .A(B[88]), .Z(n1116) );
  IV U70 ( .A(B[89]), .Z(n1117) );
  IV U71 ( .A(B[90]), .Z(n1118) );
  IV U72 ( .A(B[91]), .Z(n1119) );
  IV U73 ( .A(B[92]), .Z(n1120) );
  IV U74 ( .A(B[93]), .Z(n1121) );
  IV U75 ( .A(B[94]), .Z(n1122) );
  IV U76 ( .A(B[95]), .Z(n1123) );
  IV U77 ( .A(B[96]), .Z(n1124) );
  IV U78 ( .A(B[933]), .Z(n1961) );
  IV U79 ( .A(B[97]), .Z(n1125) );
  IV U80 ( .A(B[98]), .Z(n1126) );
  IV U81 ( .A(B[99]), .Z(n1127) );
  IV U82 ( .A(B[100]), .Z(n1128) );
  IV U83 ( .A(B[101]), .Z(n1129) );
  IV U84 ( .A(B[102]), .Z(n1130) );
  IV U85 ( .A(B[103]), .Z(n1131) );
  IV U86 ( .A(B[104]), .Z(n1132) );
  IV U87 ( .A(B[105]), .Z(n1133) );
  IV U88 ( .A(B[106]), .Z(n1134) );
  IV U89 ( .A(B[934]), .Z(n1962) );
  IV U90 ( .A(B[107]), .Z(n1135) );
  IV U91 ( .A(B[108]), .Z(n1136) );
  IV U92 ( .A(B[109]), .Z(n1137) );
  IV U93 ( .A(B[110]), .Z(n1138) );
  IV U94 ( .A(B[111]), .Z(n1139) );
  IV U95 ( .A(B[112]), .Z(n1140) );
  IV U96 ( .A(B[113]), .Z(n1141) );
  IV U97 ( .A(B[114]), .Z(n1142) );
  IV U98 ( .A(B[115]), .Z(n1143) );
  IV U99 ( .A(B[116]), .Z(n1144) );
  IV U100 ( .A(B[935]), .Z(n1963) );
  IV U101 ( .A(B[117]), .Z(n1145) );
  IV U102 ( .A(B[118]), .Z(n1146) );
  IV U103 ( .A(B[119]), .Z(n1147) );
  IV U104 ( .A(B[120]), .Z(n1148) );
  IV U105 ( .A(B[121]), .Z(n1149) );
  IV U106 ( .A(B[122]), .Z(n1150) );
  IV U107 ( .A(B[123]), .Z(n1151) );
  IV U108 ( .A(B[124]), .Z(n1152) );
  IV U109 ( .A(B[125]), .Z(n1153) );
  IV U110 ( .A(B[126]), .Z(n1154) );
  IV U111 ( .A(B[936]), .Z(n1964) );
  IV U112 ( .A(B[1017]), .Z(n2045) );
  IV U113 ( .A(B[127]), .Z(n1155) );
  IV U114 ( .A(B[128]), .Z(n1156) );
  IV U115 ( .A(B[129]), .Z(n1157) );
  IV U116 ( .A(B[130]), .Z(n1158) );
  IV U117 ( .A(B[131]), .Z(n1159) );
  IV U118 ( .A(B[132]), .Z(n1160) );
  IV U119 ( .A(B[133]), .Z(n1161) );
  IV U120 ( .A(B[134]), .Z(n1162) );
  IV U121 ( .A(B[135]), .Z(n1163) );
  IV U122 ( .A(B[136]), .Z(n1164) );
  IV U123 ( .A(B[937]), .Z(n1965) );
  IV U124 ( .A(B[137]), .Z(n1165) );
  IV U125 ( .A(B[138]), .Z(n1166) );
  IV U126 ( .A(B[139]), .Z(n1167) );
  IV U127 ( .A(B[140]), .Z(n1168) );
  IV U128 ( .A(B[141]), .Z(n1169) );
  IV U129 ( .A(B[142]), .Z(n1170) );
  IV U130 ( .A(B[143]), .Z(n1171) );
  IV U131 ( .A(B[144]), .Z(n1172) );
  IV U132 ( .A(B[145]), .Z(n1173) );
  IV U133 ( .A(B[146]), .Z(n1174) );
  IV U134 ( .A(B[938]), .Z(n1966) );
  IV U135 ( .A(B[147]), .Z(n1175) );
  IV U136 ( .A(B[148]), .Z(n1176) );
  IV U137 ( .A(B[149]), .Z(n1177) );
  IV U138 ( .A(B[150]), .Z(n1178) );
  IV U139 ( .A(B[151]), .Z(n1179) );
  IV U140 ( .A(B[152]), .Z(n1180) );
  IV U141 ( .A(B[153]), .Z(n1181) );
  IV U142 ( .A(B[154]), .Z(n1182) );
  IV U143 ( .A(B[155]), .Z(n1183) );
  IV U144 ( .A(B[156]), .Z(n1184) );
  IV U145 ( .A(B[939]), .Z(n1967) );
  IV U146 ( .A(B[157]), .Z(n1185) );
  IV U147 ( .A(B[158]), .Z(n1186) );
  IV U148 ( .A(B[159]), .Z(n1187) );
  IV U149 ( .A(B[160]), .Z(n1188) );
  IV U150 ( .A(B[161]), .Z(n1189) );
  IV U151 ( .A(B[162]), .Z(n1190) );
  IV U152 ( .A(B[163]), .Z(n1191) );
  IV U153 ( .A(B[164]), .Z(n1192) );
  IV U154 ( .A(B[165]), .Z(n1193) );
  IV U155 ( .A(B[166]), .Z(n1194) );
  IV U156 ( .A(B[940]), .Z(n1968) );
  IV U157 ( .A(B[167]), .Z(n1195) );
  IV U158 ( .A(B[168]), .Z(n1196) );
  IV U159 ( .A(B[169]), .Z(n1197) );
  IV U160 ( .A(B[170]), .Z(n1198) );
  IV U161 ( .A(B[171]), .Z(n1199) );
  IV U162 ( .A(B[172]), .Z(n1200) );
  IV U163 ( .A(B[173]), .Z(n1201) );
  IV U164 ( .A(B[174]), .Z(n1202) );
  IV U165 ( .A(B[175]), .Z(n1203) );
  IV U166 ( .A(B[176]), .Z(n1204) );
  IV U167 ( .A(B[941]), .Z(n1969) );
  IV U168 ( .A(B[177]), .Z(n1205) );
  IV U169 ( .A(B[178]), .Z(n1206) );
  IV U170 ( .A(B[179]), .Z(n1207) );
  IV U171 ( .A(B[180]), .Z(n1208) );
  IV U172 ( .A(B[181]), .Z(n1209) );
  IV U173 ( .A(B[182]), .Z(n1210) );
  IV U174 ( .A(B[183]), .Z(n1211) );
  IV U175 ( .A(B[184]), .Z(n1212) );
  IV U176 ( .A(B[185]), .Z(n1213) );
  IV U177 ( .A(B[186]), .Z(n1214) );
  IV U178 ( .A(B[942]), .Z(n1970) );
  IV U179 ( .A(B[187]), .Z(n1215) );
  IV U180 ( .A(B[188]), .Z(n1216) );
  IV U181 ( .A(B[189]), .Z(n1217) );
  IV U182 ( .A(B[190]), .Z(n1218) );
  IV U183 ( .A(B[191]), .Z(n1219) );
  IV U184 ( .A(B[192]), .Z(n1220) );
  IV U185 ( .A(B[193]), .Z(n1221) );
  IV U186 ( .A(B[194]), .Z(n1222) );
  IV U187 ( .A(B[195]), .Z(n1223) );
  IV U188 ( .A(B[196]), .Z(n1224) );
  IV U189 ( .A(B[943]), .Z(n1971) );
  IV U190 ( .A(B[197]), .Z(n1225) );
  IV U191 ( .A(B[198]), .Z(n1226) );
  IV U192 ( .A(B[199]), .Z(n1227) );
  IV U193 ( .A(B[200]), .Z(n1228) );
  IV U194 ( .A(B[201]), .Z(n1229) );
  IV U195 ( .A(B[202]), .Z(n1230) );
  IV U196 ( .A(B[203]), .Z(n1231) );
  IV U197 ( .A(B[204]), .Z(n1232) );
  IV U198 ( .A(B[205]), .Z(n1233) );
  IV U199 ( .A(B[206]), .Z(n1234) );
  IV U200 ( .A(B[944]), .Z(n1972) );
  IV U201 ( .A(B[207]), .Z(n1235) );
  IV U202 ( .A(B[208]), .Z(n1236) );
  IV U203 ( .A(B[209]), .Z(n1237) );
  IV U204 ( .A(B[210]), .Z(n1238) );
  IV U205 ( .A(B[211]), .Z(n1239) );
  IV U206 ( .A(B[212]), .Z(n1240) );
  IV U207 ( .A(B[213]), .Z(n1241) );
  IV U208 ( .A(B[214]), .Z(n1242) );
  IV U209 ( .A(B[215]), .Z(n1243) );
  IV U210 ( .A(B[216]), .Z(n1244) );
  IV U211 ( .A(B[945]), .Z(n1973) );
  IV U212 ( .A(B[217]), .Z(n1245) );
  IV U213 ( .A(B[218]), .Z(n1246) );
  IV U214 ( .A(B[219]), .Z(n1247) );
  IV U215 ( .A(B[220]), .Z(n1248) );
  IV U216 ( .A(B[221]), .Z(n1249) );
  IV U217 ( .A(B[222]), .Z(n1250) );
  IV U218 ( .A(B[223]), .Z(n1251) );
  IV U219 ( .A(B[224]), .Z(n1252) );
  IV U220 ( .A(B[225]), .Z(n1253) );
  IV U221 ( .A(B[226]), .Z(n1254) );
  IV U222 ( .A(B[946]), .Z(n1974) );
  IV U223 ( .A(B[1018]), .Z(n2046) );
  IV U224 ( .A(B[227]), .Z(n1255) );
  IV U225 ( .A(B[228]), .Z(n1256) );
  IV U226 ( .A(B[229]), .Z(n1257) );
  IV U227 ( .A(B[230]), .Z(n1258) );
  IV U228 ( .A(B[231]), .Z(n1259) );
  IV U229 ( .A(B[232]), .Z(n1260) );
  IV U230 ( .A(B[233]), .Z(n1261) );
  IV U231 ( .A(B[234]), .Z(n1262) );
  IV U232 ( .A(B[235]), .Z(n1263) );
  IV U233 ( .A(B[236]), .Z(n1264) );
  IV U234 ( .A(B[947]), .Z(n1975) );
  IV U235 ( .A(B[237]), .Z(n1265) );
  IV U236 ( .A(B[238]), .Z(n1266) );
  IV U237 ( .A(B[239]), .Z(n1267) );
  IV U238 ( .A(B[240]), .Z(n1268) );
  IV U239 ( .A(B[241]), .Z(n1269) );
  IV U240 ( .A(B[242]), .Z(n1270) );
  IV U241 ( .A(B[243]), .Z(n1271) );
  IV U242 ( .A(B[244]), .Z(n1272) );
  IV U243 ( .A(B[245]), .Z(n1273) );
  IV U244 ( .A(B[246]), .Z(n1274) );
  IV U245 ( .A(B[948]), .Z(n1976) );
  IV U246 ( .A(B[247]), .Z(n1275) );
  IV U247 ( .A(B[248]), .Z(n1276) );
  IV U248 ( .A(B[249]), .Z(n1277) );
  IV U249 ( .A(B[250]), .Z(n1278) );
  IV U250 ( .A(B[251]), .Z(n1279) );
  IV U251 ( .A(B[252]), .Z(n1280) );
  IV U252 ( .A(B[253]), .Z(n1281) );
  IV U253 ( .A(B[254]), .Z(n1282) );
  IV U254 ( .A(B[255]), .Z(n1283) );
  IV U255 ( .A(B[256]), .Z(n1284) );
  IV U256 ( .A(B[949]), .Z(n1977) );
  IV U257 ( .A(B[257]), .Z(n1285) );
  IV U258 ( .A(B[258]), .Z(n1286) );
  IV U259 ( .A(B[259]), .Z(n1287) );
  IV U260 ( .A(B[260]), .Z(n1288) );
  IV U261 ( .A(B[261]), .Z(n1289) );
  IV U262 ( .A(B[262]), .Z(n1290) );
  IV U263 ( .A(B[263]), .Z(n1291) );
  IV U264 ( .A(B[264]), .Z(n1292) );
  IV U265 ( .A(B[265]), .Z(n1293) );
  IV U266 ( .A(B[266]), .Z(n1294) );
  IV U267 ( .A(B[950]), .Z(n1978) );
  IV U268 ( .A(B[267]), .Z(n1295) );
  IV U269 ( .A(B[268]), .Z(n1296) );
  IV U270 ( .A(B[269]), .Z(n1297) );
  IV U271 ( .A(B[270]), .Z(n1298) );
  IV U272 ( .A(B[271]), .Z(n1299) );
  IV U273 ( .A(B[272]), .Z(n1300) );
  IV U274 ( .A(B[273]), .Z(n1301) );
  IV U275 ( .A(B[274]), .Z(n1302) );
  IV U276 ( .A(B[275]), .Z(n1303) );
  IV U277 ( .A(B[276]), .Z(n1304) );
  IV U278 ( .A(B[951]), .Z(n1979) );
  IV U279 ( .A(B[277]), .Z(n1305) );
  IV U280 ( .A(B[278]), .Z(n1306) );
  IV U281 ( .A(B[279]), .Z(n1307) );
  IV U282 ( .A(B[280]), .Z(n1308) );
  IV U283 ( .A(B[281]), .Z(n1309) );
  IV U284 ( .A(B[282]), .Z(n1310) );
  IV U285 ( .A(B[283]), .Z(n1311) );
  IV U286 ( .A(B[284]), .Z(n1312) );
  IV U287 ( .A(B[285]), .Z(n1313) );
  IV U288 ( .A(B[286]), .Z(n1314) );
  IV U289 ( .A(B[952]), .Z(n1980) );
  IV U290 ( .A(B[287]), .Z(n1315) );
  IV U291 ( .A(B[288]), .Z(n1316) );
  IV U292 ( .A(B[289]), .Z(n1317) );
  IV U293 ( .A(B[290]), .Z(n1318) );
  IV U294 ( .A(B[291]), .Z(n1319) );
  IV U295 ( .A(B[292]), .Z(n1320) );
  IV U296 ( .A(B[293]), .Z(n1321) );
  IV U297 ( .A(B[294]), .Z(n1322) );
  IV U298 ( .A(B[295]), .Z(n1323) );
  IV U299 ( .A(B[296]), .Z(n1324) );
  IV U300 ( .A(B[953]), .Z(n1981) );
  IV U301 ( .A(B[297]), .Z(n1325) );
  IV U302 ( .A(B[298]), .Z(n1326) );
  IV U303 ( .A(B[299]), .Z(n1327) );
  IV U304 ( .A(B[300]), .Z(n1328) );
  IV U305 ( .A(B[301]), .Z(n1329) );
  IV U306 ( .A(B[302]), .Z(n1330) );
  IV U307 ( .A(B[303]), .Z(n1331) );
  IV U308 ( .A(B[304]), .Z(n1332) );
  IV U309 ( .A(B[305]), .Z(n1333) );
  IV U310 ( .A(B[306]), .Z(n1334) );
  IV U311 ( .A(B[954]), .Z(n1982) );
  IV U312 ( .A(B[307]), .Z(n1335) );
  IV U313 ( .A(B[308]), .Z(n1336) );
  IV U314 ( .A(B[309]), .Z(n1337) );
  IV U315 ( .A(B[310]), .Z(n1338) );
  IV U316 ( .A(B[311]), .Z(n1339) );
  IV U317 ( .A(B[312]), .Z(n1340) );
  IV U318 ( .A(B[313]), .Z(n1341) );
  IV U319 ( .A(B[314]), .Z(n1342) );
  IV U320 ( .A(B[315]), .Z(n1343) );
  IV U321 ( .A(B[316]), .Z(n1344) );
  IV U322 ( .A(B[955]), .Z(n1983) );
  IV U323 ( .A(B[317]), .Z(n1345) );
  IV U324 ( .A(B[318]), .Z(n1346) );
  IV U325 ( .A(B[319]), .Z(n1347) );
  IV U326 ( .A(B[320]), .Z(n1348) );
  IV U327 ( .A(B[321]), .Z(n1349) );
  IV U328 ( .A(B[322]), .Z(n1350) );
  IV U329 ( .A(B[323]), .Z(n1351) );
  IV U330 ( .A(B[324]), .Z(n1352) );
  IV U331 ( .A(B[325]), .Z(n1353) );
  IV U332 ( .A(B[326]), .Z(n1354) );
  IV U333 ( .A(B[956]), .Z(n1984) );
  IV U334 ( .A(B[1019]), .Z(n2047) );
  IV U335 ( .A(B[327]), .Z(n1355) );
  IV U336 ( .A(B[328]), .Z(n1356) );
  IV U337 ( .A(B[329]), .Z(n1357) );
  IV U338 ( .A(B[330]), .Z(n1358) );
  IV U339 ( .A(B[331]), .Z(n1359) );
  IV U340 ( .A(B[332]), .Z(n1360) );
  IV U341 ( .A(B[333]), .Z(n1361) );
  IV U342 ( .A(B[334]), .Z(n1362) );
  IV U343 ( .A(B[335]), .Z(n1363) );
  IV U344 ( .A(B[336]), .Z(n1364) );
  IV U345 ( .A(B[957]), .Z(n1985) );
  IV U346 ( .A(B[337]), .Z(n1365) );
  IV U347 ( .A(B[338]), .Z(n1366) );
  IV U348 ( .A(B[339]), .Z(n1367) );
  IV U349 ( .A(B[340]), .Z(n1368) );
  IV U350 ( .A(B[341]), .Z(n1369) );
  IV U351 ( .A(B[342]), .Z(n1370) );
  IV U352 ( .A(B[343]), .Z(n1371) );
  IV U353 ( .A(B[344]), .Z(n1372) );
  IV U354 ( .A(B[345]), .Z(n1373) );
  IV U355 ( .A(B[346]), .Z(n1374) );
  IV U356 ( .A(B[958]), .Z(n1986) );
  IV U357 ( .A(B[347]), .Z(n1375) );
  IV U358 ( .A(B[348]), .Z(n1376) );
  IV U359 ( .A(B[349]), .Z(n1377) );
  IV U360 ( .A(B[350]), .Z(n1378) );
  IV U361 ( .A(B[351]), .Z(n1379) );
  IV U362 ( .A(B[352]), .Z(n1380) );
  IV U363 ( .A(B[353]), .Z(n1381) );
  IV U364 ( .A(B[354]), .Z(n1382) );
  IV U365 ( .A(B[355]), .Z(n1383) );
  IV U366 ( .A(B[356]), .Z(n1384) );
  IV U367 ( .A(B[959]), .Z(n1987) );
  IV U368 ( .A(B[357]), .Z(n1385) );
  IV U369 ( .A(B[358]), .Z(n1386) );
  IV U370 ( .A(B[359]), .Z(n1387) );
  IV U371 ( .A(B[360]), .Z(n1388) );
  IV U372 ( .A(B[361]), .Z(n1389) );
  IV U373 ( .A(B[362]), .Z(n1390) );
  IV U374 ( .A(B[363]), .Z(n1391) );
  IV U375 ( .A(B[364]), .Z(n1392) );
  IV U376 ( .A(B[365]), .Z(n1393) );
  IV U377 ( .A(B[366]), .Z(n1394) );
  IV U378 ( .A(B[960]), .Z(n1988) );
  IV U379 ( .A(B[367]), .Z(n1395) );
  IV U380 ( .A(B[368]), .Z(n1396) );
  IV U381 ( .A(B[369]), .Z(n1397) );
  IV U382 ( .A(B[370]), .Z(n1398) );
  IV U383 ( .A(B[371]), .Z(n1399) );
  IV U384 ( .A(B[372]), .Z(n1400) );
  IV U385 ( .A(B[373]), .Z(n1401) );
  IV U386 ( .A(B[374]), .Z(n1402) );
  IV U387 ( .A(B[375]), .Z(n1403) );
  IV U388 ( .A(B[376]), .Z(n1404) );
  IV U389 ( .A(B[961]), .Z(n1989) );
  IV U390 ( .A(B[377]), .Z(n1405) );
  IV U391 ( .A(B[378]), .Z(n1406) );
  IV U392 ( .A(B[379]), .Z(n1407) );
  IV U393 ( .A(B[380]), .Z(n1408) );
  IV U394 ( .A(B[381]), .Z(n1409) );
  IV U395 ( .A(B[382]), .Z(n1410) );
  IV U396 ( .A(B[383]), .Z(n1411) );
  IV U397 ( .A(B[384]), .Z(n1412) );
  IV U398 ( .A(B[385]), .Z(n1413) );
  IV U399 ( .A(B[386]), .Z(n1414) );
  IV U400 ( .A(B[962]), .Z(n1990) );
  IV U401 ( .A(B[387]), .Z(n1415) );
  IV U402 ( .A(B[388]), .Z(n1416) );
  IV U403 ( .A(B[389]), .Z(n1417) );
  IV U404 ( .A(B[390]), .Z(n1418) );
  IV U405 ( .A(B[391]), .Z(n1419) );
  IV U406 ( .A(B[392]), .Z(n1420) );
  IV U407 ( .A(B[393]), .Z(n1421) );
  IV U408 ( .A(B[394]), .Z(n1422) );
  IV U409 ( .A(B[395]), .Z(n1423) );
  IV U410 ( .A(B[396]), .Z(n1424) );
  IV U411 ( .A(B[963]), .Z(n1991) );
  IV U412 ( .A(B[397]), .Z(n1425) );
  IV U413 ( .A(B[398]), .Z(n1426) );
  IV U414 ( .A(B[399]), .Z(n1427) );
  IV U415 ( .A(B[400]), .Z(n1428) );
  IV U416 ( .A(B[401]), .Z(n1429) );
  IV U417 ( .A(B[402]), .Z(n1430) );
  IV U418 ( .A(B[403]), .Z(n1431) );
  IV U419 ( .A(B[404]), .Z(n1432) );
  IV U420 ( .A(B[405]), .Z(n1433) );
  IV U421 ( .A(B[406]), .Z(n1434) );
  IV U422 ( .A(B[964]), .Z(n1992) );
  IV U423 ( .A(B[407]), .Z(n1435) );
  IV U424 ( .A(B[408]), .Z(n1436) );
  IV U425 ( .A(B[409]), .Z(n1437) );
  IV U426 ( .A(B[410]), .Z(n1438) );
  IV U427 ( .A(B[411]), .Z(n1439) );
  IV U428 ( .A(B[412]), .Z(n1440) );
  IV U429 ( .A(B[413]), .Z(n1441) );
  IV U430 ( .A(B[414]), .Z(n1442) );
  IV U431 ( .A(B[415]), .Z(n1443) );
  IV U432 ( .A(B[416]), .Z(n1444) );
  IV U433 ( .A(B[965]), .Z(n1993) );
  IV U434 ( .A(B[417]), .Z(n1445) );
  IV U435 ( .A(B[418]), .Z(n1446) );
  IV U436 ( .A(B[419]), .Z(n1447) );
  IV U437 ( .A(B[420]), .Z(n1448) );
  IV U438 ( .A(B[421]), .Z(n1449) );
  IV U439 ( .A(B[422]), .Z(n1450) );
  IV U440 ( .A(B[423]), .Z(n1451) );
  IV U441 ( .A(B[424]), .Z(n1452) );
  IV U442 ( .A(B[425]), .Z(n1453) );
  IV U443 ( .A(B[426]), .Z(n1454) );
  IV U444 ( .A(B[966]), .Z(n1994) );
  IV U445 ( .A(B[1020]), .Z(n2048) );
  IV U446 ( .A(B[427]), .Z(n1455) );
  IV U447 ( .A(B[428]), .Z(n1456) );
  IV U448 ( .A(B[429]), .Z(n1457) );
  IV U449 ( .A(B[430]), .Z(n1458) );
  IV U450 ( .A(B[431]), .Z(n1459) );
  IV U451 ( .A(B[432]), .Z(n1460) );
  IV U452 ( .A(B[433]), .Z(n1461) );
  IV U453 ( .A(B[434]), .Z(n1462) );
  IV U454 ( .A(B[435]), .Z(n1463) );
  IV U455 ( .A(B[436]), .Z(n1464) );
  IV U456 ( .A(B[967]), .Z(n1995) );
  IV U457 ( .A(B[437]), .Z(n1465) );
  IV U458 ( .A(B[438]), .Z(n1466) );
  IV U459 ( .A(B[439]), .Z(n1467) );
  IV U460 ( .A(B[440]), .Z(n1468) );
  IV U461 ( .A(B[441]), .Z(n1469) );
  IV U462 ( .A(B[442]), .Z(n1470) );
  IV U463 ( .A(B[443]), .Z(n1471) );
  IV U464 ( .A(B[444]), .Z(n1472) );
  IV U465 ( .A(B[445]), .Z(n1473) );
  IV U466 ( .A(B[446]), .Z(n1474) );
  IV U467 ( .A(B[968]), .Z(n1996) );
  IV U468 ( .A(B[447]), .Z(n1475) );
  IV U469 ( .A(B[448]), .Z(n1476) );
  IV U470 ( .A(B[449]), .Z(n1477) );
  IV U471 ( .A(B[450]), .Z(n1478) );
  IV U472 ( .A(B[451]), .Z(n1479) );
  IV U473 ( .A(B[452]), .Z(n1480) );
  IV U474 ( .A(B[453]), .Z(n1481) );
  IV U475 ( .A(B[454]), .Z(n1482) );
  IV U476 ( .A(B[455]), .Z(n1483) );
  IV U477 ( .A(B[456]), .Z(n1484) );
  IV U478 ( .A(B[969]), .Z(n1997) );
  IV U479 ( .A(B[457]), .Z(n1485) );
  IV U480 ( .A(B[458]), .Z(n1486) );
  IV U481 ( .A(B[459]), .Z(n1487) );
  IV U482 ( .A(B[460]), .Z(n1488) );
  IV U483 ( .A(B[461]), .Z(n1489) );
  IV U484 ( .A(B[462]), .Z(n1490) );
  IV U485 ( .A(B[463]), .Z(n1491) );
  IV U486 ( .A(B[464]), .Z(n1492) );
  IV U487 ( .A(B[465]), .Z(n1493) );
  IV U488 ( .A(B[466]), .Z(n1494) );
  IV U489 ( .A(B[970]), .Z(n1998) );
  IV U490 ( .A(B[467]), .Z(n1495) );
  IV U491 ( .A(B[468]), .Z(n1496) );
  IV U492 ( .A(B[469]), .Z(n1497) );
  IV U493 ( .A(B[470]), .Z(n1498) );
  IV U494 ( .A(B[471]), .Z(n1499) );
  IV U495 ( .A(B[472]), .Z(n1500) );
  IV U496 ( .A(B[473]), .Z(n1501) );
  IV U497 ( .A(B[474]), .Z(n1502) );
  IV U498 ( .A(B[475]), .Z(n1503) );
  IV U499 ( .A(B[476]), .Z(n1504) );
  IV U500 ( .A(B[971]), .Z(n1999) );
  IV U501 ( .A(B[477]), .Z(n1505) );
  IV U502 ( .A(B[478]), .Z(n1506) );
  IV U503 ( .A(B[479]), .Z(n1507) );
  IV U504 ( .A(B[480]), .Z(n1508) );
  IV U505 ( .A(B[481]), .Z(n1509) );
  IV U506 ( .A(B[482]), .Z(n1510) );
  IV U507 ( .A(B[483]), .Z(n1511) );
  IV U508 ( .A(B[484]), .Z(n1512) );
  IV U509 ( .A(B[485]), .Z(n1513) );
  IV U510 ( .A(B[486]), .Z(n1514) );
  IV U511 ( .A(B[972]), .Z(n2000) );
  IV U512 ( .A(B[487]), .Z(n1515) );
  IV U513 ( .A(B[488]), .Z(n1516) );
  IV U514 ( .A(B[489]), .Z(n1517) );
  IV U515 ( .A(B[490]), .Z(n1518) );
  IV U516 ( .A(B[491]), .Z(n1519) );
  IV U517 ( .A(B[492]), .Z(n1520) );
  IV U518 ( .A(B[493]), .Z(n1521) );
  IV U519 ( .A(B[494]), .Z(n1522) );
  IV U520 ( .A(B[495]), .Z(n1523) );
  IV U521 ( .A(B[496]), .Z(n1524) );
  IV U522 ( .A(B[973]), .Z(n2001) );
  IV U523 ( .A(B[497]), .Z(n1525) );
  IV U524 ( .A(B[498]), .Z(n1526) );
  IV U525 ( .A(B[499]), .Z(n1527) );
  IV U526 ( .A(B[500]), .Z(n1528) );
  IV U527 ( .A(B[501]), .Z(n1529) );
  IV U528 ( .A(B[502]), .Z(n1530) );
  IV U529 ( .A(B[503]), .Z(n1531) );
  IV U530 ( .A(B[504]), .Z(n1532) );
  IV U531 ( .A(B[505]), .Z(n1533) );
  IV U532 ( .A(B[506]), .Z(n1534) );
  IV U533 ( .A(B[974]), .Z(n2002) );
  IV U534 ( .A(B[507]), .Z(n1535) );
  IV U535 ( .A(B[508]), .Z(n1536) );
  IV U536 ( .A(B[509]), .Z(n1537) );
  IV U537 ( .A(B[510]), .Z(n1538) );
  IV U538 ( .A(B[511]), .Z(n1539) );
  IV U539 ( .A(B[512]), .Z(n1540) );
  IV U540 ( .A(B[513]), .Z(n1541) );
  IV U541 ( .A(B[514]), .Z(n1542) );
  IV U542 ( .A(B[515]), .Z(n1543) );
  IV U543 ( .A(B[516]), .Z(n1544) );
  IV U544 ( .A(B[975]), .Z(n2003) );
  IV U545 ( .A(B[517]), .Z(n1545) );
  IV U546 ( .A(B[518]), .Z(n1546) );
  IV U547 ( .A(B[519]), .Z(n1547) );
  IV U548 ( .A(B[520]), .Z(n1548) );
  IV U549 ( .A(B[521]), .Z(n1549) );
  IV U550 ( .A(B[522]), .Z(n1550) );
  IV U551 ( .A(B[523]), .Z(n1551) );
  IV U552 ( .A(B[524]), .Z(n1552) );
  IV U553 ( .A(B[525]), .Z(n1553) );
  IV U554 ( .A(B[526]), .Z(n1554) );
  IV U555 ( .A(B[976]), .Z(n2004) );
  IV U556 ( .A(B[1021]), .Z(n2049) );
  IV U557 ( .A(B[527]), .Z(n1555) );
  IV U558 ( .A(B[528]), .Z(n1556) );
  IV U559 ( .A(B[529]), .Z(n1557) );
  IV U560 ( .A(B[530]), .Z(n1558) );
  IV U561 ( .A(B[531]), .Z(n1559) );
  IV U562 ( .A(B[532]), .Z(n1560) );
  IV U563 ( .A(B[533]), .Z(n1561) );
  IV U564 ( .A(B[534]), .Z(n1562) );
  IV U565 ( .A(B[535]), .Z(n1563) );
  IV U566 ( .A(B[536]), .Z(n1564) );
  IV U567 ( .A(B[977]), .Z(n2005) );
  IV U568 ( .A(B[537]), .Z(n1565) );
  IV U569 ( .A(B[538]), .Z(n1566) );
  IV U570 ( .A(B[539]), .Z(n1567) );
  IV U571 ( .A(B[540]), .Z(n1568) );
  IV U572 ( .A(B[541]), .Z(n1569) );
  IV U573 ( .A(B[542]), .Z(n1570) );
  IV U574 ( .A(B[543]), .Z(n1571) );
  IV U575 ( .A(B[544]), .Z(n1572) );
  IV U576 ( .A(B[545]), .Z(n1573) );
  IV U577 ( .A(B[546]), .Z(n1574) );
  IV U578 ( .A(B[978]), .Z(n2006) );
  IV U579 ( .A(B[547]), .Z(n1575) );
  IV U580 ( .A(B[548]), .Z(n1576) );
  IV U581 ( .A(B[549]), .Z(n1577) );
  IV U582 ( .A(B[550]), .Z(n1578) );
  IV U583 ( .A(B[551]), .Z(n1579) );
  IV U584 ( .A(B[552]), .Z(n1580) );
  IV U585 ( .A(B[553]), .Z(n1581) );
  IV U586 ( .A(B[554]), .Z(n1582) );
  IV U587 ( .A(B[555]), .Z(n1583) );
  IV U588 ( .A(B[556]), .Z(n1584) );
  IV U589 ( .A(B[979]), .Z(n2007) );
  IV U590 ( .A(B[557]), .Z(n1585) );
  IV U591 ( .A(B[558]), .Z(n1586) );
  IV U592 ( .A(B[559]), .Z(n1587) );
  IV U593 ( .A(B[560]), .Z(n1588) );
  IV U594 ( .A(B[561]), .Z(n1589) );
  IV U595 ( .A(B[562]), .Z(n1590) );
  IV U596 ( .A(B[563]), .Z(n1591) );
  IV U597 ( .A(B[564]), .Z(n1592) );
  IV U598 ( .A(B[565]), .Z(n1593) );
  IV U599 ( .A(B[566]), .Z(n1594) );
  IV U600 ( .A(B[980]), .Z(n2008) );
  IV U601 ( .A(B[567]), .Z(n1595) );
  IV U602 ( .A(B[568]), .Z(n1596) );
  IV U603 ( .A(B[569]), .Z(n1597) );
  IV U604 ( .A(B[570]), .Z(n1598) );
  IV U605 ( .A(B[571]), .Z(n1599) );
  IV U606 ( .A(B[572]), .Z(n1600) );
  IV U607 ( .A(B[573]), .Z(n1601) );
  IV U608 ( .A(B[574]), .Z(n1602) );
  IV U609 ( .A(B[575]), .Z(n1603) );
  IV U610 ( .A(B[576]), .Z(n1604) );
  IV U611 ( .A(B[981]), .Z(n2009) );
  IV U612 ( .A(B[577]), .Z(n1605) );
  IV U613 ( .A(B[578]), .Z(n1606) );
  IV U614 ( .A(B[579]), .Z(n1607) );
  IV U615 ( .A(B[580]), .Z(n1608) );
  IV U616 ( .A(B[581]), .Z(n1609) );
  IV U617 ( .A(B[582]), .Z(n1610) );
  IV U618 ( .A(B[583]), .Z(n1611) );
  IV U619 ( .A(B[584]), .Z(n1612) );
  IV U620 ( .A(B[585]), .Z(n1613) );
  IV U621 ( .A(B[586]), .Z(n1614) );
  IV U622 ( .A(B[982]), .Z(n2010) );
  IV U623 ( .A(B[587]), .Z(n1615) );
  IV U624 ( .A(B[588]), .Z(n1616) );
  IV U625 ( .A(B[589]), .Z(n1617) );
  IV U626 ( .A(B[590]), .Z(n1618) );
  IV U627 ( .A(B[591]), .Z(n1619) );
  IV U628 ( .A(B[592]), .Z(n1620) );
  IV U629 ( .A(B[593]), .Z(n1621) );
  IV U630 ( .A(B[594]), .Z(n1622) );
  IV U631 ( .A(B[595]), .Z(n1623) );
  IV U632 ( .A(B[596]), .Z(n1624) );
  IV U633 ( .A(B[983]), .Z(n2011) );
  IV U634 ( .A(B[597]), .Z(n1625) );
  IV U635 ( .A(B[598]), .Z(n1626) );
  IV U636 ( .A(B[599]), .Z(n1627) );
  IV U637 ( .A(B[600]), .Z(n1628) );
  IV U638 ( .A(B[601]), .Z(n1629) );
  IV U639 ( .A(B[602]), .Z(n1630) );
  IV U640 ( .A(B[603]), .Z(n1631) );
  IV U641 ( .A(B[604]), .Z(n1632) );
  IV U642 ( .A(B[605]), .Z(n1633) );
  IV U643 ( .A(B[606]), .Z(n1634) );
  IV U644 ( .A(B[984]), .Z(n2012) );
  IV U645 ( .A(B[607]), .Z(n1635) );
  IV U646 ( .A(B[608]), .Z(n1636) );
  IV U647 ( .A(B[609]), .Z(n1637) );
  IV U648 ( .A(B[610]), .Z(n1638) );
  IV U649 ( .A(B[611]), .Z(n1639) );
  IV U650 ( .A(B[612]), .Z(n1640) );
  IV U651 ( .A(B[613]), .Z(n1641) );
  IV U652 ( .A(B[614]), .Z(n1642) );
  IV U653 ( .A(B[615]), .Z(n1643) );
  IV U654 ( .A(B[616]), .Z(n1644) );
  IV U655 ( .A(B[985]), .Z(n2013) );
  IV U656 ( .A(B[617]), .Z(n1645) );
  IV U657 ( .A(B[618]), .Z(n1646) );
  IV U658 ( .A(B[619]), .Z(n1647) );
  IV U659 ( .A(B[620]), .Z(n1648) );
  IV U660 ( .A(B[621]), .Z(n1649) );
  IV U661 ( .A(B[622]), .Z(n1650) );
  IV U662 ( .A(B[623]), .Z(n1651) );
  IV U663 ( .A(B[624]), .Z(n1652) );
  IV U664 ( .A(B[625]), .Z(n1653) );
  IV U665 ( .A(B[626]), .Z(n1654) );
  IV U666 ( .A(B[986]), .Z(n2014) );
  IV U667 ( .A(B[1022]), .Z(n2050) );
  IV U668 ( .A(B[627]), .Z(n1655) );
  IV U669 ( .A(B[628]), .Z(n1656) );
  IV U670 ( .A(B[629]), .Z(n1657) );
  IV U671 ( .A(B[630]), .Z(n1658) );
  IV U672 ( .A(B[631]), .Z(n1659) );
  IV U673 ( .A(B[632]), .Z(n1660) );
  IV U674 ( .A(B[633]), .Z(n1661) );
  IV U675 ( .A(B[634]), .Z(n1662) );
  IV U676 ( .A(B[635]), .Z(n1663) );
  IV U677 ( .A(B[636]), .Z(n1664) );
  IV U678 ( .A(B[987]), .Z(n2015) );
  IV U679 ( .A(B[637]), .Z(n1665) );
  IV U680 ( .A(B[638]), .Z(n1666) );
  IV U681 ( .A(B[639]), .Z(n1667) );
  IV U682 ( .A(B[640]), .Z(n1668) );
  IV U683 ( .A(B[641]), .Z(n1669) );
  IV U684 ( .A(B[642]), .Z(n1670) );
  IV U685 ( .A(B[643]), .Z(n1671) );
  IV U686 ( .A(B[644]), .Z(n1672) );
  IV U687 ( .A(B[645]), .Z(n1673) );
  IV U688 ( .A(B[646]), .Z(n1674) );
  IV U689 ( .A(B[988]), .Z(n2016) );
  IV U690 ( .A(B[647]), .Z(n1675) );
  IV U691 ( .A(B[648]), .Z(n1676) );
  IV U692 ( .A(B[649]), .Z(n1677) );
  IV U693 ( .A(B[650]), .Z(n1678) );
  IV U694 ( .A(B[651]), .Z(n1679) );
  IV U695 ( .A(B[652]), .Z(n1680) );
  IV U696 ( .A(B[653]), .Z(n1681) );
  IV U697 ( .A(B[654]), .Z(n1682) );
  IV U698 ( .A(B[655]), .Z(n1683) );
  IV U699 ( .A(B[656]), .Z(n1684) );
  IV U700 ( .A(B[989]), .Z(n2017) );
  IV U701 ( .A(B[657]), .Z(n1685) );
  IV U702 ( .A(B[658]), .Z(n1686) );
  IV U703 ( .A(B[659]), .Z(n1687) );
  IV U704 ( .A(B[660]), .Z(n1688) );
  IV U705 ( .A(B[661]), .Z(n1689) );
  IV U706 ( .A(B[662]), .Z(n1690) );
  IV U707 ( .A(B[663]), .Z(n1691) );
  IV U708 ( .A(B[664]), .Z(n1692) );
  IV U709 ( .A(B[665]), .Z(n1693) );
  IV U710 ( .A(B[666]), .Z(n1694) );
  IV U711 ( .A(B[990]), .Z(n2018) );
  IV U712 ( .A(B[667]), .Z(n1695) );
  IV U713 ( .A(B[668]), .Z(n1696) );
  IV U714 ( .A(B[669]), .Z(n1697) );
  IV U715 ( .A(B[670]), .Z(n1698) );
  IV U716 ( .A(B[671]), .Z(n1699) );
  IV U717 ( .A(B[672]), .Z(n1700) );
  IV U718 ( .A(B[673]), .Z(n1701) );
  IV U719 ( .A(B[674]), .Z(n1702) );
  IV U720 ( .A(B[675]), .Z(n1703) );
  IV U721 ( .A(B[676]), .Z(n1704) );
  IV U722 ( .A(B[991]), .Z(n2019) );
  IV U723 ( .A(B[677]), .Z(n1705) );
  IV U724 ( .A(B[678]), .Z(n1706) );
  IV U725 ( .A(B[679]), .Z(n1707) );
  IV U726 ( .A(B[680]), .Z(n1708) );
  IV U727 ( .A(B[681]), .Z(n1709) );
  IV U728 ( .A(B[682]), .Z(n1710) );
  IV U729 ( .A(B[683]), .Z(n1711) );
  IV U730 ( .A(B[684]), .Z(n1712) );
  IV U731 ( .A(B[685]), .Z(n1713) );
  IV U732 ( .A(B[686]), .Z(n1714) );
  IV U733 ( .A(B[992]), .Z(n2020) );
  IV U734 ( .A(B[687]), .Z(n1715) );
  IV U735 ( .A(B[688]), .Z(n1716) );
  IV U736 ( .A(B[689]), .Z(n1717) );
  IV U737 ( .A(B[690]), .Z(n1718) );
  IV U738 ( .A(B[691]), .Z(n1719) );
  IV U739 ( .A(B[692]), .Z(n1720) );
  IV U740 ( .A(B[693]), .Z(n1721) );
  IV U741 ( .A(B[694]), .Z(n1722) );
  IV U742 ( .A(B[695]), .Z(n1723) );
  IV U743 ( .A(B[696]), .Z(n1724) );
  IV U744 ( .A(B[993]), .Z(n2021) );
  IV U745 ( .A(B[697]), .Z(n1725) );
  IV U746 ( .A(B[698]), .Z(n1726) );
  IV U747 ( .A(B[699]), .Z(n1727) );
  IV U748 ( .A(B[700]), .Z(n1728) );
  IV U749 ( .A(B[701]), .Z(n1729) );
  IV U750 ( .A(B[702]), .Z(n1730) );
  IV U751 ( .A(B[703]), .Z(n1731) );
  IV U752 ( .A(B[704]), .Z(n1732) );
  IV U753 ( .A(B[705]), .Z(n1733) );
  IV U754 ( .A(B[706]), .Z(n1734) );
  IV U755 ( .A(B[994]), .Z(n2022) );
  IV U756 ( .A(B[707]), .Z(n1735) );
  IV U757 ( .A(B[708]), .Z(n1736) );
  IV U758 ( .A(B[709]), .Z(n1737) );
  IV U759 ( .A(B[710]), .Z(n1738) );
  IV U760 ( .A(B[711]), .Z(n1739) );
  IV U761 ( .A(B[712]), .Z(n1740) );
  IV U762 ( .A(B[713]), .Z(n1741) );
  IV U763 ( .A(B[714]), .Z(n1742) );
  IV U764 ( .A(B[715]), .Z(n1743) );
  IV U765 ( .A(B[716]), .Z(n1744) );
  IV U766 ( .A(B[995]), .Z(n2023) );
  IV U767 ( .A(B[717]), .Z(n1745) );
  IV U768 ( .A(B[718]), .Z(n1746) );
  IV U769 ( .A(B[719]), .Z(n1747) );
  IV U770 ( .A(B[720]), .Z(n1748) );
  IV U771 ( .A(B[721]), .Z(n1749) );
  IV U772 ( .A(B[722]), .Z(n1750) );
  IV U773 ( .A(B[723]), .Z(n1751) );
  IV U774 ( .A(B[724]), .Z(n1752) );
  IV U775 ( .A(B[725]), .Z(n1753) );
  IV U776 ( .A(B[726]), .Z(n1754) );
  IV U777 ( .A(B[996]), .Z(n2024) );
  IV U778 ( .A(B[1023]), .Z(n2051) );
  IV U779 ( .A(B[727]), .Z(n1755) );
  IV U780 ( .A(B[728]), .Z(n1756) );
  IV U781 ( .A(B[729]), .Z(n1757) );
  IV U782 ( .A(B[730]), .Z(n1758) );
  IV U783 ( .A(B[731]), .Z(n1759) );
  IV U784 ( .A(B[732]), .Z(n1760) );
  IV U785 ( .A(B[733]), .Z(n1761) );
  IV U786 ( .A(B[734]), .Z(n1762) );
  IV U787 ( .A(B[735]), .Z(n1763) );
  IV U788 ( .A(B[736]), .Z(n1764) );
  IV U789 ( .A(B[997]), .Z(n2025) );
  IV U790 ( .A(B[737]), .Z(n1765) );
  IV U791 ( .A(B[738]), .Z(n1766) );
  IV U792 ( .A(B[739]), .Z(n1767) );
  IV U793 ( .A(B[740]), .Z(n1768) );
  IV U794 ( .A(B[741]), .Z(n1769) );
  IV U795 ( .A(B[742]), .Z(n1770) );
  IV U796 ( .A(B[743]), .Z(n1771) );
  IV U797 ( .A(B[744]), .Z(n1772) );
  IV U798 ( .A(B[745]), .Z(n1773) );
  IV U799 ( .A(B[746]), .Z(n1774) );
  IV U800 ( .A(B[998]), .Z(n2026) );
  IV U801 ( .A(B[747]), .Z(n1775) );
  IV U802 ( .A(B[748]), .Z(n1776) );
  IV U803 ( .A(B[749]), .Z(n1777) );
  IV U804 ( .A(B[750]), .Z(n1778) );
  IV U805 ( .A(B[751]), .Z(n1779) );
  IV U806 ( .A(B[752]), .Z(n1780) );
  IV U807 ( .A(B[753]), .Z(n1781) );
  IV U808 ( .A(B[754]), .Z(n1782) );
  IV U809 ( .A(B[755]), .Z(n1783) );
  IV U810 ( .A(B[756]), .Z(n1784) );
  IV U811 ( .A(B[999]), .Z(n2027) );
  IV U812 ( .A(B[757]), .Z(n1785) );
  IV U813 ( .A(B[758]), .Z(n1786) );
  IV U814 ( .A(B[759]), .Z(n1787) );
  IV U815 ( .A(B[760]), .Z(n1788) );
  IV U816 ( .A(B[761]), .Z(n1789) );
  IV U817 ( .A(B[762]), .Z(n1790) );
  IV U818 ( .A(B[763]), .Z(n1791) );
  IV U819 ( .A(B[764]), .Z(n1792) );
  IV U820 ( .A(B[765]), .Z(n1793) );
  IV U821 ( .A(B[766]), .Z(n1794) );
  IV U822 ( .A(B[1000]), .Z(n2028) );
  IV U823 ( .A(B[767]), .Z(n1795) );
  IV U824 ( .A(B[768]), .Z(n1796) );
  IV U825 ( .A(B[769]), .Z(n1797) );
  IV U826 ( .A(B[770]), .Z(n1798) );
  IV U827 ( .A(B[771]), .Z(n1799) );
  IV U828 ( .A(B[772]), .Z(n1800) );
  IV U829 ( .A(B[773]), .Z(n1801) );
  IV U830 ( .A(B[774]), .Z(n1802) );
  IV U831 ( .A(B[775]), .Z(n1803) );
  IV U832 ( .A(B[776]), .Z(n1804) );
  IV U833 ( .A(B[1001]), .Z(n2029) );
  IV U834 ( .A(B[777]), .Z(n1805) );
  IV U835 ( .A(B[778]), .Z(n1806) );
  IV U836 ( .A(B[779]), .Z(n1807) );
  IV U837 ( .A(B[780]), .Z(n1808) );
  IV U838 ( .A(B[781]), .Z(n1809) );
  IV U839 ( .A(B[782]), .Z(n1810) );
  IV U840 ( .A(B[783]), .Z(n1811) );
  IV U841 ( .A(B[784]), .Z(n1812) );
  IV U842 ( .A(B[785]), .Z(n1813) );
  IV U843 ( .A(B[786]), .Z(n1814) );
  IV U844 ( .A(B[1002]), .Z(n2030) );
  IV U845 ( .A(B[787]), .Z(n1815) );
  IV U846 ( .A(B[788]), .Z(n1816) );
  IV U847 ( .A(B[789]), .Z(n1817) );
  IV U848 ( .A(B[790]), .Z(n1818) );
  IV U849 ( .A(B[791]), .Z(n1819) );
  IV U850 ( .A(B[792]), .Z(n1820) );
  IV U851 ( .A(B[793]), .Z(n1821) );
  IV U852 ( .A(B[794]), .Z(n1822) );
  IV U853 ( .A(B[795]), .Z(n1823) );
  IV U854 ( .A(B[796]), .Z(n1824) );
  IV U855 ( .A(B[1003]), .Z(n2031) );
  IV U856 ( .A(B[797]), .Z(n1825) );
  IV U857 ( .A(B[798]), .Z(n1826) );
  IV U858 ( .A(B[799]), .Z(n1827) );
  IV U859 ( .A(B[800]), .Z(n1828) );
  IV U860 ( .A(B[801]), .Z(n1829) );
  IV U861 ( .A(B[802]), .Z(n1830) );
  IV U862 ( .A(B[803]), .Z(n1831) );
  IV U863 ( .A(B[804]), .Z(n1832) );
  IV U864 ( .A(B[805]), .Z(n1833) );
  IV U865 ( .A(B[806]), .Z(n1834) );
  IV U866 ( .A(B[1004]), .Z(n2032) );
  IV U867 ( .A(B[807]), .Z(n1835) );
  IV U868 ( .A(B[808]), .Z(n1836) );
  IV U869 ( .A(B[809]), .Z(n1837) );
  IV U870 ( .A(B[810]), .Z(n1838) );
  IV U871 ( .A(B[811]), .Z(n1839) );
  IV U872 ( .A(B[812]), .Z(n1840) );
  IV U873 ( .A(B[813]), .Z(n1841) );
  IV U874 ( .A(B[814]), .Z(n1842) );
  IV U875 ( .A(B[815]), .Z(n1843) );
  IV U876 ( .A(B[816]), .Z(n1844) );
  IV U877 ( .A(B[1005]), .Z(n2033) );
  IV U878 ( .A(B[817]), .Z(n1845) );
  IV U879 ( .A(B[818]), .Z(n1846) );
  IV U880 ( .A(B[819]), .Z(n1847) );
  IV U881 ( .A(B[820]), .Z(n1848) );
  IV U882 ( .A(B[821]), .Z(n1849) );
  IV U883 ( .A(B[822]), .Z(n1850) );
  IV U884 ( .A(B[823]), .Z(n1851) );
  IV U885 ( .A(B[824]), .Z(n1852) );
  IV U886 ( .A(B[825]), .Z(n1853) );
  IV U887 ( .A(B[826]), .Z(n1854) );
  IV U888 ( .A(B[1006]), .Z(n2034) );
  IV U889 ( .A(B[1024]), .Z(n2052) );
  IV U890 ( .A(B[827]), .Z(n1855) );
  IV U891 ( .A(B[828]), .Z(n1856) );
  IV U892 ( .A(B[829]), .Z(n1857) );
  IV U893 ( .A(B[830]), .Z(n1858) );
  IV U894 ( .A(B[831]), .Z(n1859) );
  IV U895 ( .A(B[832]), .Z(n1860) );
  IV U896 ( .A(B[833]), .Z(n1861) );
  IV U897 ( .A(B[834]), .Z(n1862) );
  IV U898 ( .A(B[835]), .Z(n1863) );
  IV U899 ( .A(B[836]), .Z(n1864) );
  IV U900 ( .A(B[1007]), .Z(n2035) );
  IV U901 ( .A(B[837]), .Z(n1865) );
  IV U902 ( .A(B[838]), .Z(n1866) );
  IV U903 ( .A(B[839]), .Z(n1867) );
  IV U904 ( .A(B[840]), .Z(n1868) );
  IV U905 ( .A(B[841]), .Z(n1869) );
  IV U906 ( .A(B[842]), .Z(n1870) );
  IV U907 ( .A(B[843]), .Z(n1871) );
  IV U908 ( .A(B[844]), .Z(n1872) );
  IV U909 ( .A(B[845]), .Z(n1873) );
  IV U910 ( .A(B[846]), .Z(n1874) );
  IV U911 ( .A(B[1008]), .Z(n2036) );
  IV U912 ( .A(B[847]), .Z(n1875) );
  IV U913 ( .A(B[848]), .Z(n1876) );
  IV U914 ( .A(B[849]), .Z(n1877) );
  IV U915 ( .A(B[850]), .Z(n1878) );
  IV U916 ( .A(B[851]), .Z(n1879) );
  IV U917 ( .A(B[852]), .Z(n1880) );
  IV U918 ( .A(B[853]), .Z(n1881) );
  IV U919 ( .A(B[854]), .Z(n1882) );
  IV U920 ( .A(B[855]), .Z(n1883) );
  IV U921 ( .A(B[856]), .Z(n1884) );
  IV U922 ( .A(B[1009]), .Z(n2037) );
  IV U923 ( .A(B[857]), .Z(n1885) );
  IV U924 ( .A(B[858]), .Z(n1886) );
  IV U925 ( .A(B[859]), .Z(n1887) );
  IV U926 ( .A(B[860]), .Z(n1888) );
  IV U927 ( .A(B[861]), .Z(n1889) );
  IV U928 ( .A(B[862]), .Z(n1890) );
  IV U929 ( .A(B[863]), .Z(n1891) );
  IV U930 ( .A(B[864]), .Z(n1892) );
  IV U931 ( .A(B[865]), .Z(n1893) );
  IV U932 ( .A(B[866]), .Z(n1894) );
  IV U933 ( .A(B[1010]), .Z(n2038) );
  IV U934 ( .A(B[867]), .Z(n1895) );
  IV U935 ( .A(B[868]), .Z(n1896) );
  IV U936 ( .A(B[869]), .Z(n1897) );
  IV U937 ( .A(B[870]), .Z(n1898) );
  IV U938 ( .A(B[871]), .Z(n1899) );
  IV U939 ( .A(B[872]), .Z(n1900) );
  IV U940 ( .A(B[873]), .Z(n1901) );
  IV U941 ( .A(B[874]), .Z(n1902) );
  IV U942 ( .A(B[875]), .Z(n1903) );
  IV U943 ( .A(B[876]), .Z(n1904) );
  IV U944 ( .A(B[1011]), .Z(n2039) );
  IV U945 ( .A(B[877]), .Z(n1905) );
  IV U946 ( .A(B[878]), .Z(n1906) );
  IV U947 ( .A(B[879]), .Z(n1907) );
  IV U948 ( .A(B[880]), .Z(n1908) );
  IV U949 ( .A(B[881]), .Z(n1909) );
  IV U950 ( .A(B[882]), .Z(n1910) );
  IV U951 ( .A(B[883]), .Z(n1911) );
  IV U952 ( .A(B[884]), .Z(n1912) );
  IV U953 ( .A(B[885]), .Z(n1913) );
  IV U954 ( .A(B[886]), .Z(n1914) );
  IV U955 ( .A(B[1012]), .Z(n2040) );
  IV U956 ( .A(B[887]), .Z(n1915) );
  IV U957 ( .A(B[888]), .Z(n1916) );
  IV U958 ( .A(B[889]), .Z(n1917) );
  IV U959 ( .A(B[890]), .Z(n1918) );
  IV U960 ( .A(B[891]), .Z(n1919) );
  IV U961 ( .A(B[892]), .Z(n1920) );
  IV U962 ( .A(B[893]), .Z(n1921) );
  IV U963 ( .A(B[894]), .Z(n1922) );
  IV U964 ( .A(B[895]), .Z(n1923) );
  IV U965 ( .A(B[896]), .Z(n1924) );
  IV U966 ( .A(B[1013]), .Z(n2041) );
  IV U967 ( .A(B[897]), .Z(n1925) );
  IV U968 ( .A(B[898]), .Z(n1926) );
  IV U969 ( .A(B[899]), .Z(n1927) );
  IV U970 ( .A(B[900]), .Z(n1928) );
  IV U971 ( .A(B[901]), .Z(n1929) );
  IV U972 ( .A(B[902]), .Z(n1930) );
  IV U973 ( .A(B[903]), .Z(n1931) );
  IV U974 ( .A(B[904]), .Z(n1932) );
  IV U975 ( .A(B[905]), .Z(n1933) );
  IV U976 ( .A(B[906]), .Z(n1934) );
  IV U977 ( .A(B[1014]), .Z(n2042) );
  IV U978 ( .A(B[907]), .Z(n1935) );
  IV U979 ( .A(B[908]), .Z(n1936) );
  IV U980 ( .A(B[909]), .Z(n1937) );
  IV U981 ( .A(B[910]), .Z(n1938) );
  IV U982 ( .A(B[911]), .Z(n1939) );
  IV U983 ( .A(B[912]), .Z(n1940) );
  IV U984 ( .A(B[913]), .Z(n1941) );
  IV U985 ( .A(B[914]), .Z(n1942) );
  IV U986 ( .A(B[915]), .Z(n1943) );
  IV U987 ( .A(B[916]), .Z(n1944) );
  IV U988 ( .A(B[1015]), .Z(n2043) );
  IV U989 ( .A(B[917]), .Z(n1945) );
  IV U990 ( .A(B[918]), .Z(n1946) );
  IV U991 ( .A(B[919]), .Z(n1947) );
  IV U992 ( .A(B[920]), .Z(n1948) );
  IV U993 ( .A(B[921]), .Z(n1949) );
  IV U994 ( .A(B[922]), .Z(n1950) );
  IV U995 ( .A(B[923]), .Z(n1951) );
  IV U996 ( .A(B[0]), .Z(n1028) );
  IV U997 ( .A(B[1]), .Z(n1029) );
  IV U998 ( .A(B[2]), .Z(n1030) );
  IV U999 ( .A(B[3]), .Z(n1031) );
  IV U1000 ( .A(B[4]), .Z(n1032) );
  IV U1001 ( .A(B[5]), .Z(n1033) );
  IV U1002 ( .A(B[6]), .Z(n1034) );
  IV U1003 ( .A(B[924]), .Z(n1952) );
  IV U1004 ( .A(B[7]), .Z(n1035) );
  IV U1005 ( .A(B[8]), .Z(n1036) );
  IV U1006 ( .A(B[9]), .Z(n1037) );
  IV U1007 ( .A(B[10]), .Z(n1038) );
  IV U1008 ( .A(B[11]), .Z(n1039) );
  IV U1009 ( .A(B[12]), .Z(n1040) );
  IV U1010 ( .A(B[13]), .Z(n1041) );
  IV U1011 ( .A(B[14]), .Z(n1042) );
  IV U1012 ( .A(B[15]), .Z(n1043) );
  IV U1013 ( .A(B[16]), .Z(n1044) );
  IV U1014 ( .A(B[925]), .Z(n1953) );
  IV U1015 ( .A(B[17]), .Z(n1045) );
  IV U1016 ( .A(B[18]), .Z(n1046) );
  IV U1017 ( .A(B[19]), .Z(n1047) );
  IV U1018 ( .A(B[20]), .Z(n1048) );
  IV U1019 ( .A(B[21]), .Z(n1049) );
  IV U1020 ( .A(B[22]), .Z(n1050) );
  IV U1021 ( .A(B[23]), .Z(n1051) );
  IV U1022 ( .A(B[24]), .Z(n1052) );
  IV U1023 ( .A(B[25]), .Z(n1053) );
  IV U1024 ( .A(B[26]), .Z(n1054) );
  IV U1025 ( .A(B[926]), .Z(n1954) );
  IV U1026 ( .A(B[1016]), .Z(n2044) );
  IV U1027 ( .A(B[1025]), .Z(n2053) );
endmodule


module FA_11576 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XNOR U1 ( .A(CI), .B(A), .Z(S) );
endmodule


module FA_11577 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11578 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11579 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11580 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11581 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11582 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11583 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11584 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11585 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11586 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11587 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11588 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11589 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11590 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11591 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11592 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11593 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11594 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11595 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11596 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11597 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11598 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11599 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11600 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11601 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11602 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11603 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11604 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11605 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11606 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11607 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11608 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11609 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11610 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11611 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11612 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11613 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11614 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11615 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11616 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11617 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11618 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11619 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11620 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11621 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11622 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11623 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11624 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11625 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11626 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11627 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11628 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11629 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11630 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11631 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11632 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11633 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11634 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11635 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11636 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11637 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11638 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11639 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11640 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11641 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11642 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11643 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11644 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11645 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11646 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11647 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11648 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11649 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11650 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11651 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11652 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11653 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11654 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11655 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11656 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11657 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11658 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11659 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11660 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11661 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11662 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11663 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11664 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11665 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11666 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11667 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11668 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11669 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11670 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11671 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11672 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11673 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11674 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11675 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11676 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11677 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11678 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11679 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11680 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11681 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11682 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11683 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11684 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11685 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11686 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11687 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11688 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11689 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11690 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11691 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11692 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11693 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11694 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11695 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11696 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11697 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11698 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11699 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11700 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11701 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11702 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11703 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11704 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11705 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11706 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11707 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11708 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11709 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11710 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11711 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11712 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11713 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11714 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11715 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11716 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11717 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11718 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11719 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11720 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11721 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11722 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11723 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11724 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11725 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11726 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11727 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11728 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11729 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11730 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11731 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11732 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11733 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11734 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11735 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11736 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11737 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11738 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11739 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11740 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11741 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11742 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11743 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11744 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11745 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11746 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11747 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11748 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11749 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11750 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11751 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11752 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11753 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11754 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11755 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11756 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11757 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11758 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11759 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11760 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11761 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11762 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11763 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11764 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11765 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11766 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11767 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11768 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11769 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11770 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11771 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11772 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11773 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11774 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11775 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11776 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11777 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11778 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11779 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11780 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11781 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11782 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11783 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11784 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11785 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11786 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11787 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11788 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11789 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11790 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11791 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11792 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11793 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11794 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11795 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11796 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11797 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11798 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11799 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11800 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11801 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11802 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11803 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11804 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11805 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11806 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11807 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11808 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11809 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11810 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11811 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11812 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11813 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11814 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11815 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11816 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11817 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11818 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11819 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11820 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11821 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11822 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11823 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11824 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11825 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11826 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11827 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11828 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11829 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11830 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11831 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11832 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11833 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11834 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11835 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11836 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11837 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11838 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11839 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11840 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11841 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11842 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11843 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11844 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11845 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11846 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11847 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11848 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11849 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11850 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11851 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11852 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11853 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11854 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11855 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11856 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11857 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11858 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11859 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11860 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11861 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11862 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11863 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11864 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11865 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11866 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11867 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11868 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11869 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11870 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11871 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11872 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11873 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11874 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11875 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11876 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11877 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11878 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11879 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11880 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11881 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11882 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11883 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11884 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11885 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11886 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11887 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11888 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11889 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11890 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11891 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11892 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11893 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11894 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11895 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11896 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11897 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11898 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11899 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11900 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11901 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11902 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11903 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11904 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11905 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11906 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11907 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11908 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11909 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11910 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11911 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11912 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11913 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11914 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11915 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11916 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11917 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11918 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11919 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11920 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11921 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11922 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11923 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11924 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11925 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11926 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11927 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11928 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11929 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11930 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11931 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11932 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11933 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11934 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11935 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11936 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11937 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11938 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11939 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11940 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11941 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11942 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11943 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11944 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11945 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11946 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11947 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11948 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11949 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11950 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11951 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11952 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11953 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11954 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11955 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11956 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11957 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11958 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11959 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11960 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11961 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11962 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11963 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11964 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11965 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11966 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11967 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11968 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11969 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11970 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11971 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11972 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11973 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11974 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11975 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11976 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11977 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11978 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11979 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11980 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11981 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11982 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11983 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11984 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11985 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11986 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11987 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11988 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11989 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11990 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11991 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11992 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11993 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11994 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11995 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11996 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11997 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11998 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11999 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12000 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12001 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12002 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12003 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12004 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12005 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12006 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12007 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12008 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12009 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12010 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12011 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12012 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12013 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12014 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12015 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12016 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12017 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12018 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12019 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12020 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12021 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12022 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12023 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12024 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12025 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12026 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12027 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12028 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12029 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12030 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12031 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12032 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12033 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12034 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12035 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12036 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12037 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12038 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12039 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12040 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12041 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12042 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12043 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12044 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12045 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12046 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12047 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12048 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12049 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12050 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12051 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12052 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12053 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12054 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12055 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12056 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12057 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12058 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12059 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12060 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12061 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12062 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12063 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12064 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12065 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12066 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12067 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12068 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12069 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12070 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12071 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12072 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12073 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12074 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12075 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12076 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12077 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12078 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12079 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12080 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12081 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12082 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12083 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12084 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12085 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12086 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12087 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12088 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12089 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12090 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12091 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12092 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12093 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12094 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12095 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12096 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12097 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12098 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12099 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12100 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12101 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12102 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12103 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12104 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12105 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12106 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12107 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12108 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12109 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12110 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12111 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12112 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12113 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12114 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12115 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12116 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12117 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12118 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12119 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12120 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12121 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12122 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12123 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12124 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12125 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12126 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12127 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12128 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12129 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12130 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12131 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12132 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12133 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12134 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12135 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12136 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12137 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12138 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12139 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12140 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12141 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12142 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12143 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12144 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12145 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12146 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12147 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12148 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12149 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12150 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12151 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12152 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12153 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12154 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12155 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12156 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12157 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12158 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12159 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12160 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12161 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12162 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12163 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12164 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12165 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12166 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12167 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12168 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12169 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12170 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12171 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12172 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12173 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12174 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12175 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12176 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12177 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12178 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12179 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12180 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12181 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12182 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12183 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12184 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12185 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12186 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12187 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12188 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12189 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12190 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12191 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12192 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12193 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12194 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12195 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12196 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12197 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12198 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12199 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12200 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12201 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12202 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12203 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12204 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12205 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12206 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12207 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12208 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12209 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12210 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12211 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12212 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12213 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12214 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12215 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12216 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12217 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12218 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12219 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12220 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12221 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12222 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12223 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12224 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12225 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12226 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12227 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12228 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12229 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12230 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12231 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12232 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12233 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12234 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12235 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12236 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12237 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12238 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12239 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12240 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12241 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12242 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12243 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12244 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12245 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12246 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12247 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12248 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12249 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12250 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12251 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12252 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12253 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12254 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12255 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12256 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12257 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12258 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12259 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12260 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12261 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12262 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12263 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12264 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12265 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12266 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12267 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12268 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12269 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12270 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12271 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12272 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12273 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12274 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12275 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12276 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12277 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12278 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12279 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12280 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12281 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12282 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12283 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12284 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12285 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12286 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12287 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12288 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12289 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12290 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12291 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12292 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12293 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12294 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12295 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12296 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12297 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12298 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12299 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12300 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12301 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12302 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12303 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12304 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12305 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12306 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12307 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12308 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12309 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12310 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12311 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12312 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12313 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12314 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12315 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12316 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12317 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12318 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12319 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12320 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12321 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12322 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12323 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12324 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12325 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12326 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12327 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12328 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12329 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12330 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12331 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12332 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12333 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12334 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12335 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12336 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12337 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12338 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12339 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12340 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12341 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12342 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12343 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12344 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12345 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12346 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12347 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12348 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12349 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12350 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12351 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12352 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12353 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12354 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12355 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12356 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12357 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12358 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12359 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12360 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12361 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12362 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12363 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12364 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12365 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12366 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12367 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12368 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12369 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12370 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12371 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12372 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12373 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12374 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12375 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12376 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12377 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12378 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12379 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12380 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12381 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12382 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12383 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12384 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12385 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12386 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12387 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12388 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12389 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12390 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12391 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12392 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12393 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12394 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12395 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12396 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12397 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12398 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12399 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12400 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12401 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12402 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12403 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12404 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12405 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12406 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12407 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12408 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12409 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12410 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12411 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12412 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12413 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12414 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12415 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12416 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12417 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12418 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12419 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12420 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12421 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12422 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12423 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12424 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12425 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12426 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12427 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12428 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12429 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12430 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12431 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12432 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12433 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12434 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12435 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12436 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12437 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12438 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12439 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12440 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12441 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12442 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12443 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12444 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12445 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12446 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12447 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12448 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12449 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12450 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12451 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12452 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12453 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12454 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12455 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12456 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12457 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12458 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12459 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12460 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12461 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12462 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12463 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12464 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12465 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12466 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12467 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12468 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12469 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12470 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12471 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12472 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12473 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12474 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12475 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12476 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12477 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12478 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12479 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12480 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12481 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12482 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12483 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12484 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12485 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12486 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12487 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12488 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12489 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12490 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12491 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12492 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12493 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12494 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12495 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12496 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12497 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12498 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12499 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12500 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12501 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12502 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12503 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12504 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12505 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12506 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12507 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12508 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12509 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12510 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12511 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12512 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12513 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12514 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12515 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12516 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12517 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12518 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12519 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12520 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12521 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12522 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12523 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12524 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12525 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12526 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12527 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12528 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12529 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12530 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12531 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12532 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12533 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12534 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12535 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12536 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12537 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12538 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12539 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12540 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12541 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12542 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12543 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12544 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12545 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12546 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12547 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12548 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12549 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12550 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12551 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12552 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12553 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12554 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12555 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12556 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12557 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12558 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12559 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12560 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12561 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12562 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12563 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12564 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12565 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12566 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12567 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12568 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12569 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12570 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12571 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12572 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12573 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12574 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12575 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12576 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12577 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12578 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12579 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12580 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12581 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12582 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12583 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12584 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12585 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12586 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12587 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12588 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12589 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12590 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12591 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12592 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12593 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12594 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12595 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12596 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12597 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12598 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12599 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12600 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XNOR U1 ( .A(B), .B(A), .Z(S) );
  OR U2 ( .A(B), .B(A), .Z(CO) );
endmodule


module SUB_N1026_1 ( A, B, S, CO );
  input [1025:0] A;
  input [1025:0] B;
  output [1025:0] S;
  output CO;
  wire   n2, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048;
  wire   [1025:1] C;

  FA_12600 \FA_INST_0[0].FA_INST_1[0].FA_  ( .A(A[0]), .B(n2), .CI(1'b1), .S(
        S[0]), .CO(C[1]) );
  FA_12599 \FA_INST_0[0].FA_INST_1[1].FA_  ( .A(A[1]), .B(n1026), .CI(C[1]), 
        .S(S[1]), .CO(C[2]) );
  FA_12598 \FA_INST_0[0].FA_INST_1[2].FA_  ( .A(A[2]), .B(n1027), .CI(C[2]), 
        .S(S[2]), .CO(C[3]) );
  FA_12597 \FA_INST_0[0].FA_INST_1[3].FA_  ( .A(A[3]), .B(n1028), .CI(C[3]), 
        .S(S[3]), .CO(C[4]) );
  FA_12596 \FA_INST_0[0].FA_INST_1[4].FA_  ( .A(A[4]), .B(n1029), .CI(C[4]), 
        .S(S[4]), .CO(C[5]) );
  FA_12595 \FA_INST_0[0].FA_INST_1[5].FA_  ( .A(A[5]), .B(n1030), .CI(C[5]), 
        .S(S[5]), .CO(C[6]) );
  FA_12594 \FA_INST_0[0].FA_INST_1[6].FA_  ( .A(A[6]), .B(n1031), .CI(C[6]), 
        .S(S[6]), .CO(C[7]) );
  FA_12593 \FA_INST_0[0].FA_INST_1[7].FA_  ( .A(A[7]), .B(n1032), .CI(C[7]), 
        .S(S[7]), .CO(C[8]) );
  FA_12592 \FA_INST_0[0].FA_INST_1[8].FA_  ( .A(A[8]), .B(n1033), .CI(C[8]), 
        .S(S[8]), .CO(C[9]) );
  FA_12591 \FA_INST_0[0].FA_INST_1[9].FA_  ( .A(A[9]), .B(n1034), .CI(C[9]), 
        .S(S[9]), .CO(C[10]) );
  FA_12590 \FA_INST_0[0].FA_INST_1[10].FA_  ( .A(A[10]), .B(n1035), .CI(C[10]), 
        .S(S[10]), .CO(C[11]) );
  FA_12589 \FA_INST_0[0].FA_INST_1[11].FA_  ( .A(A[11]), .B(n1036), .CI(C[11]), 
        .S(S[11]), .CO(C[12]) );
  FA_12588 \FA_INST_0[0].FA_INST_1[12].FA_  ( .A(A[12]), .B(n1037), .CI(C[12]), 
        .S(S[12]), .CO(C[13]) );
  FA_12587 \FA_INST_0[0].FA_INST_1[13].FA_  ( .A(A[13]), .B(n1038), .CI(C[13]), 
        .S(S[13]), .CO(C[14]) );
  FA_12586 \FA_INST_0[0].FA_INST_1[14].FA_  ( .A(A[14]), .B(n1039), .CI(C[14]), 
        .S(S[14]), .CO(C[15]) );
  FA_12585 \FA_INST_0[0].FA_INST_1[15].FA_  ( .A(A[15]), .B(n1040), .CI(C[15]), 
        .S(S[15]), .CO(C[16]) );
  FA_12584 \FA_INST_0[0].FA_INST_1[16].FA_  ( .A(A[16]), .B(n1041), .CI(C[16]), 
        .S(S[16]), .CO(C[17]) );
  FA_12583 \FA_INST_0[0].FA_INST_1[17].FA_  ( .A(A[17]), .B(n1042), .CI(C[17]), 
        .S(S[17]), .CO(C[18]) );
  FA_12582 \FA_INST_0[0].FA_INST_1[18].FA_  ( .A(A[18]), .B(n1043), .CI(C[18]), 
        .S(S[18]), .CO(C[19]) );
  FA_12581 \FA_INST_0[0].FA_INST_1[19].FA_  ( .A(A[19]), .B(n1044), .CI(C[19]), 
        .S(S[19]), .CO(C[20]) );
  FA_12580 \FA_INST_0[0].FA_INST_1[20].FA_  ( .A(A[20]), .B(n1045), .CI(C[20]), 
        .S(S[20]), .CO(C[21]) );
  FA_12579 \FA_INST_0[0].FA_INST_1[21].FA_  ( .A(A[21]), .B(n1046), .CI(C[21]), 
        .S(S[21]), .CO(C[22]) );
  FA_12578 \FA_INST_0[0].FA_INST_1[22].FA_  ( .A(A[22]), .B(n1047), .CI(C[22]), 
        .S(S[22]), .CO(C[23]) );
  FA_12577 \FA_INST_0[0].FA_INST_1[23].FA_  ( .A(A[23]), .B(n1048), .CI(C[23]), 
        .S(S[23]), .CO(C[24]) );
  FA_12576 \FA_INST_0[0].FA_INST_1[24].FA_  ( .A(A[24]), .B(n1049), .CI(C[24]), 
        .S(S[24]), .CO(C[25]) );
  FA_12575 \FA_INST_0[0].FA_INST_1[25].FA_  ( .A(A[25]), .B(n1050), .CI(C[25]), 
        .S(S[25]), .CO(C[26]) );
  FA_12574 \FA_INST_0[0].FA_INST_1[26].FA_  ( .A(A[26]), .B(n1051), .CI(C[26]), 
        .S(S[26]), .CO(C[27]) );
  FA_12573 \FA_INST_0[0].FA_INST_1[27].FA_  ( .A(A[27]), .B(n1052), .CI(C[27]), 
        .S(S[27]), .CO(C[28]) );
  FA_12572 \FA_INST_0[0].FA_INST_1[28].FA_  ( .A(A[28]), .B(n1053), .CI(C[28]), 
        .S(S[28]), .CO(C[29]) );
  FA_12571 \FA_INST_0[0].FA_INST_1[29].FA_  ( .A(A[29]), .B(n1054), .CI(C[29]), 
        .S(S[29]), .CO(C[30]) );
  FA_12570 \FA_INST_0[0].FA_INST_1[30].FA_  ( .A(A[30]), .B(n1055), .CI(C[30]), 
        .S(S[30]), .CO(C[31]) );
  FA_12569 \FA_INST_0[0].FA_INST_1[31].FA_  ( .A(A[31]), .B(n1056), .CI(C[31]), 
        .S(S[31]), .CO(C[32]) );
  FA_12568 \FA_INST_0[0].FA_INST_1[32].FA_  ( .A(A[32]), .B(n1057), .CI(C[32]), 
        .S(S[32]), .CO(C[33]) );
  FA_12567 \FA_INST_0[0].FA_INST_1[33].FA_  ( .A(A[33]), .B(n1058), .CI(C[33]), 
        .S(S[33]), .CO(C[34]) );
  FA_12566 \FA_INST_0[0].FA_INST_1[34].FA_  ( .A(A[34]), .B(n1059), .CI(C[34]), 
        .S(S[34]), .CO(C[35]) );
  FA_12565 \FA_INST_0[0].FA_INST_1[35].FA_  ( .A(A[35]), .B(n1060), .CI(C[35]), 
        .S(S[35]), .CO(C[36]) );
  FA_12564 \FA_INST_0[0].FA_INST_1[36].FA_  ( .A(A[36]), .B(n1061), .CI(C[36]), 
        .S(S[36]), .CO(C[37]) );
  FA_12563 \FA_INST_0[0].FA_INST_1[37].FA_  ( .A(A[37]), .B(n1062), .CI(C[37]), 
        .S(S[37]), .CO(C[38]) );
  FA_12562 \FA_INST_0[0].FA_INST_1[38].FA_  ( .A(A[38]), .B(n1063), .CI(C[38]), 
        .S(S[38]), .CO(C[39]) );
  FA_12561 \FA_INST_0[0].FA_INST_1[39].FA_  ( .A(A[39]), .B(n1064), .CI(C[39]), 
        .S(S[39]), .CO(C[40]) );
  FA_12560 \FA_INST_0[0].FA_INST_1[40].FA_  ( .A(A[40]), .B(n1065), .CI(C[40]), 
        .S(S[40]), .CO(C[41]) );
  FA_12559 \FA_INST_0[0].FA_INST_1[41].FA_  ( .A(A[41]), .B(n1066), .CI(C[41]), 
        .S(S[41]), .CO(C[42]) );
  FA_12558 \FA_INST_0[0].FA_INST_1[42].FA_  ( .A(A[42]), .B(n1067), .CI(C[42]), 
        .S(S[42]), .CO(C[43]) );
  FA_12557 \FA_INST_0[0].FA_INST_1[43].FA_  ( .A(A[43]), .B(n1068), .CI(C[43]), 
        .S(S[43]), .CO(C[44]) );
  FA_12556 \FA_INST_0[0].FA_INST_1[44].FA_  ( .A(A[44]), .B(n1069), .CI(C[44]), 
        .S(S[44]), .CO(C[45]) );
  FA_12555 \FA_INST_0[0].FA_INST_1[45].FA_  ( .A(A[45]), .B(n1070), .CI(C[45]), 
        .S(S[45]), .CO(C[46]) );
  FA_12554 \FA_INST_0[0].FA_INST_1[46].FA_  ( .A(A[46]), .B(n1071), .CI(C[46]), 
        .S(S[46]), .CO(C[47]) );
  FA_12553 \FA_INST_0[0].FA_INST_1[47].FA_  ( .A(A[47]), .B(n1072), .CI(C[47]), 
        .S(S[47]), .CO(C[48]) );
  FA_12552 \FA_INST_0[0].FA_INST_1[48].FA_  ( .A(A[48]), .B(n1073), .CI(C[48]), 
        .S(S[48]), .CO(C[49]) );
  FA_12551 \FA_INST_0[0].FA_INST_1[49].FA_  ( .A(A[49]), .B(n1074), .CI(C[49]), 
        .S(S[49]), .CO(C[50]) );
  FA_12550 \FA_INST_0[0].FA_INST_1[50].FA_  ( .A(A[50]), .B(n1075), .CI(C[50]), 
        .S(S[50]), .CO(C[51]) );
  FA_12549 \FA_INST_0[0].FA_INST_1[51].FA_  ( .A(A[51]), .B(n1076), .CI(C[51]), 
        .S(S[51]), .CO(C[52]) );
  FA_12548 \FA_INST_0[0].FA_INST_1[52].FA_  ( .A(A[52]), .B(n1077), .CI(C[52]), 
        .S(S[52]), .CO(C[53]) );
  FA_12547 \FA_INST_0[0].FA_INST_1[53].FA_  ( .A(A[53]), .B(n1078), .CI(C[53]), 
        .S(S[53]), .CO(C[54]) );
  FA_12546 \FA_INST_0[0].FA_INST_1[54].FA_  ( .A(A[54]), .B(n1079), .CI(C[54]), 
        .S(S[54]), .CO(C[55]) );
  FA_12545 \FA_INST_0[0].FA_INST_1[55].FA_  ( .A(A[55]), .B(n1080), .CI(C[55]), 
        .S(S[55]), .CO(C[56]) );
  FA_12544 \FA_INST_0[0].FA_INST_1[56].FA_  ( .A(A[56]), .B(n1081), .CI(C[56]), 
        .S(S[56]), .CO(C[57]) );
  FA_12543 \FA_INST_0[0].FA_INST_1[57].FA_  ( .A(A[57]), .B(n1082), .CI(C[57]), 
        .S(S[57]), .CO(C[58]) );
  FA_12542 \FA_INST_0[0].FA_INST_1[58].FA_  ( .A(A[58]), .B(n1083), .CI(C[58]), 
        .S(S[58]), .CO(C[59]) );
  FA_12541 \FA_INST_0[0].FA_INST_1[59].FA_  ( .A(A[59]), .B(n1084), .CI(C[59]), 
        .S(S[59]), .CO(C[60]) );
  FA_12540 \FA_INST_0[0].FA_INST_1[60].FA_  ( .A(A[60]), .B(n1085), .CI(C[60]), 
        .S(S[60]), .CO(C[61]) );
  FA_12539 \FA_INST_0[0].FA_INST_1[61].FA_  ( .A(A[61]), .B(n1086), .CI(C[61]), 
        .S(S[61]), .CO(C[62]) );
  FA_12538 \FA_INST_0[0].FA_INST_1[62].FA_  ( .A(A[62]), .B(n1087), .CI(C[62]), 
        .S(S[62]), .CO(C[63]) );
  FA_12537 \FA_INST_0[0].FA_INST_1[63].FA_  ( .A(A[63]), .B(n1088), .CI(C[63]), 
        .S(S[63]), .CO(C[64]) );
  FA_12536 \FA_INST_0[0].FA_INST_1[64].FA_  ( .A(A[64]), .B(n1089), .CI(C[64]), 
        .S(S[64]), .CO(C[65]) );
  FA_12535 \FA_INST_0[0].FA_INST_1[65].FA_  ( .A(A[65]), .B(n1090), .CI(C[65]), 
        .S(S[65]), .CO(C[66]) );
  FA_12534 \FA_INST_0[0].FA_INST_1[66].FA_  ( .A(A[66]), .B(n1091), .CI(C[66]), 
        .S(S[66]), .CO(C[67]) );
  FA_12533 \FA_INST_0[0].FA_INST_1[67].FA_  ( .A(A[67]), .B(n1092), .CI(C[67]), 
        .S(S[67]), .CO(C[68]) );
  FA_12532 \FA_INST_0[0].FA_INST_1[68].FA_  ( .A(A[68]), .B(n1093), .CI(C[68]), 
        .S(S[68]), .CO(C[69]) );
  FA_12531 \FA_INST_0[0].FA_INST_1[69].FA_  ( .A(A[69]), .B(n1094), .CI(C[69]), 
        .S(S[69]), .CO(C[70]) );
  FA_12530 \FA_INST_0[0].FA_INST_1[70].FA_  ( .A(A[70]), .B(n1095), .CI(C[70]), 
        .S(S[70]), .CO(C[71]) );
  FA_12529 \FA_INST_0[0].FA_INST_1[71].FA_  ( .A(A[71]), .B(n1096), .CI(C[71]), 
        .S(S[71]), .CO(C[72]) );
  FA_12528 \FA_INST_0[0].FA_INST_1[72].FA_  ( .A(A[72]), .B(n1097), .CI(C[72]), 
        .S(S[72]), .CO(C[73]) );
  FA_12527 \FA_INST_0[0].FA_INST_1[73].FA_  ( .A(A[73]), .B(n1098), .CI(C[73]), 
        .S(S[73]), .CO(C[74]) );
  FA_12526 \FA_INST_0[0].FA_INST_1[74].FA_  ( .A(A[74]), .B(n1099), .CI(C[74]), 
        .S(S[74]), .CO(C[75]) );
  FA_12525 \FA_INST_0[0].FA_INST_1[75].FA_  ( .A(A[75]), .B(n1100), .CI(C[75]), 
        .S(S[75]), .CO(C[76]) );
  FA_12524 \FA_INST_0[0].FA_INST_1[76].FA_  ( .A(A[76]), .B(n1101), .CI(C[76]), 
        .S(S[76]), .CO(C[77]) );
  FA_12523 \FA_INST_0[0].FA_INST_1[77].FA_  ( .A(A[77]), .B(n1102), .CI(C[77]), 
        .S(S[77]), .CO(C[78]) );
  FA_12522 \FA_INST_0[0].FA_INST_1[78].FA_  ( .A(A[78]), .B(n1103), .CI(C[78]), 
        .S(S[78]), .CO(C[79]) );
  FA_12521 \FA_INST_0[0].FA_INST_1[79].FA_  ( .A(A[79]), .B(n1104), .CI(C[79]), 
        .S(S[79]), .CO(C[80]) );
  FA_12520 \FA_INST_0[0].FA_INST_1[80].FA_  ( .A(A[80]), .B(n1105), .CI(C[80]), 
        .S(S[80]), .CO(C[81]) );
  FA_12519 \FA_INST_0[0].FA_INST_1[81].FA_  ( .A(A[81]), .B(n1106), .CI(C[81]), 
        .S(S[81]), .CO(C[82]) );
  FA_12518 \FA_INST_0[0].FA_INST_1[82].FA_  ( .A(A[82]), .B(n1107), .CI(C[82]), 
        .S(S[82]), .CO(C[83]) );
  FA_12517 \FA_INST_0[0].FA_INST_1[83].FA_  ( .A(A[83]), .B(n1108), .CI(C[83]), 
        .S(S[83]), .CO(C[84]) );
  FA_12516 \FA_INST_0[0].FA_INST_1[84].FA_  ( .A(A[84]), .B(n1109), .CI(C[84]), 
        .S(S[84]), .CO(C[85]) );
  FA_12515 \FA_INST_0[0].FA_INST_1[85].FA_  ( .A(A[85]), .B(n1110), .CI(C[85]), 
        .S(S[85]), .CO(C[86]) );
  FA_12514 \FA_INST_0[0].FA_INST_1[86].FA_  ( .A(A[86]), .B(n1111), .CI(C[86]), 
        .S(S[86]), .CO(C[87]) );
  FA_12513 \FA_INST_0[0].FA_INST_1[87].FA_  ( .A(A[87]), .B(n1112), .CI(C[87]), 
        .S(S[87]), .CO(C[88]) );
  FA_12512 \FA_INST_0[0].FA_INST_1[88].FA_  ( .A(A[88]), .B(n1113), .CI(C[88]), 
        .S(S[88]), .CO(C[89]) );
  FA_12511 \FA_INST_0[0].FA_INST_1[89].FA_  ( .A(A[89]), .B(n1114), .CI(C[89]), 
        .S(S[89]), .CO(C[90]) );
  FA_12510 \FA_INST_0[0].FA_INST_1[90].FA_  ( .A(A[90]), .B(n1115), .CI(C[90]), 
        .S(S[90]), .CO(C[91]) );
  FA_12509 \FA_INST_0[0].FA_INST_1[91].FA_  ( .A(A[91]), .B(n1116), .CI(C[91]), 
        .S(S[91]), .CO(C[92]) );
  FA_12508 \FA_INST_0[0].FA_INST_1[92].FA_  ( .A(A[92]), .B(n1117), .CI(C[92]), 
        .S(S[92]), .CO(C[93]) );
  FA_12507 \FA_INST_0[0].FA_INST_1[93].FA_  ( .A(A[93]), .B(n1118), .CI(C[93]), 
        .S(S[93]), .CO(C[94]) );
  FA_12506 \FA_INST_0[0].FA_INST_1[94].FA_  ( .A(A[94]), .B(n1119), .CI(C[94]), 
        .S(S[94]), .CO(C[95]) );
  FA_12505 \FA_INST_0[0].FA_INST_1[95].FA_  ( .A(A[95]), .B(n1120), .CI(C[95]), 
        .S(S[95]), .CO(C[96]) );
  FA_12504 \FA_INST_0[0].FA_INST_1[96].FA_  ( .A(A[96]), .B(n1121), .CI(C[96]), 
        .S(S[96]), .CO(C[97]) );
  FA_12503 \FA_INST_0[0].FA_INST_1[97].FA_  ( .A(A[97]), .B(n1122), .CI(C[97]), 
        .S(S[97]), .CO(C[98]) );
  FA_12502 \FA_INST_0[0].FA_INST_1[98].FA_  ( .A(A[98]), .B(n1123), .CI(C[98]), 
        .S(S[98]), .CO(C[99]) );
  FA_12501 \FA_INST_0[0].FA_INST_1[99].FA_  ( .A(A[99]), .B(n1124), .CI(C[99]), 
        .S(S[99]), .CO(C[100]) );
  FA_12500 \FA_INST_0[0].FA_INST_1[100].FA_  ( .A(A[100]), .B(n1125), .CI(
        C[100]), .S(S[100]), .CO(C[101]) );
  FA_12499 \FA_INST_0[0].FA_INST_1[101].FA_  ( .A(A[101]), .B(n1126), .CI(
        C[101]), .S(S[101]), .CO(C[102]) );
  FA_12498 \FA_INST_0[0].FA_INST_1[102].FA_  ( .A(A[102]), .B(n1127), .CI(
        C[102]), .S(S[102]), .CO(C[103]) );
  FA_12497 \FA_INST_0[0].FA_INST_1[103].FA_  ( .A(A[103]), .B(n1128), .CI(
        C[103]), .S(S[103]), .CO(C[104]) );
  FA_12496 \FA_INST_0[0].FA_INST_1[104].FA_  ( .A(A[104]), .B(n1129), .CI(
        C[104]), .S(S[104]), .CO(C[105]) );
  FA_12495 \FA_INST_0[0].FA_INST_1[105].FA_  ( .A(A[105]), .B(n1130), .CI(
        C[105]), .S(S[105]), .CO(C[106]) );
  FA_12494 \FA_INST_0[0].FA_INST_1[106].FA_  ( .A(A[106]), .B(n1131), .CI(
        C[106]), .S(S[106]), .CO(C[107]) );
  FA_12493 \FA_INST_0[0].FA_INST_1[107].FA_  ( .A(A[107]), .B(n1132), .CI(
        C[107]), .S(S[107]), .CO(C[108]) );
  FA_12492 \FA_INST_0[0].FA_INST_1[108].FA_  ( .A(A[108]), .B(n1133), .CI(
        C[108]), .S(S[108]), .CO(C[109]) );
  FA_12491 \FA_INST_0[0].FA_INST_1[109].FA_  ( .A(A[109]), .B(n1134), .CI(
        C[109]), .S(S[109]), .CO(C[110]) );
  FA_12490 \FA_INST_0[0].FA_INST_1[110].FA_  ( .A(A[110]), .B(n1135), .CI(
        C[110]), .S(S[110]), .CO(C[111]) );
  FA_12489 \FA_INST_0[0].FA_INST_1[111].FA_  ( .A(A[111]), .B(n1136), .CI(
        C[111]), .S(S[111]), .CO(C[112]) );
  FA_12488 \FA_INST_0[0].FA_INST_1[112].FA_  ( .A(A[112]), .B(n1137), .CI(
        C[112]), .S(S[112]), .CO(C[113]) );
  FA_12487 \FA_INST_0[0].FA_INST_1[113].FA_  ( .A(A[113]), .B(n1138), .CI(
        C[113]), .S(S[113]), .CO(C[114]) );
  FA_12486 \FA_INST_0[0].FA_INST_1[114].FA_  ( .A(A[114]), .B(n1139), .CI(
        C[114]), .S(S[114]), .CO(C[115]) );
  FA_12485 \FA_INST_0[0].FA_INST_1[115].FA_  ( .A(A[115]), .B(n1140), .CI(
        C[115]), .S(S[115]), .CO(C[116]) );
  FA_12484 \FA_INST_0[0].FA_INST_1[116].FA_  ( .A(A[116]), .B(n1141), .CI(
        C[116]), .S(S[116]), .CO(C[117]) );
  FA_12483 \FA_INST_0[0].FA_INST_1[117].FA_  ( .A(A[117]), .B(n1142), .CI(
        C[117]), .S(S[117]), .CO(C[118]) );
  FA_12482 \FA_INST_0[0].FA_INST_1[118].FA_  ( .A(A[118]), .B(n1143), .CI(
        C[118]), .S(S[118]), .CO(C[119]) );
  FA_12481 \FA_INST_0[0].FA_INST_1[119].FA_  ( .A(A[119]), .B(n1144), .CI(
        C[119]), .S(S[119]), .CO(C[120]) );
  FA_12480 \FA_INST_0[0].FA_INST_1[120].FA_  ( .A(A[120]), .B(n1145), .CI(
        C[120]), .S(S[120]), .CO(C[121]) );
  FA_12479 \FA_INST_0[0].FA_INST_1[121].FA_  ( .A(A[121]), .B(n1146), .CI(
        C[121]), .S(S[121]), .CO(C[122]) );
  FA_12478 \FA_INST_0[0].FA_INST_1[122].FA_  ( .A(A[122]), .B(n1147), .CI(
        C[122]), .S(S[122]), .CO(C[123]) );
  FA_12477 \FA_INST_0[0].FA_INST_1[123].FA_  ( .A(A[123]), .B(n1148), .CI(
        C[123]), .S(S[123]), .CO(C[124]) );
  FA_12476 \FA_INST_0[0].FA_INST_1[124].FA_  ( .A(A[124]), .B(n1149), .CI(
        C[124]), .S(S[124]), .CO(C[125]) );
  FA_12475 \FA_INST_0[0].FA_INST_1[125].FA_  ( .A(A[125]), .B(n1150), .CI(
        C[125]), .S(S[125]), .CO(C[126]) );
  FA_12474 \FA_INST_0[0].FA_INST_1[126].FA_  ( .A(A[126]), .B(n1151), .CI(
        C[126]), .S(S[126]), .CO(C[127]) );
  FA_12473 \FA_INST_0[0].FA_INST_1[127].FA_  ( .A(A[127]), .B(n1152), .CI(
        C[127]), .S(S[127]), .CO(C[128]) );
  FA_12472 \FA_INST_0[0].FA_INST_1[128].FA_  ( .A(A[128]), .B(n1153), .CI(
        C[128]), .S(S[128]), .CO(C[129]) );
  FA_12471 \FA_INST_0[0].FA_INST_1[129].FA_  ( .A(A[129]), .B(n1154), .CI(
        C[129]), .S(S[129]), .CO(C[130]) );
  FA_12470 \FA_INST_0[0].FA_INST_1[130].FA_  ( .A(A[130]), .B(n1155), .CI(
        C[130]), .S(S[130]), .CO(C[131]) );
  FA_12469 \FA_INST_0[0].FA_INST_1[131].FA_  ( .A(A[131]), .B(n1156), .CI(
        C[131]), .S(S[131]), .CO(C[132]) );
  FA_12468 \FA_INST_0[0].FA_INST_1[132].FA_  ( .A(A[132]), .B(n1157), .CI(
        C[132]), .S(S[132]), .CO(C[133]) );
  FA_12467 \FA_INST_0[0].FA_INST_1[133].FA_  ( .A(A[133]), .B(n1158), .CI(
        C[133]), .S(S[133]), .CO(C[134]) );
  FA_12466 \FA_INST_0[0].FA_INST_1[134].FA_  ( .A(A[134]), .B(n1159), .CI(
        C[134]), .S(S[134]), .CO(C[135]) );
  FA_12465 \FA_INST_0[0].FA_INST_1[135].FA_  ( .A(A[135]), .B(n1160), .CI(
        C[135]), .S(S[135]), .CO(C[136]) );
  FA_12464 \FA_INST_0[0].FA_INST_1[136].FA_  ( .A(A[136]), .B(n1161), .CI(
        C[136]), .S(S[136]), .CO(C[137]) );
  FA_12463 \FA_INST_0[0].FA_INST_1[137].FA_  ( .A(A[137]), .B(n1162), .CI(
        C[137]), .S(S[137]), .CO(C[138]) );
  FA_12462 \FA_INST_0[0].FA_INST_1[138].FA_  ( .A(A[138]), .B(n1163), .CI(
        C[138]), .S(S[138]), .CO(C[139]) );
  FA_12461 \FA_INST_0[0].FA_INST_1[139].FA_  ( .A(A[139]), .B(n1164), .CI(
        C[139]), .S(S[139]), .CO(C[140]) );
  FA_12460 \FA_INST_0[0].FA_INST_1[140].FA_  ( .A(A[140]), .B(n1165), .CI(
        C[140]), .S(S[140]), .CO(C[141]) );
  FA_12459 \FA_INST_0[0].FA_INST_1[141].FA_  ( .A(A[141]), .B(n1166), .CI(
        C[141]), .S(S[141]), .CO(C[142]) );
  FA_12458 \FA_INST_0[0].FA_INST_1[142].FA_  ( .A(A[142]), .B(n1167), .CI(
        C[142]), .S(S[142]), .CO(C[143]) );
  FA_12457 \FA_INST_0[0].FA_INST_1[143].FA_  ( .A(A[143]), .B(n1168), .CI(
        C[143]), .S(S[143]), .CO(C[144]) );
  FA_12456 \FA_INST_0[0].FA_INST_1[144].FA_  ( .A(A[144]), .B(n1169), .CI(
        C[144]), .S(S[144]), .CO(C[145]) );
  FA_12455 \FA_INST_0[0].FA_INST_1[145].FA_  ( .A(A[145]), .B(n1170), .CI(
        C[145]), .S(S[145]), .CO(C[146]) );
  FA_12454 \FA_INST_0[0].FA_INST_1[146].FA_  ( .A(A[146]), .B(n1171), .CI(
        C[146]), .S(S[146]), .CO(C[147]) );
  FA_12453 \FA_INST_0[0].FA_INST_1[147].FA_  ( .A(A[147]), .B(n1172), .CI(
        C[147]), .S(S[147]), .CO(C[148]) );
  FA_12452 \FA_INST_0[0].FA_INST_1[148].FA_  ( .A(A[148]), .B(n1173), .CI(
        C[148]), .S(S[148]), .CO(C[149]) );
  FA_12451 \FA_INST_0[0].FA_INST_1[149].FA_  ( .A(A[149]), .B(n1174), .CI(
        C[149]), .S(S[149]), .CO(C[150]) );
  FA_12450 \FA_INST_0[0].FA_INST_1[150].FA_  ( .A(A[150]), .B(n1175), .CI(
        C[150]), .S(S[150]), .CO(C[151]) );
  FA_12449 \FA_INST_0[0].FA_INST_1[151].FA_  ( .A(A[151]), .B(n1176), .CI(
        C[151]), .S(S[151]), .CO(C[152]) );
  FA_12448 \FA_INST_0[0].FA_INST_1[152].FA_  ( .A(A[152]), .B(n1177), .CI(
        C[152]), .S(S[152]), .CO(C[153]) );
  FA_12447 \FA_INST_0[0].FA_INST_1[153].FA_  ( .A(A[153]), .B(n1178), .CI(
        C[153]), .S(S[153]), .CO(C[154]) );
  FA_12446 \FA_INST_0[0].FA_INST_1[154].FA_  ( .A(A[154]), .B(n1179), .CI(
        C[154]), .S(S[154]), .CO(C[155]) );
  FA_12445 \FA_INST_0[0].FA_INST_1[155].FA_  ( .A(A[155]), .B(n1180), .CI(
        C[155]), .S(S[155]), .CO(C[156]) );
  FA_12444 \FA_INST_0[0].FA_INST_1[156].FA_  ( .A(A[156]), .B(n1181), .CI(
        C[156]), .S(S[156]), .CO(C[157]) );
  FA_12443 \FA_INST_0[0].FA_INST_1[157].FA_  ( .A(A[157]), .B(n1182), .CI(
        C[157]), .S(S[157]), .CO(C[158]) );
  FA_12442 \FA_INST_0[0].FA_INST_1[158].FA_  ( .A(A[158]), .B(n1183), .CI(
        C[158]), .S(S[158]), .CO(C[159]) );
  FA_12441 \FA_INST_0[0].FA_INST_1[159].FA_  ( .A(A[159]), .B(n1184), .CI(
        C[159]), .S(S[159]), .CO(C[160]) );
  FA_12440 \FA_INST_0[0].FA_INST_1[160].FA_  ( .A(A[160]), .B(n1185), .CI(
        C[160]), .S(S[160]), .CO(C[161]) );
  FA_12439 \FA_INST_0[0].FA_INST_1[161].FA_  ( .A(A[161]), .B(n1186), .CI(
        C[161]), .S(S[161]), .CO(C[162]) );
  FA_12438 \FA_INST_0[0].FA_INST_1[162].FA_  ( .A(A[162]), .B(n1187), .CI(
        C[162]), .S(S[162]), .CO(C[163]) );
  FA_12437 \FA_INST_0[0].FA_INST_1[163].FA_  ( .A(A[163]), .B(n1188), .CI(
        C[163]), .S(S[163]), .CO(C[164]) );
  FA_12436 \FA_INST_0[0].FA_INST_1[164].FA_  ( .A(A[164]), .B(n1189), .CI(
        C[164]), .S(S[164]), .CO(C[165]) );
  FA_12435 \FA_INST_0[0].FA_INST_1[165].FA_  ( .A(A[165]), .B(n1190), .CI(
        C[165]), .S(S[165]), .CO(C[166]) );
  FA_12434 \FA_INST_0[0].FA_INST_1[166].FA_  ( .A(A[166]), .B(n1191), .CI(
        C[166]), .S(S[166]), .CO(C[167]) );
  FA_12433 \FA_INST_0[0].FA_INST_1[167].FA_  ( .A(A[167]), .B(n1192), .CI(
        C[167]), .S(S[167]), .CO(C[168]) );
  FA_12432 \FA_INST_0[0].FA_INST_1[168].FA_  ( .A(A[168]), .B(n1193), .CI(
        C[168]), .S(S[168]), .CO(C[169]) );
  FA_12431 \FA_INST_0[0].FA_INST_1[169].FA_  ( .A(A[169]), .B(n1194), .CI(
        C[169]), .S(S[169]), .CO(C[170]) );
  FA_12430 \FA_INST_0[0].FA_INST_1[170].FA_  ( .A(A[170]), .B(n1195), .CI(
        C[170]), .S(S[170]), .CO(C[171]) );
  FA_12429 \FA_INST_0[0].FA_INST_1[171].FA_  ( .A(A[171]), .B(n1196), .CI(
        C[171]), .S(S[171]), .CO(C[172]) );
  FA_12428 \FA_INST_0[0].FA_INST_1[172].FA_  ( .A(A[172]), .B(n1197), .CI(
        C[172]), .S(S[172]), .CO(C[173]) );
  FA_12427 \FA_INST_0[0].FA_INST_1[173].FA_  ( .A(A[173]), .B(n1198), .CI(
        C[173]), .S(S[173]), .CO(C[174]) );
  FA_12426 \FA_INST_0[0].FA_INST_1[174].FA_  ( .A(A[174]), .B(n1199), .CI(
        C[174]), .S(S[174]), .CO(C[175]) );
  FA_12425 \FA_INST_0[0].FA_INST_1[175].FA_  ( .A(A[175]), .B(n1200), .CI(
        C[175]), .S(S[175]), .CO(C[176]) );
  FA_12424 \FA_INST_0[0].FA_INST_1[176].FA_  ( .A(A[176]), .B(n1201), .CI(
        C[176]), .S(S[176]), .CO(C[177]) );
  FA_12423 \FA_INST_0[0].FA_INST_1[177].FA_  ( .A(A[177]), .B(n1202), .CI(
        C[177]), .S(S[177]), .CO(C[178]) );
  FA_12422 \FA_INST_0[0].FA_INST_1[178].FA_  ( .A(A[178]), .B(n1203), .CI(
        C[178]), .S(S[178]), .CO(C[179]) );
  FA_12421 \FA_INST_0[0].FA_INST_1[179].FA_  ( .A(A[179]), .B(n1204), .CI(
        C[179]), .S(S[179]), .CO(C[180]) );
  FA_12420 \FA_INST_0[0].FA_INST_1[180].FA_  ( .A(A[180]), .B(n1205), .CI(
        C[180]), .S(S[180]), .CO(C[181]) );
  FA_12419 \FA_INST_0[0].FA_INST_1[181].FA_  ( .A(A[181]), .B(n1206), .CI(
        C[181]), .S(S[181]), .CO(C[182]) );
  FA_12418 \FA_INST_0[0].FA_INST_1[182].FA_  ( .A(A[182]), .B(n1207), .CI(
        C[182]), .S(S[182]), .CO(C[183]) );
  FA_12417 \FA_INST_0[0].FA_INST_1[183].FA_  ( .A(A[183]), .B(n1208), .CI(
        C[183]), .S(S[183]), .CO(C[184]) );
  FA_12416 \FA_INST_0[0].FA_INST_1[184].FA_  ( .A(A[184]), .B(n1209), .CI(
        C[184]), .S(S[184]), .CO(C[185]) );
  FA_12415 \FA_INST_0[0].FA_INST_1[185].FA_  ( .A(A[185]), .B(n1210), .CI(
        C[185]), .S(S[185]), .CO(C[186]) );
  FA_12414 \FA_INST_0[0].FA_INST_1[186].FA_  ( .A(A[186]), .B(n1211), .CI(
        C[186]), .S(S[186]), .CO(C[187]) );
  FA_12413 \FA_INST_0[0].FA_INST_1[187].FA_  ( .A(A[187]), .B(n1212), .CI(
        C[187]), .S(S[187]), .CO(C[188]) );
  FA_12412 \FA_INST_0[0].FA_INST_1[188].FA_  ( .A(A[188]), .B(n1213), .CI(
        C[188]), .S(S[188]), .CO(C[189]) );
  FA_12411 \FA_INST_0[0].FA_INST_1[189].FA_  ( .A(A[189]), .B(n1214), .CI(
        C[189]), .S(S[189]), .CO(C[190]) );
  FA_12410 \FA_INST_0[0].FA_INST_1[190].FA_  ( .A(A[190]), .B(n1215), .CI(
        C[190]), .S(S[190]), .CO(C[191]) );
  FA_12409 \FA_INST_0[0].FA_INST_1[191].FA_  ( .A(A[191]), .B(n1216), .CI(
        C[191]), .S(S[191]), .CO(C[192]) );
  FA_12408 \FA_INST_0[0].FA_INST_1[192].FA_  ( .A(A[192]), .B(n1217), .CI(
        C[192]), .S(S[192]), .CO(C[193]) );
  FA_12407 \FA_INST_0[0].FA_INST_1[193].FA_  ( .A(A[193]), .B(n1218), .CI(
        C[193]), .S(S[193]), .CO(C[194]) );
  FA_12406 \FA_INST_0[0].FA_INST_1[194].FA_  ( .A(A[194]), .B(n1219), .CI(
        C[194]), .S(S[194]), .CO(C[195]) );
  FA_12405 \FA_INST_0[0].FA_INST_1[195].FA_  ( .A(A[195]), .B(n1220), .CI(
        C[195]), .S(S[195]), .CO(C[196]) );
  FA_12404 \FA_INST_0[0].FA_INST_1[196].FA_  ( .A(A[196]), .B(n1221), .CI(
        C[196]), .S(S[196]), .CO(C[197]) );
  FA_12403 \FA_INST_0[0].FA_INST_1[197].FA_  ( .A(A[197]), .B(n1222), .CI(
        C[197]), .S(S[197]), .CO(C[198]) );
  FA_12402 \FA_INST_0[0].FA_INST_1[198].FA_  ( .A(A[198]), .B(n1223), .CI(
        C[198]), .S(S[198]), .CO(C[199]) );
  FA_12401 \FA_INST_0[0].FA_INST_1[199].FA_  ( .A(A[199]), .B(n1224), .CI(
        C[199]), .S(S[199]), .CO(C[200]) );
  FA_12400 \FA_INST_0[0].FA_INST_1[200].FA_  ( .A(A[200]), .B(n1225), .CI(
        C[200]), .S(S[200]), .CO(C[201]) );
  FA_12399 \FA_INST_0[0].FA_INST_1[201].FA_  ( .A(A[201]), .B(n1226), .CI(
        C[201]), .S(S[201]), .CO(C[202]) );
  FA_12398 \FA_INST_0[0].FA_INST_1[202].FA_  ( .A(A[202]), .B(n1227), .CI(
        C[202]), .S(S[202]), .CO(C[203]) );
  FA_12397 \FA_INST_0[0].FA_INST_1[203].FA_  ( .A(A[203]), .B(n1228), .CI(
        C[203]), .S(S[203]), .CO(C[204]) );
  FA_12396 \FA_INST_0[0].FA_INST_1[204].FA_  ( .A(A[204]), .B(n1229), .CI(
        C[204]), .S(S[204]), .CO(C[205]) );
  FA_12395 \FA_INST_0[0].FA_INST_1[205].FA_  ( .A(A[205]), .B(n1230), .CI(
        C[205]), .S(S[205]), .CO(C[206]) );
  FA_12394 \FA_INST_0[0].FA_INST_1[206].FA_  ( .A(A[206]), .B(n1231), .CI(
        C[206]), .S(S[206]), .CO(C[207]) );
  FA_12393 \FA_INST_0[0].FA_INST_1[207].FA_  ( .A(A[207]), .B(n1232), .CI(
        C[207]), .S(S[207]), .CO(C[208]) );
  FA_12392 \FA_INST_0[0].FA_INST_1[208].FA_  ( .A(A[208]), .B(n1233), .CI(
        C[208]), .S(S[208]), .CO(C[209]) );
  FA_12391 \FA_INST_0[0].FA_INST_1[209].FA_  ( .A(A[209]), .B(n1234), .CI(
        C[209]), .S(S[209]), .CO(C[210]) );
  FA_12390 \FA_INST_0[0].FA_INST_1[210].FA_  ( .A(A[210]), .B(n1235), .CI(
        C[210]), .S(S[210]), .CO(C[211]) );
  FA_12389 \FA_INST_0[0].FA_INST_1[211].FA_  ( .A(A[211]), .B(n1236), .CI(
        C[211]), .S(S[211]), .CO(C[212]) );
  FA_12388 \FA_INST_0[0].FA_INST_1[212].FA_  ( .A(A[212]), .B(n1237), .CI(
        C[212]), .S(S[212]), .CO(C[213]) );
  FA_12387 \FA_INST_0[0].FA_INST_1[213].FA_  ( .A(A[213]), .B(n1238), .CI(
        C[213]), .S(S[213]), .CO(C[214]) );
  FA_12386 \FA_INST_0[0].FA_INST_1[214].FA_  ( .A(A[214]), .B(n1239), .CI(
        C[214]), .S(S[214]), .CO(C[215]) );
  FA_12385 \FA_INST_0[0].FA_INST_1[215].FA_  ( .A(A[215]), .B(n1240), .CI(
        C[215]), .S(S[215]), .CO(C[216]) );
  FA_12384 \FA_INST_0[0].FA_INST_1[216].FA_  ( .A(A[216]), .B(n1241), .CI(
        C[216]), .S(S[216]), .CO(C[217]) );
  FA_12383 \FA_INST_0[0].FA_INST_1[217].FA_  ( .A(A[217]), .B(n1242), .CI(
        C[217]), .S(S[217]), .CO(C[218]) );
  FA_12382 \FA_INST_0[0].FA_INST_1[218].FA_  ( .A(A[218]), .B(n1243), .CI(
        C[218]), .S(S[218]), .CO(C[219]) );
  FA_12381 \FA_INST_0[0].FA_INST_1[219].FA_  ( .A(A[219]), .B(n1244), .CI(
        C[219]), .S(S[219]), .CO(C[220]) );
  FA_12380 \FA_INST_0[0].FA_INST_1[220].FA_  ( .A(A[220]), .B(n1245), .CI(
        C[220]), .S(S[220]), .CO(C[221]) );
  FA_12379 \FA_INST_0[0].FA_INST_1[221].FA_  ( .A(A[221]), .B(n1246), .CI(
        C[221]), .S(S[221]), .CO(C[222]) );
  FA_12378 \FA_INST_0[0].FA_INST_1[222].FA_  ( .A(A[222]), .B(n1247), .CI(
        C[222]), .S(S[222]), .CO(C[223]) );
  FA_12377 \FA_INST_0[0].FA_INST_1[223].FA_  ( .A(A[223]), .B(n1248), .CI(
        C[223]), .S(S[223]), .CO(C[224]) );
  FA_12376 \FA_INST_0[0].FA_INST_1[224].FA_  ( .A(A[224]), .B(n1249), .CI(
        C[224]), .S(S[224]), .CO(C[225]) );
  FA_12375 \FA_INST_0[0].FA_INST_1[225].FA_  ( .A(A[225]), .B(n1250), .CI(
        C[225]), .S(S[225]), .CO(C[226]) );
  FA_12374 \FA_INST_0[0].FA_INST_1[226].FA_  ( .A(A[226]), .B(n1251), .CI(
        C[226]), .S(S[226]), .CO(C[227]) );
  FA_12373 \FA_INST_0[0].FA_INST_1[227].FA_  ( .A(A[227]), .B(n1252), .CI(
        C[227]), .S(S[227]), .CO(C[228]) );
  FA_12372 \FA_INST_0[0].FA_INST_1[228].FA_  ( .A(A[228]), .B(n1253), .CI(
        C[228]), .S(S[228]), .CO(C[229]) );
  FA_12371 \FA_INST_0[0].FA_INST_1[229].FA_  ( .A(A[229]), .B(n1254), .CI(
        C[229]), .S(S[229]), .CO(C[230]) );
  FA_12370 \FA_INST_0[0].FA_INST_1[230].FA_  ( .A(A[230]), .B(n1255), .CI(
        C[230]), .S(S[230]), .CO(C[231]) );
  FA_12369 \FA_INST_0[0].FA_INST_1[231].FA_  ( .A(A[231]), .B(n1256), .CI(
        C[231]), .S(S[231]), .CO(C[232]) );
  FA_12368 \FA_INST_0[0].FA_INST_1[232].FA_  ( .A(A[232]), .B(n1257), .CI(
        C[232]), .S(S[232]), .CO(C[233]) );
  FA_12367 \FA_INST_0[0].FA_INST_1[233].FA_  ( .A(A[233]), .B(n1258), .CI(
        C[233]), .S(S[233]), .CO(C[234]) );
  FA_12366 \FA_INST_0[0].FA_INST_1[234].FA_  ( .A(A[234]), .B(n1259), .CI(
        C[234]), .S(S[234]), .CO(C[235]) );
  FA_12365 \FA_INST_0[0].FA_INST_1[235].FA_  ( .A(A[235]), .B(n1260), .CI(
        C[235]), .S(S[235]), .CO(C[236]) );
  FA_12364 \FA_INST_0[0].FA_INST_1[236].FA_  ( .A(A[236]), .B(n1261), .CI(
        C[236]), .S(S[236]), .CO(C[237]) );
  FA_12363 \FA_INST_0[0].FA_INST_1[237].FA_  ( .A(A[237]), .B(n1262), .CI(
        C[237]), .S(S[237]), .CO(C[238]) );
  FA_12362 \FA_INST_0[0].FA_INST_1[238].FA_  ( .A(A[238]), .B(n1263), .CI(
        C[238]), .S(S[238]), .CO(C[239]) );
  FA_12361 \FA_INST_0[0].FA_INST_1[239].FA_  ( .A(A[239]), .B(n1264), .CI(
        C[239]), .S(S[239]), .CO(C[240]) );
  FA_12360 \FA_INST_0[0].FA_INST_1[240].FA_  ( .A(A[240]), .B(n1265), .CI(
        C[240]), .S(S[240]), .CO(C[241]) );
  FA_12359 \FA_INST_0[0].FA_INST_1[241].FA_  ( .A(A[241]), .B(n1266), .CI(
        C[241]), .S(S[241]), .CO(C[242]) );
  FA_12358 \FA_INST_0[0].FA_INST_1[242].FA_  ( .A(A[242]), .B(n1267), .CI(
        C[242]), .S(S[242]), .CO(C[243]) );
  FA_12357 \FA_INST_0[0].FA_INST_1[243].FA_  ( .A(A[243]), .B(n1268), .CI(
        C[243]), .S(S[243]), .CO(C[244]) );
  FA_12356 \FA_INST_0[0].FA_INST_1[244].FA_  ( .A(A[244]), .B(n1269), .CI(
        C[244]), .S(S[244]), .CO(C[245]) );
  FA_12355 \FA_INST_0[0].FA_INST_1[245].FA_  ( .A(A[245]), .B(n1270), .CI(
        C[245]), .S(S[245]), .CO(C[246]) );
  FA_12354 \FA_INST_0[0].FA_INST_1[246].FA_  ( .A(A[246]), .B(n1271), .CI(
        C[246]), .S(S[246]), .CO(C[247]) );
  FA_12353 \FA_INST_0[0].FA_INST_1[247].FA_  ( .A(A[247]), .B(n1272), .CI(
        C[247]), .S(S[247]), .CO(C[248]) );
  FA_12352 \FA_INST_0[0].FA_INST_1[248].FA_  ( .A(A[248]), .B(n1273), .CI(
        C[248]), .S(S[248]), .CO(C[249]) );
  FA_12351 \FA_INST_0[0].FA_INST_1[249].FA_  ( .A(A[249]), .B(n1274), .CI(
        C[249]), .S(S[249]), .CO(C[250]) );
  FA_12350 \FA_INST_0[0].FA_INST_1[250].FA_  ( .A(A[250]), .B(n1275), .CI(
        C[250]), .S(S[250]), .CO(C[251]) );
  FA_12349 \FA_INST_0[0].FA_INST_1[251].FA_  ( .A(A[251]), .B(n1276), .CI(
        C[251]), .S(S[251]), .CO(C[252]) );
  FA_12348 \FA_INST_0[0].FA_INST_1[252].FA_  ( .A(A[252]), .B(n1277), .CI(
        C[252]), .S(S[252]), .CO(C[253]) );
  FA_12347 \FA_INST_0[0].FA_INST_1[253].FA_  ( .A(A[253]), .B(n1278), .CI(
        C[253]), .S(S[253]), .CO(C[254]) );
  FA_12346 \FA_INST_0[0].FA_INST_1[254].FA_  ( .A(A[254]), .B(n1279), .CI(
        C[254]), .S(S[254]), .CO(C[255]) );
  FA_12345 \FA_INST_0[0].FA_INST_1[255].FA_  ( .A(A[255]), .B(n1280), .CI(
        C[255]), .S(S[255]), .CO(C[256]) );
  FA_12344 \FA_INST_0[0].FA_INST_1[256].FA_  ( .A(A[256]), .B(n1281), .CI(
        C[256]), .S(S[256]), .CO(C[257]) );
  FA_12343 \FA_INST_0[0].FA_INST_1[257].FA_  ( .A(A[257]), .B(n1282), .CI(
        C[257]), .S(S[257]), .CO(C[258]) );
  FA_12342 \FA_INST_0[0].FA_INST_1[258].FA_  ( .A(A[258]), .B(n1283), .CI(
        C[258]), .S(S[258]), .CO(C[259]) );
  FA_12341 \FA_INST_0[0].FA_INST_1[259].FA_  ( .A(A[259]), .B(n1284), .CI(
        C[259]), .S(S[259]), .CO(C[260]) );
  FA_12340 \FA_INST_0[0].FA_INST_1[260].FA_  ( .A(A[260]), .B(n1285), .CI(
        C[260]), .S(S[260]), .CO(C[261]) );
  FA_12339 \FA_INST_0[0].FA_INST_1[261].FA_  ( .A(A[261]), .B(n1286), .CI(
        C[261]), .S(S[261]), .CO(C[262]) );
  FA_12338 \FA_INST_0[0].FA_INST_1[262].FA_  ( .A(A[262]), .B(n1287), .CI(
        C[262]), .S(S[262]), .CO(C[263]) );
  FA_12337 \FA_INST_0[0].FA_INST_1[263].FA_  ( .A(A[263]), .B(n1288), .CI(
        C[263]), .S(S[263]), .CO(C[264]) );
  FA_12336 \FA_INST_0[0].FA_INST_1[264].FA_  ( .A(A[264]), .B(n1289), .CI(
        C[264]), .S(S[264]), .CO(C[265]) );
  FA_12335 \FA_INST_0[0].FA_INST_1[265].FA_  ( .A(A[265]), .B(n1290), .CI(
        C[265]), .S(S[265]), .CO(C[266]) );
  FA_12334 \FA_INST_0[0].FA_INST_1[266].FA_  ( .A(A[266]), .B(n1291), .CI(
        C[266]), .S(S[266]), .CO(C[267]) );
  FA_12333 \FA_INST_0[0].FA_INST_1[267].FA_  ( .A(A[267]), .B(n1292), .CI(
        C[267]), .S(S[267]), .CO(C[268]) );
  FA_12332 \FA_INST_0[0].FA_INST_1[268].FA_  ( .A(A[268]), .B(n1293), .CI(
        C[268]), .S(S[268]), .CO(C[269]) );
  FA_12331 \FA_INST_0[0].FA_INST_1[269].FA_  ( .A(A[269]), .B(n1294), .CI(
        C[269]), .S(S[269]), .CO(C[270]) );
  FA_12330 \FA_INST_0[0].FA_INST_1[270].FA_  ( .A(A[270]), .B(n1295), .CI(
        C[270]), .S(S[270]), .CO(C[271]) );
  FA_12329 \FA_INST_0[0].FA_INST_1[271].FA_  ( .A(A[271]), .B(n1296), .CI(
        C[271]), .S(S[271]), .CO(C[272]) );
  FA_12328 \FA_INST_0[0].FA_INST_1[272].FA_  ( .A(A[272]), .B(n1297), .CI(
        C[272]), .S(S[272]), .CO(C[273]) );
  FA_12327 \FA_INST_0[0].FA_INST_1[273].FA_  ( .A(A[273]), .B(n1298), .CI(
        C[273]), .S(S[273]), .CO(C[274]) );
  FA_12326 \FA_INST_0[0].FA_INST_1[274].FA_  ( .A(A[274]), .B(n1299), .CI(
        C[274]), .S(S[274]), .CO(C[275]) );
  FA_12325 \FA_INST_0[0].FA_INST_1[275].FA_  ( .A(A[275]), .B(n1300), .CI(
        C[275]), .S(S[275]), .CO(C[276]) );
  FA_12324 \FA_INST_0[0].FA_INST_1[276].FA_  ( .A(A[276]), .B(n1301), .CI(
        C[276]), .S(S[276]), .CO(C[277]) );
  FA_12323 \FA_INST_0[0].FA_INST_1[277].FA_  ( .A(A[277]), .B(n1302), .CI(
        C[277]), .S(S[277]), .CO(C[278]) );
  FA_12322 \FA_INST_0[0].FA_INST_1[278].FA_  ( .A(A[278]), .B(n1303), .CI(
        C[278]), .S(S[278]), .CO(C[279]) );
  FA_12321 \FA_INST_0[0].FA_INST_1[279].FA_  ( .A(A[279]), .B(n1304), .CI(
        C[279]), .S(S[279]), .CO(C[280]) );
  FA_12320 \FA_INST_0[0].FA_INST_1[280].FA_  ( .A(A[280]), .B(n1305), .CI(
        C[280]), .S(S[280]), .CO(C[281]) );
  FA_12319 \FA_INST_0[0].FA_INST_1[281].FA_  ( .A(A[281]), .B(n1306), .CI(
        C[281]), .S(S[281]), .CO(C[282]) );
  FA_12318 \FA_INST_0[0].FA_INST_1[282].FA_  ( .A(A[282]), .B(n1307), .CI(
        C[282]), .S(S[282]), .CO(C[283]) );
  FA_12317 \FA_INST_0[0].FA_INST_1[283].FA_  ( .A(A[283]), .B(n1308), .CI(
        C[283]), .S(S[283]), .CO(C[284]) );
  FA_12316 \FA_INST_0[0].FA_INST_1[284].FA_  ( .A(A[284]), .B(n1309), .CI(
        C[284]), .S(S[284]), .CO(C[285]) );
  FA_12315 \FA_INST_0[0].FA_INST_1[285].FA_  ( .A(A[285]), .B(n1310), .CI(
        C[285]), .S(S[285]), .CO(C[286]) );
  FA_12314 \FA_INST_0[0].FA_INST_1[286].FA_  ( .A(A[286]), .B(n1311), .CI(
        C[286]), .S(S[286]), .CO(C[287]) );
  FA_12313 \FA_INST_0[0].FA_INST_1[287].FA_  ( .A(A[287]), .B(n1312), .CI(
        C[287]), .S(S[287]), .CO(C[288]) );
  FA_12312 \FA_INST_0[0].FA_INST_1[288].FA_  ( .A(A[288]), .B(n1313), .CI(
        C[288]), .S(S[288]), .CO(C[289]) );
  FA_12311 \FA_INST_0[0].FA_INST_1[289].FA_  ( .A(A[289]), .B(n1314), .CI(
        C[289]), .S(S[289]), .CO(C[290]) );
  FA_12310 \FA_INST_0[0].FA_INST_1[290].FA_  ( .A(A[290]), .B(n1315), .CI(
        C[290]), .S(S[290]), .CO(C[291]) );
  FA_12309 \FA_INST_0[0].FA_INST_1[291].FA_  ( .A(A[291]), .B(n1316), .CI(
        C[291]), .S(S[291]), .CO(C[292]) );
  FA_12308 \FA_INST_0[0].FA_INST_1[292].FA_  ( .A(A[292]), .B(n1317), .CI(
        C[292]), .S(S[292]), .CO(C[293]) );
  FA_12307 \FA_INST_0[0].FA_INST_1[293].FA_  ( .A(A[293]), .B(n1318), .CI(
        C[293]), .S(S[293]), .CO(C[294]) );
  FA_12306 \FA_INST_0[0].FA_INST_1[294].FA_  ( .A(A[294]), .B(n1319), .CI(
        C[294]), .S(S[294]), .CO(C[295]) );
  FA_12305 \FA_INST_0[0].FA_INST_1[295].FA_  ( .A(A[295]), .B(n1320), .CI(
        C[295]), .S(S[295]), .CO(C[296]) );
  FA_12304 \FA_INST_0[0].FA_INST_1[296].FA_  ( .A(A[296]), .B(n1321), .CI(
        C[296]), .S(S[296]), .CO(C[297]) );
  FA_12303 \FA_INST_0[0].FA_INST_1[297].FA_  ( .A(A[297]), .B(n1322), .CI(
        C[297]), .S(S[297]), .CO(C[298]) );
  FA_12302 \FA_INST_0[0].FA_INST_1[298].FA_  ( .A(A[298]), .B(n1323), .CI(
        C[298]), .S(S[298]), .CO(C[299]) );
  FA_12301 \FA_INST_0[0].FA_INST_1[299].FA_  ( .A(A[299]), .B(n1324), .CI(
        C[299]), .S(S[299]), .CO(C[300]) );
  FA_12300 \FA_INST_0[0].FA_INST_1[300].FA_  ( .A(A[300]), .B(n1325), .CI(
        C[300]), .S(S[300]), .CO(C[301]) );
  FA_12299 \FA_INST_0[0].FA_INST_1[301].FA_  ( .A(A[301]), .B(n1326), .CI(
        C[301]), .S(S[301]), .CO(C[302]) );
  FA_12298 \FA_INST_0[0].FA_INST_1[302].FA_  ( .A(A[302]), .B(n1327), .CI(
        C[302]), .S(S[302]), .CO(C[303]) );
  FA_12297 \FA_INST_0[0].FA_INST_1[303].FA_  ( .A(A[303]), .B(n1328), .CI(
        C[303]), .S(S[303]), .CO(C[304]) );
  FA_12296 \FA_INST_0[0].FA_INST_1[304].FA_  ( .A(A[304]), .B(n1329), .CI(
        C[304]), .S(S[304]), .CO(C[305]) );
  FA_12295 \FA_INST_0[0].FA_INST_1[305].FA_  ( .A(A[305]), .B(n1330), .CI(
        C[305]), .S(S[305]), .CO(C[306]) );
  FA_12294 \FA_INST_0[0].FA_INST_1[306].FA_  ( .A(A[306]), .B(n1331), .CI(
        C[306]), .S(S[306]), .CO(C[307]) );
  FA_12293 \FA_INST_0[0].FA_INST_1[307].FA_  ( .A(A[307]), .B(n1332), .CI(
        C[307]), .S(S[307]), .CO(C[308]) );
  FA_12292 \FA_INST_0[0].FA_INST_1[308].FA_  ( .A(A[308]), .B(n1333), .CI(
        C[308]), .S(S[308]), .CO(C[309]) );
  FA_12291 \FA_INST_0[0].FA_INST_1[309].FA_  ( .A(A[309]), .B(n1334), .CI(
        C[309]), .S(S[309]), .CO(C[310]) );
  FA_12290 \FA_INST_0[0].FA_INST_1[310].FA_  ( .A(A[310]), .B(n1335), .CI(
        C[310]), .S(S[310]), .CO(C[311]) );
  FA_12289 \FA_INST_0[0].FA_INST_1[311].FA_  ( .A(A[311]), .B(n1336), .CI(
        C[311]), .S(S[311]), .CO(C[312]) );
  FA_12288 \FA_INST_0[0].FA_INST_1[312].FA_  ( .A(A[312]), .B(n1337), .CI(
        C[312]), .S(S[312]), .CO(C[313]) );
  FA_12287 \FA_INST_0[0].FA_INST_1[313].FA_  ( .A(A[313]), .B(n1338), .CI(
        C[313]), .S(S[313]), .CO(C[314]) );
  FA_12286 \FA_INST_0[0].FA_INST_1[314].FA_  ( .A(A[314]), .B(n1339), .CI(
        C[314]), .S(S[314]), .CO(C[315]) );
  FA_12285 \FA_INST_0[0].FA_INST_1[315].FA_  ( .A(A[315]), .B(n1340), .CI(
        C[315]), .S(S[315]), .CO(C[316]) );
  FA_12284 \FA_INST_0[0].FA_INST_1[316].FA_  ( .A(A[316]), .B(n1341), .CI(
        C[316]), .S(S[316]), .CO(C[317]) );
  FA_12283 \FA_INST_0[0].FA_INST_1[317].FA_  ( .A(A[317]), .B(n1342), .CI(
        C[317]), .S(S[317]), .CO(C[318]) );
  FA_12282 \FA_INST_0[0].FA_INST_1[318].FA_  ( .A(A[318]), .B(n1343), .CI(
        C[318]), .S(S[318]), .CO(C[319]) );
  FA_12281 \FA_INST_0[0].FA_INST_1[319].FA_  ( .A(A[319]), .B(n1344), .CI(
        C[319]), .S(S[319]), .CO(C[320]) );
  FA_12280 \FA_INST_0[0].FA_INST_1[320].FA_  ( .A(A[320]), .B(n1345), .CI(
        C[320]), .S(S[320]), .CO(C[321]) );
  FA_12279 \FA_INST_0[0].FA_INST_1[321].FA_  ( .A(A[321]), .B(n1346), .CI(
        C[321]), .S(S[321]), .CO(C[322]) );
  FA_12278 \FA_INST_0[0].FA_INST_1[322].FA_  ( .A(A[322]), .B(n1347), .CI(
        C[322]), .S(S[322]), .CO(C[323]) );
  FA_12277 \FA_INST_0[0].FA_INST_1[323].FA_  ( .A(A[323]), .B(n1348), .CI(
        C[323]), .S(S[323]), .CO(C[324]) );
  FA_12276 \FA_INST_0[0].FA_INST_1[324].FA_  ( .A(A[324]), .B(n1349), .CI(
        C[324]), .S(S[324]), .CO(C[325]) );
  FA_12275 \FA_INST_0[0].FA_INST_1[325].FA_  ( .A(A[325]), .B(n1350), .CI(
        C[325]), .S(S[325]), .CO(C[326]) );
  FA_12274 \FA_INST_0[0].FA_INST_1[326].FA_  ( .A(A[326]), .B(n1351), .CI(
        C[326]), .S(S[326]), .CO(C[327]) );
  FA_12273 \FA_INST_0[0].FA_INST_1[327].FA_  ( .A(A[327]), .B(n1352), .CI(
        C[327]), .S(S[327]), .CO(C[328]) );
  FA_12272 \FA_INST_0[0].FA_INST_1[328].FA_  ( .A(A[328]), .B(n1353), .CI(
        C[328]), .S(S[328]), .CO(C[329]) );
  FA_12271 \FA_INST_0[0].FA_INST_1[329].FA_  ( .A(A[329]), .B(n1354), .CI(
        C[329]), .S(S[329]), .CO(C[330]) );
  FA_12270 \FA_INST_0[0].FA_INST_1[330].FA_  ( .A(A[330]), .B(n1355), .CI(
        C[330]), .S(S[330]), .CO(C[331]) );
  FA_12269 \FA_INST_0[0].FA_INST_1[331].FA_  ( .A(A[331]), .B(n1356), .CI(
        C[331]), .S(S[331]), .CO(C[332]) );
  FA_12268 \FA_INST_0[0].FA_INST_1[332].FA_  ( .A(A[332]), .B(n1357), .CI(
        C[332]), .S(S[332]), .CO(C[333]) );
  FA_12267 \FA_INST_0[0].FA_INST_1[333].FA_  ( .A(A[333]), .B(n1358), .CI(
        C[333]), .S(S[333]), .CO(C[334]) );
  FA_12266 \FA_INST_0[0].FA_INST_1[334].FA_  ( .A(A[334]), .B(n1359), .CI(
        C[334]), .S(S[334]), .CO(C[335]) );
  FA_12265 \FA_INST_0[0].FA_INST_1[335].FA_  ( .A(A[335]), .B(n1360), .CI(
        C[335]), .S(S[335]), .CO(C[336]) );
  FA_12264 \FA_INST_0[0].FA_INST_1[336].FA_  ( .A(A[336]), .B(n1361), .CI(
        C[336]), .S(S[336]), .CO(C[337]) );
  FA_12263 \FA_INST_0[0].FA_INST_1[337].FA_  ( .A(A[337]), .B(n1362), .CI(
        C[337]), .S(S[337]), .CO(C[338]) );
  FA_12262 \FA_INST_0[0].FA_INST_1[338].FA_  ( .A(A[338]), .B(n1363), .CI(
        C[338]), .S(S[338]), .CO(C[339]) );
  FA_12261 \FA_INST_0[0].FA_INST_1[339].FA_  ( .A(A[339]), .B(n1364), .CI(
        C[339]), .S(S[339]), .CO(C[340]) );
  FA_12260 \FA_INST_0[0].FA_INST_1[340].FA_  ( .A(A[340]), .B(n1365), .CI(
        C[340]), .S(S[340]), .CO(C[341]) );
  FA_12259 \FA_INST_0[0].FA_INST_1[341].FA_  ( .A(A[341]), .B(n1366), .CI(
        C[341]), .S(S[341]), .CO(C[342]) );
  FA_12258 \FA_INST_0[0].FA_INST_1[342].FA_  ( .A(A[342]), .B(n1367), .CI(
        C[342]), .S(S[342]), .CO(C[343]) );
  FA_12257 \FA_INST_0[0].FA_INST_1[343].FA_  ( .A(A[343]), .B(n1368), .CI(
        C[343]), .S(S[343]), .CO(C[344]) );
  FA_12256 \FA_INST_0[0].FA_INST_1[344].FA_  ( .A(A[344]), .B(n1369), .CI(
        C[344]), .S(S[344]), .CO(C[345]) );
  FA_12255 \FA_INST_0[0].FA_INST_1[345].FA_  ( .A(A[345]), .B(n1370), .CI(
        C[345]), .S(S[345]), .CO(C[346]) );
  FA_12254 \FA_INST_0[0].FA_INST_1[346].FA_  ( .A(A[346]), .B(n1371), .CI(
        C[346]), .S(S[346]), .CO(C[347]) );
  FA_12253 \FA_INST_0[0].FA_INST_1[347].FA_  ( .A(A[347]), .B(n1372), .CI(
        C[347]), .S(S[347]), .CO(C[348]) );
  FA_12252 \FA_INST_0[0].FA_INST_1[348].FA_  ( .A(A[348]), .B(n1373), .CI(
        C[348]), .S(S[348]), .CO(C[349]) );
  FA_12251 \FA_INST_0[0].FA_INST_1[349].FA_  ( .A(A[349]), .B(n1374), .CI(
        C[349]), .S(S[349]), .CO(C[350]) );
  FA_12250 \FA_INST_0[0].FA_INST_1[350].FA_  ( .A(A[350]), .B(n1375), .CI(
        C[350]), .S(S[350]), .CO(C[351]) );
  FA_12249 \FA_INST_0[0].FA_INST_1[351].FA_  ( .A(A[351]), .B(n1376), .CI(
        C[351]), .S(S[351]), .CO(C[352]) );
  FA_12248 \FA_INST_0[0].FA_INST_1[352].FA_  ( .A(A[352]), .B(n1377), .CI(
        C[352]), .S(S[352]), .CO(C[353]) );
  FA_12247 \FA_INST_0[0].FA_INST_1[353].FA_  ( .A(A[353]), .B(n1378), .CI(
        C[353]), .S(S[353]), .CO(C[354]) );
  FA_12246 \FA_INST_0[0].FA_INST_1[354].FA_  ( .A(A[354]), .B(n1379), .CI(
        C[354]), .S(S[354]), .CO(C[355]) );
  FA_12245 \FA_INST_0[0].FA_INST_1[355].FA_  ( .A(A[355]), .B(n1380), .CI(
        C[355]), .S(S[355]), .CO(C[356]) );
  FA_12244 \FA_INST_0[0].FA_INST_1[356].FA_  ( .A(A[356]), .B(n1381), .CI(
        C[356]), .S(S[356]), .CO(C[357]) );
  FA_12243 \FA_INST_0[0].FA_INST_1[357].FA_  ( .A(A[357]), .B(n1382), .CI(
        C[357]), .S(S[357]), .CO(C[358]) );
  FA_12242 \FA_INST_0[0].FA_INST_1[358].FA_  ( .A(A[358]), .B(n1383), .CI(
        C[358]), .S(S[358]), .CO(C[359]) );
  FA_12241 \FA_INST_0[0].FA_INST_1[359].FA_  ( .A(A[359]), .B(n1384), .CI(
        C[359]), .S(S[359]), .CO(C[360]) );
  FA_12240 \FA_INST_0[0].FA_INST_1[360].FA_  ( .A(A[360]), .B(n1385), .CI(
        C[360]), .S(S[360]), .CO(C[361]) );
  FA_12239 \FA_INST_0[0].FA_INST_1[361].FA_  ( .A(A[361]), .B(n1386), .CI(
        C[361]), .S(S[361]), .CO(C[362]) );
  FA_12238 \FA_INST_0[0].FA_INST_1[362].FA_  ( .A(A[362]), .B(n1387), .CI(
        C[362]), .S(S[362]), .CO(C[363]) );
  FA_12237 \FA_INST_0[0].FA_INST_1[363].FA_  ( .A(A[363]), .B(n1388), .CI(
        C[363]), .S(S[363]), .CO(C[364]) );
  FA_12236 \FA_INST_0[0].FA_INST_1[364].FA_  ( .A(A[364]), .B(n1389), .CI(
        C[364]), .S(S[364]), .CO(C[365]) );
  FA_12235 \FA_INST_0[0].FA_INST_1[365].FA_  ( .A(A[365]), .B(n1390), .CI(
        C[365]), .S(S[365]), .CO(C[366]) );
  FA_12234 \FA_INST_0[0].FA_INST_1[366].FA_  ( .A(A[366]), .B(n1391), .CI(
        C[366]), .S(S[366]), .CO(C[367]) );
  FA_12233 \FA_INST_0[0].FA_INST_1[367].FA_  ( .A(A[367]), .B(n1392), .CI(
        C[367]), .S(S[367]), .CO(C[368]) );
  FA_12232 \FA_INST_0[0].FA_INST_1[368].FA_  ( .A(A[368]), .B(n1393), .CI(
        C[368]), .S(S[368]), .CO(C[369]) );
  FA_12231 \FA_INST_0[0].FA_INST_1[369].FA_  ( .A(A[369]), .B(n1394), .CI(
        C[369]), .S(S[369]), .CO(C[370]) );
  FA_12230 \FA_INST_0[0].FA_INST_1[370].FA_  ( .A(A[370]), .B(n1395), .CI(
        C[370]), .S(S[370]), .CO(C[371]) );
  FA_12229 \FA_INST_0[0].FA_INST_1[371].FA_  ( .A(A[371]), .B(n1396), .CI(
        C[371]), .S(S[371]), .CO(C[372]) );
  FA_12228 \FA_INST_0[0].FA_INST_1[372].FA_  ( .A(A[372]), .B(n1397), .CI(
        C[372]), .S(S[372]), .CO(C[373]) );
  FA_12227 \FA_INST_0[0].FA_INST_1[373].FA_  ( .A(A[373]), .B(n1398), .CI(
        C[373]), .S(S[373]), .CO(C[374]) );
  FA_12226 \FA_INST_0[0].FA_INST_1[374].FA_  ( .A(A[374]), .B(n1399), .CI(
        C[374]), .S(S[374]), .CO(C[375]) );
  FA_12225 \FA_INST_0[0].FA_INST_1[375].FA_  ( .A(A[375]), .B(n1400), .CI(
        C[375]), .S(S[375]), .CO(C[376]) );
  FA_12224 \FA_INST_0[0].FA_INST_1[376].FA_  ( .A(A[376]), .B(n1401), .CI(
        C[376]), .S(S[376]), .CO(C[377]) );
  FA_12223 \FA_INST_0[0].FA_INST_1[377].FA_  ( .A(A[377]), .B(n1402), .CI(
        C[377]), .S(S[377]), .CO(C[378]) );
  FA_12222 \FA_INST_0[0].FA_INST_1[378].FA_  ( .A(A[378]), .B(n1403), .CI(
        C[378]), .S(S[378]), .CO(C[379]) );
  FA_12221 \FA_INST_0[0].FA_INST_1[379].FA_  ( .A(A[379]), .B(n1404), .CI(
        C[379]), .S(S[379]), .CO(C[380]) );
  FA_12220 \FA_INST_0[0].FA_INST_1[380].FA_  ( .A(A[380]), .B(n1405), .CI(
        C[380]), .S(S[380]), .CO(C[381]) );
  FA_12219 \FA_INST_0[0].FA_INST_1[381].FA_  ( .A(A[381]), .B(n1406), .CI(
        C[381]), .S(S[381]), .CO(C[382]) );
  FA_12218 \FA_INST_0[0].FA_INST_1[382].FA_  ( .A(A[382]), .B(n1407), .CI(
        C[382]), .S(S[382]), .CO(C[383]) );
  FA_12217 \FA_INST_0[0].FA_INST_1[383].FA_  ( .A(A[383]), .B(n1408), .CI(
        C[383]), .S(S[383]), .CO(C[384]) );
  FA_12216 \FA_INST_0[0].FA_INST_1[384].FA_  ( .A(A[384]), .B(n1409), .CI(
        C[384]), .S(S[384]), .CO(C[385]) );
  FA_12215 \FA_INST_0[0].FA_INST_1[385].FA_  ( .A(A[385]), .B(n1410), .CI(
        C[385]), .S(S[385]), .CO(C[386]) );
  FA_12214 \FA_INST_0[0].FA_INST_1[386].FA_  ( .A(A[386]), .B(n1411), .CI(
        C[386]), .S(S[386]), .CO(C[387]) );
  FA_12213 \FA_INST_0[0].FA_INST_1[387].FA_  ( .A(A[387]), .B(n1412), .CI(
        C[387]), .S(S[387]), .CO(C[388]) );
  FA_12212 \FA_INST_0[0].FA_INST_1[388].FA_  ( .A(A[388]), .B(n1413), .CI(
        C[388]), .S(S[388]), .CO(C[389]) );
  FA_12211 \FA_INST_0[0].FA_INST_1[389].FA_  ( .A(A[389]), .B(n1414), .CI(
        C[389]), .S(S[389]), .CO(C[390]) );
  FA_12210 \FA_INST_0[0].FA_INST_1[390].FA_  ( .A(A[390]), .B(n1415), .CI(
        C[390]), .S(S[390]), .CO(C[391]) );
  FA_12209 \FA_INST_0[0].FA_INST_1[391].FA_  ( .A(A[391]), .B(n1416), .CI(
        C[391]), .S(S[391]), .CO(C[392]) );
  FA_12208 \FA_INST_0[0].FA_INST_1[392].FA_  ( .A(A[392]), .B(n1417), .CI(
        C[392]), .S(S[392]), .CO(C[393]) );
  FA_12207 \FA_INST_0[0].FA_INST_1[393].FA_  ( .A(A[393]), .B(n1418), .CI(
        C[393]), .S(S[393]), .CO(C[394]) );
  FA_12206 \FA_INST_0[0].FA_INST_1[394].FA_  ( .A(A[394]), .B(n1419), .CI(
        C[394]), .S(S[394]), .CO(C[395]) );
  FA_12205 \FA_INST_0[0].FA_INST_1[395].FA_  ( .A(A[395]), .B(n1420), .CI(
        C[395]), .S(S[395]), .CO(C[396]) );
  FA_12204 \FA_INST_0[0].FA_INST_1[396].FA_  ( .A(A[396]), .B(n1421), .CI(
        C[396]), .S(S[396]), .CO(C[397]) );
  FA_12203 \FA_INST_0[0].FA_INST_1[397].FA_  ( .A(A[397]), .B(n1422), .CI(
        C[397]), .S(S[397]), .CO(C[398]) );
  FA_12202 \FA_INST_0[0].FA_INST_1[398].FA_  ( .A(A[398]), .B(n1423), .CI(
        C[398]), .S(S[398]), .CO(C[399]) );
  FA_12201 \FA_INST_0[0].FA_INST_1[399].FA_  ( .A(A[399]), .B(n1424), .CI(
        C[399]), .S(S[399]), .CO(C[400]) );
  FA_12200 \FA_INST_0[0].FA_INST_1[400].FA_  ( .A(A[400]), .B(n1425), .CI(
        C[400]), .S(S[400]), .CO(C[401]) );
  FA_12199 \FA_INST_0[0].FA_INST_1[401].FA_  ( .A(A[401]), .B(n1426), .CI(
        C[401]), .S(S[401]), .CO(C[402]) );
  FA_12198 \FA_INST_0[0].FA_INST_1[402].FA_  ( .A(A[402]), .B(n1427), .CI(
        C[402]), .S(S[402]), .CO(C[403]) );
  FA_12197 \FA_INST_0[0].FA_INST_1[403].FA_  ( .A(A[403]), .B(n1428), .CI(
        C[403]), .S(S[403]), .CO(C[404]) );
  FA_12196 \FA_INST_0[0].FA_INST_1[404].FA_  ( .A(A[404]), .B(n1429), .CI(
        C[404]), .S(S[404]), .CO(C[405]) );
  FA_12195 \FA_INST_0[0].FA_INST_1[405].FA_  ( .A(A[405]), .B(n1430), .CI(
        C[405]), .S(S[405]), .CO(C[406]) );
  FA_12194 \FA_INST_0[0].FA_INST_1[406].FA_  ( .A(A[406]), .B(n1431), .CI(
        C[406]), .S(S[406]), .CO(C[407]) );
  FA_12193 \FA_INST_0[0].FA_INST_1[407].FA_  ( .A(A[407]), .B(n1432), .CI(
        C[407]), .S(S[407]), .CO(C[408]) );
  FA_12192 \FA_INST_0[0].FA_INST_1[408].FA_  ( .A(A[408]), .B(n1433), .CI(
        C[408]), .S(S[408]), .CO(C[409]) );
  FA_12191 \FA_INST_0[0].FA_INST_1[409].FA_  ( .A(A[409]), .B(n1434), .CI(
        C[409]), .S(S[409]), .CO(C[410]) );
  FA_12190 \FA_INST_0[0].FA_INST_1[410].FA_  ( .A(A[410]), .B(n1435), .CI(
        C[410]), .S(S[410]), .CO(C[411]) );
  FA_12189 \FA_INST_0[0].FA_INST_1[411].FA_  ( .A(A[411]), .B(n1436), .CI(
        C[411]), .S(S[411]), .CO(C[412]) );
  FA_12188 \FA_INST_0[0].FA_INST_1[412].FA_  ( .A(A[412]), .B(n1437), .CI(
        C[412]), .S(S[412]), .CO(C[413]) );
  FA_12187 \FA_INST_0[0].FA_INST_1[413].FA_  ( .A(A[413]), .B(n1438), .CI(
        C[413]), .S(S[413]), .CO(C[414]) );
  FA_12186 \FA_INST_0[0].FA_INST_1[414].FA_  ( .A(A[414]), .B(n1439), .CI(
        C[414]), .S(S[414]), .CO(C[415]) );
  FA_12185 \FA_INST_0[0].FA_INST_1[415].FA_  ( .A(A[415]), .B(n1440), .CI(
        C[415]), .S(S[415]), .CO(C[416]) );
  FA_12184 \FA_INST_0[0].FA_INST_1[416].FA_  ( .A(A[416]), .B(n1441), .CI(
        C[416]), .S(S[416]), .CO(C[417]) );
  FA_12183 \FA_INST_0[0].FA_INST_1[417].FA_  ( .A(A[417]), .B(n1442), .CI(
        C[417]), .S(S[417]), .CO(C[418]) );
  FA_12182 \FA_INST_0[0].FA_INST_1[418].FA_  ( .A(A[418]), .B(n1443), .CI(
        C[418]), .S(S[418]), .CO(C[419]) );
  FA_12181 \FA_INST_0[0].FA_INST_1[419].FA_  ( .A(A[419]), .B(n1444), .CI(
        C[419]), .S(S[419]), .CO(C[420]) );
  FA_12180 \FA_INST_0[0].FA_INST_1[420].FA_  ( .A(A[420]), .B(n1445), .CI(
        C[420]), .S(S[420]), .CO(C[421]) );
  FA_12179 \FA_INST_0[0].FA_INST_1[421].FA_  ( .A(A[421]), .B(n1446), .CI(
        C[421]), .S(S[421]), .CO(C[422]) );
  FA_12178 \FA_INST_0[0].FA_INST_1[422].FA_  ( .A(A[422]), .B(n1447), .CI(
        C[422]), .S(S[422]), .CO(C[423]) );
  FA_12177 \FA_INST_0[0].FA_INST_1[423].FA_  ( .A(A[423]), .B(n1448), .CI(
        C[423]), .S(S[423]), .CO(C[424]) );
  FA_12176 \FA_INST_0[0].FA_INST_1[424].FA_  ( .A(A[424]), .B(n1449), .CI(
        C[424]), .S(S[424]), .CO(C[425]) );
  FA_12175 \FA_INST_0[0].FA_INST_1[425].FA_  ( .A(A[425]), .B(n1450), .CI(
        C[425]), .S(S[425]), .CO(C[426]) );
  FA_12174 \FA_INST_0[0].FA_INST_1[426].FA_  ( .A(A[426]), .B(n1451), .CI(
        C[426]), .S(S[426]), .CO(C[427]) );
  FA_12173 \FA_INST_0[0].FA_INST_1[427].FA_  ( .A(A[427]), .B(n1452), .CI(
        C[427]), .S(S[427]), .CO(C[428]) );
  FA_12172 \FA_INST_0[0].FA_INST_1[428].FA_  ( .A(A[428]), .B(n1453), .CI(
        C[428]), .S(S[428]), .CO(C[429]) );
  FA_12171 \FA_INST_0[0].FA_INST_1[429].FA_  ( .A(A[429]), .B(n1454), .CI(
        C[429]), .S(S[429]), .CO(C[430]) );
  FA_12170 \FA_INST_0[0].FA_INST_1[430].FA_  ( .A(A[430]), .B(n1455), .CI(
        C[430]), .S(S[430]), .CO(C[431]) );
  FA_12169 \FA_INST_0[0].FA_INST_1[431].FA_  ( .A(A[431]), .B(n1456), .CI(
        C[431]), .S(S[431]), .CO(C[432]) );
  FA_12168 \FA_INST_0[0].FA_INST_1[432].FA_  ( .A(A[432]), .B(n1457), .CI(
        C[432]), .S(S[432]), .CO(C[433]) );
  FA_12167 \FA_INST_0[0].FA_INST_1[433].FA_  ( .A(A[433]), .B(n1458), .CI(
        C[433]), .S(S[433]), .CO(C[434]) );
  FA_12166 \FA_INST_0[0].FA_INST_1[434].FA_  ( .A(A[434]), .B(n1459), .CI(
        C[434]), .S(S[434]), .CO(C[435]) );
  FA_12165 \FA_INST_0[0].FA_INST_1[435].FA_  ( .A(A[435]), .B(n1460), .CI(
        C[435]), .S(S[435]), .CO(C[436]) );
  FA_12164 \FA_INST_0[0].FA_INST_1[436].FA_  ( .A(A[436]), .B(n1461), .CI(
        C[436]), .S(S[436]), .CO(C[437]) );
  FA_12163 \FA_INST_0[0].FA_INST_1[437].FA_  ( .A(A[437]), .B(n1462), .CI(
        C[437]), .S(S[437]), .CO(C[438]) );
  FA_12162 \FA_INST_0[0].FA_INST_1[438].FA_  ( .A(A[438]), .B(n1463), .CI(
        C[438]), .S(S[438]), .CO(C[439]) );
  FA_12161 \FA_INST_0[0].FA_INST_1[439].FA_  ( .A(A[439]), .B(n1464), .CI(
        C[439]), .S(S[439]), .CO(C[440]) );
  FA_12160 \FA_INST_0[0].FA_INST_1[440].FA_  ( .A(A[440]), .B(n1465), .CI(
        C[440]), .S(S[440]), .CO(C[441]) );
  FA_12159 \FA_INST_0[0].FA_INST_1[441].FA_  ( .A(A[441]), .B(n1466), .CI(
        C[441]), .S(S[441]), .CO(C[442]) );
  FA_12158 \FA_INST_0[0].FA_INST_1[442].FA_  ( .A(A[442]), .B(n1467), .CI(
        C[442]), .S(S[442]), .CO(C[443]) );
  FA_12157 \FA_INST_0[0].FA_INST_1[443].FA_  ( .A(A[443]), .B(n1468), .CI(
        C[443]), .S(S[443]), .CO(C[444]) );
  FA_12156 \FA_INST_0[0].FA_INST_1[444].FA_  ( .A(A[444]), .B(n1469), .CI(
        C[444]), .S(S[444]), .CO(C[445]) );
  FA_12155 \FA_INST_0[0].FA_INST_1[445].FA_  ( .A(A[445]), .B(n1470), .CI(
        C[445]), .S(S[445]), .CO(C[446]) );
  FA_12154 \FA_INST_0[0].FA_INST_1[446].FA_  ( .A(A[446]), .B(n1471), .CI(
        C[446]), .S(S[446]), .CO(C[447]) );
  FA_12153 \FA_INST_0[0].FA_INST_1[447].FA_  ( .A(A[447]), .B(n1472), .CI(
        C[447]), .S(S[447]), .CO(C[448]) );
  FA_12152 \FA_INST_0[0].FA_INST_1[448].FA_  ( .A(A[448]), .B(n1473), .CI(
        C[448]), .S(S[448]), .CO(C[449]) );
  FA_12151 \FA_INST_0[0].FA_INST_1[449].FA_  ( .A(A[449]), .B(n1474), .CI(
        C[449]), .S(S[449]), .CO(C[450]) );
  FA_12150 \FA_INST_0[0].FA_INST_1[450].FA_  ( .A(A[450]), .B(n1475), .CI(
        C[450]), .S(S[450]), .CO(C[451]) );
  FA_12149 \FA_INST_0[0].FA_INST_1[451].FA_  ( .A(A[451]), .B(n1476), .CI(
        C[451]), .S(S[451]), .CO(C[452]) );
  FA_12148 \FA_INST_0[0].FA_INST_1[452].FA_  ( .A(A[452]), .B(n1477), .CI(
        C[452]), .S(S[452]), .CO(C[453]) );
  FA_12147 \FA_INST_0[0].FA_INST_1[453].FA_  ( .A(A[453]), .B(n1478), .CI(
        C[453]), .S(S[453]), .CO(C[454]) );
  FA_12146 \FA_INST_0[0].FA_INST_1[454].FA_  ( .A(A[454]), .B(n1479), .CI(
        C[454]), .S(S[454]), .CO(C[455]) );
  FA_12145 \FA_INST_0[0].FA_INST_1[455].FA_  ( .A(A[455]), .B(n1480), .CI(
        C[455]), .S(S[455]), .CO(C[456]) );
  FA_12144 \FA_INST_0[0].FA_INST_1[456].FA_  ( .A(A[456]), .B(n1481), .CI(
        C[456]), .S(S[456]), .CO(C[457]) );
  FA_12143 \FA_INST_0[0].FA_INST_1[457].FA_  ( .A(A[457]), .B(n1482), .CI(
        C[457]), .S(S[457]), .CO(C[458]) );
  FA_12142 \FA_INST_0[0].FA_INST_1[458].FA_  ( .A(A[458]), .B(n1483), .CI(
        C[458]), .S(S[458]), .CO(C[459]) );
  FA_12141 \FA_INST_0[0].FA_INST_1[459].FA_  ( .A(A[459]), .B(n1484), .CI(
        C[459]), .S(S[459]), .CO(C[460]) );
  FA_12140 \FA_INST_0[0].FA_INST_1[460].FA_  ( .A(A[460]), .B(n1485), .CI(
        C[460]), .S(S[460]), .CO(C[461]) );
  FA_12139 \FA_INST_0[0].FA_INST_1[461].FA_  ( .A(A[461]), .B(n1486), .CI(
        C[461]), .S(S[461]), .CO(C[462]) );
  FA_12138 \FA_INST_0[0].FA_INST_1[462].FA_  ( .A(A[462]), .B(n1487), .CI(
        C[462]), .S(S[462]), .CO(C[463]) );
  FA_12137 \FA_INST_0[0].FA_INST_1[463].FA_  ( .A(A[463]), .B(n1488), .CI(
        C[463]), .S(S[463]), .CO(C[464]) );
  FA_12136 \FA_INST_0[0].FA_INST_1[464].FA_  ( .A(A[464]), .B(n1489), .CI(
        C[464]), .S(S[464]), .CO(C[465]) );
  FA_12135 \FA_INST_0[0].FA_INST_1[465].FA_  ( .A(A[465]), .B(n1490), .CI(
        C[465]), .S(S[465]), .CO(C[466]) );
  FA_12134 \FA_INST_0[0].FA_INST_1[466].FA_  ( .A(A[466]), .B(n1491), .CI(
        C[466]), .S(S[466]), .CO(C[467]) );
  FA_12133 \FA_INST_0[0].FA_INST_1[467].FA_  ( .A(A[467]), .B(n1492), .CI(
        C[467]), .S(S[467]), .CO(C[468]) );
  FA_12132 \FA_INST_0[0].FA_INST_1[468].FA_  ( .A(A[468]), .B(n1493), .CI(
        C[468]), .S(S[468]), .CO(C[469]) );
  FA_12131 \FA_INST_0[0].FA_INST_1[469].FA_  ( .A(A[469]), .B(n1494), .CI(
        C[469]), .S(S[469]), .CO(C[470]) );
  FA_12130 \FA_INST_0[0].FA_INST_1[470].FA_  ( .A(A[470]), .B(n1495), .CI(
        C[470]), .S(S[470]), .CO(C[471]) );
  FA_12129 \FA_INST_0[0].FA_INST_1[471].FA_  ( .A(A[471]), .B(n1496), .CI(
        C[471]), .S(S[471]), .CO(C[472]) );
  FA_12128 \FA_INST_0[0].FA_INST_1[472].FA_  ( .A(A[472]), .B(n1497), .CI(
        C[472]), .S(S[472]), .CO(C[473]) );
  FA_12127 \FA_INST_0[0].FA_INST_1[473].FA_  ( .A(A[473]), .B(n1498), .CI(
        C[473]), .S(S[473]), .CO(C[474]) );
  FA_12126 \FA_INST_0[0].FA_INST_1[474].FA_  ( .A(A[474]), .B(n1499), .CI(
        C[474]), .S(S[474]), .CO(C[475]) );
  FA_12125 \FA_INST_0[0].FA_INST_1[475].FA_  ( .A(A[475]), .B(n1500), .CI(
        C[475]), .S(S[475]), .CO(C[476]) );
  FA_12124 \FA_INST_0[0].FA_INST_1[476].FA_  ( .A(A[476]), .B(n1501), .CI(
        C[476]), .S(S[476]), .CO(C[477]) );
  FA_12123 \FA_INST_0[0].FA_INST_1[477].FA_  ( .A(A[477]), .B(n1502), .CI(
        C[477]), .S(S[477]), .CO(C[478]) );
  FA_12122 \FA_INST_0[0].FA_INST_1[478].FA_  ( .A(A[478]), .B(n1503), .CI(
        C[478]), .S(S[478]), .CO(C[479]) );
  FA_12121 \FA_INST_0[0].FA_INST_1[479].FA_  ( .A(A[479]), .B(n1504), .CI(
        C[479]), .S(S[479]), .CO(C[480]) );
  FA_12120 \FA_INST_0[0].FA_INST_1[480].FA_  ( .A(A[480]), .B(n1505), .CI(
        C[480]), .S(S[480]), .CO(C[481]) );
  FA_12119 \FA_INST_0[0].FA_INST_1[481].FA_  ( .A(A[481]), .B(n1506), .CI(
        C[481]), .S(S[481]), .CO(C[482]) );
  FA_12118 \FA_INST_0[0].FA_INST_1[482].FA_  ( .A(A[482]), .B(n1507), .CI(
        C[482]), .S(S[482]), .CO(C[483]) );
  FA_12117 \FA_INST_0[0].FA_INST_1[483].FA_  ( .A(A[483]), .B(n1508), .CI(
        C[483]), .S(S[483]), .CO(C[484]) );
  FA_12116 \FA_INST_0[0].FA_INST_1[484].FA_  ( .A(A[484]), .B(n1509), .CI(
        C[484]), .S(S[484]), .CO(C[485]) );
  FA_12115 \FA_INST_0[0].FA_INST_1[485].FA_  ( .A(A[485]), .B(n1510), .CI(
        C[485]), .S(S[485]), .CO(C[486]) );
  FA_12114 \FA_INST_0[0].FA_INST_1[486].FA_  ( .A(A[486]), .B(n1511), .CI(
        C[486]), .S(S[486]), .CO(C[487]) );
  FA_12113 \FA_INST_0[0].FA_INST_1[487].FA_  ( .A(A[487]), .B(n1512), .CI(
        C[487]), .S(S[487]), .CO(C[488]) );
  FA_12112 \FA_INST_0[0].FA_INST_1[488].FA_  ( .A(A[488]), .B(n1513), .CI(
        C[488]), .S(S[488]), .CO(C[489]) );
  FA_12111 \FA_INST_0[0].FA_INST_1[489].FA_  ( .A(A[489]), .B(n1514), .CI(
        C[489]), .S(S[489]), .CO(C[490]) );
  FA_12110 \FA_INST_0[0].FA_INST_1[490].FA_  ( .A(A[490]), .B(n1515), .CI(
        C[490]), .S(S[490]), .CO(C[491]) );
  FA_12109 \FA_INST_0[0].FA_INST_1[491].FA_  ( .A(A[491]), .B(n1516), .CI(
        C[491]), .S(S[491]), .CO(C[492]) );
  FA_12108 \FA_INST_0[0].FA_INST_1[492].FA_  ( .A(A[492]), .B(n1517), .CI(
        C[492]), .S(S[492]), .CO(C[493]) );
  FA_12107 \FA_INST_0[0].FA_INST_1[493].FA_  ( .A(A[493]), .B(n1518), .CI(
        C[493]), .S(S[493]), .CO(C[494]) );
  FA_12106 \FA_INST_0[0].FA_INST_1[494].FA_  ( .A(A[494]), .B(n1519), .CI(
        C[494]), .S(S[494]), .CO(C[495]) );
  FA_12105 \FA_INST_0[0].FA_INST_1[495].FA_  ( .A(A[495]), .B(n1520), .CI(
        C[495]), .S(S[495]), .CO(C[496]) );
  FA_12104 \FA_INST_0[0].FA_INST_1[496].FA_  ( .A(A[496]), .B(n1521), .CI(
        C[496]), .S(S[496]), .CO(C[497]) );
  FA_12103 \FA_INST_0[0].FA_INST_1[497].FA_  ( .A(A[497]), .B(n1522), .CI(
        C[497]), .S(S[497]), .CO(C[498]) );
  FA_12102 \FA_INST_0[0].FA_INST_1[498].FA_  ( .A(A[498]), .B(n1523), .CI(
        C[498]), .S(S[498]), .CO(C[499]) );
  FA_12101 \FA_INST_0[0].FA_INST_1[499].FA_  ( .A(A[499]), .B(n1524), .CI(
        C[499]), .S(S[499]), .CO(C[500]) );
  FA_12100 \FA_INST_0[0].FA_INST_1[500].FA_  ( .A(A[500]), .B(n1525), .CI(
        C[500]), .S(S[500]), .CO(C[501]) );
  FA_12099 \FA_INST_0[0].FA_INST_1[501].FA_  ( .A(A[501]), .B(n1526), .CI(
        C[501]), .S(S[501]), .CO(C[502]) );
  FA_12098 \FA_INST_0[0].FA_INST_1[502].FA_  ( .A(A[502]), .B(n1527), .CI(
        C[502]), .S(S[502]), .CO(C[503]) );
  FA_12097 \FA_INST_0[0].FA_INST_1[503].FA_  ( .A(A[503]), .B(n1528), .CI(
        C[503]), .S(S[503]), .CO(C[504]) );
  FA_12096 \FA_INST_0[0].FA_INST_1[504].FA_  ( .A(A[504]), .B(n1529), .CI(
        C[504]), .S(S[504]), .CO(C[505]) );
  FA_12095 \FA_INST_0[0].FA_INST_1[505].FA_  ( .A(A[505]), .B(n1530), .CI(
        C[505]), .S(S[505]), .CO(C[506]) );
  FA_12094 \FA_INST_0[0].FA_INST_1[506].FA_  ( .A(A[506]), .B(n1531), .CI(
        C[506]), .S(S[506]), .CO(C[507]) );
  FA_12093 \FA_INST_0[0].FA_INST_1[507].FA_  ( .A(A[507]), .B(n1532), .CI(
        C[507]), .S(S[507]), .CO(C[508]) );
  FA_12092 \FA_INST_0[0].FA_INST_1[508].FA_  ( .A(A[508]), .B(n1533), .CI(
        C[508]), .S(S[508]), .CO(C[509]) );
  FA_12091 \FA_INST_0[0].FA_INST_1[509].FA_  ( .A(A[509]), .B(n1534), .CI(
        C[509]), .S(S[509]), .CO(C[510]) );
  FA_12090 \FA_INST_0[0].FA_INST_1[510].FA_  ( .A(A[510]), .B(n1535), .CI(
        C[510]), .S(S[510]), .CO(C[511]) );
  FA_12089 \FA_INST_0[0].FA_INST_1[511].FA_  ( .A(A[511]), .B(n1536), .CI(
        C[511]), .S(S[511]), .CO(C[512]) );
  FA_12088 \FA_INST_0[1].FA_INST_1[0].FA_  ( .A(A[512]), .B(n1537), .CI(C[512]), .S(S[512]), .CO(C[513]) );
  FA_12087 \FA_INST_0[1].FA_INST_1[1].FA_  ( .A(A[513]), .B(n1538), .CI(C[513]), .S(S[513]), .CO(C[514]) );
  FA_12086 \FA_INST_0[1].FA_INST_1[2].FA_  ( .A(A[514]), .B(n1539), .CI(C[514]), .S(S[514]), .CO(C[515]) );
  FA_12085 \FA_INST_0[1].FA_INST_1[3].FA_  ( .A(A[515]), .B(n1540), .CI(C[515]), .S(S[515]), .CO(C[516]) );
  FA_12084 \FA_INST_0[1].FA_INST_1[4].FA_  ( .A(A[516]), .B(n1541), .CI(C[516]), .S(S[516]), .CO(C[517]) );
  FA_12083 \FA_INST_0[1].FA_INST_1[5].FA_  ( .A(A[517]), .B(n1542), .CI(C[517]), .S(S[517]), .CO(C[518]) );
  FA_12082 \FA_INST_0[1].FA_INST_1[6].FA_  ( .A(A[518]), .B(n1543), .CI(C[518]), .S(S[518]), .CO(C[519]) );
  FA_12081 \FA_INST_0[1].FA_INST_1[7].FA_  ( .A(A[519]), .B(n1544), .CI(C[519]), .S(S[519]), .CO(C[520]) );
  FA_12080 \FA_INST_0[1].FA_INST_1[8].FA_  ( .A(A[520]), .B(n1545), .CI(C[520]), .S(S[520]), .CO(C[521]) );
  FA_12079 \FA_INST_0[1].FA_INST_1[9].FA_  ( .A(A[521]), .B(n1546), .CI(C[521]), .S(S[521]), .CO(C[522]) );
  FA_12078 \FA_INST_0[1].FA_INST_1[10].FA_  ( .A(A[522]), .B(n1547), .CI(
        C[522]), .S(S[522]), .CO(C[523]) );
  FA_12077 \FA_INST_0[1].FA_INST_1[11].FA_  ( .A(A[523]), .B(n1548), .CI(
        C[523]), .S(S[523]), .CO(C[524]) );
  FA_12076 \FA_INST_0[1].FA_INST_1[12].FA_  ( .A(A[524]), .B(n1549), .CI(
        C[524]), .S(S[524]), .CO(C[525]) );
  FA_12075 \FA_INST_0[1].FA_INST_1[13].FA_  ( .A(A[525]), .B(n1550), .CI(
        C[525]), .S(S[525]), .CO(C[526]) );
  FA_12074 \FA_INST_0[1].FA_INST_1[14].FA_  ( .A(A[526]), .B(n1551), .CI(
        C[526]), .S(S[526]), .CO(C[527]) );
  FA_12073 \FA_INST_0[1].FA_INST_1[15].FA_  ( .A(A[527]), .B(n1552), .CI(
        C[527]), .S(S[527]), .CO(C[528]) );
  FA_12072 \FA_INST_0[1].FA_INST_1[16].FA_  ( .A(A[528]), .B(n1553), .CI(
        C[528]), .S(S[528]), .CO(C[529]) );
  FA_12071 \FA_INST_0[1].FA_INST_1[17].FA_  ( .A(A[529]), .B(n1554), .CI(
        C[529]), .S(S[529]), .CO(C[530]) );
  FA_12070 \FA_INST_0[1].FA_INST_1[18].FA_  ( .A(A[530]), .B(n1555), .CI(
        C[530]), .S(S[530]), .CO(C[531]) );
  FA_12069 \FA_INST_0[1].FA_INST_1[19].FA_  ( .A(A[531]), .B(n1556), .CI(
        C[531]), .S(S[531]), .CO(C[532]) );
  FA_12068 \FA_INST_0[1].FA_INST_1[20].FA_  ( .A(A[532]), .B(n1557), .CI(
        C[532]), .S(S[532]), .CO(C[533]) );
  FA_12067 \FA_INST_0[1].FA_INST_1[21].FA_  ( .A(A[533]), .B(n1558), .CI(
        C[533]), .S(S[533]), .CO(C[534]) );
  FA_12066 \FA_INST_0[1].FA_INST_1[22].FA_  ( .A(A[534]), .B(n1559), .CI(
        C[534]), .S(S[534]), .CO(C[535]) );
  FA_12065 \FA_INST_0[1].FA_INST_1[23].FA_  ( .A(A[535]), .B(n1560), .CI(
        C[535]), .S(S[535]), .CO(C[536]) );
  FA_12064 \FA_INST_0[1].FA_INST_1[24].FA_  ( .A(A[536]), .B(n1561), .CI(
        C[536]), .S(S[536]), .CO(C[537]) );
  FA_12063 \FA_INST_0[1].FA_INST_1[25].FA_  ( .A(A[537]), .B(n1562), .CI(
        C[537]), .S(S[537]), .CO(C[538]) );
  FA_12062 \FA_INST_0[1].FA_INST_1[26].FA_  ( .A(A[538]), .B(n1563), .CI(
        C[538]), .S(S[538]), .CO(C[539]) );
  FA_12061 \FA_INST_0[1].FA_INST_1[27].FA_  ( .A(A[539]), .B(n1564), .CI(
        C[539]), .S(S[539]), .CO(C[540]) );
  FA_12060 \FA_INST_0[1].FA_INST_1[28].FA_  ( .A(A[540]), .B(n1565), .CI(
        C[540]), .S(S[540]), .CO(C[541]) );
  FA_12059 \FA_INST_0[1].FA_INST_1[29].FA_  ( .A(A[541]), .B(n1566), .CI(
        C[541]), .S(S[541]), .CO(C[542]) );
  FA_12058 \FA_INST_0[1].FA_INST_1[30].FA_  ( .A(A[542]), .B(n1567), .CI(
        C[542]), .S(S[542]), .CO(C[543]) );
  FA_12057 \FA_INST_0[1].FA_INST_1[31].FA_  ( .A(A[543]), .B(n1568), .CI(
        C[543]), .S(S[543]), .CO(C[544]) );
  FA_12056 \FA_INST_0[1].FA_INST_1[32].FA_  ( .A(A[544]), .B(n1569), .CI(
        C[544]), .S(S[544]), .CO(C[545]) );
  FA_12055 \FA_INST_0[1].FA_INST_1[33].FA_  ( .A(A[545]), .B(n1570), .CI(
        C[545]), .S(S[545]), .CO(C[546]) );
  FA_12054 \FA_INST_0[1].FA_INST_1[34].FA_  ( .A(A[546]), .B(n1571), .CI(
        C[546]), .S(S[546]), .CO(C[547]) );
  FA_12053 \FA_INST_0[1].FA_INST_1[35].FA_  ( .A(A[547]), .B(n1572), .CI(
        C[547]), .S(S[547]), .CO(C[548]) );
  FA_12052 \FA_INST_0[1].FA_INST_1[36].FA_  ( .A(A[548]), .B(n1573), .CI(
        C[548]), .S(S[548]), .CO(C[549]) );
  FA_12051 \FA_INST_0[1].FA_INST_1[37].FA_  ( .A(A[549]), .B(n1574), .CI(
        C[549]), .S(S[549]), .CO(C[550]) );
  FA_12050 \FA_INST_0[1].FA_INST_1[38].FA_  ( .A(A[550]), .B(n1575), .CI(
        C[550]), .S(S[550]), .CO(C[551]) );
  FA_12049 \FA_INST_0[1].FA_INST_1[39].FA_  ( .A(A[551]), .B(n1576), .CI(
        C[551]), .S(S[551]), .CO(C[552]) );
  FA_12048 \FA_INST_0[1].FA_INST_1[40].FA_  ( .A(A[552]), .B(n1577), .CI(
        C[552]), .S(S[552]), .CO(C[553]) );
  FA_12047 \FA_INST_0[1].FA_INST_1[41].FA_  ( .A(A[553]), .B(n1578), .CI(
        C[553]), .S(S[553]), .CO(C[554]) );
  FA_12046 \FA_INST_0[1].FA_INST_1[42].FA_  ( .A(A[554]), .B(n1579), .CI(
        C[554]), .S(S[554]), .CO(C[555]) );
  FA_12045 \FA_INST_0[1].FA_INST_1[43].FA_  ( .A(A[555]), .B(n1580), .CI(
        C[555]), .S(S[555]), .CO(C[556]) );
  FA_12044 \FA_INST_0[1].FA_INST_1[44].FA_  ( .A(A[556]), .B(n1581), .CI(
        C[556]), .S(S[556]), .CO(C[557]) );
  FA_12043 \FA_INST_0[1].FA_INST_1[45].FA_  ( .A(A[557]), .B(n1582), .CI(
        C[557]), .S(S[557]), .CO(C[558]) );
  FA_12042 \FA_INST_0[1].FA_INST_1[46].FA_  ( .A(A[558]), .B(n1583), .CI(
        C[558]), .S(S[558]), .CO(C[559]) );
  FA_12041 \FA_INST_0[1].FA_INST_1[47].FA_  ( .A(A[559]), .B(n1584), .CI(
        C[559]), .S(S[559]), .CO(C[560]) );
  FA_12040 \FA_INST_0[1].FA_INST_1[48].FA_  ( .A(A[560]), .B(n1585), .CI(
        C[560]), .S(S[560]), .CO(C[561]) );
  FA_12039 \FA_INST_0[1].FA_INST_1[49].FA_  ( .A(A[561]), .B(n1586), .CI(
        C[561]), .S(S[561]), .CO(C[562]) );
  FA_12038 \FA_INST_0[1].FA_INST_1[50].FA_  ( .A(A[562]), .B(n1587), .CI(
        C[562]), .S(S[562]), .CO(C[563]) );
  FA_12037 \FA_INST_0[1].FA_INST_1[51].FA_  ( .A(A[563]), .B(n1588), .CI(
        C[563]), .S(S[563]), .CO(C[564]) );
  FA_12036 \FA_INST_0[1].FA_INST_1[52].FA_  ( .A(A[564]), .B(n1589), .CI(
        C[564]), .S(S[564]), .CO(C[565]) );
  FA_12035 \FA_INST_0[1].FA_INST_1[53].FA_  ( .A(A[565]), .B(n1590), .CI(
        C[565]), .S(S[565]), .CO(C[566]) );
  FA_12034 \FA_INST_0[1].FA_INST_1[54].FA_  ( .A(A[566]), .B(n1591), .CI(
        C[566]), .S(S[566]), .CO(C[567]) );
  FA_12033 \FA_INST_0[1].FA_INST_1[55].FA_  ( .A(A[567]), .B(n1592), .CI(
        C[567]), .S(S[567]), .CO(C[568]) );
  FA_12032 \FA_INST_0[1].FA_INST_1[56].FA_  ( .A(A[568]), .B(n1593), .CI(
        C[568]), .S(S[568]), .CO(C[569]) );
  FA_12031 \FA_INST_0[1].FA_INST_1[57].FA_  ( .A(A[569]), .B(n1594), .CI(
        C[569]), .S(S[569]), .CO(C[570]) );
  FA_12030 \FA_INST_0[1].FA_INST_1[58].FA_  ( .A(A[570]), .B(n1595), .CI(
        C[570]), .S(S[570]), .CO(C[571]) );
  FA_12029 \FA_INST_0[1].FA_INST_1[59].FA_  ( .A(A[571]), .B(n1596), .CI(
        C[571]), .S(S[571]), .CO(C[572]) );
  FA_12028 \FA_INST_0[1].FA_INST_1[60].FA_  ( .A(A[572]), .B(n1597), .CI(
        C[572]), .S(S[572]), .CO(C[573]) );
  FA_12027 \FA_INST_0[1].FA_INST_1[61].FA_  ( .A(A[573]), .B(n1598), .CI(
        C[573]), .S(S[573]), .CO(C[574]) );
  FA_12026 \FA_INST_0[1].FA_INST_1[62].FA_  ( .A(A[574]), .B(n1599), .CI(
        C[574]), .S(S[574]), .CO(C[575]) );
  FA_12025 \FA_INST_0[1].FA_INST_1[63].FA_  ( .A(A[575]), .B(n1600), .CI(
        C[575]), .S(S[575]), .CO(C[576]) );
  FA_12024 \FA_INST_0[1].FA_INST_1[64].FA_  ( .A(A[576]), .B(n1601), .CI(
        C[576]), .S(S[576]), .CO(C[577]) );
  FA_12023 \FA_INST_0[1].FA_INST_1[65].FA_  ( .A(A[577]), .B(n1602), .CI(
        C[577]), .S(S[577]), .CO(C[578]) );
  FA_12022 \FA_INST_0[1].FA_INST_1[66].FA_  ( .A(A[578]), .B(n1603), .CI(
        C[578]), .S(S[578]), .CO(C[579]) );
  FA_12021 \FA_INST_0[1].FA_INST_1[67].FA_  ( .A(A[579]), .B(n1604), .CI(
        C[579]), .S(S[579]), .CO(C[580]) );
  FA_12020 \FA_INST_0[1].FA_INST_1[68].FA_  ( .A(A[580]), .B(n1605), .CI(
        C[580]), .S(S[580]), .CO(C[581]) );
  FA_12019 \FA_INST_0[1].FA_INST_1[69].FA_  ( .A(A[581]), .B(n1606), .CI(
        C[581]), .S(S[581]), .CO(C[582]) );
  FA_12018 \FA_INST_0[1].FA_INST_1[70].FA_  ( .A(A[582]), .B(n1607), .CI(
        C[582]), .S(S[582]), .CO(C[583]) );
  FA_12017 \FA_INST_0[1].FA_INST_1[71].FA_  ( .A(A[583]), .B(n1608), .CI(
        C[583]), .S(S[583]), .CO(C[584]) );
  FA_12016 \FA_INST_0[1].FA_INST_1[72].FA_  ( .A(A[584]), .B(n1609), .CI(
        C[584]), .S(S[584]), .CO(C[585]) );
  FA_12015 \FA_INST_0[1].FA_INST_1[73].FA_  ( .A(A[585]), .B(n1610), .CI(
        C[585]), .S(S[585]), .CO(C[586]) );
  FA_12014 \FA_INST_0[1].FA_INST_1[74].FA_  ( .A(A[586]), .B(n1611), .CI(
        C[586]), .S(S[586]), .CO(C[587]) );
  FA_12013 \FA_INST_0[1].FA_INST_1[75].FA_  ( .A(A[587]), .B(n1612), .CI(
        C[587]), .S(S[587]), .CO(C[588]) );
  FA_12012 \FA_INST_0[1].FA_INST_1[76].FA_  ( .A(A[588]), .B(n1613), .CI(
        C[588]), .S(S[588]), .CO(C[589]) );
  FA_12011 \FA_INST_0[1].FA_INST_1[77].FA_  ( .A(A[589]), .B(n1614), .CI(
        C[589]), .S(S[589]), .CO(C[590]) );
  FA_12010 \FA_INST_0[1].FA_INST_1[78].FA_  ( .A(A[590]), .B(n1615), .CI(
        C[590]), .S(S[590]), .CO(C[591]) );
  FA_12009 \FA_INST_0[1].FA_INST_1[79].FA_  ( .A(A[591]), .B(n1616), .CI(
        C[591]), .S(S[591]), .CO(C[592]) );
  FA_12008 \FA_INST_0[1].FA_INST_1[80].FA_  ( .A(A[592]), .B(n1617), .CI(
        C[592]), .S(S[592]), .CO(C[593]) );
  FA_12007 \FA_INST_0[1].FA_INST_1[81].FA_  ( .A(A[593]), .B(n1618), .CI(
        C[593]), .S(S[593]), .CO(C[594]) );
  FA_12006 \FA_INST_0[1].FA_INST_1[82].FA_  ( .A(A[594]), .B(n1619), .CI(
        C[594]), .S(S[594]), .CO(C[595]) );
  FA_12005 \FA_INST_0[1].FA_INST_1[83].FA_  ( .A(A[595]), .B(n1620), .CI(
        C[595]), .S(S[595]), .CO(C[596]) );
  FA_12004 \FA_INST_0[1].FA_INST_1[84].FA_  ( .A(A[596]), .B(n1621), .CI(
        C[596]), .S(S[596]), .CO(C[597]) );
  FA_12003 \FA_INST_0[1].FA_INST_1[85].FA_  ( .A(A[597]), .B(n1622), .CI(
        C[597]), .S(S[597]), .CO(C[598]) );
  FA_12002 \FA_INST_0[1].FA_INST_1[86].FA_  ( .A(A[598]), .B(n1623), .CI(
        C[598]), .S(S[598]), .CO(C[599]) );
  FA_12001 \FA_INST_0[1].FA_INST_1[87].FA_  ( .A(A[599]), .B(n1624), .CI(
        C[599]), .S(S[599]), .CO(C[600]) );
  FA_12000 \FA_INST_0[1].FA_INST_1[88].FA_  ( .A(A[600]), .B(n1625), .CI(
        C[600]), .S(S[600]), .CO(C[601]) );
  FA_11999 \FA_INST_0[1].FA_INST_1[89].FA_  ( .A(A[601]), .B(n1626), .CI(
        C[601]), .S(S[601]), .CO(C[602]) );
  FA_11998 \FA_INST_0[1].FA_INST_1[90].FA_  ( .A(A[602]), .B(n1627), .CI(
        C[602]), .S(S[602]), .CO(C[603]) );
  FA_11997 \FA_INST_0[1].FA_INST_1[91].FA_  ( .A(A[603]), .B(n1628), .CI(
        C[603]), .S(S[603]), .CO(C[604]) );
  FA_11996 \FA_INST_0[1].FA_INST_1[92].FA_  ( .A(A[604]), .B(n1629), .CI(
        C[604]), .S(S[604]), .CO(C[605]) );
  FA_11995 \FA_INST_0[1].FA_INST_1[93].FA_  ( .A(A[605]), .B(n1630), .CI(
        C[605]), .S(S[605]), .CO(C[606]) );
  FA_11994 \FA_INST_0[1].FA_INST_1[94].FA_  ( .A(A[606]), .B(n1631), .CI(
        C[606]), .S(S[606]), .CO(C[607]) );
  FA_11993 \FA_INST_0[1].FA_INST_1[95].FA_  ( .A(A[607]), .B(n1632), .CI(
        C[607]), .S(S[607]), .CO(C[608]) );
  FA_11992 \FA_INST_0[1].FA_INST_1[96].FA_  ( .A(A[608]), .B(n1633), .CI(
        C[608]), .S(S[608]), .CO(C[609]) );
  FA_11991 \FA_INST_0[1].FA_INST_1[97].FA_  ( .A(A[609]), .B(n1634), .CI(
        C[609]), .S(S[609]), .CO(C[610]) );
  FA_11990 \FA_INST_0[1].FA_INST_1[98].FA_  ( .A(A[610]), .B(n1635), .CI(
        C[610]), .S(S[610]), .CO(C[611]) );
  FA_11989 \FA_INST_0[1].FA_INST_1[99].FA_  ( .A(A[611]), .B(n1636), .CI(
        C[611]), .S(S[611]), .CO(C[612]) );
  FA_11988 \FA_INST_0[1].FA_INST_1[100].FA_  ( .A(A[612]), .B(n1637), .CI(
        C[612]), .S(S[612]), .CO(C[613]) );
  FA_11987 \FA_INST_0[1].FA_INST_1[101].FA_  ( .A(A[613]), .B(n1638), .CI(
        C[613]), .S(S[613]), .CO(C[614]) );
  FA_11986 \FA_INST_0[1].FA_INST_1[102].FA_  ( .A(A[614]), .B(n1639), .CI(
        C[614]), .S(S[614]), .CO(C[615]) );
  FA_11985 \FA_INST_0[1].FA_INST_1[103].FA_  ( .A(A[615]), .B(n1640), .CI(
        C[615]), .S(S[615]), .CO(C[616]) );
  FA_11984 \FA_INST_0[1].FA_INST_1[104].FA_  ( .A(A[616]), .B(n1641), .CI(
        C[616]), .S(S[616]), .CO(C[617]) );
  FA_11983 \FA_INST_0[1].FA_INST_1[105].FA_  ( .A(A[617]), .B(n1642), .CI(
        C[617]), .S(S[617]), .CO(C[618]) );
  FA_11982 \FA_INST_0[1].FA_INST_1[106].FA_  ( .A(A[618]), .B(n1643), .CI(
        C[618]), .S(S[618]), .CO(C[619]) );
  FA_11981 \FA_INST_0[1].FA_INST_1[107].FA_  ( .A(A[619]), .B(n1644), .CI(
        C[619]), .S(S[619]), .CO(C[620]) );
  FA_11980 \FA_INST_0[1].FA_INST_1[108].FA_  ( .A(A[620]), .B(n1645), .CI(
        C[620]), .S(S[620]), .CO(C[621]) );
  FA_11979 \FA_INST_0[1].FA_INST_1[109].FA_  ( .A(A[621]), .B(n1646), .CI(
        C[621]), .S(S[621]), .CO(C[622]) );
  FA_11978 \FA_INST_0[1].FA_INST_1[110].FA_  ( .A(A[622]), .B(n1647), .CI(
        C[622]), .S(S[622]), .CO(C[623]) );
  FA_11977 \FA_INST_0[1].FA_INST_1[111].FA_  ( .A(A[623]), .B(n1648), .CI(
        C[623]), .S(S[623]), .CO(C[624]) );
  FA_11976 \FA_INST_0[1].FA_INST_1[112].FA_  ( .A(A[624]), .B(n1649), .CI(
        C[624]), .S(S[624]), .CO(C[625]) );
  FA_11975 \FA_INST_0[1].FA_INST_1[113].FA_  ( .A(A[625]), .B(n1650), .CI(
        C[625]), .S(S[625]), .CO(C[626]) );
  FA_11974 \FA_INST_0[1].FA_INST_1[114].FA_  ( .A(A[626]), .B(n1651), .CI(
        C[626]), .S(S[626]), .CO(C[627]) );
  FA_11973 \FA_INST_0[1].FA_INST_1[115].FA_  ( .A(A[627]), .B(n1652), .CI(
        C[627]), .S(S[627]), .CO(C[628]) );
  FA_11972 \FA_INST_0[1].FA_INST_1[116].FA_  ( .A(A[628]), .B(n1653), .CI(
        C[628]), .S(S[628]), .CO(C[629]) );
  FA_11971 \FA_INST_0[1].FA_INST_1[117].FA_  ( .A(A[629]), .B(n1654), .CI(
        C[629]), .S(S[629]), .CO(C[630]) );
  FA_11970 \FA_INST_0[1].FA_INST_1[118].FA_  ( .A(A[630]), .B(n1655), .CI(
        C[630]), .S(S[630]), .CO(C[631]) );
  FA_11969 \FA_INST_0[1].FA_INST_1[119].FA_  ( .A(A[631]), .B(n1656), .CI(
        C[631]), .S(S[631]), .CO(C[632]) );
  FA_11968 \FA_INST_0[1].FA_INST_1[120].FA_  ( .A(A[632]), .B(n1657), .CI(
        C[632]), .S(S[632]), .CO(C[633]) );
  FA_11967 \FA_INST_0[1].FA_INST_1[121].FA_  ( .A(A[633]), .B(n1658), .CI(
        C[633]), .S(S[633]), .CO(C[634]) );
  FA_11966 \FA_INST_0[1].FA_INST_1[122].FA_  ( .A(A[634]), .B(n1659), .CI(
        C[634]), .S(S[634]), .CO(C[635]) );
  FA_11965 \FA_INST_0[1].FA_INST_1[123].FA_  ( .A(A[635]), .B(n1660), .CI(
        C[635]), .S(S[635]), .CO(C[636]) );
  FA_11964 \FA_INST_0[1].FA_INST_1[124].FA_  ( .A(A[636]), .B(n1661), .CI(
        C[636]), .S(S[636]), .CO(C[637]) );
  FA_11963 \FA_INST_0[1].FA_INST_1[125].FA_  ( .A(A[637]), .B(n1662), .CI(
        C[637]), .S(S[637]), .CO(C[638]) );
  FA_11962 \FA_INST_0[1].FA_INST_1[126].FA_  ( .A(A[638]), .B(n1663), .CI(
        C[638]), .S(S[638]), .CO(C[639]) );
  FA_11961 \FA_INST_0[1].FA_INST_1[127].FA_  ( .A(A[639]), .B(n1664), .CI(
        C[639]), .S(S[639]), .CO(C[640]) );
  FA_11960 \FA_INST_0[1].FA_INST_1[128].FA_  ( .A(A[640]), .B(n1665), .CI(
        C[640]), .S(S[640]), .CO(C[641]) );
  FA_11959 \FA_INST_0[1].FA_INST_1[129].FA_  ( .A(A[641]), .B(n1666), .CI(
        C[641]), .S(S[641]), .CO(C[642]) );
  FA_11958 \FA_INST_0[1].FA_INST_1[130].FA_  ( .A(A[642]), .B(n1667), .CI(
        C[642]), .S(S[642]), .CO(C[643]) );
  FA_11957 \FA_INST_0[1].FA_INST_1[131].FA_  ( .A(A[643]), .B(n1668), .CI(
        C[643]), .S(S[643]), .CO(C[644]) );
  FA_11956 \FA_INST_0[1].FA_INST_1[132].FA_  ( .A(A[644]), .B(n1669), .CI(
        C[644]), .S(S[644]), .CO(C[645]) );
  FA_11955 \FA_INST_0[1].FA_INST_1[133].FA_  ( .A(A[645]), .B(n1670), .CI(
        C[645]), .S(S[645]), .CO(C[646]) );
  FA_11954 \FA_INST_0[1].FA_INST_1[134].FA_  ( .A(A[646]), .B(n1671), .CI(
        C[646]), .S(S[646]), .CO(C[647]) );
  FA_11953 \FA_INST_0[1].FA_INST_1[135].FA_  ( .A(A[647]), .B(n1672), .CI(
        C[647]), .S(S[647]), .CO(C[648]) );
  FA_11952 \FA_INST_0[1].FA_INST_1[136].FA_  ( .A(A[648]), .B(n1673), .CI(
        C[648]), .S(S[648]), .CO(C[649]) );
  FA_11951 \FA_INST_0[1].FA_INST_1[137].FA_  ( .A(A[649]), .B(n1674), .CI(
        C[649]), .S(S[649]), .CO(C[650]) );
  FA_11950 \FA_INST_0[1].FA_INST_1[138].FA_  ( .A(A[650]), .B(n1675), .CI(
        C[650]), .S(S[650]), .CO(C[651]) );
  FA_11949 \FA_INST_0[1].FA_INST_1[139].FA_  ( .A(A[651]), .B(n1676), .CI(
        C[651]), .S(S[651]), .CO(C[652]) );
  FA_11948 \FA_INST_0[1].FA_INST_1[140].FA_  ( .A(A[652]), .B(n1677), .CI(
        C[652]), .S(S[652]), .CO(C[653]) );
  FA_11947 \FA_INST_0[1].FA_INST_1[141].FA_  ( .A(A[653]), .B(n1678), .CI(
        C[653]), .S(S[653]), .CO(C[654]) );
  FA_11946 \FA_INST_0[1].FA_INST_1[142].FA_  ( .A(A[654]), .B(n1679), .CI(
        C[654]), .S(S[654]), .CO(C[655]) );
  FA_11945 \FA_INST_0[1].FA_INST_1[143].FA_  ( .A(A[655]), .B(n1680), .CI(
        C[655]), .S(S[655]), .CO(C[656]) );
  FA_11944 \FA_INST_0[1].FA_INST_1[144].FA_  ( .A(A[656]), .B(n1681), .CI(
        C[656]), .S(S[656]), .CO(C[657]) );
  FA_11943 \FA_INST_0[1].FA_INST_1[145].FA_  ( .A(A[657]), .B(n1682), .CI(
        C[657]), .S(S[657]), .CO(C[658]) );
  FA_11942 \FA_INST_0[1].FA_INST_1[146].FA_  ( .A(A[658]), .B(n1683), .CI(
        C[658]), .S(S[658]), .CO(C[659]) );
  FA_11941 \FA_INST_0[1].FA_INST_1[147].FA_  ( .A(A[659]), .B(n1684), .CI(
        C[659]), .S(S[659]), .CO(C[660]) );
  FA_11940 \FA_INST_0[1].FA_INST_1[148].FA_  ( .A(A[660]), .B(n1685), .CI(
        C[660]), .S(S[660]), .CO(C[661]) );
  FA_11939 \FA_INST_0[1].FA_INST_1[149].FA_  ( .A(A[661]), .B(n1686), .CI(
        C[661]), .S(S[661]), .CO(C[662]) );
  FA_11938 \FA_INST_0[1].FA_INST_1[150].FA_  ( .A(A[662]), .B(n1687), .CI(
        C[662]), .S(S[662]), .CO(C[663]) );
  FA_11937 \FA_INST_0[1].FA_INST_1[151].FA_  ( .A(A[663]), .B(n1688), .CI(
        C[663]), .S(S[663]), .CO(C[664]) );
  FA_11936 \FA_INST_0[1].FA_INST_1[152].FA_  ( .A(A[664]), .B(n1689), .CI(
        C[664]), .S(S[664]), .CO(C[665]) );
  FA_11935 \FA_INST_0[1].FA_INST_1[153].FA_  ( .A(A[665]), .B(n1690), .CI(
        C[665]), .S(S[665]), .CO(C[666]) );
  FA_11934 \FA_INST_0[1].FA_INST_1[154].FA_  ( .A(A[666]), .B(n1691), .CI(
        C[666]), .S(S[666]), .CO(C[667]) );
  FA_11933 \FA_INST_0[1].FA_INST_1[155].FA_  ( .A(A[667]), .B(n1692), .CI(
        C[667]), .S(S[667]), .CO(C[668]) );
  FA_11932 \FA_INST_0[1].FA_INST_1[156].FA_  ( .A(A[668]), .B(n1693), .CI(
        C[668]), .S(S[668]), .CO(C[669]) );
  FA_11931 \FA_INST_0[1].FA_INST_1[157].FA_  ( .A(A[669]), .B(n1694), .CI(
        C[669]), .S(S[669]), .CO(C[670]) );
  FA_11930 \FA_INST_0[1].FA_INST_1[158].FA_  ( .A(A[670]), .B(n1695), .CI(
        C[670]), .S(S[670]), .CO(C[671]) );
  FA_11929 \FA_INST_0[1].FA_INST_1[159].FA_  ( .A(A[671]), .B(n1696), .CI(
        C[671]), .S(S[671]), .CO(C[672]) );
  FA_11928 \FA_INST_0[1].FA_INST_1[160].FA_  ( .A(A[672]), .B(n1697), .CI(
        C[672]), .S(S[672]), .CO(C[673]) );
  FA_11927 \FA_INST_0[1].FA_INST_1[161].FA_  ( .A(A[673]), .B(n1698), .CI(
        C[673]), .S(S[673]), .CO(C[674]) );
  FA_11926 \FA_INST_0[1].FA_INST_1[162].FA_  ( .A(A[674]), .B(n1699), .CI(
        C[674]), .S(S[674]), .CO(C[675]) );
  FA_11925 \FA_INST_0[1].FA_INST_1[163].FA_  ( .A(A[675]), .B(n1700), .CI(
        C[675]), .S(S[675]), .CO(C[676]) );
  FA_11924 \FA_INST_0[1].FA_INST_1[164].FA_  ( .A(A[676]), .B(n1701), .CI(
        C[676]), .S(S[676]), .CO(C[677]) );
  FA_11923 \FA_INST_0[1].FA_INST_1[165].FA_  ( .A(A[677]), .B(n1702), .CI(
        C[677]), .S(S[677]), .CO(C[678]) );
  FA_11922 \FA_INST_0[1].FA_INST_1[166].FA_  ( .A(A[678]), .B(n1703), .CI(
        C[678]), .S(S[678]), .CO(C[679]) );
  FA_11921 \FA_INST_0[1].FA_INST_1[167].FA_  ( .A(A[679]), .B(n1704), .CI(
        C[679]), .S(S[679]), .CO(C[680]) );
  FA_11920 \FA_INST_0[1].FA_INST_1[168].FA_  ( .A(A[680]), .B(n1705), .CI(
        C[680]), .S(S[680]), .CO(C[681]) );
  FA_11919 \FA_INST_0[1].FA_INST_1[169].FA_  ( .A(A[681]), .B(n1706), .CI(
        C[681]), .S(S[681]), .CO(C[682]) );
  FA_11918 \FA_INST_0[1].FA_INST_1[170].FA_  ( .A(A[682]), .B(n1707), .CI(
        C[682]), .S(S[682]), .CO(C[683]) );
  FA_11917 \FA_INST_0[1].FA_INST_1[171].FA_  ( .A(A[683]), .B(n1708), .CI(
        C[683]), .S(S[683]), .CO(C[684]) );
  FA_11916 \FA_INST_0[1].FA_INST_1[172].FA_  ( .A(A[684]), .B(n1709), .CI(
        C[684]), .S(S[684]), .CO(C[685]) );
  FA_11915 \FA_INST_0[1].FA_INST_1[173].FA_  ( .A(A[685]), .B(n1710), .CI(
        C[685]), .S(S[685]), .CO(C[686]) );
  FA_11914 \FA_INST_0[1].FA_INST_1[174].FA_  ( .A(A[686]), .B(n1711), .CI(
        C[686]), .S(S[686]), .CO(C[687]) );
  FA_11913 \FA_INST_0[1].FA_INST_1[175].FA_  ( .A(A[687]), .B(n1712), .CI(
        C[687]), .S(S[687]), .CO(C[688]) );
  FA_11912 \FA_INST_0[1].FA_INST_1[176].FA_  ( .A(A[688]), .B(n1713), .CI(
        C[688]), .S(S[688]), .CO(C[689]) );
  FA_11911 \FA_INST_0[1].FA_INST_1[177].FA_  ( .A(A[689]), .B(n1714), .CI(
        C[689]), .S(S[689]), .CO(C[690]) );
  FA_11910 \FA_INST_0[1].FA_INST_1[178].FA_  ( .A(A[690]), .B(n1715), .CI(
        C[690]), .S(S[690]), .CO(C[691]) );
  FA_11909 \FA_INST_0[1].FA_INST_1[179].FA_  ( .A(A[691]), .B(n1716), .CI(
        C[691]), .S(S[691]), .CO(C[692]) );
  FA_11908 \FA_INST_0[1].FA_INST_1[180].FA_  ( .A(A[692]), .B(n1717), .CI(
        C[692]), .S(S[692]), .CO(C[693]) );
  FA_11907 \FA_INST_0[1].FA_INST_1[181].FA_  ( .A(A[693]), .B(n1718), .CI(
        C[693]), .S(S[693]), .CO(C[694]) );
  FA_11906 \FA_INST_0[1].FA_INST_1[182].FA_  ( .A(A[694]), .B(n1719), .CI(
        C[694]), .S(S[694]), .CO(C[695]) );
  FA_11905 \FA_INST_0[1].FA_INST_1[183].FA_  ( .A(A[695]), .B(n1720), .CI(
        C[695]), .S(S[695]), .CO(C[696]) );
  FA_11904 \FA_INST_0[1].FA_INST_1[184].FA_  ( .A(A[696]), .B(n1721), .CI(
        C[696]), .S(S[696]), .CO(C[697]) );
  FA_11903 \FA_INST_0[1].FA_INST_1[185].FA_  ( .A(A[697]), .B(n1722), .CI(
        C[697]), .S(S[697]), .CO(C[698]) );
  FA_11902 \FA_INST_0[1].FA_INST_1[186].FA_  ( .A(A[698]), .B(n1723), .CI(
        C[698]), .S(S[698]), .CO(C[699]) );
  FA_11901 \FA_INST_0[1].FA_INST_1[187].FA_  ( .A(A[699]), .B(n1724), .CI(
        C[699]), .S(S[699]), .CO(C[700]) );
  FA_11900 \FA_INST_0[1].FA_INST_1[188].FA_  ( .A(A[700]), .B(n1725), .CI(
        C[700]), .S(S[700]), .CO(C[701]) );
  FA_11899 \FA_INST_0[1].FA_INST_1[189].FA_  ( .A(A[701]), .B(n1726), .CI(
        C[701]), .S(S[701]), .CO(C[702]) );
  FA_11898 \FA_INST_0[1].FA_INST_1[190].FA_  ( .A(A[702]), .B(n1727), .CI(
        C[702]), .S(S[702]), .CO(C[703]) );
  FA_11897 \FA_INST_0[1].FA_INST_1[191].FA_  ( .A(A[703]), .B(n1728), .CI(
        C[703]), .S(S[703]), .CO(C[704]) );
  FA_11896 \FA_INST_0[1].FA_INST_1[192].FA_  ( .A(A[704]), .B(n1729), .CI(
        C[704]), .S(S[704]), .CO(C[705]) );
  FA_11895 \FA_INST_0[1].FA_INST_1[193].FA_  ( .A(A[705]), .B(n1730), .CI(
        C[705]), .S(S[705]), .CO(C[706]) );
  FA_11894 \FA_INST_0[1].FA_INST_1[194].FA_  ( .A(A[706]), .B(n1731), .CI(
        C[706]), .S(S[706]), .CO(C[707]) );
  FA_11893 \FA_INST_0[1].FA_INST_1[195].FA_  ( .A(A[707]), .B(n1732), .CI(
        C[707]), .S(S[707]), .CO(C[708]) );
  FA_11892 \FA_INST_0[1].FA_INST_1[196].FA_  ( .A(A[708]), .B(n1733), .CI(
        C[708]), .S(S[708]), .CO(C[709]) );
  FA_11891 \FA_INST_0[1].FA_INST_1[197].FA_  ( .A(A[709]), .B(n1734), .CI(
        C[709]), .S(S[709]), .CO(C[710]) );
  FA_11890 \FA_INST_0[1].FA_INST_1[198].FA_  ( .A(A[710]), .B(n1735), .CI(
        C[710]), .S(S[710]), .CO(C[711]) );
  FA_11889 \FA_INST_0[1].FA_INST_1[199].FA_  ( .A(A[711]), .B(n1736), .CI(
        C[711]), .S(S[711]), .CO(C[712]) );
  FA_11888 \FA_INST_0[1].FA_INST_1[200].FA_  ( .A(A[712]), .B(n1737), .CI(
        C[712]), .S(S[712]), .CO(C[713]) );
  FA_11887 \FA_INST_0[1].FA_INST_1[201].FA_  ( .A(A[713]), .B(n1738), .CI(
        C[713]), .S(S[713]), .CO(C[714]) );
  FA_11886 \FA_INST_0[1].FA_INST_1[202].FA_  ( .A(A[714]), .B(n1739), .CI(
        C[714]), .S(S[714]), .CO(C[715]) );
  FA_11885 \FA_INST_0[1].FA_INST_1[203].FA_  ( .A(A[715]), .B(n1740), .CI(
        C[715]), .S(S[715]), .CO(C[716]) );
  FA_11884 \FA_INST_0[1].FA_INST_1[204].FA_  ( .A(A[716]), .B(n1741), .CI(
        C[716]), .S(S[716]), .CO(C[717]) );
  FA_11883 \FA_INST_0[1].FA_INST_1[205].FA_  ( .A(A[717]), .B(n1742), .CI(
        C[717]), .S(S[717]), .CO(C[718]) );
  FA_11882 \FA_INST_0[1].FA_INST_1[206].FA_  ( .A(A[718]), .B(n1743), .CI(
        C[718]), .S(S[718]), .CO(C[719]) );
  FA_11881 \FA_INST_0[1].FA_INST_1[207].FA_  ( .A(A[719]), .B(n1744), .CI(
        C[719]), .S(S[719]), .CO(C[720]) );
  FA_11880 \FA_INST_0[1].FA_INST_1[208].FA_  ( .A(A[720]), .B(n1745), .CI(
        C[720]), .S(S[720]), .CO(C[721]) );
  FA_11879 \FA_INST_0[1].FA_INST_1[209].FA_  ( .A(A[721]), .B(n1746), .CI(
        C[721]), .S(S[721]), .CO(C[722]) );
  FA_11878 \FA_INST_0[1].FA_INST_1[210].FA_  ( .A(A[722]), .B(n1747), .CI(
        C[722]), .S(S[722]), .CO(C[723]) );
  FA_11877 \FA_INST_0[1].FA_INST_1[211].FA_  ( .A(A[723]), .B(n1748), .CI(
        C[723]), .S(S[723]), .CO(C[724]) );
  FA_11876 \FA_INST_0[1].FA_INST_1[212].FA_  ( .A(A[724]), .B(n1749), .CI(
        C[724]), .S(S[724]), .CO(C[725]) );
  FA_11875 \FA_INST_0[1].FA_INST_1[213].FA_  ( .A(A[725]), .B(n1750), .CI(
        C[725]), .S(S[725]), .CO(C[726]) );
  FA_11874 \FA_INST_0[1].FA_INST_1[214].FA_  ( .A(A[726]), .B(n1751), .CI(
        C[726]), .S(S[726]), .CO(C[727]) );
  FA_11873 \FA_INST_0[1].FA_INST_1[215].FA_  ( .A(A[727]), .B(n1752), .CI(
        C[727]), .S(S[727]), .CO(C[728]) );
  FA_11872 \FA_INST_0[1].FA_INST_1[216].FA_  ( .A(A[728]), .B(n1753), .CI(
        C[728]), .S(S[728]), .CO(C[729]) );
  FA_11871 \FA_INST_0[1].FA_INST_1[217].FA_  ( .A(A[729]), .B(n1754), .CI(
        C[729]), .S(S[729]), .CO(C[730]) );
  FA_11870 \FA_INST_0[1].FA_INST_1[218].FA_  ( .A(A[730]), .B(n1755), .CI(
        C[730]), .S(S[730]), .CO(C[731]) );
  FA_11869 \FA_INST_0[1].FA_INST_1[219].FA_  ( .A(A[731]), .B(n1756), .CI(
        C[731]), .S(S[731]), .CO(C[732]) );
  FA_11868 \FA_INST_0[1].FA_INST_1[220].FA_  ( .A(A[732]), .B(n1757), .CI(
        C[732]), .S(S[732]), .CO(C[733]) );
  FA_11867 \FA_INST_0[1].FA_INST_1[221].FA_  ( .A(A[733]), .B(n1758), .CI(
        C[733]), .S(S[733]), .CO(C[734]) );
  FA_11866 \FA_INST_0[1].FA_INST_1[222].FA_  ( .A(A[734]), .B(n1759), .CI(
        C[734]), .S(S[734]), .CO(C[735]) );
  FA_11865 \FA_INST_0[1].FA_INST_1[223].FA_  ( .A(A[735]), .B(n1760), .CI(
        C[735]), .S(S[735]), .CO(C[736]) );
  FA_11864 \FA_INST_0[1].FA_INST_1[224].FA_  ( .A(A[736]), .B(n1761), .CI(
        C[736]), .S(S[736]), .CO(C[737]) );
  FA_11863 \FA_INST_0[1].FA_INST_1[225].FA_  ( .A(A[737]), .B(n1762), .CI(
        C[737]), .S(S[737]), .CO(C[738]) );
  FA_11862 \FA_INST_0[1].FA_INST_1[226].FA_  ( .A(A[738]), .B(n1763), .CI(
        C[738]), .S(S[738]), .CO(C[739]) );
  FA_11861 \FA_INST_0[1].FA_INST_1[227].FA_  ( .A(A[739]), .B(n1764), .CI(
        C[739]), .S(S[739]), .CO(C[740]) );
  FA_11860 \FA_INST_0[1].FA_INST_1[228].FA_  ( .A(A[740]), .B(n1765), .CI(
        C[740]), .S(S[740]), .CO(C[741]) );
  FA_11859 \FA_INST_0[1].FA_INST_1[229].FA_  ( .A(A[741]), .B(n1766), .CI(
        C[741]), .S(S[741]), .CO(C[742]) );
  FA_11858 \FA_INST_0[1].FA_INST_1[230].FA_  ( .A(A[742]), .B(n1767), .CI(
        C[742]), .S(S[742]), .CO(C[743]) );
  FA_11857 \FA_INST_0[1].FA_INST_1[231].FA_  ( .A(A[743]), .B(n1768), .CI(
        C[743]), .S(S[743]), .CO(C[744]) );
  FA_11856 \FA_INST_0[1].FA_INST_1[232].FA_  ( .A(A[744]), .B(n1769), .CI(
        C[744]), .S(S[744]), .CO(C[745]) );
  FA_11855 \FA_INST_0[1].FA_INST_1[233].FA_  ( .A(A[745]), .B(n1770), .CI(
        C[745]), .S(S[745]), .CO(C[746]) );
  FA_11854 \FA_INST_0[1].FA_INST_1[234].FA_  ( .A(A[746]), .B(n1771), .CI(
        C[746]), .S(S[746]), .CO(C[747]) );
  FA_11853 \FA_INST_0[1].FA_INST_1[235].FA_  ( .A(A[747]), .B(n1772), .CI(
        C[747]), .S(S[747]), .CO(C[748]) );
  FA_11852 \FA_INST_0[1].FA_INST_1[236].FA_  ( .A(A[748]), .B(n1773), .CI(
        C[748]), .S(S[748]), .CO(C[749]) );
  FA_11851 \FA_INST_0[1].FA_INST_1[237].FA_  ( .A(A[749]), .B(n1774), .CI(
        C[749]), .S(S[749]), .CO(C[750]) );
  FA_11850 \FA_INST_0[1].FA_INST_1[238].FA_  ( .A(A[750]), .B(n1775), .CI(
        C[750]), .S(S[750]), .CO(C[751]) );
  FA_11849 \FA_INST_0[1].FA_INST_1[239].FA_  ( .A(A[751]), .B(n1776), .CI(
        C[751]), .S(S[751]), .CO(C[752]) );
  FA_11848 \FA_INST_0[1].FA_INST_1[240].FA_  ( .A(A[752]), .B(n1777), .CI(
        C[752]), .S(S[752]), .CO(C[753]) );
  FA_11847 \FA_INST_0[1].FA_INST_1[241].FA_  ( .A(A[753]), .B(n1778), .CI(
        C[753]), .S(S[753]), .CO(C[754]) );
  FA_11846 \FA_INST_0[1].FA_INST_1[242].FA_  ( .A(A[754]), .B(n1779), .CI(
        C[754]), .S(S[754]), .CO(C[755]) );
  FA_11845 \FA_INST_0[1].FA_INST_1[243].FA_  ( .A(A[755]), .B(n1780), .CI(
        C[755]), .S(S[755]), .CO(C[756]) );
  FA_11844 \FA_INST_0[1].FA_INST_1[244].FA_  ( .A(A[756]), .B(n1781), .CI(
        C[756]), .S(S[756]), .CO(C[757]) );
  FA_11843 \FA_INST_0[1].FA_INST_1[245].FA_  ( .A(A[757]), .B(n1782), .CI(
        C[757]), .S(S[757]), .CO(C[758]) );
  FA_11842 \FA_INST_0[1].FA_INST_1[246].FA_  ( .A(A[758]), .B(n1783), .CI(
        C[758]), .S(S[758]), .CO(C[759]) );
  FA_11841 \FA_INST_0[1].FA_INST_1[247].FA_  ( .A(A[759]), .B(n1784), .CI(
        C[759]), .S(S[759]), .CO(C[760]) );
  FA_11840 \FA_INST_0[1].FA_INST_1[248].FA_  ( .A(A[760]), .B(n1785), .CI(
        C[760]), .S(S[760]), .CO(C[761]) );
  FA_11839 \FA_INST_0[1].FA_INST_1[249].FA_  ( .A(A[761]), .B(n1786), .CI(
        C[761]), .S(S[761]), .CO(C[762]) );
  FA_11838 \FA_INST_0[1].FA_INST_1[250].FA_  ( .A(A[762]), .B(n1787), .CI(
        C[762]), .S(S[762]), .CO(C[763]) );
  FA_11837 \FA_INST_0[1].FA_INST_1[251].FA_  ( .A(A[763]), .B(n1788), .CI(
        C[763]), .S(S[763]), .CO(C[764]) );
  FA_11836 \FA_INST_0[1].FA_INST_1[252].FA_  ( .A(A[764]), .B(n1789), .CI(
        C[764]), .S(S[764]), .CO(C[765]) );
  FA_11835 \FA_INST_0[1].FA_INST_1[253].FA_  ( .A(A[765]), .B(n1790), .CI(
        C[765]), .S(S[765]), .CO(C[766]) );
  FA_11834 \FA_INST_0[1].FA_INST_1[254].FA_  ( .A(A[766]), .B(n1791), .CI(
        C[766]), .S(S[766]), .CO(C[767]) );
  FA_11833 \FA_INST_0[1].FA_INST_1[255].FA_  ( .A(A[767]), .B(n1792), .CI(
        C[767]), .S(S[767]), .CO(C[768]) );
  FA_11832 \FA_INST_0[1].FA_INST_1[256].FA_  ( .A(A[768]), .B(n1793), .CI(
        C[768]), .S(S[768]), .CO(C[769]) );
  FA_11831 \FA_INST_0[1].FA_INST_1[257].FA_  ( .A(A[769]), .B(n1794), .CI(
        C[769]), .S(S[769]), .CO(C[770]) );
  FA_11830 \FA_INST_0[1].FA_INST_1[258].FA_  ( .A(A[770]), .B(n1795), .CI(
        C[770]), .S(S[770]), .CO(C[771]) );
  FA_11829 \FA_INST_0[1].FA_INST_1[259].FA_  ( .A(A[771]), .B(n1796), .CI(
        C[771]), .S(S[771]), .CO(C[772]) );
  FA_11828 \FA_INST_0[1].FA_INST_1[260].FA_  ( .A(A[772]), .B(n1797), .CI(
        C[772]), .S(S[772]), .CO(C[773]) );
  FA_11827 \FA_INST_0[1].FA_INST_1[261].FA_  ( .A(A[773]), .B(n1798), .CI(
        C[773]), .S(S[773]), .CO(C[774]) );
  FA_11826 \FA_INST_0[1].FA_INST_1[262].FA_  ( .A(A[774]), .B(n1799), .CI(
        C[774]), .S(S[774]), .CO(C[775]) );
  FA_11825 \FA_INST_0[1].FA_INST_1[263].FA_  ( .A(A[775]), .B(n1800), .CI(
        C[775]), .S(S[775]), .CO(C[776]) );
  FA_11824 \FA_INST_0[1].FA_INST_1[264].FA_  ( .A(A[776]), .B(n1801), .CI(
        C[776]), .S(S[776]), .CO(C[777]) );
  FA_11823 \FA_INST_0[1].FA_INST_1[265].FA_  ( .A(A[777]), .B(n1802), .CI(
        C[777]), .S(S[777]), .CO(C[778]) );
  FA_11822 \FA_INST_0[1].FA_INST_1[266].FA_  ( .A(A[778]), .B(n1803), .CI(
        C[778]), .S(S[778]), .CO(C[779]) );
  FA_11821 \FA_INST_0[1].FA_INST_1[267].FA_  ( .A(A[779]), .B(n1804), .CI(
        C[779]), .S(S[779]), .CO(C[780]) );
  FA_11820 \FA_INST_0[1].FA_INST_1[268].FA_  ( .A(A[780]), .B(n1805), .CI(
        C[780]), .S(S[780]), .CO(C[781]) );
  FA_11819 \FA_INST_0[1].FA_INST_1[269].FA_  ( .A(A[781]), .B(n1806), .CI(
        C[781]), .S(S[781]), .CO(C[782]) );
  FA_11818 \FA_INST_0[1].FA_INST_1[270].FA_  ( .A(A[782]), .B(n1807), .CI(
        C[782]), .S(S[782]), .CO(C[783]) );
  FA_11817 \FA_INST_0[1].FA_INST_1[271].FA_  ( .A(A[783]), .B(n1808), .CI(
        C[783]), .S(S[783]), .CO(C[784]) );
  FA_11816 \FA_INST_0[1].FA_INST_1[272].FA_  ( .A(A[784]), .B(n1809), .CI(
        C[784]), .S(S[784]), .CO(C[785]) );
  FA_11815 \FA_INST_0[1].FA_INST_1[273].FA_  ( .A(A[785]), .B(n1810), .CI(
        C[785]), .S(S[785]), .CO(C[786]) );
  FA_11814 \FA_INST_0[1].FA_INST_1[274].FA_  ( .A(A[786]), .B(n1811), .CI(
        C[786]), .S(S[786]), .CO(C[787]) );
  FA_11813 \FA_INST_0[1].FA_INST_1[275].FA_  ( .A(A[787]), .B(n1812), .CI(
        C[787]), .S(S[787]), .CO(C[788]) );
  FA_11812 \FA_INST_0[1].FA_INST_1[276].FA_  ( .A(A[788]), .B(n1813), .CI(
        C[788]), .S(S[788]), .CO(C[789]) );
  FA_11811 \FA_INST_0[1].FA_INST_1[277].FA_  ( .A(A[789]), .B(n1814), .CI(
        C[789]), .S(S[789]), .CO(C[790]) );
  FA_11810 \FA_INST_0[1].FA_INST_1[278].FA_  ( .A(A[790]), .B(n1815), .CI(
        C[790]), .S(S[790]), .CO(C[791]) );
  FA_11809 \FA_INST_0[1].FA_INST_1[279].FA_  ( .A(A[791]), .B(n1816), .CI(
        C[791]), .S(S[791]), .CO(C[792]) );
  FA_11808 \FA_INST_0[1].FA_INST_1[280].FA_  ( .A(A[792]), .B(n1817), .CI(
        C[792]), .S(S[792]), .CO(C[793]) );
  FA_11807 \FA_INST_0[1].FA_INST_1[281].FA_  ( .A(A[793]), .B(n1818), .CI(
        C[793]), .S(S[793]), .CO(C[794]) );
  FA_11806 \FA_INST_0[1].FA_INST_1[282].FA_  ( .A(A[794]), .B(n1819), .CI(
        C[794]), .S(S[794]), .CO(C[795]) );
  FA_11805 \FA_INST_0[1].FA_INST_1[283].FA_  ( .A(A[795]), .B(n1820), .CI(
        C[795]), .S(S[795]), .CO(C[796]) );
  FA_11804 \FA_INST_0[1].FA_INST_1[284].FA_  ( .A(A[796]), .B(n1821), .CI(
        C[796]), .S(S[796]), .CO(C[797]) );
  FA_11803 \FA_INST_0[1].FA_INST_1[285].FA_  ( .A(A[797]), .B(n1822), .CI(
        C[797]), .S(S[797]), .CO(C[798]) );
  FA_11802 \FA_INST_0[1].FA_INST_1[286].FA_  ( .A(A[798]), .B(n1823), .CI(
        C[798]), .S(S[798]), .CO(C[799]) );
  FA_11801 \FA_INST_0[1].FA_INST_1[287].FA_  ( .A(A[799]), .B(n1824), .CI(
        C[799]), .S(S[799]), .CO(C[800]) );
  FA_11800 \FA_INST_0[1].FA_INST_1[288].FA_  ( .A(A[800]), .B(n1825), .CI(
        C[800]), .S(S[800]), .CO(C[801]) );
  FA_11799 \FA_INST_0[1].FA_INST_1[289].FA_  ( .A(A[801]), .B(n1826), .CI(
        C[801]), .S(S[801]), .CO(C[802]) );
  FA_11798 \FA_INST_0[1].FA_INST_1[290].FA_  ( .A(A[802]), .B(n1827), .CI(
        C[802]), .S(S[802]), .CO(C[803]) );
  FA_11797 \FA_INST_0[1].FA_INST_1[291].FA_  ( .A(A[803]), .B(n1828), .CI(
        C[803]), .S(S[803]), .CO(C[804]) );
  FA_11796 \FA_INST_0[1].FA_INST_1[292].FA_  ( .A(A[804]), .B(n1829), .CI(
        C[804]), .S(S[804]), .CO(C[805]) );
  FA_11795 \FA_INST_0[1].FA_INST_1[293].FA_  ( .A(A[805]), .B(n1830), .CI(
        C[805]), .S(S[805]), .CO(C[806]) );
  FA_11794 \FA_INST_0[1].FA_INST_1[294].FA_  ( .A(A[806]), .B(n1831), .CI(
        C[806]), .S(S[806]), .CO(C[807]) );
  FA_11793 \FA_INST_0[1].FA_INST_1[295].FA_  ( .A(A[807]), .B(n1832), .CI(
        C[807]), .S(S[807]), .CO(C[808]) );
  FA_11792 \FA_INST_0[1].FA_INST_1[296].FA_  ( .A(A[808]), .B(n1833), .CI(
        C[808]), .S(S[808]), .CO(C[809]) );
  FA_11791 \FA_INST_0[1].FA_INST_1[297].FA_  ( .A(A[809]), .B(n1834), .CI(
        C[809]), .S(S[809]), .CO(C[810]) );
  FA_11790 \FA_INST_0[1].FA_INST_1[298].FA_  ( .A(A[810]), .B(n1835), .CI(
        C[810]), .S(S[810]), .CO(C[811]) );
  FA_11789 \FA_INST_0[1].FA_INST_1[299].FA_  ( .A(A[811]), .B(n1836), .CI(
        C[811]), .S(S[811]), .CO(C[812]) );
  FA_11788 \FA_INST_0[1].FA_INST_1[300].FA_  ( .A(A[812]), .B(n1837), .CI(
        C[812]), .S(S[812]), .CO(C[813]) );
  FA_11787 \FA_INST_0[1].FA_INST_1[301].FA_  ( .A(A[813]), .B(n1838), .CI(
        C[813]), .S(S[813]), .CO(C[814]) );
  FA_11786 \FA_INST_0[1].FA_INST_1[302].FA_  ( .A(A[814]), .B(n1839), .CI(
        C[814]), .S(S[814]), .CO(C[815]) );
  FA_11785 \FA_INST_0[1].FA_INST_1[303].FA_  ( .A(A[815]), .B(n1840), .CI(
        C[815]), .S(S[815]), .CO(C[816]) );
  FA_11784 \FA_INST_0[1].FA_INST_1[304].FA_  ( .A(A[816]), .B(n1841), .CI(
        C[816]), .S(S[816]), .CO(C[817]) );
  FA_11783 \FA_INST_0[1].FA_INST_1[305].FA_  ( .A(A[817]), .B(n1842), .CI(
        C[817]), .S(S[817]), .CO(C[818]) );
  FA_11782 \FA_INST_0[1].FA_INST_1[306].FA_  ( .A(A[818]), .B(n1843), .CI(
        C[818]), .S(S[818]), .CO(C[819]) );
  FA_11781 \FA_INST_0[1].FA_INST_1[307].FA_  ( .A(A[819]), .B(n1844), .CI(
        C[819]), .S(S[819]), .CO(C[820]) );
  FA_11780 \FA_INST_0[1].FA_INST_1[308].FA_  ( .A(A[820]), .B(n1845), .CI(
        C[820]), .S(S[820]), .CO(C[821]) );
  FA_11779 \FA_INST_0[1].FA_INST_1[309].FA_  ( .A(A[821]), .B(n1846), .CI(
        C[821]), .S(S[821]), .CO(C[822]) );
  FA_11778 \FA_INST_0[1].FA_INST_1[310].FA_  ( .A(A[822]), .B(n1847), .CI(
        C[822]), .S(S[822]), .CO(C[823]) );
  FA_11777 \FA_INST_0[1].FA_INST_1[311].FA_  ( .A(A[823]), .B(n1848), .CI(
        C[823]), .S(S[823]), .CO(C[824]) );
  FA_11776 \FA_INST_0[1].FA_INST_1[312].FA_  ( .A(A[824]), .B(n1849), .CI(
        C[824]), .S(S[824]), .CO(C[825]) );
  FA_11775 \FA_INST_0[1].FA_INST_1[313].FA_  ( .A(A[825]), .B(n1850), .CI(
        C[825]), .S(S[825]), .CO(C[826]) );
  FA_11774 \FA_INST_0[1].FA_INST_1[314].FA_  ( .A(A[826]), .B(n1851), .CI(
        C[826]), .S(S[826]), .CO(C[827]) );
  FA_11773 \FA_INST_0[1].FA_INST_1[315].FA_  ( .A(A[827]), .B(n1852), .CI(
        C[827]), .S(S[827]), .CO(C[828]) );
  FA_11772 \FA_INST_0[1].FA_INST_1[316].FA_  ( .A(A[828]), .B(n1853), .CI(
        C[828]), .S(S[828]), .CO(C[829]) );
  FA_11771 \FA_INST_0[1].FA_INST_1[317].FA_  ( .A(A[829]), .B(n1854), .CI(
        C[829]), .S(S[829]), .CO(C[830]) );
  FA_11770 \FA_INST_0[1].FA_INST_1[318].FA_  ( .A(A[830]), .B(n1855), .CI(
        C[830]), .S(S[830]), .CO(C[831]) );
  FA_11769 \FA_INST_0[1].FA_INST_1[319].FA_  ( .A(A[831]), .B(n1856), .CI(
        C[831]), .S(S[831]), .CO(C[832]) );
  FA_11768 \FA_INST_0[1].FA_INST_1[320].FA_  ( .A(A[832]), .B(n1857), .CI(
        C[832]), .S(S[832]), .CO(C[833]) );
  FA_11767 \FA_INST_0[1].FA_INST_1[321].FA_  ( .A(A[833]), .B(n1858), .CI(
        C[833]), .S(S[833]), .CO(C[834]) );
  FA_11766 \FA_INST_0[1].FA_INST_1[322].FA_  ( .A(A[834]), .B(n1859), .CI(
        C[834]), .S(S[834]), .CO(C[835]) );
  FA_11765 \FA_INST_0[1].FA_INST_1[323].FA_  ( .A(A[835]), .B(n1860), .CI(
        C[835]), .S(S[835]), .CO(C[836]) );
  FA_11764 \FA_INST_0[1].FA_INST_1[324].FA_  ( .A(A[836]), .B(n1861), .CI(
        C[836]), .S(S[836]), .CO(C[837]) );
  FA_11763 \FA_INST_0[1].FA_INST_1[325].FA_  ( .A(A[837]), .B(n1862), .CI(
        C[837]), .S(S[837]), .CO(C[838]) );
  FA_11762 \FA_INST_0[1].FA_INST_1[326].FA_  ( .A(A[838]), .B(n1863), .CI(
        C[838]), .S(S[838]), .CO(C[839]) );
  FA_11761 \FA_INST_0[1].FA_INST_1[327].FA_  ( .A(A[839]), .B(n1864), .CI(
        C[839]), .S(S[839]), .CO(C[840]) );
  FA_11760 \FA_INST_0[1].FA_INST_1[328].FA_  ( .A(A[840]), .B(n1865), .CI(
        C[840]), .S(S[840]), .CO(C[841]) );
  FA_11759 \FA_INST_0[1].FA_INST_1[329].FA_  ( .A(A[841]), .B(n1866), .CI(
        C[841]), .S(S[841]), .CO(C[842]) );
  FA_11758 \FA_INST_0[1].FA_INST_1[330].FA_  ( .A(A[842]), .B(n1867), .CI(
        C[842]), .S(S[842]), .CO(C[843]) );
  FA_11757 \FA_INST_0[1].FA_INST_1[331].FA_  ( .A(A[843]), .B(n1868), .CI(
        C[843]), .S(S[843]), .CO(C[844]) );
  FA_11756 \FA_INST_0[1].FA_INST_1[332].FA_  ( .A(A[844]), .B(n1869), .CI(
        C[844]), .S(S[844]), .CO(C[845]) );
  FA_11755 \FA_INST_0[1].FA_INST_1[333].FA_  ( .A(A[845]), .B(n1870), .CI(
        C[845]), .S(S[845]), .CO(C[846]) );
  FA_11754 \FA_INST_0[1].FA_INST_1[334].FA_  ( .A(A[846]), .B(n1871), .CI(
        C[846]), .S(S[846]), .CO(C[847]) );
  FA_11753 \FA_INST_0[1].FA_INST_1[335].FA_  ( .A(A[847]), .B(n1872), .CI(
        C[847]), .S(S[847]), .CO(C[848]) );
  FA_11752 \FA_INST_0[1].FA_INST_1[336].FA_  ( .A(A[848]), .B(n1873), .CI(
        C[848]), .S(S[848]), .CO(C[849]) );
  FA_11751 \FA_INST_0[1].FA_INST_1[337].FA_  ( .A(A[849]), .B(n1874), .CI(
        C[849]), .S(S[849]), .CO(C[850]) );
  FA_11750 \FA_INST_0[1].FA_INST_1[338].FA_  ( .A(A[850]), .B(n1875), .CI(
        C[850]), .S(S[850]), .CO(C[851]) );
  FA_11749 \FA_INST_0[1].FA_INST_1[339].FA_  ( .A(A[851]), .B(n1876), .CI(
        C[851]), .S(S[851]), .CO(C[852]) );
  FA_11748 \FA_INST_0[1].FA_INST_1[340].FA_  ( .A(A[852]), .B(n1877), .CI(
        C[852]), .S(S[852]), .CO(C[853]) );
  FA_11747 \FA_INST_0[1].FA_INST_1[341].FA_  ( .A(A[853]), .B(n1878), .CI(
        C[853]), .S(S[853]), .CO(C[854]) );
  FA_11746 \FA_INST_0[1].FA_INST_1[342].FA_  ( .A(A[854]), .B(n1879), .CI(
        C[854]), .S(S[854]), .CO(C[855]) );
  FA_11745 \FA_INST_0[1].FA_INST_1[343].FA_  ( .A(A[855]), .B(n1880), .CI(
        C[855]), .S(S[855]), .CO(C[856]) );
  FA_11744 \FA_INST_0[1].FA_INST_1[344].FA_  ( .A(A[856]), .B(n1881), .CI(
        C[856]), .S(S[856]), .CO(C[857]) );
  FA_11743 \FA_INST_0[1].FA_INST_1[345].FA_  ( .A(A[857]), .B(n1882), .CI(
        C[857]), .S(S[857]), .CO(C[858]) );
  FA_11742 \FA_INST_0[1].FA_INST_1[346].FA_  ( .A(A[858]), .B(n1883), .CI(
        C[858]), .S(S[858]), .CO(C[859]) );
  FA_11741 \FA_INST_0[1].FA_INST_1[347].FA_  ( .A(A[859]), .B(n1884), .CI(
        C[859]), .S(S[859]), .CO(C[860]) );
  FA_11740 \FA_INST_0[1].FA_INST_1[348].FA_  ( .A(A[860]), .B(n1885), .CI(
        C[860]), .S(S[860]), .CO(C[861]) );
  FA_11739 \FA_INST_0[1].FA_INST_1[349].FA_  ( .A(A[861]), .B(n1886), .CI(
        C[861]), .S(S[861]), .CO(C[862]) );
  FA_11738 \FA_INST_0[1].FA_INST_1[350].FA_  ( .A(A[862]), .B(n1887), .CI(
        C[862]), .S(S[862]), .CO(C[863]) );
  FA_11737 \FA_INST_0[1].FA_INST_1[351].FA_  ( .A(A[863]), .B(n1888), .CI(
        C[863]), .S(S[863]), .CO(C[864]) );
  FA_11736 \FA_INST_0[1].FA_INST_1[352].FA_  ( .A(A[864]), .B(n1889), .CI(
        C[864]), .S(S[864]), .CO(C[865]) );
  FA_11735 \FA_INST_0[1].FA_INST_1[353].FA_  ( .A(A[865]), .B(n1890), .CI(
        C[865]), .S(S[865]), .CO(C[866]) );
  FA_11734 \FA_INST_0[1].FA_INST_1[354].FA_  ( .A(A[866]), .B(n1891), .CI(
        C[866]), .S(S[866]), .CO(C[867]) );
  FA_11733 \FA_INST_0[1].FA_INST_1[355].FA_  ( .A(A[867]), .B(n1892), .CI(
        C[867]), .S(S[867]), .CO(C[868]) );
  FA_11732 \FA_INST_0[1].FA_INST_1[356].FA_  ( .A(A[868]), .B(n1893), .CI(
        C[868]), .S(S[868]), .CO(C[869]) );
  FA_11731 \FA_INST_0[1].FA_INST_1[357].FA_  ( .A(A[869]), .B(n1894), .CI(
        C[869]), .S(S[869]), .CO(C[870]) );
  FA_11730 \FA_INST_0[1].FA_INST_1[358].FA_  ( .A(A[870]), .B(n1895), .CI(
        C[870]), .S(S[870]), .CO(C[871]) );
  FA_11729 \FA_INST_0[1].FA_INST_1[359].FA_  ( .A(A[871]), .B(n1896), .CI(
        C[871]), .S(S[871]), .CO(C[872]) );
  FA_11728 \FA_INST_0[1].FA_INST_1[360].FA_  ( .A(A[872]), .B(n1897), .CI(
        C[872]), .S(S[872]), .CO(C[873]) );
  FA_11727 \FA_INST_0[1].FA_INST_1[361].FA_  ( .A(A[873]), .B(n1898), .CI(
        C[873]), .S(S[873]), .CO(C[874]) );
  FA_11726 \FA_INST_0[1].FA_INST_1[362].FA_  ( .A(A[874]), .B(n1899), .CI(
        C[874]), .S(S[874]), .CO(C[875]) );
  FA_11725 \FA_INST_0[1].FA_INST_1[363].FA_  ( .A(A[875]), .B(n1900), .CI(
        C[875]), .S(S[875]), .CO(C[876]) );
  FA_11724 \FA_INST_0[1].FA_INST_1[364].FA_  ( .A(A[876]), .B(n1901), .CI(
        C[876]), .S(S[876]), .CO(C[877]) );
  FA_11723 \FA_INST_0[1].FA_INST_1[365].FA_  ( .A(A[877]), .B(n1902), .CI(
        C[877]), .S(S[877]), .CO(C[878]) );
  FA_11722 \FA_INST_0[1].FA_INST_1[366].FA_  ( .A(A[878]), .B(n1903), .CI(
        C[878]), .S(S[878]), .CO(C[879]) );
  FA_11721 \FA_INST_0[1].FA_INST_1[367].FA_  ( .A(A[879]), .B(n1904), .CI(
        C[879]), .S(S[879]), .CO(C[880]) );
  FA_11720 \FA_INST_0[1].FA_INST_1[368].FA_  ( .A(A[880]), .B(n1905), .CI(
        C[880]), .S(S[880]), .CO(C[881]) );
  FA_11719 \FA_INST_0[1].FA_INST_1[369].FA_  ( .A(A[881]), .B(n1906), .CI(
        C[881]), .S(S[881]), .CO(C[882]) );
  FA_11718 \FA_INST_0[1].FA_INST_1[370].FA_  ( .A(A[882]), .B(n1907), .CI(
        C[882]), .S(S[882]), .CO(C[883]) );
  FA_11717 \FA_INST_0[1].FA_INST_1[371].FA_  ( .A(A[883]), .B(n1908), .CI(
        C[883]), .S(S[883]), .CO(C[884]) );
  FA_11716 \FA_INST_0[1].FA_INST_1[372].FA_  ( .A(A[884]), .B(n1909), .CI(
        C[884]), .S(S[884]), .CO(C[885]) );
  FA_11715 \FA_INST_0[1].FA_INST_1[373].FA_  ( .A(A[885]), .B(n1910), .CI(
        C[885]), .S(S[885]), .CO(C[886]) );
  FA_11714 \FA_INST_0[1].FA_INST_1[374].FA_  ( .A(A[886]), .B(n1911), .CI(
        C[886]), .S(S[886]), .CO(C[887]) );
  FA_11713 \FA_INST_0[1].FA_INST_1[375].FA_  ( .A(A[887]), .B(n1912), .CI(
        C[887]), .S(S[887]), .CO(C[888]) );
  FA_11712 \FA_INST_0[1].FA_INST_1[376].FA_  ( .A(A[888]), .B(n1913), .CI(
        C[888]), .S(S[888]), .CO(C[889]) );
  FA_11711 \FA_INST_0[1].FA_INST_1[377].FA_  ( .A(A[889]), .B(n1914), .CI(
        C[889]), .S(S[889]), .CO(C[890]) );
  FA_11710 \FA_INST_0[1].FA_INST_1[378].FA_  ( .A(A[890]), .B(n1915), .CI(
        C[890]), .S(S[890]), .CO(C[891]) );
  FA_11709 \FA_INST_0[1].FA_INST_1[379].FA_  ( .A(A[891]), .B(n1916), .CI(
        C[891]), .S(S[891]), .CO(C[892]) );
  FA_11708 \FA_INST_0[1].FA_INST_1[380].FA_  ( .A(A[892]), .B(n1917), .CI(
        C[892]), .S(S[892]), .CO(C[893]) );
  FA_11707 \FA_INST_0[1].FA_INST_1[381].FA_  ( .A(A[893]), .B(n1918), .CI(
        C[893]), .S(S[893]), .CO(C[894]) );
  FA_11706 \FA_INST_0[1].FA_INST_1[382].FA_  ( .A(A[894]), .B(n1919), .CI(
        C[894]), .S(S[894]), .CO(C[895]) );
  FA_11705 \FA_INST_0[1].FA_INST_1[383].FA_  ( .A(A[895]), .B(n1920), .CI(
        C[895]), .S(S[895]), .CO(C[896]) );
  FA_11704 \FA_INST_0[1].FA_INST_1[384].FA_  ( .A(A[896]), .B(n1921), .CI(
        C[896]), .S(S[896]), .CO(C[897]) );
  FA_11703 \FA_INST_0[1].FA_INST_1[385].FA_  ( .A(A[897]), .B(n1922), .CI(
        C[897]), .S(S[897]), .CO(C[898]) );
  FA_11702 \FA_INST_0[1].FA_INST_1[386].FA_  ( .A(A[898]), .B(n1923), .CI(
        C[898]), .S(S[898]), .CO(C[899]) );
  FA_11701 \FA_INST_0[1].FA_INST_1[387].FA_  ( .A(A[899]), .B(n1924), .CI(
        C[899]), .S(S[899]), .CO(C[900]) );
  FA_11700 \FA_INST_0[1].FA_INST_1[388].FA_  ( .A(A[900]), .B(n1925), .CI(
        C[900]), .S(S[900]), .CO(C[901]) );
  FA_11699 \FA_INST_0[1].FA_INST_1[389].FA_  ( .A(A[901]), .B(n1926), .CI(
        C[901]), .S(S[901]), .CO(C[902]) );
  FA_11698 \FA_INST_0[1].FA_INST_1[390].FA_  ( .A(A[902]), .B(n1927), .CI(
        C[902]), .S(S[902]), .CO(C[903]) );
  FA_11697 \FA_INST_0[1].FA_INST_1[391].FA_  ( .A(A[903]), .B(n1928), .CI(
        C[903]), .S(S[903]), .CO(C[904]) );
  FA_11696 \FA_INST_0[1].FA_INST_1[392].FA_  ( .A(A[904]), .B(n1929), .CI(
        C[904]), .S(S[904]), .CO(C[905]) );
  FA_11695 \FA_INST_0[1].FA_INST_1[393].FA_  ( .A(A[905]), .B(n1930), .CI(
        C[905]), .S(S[905]), .CO(C[906]) );
  FA_11694 \FA_INST_0[1].FA_INST_1[394].FA_  ( .A(A[906]), .B(n1931), .CI(
        C[906]), .S(S[906]), .CO(C[907]) );
  FA_11693 \FA_INST_0[1].FA_INST_1[395].FA_  ( .A(A[907]), .B(n1932), .CI(
        C[907]), .S(S[907]), .CO(C[908]) );
  FA_11692 \FA_INST_0[1].FA_INST_1[396].FA_  ( .A(A[908]), .B(n1933), .CI(
        C[908]), .S(S[908]), .CO(C[909]) );
  FA_11691 \FA_INST_0[1].FA_INST_1[397].FA_  ( .A(A[909]), .B(n1934), .CI(
        C[909]), .S(S[909]), .CO(C[910]) );
  FA_11690 \FA_INST_0[1].FA_INST_1[398].FA_  ( .A(A[910]), .B(n1935), .CI(
        C[910]), .S(S[910]), .CO(C[911]) );
  FA_11689 \FA_INST_0[1].FA_INST_1[399].FA_  ( .A(A[911]), .B(n1936), .CI(
        C[911]), .S(S[911]), .CO(C[912]) );
  FA_11688 \FA_INST_0[1].FA_INST_1[400].FA_  ( .A(A[912]), .B(n1937), .CI(
        C[912]), .S(S[912]), .CO(C[913]) );
  FA_11687 \FA_INST_0[1].FA_INST_1[401].FA_  ( .A(A[913]), .B(n1938), .CI(
        C[913]), .S(S[913]), .CO(C[914]) );
  FA_11686 \FA_INST_0[1].FA_INST_1[402].FA_  ( .A(A[914]), .B(n1939), .CI(
        C[914]), .S(S[914]), .CO(C[915]) );
  FA_11685 \FA_INST_0[1].FA_INST_1[403].FA_  ( .A(A[915]), .B(n1940), .CI(
        C[915]), .S(S[915]), .CO(C[916]) );
  FA_11684 \FA_INST_0[1].FA_INST_1[404].FA_  ( .A(A[916]), .B(n1941), .CI(
        C[916]), .S(S[916]), .CO(C[917]) );
  FA_11683 \FA_INST_0[1].FA_INST_1[405].FA_  ( .A(A[917]), .B(n1942), .CI(
        C[917]), .S(S[917]), .CO(C[918]) );
  FA_11682 \FA_INST_0[1].FA_INST_1[406].FA_  ( .A(A[918]), .B(n1943), .CI(
        C[918]), .S(S[918]), .CO(C[919]) );
  FA_11681 \FA_INST_0[1].FA_INST_1[407].FA_  ( .A(A[919]), .B(n1944), .CI(
        C[919]), .S(S[919]), .CO(C[920]) );
  FA_11680 \FA_INST_0[1].FA_INST_1[408].FA_  ( .A(A[920]), .B(n1945), .CI(
        C[920]), .S(S[920]), .CO(C[921]) );
  FA_11679 \FA_INST_0[1].FA_INST_1[409].FA_  ( .A(A[921]), .B(n1946), .CI(
        C[921]), .S(S[921]), .CO(C[922]) );
  FA_11678 \FA_INST_0[1].FA_INST_1[410].FA_  ( .A(A[922]), .B(n1947), .CI(
        C[922]), .S(S[922]), .CO(C[923]) );
  FA_11677 \FA_INST_0[1].FA_INST_1[411].FA_  ( .A(A[923]), .B(n1948), .CI(
        C[923]), .S(S[923]), .CO(C[924]) );
  FA_11676 \FA_INST_0[1].FA_INST_1[412].FA_  ( .A(A[924]), .B(n1949), .CI(
        C[924]), .S(S[924]), .CO(C[925]) );
  FA_11675 \FA_INST_0[1].FA_INST_1[413].FA_  ( .A(A[925]), .B(n1950), .CI(
        C[925]), .S(S[925]), .CO(C[926]) );
  FA_11674 \FA_INST_0[1].FA_INST_1[414].FA_  ( .A(A[926]), .B(n1951), .CI(
        C[926]), .S(S[926]), .CO(C[927]) );
  FA_11673 \FA_INST_0[1].FA_INST_1[415].FA_  ( .A(A[927]), .B(n1952), .CI(
        C[927]), .S(S[927]), .CO(C[928]) );
  FA_11672 \FA_INST_0[1].FA_INST_1[416].FA_  ( .A(A[928]), .B(n1953), .CI(
        C[928]), .S(S[928]), .CO(C[929]) );
  FA_11671 \FA_INST_0[1].FA_INST_1[417].FA_  ( .A(A[929]), .B(n1954), .CI(
        C[929]), .S(S[929]), .CO(C[930]) );
  FA_11670 \FA_INST_0[1].FA_INST_1[418].FA_  ( .A(A[930]), .B(n1955), .CI(
        C[930]), .S(S[930]), .CO(C[931]) );
  FA_11669 \FA_INST_0[1].FA_INST_1[419].FA_  ( .A(A[931]), .B(n1956), .CI(
        C[931]), .S(S[931]), .CO(C[932]) );
  FA_11668 \FA_INST_0[1].FA_INST_1[420].FA_  ( .A(A[932]), .B(n1957), .CI(
        C[932]), .S(S[932]), .CO(C[933]) );
  FA_11667 \FA_INST_0[1].FA_INST_1[421].FA_  ( .A(A[933]), .B(n1958), .CI(
        C[933]), .S(S[933]), .CO(C[934]) );
  FA_11666 \FA_INST_0[1].FA_INST_1[422].FA_  ( .A(A[934]), .B(n1959), .CI(
        C[934]), .S(S[934]), .CO(C[935]) );
  FA_11665 \FA_INST_0[1].FA_INST_1[423].FA_  ( .A(A[935]), .B(n1960), .CI(
        C[935]), .S(S[935]), .CO(C[936]) );
  FA_11664 \FA_INST_0[1].FA_INST_1[424].FA_  ( .A(A[936]), .B(n1961), .CI(
        C[936]), .S(S[936]), .CO(C[937]) );
  FA_11663 \FA_INST_0[1].FA_INST_1[425].FA_  ( .A(A[937]), .B(n1962), .CI(
        C[937]), .S(S[937]), .CO(C[938]) );
  FA_11662 \FA_INST_0[1].FA_INST_1[426].FA_  ( .A(A[938]), .B(n1963), .CI(
        C[938]), .S(S[938]), .CO(C[939]) );
  FA_11661 \FA_INST_0[1].FA_INST_1[427].FA_  ( .A(A[939]), .B(n1964), .CI(
        C[939]), .S(S[939]), .CO(C[940]) );
  FA_11660 \FA_INST_0[1].FA_INST_1[428].FA_  ( .A(A[940]), .B(n1965), .CI(
        C[940]), .S(S[940]), .CO(C[941]) );
  FA_11659 \FA_INST_0[1].FA_INST_1[429].FA_  ( .A(A[941]), .B(n1966), .CI(
        C[941]), .S(S[941]), .CO(C[942]) );
  FA_11658 \FA_INST_0[1].FA_INST_1[430].FA_  ( .A(A[942]), .B(n1967), .CI(
        C[942]), .S(S[942]), .CO(C[943]) );
  FA_11657 \FA_INST_0[1].FA_INST_1[431].FA_  ( .A(A[943]), .B(n1968), .CI(
        C[943]), .S(S[943]), .CO(C[944]) );
  FA_11656 \FA_INST_0[1].FA_INST_1[432].FA_  ( .A(A[944]), .B(n1969), .CI(
        C[944]), .S(S[944]), .CO(C[945]) );
  FA_11655 \FA_INST_0[1].FA_INST_1[433].FA_  ( .A(A[945]), .B(n1970), .CI(
        C[945]), .S(S[945]), .CO(C[946]) );
  FA_11654 \FA_INST_0[1].FA_INST_1[434].FA_  ( .A(A[946]), .B(n1971), .CI(
        C[946]), .S(S[946]), .CO(C[947]) );
  FA_11653 \FA_INST_0[1].FA_INST_1[435].FA_  ( .A(A[947]), .B(n1972), .CI(
        C[947]), .S(S[947]), .CO(C[948]) );
  FA_11652 \FA_INST_0[1].FA_INST_1[436].FA_  ( .A(A[948]), .B(n1973), .CI(
        C[948]), .S(S[948]), .CO(C[949]) );
  FA_11651 \FA_INST_0[1].FA_INST_1[437].FA_  ( .A(A[949]), .B(n1974), .CI(
        C[949]), .S(S[949]), .CO(C[950]) );
  FA_11650 \FA_INST_0[1].FA_INST_1[438].FA_  ( .A(A[950]), .B(n1975), .CI(
        C[950]), .S(S[950]), .CO(C[951]) );
  FA_11649 \FA_INST_0[1].FA_INST_1[439].FA_  ( .A(A[951]), .B(n1976), .CI(
        C[951]), .S(S[951]), .CO(C[952]) );
  FA_11648 \FA_INST_0[1].FA_INST_1[440].FA_  ( .A(A[952]), .B(n1977), .CI(
        C[952]), .S(S[952]), .CO(C[953]) );
  FA_11647 \FA_INST_0[1].FA_INST_1[441].FA_  ( .A(A[953]), .B(n1978), .CI(
        C[953]), .S(S[953]), .CO(C[954]) );
  FA_11646 \FA_INST_0[1].FA_INST_1[442].FA_  ( .A(A[954]), .B(n1979), .CI(
        C[954]), .S(S[954]), .CO(C[955]) );
  FA_11645 \FA_INST_0[1].FA_INST_1[443].FA_  ( .A(A[955]), .B(n1980), .CI(
        C[955]), .S(S[955]), .CO(C[956]) );
  FA_11644 \FA_INST_0[1].FA_INST_1[444].FA_  ( .A(A[956]), .B(n1981), .CI(
        C[956]), .S(S[956]), .CO(C[957]) );
  FA_11643 \FA_INST_0[1].FA_INST_1[445].FA_  ( .A(A[957]), .B(n1982), .CI(
        C[957]), .S(S[957]), .CO(C[958]) );
  FA_11642 \FA_INST_0[1].FA_INST_1[446].FA_  ( .A(A[958]), .B(n1983), .CI(
        C[958]), .S(S[958]), .CO(C[959]) );
  FA_11641 \FA_INST_0[1].FA_INST_1[447].FA_  ( .A(A[959]), .B(n1984), .CI(
        C[959]), .S(S[959]), .CO(C[960]) );
  FA_11640 \FA_INST_0[1].FA_INST_1[448].FA_  ( .A(A[960]), .B(n1985), .CI(
        C[960]), .S(S[960]), .CO(C[961]) );
  FA_11639 \FA_INST_0[1].FA_INST_1[449].FA_  ( .A(A[961]), .B(n1986), .CI(
        C[961]), .S(S[961]), .CO(C[962]) );
  FA_11638 \FA_INST_0[1].FA_INST_1[450].FA_  ( .A(A[962]), .B(n1987), .CI(
        C[962]), .S(S[962]), .CO(C[963]) );
  FA_11637 \FA_INST_0[1].FA_INST_1[451].FA_  ( .A(A[963]), .B(n1988), .CI(
        C[963]), .S(S[963]), .CO(C[964]) );
  FA_11636 \FA_INST_0[1].FA_INST_1[452].FA_  ( .A(A[964]), .B(n1989), .CI(
        C[964]), .S(S[964]), .CO(C[965]) );
  FA_11635 \FA_INST_0[1].FA_INST_1[453].FA_  ( .A(A[965]), .B(n1990), .CI(
        C[965]), .S(S[965]), .CO(C[966]) );
  FA_11634 \FA_INST_0[1].FA_INST_1[454].FA_  ( .A(A[966]), .B(n1991), .CI(
        C[966]), .S(S[966]), .CO(C[967]) );
  FA_11633 \FA_INST_0[1].FA_INST_1[455].FA_  ( .A(A[967]), .B(n1992), .CI(
        C[967]), .S(S[967]), .CO(C[968]) );
  FA_11632 \FA_INST_0[1].FA_INST_1[456].FA_  ( .A(A[968]), .B(n1993), .CI(
        C[968]), .S(S[968]), .CO(C[969]) );
  FA_11631 \FA_INST_0[1].FA_INST_1[457].FA_  ( .A(A[969]), .B(n1994), .CI(
        C[969]), .S(S[969]), .CO(C[970]) );
  FA_11630 \FA_INST_0[1].FA_INST_1[458].FA_  ( .A(A[970]), .B(n1995), .CI(
        C[970]), .S(S[970]), .CO(C[971]) );
  FA_11629 \FA_INST_0[1].FA_INST_1[459].FA_  ( .A(A[971]), .B(n1996), .CI(
        C[971]), .S(S[971]), .CO(C[972]) );
  FA_11628 \FA_INST_0[1].FA_INST_1[460].FA_  ( .A(A[972]), .B(n1997), .CI(
        C[972]), .S(S[972]), .CO(C[973]) );
  FA_11627 \FA_INST_0[1].FA_INST_1[461].FA_  ( .A(A[973]), .B(n1998), .CI(
        C[973]), .S(S[973]), .CO(C[974]) );
  FA_11626 \FA_INST_0[1].FA_INST_1[462].FA_  ( .A(A[974]), .B(n1999), .CI(
        C[974]), .S(S[974]), .CO(C[975]) );
  FA_11625 \FA_INST_0[1].FA_INST_1[463].FA_  ( .A(A[975]), .B(n2000), .CI(
        C[975]), .S(S[975]), .CO(C[976]) );
  FA_11624 \FA_INST_0[1].FA_INST_1[464].FA_  ( .A(A[976]), .B(n2001), .CI(
        C[976]), .S(S[976]), .CO(C[977]) );
  FA_11623 \FA_INST_0[1].FA_INST_1[465].FA_  ( .A(A[977]), .B(n2002), .CI(
        C[977]), .S(S[977]), .CO(C[978]) );
  FA_11622 \FA_INST_0[1].FA_INST_1[466].FA_  ( .A(A[978]), .B(n2003), .CI(
        C[978]), .S(S[978]), .CO(C[979]) );
  FA_11621 \FA_INST_0[1].FA_INST_1[467].FA_  ( .A(A[979]), .B(n2004), .CI(
        C[979]), .S(S[979]), .CO(C[980]) );
  FA_11620 \FA_INST_0[1].FA_INST_1[468].FA_  ( .A(A[980]), .B(n2005), .CI(
        C[980]), .S(S[980]), .CO(C[981]) );
  FA_11619 \FA_INST_0[1].FA_INST_1[469].FA_  ( .A(A[981]), .B(n2006), .CI(
        C[981]), .S(S[981]), .CO(C[982]) );
  FA_11618 \FA_INST_0[1].FA_INST_1[470].FA_  ( .A(A[982]), .B(n2007), .CI(
        C[982]), .S(S[982]), .CO(C[983]) );
  FA_11617 \FA_INST_0[1].FA_INST_1[471].FA_  ( .A(A[983]), .B(n2008), .CI(
        C[983]), .S(S[983]), .CO(C[984]) );
  FA_11616 \FA_INST_0[1].FA_INST_1[472].FA_  ( .A(A[984]), .B(n2009), .CI(
        C[984]), .S(S[984]), .CO(C[985]) );
  FA_11615 \FA_INST_0[1].FA_INST_1[473].FA_  ( .A(A[985]), .B(n2010), .CI(
        C[985]), .S(S[985]), .CO(C[986]) );
  FA_11614 \FA_INST_0[1].FA_INST_1[474].FA_  ( .A(A[986]), .B(n2011), .CI(
        C[986]), .S(S[986]), .CO(C[987]) );
  FA_11613 \FA_INST_0[1].FA_INST_1[475].FA_  ( .A(A[987]), .B(n2012), .CI(
        C[987]), .S(S[987]), .CO(C[988]) );
  FA_11612 \FA_INST_0[1].FA_INST_1[476].FA_  ( .A(A[988]), .B(n2013), .CI(
        C[988]), .S(S[988]), .CO(C[989]) );
  FA_11611 \FA_INST_0[1].FA_INST_1[477].FA_  ( .A(A[989]), .B(n2014), .CI(
        C[989]), .S(S[989]), .CO(C[990]) );
  FA_11610 \FA_INST_0[1].FA_INST_1[478].FA_  ( .A(A[990]), .B(n2015), .CI(
        C[990]), .S(S[990]), .CO(C[991]) );
  FA_11609 \FA_INST_0[1].FA_INST_1[479].FA_  ( .A(A[991]), .B(n2016), .CI(
        C[991]), .S(S[991]), .CO(C[992]) );
  FA_11608 \FA_INST_0[1].FA_INST_1[480].FA_  ( .A(A[992]), .B(n2017), .CI(
        C[992]), .S(S[992]), .CO(C[993]) );
  FA_11607 \FA_INST_0[1].FA_INST_1[481].FA_  ( .A(A[993]), .B(n2018), .CI(
        C[993]), .S(S[993]), .CO(C[994]) );
  FA_11606 \FA_INST_0[1].FA_INST_1[482].FA_  ( .A(A[994]), .B(n2019), .CI(
        C[994]), .S(S[994]), .CO(C[995]) );
  FA_11605 \FA_INST_0[1].FA_INST_1[483].FA_  ( .A(A[995]), .B(n2020), .CI(
        C[995]), .S(S[995]), .CO(C[996]) );
  FA_11604 \FA_INST_0[1].FA_INST_1[484].FA_  ( .A(A[996]), .B(n2021), .CI(
        C[996]), .S(S[996]), .CO(C[997]) );
  FA_11603 \FA_INST_0[1].FA_INST_1[485].FA_  ( .A(A[997]), .B(n2022), .CI(
        C[997]), .S(S[997]), .CO(C[998]) );
  FA_11602 \FA_INST_0[1].FA_INST_1[486].FA_  ( .A(A[998]), .B(n2023), .CI(
        C[998]), .S(S[998]), .CO(C[999]) );
  FA_11601 \FA_INST_0[1].FA_INST_1[487].FA_  ( .A(A[999]), .B(n2024), .CI(
        C[999]), .S(S[999]), .CO(C[1000]) );
  FA_11600 \FA_INST_0[1].FA_INST_1[488].FA_  ( .A(A[1000]), .B(n2025), .CI(
        C[1000]), .S(S[1000]), .CO(C[1001]) );
  FA_11599 \FA_INST_0[1].FA_INST_1[489].FA_  ( .A(A[1001]), .B(n2026), .CI(
        C[1001]), .S(S[1001]), .CO(C[1002]) );
  FA_11598 \FA_INST_0[1].FA_INST_1[490].FA_  ( .A(A[1002]), .B(n2027), .CI(
        C[1002]), .S(S[1002]), .CO(C[1003]) );
  FA_11597 \FA_INST_0[1].FA_INST_1[491].FA_  ( .A(A[1003]), .B(n2028), .CI(
        C[1003]), .S(S[1003]), .CO(C[1004]) );
  FA_11596 \FA_INST_0[1].FA_INST_1[492].FA_  ( .A(A[1004]), .B(n2029), .CI(
        C[1004]), .S(S[1004]), .CO(C[1005]) );
  FA_11595 \FA_INST_0[1].FA_INST_1[493].FA_  ( .A(A[1005]), .B(n2030), .CI(
        C[1005]), .S(S[1005]), .CO(C[1006]) );
  FA_11594 \FA_INST_0[1].FA_INST_1[494].FA_  ( .A(A[1006]), .B(n2031), .CI(
        C[1006]), .S(S[1006]), .CO(C[1007]) );
  FA_11593 \FA_INST_0[1].FA_INST_1[495].FA_  ( .A(A[1007]), .B(n2032), .CI(
        C[1007]), .S(S[1007]), .CO(C[1008]) );
  FA_11592 \FA_INST_0[1].FA_INST_1[496].FA_  ( .A(A[1008]), .B(n2033), .CI(
        C[1008]), .S(S[1008]), .CO(C[1009]) );
  FA_11591 \FA_INST_0[1].FA_INST_1[497].FA_  ( .A(A[1009]), .B(n2034), .CI(
        C[1009]), .S(S[1009]), .CO(C[1010]) );
  FA_11590 \FA_INST_0[1].FA_INST_1[498].FA_  ( .A(A[1010]), .B(n2035), .CI(
        C[1010]), .S(S[1010]), .CO(C[1011]) );
  FA_11589 \FA_INST_0[1].FA_INST_1[499].FA_  ( .A(A[1011]), .B(n2036), .CI(
        C[1011]), .S(S[1011]), .CO(C[1012]) );
  FA_11588 \FA_INST_0[1].FA_INST_1[500].FA_  ( .A(A[1012]), .B(n2037), .CI(
        C[1012]), .S(S[1012]), .CO(C[1013]) );
  FA_11587 \FA_INST_0[1].FA_INST_1[501].FA_  ( .A(A[1013]), .B(n2038), .CI(
        C[1013]), .S(S[1013]), .CO(C[1014]) );
  FA_11586 \FA_INST_0[1].FA_INST_1[502].FA_  ( .A(A[1014]), .B(n2039), .CI(
        C[1014]), .S(S[1014]), .CO(C[1015]) );
  FA_11585 \FA_INST_0[1].FA_INST_1[503].FA_  ( .A(A[1015]), .B(n2040), .CI(
        C[1015]), .S(S[1015]), .CO(C[1016]) );
  FA_11584 \FA_INST_0[1].FA_INST_1[504].FA_  ( .A(A[1016]), .B(n2041), .CI(
        C[1016]), .S(S[1016]), .CO(C[1017]) );
  FA_11583 \FA_INST_0[1].FA_INST_1[505].FA_  ( .A(A[1017]), .B(n2042), .CI(
        C[1017]), .S(S[1017]), .CO(C[1018]) );
  FA_11582 \FA_INST_0[1].FA_INST_1[506].FA_  ( .A(A[1018]), .B(n2043), .CI(
        C[1018]), .S(S[1018]), .CO(C[1019]) );
  FA_11581 \FA_INST_0[1].FA_INST_1[507].FA_  ( .A(A[1019]), .B(n2044), .CI(
        C[1019]), .S(S[1019]), .CO(C[1020]) );
  FA_11580 \FA_INST_0[1].FA_INST_1[508].FA_  ( .A(A[1020]), .B(n2045), .CI(
        C[1020]), .S(S[1020]), .CO(C[1021]) );
  FA_11579 \FA_INST_0[1].FA_INST_1[509].FA_  ( .A(A[1021]), .B(n2046), .CI(
        C[1021]), .S(S[1021]), .CO(C[1022]) );
  FA_11578 \FA_INST_0[1].FA_INST_1[510].FA_  ( .A(A[1022]), .B(n2047), .CI(
        C[1022]), .S(S[1022]), .CO(C[1023]) );
  FA_11577 \FA_INST_0[1].FA_INST_1[511].FA_  ( .A(A[1023]), .B(n2048), .CI(
        C[1023]), .S(S[1023]), .CO(C[1024]) );
  FA_11576 \FA_INST_1[1024].FA_  ( .A(A[1024]), .B(1'b1), .CI(C[1024]), .S(
        S[1024]) );
  IV U2 ( .A(B[27]), .Z(n1052) );
  IV U3 ( .A(B[28]), .Z(n1053) );
  IV U4 ( .A(B[29]), .Z(n1054) );
  IV U5 ( .A(B[30]), .Z(n1055) );
  IV U6 ( .A(B[31]), .Z(n1056) );
  IV U7 ( .A(B[32]), .Z(n1057) );
  IV U8 ( .A(B[33]), .Z(n1058) );
  IV U9 ( .A(B[34]), .Z(n1059) );
  IV U10 ( .A(B[35]), .Z(n1060) );
  IV U11 ( .A(B[36]), .Z(n1061) );
  IV U12 ( .A(B[927]), .Z(n1952) );
  IV U13 ( .A(B[37]), .Z(n1062) );
  IV U14 ( .A(B[38]), .Z(n1063) );
  IV U15 ( .A(B[39]), .Z(n1064) );
  IV U16 ( .A(B[40]), .Z(n1065) );
  IV U17 ( .A(B[41]), .Z(n1066) );
  IV U18 ( .A(B[42]), .Z(n1067) );
  IV U19 ( .A(B[43]), .Z(n1068) );
  IV U20 ( .A(B[44]), .Z(n1069) );
  IV U21 ( .A(B[45]), .Z(n1070) );
  IV U22 ( .A(B[46]), .Z(n1071) );
  IV U23 ( .A(B[928]), .Z(n1953) );
  IV U24 ( .A(B[47]), .Z(n1072) );
  IV U25 ( .A(B[48]), .Z(n1073) );
  IV U26 ( .A(B[49]), .Z(n1074) );
  IV U27 ( .A(B[50]), .Z(n1075) );
  IV U28 ( .A(B[51]), .Z(n1076) );
  IV U29 ( .A(B[52]), .Z(n1077) );
  IV U30 ( .A(B[53]), .Z(n1078) );
  IV U31 ( .A(B[54]), .Z(n1079) );
  IV U32 ( .A(B[55]), .Z(n1080) );
  IV U33 ( .A(B[56]), .Z(n1081) );
  IV U34 ( .A(B[929]), .Z(n1954) );
  IV U35 ( .A(B[57]), .Z(n1082) );
  IV U36 ( .A(B[58]), .Z(n1083) );
  IV U37 ( .A(B[59]), .Z(n1084) );
  IV U38 ( .A(B[60]), .Z(n1085) );
  IV U39 ( .A(B[61]), .Z(n1086) );
  IV U40 ( .A(B[62]), .Z(n1087) );
  IV U41 ( .A(B[63]), .Z(n1088) );
  IV U42 ( .A(B[64]), .Z(n1089) );
  IV U43 ( .A(B[65]), .Z(n1090) );
  IV U44 ( .A(B[66]), .Z(n1091) );
  IV U45 ( .A(B[930]), .Z(n1955) );
  IV U46 ( .A(B[67]), .Z(n1092) );
  IV U47 ( .A(B[68]), .Z(n1093) );
  IV U48 ( .A(B[69]), .Z(n1094) );
  IV U49 ( .A(B[70]), .Z(n1095) );
  IV U50 ( .A(B[71]), .Z(n1096) );
  IV U51 ( .A(B[72]), .Z(n1097) );
  IV U52 ( .A(B[73]), .Z(n1098) );
  IV U53 ( .A(B[74]), .Z(n1099) );
  IV U54 ( .A(B[75]), .Z(n1100) );
  IV U55 ( .A(B[76]), .Z(n1101) );
  IV U56 ( .A(B[931]), .Z(n1956) );
  IV U57 ( .A(B[77]), .Z(n1102) );
  IV U58 ( .A(B[78]), .Z(n1103) );
  IV U59 ( .A(B[79]), .Z(n1104) );
  IV U60 ( .A(B[80]), .Z(n1105) );
  IV U61 ( .A(B[81]), .Z(n1106) );
  IV U62 ( .A(B[82]), .Z(n1107) );
  IV U63 ( .A(B[83]), .Z(n1108) );
  IV U64 ( .A(B[84]), .Z(n1109) );
  IV U65 ( .A(B[85]), .Z(n1110) );
  IV U66 ( .A(B[86]), .Z(n1111) );
  IV U67 ( .A(B[932]), .Z(n1957) );
  IV U68 ( .A(B[87]), .Z(n1112) );
  IV U69 ( .A(B[88]), .Z(n1113) );
  IV U70 ( .A(B[89]), .Z(n1114) );
  IV U71 ( .A(B[90]), .Z(n1115) );
  IV U72 ( .A(B[91]), .Z(n1116) );
  IV U73 ( .A(B[92]), .Z(n1117) );
  IV U74 ( .A(B[93]), .Z(n1118) );
  IV U75 ( .A(B[94]), .Z(n1119) );
  IV U76 ( .A(B[95]), .Z(n1120) );
  IV U77 ( .A(B[96]), .Z(n1121) );
  IV U78 ( .A(B[933]), .Z(n1958) );
  IV U79 ( .A(B[97]), .Z(n1122) );
  IV U80 ( .A(B[98]), .Z(n1123) );
  IV U81 ( .A(B[99]), .Z(n1124) );
  IV U82 ( .A(B[100]), .Z(n1125) );
  IV U83 ( .A(B[101]), .Z(n1126) );
  IV U84 ( .A(B[102]), .Z(n1127) );
  IV U85 ( .A(B[103]), .Z(n1128) );
  IV U86 ( .A(B[104]), .Z(n1129) );
  IV U87 ( .A(B[105]), .Z(n1130) );
  IV U88 ( .A(B[106]), .Z(n1131) );
  IV U89 ( .A(B[934]), .Z(n1959) );
  IV U90 ( .A(B[107]), .Z(n1132) );
  IV U91 ( .A(B[108]), .Z(n1133) );
  IV U92 ( .A(B[109]), .Z(n1134) );
  IV U93 ( .A(B[110]), .Z(n1135) );
  IV U94 ( .A(B[111]), .Z(n1136) );
  IV U95 ( .A(B[112]), .Z(n1137) );
  IV U96 ( .A(B[113]), .Z(n1138) );
  IV U97 ( .A(B[114]), .Z(n1139) );
  IV U98 ( .A(B[115]), .Z(n1140) );
  IV U99 ( .A(B[116]), .Z(n1141) );
  IV U100 ( .A(B[935]), .Z(n1960) );
  IV U101 ( .A(B[117]), .Z(n1142) );
  IV U102 ( .A(B[118]), .Z(n1143) );
  IV U103 ( .A(B[119]), .Z(n1144) );
  IV U104 ( .A(B[120]), .Z(n1145) );
  IV U105 ( .A(B[121]), .Z(n1146) );
  IV U106 ( .A(B[122]), .Z(n1147) );
  IV U107 ( .A(B[123]), .Z(n1148) );
  IV U108 ( .A(B[124]), .Z(n1149) );
  IV U109 ( .A(B[125]), .Z(n1150) );
  IV U110 ( .A(B[126]), .Z(n1151) );
  IV U111 ( .A(B[936]), .Z(n1961) );
  IV U112 ( .A(B[1017]), .Z(n2042) );
  IV U113 ( .A(B[127]), .Z(n1152) );
  IV U114 ( .A(B[128]), .Z(n1153) );
  IV U115 ( .A(B[129]), .Z(n1154) );
  IV U116 ( .A(B[130]), .Z(n1155) );
  IV U117 ( .A(B[131]), .Z(n1156) );
  IV U118 ( .A(B[132]), .Z(n1157) );
  IV U119 ( .A(B[133]), .Z(n1158) );
  IV U120 ( .A(B[134]), .Z(n1159) );
  IV U121 ( .A(B[135]), .Z(n1160) );
  IV U122 ( .A(B[136]), .Z(n1161) );
  IV U123 ( .A(B[937]), .Z(n1962) );
  IV U124 ( .A(B[137]), .Z(n1162) );
  IV U125 ( .A(B[138]), .Z(n1163) );
  IV U126 ( .A(B[139]), .Z(n1164) );
  IV U127 ( .A(B[140]), .Z(n1165) );
  IV U128 ( .A(B[141]), .Z(n1166) );
  IV U129 ( .A(B[142]), .Z(n1167) );
  IV U130 ( .A(B[143]), .Z(n1168) );
  IV U131 ( .A(B[144]), .Z(n1169) );
  IV U132 ( .A(B[145]), .Z(n1170) );
  IV U133 ( .A(B[146]), .Z(n1171) );
  IV U134 ( .A(B[938]), .Z(n1963) );
  IV U135 ( .A(B[147]), .Z(n1172) );
  IV U136 ( .A(B[148]), .Z(n1173) );
  IV U137 ( .A(B[149]), .Z(n1174) );
  IV U138 ( .A(B[150]), .Z(n1175) );
  IV U139 ( .A(B[151]), .Z(n1176) );
  IV U140 ( .A(B[152]), .Z(n1177) );
  IV U141 ( .A(B[153]), .Z(n1178) );
  IV U142 ( .A(B[154]), .Z(n1179) );
  IV U143 ( .A(B[155]), .Z(n1180) );
  IV U144 ( .A(B[156]), .Z(n1181) );
  IV U145 ( .A(B[939]), .Z(n1964) );
  IV U146 ( .A(B[157]), .Z(n1182) );
  IV U147 ( .A(B[158]), .Z(n1183) );
  IV U148 ( .A(B[159]), .Z(n1184) );
  IV U149 ( .A(B[160]), .Z(n1185) );
  IV U150 ( .A(B[161]), .Z(n1186) );
  IV U151 ( .A(B[162]), .Z(n1187) );
  IV U152 ( .A(B[163]), .Z(n1188) );
  IV U153 ( .A(B[164]), .Z(n1189) );
  IV U154 ( .A(B[165]), .Z(n1190) );
  IV U155 ( .A(B[166]), .Z(n1191) );
  IV U156 ( .A(B[940]), .Z(n1965) );
  IV U157 ( .A(B[167]), .Z(n1192) );
  IV U158 ( .A(B[168]), .Z(n1193) );
  IV U159 ( .A(B[169]), .Z(n1194) );
  IV U160 ( .A(B[170]), .Z(n1195) );
  IV U161 ( .A(B[171]), .Z(n1196) );
  IV U162 ( .A(B[172]), .Z(n1197) );
  IV U163 ( .A(B[173]), .Z(n1198) );
  IV U164 ( .A(B[174]), .Z(n1199) );
  IV U165 ( .A(B[175]), .Z(n1200) );
  IV U166 ( .A(B[176]), .Z(n1201) );
  IV U167 ( .A(B[941]), .Z(n1966) );
  IV U168 ( .A(B[177]), .Z(n1202) );
  IV U169 ( .A(B[178]), .Z(n1203) );
  IV U170 ( .A(B[179]), .Z(n1204) );
  IV U171 ( .A(B[180]), .Z(n1205) );
  IV U172 ( .A(B[181]), .Z(n1206) );
  IV U173 ( .A(B[182]), .Z(n1207) );
  IV U174 ( .A(B[183]), .Z(n1208) );
  IV U175 ( .A(B[184]), .Z(n1209) );
  IV U176 ( .A(B[185]), .Z(n1210) );
  IV U177 ( .A(B[186]), .Z(n1211) );
  IV U178 ( .A(B[942]), .Z(n1967) );
  IV U179 ( .A(B[187]), .Z(n1212) );
  IV U180 ( .A(B[188]), .Z(n1213) );
  IV U181 ( .A(B[189]), .Z(n1214) );
  IV U182 ( .A(B[190]), .Z(n1215) );
  IV U183 ( .A(B[191]), .Z(n1216) );
  IV U184 ( .A(B[192]), .Z(n1217) );
  IV U185 ( .A(B[193]), .Z(n1218) );
  IV U186 ( .A(B[194]), .Z(n1219) );
  IV U187 ( .A(B[195]), .Z(n1220) );
  IV U188 ( .A(B[196]), .Z(n1221) );
  IV U189 ( .A(B[943]), .Z(n1968) );
  IV U190 ( .A(B[197]), .Z(n1222) );
  IV U191 ( .A(B[198]), .Z(n1223) );
  IV U192 ( .A(B[199]), .Z(n1224) );
  IV U193 ( .A(B[200]), .Z(n1225) );
  IV U194 ( .A(B[201]), .Z(n1226) );
  IV U195 ( .A(B[202]), .Z(n1227) );
  IV U196 ( .A(B[203]), .Z(n1228) );
  IV U197 ( .A(B[204]), .Z(n1229) );
  IV U198 ( .A(B[205]), .Z(n1230) );
  IV U199 ( .A(B[206]), .Z(n1231) );
  IV U200 ( .A(B[944]), .Z(n1969) );
  IV U201 ( .A(B[207]), .Z(n1232) );
  IV U202 ( .A(B[208]), .Z(n1233) );
  IV U203 ( .A(B[209]), .Z(n1234) );
  IV U204 ( .A(B[210]), .Z(n1235) );
  IV U205 ( .A(B[211]), .Z(n1236) );
  IV U206 ( .A(B[212]), .Z(n1237) );
  IV U207 ( .A(B[213]), .Z(n1238) );
  IV U208 ( .A(B[214]), .Z(n1239) );
  IV U209 ( .A(B[215]), .Z(n1240) );
  IV U210 ( .A(B[216]), .Z(n1241) );
  IV U211 ( .A(B[945]), .Z(n1970) );
  IV U212 ( .A(B[217]), .Z(n1242) );
  IV U213 ( .A(B[218]), .Z(n1243) );
  IV U214 ( .A(B[219]), .Z(n1244) );
  IV U215 ( .A(B[220]), .Z(n1245) );
  IV U216 ( .A(B[221]), .Z(n1246) );
  IV U217 ( .A(B[222]), .Z(n1247) );
  IV U218 ( .A(B[223]), .Z(n1248) );
  IV U219 ( .A(B[224]), .Z(n1249) );
  IV U220 ( .A(B[225]), .Z(n1250) );
  IV U221 ( .A(B[226]), .Z(n1251) );
  IV U222 ( .A(B[946]), .Z(n1971) );
  IV U223 ( .A(B[1018]), .Z(n2043) );
  IV U224 ( .A(B[227]), .Z(n1252) );
  IV U225 ( .A(B[228]), .Z(n1253) );
  IV U226 ( .A(B[229]), .Z(n1254) );
  IV U227 ( .A(B[230]), .Z(n1255) );
  IV U228 ( .A(B[231]), .Z(n1256) );
  IV U229 ( .A(B[232]), .Z(n1257) );
  IV U230 ( .A(B[233]), .Z(n1258) );
  IV U231 ( .A(B[234]), .Z(n1259) );
  IV U232 ( .A(B[235]), .Z(n1260) );
  IV U233 ( .A(B[236]), .Z(n1261) );
  IV U234 ( .A(B[947]), .Z(n1972) );
  IV U235 ( .A(B[237]), .Z(n1262) );
  IV U236 ( .A(B[238]), .Z(n1263) );
  IV U237 ( .A(B[239]), .Z(n1264) );
  IV U238 ( .A(B[240]), .Z(n1265) );
  IV U239 ( .A(B[241]), .Z(n1266) );
  IV U240 ( .A(B[242]), .Z(n1267) );
  IV U241 ( .A(B[243]), .Z(n1268) );
  IV U242 ( .A(B[244]), .Z(n1269) );
  IV U243 ( .A(B[245]), .Z(n1270) );
  IV U244 ( .A(B[246]), .Z(n1271) );
  IV U245 ( .A(B[948]), .Z(n1973) );
  IV U246 ( .A(B[247]), .Z(n1272) );
  IV U247 ( .A(B[248]), .Z(n1273) );
  IV U248 ( .A(B[249]), .Z(n1274) );
  IV U249 ( .A(B[250]), .Z(n1275) );
  IV U250 ( .A(B[251]), .Z(n1276) );
  IV U251 ( .A(B[252]), .Z(n1277) );
  IV U252 ( .A(B[253]), .Z(n1278) );
  IV U253 ( .A(B[254]), .Z(n1279) );
  IV U254 ( .A(B[255]), .Z(n1280) );
  IV U255 ( .A(B[256]), .Z(n1281) );
  IV U256 ( .A(B[949]), .Z(n1974) );
  IV U257 ( .A(B[257]), .Z(n1282) );
  IV U258 ( .A(B[258]), .Z(n1283) );
  IV U259 ( .A(B[259]), .Z(n1284) );
  IV U260 ( .A(B[260]), .Z(n1285) );
  IV U261 ( .A(B[261]), .Z(n1286) );
  IV U262 ( .A(B[262]), .Z(n1287) );
  IV U263 ( .A(B[263]), .Z(n1288) );
  IV U264 ( .A(B[264]), .Z(n1289) );
  IV U265 ( .A(B[265]), .Z(n1290) );
  IV U266 ( .A(B[266]), .Z(n1291) );
  IV U267 ( .A(B[950]), .Z(n1975) );
  IV U268 ( .A(B[267]), .Z(n1292) );
  IV U269 ( .A(B[268]), .Z(n1293) );
  IV U270 ( .A(B[269]), .Z(n1294) );
  IV U271 ( .A(B[270]), .Z(n1295) );
  IV U272 ( .A(B[271]), .Z(n1296) );
  IV U273 ( .A(B[272]), .Z(n1297) );
  IV U274 ( .A(B[273]), .Z(n1298) );
  IV U275 ( .A(B[274]), .Z(n1299) );
  IV U276 ( .A(B[275]), .Z(n1300) );
  IV U277 ( .A(B[276]), .Z(n1301) );
  IV U278 ( .A(B[951]), .Z(n1976) );
  IV U279 ( .A(B[277]), .Z(n1302) );
  IV U280 ( .A(B[278]), .Z(n1303) );
  IV U281 ( .A(B[279]), .Z(n1304) );
  IV U282 ( .A(B[280]), .Z(n1305) );
  IV U283 ( .A(B[281]), .Z(n1306) );
  IV U284 ( .A(B[282]), .Z(n1307) );
  IV U285 ( .A(B[283]), .Z(n1308) );
  IV U286 ( .A(B[284]), .Z(n1309) );
  IV U287 ( .A(B[285]), .Z(n1310) );
  IV U288 ( .A(B[286]), .Z(n1311) );
  IV U289 ( .A(B[952]), .Z(n1977) );
  IV U290 ( .A(B[287]), .Z(n1312) );
  IV U291 ( .A(B[288]), .Z(n1313) );
  IV U292 ( .A(B[289]), .Z(n1314) );
  IV U293 ( .A(B[290]), .Z(n1315) );
  IV U294 ( .A(B[291]), .Z(n1316) );
  IV U295 ( .A(B[292]), .Z(n1317) );
  IV U296 ( .A(B[293]), .Z(n1318) );
  IV U297 ( .A(B[294]), .Z(n1319) );
  IV U298 ( .A(B[295]), .Z(n1320) );
  IV U299 ( .A(B[296]), .Z(n1321) );
  IV U300 ( .A(B[953]), .Z(n1978) );
  IV U301 ( .A(B[297]), .Z(n1322) );
  IV U302 ( .A(B[298]), .Z(n1323) );
  IV U303 ( .A(B[299]), .Z(n1324) );
  IV U304 ( .A(B[300]), .Z(n1325) );
  IV U305 ( .A(B[301]), .Z(n1326) );
  IV U306 ( .A(B[302]), .Z(n1327) );
  IV U307 ( .A(B[303]), .Z(n1328) );
  IV U308 ( .A(B[304]), .Z(n1329) );
  IV U309 ( .A(B[305]), .Z(n1330) );
  IV U310 ( .A(B[306]), .Z(n1331) );
  IV U311 ( .A(B[954]), .Z(n1979) );
  IV U312 ( .A(B[307]), .Z(n1332) );
  IV U313 ( .A(B[308]), .Z(n1333) );
  IV U314 ( .A(B[309]), .Z(n1334) );
  IV U315 ( .A(B[310]), .Z(n1335) );
  IV U316 ( .A(B[311]), .Z(n1336) );
  IV U317 ( .A(B[312]), .Z(n1337) );
  IV U318 ( .A(B[313]), .Z(n1338) );
  IV U319 ( .A(B[314]), .Z(n1339) );
  IV U320 ( .A(B[315]), .Z(n1340) );
  IV U321 ( .A(B[316]), .Z(n1341) );
  IV U322 ( .A(B[955]), .Z(n1980) );
  IV U323 ( .A(B[317]), .Z(n1342) );
  IV U324 ( .A(B[318]), .Z(n1343) );
  IV U325 ( .A(B[319]), .Z(n1344) );
  IV U326 ( .A(B[320]), .Z(n1345) );
  IV U327 ( .A(B[321]), .Z(n1346) );
  IV U328 ( .A(B[322]), .Z(n1347) );
  IV U329 ( .A(B[323]), .Z(n1348) );
  IV U330 ( .A(B[324]), .Z(n1349) );
  IV U331 ( .A(B[325]), .Z(n1350) );
  IV U332 ( .A(B[326]), .Z(n1351) );
  IV U333 ( .A(B[956]), .Z(n1981) );
  IV U334 ( .A(B[1019]), .Z(n2044) );
  IV U335 ( .A(B[327]), .Z(n1352) );
  IV U336 ( .A(B[328]), .Z(n1353) );
  IV U337 ( .A(B[329]), .Z(n1354) );
  IV U338 ( .A(B[330]), .Z(n1355) );
  IV U339 ( .A(B[331]), .Z(n1356) );
  IV U340 ( .A(B[332]), .Z(n1357) );
  IV U341 ( .A(B[333]), .Z(n1358) );
  IV U342 ( .A(B[334]), .Z(n1359) );
  IV U343 ( .A(B[335]), .Z(n1360) );
  IV U344 ( .A(B[336]), .Z(n1361) );
  IV U345 ( .A(B[957]), .Z(n1982) );
  IV U346 ( .A(B[337]), .Z(n1362) );
  IV U347 ( .A(B[338]), .Z(n1363) );
  IV U348 ( .A(B[339]), .Z(n1364) );
  IV U349 ( .A(B[340]), .Z(n1365) );
  IV U350 ( .A(B[341]), .Z(n1366) );
  IV U351 ( .A(B[342]), .Z(n1367) );
  IV U352 ( .A(B[343]), .Z(n1368) );
  IV U353 ( .A(B[344]), .Z(n1369) );
  IV U354 ( .A(B[345]), .Z(n1370) );
  IV U355 ( .A(B[346]), .Z(n1371) );
  IV U356 ( .A(B[958]), .Z(n1983) );
  IV U357 ( .A(B[347]), .Z(n1372) );
  IV U358 ( .A(B[348]), .Z(n1373) );
  IV U359 ( .A(B[349]), .Z(n1374) );
  IV U360 ( .A(B[350]), .Z(n1375) );
  IV U361 ( .A(B[351]), .Z(n1376) );
  IV U362 ( .A(B[352]), .Z(n1377) );
  IV U363 ( .A(B[353]), .Z(n1378) );
  IV U364 ( .A(B[354]), .Z(n1379) );
  IV U365 ( .A(B[355]), .Z(n1380) );
  IV U366 ( .A(B[356]), .Z(n1381) );
  IV U367 ( .A(B[959]), .Z(n1984) );
  IV U368 ( .A(B[357]), .Z(n1382) );
  IV U369 ( .A(B[358]), .Z(n1383) );
  IV U370 ( .A(B[359]), .Z(n1384) );
  IV U371 ( .A(B[360]), .Z(n1385) );
  IV U372 ( .A(B[361]), .Z(n1386) );
  IV U373 ( .A(B[362]), .Z(n1387) );
  IV U374 ( .A(B[363]), .Z(n1388) );
  IV U375 ( .A(B[364]), .Z(n1389) );
  IV U376 ( .A(B[365]), .Z(n1390) );
  IV U377 ( .A(B[366]), .Z(n1391) );
  IV U378 ( .A(B[960]), .Z(n1985) );
  IV U379 ( .A(B[367]), .Z(n1392) );
  IV U380 ( .A(B[368]), .Z(n1393) );
  IV U381 ( .A(B[369]), .Z(n1394) );
  IV U382 ( .A(B[370]), .Z(n1395) );
  IV U383 ( .A(B[371]), .Z(n1396) );
  IV U384 ( .A(B[372]), .Z(n1397) );
  IV U385 ( .A(B[373]), .Z(n1398) );
  IV U386 ( .A(B[374]), .Z(n1399) );
  IV U387 ( .A(B[375]), .Z(n1400) );
  IV U388 ( .A(B[376]), .Z(n1401) );
  IV U389 ( .A(B[961]), .Z(n1986) );
  IV U390 ( .A(B[377]), .Z(n1402) );
  IV U391 ( .A(B[378]), .Z(n1403) );
  IV U392 ( .A(B[379]), .Z(n1404) );
  IV U393 ( .A(B[380]), .Z(n1405) );
  IV U394 ( .A(B[381]), .Z(n1406) );
  IV U395 ( .A(B[382]), .Z(n1407) );
  IV U396 ( .A(B[383]), .Z(n1408) );
  IV U397 ( .A(B[384]), .Z(n1409) );
  IV U398 ( .A(B[385]), .Z(n1410) );
  IV U399 ( .A(B[386]), .Z(n1411) );
  IV U400 ( .A(B[962]), .Z(n1987) );
  IV U401 ( .A(B[387]), .Z(n1412) );
  IV U402 ( .A(B[388]), .Z(n1413) );
  IV U403 ( .A(B[389]), .Z(n1414) );
  IV U404 ( .A(B[390]), .Z(n1415) );
  IV U405 ( .A(B[391]), .Z(n1416) );
  IV U406 ( .A(B[392]), .Z(n1417) );
  IV U407 ( .A(B[393]), .Z(n1418) );
  IV U408 ( .A(B[394]), .Z(n1419) );
  IV U409 ( .A(B[395]), .Z(n1420) );
  IV U410 ( .A(B[396]), .Z(n1421) );
  IV U411 ( .A(B[963]), .Z(n1988) );
  IV U412 ( .A(B[397]), .Z(n1422) );
  IV U413 ( .A(B[398]), .Z(n1423) );
  IV U414 ( .A(B[399]), .Z(n1424) );
  IV U415 ( .A(B[400]), .Z(n1425) );
  IV U416 ( .A(B[401]), .Z(n1426) );
  IV U417 ( .A(B[402]), .Z(n1427) );
  IV U418 ( .A(B[403]), .Z(n1428) );
  IV U419 ( .A(B[404]), .Z(n1429) );
  IV U420 ( .A(B[405]), .Z(n1430) );
  IV U421 ( .A(B[406]), .Z(n1431) );
  IV U422 ( .A(B[964]), .Z(n1989) );
  IV U423 ( .A(B[407]), .Z(n1432) );
  IV U424 ( .A(B[408]), .Z(n1433) );
  IV U425 ( .A(B[409]), .Z(n1434) );
  IV U426 ( .A(B[410]), .Z(n1435) );
  IV U427 ( .A(B[411]), .Z(n1436) );
  IV U428 ( .A(B[412]), .Z(n1437) );
  IV U429 ( .A(B[413]), .Z(n1438) );
  IV U430 ( .A(B[414]), .Z(n1439) );
  IV U431 ( .A(B[415]), .Z(n1440) );
  IV U432 ( .A(B[416]), .Z(n1441) );
  IV U433 ( .A(B[965]), .Z(n1990) );
  IV U434 ( .A(B[417]), .Z(n1442) );
  IV U435 ( .A(B[418]), .Z(n1443) );
  IV U436 ( .A(B[419]), .Z(n1444) );
  IV U437 ( .A(B[420]), .Z(n1445) );
  IV U438 ( .A(B[421]), .Z(n1446) );
  IV U439 ( .A(B[422]), .Z(n1447) );
  IV U440 ( .A(B[423]), .Z(n1448) );
  IV U441 ( .A(B[424]), .Z(n1449) );
  IV U442 ( .A(B[425]), .Z(n1450) );
  IV U443 ( .A(B[426]), .Z(n1451) );
  IV U444 ( .A(B[966]), .Z(n1991) );
  IV U445 ( .A(B[1020]), .Z(n2045) );
  IV U446 ( .A(B[427]), .Z(n1452) );
  IV U447 ( .A(B[428]), .Z(n1453) );
  IV U448 ( .A(B[429]), .Z(n1454) );
  IV U449 ( .A(B[430]), .Z(n1455) );
  IV U450 ( .A(B[431]), .Z(n1456) );
  IV U451 ( .A(B[432]), .Z(n1457) );
  IV U452 ( .A(B[433]), .Z(n1458) );
  IV U453 ( .A(B[434]), .Z(n1459) );
  IV U454 ( .A(B[435]), .Z(n1460) );
  IV U455 ( .A(B[436]), .Z(n1461) );
  IV U456 ( .A(B[967]), .Z(n1992) );
  IV U457 ( .A(B[437]), .Z(n1462) );
  IV U458 ( .A(B[438]), .Z(n1463) );
  IV U459 ( .A(B[439]), .Z(n1464) );
  IV U460 ( .A(B[440]), .Z(n1465) );
  IV U461 ( .A(B[441]), .Z(n1466) );
  IV U462 ( .A(B[442]), .Z(n1467) );
  IV U463 ( .A(B[443]), .Z(n1468) );
  IV U464 ( .A(B[444]), .Z(n1469) );
  IV U465 ( .A(B[445]), .Z(n1470) );
  IV U466 ( .A(B[446]), .Z(n1471) );
  IV U467 ( .A(B[968]), .Z(n1993) );
  IV U468 ( .A(B[447]), .Z(n1472) );
  IV U469 ( .A(B[448]), .Z(n1473) );
  IV U470 ( .A(B[449]), .Z(n1474) );
  IV U471 ( .A(B[450]), .Z(n1475) );
  IV U472 ( .A(B[451]), .Z(n1476) );
  IV U473 ( .A(B[452]), .Z(n1477) );
  IV U474 ( .A(B[453]), .Z(n1478) );
  IV U475 ( .A(B[454]), .Z(n1479) );
  IV U476 ( .A(B[455]), .Z(n1480) );
  IV U477 ( .A(B[456]), .Z(n1481) );
  IV U478 ( .A(B[969]), .Z(n1994) );
  IV U479 ( .A(B[457]), .Z(n1482) );
  IV U480 ( .A(B[458]), .Z(n1483) );
  IV U481 ( .A(B[459]), .Z(n1484) );
  IV U482 ( .A(B[460]), .Z(n1485) );
  IV U483 ( .A(B[461]), .Z(n1486) );
  IV U484 ( .A(B[462]), .Z(n1487) );
  IV U485 ( .A(B[463]), .Z(n1488) );
  IV U486 ( .A(B[464]), .Z(n1489) );
  IV U487 ( .A(B[465]), .Z(n1490) );
  IV U488 ( .A(B[466]), .Z(n1491) );
  IV U489 ( .A(B[970]), .Z(n1995) );
  IV U490 ( .A(B[467]), .Z(n1492) );
  IV U491 ( .A(B[468]), .Z(n1493) );
  IV U492 ( .A(B[469]), .Z(n1494) );
  IV U493 ( .A(B[470]), .Z(n1495) );
  IV U494 ( .A(B[471]), .Z(n1496) );
  IV U495 ( .A(B[472]), .Z(n1497) );
  IV U496 ( .A(B[473]), .Z(n1498) );
  IV U497 ( .A(B[474]), .Z(n1499) );
  IV U498 ( .A(B[475]), .Z(n1500) );
  IV U499 ( .A(B[476]), .Z(n1501) );
  IV U500 ( .A(B[971]), .Z(n1996) );
  IV U501 ( .A(B[477]), .Z(n1502) );
  IV U502 ( .A(B[478]), .Z(n1503) );
  IV U503 ( .A(B[479]), .Z(n1504) );
  IV U504 ( .A(B[480]), .Z(n1505) );
  IV U505 ( .A(B[481]), .Z(n1506) );
  IV U506 ( .A(B[482]), .Z(n1507) );
  IV U507 ( .A(B[483]), .Z(n1508) );
  IV U508 ( .A(B[484]), .Z(n1509) );
  IV U509 ( .A(B[485]), .Z(n1510) );
  IV U510 ( .A(B[486]), .Z(n1511) );
  IV U511 ( .A(B[972]), .Z(n1997) );
  IV U512 ( .A(B[487]), .Z(n1512) );
  IV U513 ( .A(B[488]), .Z(n1513) );
  IV U514 ( .A(B[489]), .Z(n1514) );
  IV U515 ( .A(B[490]), .Z(n1515) );
  IV U516 ( .A(B[491]), .Z(n1516) );
  IV U517 ( .A(B[492]), .Z(n1517) );
  IV U518 ( .A(B[493]), .Z(n1518) );
  IV U519 ( .A(B[494]), .Z(n1519) );
  IV U520 ( .A(B[495]), .Z(n1520) );
  IV U521 ( .A(B[496]), .Z(n1521) );
  IV U522 ( .A(B[973]), .Z(n1998) );
  IV U523 ( .A(B[497]), .Z(n1522) );
  IV U524 ( .A(B[498]), .Z(n1523) );
  IV U525 ( .A(B[499]), .Z(n1524) );
  IV U526 ( .A(B[500]), .Z(n1525) );
  IV U527 ( .A(B[501]), .Z(n1526) );
  IV U528 ( .A(B[502]), .Z(n1527) );
  IV U529 ( .A(B[503]), .Z(n1528) );
  IV U530 ( .A(B[504]), .Z(n1529) );
  IV U531 ( .A(B[505]), .Z(n1530) );
  IV U532 ( .A(B[506]), .Z(n1531) );
  IV U533 ( .A(B[974]), .Z(n1999) );
  IV U534 ( .A(B[507]), .Z(n1532) );
  IV U535 ( .A(B[508]), .Z(n1533) );
  IV U536 ( .A(B[509]), .Z(n1534) );
  IV U537 ( .A(B[510]), .Z(n1535) );
  IV U538 ( .A(B[511]), .Z(n1536) );
  IV U539 ( .A(B[512]), .Z(n1537) );
  IV U540 ( .A(B[513]), .Z(n1538) );
  IV U541 ( .A(B[514]), .Z(n1539) );
  IV U542 ( .A(B[515]), .Z(n1540) );
  IV U543 ( .A(B[516]), .Z(n1541) );
  IV U544 ( .A(B[975]), .Z(n2000) );
  IV U545 ( .A(B[517]), .Z(n1542) );
  IV U546 ( .A(B[518]), .Z(n1543) );
  IV U547 ( .A(B[519]), .Z(n1544) );
  IV U548 ( .A(B[520]), .Z(n1545) );
  IV U549 ( .A(B[521]), .Z(n1546) );
  IV U550 ( .A(B[522]), .Z(n1547) );
  IV U551 ( .A(B[523]), .Z(n1548) );
  IV U552 ( .A(B[524]), .Z(n1549) );
  IV U553 ( .A(B[525]), .Z(n1550) );
  IV U554 ( .A(B[526]), .Z(n1551) );
  IV U555 ( .A(B[976]), .Z(n2001) );
  IV U556 ( .A(B[1021]), .Z(n2046) );
  IV U557 ( .A(B[527]), .Z(n1552) );
  IV U558 ( .A(B[528]), .Z(n1553) );
  IV U559 ( .A(B[529]), .Z(n1554) );
  IV U560 ( .A(B[530]), .Z(n1555) );
  IV U561 ( .A(B[531]), .Z(n1556) );
  IV U562 ( .A(B[532]), .Z(n1557) );
  IV U563 ( .A(B[533]), .Z(n1558) );
  IV U564 ( .A(B[534]), .Z(n1559) );
  IV U565 ( .A(B[535]), .Z(n1560) );
  IV U566 ( .A(B[536]), .Z(n1561) );
  IV U567 ( .A(B[977]), .Z(n2002) );
  IV U568 ( .A(B[537]), .Z(n1562) );
  IV U569 ( .A(B[538]), .Z(n1563) );
  IV U570 ( .A(B[539]), .Z(n1564) );
  IV U571 ( .A(B[540]), .Z(n1565) );
  IV U572 ( .A(B[541]), .Z(n1566) );
  IV U573 ( .A(B[542]), .Z(n1567) );
  IV U574 ( .A(B[543]), .Z(n1568) );
  IV U575 ( .A(B[544]), .Z(n1569) );
  IV U576 ( .A(B[545]), .Z(n1570) );
  IV U577 ( .A(B[546]), .Z(n1571) );
  IV U578 ( .A(B[978]), .Z(n2003) );
  IV U579 ( .A(B[547]), .Z(n1572) );
  IV U580 ( .A(B[548]), .Z(n1573) );
  IV U581 ( .A(B[549]), .Z(n1574) );
  IV U582 ( .A(B[550]), .Z(n1575) );
  IV U583 ( .A(B[551]), .Z(n1576) );
  IV U584 ( .A(B[552]), .Z(n1577) );
  IV U585 ( .A(B[553]), .Z(n1578) );
  IV U586 ( .A(B[554]), .Z(n1579) );
  IV U587 ( .A(B[555]), .Z(n1580) );
  IV U588 ( .A(B[556]), .Z(n1581) );
  IV U589 ( .A(B[979]), .Z(n2004) );
  IV U590 ( .A(B[557]), .Z(n1582) );
  IV U591 ( .A(B[558]), .Z(n1583) );
  IV U592 ( .A(B[559]), .Z(n1584) );
  IV U593 ( .A(B[560]), .Z(n1585) );
  IV U594 ( .A(B[561]), .Z(n1586) );
  IV U595 ( .A(B[562]), .Z(n1587) );
  IV U596 ( .A(B[563]), .Z(n1588) );
  IV U597 ( .A(B[564]), .Z(n1589) );
  IV U598 ( .A(B[565]), .Z(n1590) );
  IV U599 ( .A(B[566]), .Z(n1591) );
  IV U600 ( .A(B[980]), .Z(n2005) );
  IV U601 ( .A(B[567]), .Z(n1592) );
  IV U602 ( .A(B[568]), .Z(n1593) );
  IV U603 ( .A(B[569]), .Z(n1594) );
  IV U604 ( .A(B[570]), .Z(n1595) );
  IV U605 ( .A(B[571]), .Z(n1596) );
  IV U606 ( .A(B[572]), .Z(n1597) );
  IV U607 ( .A(B[573]), .Z(n1598) );
  IV U608 ( .A(B[574]), .Z(n1599) );
  IV U609 ( .A(B[575]), .Z(n1600) );
  IV U610 ( .A(B[576]), .Z(n1601) );
  IV U611 ( .A(B[981]), .Z(n2006) );
  IV U612 ( .A(B[577]), .Z(n1602) );
  IV U613 ( .A(B[578]), .Z(n1603) );
  IV U614 ( .A(B[579]), .Z(n1604) );
  IV U615 ( .A(B[580]), .Z(n1605) );
  IV U616 ( .A(B[581]), .Z(n1606) );
  IV U617 ( .A(B[582]), .Z(n1607) );
  IV U618 ( .A(B[583]), .Z(n1608) );
  IV U619 ( .A(B[584]), .Z(n1609) );
  IV U620 ( .A(B[585]), .Z(n1610) );
  IV U621 ( .A(B[586]), .Z(n1611) );
  IV U622 ( .A(B[982]), .Z(n2007) );
  IV U623 ( .A(B[587]), .Z(n1612) );
  IV U624 ( .A(B[588]), .Z(n1613) );
  IV U625 ( .A(B[589]), .Z(n1614) );
  IV U626 ( .A(B[590]), .Z(n1615) );
  IV U627 ( .A(B[591]), .Z(n1616) );
  IV U628 ( .A(B[592]), .Z(n1617) );
  IV U629 ( .A(B[593]), .Z(n1618) );
  IV U630 ( .A(B[594]), .Z(n1619) );
  IV U631 ( .A(B[595]), .Z(n1620) );
  IV U632 ( .A(B[596]), .Z(n1621) );
  IV U633 ( .A(B[983]), .Z(n2008) );
  IV U634 ( .A(B[597]), .Z(n1622) );
  IV U635 ( .A(B[598]), .Z(n1623) );
  IV U636 ( .A(B[599]), .Z(n1624) );
  IV U637 ( .A(B[600]), .Z(n1625) );
  IV U638 ( .A(B[601]), .Z(n1626) );
  IV U639 ( .A(B[602]), .Z(n1627) );
  IV U640 ( .A(B[603]), .Z(n1628) );
  IV U641 ( .A(B[604]), .Z(n1629) );
  IV U642 ( .A(B[605]), .Z(n1630) );
  IV U643 ( .A(B[606]), .Z(n1631) );
  IV U644 ( .A(B[984]), .Z(n2009) );
  IV U645 ( .A(B[607]), .Z(n1632) );
  IV U646 ( .A(B[608]), .Z(n1633) );
  IV U647 ( .A(B[609]), .Z(n1634) );
  IV U648 ( .A(B[610]), .Z(n1635) );
  IV U649 ( .A(B[611]), .Z(n1636) );
  IV U650 ( .A(B[612]), .Z(n1637) );
  IV U651 ( .A(B[613]), .Z(n1638) );
  IV U652 ( .A(B[614]), .Z(n1639) );
  IV U653 ( .A(B[615]), .Z(n1640) );
  IV U654 ( .A(B[616]), .Z(n1641) );
  IV U655 ( .A(B[985]), .Z(n2010) );
  IV U656 ( .A(B[617]), .Z(n1642) );
  IV U657 ( .A(B[618]), .Z(n1643) );
  IV U658 ( .A(B[619]), .Z(n1644) );
  IV U659 ( .A(B[620]), .Z(n1645) );
  IV U660 ( .A(B[621]), .Z(n1646) );
  IV U661 ( .A(B[622]), .Z(n1647) );
  IV U662 ( .A(B[623]), .Z(n1648) );
  IV U663 ( .A(B[624]), .Z(n1649) );
  IV U664 ( .A(B[625]), .Z(n1650) );
  IV U665 ( .A(B[626]), .Z(n1651) );
  IV U666 ( .A(B[986]), .Z(n2011) );
  IV U667 ( .A(B[1022]), .Z(n2047) );
  IV U668 ( .A(B[627]), .Z(n1652) );
  IV U669 ( .A(B[628]), .Z(n1653) );
  IV U670 ( .A(B[629]), .Z(n1654) );
  IV U671 ( .A(B[630]), .Z(n1655) );
  IV U672 ( .A(B[631]), .Z(n1656) );
  IV U673 ( .A(B[632]), .Z(n1657) );
  IV U674 ( .A(B[633]), .Z(n1658) );
  IV U675 ( .A(B[634]), .Z(n1659) );
  IV U676 ( .A(B[635]), .Z(n1660) );
  IV U677 ( .A(B[636]), .Z(n1661) );
  IV U678 ( .A(B[987]), .Z(n2012) );
  IV U679 ( .A(B[637]), .Z(n1662) );
  IV U680 ( .A(B[638]), .Z(n1663) );
  IV U681 ( .A(B[639]), .Z(n1664) );
  IV U682 ( .A(B[640]), .Z(n1665) );
  IV U683 ( .A(B[641]), .Z(n1666) );
  IV U684 ( .A(B[642]), .Z(n1667) );
  IV U685 ( .A(B[643]), .Z(n1668) );
  IV U686 ( .A(B[644]), .Z(n1669) );
  IV U687 ( .A(B[645]), .Z(n1670) );
  IV U688 ( .A(B[646]), .Z(n1671) );
  IV U689 ( .A(B[988]), .Z(n2013) );
  IV U690 ( .A(B[647]), .Z(n1672) );
  IV U691 ( .A(B[648]), .Z(n1673) );
  IV U692 ( .A(B[649]), .Z(n1674) );
  IV U693 ( .A(B[650]), .Z(n1675) );
  IV U694 ( .A(B[651]), .Z(n1676) );
  IV U695 ( .A(B[652]), .Z(n1677) );
  IV U696 ( .A(B[653]), .Z(n1678) );
  IV U697 ( .A(B[654]), .Z(n1679) );
  IV U698 ( .A(B[655]), .Z(n1680) );
  IV U699 ( .A(B[656]), .Z(n1681) );
  IV U700 ( .A(B[989]), .Z(n2014) );
  IV U701 ( .A(B[657]), .Z(n1682) );
  IV U702 ( .A(B[658]), .Z(n1683) );
  IV U703 ( .A(B[659]), .Z(n1684) );
  IV U704 ( .A(B[660]), .Z(n1685) );
  IV U705 ( .A(B[661]), .Z(n1686) );
  IV U706 ( .A(B[662]), .Z(n1687) );
  IV U707 ( .A(B[663]), .Z(n1688) );
  IV U708 ( .A(B[664]), .Z(n1689) );
  IV U709 ( .A(B[665]), .Z(n1690) );
  IV U710 ( .A(B[666]), .Z(n1691) );
  IV U711 ( .A(B[990]), .Z(n2015) );
  IV U712 ( .A(B[667]), .Z(n1692) );
  IV U713 ( .A(B[668]), .Z(n1693) );
  IV U714 ( .A(B[669]), .Z(n1694) );
  IV U715 ( .A(B[670]), .Z(n1695) );
  IV U716 ( .A(B[671]), .Z(n1696) );
  IV U717 ( .A(B[672]), .Z(n1697) );
  IV U718 ( .A(B[673]), .Z(n1698) );
  IV U719 ( .A(B[674]), .Z(n1699) );
  IV U720 ( .A(B[675]), .Z(n1700) );
  IV U721 ( .A(B[676]), .Z(n1701) );
  IV U722 ( .A(B[991]), .Z(n2016) );
  IV U723 ( .A(B[677]), .Z(n1702) );
  IV U724 ( .A(B[678]), .Z(n1703) );
  IV U725 ( .A(B[679]), .Z(n1704) );
  IV U726 ( .A(B[680]), .Z(n1705) );
  IV U727 ( .A(B[681]), .Z(n1706) );
  IV U728 ( .A(B[682]), .Z(n1707) );
  IV U729 ( .A(B[683]), .Z(n1708) );
  IV U730 ( .A(B[684]), .Z(n1709) );
  IV U731 ( .A(B[685]), .Z(n1710) );
  IV U732 ( .A(B[686]), .Z(n1711) );
  IV U733 ( .A(B[992]), .Z(n2017) );
  IV U734 ( .A(B[687]), .Z(n1712) );
  IV U735 ( .A(B[688]), .Z(n1713) );
  IV U736 ( .A(B[689]), .Z(n1714) );
  IV U737 ( .A(B[690]), .Z(n1715) );
  IV U738 ( .A(B[691]), .Z(n1716) );
  IV U739 ( .A(B[692]), .Z(n1717) );
  IV U740 ( .A(B[693]), .Z(n1718) );
  IV U741 ( .A(B[694]), .Z(n1719) );
  IV U742 ( .A(B[695]), .Z(n1720) );
  IV U743 ( .A(B[696]), .Z(n1721) );
  IV U744 ( .A(B[993]), .Z(n2018) );
  IV U745 ( .A(B[697]), .Z(n1722) );
  IV U746 ( .A(B[698]), .Z(n1723) );
  IV U747 ( .A(B[699]), .Z(n1724) );
  IV U748 ( .A(B[700]), .Z(n1725) );
  IV U749 ( .A(B[701]), .Z(n1726) );
  IV U750 ( .A(B[702]), .Z(n1727) );
  IV U751 ( .A(B[703]), .Z(n1728) );
  IV U752 ( .A(B[704]), .Z(n1729) );
  IV U753 ( .A(B[705]), .Z(n1730) );
  IV U754 ( .A(B[706]), .Z(n1731) );
  IV U755 ( .A(B[994]), .Z(n2019) );
  IV U756 ( .A(B[707]), .Z(n1732) );
  IV U757 ( .A(B[708]), .Z(n1733) );
  IV U758 ( .A(B[709]), .Z(n1734) );
  IV U759 ( .A(B[710]), .Z(n1735) );
  IV U760 ( .A(B[711]), .Z(n1736) );
  IV U761 ( .A(B[712]), .Z(n1737) );
  IV U762 ( .A(B[713]), .Z(n1738) );
  IV U763 ( .A(B[714]), .Z(n1739) );
  IV U764 ( .A(B[715]), .Z(n1740) );
  IV U765 ( .A(B[716]), .Z(n1741) );
  IV U766 ( .A(B[995]), .Z(n2020) );
  IV U767 ( .A(B[717]), .Z(n1742) );
  IV U768 ( .A(B[718]), .Z(n1743) );
  IV U769 ( .A(B[719]), .Z(n1744) );
  IV U770 ( .A(B[720]), .Z(n1745) );
  IV U771 ( .A(B[721]), .Z(n1746) );
  IV U772 ( .A(B[722]), .Z(n1747) );
  IV U773 ( .A(B[723]), .Z(n1748) );
  IV U774 ( .A(B[724]), .Z(n1749) );
  IV U775 ( .A(B[725]), .Z(n1750) );
  IV U776 ( .A(B[726]), .Z(n1751) );
  IV U777 ( .A(B[996]), .Z(n2021) );
  IV U778 ( .A(B[1023]), .Z(n2048) );
  IV U779 ( .A(B[727]), .Z(n1752) );
  IV U780 ( .A(B[728]), .Z(n1753) );
  IV U781 ( .A(B[729]), .Z(n1754) );
  IV U782 ( .A(B[730]), .Z(n1755) );
  IV U783 ( .A(B[731]), .Z(n1756) );
  IV U784 ( .A(B[732]), .Z(n1757) );
  IV U785 ( .A(B[733]), .Z(n1758) );
  IV U786 ( .A(B[734]), .Z(n1759) );
  IV U787 ( .A(B[735]), .Z(n1760) );
  IV U788 ( .A(B[736]), .Z(n1761) );
  IV U789 ( .A(B[997]), .Z(n2022) );
  IV U790 ( .A(B[737]), .Z(n1762) );
  IV U791 ( .A(B[738]), .Z(n1763) );
  IV U792 ( .A(B[739]), .Z(n1764) );
  IV U793 ( .A(B[740]), .Z(n1765) );
  IV U794 ( .A(B[741]), .Z(n1766) );
  IV U795 ( .A(B[742]), .Z(n1767) );
  IV U796 ( .A(B[743]), .Z(n1768) );
  IV U797 ( .A(B[744]), .Z(n1769) );
  IV U798 ( .A(B[745]), .Z(n1770) );
  IV U799 ( .A(B[746]), .Z(n1771) );
  IV U800 ( .A(B[998]), .Z(n2023) );
  IV U801 ( .A(B[747]), .Z(n1772) );
  IV U802 ( .A(B[748]), .Z(n1773) );
  IV U803 ( .A(B[749]), .Z(n1774) );
  IV U804 ( .A(B[750]), .Z(n1775) );
  IV U805 ( .A(B[751]), .Z(n1776) );
  IV U806 ( .A(B[752]), .Z(n1777) );
  IV U807 ( .A(B[753]), .Z(n1778) );
  IV U808 ( .A(B[754]), .Z(n1779) );
  IV U809 ( .A(B[755]), .Z(n1780) );
  IV U810 ( .A(B[756]), .Z(n1781) );
  IV U811 ( .A(B[999]), .Z(n2024) );
  IV U812 ( .A(B[757]), .Z(n1782) );
  IV U813 ( .A(B[758]), .Z(n1783) );
  IV U814 ( .A(B[759]), .Z(n1784) );
  IV U815 ( .A(B[760]), .Z(n1785) );
  IV U816 ( .A(B[761]), .Z(n1786) );
  IV U817 ( .A(B[762]), .Z(n1787) );
  IV U818 ( .A(B[763]), .Z(n1788) );
  IV U819 ( .A(B[764]), .Z(n1789) );
  IV U820 ( .A(B[765]), .Z(n1790) );
  IV U821 ( .A(B[766]), .Z(n1791) );
  IV U822 ( .A(B[1000]), .Z(n2025) );
  IV U823 ( .A(B[767]), .Z(n1792) );
  IV U824 ( .A(B[768]), .Z(n1793) );
  IV U825 ( .A(B[769]), .Z(n1794) );
  IV U826 ( .A(B[770]), .Z(n1795) );
  IV U827 ( .A(B[771]), .Z(n1796) );
  IV U828 ( .A(B[772]), .Z(n1797) );
  IV U829 ( .A(B[773]), .Z(n1798) );
  IV U830 ( .A(B[774]), .Z(n1799) );
  IV U831 ( .A(B[775]), .Z(n1800) );
  IV U832 ( .A(B[776]), .Z(n1801) );
  IV U833 ( .A(B[1001]), .Z(n2026) );
  IV U834 ( .A(B[777]), .Z(n1802) );
  IV U835 ( .A(B[778]), .Z(n1803) );
  IV U836 ( .A(B[779]), .Z(n1804) );
  IV U837 ( .A(B[780]), .Z(n1805) );
  IV U838 ( .A(B[781]), .Z(n1806) );
  IV U839 ( .A(B[782]), .Z(n1807) );
  IV U840 ( .A(B[783]), .Z(n1808) );
  IV U841 ( .A(B[784]), .Z(n1809) );
  IV U842 ( .A(B[785]), .Z(n1810) );
  IV U843 ( .A(B[786]), .Z(n1811) );
  IV U844 ( .A(B[1002]), .Z(n2027) );
  IV U845 ( .A(B[787]), .Z(n1812) );
  IV U846 ( .A(B[788]), .Z(n1813) );
  IV U847 ( .A(B[789]), .Z(n1814) );
  IV U848 ( .A(B[790]), .Z(n1815) );
  IV U849 ( .A(B[791]), .Z(n1816) );
  IV U850 ( .A(B[792]), .Z(n1817) );
  IV U851 ( .A(B[793]), .Z(n1818) );
  IV U852 ( .A(B[794]), .Z(n1819) );
  IV U853 ( .A(B[795]), .Z(n1820) );
  IV U854 ( .A(B[796]), .Z(n1821) );
  IV U855 ( .A(B[1003]), .Z(n2028) );
  IV U856 ( .A(B[797]), .Z(n1822) );
  IV U857 ( .A(B[798]), .Z(n1823) );
  IV U858 ( .A(B[799]), .Z(n1824) );
  IV U859 ( .A(B[800]), .Z(n1825) );
  IV U860 ( .A(B[801]), .Z(n1826) );
  IV U861 ( .A(B[802]), .Z(n1827) );
  IV U862 ( .A(B[803]), .Z(n1828) );
  IV U863 ( .A(B[804]), .Z(n1829) );
  IV U864 ( .A(B[805]), .Z(n1830) );
  IV U865 ( .A(B[806]), .Z(n1831) );
  IV U866 ( .A(B[1004]), .Z(n2029) );
  IV U867 ( .A(B[807]), .Z(n1832) );
  IV U868 ( .A(B[808]), .Z(n1833) );
  IV U869 ( .A(B[809]), .Z(n1834) );
  IV U870 ( .A(B[810]), .Z(n1835) );
  IV U871 ( .A(B[811]), .Z(n1836) );
  IV U872 ( .A(B[812]), .Z(n1837) );
  IV U873 ( .A(B[813]), .Z(n1838) );
  IV U874 ( .A(B[814]), .Z(n1839) );
  IV U875 ( .A(B[815]), .Z(n1840) );
  IV U876 ( .A(B[816]), .Z(n1841) );
  IV U877 ( .A(B[1005]), .Z(n2030) );
  IV U878 ( .A(B[817]), .Z(n1842) );
  IV U879 ( .A(B[818]), .Z(n1843) );
  IV U880 ( .A(B[819]), .Z(n1844) );
  IV U881 ( .A(B[820]), .Z(n1845) );
  IV U882 ( .A(B[821]), .Z(n1846) );
  IV U883 ( .A(B[822]), .Z(n1847) );
  IV U884 ( .A(B[823]), .Z(n1848) );
  IV U885 ( .A(B[824]), .Z(n1849) );
  IV U886 ( .A(B[825]), .Z(n1850) );
  IV U887 ( .A(B[826]), .Z(n1851) );
  IV U888 ( .A(B[1006]), .Z(n2031) );
  IV U889 ( .A(B[827]), .Z(n1852) );
  IV U890 ( .A(B[828]), .Z(n1853) );
  IV U891 ( .A(B[829]), .Z(n1854) );
  IV U892 ( .A(B[830]), .Z(n1855) );
  IV U893 ( .A(B[831]), .Z(n1856) );
  IV U894 ( .A(B[832]), .Z(n1857) );
  IV U895 ( .A(B[833]), .Z(n1858) );
  IV U896 ( .A(B[834]), .Z(n1859) );
  IV U897 ( .A(B[835]), .Z(n1860) );
  IV U898 ( .A(B[836]), .Z(n1861) );
  IV U899 ( .A(B[1007]), .Z(n2032) );
  IV U900 ( .A(B[837]), .Z(n1862) );
  IV U901 ( .A(B[838]), .Z(n1863) );
  IV U902 ( .A(B[839]), .Z(n1864) );
  IV U903 ( .A(B[840]), .Z(n1865) );
  IV U904 ( .A(B[841]), .Z(n1866) );
  IV U905 ( .A(B[842]), .Z(n1867) );
  IV U906 ( .A(B[843]), .Z(n1868) );
  IV U907 ( .A(B[844]), .Z(n1869) );
  IV U908 ( .A(B[845]), .Z(n1870) );
  IV U909 ( .A(B[846]), .Z(n1871) );
  IV U910 ( .A(B[1008]), .Z(n2033) );
  IV U911 ( .A(B[847]), .Z(n1872) );
  IV U912 ( .A(B[848]), .Z(n1873) );
  IV U913 ( .A(B[849]), .Z(n1874) );
  IV U914 ( .A(B[850]), .Z(n1875) );
  IV U915 ( .A(B[851]), .Z(n1876) );
  IV U916 ( .A(B[852]), .Z(n1877) );
  IV U917 ( .A(B[853]), .Z(n1878) );
  IV U918 ( .A(B[854]), .Z(n1879) );
  IV U919 ( .A(B[855]), .Z(n1880) );
  IV U920 ( .A(B[856]), .Z(n1881) );
  IV U921 ( .A(B[1009]), .Z(n2034) );
  IV U922 ( .A(B[857]), .Z(n1882) );
  IV U923 ( .A(B[858]), .Z(n1883) );
  IV U924 ( .A(B[859]), .Z(n1884) );
  IV U925 ( .A(B[860]), .Z(n1885) );
  IV U926 ( .A(B[861]), .Z(n1886) );
  IV U927 ( .A(B[862]), .Z(n1887) );
  IV U928 ( .A(B[863]), .Z(n1888) );
  IV U929 ( .A(B[864]), .Z(n1889) );
  IV U930 ( .A(B[865]), .Z(n1890) );
  IV U931 ( .A(B[866]), .Z(n1891) );
  IV U932 ( .A(B[1010]), .Z(n2035) );
  IV U933 ( .A(B[867]), .Z(n1892) );
  IV U934 ( .A(B[868]), .Z(n1893) );
  IV U935 ( .A(B[869]), .Z(n1894) );
  IV U936 ( .A(B[870]), .Z(n1895) );
  IV U937 ( .A(B[871]), .Z(n1896) );
  IV U938 ( .A(B[872]), .Z(n1897) );
  IV U939 ( .A(B[873]), .Z(n1898) );
  IV U940 ( .A(B[874]), .Z(n1899) );
  IV U941 ( .A(B[875]), .Z(n1900) );
  IV U942 ( .A(B[876]), .Z(n1901) );
  IV U943 ( .A(B[1011]), .Z(n2036) );
  IV U944 ( .A(B[877]), .Z(n1902) );
  IV U945 ( .A(B[878]), .Z(n1903) );
  IV U946 ( .A(B[879]), .Z(n1904) );
  IV U947 ( .A(B[880]), .Z(n1905) );
  IV U948 ( .A(B[881]), .Z(n1906) );
  IV U949 ( .A(B[882]), .Z(n1907) );
  IV U950 ( .A(B[883]), .Z(n1908) );
  IV U951 ( .A(B[884]), .Z(n1909) );
  IV U952 ( .A(B[885]), .Z(n1910) );
  IV U953 ( .A(B[886]), .Z(n1911) );
  IV U954 ( .A(B[1012]), .Z(n2037) );
  IV U955 ( .A(B[887]), .Z(n1912) );
  IV U956 ( .A(B[888]), .Z(n1913) );
  IV U957 ( .A(B[889]), .Z(n1914) );
  IV U958 ( .A(B[890]), .Z(n1915) );
  IV U959 ( .A(B[891]), .Z(n1916) );
  IV U960 ( .A(B[892]), .Z(n1917) );
  IV U961 ( .A(B[893]), .Z(n1918) );
  IV U962 ( .A(B[894]), .Z(n1919) );
  IV U963 ( .A(B[895]), .Z(n1920) );
  IV U964 ( .A(B[896]), .Z(n1921) );
  IV U965 ( .A(B[1013]), .Z(n2038) );
  IV U966 ( .A(B[897]), .Z(n1922) );
  IV U967 ( .A(B[898]), .Z(n1923) );
  IV U968 ( .A(B[899]), .Z(n1924) );
  IV U969 ( .A(B[900]), .Z(n1925) );
  IV U970 ( .A(B[901]), .Z(n1926) );
  IV U971 ( .A(B[902]), .Z(n1927) );
  IV U972 ( .A(B[903]), .Z(n1928) );
  IV U973 ( .A(B[904]), .Z(n1929) );
  IV U974 ( .A(B[905]), .Z(n1930) );
  IV U975 ( .A(B[906]), .Z(n1931) );
  IV U976 ( .A(B[1014]), .Z(n2039) );
  IV U977 ( .A(B[907]), .Z(n1932) );
  IV U978 ( .A(B[908]), .Z(n1933) );
  IV U979 ( .A(B[909]), .Z(n1934) );
  IV U980 ( .A(B[910]), .Z(n1935) );
  IV U981 ( .A(B[911]), .Z(n1936) );
  IV U982 ( .A(B[912]), .Z(n1937) );
  IV U983 ( .A(B[913]), .Z(n1938) );
  IV U984 ( .A(B[914]), .Z(n1939) );
  IV U985 ( .A(B[915]), .Z(n1940) );
  IV U986 ( .A(B[916]), .Z(n1941) );
  IV U987 ( .A(B[1015]), .Z(n2040) );
  IV U988 ( .A(B[917]), .Z(n1942) );
  IV U989 ( .A(B[918]), .Z(n1943) );
  IV U990 ( .A(B[919]), .Z(n1944) );
  IV U991 ( .A(B[920]), .Z(n1945) );
  IV U992 ( .A(B[921]), .Z(n1946) );
  IV U993 ( .A(B[922]), .Z(n1947) );
  IV U994 ( .A(B[923]), .Z(n1948) );
  IV U995 ( .A(B[0]), .Z(n2) );
  IV U996 ( .A(B[1]), .Z(n1026) );
  IV U997 ( .A(B[2]), .Z(n1027) );
  IV U998 ( .A(B[3]), .Z(n1028) );
  IV U999 ( .A(B[4]), .Z(n1029) );
  IV U1000 ( .A(B[5]), .Z(n1030) );
  IV U1001 ( .A(B[6]), .Z(n1031) );
  IV U1002 ( .A(B[924]), .Z(n1949) );
  IV U1003 ( .A(B[7]), .Z(n1032) );
  IV U1004 ( .A(B[8]), .Z(n1033) );
  IV U1005 ( .A(B[9]), .Z(n1034) );
  IV U1006 ( .A(B[10]), .Z(n1035) );
  IV U1007 ( .A(B[11]), .Z(n1036) );
  IV U1008 ( .A(B[12]), .Z(n1037) );
  IV U1009 ( .A(B[13]), .Z(n1038) );
  IV U1010 ( .A(B[14]), .Z(n1039) );
  IV U1011 ( .A(B[15]), .Z(n1040) );
  IV U1012 ( .A(B[16]), .Z(n1041) );
  IV U1013 ( .A(B[925]), .Z(n1950) );
  IV U1014 ( .A(B[17]), .Z(n1042) );
  IV U1015 ( .A(B[18]), .Z(n1043) );
  IV U1016 ( .A(B[19]), .Z(n1044) );
  IV U1017 ( .A(B[20]), .Z(n1045) );
  IV U1018 ( .A(B[21]), .Z(n1046) );
  IV U1019 ( .A(B[22]), .Z(n1047) );
  IV U1020 ( .A(B[23]), .Z(n1048) );
  IV U1021 ( .A(B[24]), .Z(n1049) );
  IV U1022 ( .A(B[25]), .Z(n1050) );
  IV U1023 ( .A(B[26]), .Z(n1051) );
  IV U1024 ( .A(B[926]), .Z(n1951) );
  IV U1025 ( .A(B[1016]), .Z(n2041) );
endmodule


module modmult_step_N1024 ( xregN_1, y, n, zin, zout );
  input [1023:0] y;
  input [1023:0] n;
  input [1025:0] zin;
  output [1025:0] zout;
  input xregN_1;
  wire   c1, c2, n1;
  wire   [1025:0] w1;
  wire   [1025:0] w2;
  wire   [1025:0] w3;
  wire   [1025:0] z2;
  wire   [1025:0] z3;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6;

  MUX_N1026_0 MUX_1 ( .A({1'b0, 1'b0, y}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .S(xregN_1), .O({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, w1[1023:0]}) );
  MUX_N1026_2 MUX_2 ( .A({1'b0, 1'b0, n}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .S(c1), .O({SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        w2[1023:0]}) );
  MUX_N1026_1 MUX_3 ( .A({1'b0, 1'b0, n}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .S(n1), .O({SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        w3[1023:0]}) );
  ADD_N1026 ADD_1 ( .A({zin[1024:0], 1'b0}), .B({1'b0, 1'b0, w1[1023:0]}), 
        .CI(1'b0), .S(z2) );
  COMP_N1026_0 COMP_1 ( .A(z2), .B({1'b0, 1'b0, n}), .O(c1) );
  SUB_N1026_0 SUB_1 ( .A(z2), .B({1'b0, 1'b0, w2[1023:0]}), .S(z3) );
  COMP_N1026_1 COMP_2 ( .A({1'b0, 1'b0, n}), .B(z3), .O(c2) );
  SUB_N1026_1 SUB_2 ( .A({1'b0, z3[1024:0]}), .B({1'b0, 1'b0, w3[1023:0]}), 
        .S({SYNOPSYS_UNCONNECTED__6, zout[1024:0]}) );
  IV U2 ( .A(c2), .Z(n1) );
endmodule


module modmult_N1024_CC1024 ( clk, rst, start, x, y, n, o );
  input [1023:0] x;
  input [1023:0] y;
  input [1023:0] n;
  output [1023:0] o;
  input clk, rst, start;
  wire   \zout[0][1024] , \zin[0][1024] , \zin[0][1023] , \zin[0][1022] ,
         \zin[0][1021] , \zin[0][1020] , \zin[0][1019] , \zin[0][1018] ,
         \zin[0][1017] , \zin[0][1016] , \zin[0][1015] , \zin[0][1014] ,
         \zin[0][1013] , \zin[0][1012] , \zin[0][1011] , \zin[0][1010] ,
         \zin[0][1009] , \zin[0][1008] , \zin[0][1007] , \zin[0][1006] ,
         \zin[0][1005] , \zin[0][1004] , \zin[0][1003] , \zin[0][1002] ,
         \zin[0][1001] , \zin[0][1000] , \zin[0][999] , \zin[0][998] ,
         \zin[0][997] , \zin[0][996] , \zin[0][995] , \zin[0][994] ,
         \zin[0][993] , \zin[0][992] , \zin[0][991] , \zin[0][990] ,
         \zin[0][989] , \zin[0][988] , \zin[0][987] , \zin[0][986] ,
         \zin[0][985] , \zin[0][984] , \zin[0][983] , \zin[0][982] ,
         \zin[0][981] , \zin[0][980] , \zin[0][979] , \zin[0][978] ,
         \zin[0][977] , \zin[0][976] , \zin[0][975] , \zin[0][974] ,
         \zin[0][973] , \zin[0][972] , \zin[0][971] , \zin[0][970] ,
         \zin[0][969] , \zin[0][968] , \zin[0][967] , \zin[0][966] ,
         \zin[0][965] , \zin[0][964] , \zin[0][963] , \zin[0][962] ,
         \zin[0][961] , \zin[0][960] , \zin[0][959] , \zin[0][958] ,
         \zin[0][957] , \zin[0][956] , \zin[0][955] , \zin[0][954] ,
         \zin[0][953] , \zin[0][952] , \zin[0][951] , \zin[0][950] ,
         \zin[0][949] , \zin[0][948] , \zin[0][947] , \zin[0][946] ,
         \zin[0][945] , \zin[0][944] , \zin[0][943] , \zin[0][942] ,
         \zin[0][941] , \zin[0][940] , \zin[0][939] , \zin[0][938] ,
         \zin[0][937] , \zin[0][936] , \zin[0][935] , \zin[0][934] ,
         \zin[0][933] , \zin[0][932] , \zin[0][931] , \zin[0][930] ,
         \zin[0][929] , \zin[0][928] , \zin[0][927] , \zin[0][926] ,
         \zin[0][925] , \zin[0][924] , \zin[0][923] , \zin[0][922] ,
         \zin[0][921] , \zin[0][920] , \zin[0][919] , \zin[0][918] ,
         \zin[0][917] , \zin[0][916] , \zin[0][915] , \zin[0][914] ,
         \zin[0][913] , \zin[0][912] , \zin[0][911] , \zin[0][910] ,
         \zin[0][909] , \zin[0][908] , \zin[0][907] , \zin[0][906] ,
         \zin[0][905] , \zin[0][904] , \zin[0][903] , \zin[0][902] ,
         \zin[0][901] , \zin[0][900] , \zin[0][899] , \zin[0][898] ,
         \zin[0][897] , \zin[0][896] , \zin[0][895] , \zin[0][894] ,
         \zin[0][893] , \zin[0][892] , \zin[0][891] , \zin[0][890] ,
         \zin[0][889] , \zin[0][888] , \zin[0][887] , \zin[0][886] ,
         \zin[0][885] , \zin[0][884] , \zin[0][883] , \zin[0][882] ,
         \zin[0][881] , \zin[0][880] , \zin[0][879] , \zin[0][878] ,
         \zin[0][877] , \zin[0][876] , \zin[0][875] , \zin[0][874] ,
         \zin[0][873] , \zin[0][872] , \zin[0][871] , \zin[0][870] ,
         \zin[0][869] , \zin[0][868] , \zin[0][867] , \zin[0][866] ,
         \zin[0][865] , \zin[0][864] , \zin[0][863] , \zin[0][862] ,
         \zin[0][861] , \zin[0][860] , \zin[0][859] , \zin[0][858] ,
         \zin[0][857] , \zin[0][856] , \zin[0][855] , \zin[0][854] ,
         \zin[0][853] , \zin[0][852] , \zin[0][851] , \zin[0][850] ,
         \zin[0][849] , \zin[0][848] , \zin[0][847] , \zin[0][846] ,
         \zin[0][845] , \zin[0][844] , \zin[0][843] , \zin[0][842] ,
         \zin[0][841] , \zin[0][840] , \zin[0][839] , \zin[0][838] ,
         \zin[0][837] , \zin[0][836] , \zin[0][835] , \zin[0][834] ,
         \zin[0][833] , \zin[0][832] , \zin[0][831] , \zin[0][830] ,
         \zin[0][829] , \zin[0][828] , \zin[0][827] , \zin[0][826] ,
         \zin[0][825] , \zin[0][824] , \zin[0][823] , \zin[0][822] ,
         \zin[0][821] , \zin[0][820] , \zin[0][819] , \zin[0][818] ,
         \zin[0][817] , \zin[0][816] , \zin[0][815] , \zin[0][814] ,
         \zin[0][813] , \zin[0][812] , \zin[0][811] , \zin[0][810] ,
         \zin[0][809] , \zin[0][808] , \zin[0][807] , \zin[0][806] ,
         \zin[0][805] , \zin[0][804] , \zin[0][803] , \zin[0][802] ,
         \zin[0][801] , \zin[0][800] , \zin[0][799] , \zin[0][798] ,
         \zin[0][797] , \zin[0][796] , \zin[0][795] , \zin[0][794] ,
         \zin[0][793] , \zin[0][792] , \zin[0][791] , \zin[0][790] ,
         \zin[0][789] , \zin[0][788] , \zin[0][787] , \zin[0][786] ,
         \zin[0][785] , \zin[0][784] , \zin[0][783] , \zin[0][782] ,
         \zin[0][781] , \zin[0][780] , \zin[0][779] , \zin[0][778] ,
         \zin[0][777] , \zin[0][776] , \zin[0][775] , \zin[0][774] ,
         \zin[0][773] , \zin[0][772] , \zin[0][771] , \zin[0][770] ,
         \zin[0][769] , \zin[0][768] , \zin[0][767] , \zin[0][766] ,
         \zin[0][765] , \zin[0][764] , \zin[0][763] , \zin[0][762] ,
         \zin[0][761] , \zin[0][760] , \zin[0][759] , \zin[0][758] ,
         \zin[0][757] , \zin[0][756] , \zin[0][755] , \zin[0][754] ,
         \zin[0][753] , \zin[0][752] , \zin[0][751] , \zin[0][750] ,
         \zin[0][749] , \zin[0][748] , \zin[0][747] , \zin[0][746] ,
         \zin[0][745] , \zin[0][744] , \zin[0][743] , \zin[0][742] ,
         \zin[0][741] , \zin[0][740] , \zin[0][739] , \zin[0][738] ,
         \zin[0][737] , \zin[0][736] , \zin[0][735] , \zin[0][734] ,
         \zin[0][733] , \zin[0][732] , \zin[0][731] , \zin[0][730] ,
         \zin[0][729] , \zin[0][728] , \zin[0][727] , \zin[0][726] ,
         \zin[0][725] , \zin[0][724] , \zin[0][723] , \zin[0][722] ,
         \zin[0][721] , \zin[0][720] , \zin[0][719] , \zin[0][718] ,
         \zin[0][717] , \zin[0][716] , \zin[0][715] , \zin[0][714] ,
         \zin[0][713] , \zin[0][712] , \zin[0][711] , \zin[0][710] ,
         \zin[0][709] , \zin[0][708] , \zin[0][707] , \zin[0][706] ,
         \zin[0][705] , \zin[0][704] , \zin[0][703] , \zin[0][702] ,
         \zin[0][701] , \zin[0][700] , \zin[0][699] , \zin[0][698] ,
         \zin[0][697] , \zin[0][696] , \zin[0][695] , \zin[0][694] ,
         \zin[0][693] , \zin[0][692] , \zin[0][691] , \zin[0][690] ,
         \zin[0][689] , \zin[0][688] , \zin[0][687] , \zin[0][686] ,
         \zin[0][685] , \zin[0][684] , \zin[0][683] , \zin[0][682] ,
         \zin[0][681] , \zin[0][680] , \zin[0][679] , \zin[0][678] ,
         \zin[0][677] , \zin[0][676] , \zin[0][675] , \zin[0][674] ,
         \zin[0][673] , \zin[0][672] , \zin[0][671] , \zin[0][670] ,
         \zin[0][669] , \zin[0][668] , \zin[0][667] , \zin[0][666] ,
         \zin[0][665] , \zin[0][664] , \zin[0][663] , \zin[0][662] ,
         \zin[0][661] , \zin[0][660] , \zin[0][659] , \zin[0][658] ,
         \zin[0][657] , \zin[0][656] , \zin[0][655] , \zin[0][654] ,
         \zin[0][653] , \zin[0][652] , \zin[0][651] , \zin[0][650] ,
         \zin[0][649] , \zin[0][648] , \zin[0][647] , \zin[0][646] ,
         \zin[0][645] , \zin[0][644] , \zin[0][643] , \zin[0][642] ,
         \zin[0][641] , \zin[0][640] , \zin[0][639] , \zin[0][638] ,
         \zin[0][637] , \zin[0][636] , \zin[0][635] , \zin[0][634] ,
         \zin[0][633] , \zin[0][632] , \zin[0][631] , \zin[0][630] ,
         \zin[0][629] , \zin[0][628] , \zin[0][627] , \zin[0][626] ,
         \zin[0][625] , \zin[0][624] , \zin[0][623] , \zin[0][622] ,
         \zin[0][621] , \zin[0][620] , \zin[0][619] , \zin[0][618] ,
         \zin[0][617] , \zin[0][616] , \zin[0][615] , \zin[0][614] ,
         \zin[0][613] , \zin[0][612] , \zin[0][611] , \zin[0][610] ,
         \zin[0][609] , \zin[0][608] , \zin[0][607] , \zin[0][606] ,
         \zin[0][605] , \zin[0][604] , \zin[0][603] , \zin[0][602] ,
         \zin[0][601] , \zin[0][600] , \zin[0][599] , \zin[0][598] ,
         \zin[0][597] , \zin[0][596] , \zin[0][595] , \zin[0][594] ,
         \zin[0][593] , \zin[0][592] , \zin[0][591] , \zin[0][590] ,
         \zin[0][589] , \zin[0][588] , \zin[0][587] , \zin[0][586] ,
         \zin[0][585] , \zin[0][584] , \zin[0][583] , \zin[0][582] ,
         \zin[0][581] , \zin[0][580] , \zin[0][579] , \zin[0][578] ,
         \zin[0][577] , \zin[0][576] , \zin[0][575] , \zin[0][574] ,
         \zin[0][573] , \zin[0][572] , \zin[0][571] , \zin[0][570] ,
         \zin[0][569] , \zin[0][568] , \zin[0][567] , \zin[0][566] ,
         \zin[0][565] , \zin[0][564] , \zin[0][563] , \zin[0][562] ,
         \zin[0][561] , \zin[0][560] , \zin[0][559] , \zin[0][558] ,
         \zin[0][557] , \zin[0][556] , \zin[0][555] , \zin[0][554] ,
         \zin[0][553] , \zin[0][552] , \zin[0][551] , \zin[0][550] ,
         \zin[0][549] , \zin[0][548] , \zin[0][547] , \zin[0][546] ,
         \zin[0][545] , \zin[0][544] , \zin[0][543] , \zin[0][542] ,
         \zin[0][541] , \zin[0][540] , \zin[0][539] , \zin[0][538] ,
         \zin[0][537] , \zin[0][536] , \zin[0][535] , \zin[0][534] ,
         \zin[0][533] , \zin[0][532] , \zin[0][531] , \zin[0][530] ,
         \zin[0][529] , \zin[0][528] , \zin[0][527] , \zin[0][526] ,
         \zin[0][525] , \zin[0][524] , \zin[0][523] , \zin[0][522] ,
         \zin[0][521] , \zin[0][520] , \zin[0][519] , \zin[0][518] ,
         \zin[0][517] , \zin[0][516] , \zin[0][515] , \zin[0][514] ,
         \zin[0][513] , \zin[0][512] , \zin[0][511] , \zin[0][510] ,
         \zin[0][509] , \zin[0][508] , \zin[0][507] , \zin[0][506] ,
         \zin[0][505] , \zin[0][504] , \zin[0][503] , \zin[0][502] ,
         \zin[0][501] , \zin[0][500] , \zin[0][499] , \zin[0][498] ,
         \zin[0][497] , \zin[0][496] , \zin[0][495] , \zin[0][494] ,
         \zin[0][493] , \zin[0][492] , \zin[0][491] , \zin[0][490] ,
         \zin[0][489] , \zin[0][488] , \zin[0][487] , \zin[0][486] ,
         \zin[0][485] , \zin[0][484] , \zin[0][483] , \zin[0][482] ,
         \zin[0][481] , \zin[0][480] , \zin[0][479] , \zin[0][478] ,
         \zin[0][477] , \zin[0][476] , \zin[0][475] , \zin[0][474] ,
         \zin[0][473] , \zin[0][472] , \zin[0][471] , \zin[0][470] ,
         \zin[0][469] , \zin[0][468] , \zin[0][467] , \zin[0][466] ,
         \zin[0][465] , \zin[0][464] , \zin[0][463] , \zin[0][462] ,
         \zin[0][461] , \zin[0][460] , \zin[0][459] , \zin[0][458] ,
         \zin[0][457] , \zin[0][456] , \zin[0][455] , \zin[0][454] ,
         \zin[0][453] , \zin[0][452] , \zin[0][451] , \zin[0][450] ,
         \zin[0][449] , \zin[0][448] , \zin[0][447] , \zin[0][446] ,
         \zin[0][445] , \zin[0][444] , \zin[0][443] , \zin[0][442] ,
         \zin[0][441] , \zin[0][440] , \zin[0][439] , \zin[0][438] ,
         \zin[0][437] , \zin[0][436] , \zin[0][435] , \zin[0][434] ,
         \zin[0][433] , \zin[0][432] , \zin[0][431] , \zin[0][430] ,
         \zin[0][429] , \zin[0][428] , \zin[0][427] , \zin[0][426] ,
         \zin[0][425] , \zin[0][424] , \zin[0][423] , \zin[0][422] ,
         \zin[0][421] , \zin[0][420] , \zin[0][419] , \zin[0][418] ,
         \zin[0][417] , \zin[0][416] , \zin[0][415] , \zin[0][414] ,
         \zin[0][413] , \zin[0][412] , \zin[0][411] , \zin[0][410] ,
         \zin[0][409] , \zin[0][408] , \zin[0][407] , \zin[0][406] ,
         \zin[0][405] , \zin[0][404] , \zin[0][403] , \zin[0][402] ,
         \zin[0][401] , \zin[0][400] , \zin[0][399] , \zin[0][398] ,
         \zin[0][397] , \zin[0][396] , \zin[0][395] , \zin[0][394] ,
         \zin[0][393] , \zin[0][392] , \zin[0][391] , \zin[0][390] ,
         \zin[0][389] , \zin[0][388] , \zin[0][387] , \zin[0][386] ,
         \zin[0][385] , \zin[0][384] , \zin[0][383] , \zin[0][382] ,
         \zin[0][381] , \zin[0][380] , \zin[0][379] , \zin[0][378] ,
         \zin[0][377] , \zin[0][376] , \zin[0][375] , \zin[0][374] ,
         \zin[0][373] , \zin[0][372] , \zin[0][371] , \zin[0][370] ,
         \zin[0][369] , \zin[0][368] , \zin[0][367] , \zin[0][366] ,
         \zin[0][365] , \zin[0][364] , \zin[0][363] , \zin[0][362] ,
         \zin[0][361] , \zin[0][360] , \zin[0][359] , \zin[0][358] ,
         \zin[0][357] , \zin[0][356] , \zin[0][355] , \zin[0][354] ,
         \zin[0][353] , \zin[0][352] , \zin[0][351] , \zin[0][350] ,
         \zin[0][349] , \zin[0][348] , \zin[0][347] , \zin[0][346] ,
         \zin[0][345] , \zin[0][344] , \zin[0][343] , \zin[0][342] ,
         \zin[0][341] , \zin[0][340] , \zin[0][339] , \zin[0][338] ,
         \zin[0][337] , \zin[0][336] , \zin[0][335] , \zin[0][334] ,
         \zin[0][333] , \zin[0][332] , \zin[0][331] , \zin[0][330] ,
         \zin[0][329] , \zin[0][328] , \zin[0][327] , \zin[0][326] ,
         \zin[0][325] , \zin[0][324] , \zin[0][323] , \zin[0][322] ,
         \zin[0][321] , \zin[0][320] , \zin[0][319] , \zin[0][318] ,
         \zin[0][317] , \zin[0][316] , \zin[0][315] , \zin[0][314] ,
         \zin[0][313] , \zin[0][312] , \zin[0][311] , \zin[0][310] ,
         \zin[0][309] , \zin[0][308] , \zin[0][307] , \zin[0][306] ,
         \zin[0][305] , \zin[0][304] , \zin[0][303] , \zin[0][302] ,
         \zin[0][301] , \zin[0][300] , \zin[0][299] , \zin[0][298] ,
         \zin[0][297] , \zin[0][296] , \zin[0][295] , \zin[0][294] ,
         \zin[0][293] , \zin[0][292] , \zin[0][291] , \zin[0][290] ,
         \zin[0][289] , \zin[0][288] , \zin[0][287] , \zin[0][286] ,
         \zin[0][285] , \zin[0][284] , \zin[0][283] , \zin[0][282] ,
         \zin[0][281] , \zin[0][280] , \zin[0][279] , \zin[0][278] ,
         \zin[0][277] , \zin[0][276] , \zin[0][275] , \zin[0][274] ,
         \zin[0][273] , \zin[0][272] , \zin[0][271] , \zin[0][270] ,
         \zin[0][269] , \zin[0][268] , \zin[0][267] , \zin[0][266] ,
         \zin[0][265] , \zin[0][264] , \zin[0][263] , \zin[0][262] ,
         \zin[0][261] , \zin[0][260] , \zin[0][259] , \zin[0][258] ,
         \zin[0][257] , \zin[0][256] , \zin[0][255] , \zin[0][254] ,
         \zin[0][253] , \zin[0][252] , \zin[0][251] , \zin[0][250] ,
         \zin[0][249] , \zin[0][248] , \zin[0][247] , \zin[0][246] ,
         \zin[0][245] , \zin[0][244] , \zin[0][243] , \zin[0][242] ,
         \zin[0][241] , \zin[0][240] , \zin[0][239] , \zin[0][238] ,
         \zin[0][237] , \zin[0][236] , \zin[0][235] , \zin[0][234] ,
         \zin[0][233] , \zin[0][232] , \zin[0][231] , \zin[0][230] ,
         \zin[0][229] , \zin[0][228] , \zin[0][227] , \zin[0][226] ,
         \zin[0][225] , \zin[0][224] , \zin[0][223] , \zin[0][222] ,
         \zin[0][221] , \zin[0][220] , \zin[0][219] , \zin[0][218] ,
         \zin[0][217] , \zin[0][216] , \zin[0][215] , \zin[0][214] ,
         \zin[0][213] , \zin[0][212] , \zin[0][211] , \zin[0][210] ,
         \zin[0][209] , \zin[0][208] , \zin[0][207] , \zin[0][206] ,
         \zin[0][205] , \zin[0][204] , \zin[0][203] , \zin[0][202] ,
         \zin[0][201] , \zin[0][200] , \zin[0][199] , \zin[0][198] ,
         \zin[0][197] , \zin[0][196] , \zin[0][195] , \zin[0][194] ,
         \zin[0][193] , \zin[0][192] , \zin[0][191] , \zin[0][190] ,
         \zin[0][189] , \zin[0][188] , \zin[0][187] , \zin[0][186] ,
         \zin[0][185] , \zin[0][184] , \zin[0][183] , \zin[0][182] ,
         \zin[0][181] , \zin[0][180] , \zin[0][179] , \zin[0][178] ,
         \zin[0][177] , \zin[0][176] , \zin[0][175] , \zin[0][174] ,
         \zin[0][173] , \zin[0][172] , \zin[0][171] , \zin[0][170] ,
         \zin[0][169] , \zin[0][168] , \zin[0][167] , \zin[0][166] ,
         \zin[0][165] , \zin[0][164] , \zin[0][163] , \zin[0][162] ,
         \zin[0][161] , \zin[0][160] , \zin[0][159] , \zin[0][158] ,
         \zin[0][157] , \zin[0][156] , \zin[0][155] , \zin[0][154] ,
         \zin[0][153] , \zin[0][152] , \zin[0][151] , \zin[0][150] ,
         \zin[0][149] , \zin[0][148] , \zin[0][147] , \zin[0][146] ,
         \zin[0][145] , \zin[0][144] , \zin[0][143] , \zin[0][142] ,
         \zin[0][141] , \zin[0][140] , \zin[0][139] , \zin[0][138] ,
         \zin[0][137] , \zin[0][136] , \zin[0][135] , \zin[0][134] ,
         \zin[0][133] , \zin[0][132] , \zin[0][131] , \zin[0][130] ,
         \zin[0][129] , \zin[0][128] , \zin[0][127] , \zin[0][126] ,
         \zin[0][125] , \zin[0][124] , \zin[0][123] , \zin[0][122] ,
         \zin[0][121] , \zin[0][120] , \zin[0][119] , \zin[0][118] ,
         \zin[0][117] , \zin[0][116] , \zin[0][115] , \zin[0][114] ,
         \zin[0][113] , \zin[0][112] , \zin[0][111] , \zin[0][110] ,
         \zin[0][109] , \zin[0][108] , \zin[0][107] , \zin[0][106] ,
         \zin[0][105] , \zin[0][104] , \zin[0][103] , \zin[0][102] ,
         \zin[0][101] , \zin[0][100] , \zin[0][99] , \zin[0][98] ,
         \zin[0][97] , \zin[0][96] , \zin[0][95] , \zin[0][94] , \zin[0][93] ,
         \zin[0][92] , \zin[0][91] , \zin[0][90] , \zin[0][89] , \zin[0][88] ,
         \zin[0][87] , \zin[0][86] , \zin[0][85] , \zin[0][84] , \zin[0][83] ,
         \zin[0][82] , \zin[0][81] , \zin[0][80] , \zin[0][79] , \zin[0][78] ,
         \zin[0][77] , \zin[0][76] , \zin[0][75] , \zin[0][74] , \zin[0][73] ,
         \zin[0][72] , \zin[0][71] , \zin[0][70] , \zin[0][69] , \zin[0][68] ,
         \zin[0][67] , \zin[0][66] , \zin[0][65] , \zin[0][64] , \zin[0][63] ,
         \zin[0][62] , \zin[0][61] , \zin[0][60] , \zin[0][59] , \zin[0][58] ,
         \zin[0][57] , \zin[0][56] , \zin[0][55] , \zin[0][54] , \zin[0][53] ,
         \zin[0][52] , \zin[0][51] , \zin[0][50] , \zin[0][49] , \zin[0][48] ,
         \zin[0][47] , \zin[0][46] , \zin[0][45] , \zin[0][44] , \zin[0][43] ,
         \zin[0][42] , \zin[0][41] , \zin[0][40] , \zin[0][39] , \zin[0][38] ,
         \zin[0][37] , \zin[0][36] , \zin[0][35] , \zin[0][34] , \zin[0][33] ,
         \zin[0][32] , \zin[0][31] , \zin[0][30] , \zin[0][29] , \zin[0][28] ,
         \zin[0][27] , \zin[0][26] , \zin[0][25] , \zin[0][24] , \zin[0][23] ,
         \zin[0][22] , \zin[0][21] , \zin[0][20] , \zin[0][19] , \zin[0][18] ,
         \zin[0][17] , \zin[0][16] , \zin[0][15] , \zin[0][14] , \zin[0][13] ,
         \zin[0][12] , \zin[0][11] , \zin[0][10] , \zin[0][9] , \zin[0][8] ,
         \zin[0][7] , \zin[0][6] , \zin[0][5] , \zin[0][4] , \zin[0][3] ,
         \zin[0][2] , \zin[0][1] , \zin[0][0] ;
  wire   [1023:0] xin;
  wire   SYNOPSYS_UNCONNECTED__0;

  modmult_step_N1024 \MODMULT_STEP[0].modmult_step_  ( .xregN_1(xin[1023]), 
        .y(y), .n(n), .zin({1'b0, \zin[0][1024] , \zin[0][1023] , 
        \zin[0][1022] , \zin[0][1021] , \zin[0][1020] , \zin[0][1019] , 
        \zin[0][1018] , \zin[0][1017] , \zin[0][1016] , \zin[0][1015] , 
        \zin[0][1014] , \zin[0][1013] , \zin[0][1012] , \zin[0][1011] , 
        \zin[0][1010] , \zin[0][1009] , \zin[0][1008] , \zin[0][1007] , 
        \zin[0][1006] , \zin[0][1005] , \zin[0][1004] , \zin[0][1003] , 
        \zin[0][1002] , \zin[0][1001] , \zin[0][1000] , \zin[0][999] , 
        \zin[0][998] , \zin[0][997] , \zin[0][996] , \zin[0][995] , 
        \zin[0][994] , \zin[0][993] , \zin[0][992] , \zin[0][991] , 
        \zin[0][990] , \zin[0][989] , \zin[0][988] , \zin[0][987] , 
        \zin[0][986] , \zin[0][985] , \zin[0][984] , \zin[0][983] , 
        \zin[0][982] , \zin[0][981] , \zin[0][980] , \zin[0][979] , 
        \zin[0][978] , \zin[0][977] , \zin[0][976] , \zin[0][975] , 
        \zin[0][974] , \zin[0][973] , \zin[0][972] , \zin[0][971] , 
        \zin[0][970] , \zin[0][969] , \zin[0][968] , \zin[0][967] , 
        \zin[0][966] , \zin[0][965] , \zin[0][964] , \zin[0][963] , 
        \zin[0][962] , \zin[0][961] , \zin[0][960] , \zin[0][959] , 
        \zin[0][958] , \zin[0][957] , \zin[0][956] , \zin[0][955] , 
        \zin[0][954] , \zin[0][953] , \zin[0][952] , \zin[0][951] , 
        \zin[0][950] , \zin[0][949] , \zin[0][948] , \zin[0][947] , 
        \zin[0][946] , \zin[0][945] , \zin[0][944] , \zin[0][943] , 
        \zin[0][942] , \zin[0][941] , \zin[0][940] , \zin[0][939] , 
        \zin[0][938] , \zin[0][937] , \zin[0][936] , \zin[0][935] , 
        \zin[0][934] , \zin[0][933] , \zin[0][932] , \zin[0][931] , 
        \zin[0][930] , \zin[0][929] , \zin[0][928] , \zin[0][927] , 
        \zin[0][926] , \zin[0][925] , \zin[0][924] , \zin[0][923] , 
        \zin[0][922] , \zin[0][921] , \zin[0][920] , \zin[0][919] , 
        \zin[0][918] , \zin[0][917] , \zin[0][916] , \zin[0][915] , 
        \zin[0][914] , \zin[0][913] , \zin[0][912] , \zin[0][911] , 
        \zin[0][910] , \zin[0][909] , \zin[0][908] , \zin[0][907] , 
        \zin[0][906] , \zin[0][905] , \zin[0][904] , \zin[0][903] , 
        \zin[0][902] , \zin[0][901] , \zin[0][900] , \zin[0][899] , 
        \zin[0][898] , \zin[0][897] , \zin[0][896] , \zin[0][895] , 
        \zin[0][894] , \zin[0][893] , \zin[0][892] , \zin[0][891] , 
        \zin[0][890] , \zin[0][889] , \zin[0][888] , \zin[0][887] , 
        \zin[0][886] , \zin[0][885] , \zin[0][884] , \zin[0][883] , 
        \zin[0][882] , \zin[0][881] , \zin[0][880] , \zin[0][879] , 
        \zin[0][878] , \zin[0][877] , \zin[0][876] , \zin[0][875] , 
        \zin[0][874] , \zin[0][873] , \zin[0][872] , \zin[0][871] , 
        \zin[0][870] , \zin[0][869] , \zin[0][868] , \zin[0][867] , 
        \zin[0][866] , \zin[0][865] , \zin[0][864] , \zin[0][863] , 
        \zin[0][862] , \zin[0][861] , \zin[0][860] , \zin[0][859] , 
        \zin[0][858] , \zin[0][857] , \zin[0][856] , \zin[0][855] , 
        \zin[0][854] , \zin[0][853] , \zin[0][852] , \zin[0][851] , 
        \zin[0][850] , \zin[0][849] , \zin[0][848] , \zin[0][847] , 
        \zin[0][846] , \zin[0][845] , \zin[0][844] , \zin[0][843] , 
        \zin[0][842] , \zin[0][841] , \zin[0][840] , \zin[0][839] , 
        \zin[0][838] , \zin[0][837] , \zin[0][836] , \zin[0][835] , 
        \zin[0][834] , \zin[0][833] , \zin[0][832] , \zin[0][831] , 
        \zin[0][830] , \zin[0][829] , \zin[0][828] , \zin[0][827] , 
        \zin[0][826] , \zin[0][825] , \zin[0][824] , \zin[0][823] , 
        \zin[0][822] , \zin[0][821] , \zin[0][820] , \zin[0][819] , 
        \zin[0][818] , \zin[0][817] , \zin[0][816] , \zin[0][815] , 
        \zin[0][814] , \zin[0][813] , \zin[0][812] , \zin[0][811] , 
        \zin[0][810] , \zin[0][809] , \zin[0][808] , \zin[0][807] , 
        \zin[0][806] , \zin[0][805] , \zin[0][804] , \zin[0][803] , 
        \zin[0][802] , \zin[0][801] , \zin[0][800] , \zin[0][799] , 
        \zin[0][798] , \zin[0][797] , \zin[0][796] , \zin[0][795] , 
        \zin[0][794] , \zin[0][793] , \zin[0][792] , \zin[0][791] , 
        \zin[0][790] , \zin[0][789] , \zin[0][788] , \zin[0][787] , 
        \zin[0][786] , \zin[0][785] , \zin[0][784] , \zin[0][783] , 
        \zin[0][782] , \zin[0][781] , \zin[0][780] , \zin[0][779] , 
        \zin[0][778] , \zin[0][777] , \zin[0][776] , \zin[0][775] , 
        \zin[0][774] , \zin[0][773] , \zin[0][772] , \zin[0][771] , 
        \zin[0][770] , \zin[0][769] , \zin[0][768] , \zin[0][767] , 
        \zin[0][766] , \zin[0][765] , \zin[0][764] , \zin[0][763] , 
        \zin[0][762] , \zin[0][761] , \zin[0][760] , \zin[0][759] , 
        \zin[0][758] , \zin[0][757] , \zin[0][756] , \zin[0][755] , 
        \zin[0][754] , \zin[0][753] , \zin[0][752] , \zin[0][751] , 
        \zin[0][750] , \zin[0][749] , \zin[0][748] , \zin[0][747] , 
        \zin[0][746] , \zin[0][745] , \zin[0][744] , \zin[0][743] , 
        \zin[0][742] , \zin[0][741] , \zin[0][740] , \zin[0][739] , 
        \zin[0][738] , \zin[0][737] , \zin[0][736] , \zin[0][735] , 
        \zin[0][734] , \zin[0][733] , \zin[0][732] , \zin[0][731] , 
        \zin[0][730] , \zin[0][729] , \zin[0][728] , \zin[0][727] , 
        \zin[0][726] , \zin[0][725] , \zin[0][724] , \zin[0][723] , 
        \zin[0][722] , \zin[0][721] , \zin[0][720] , \zin[0][719] , 
        \zin[0][718] , \zin[0][717] , \zin[0][716] , \zin[0][715] , 
        \zin[0][714] , \zin[0][713] , \zin[0][712] , \zin[0][711] , 
        \zin[0][710] , \zin[0][709] , \zin[0][708] , \zin[0][707] , 
        \zin[0][706] , \zin[0][705] , \zin[0][704] , \zin[0][703] , 
        \zin[0][702] , \zin[0][701] , \zin[0][700] , \zin[0][699] , 
        \zin[0][698] , \zin[0][697] , \zin[0][696] , \zin[0][695] , 
        \zin[0][694] , \zin[0][693] , \zin[0][692] , \zin[0][691] , 
        \zin[0][690] , \zin[0][689] , \zin[0][688] , \zin[0][687] , 
        \zin[0][686] , \zin[0][685] , \zin[0][684] , \zin[0][683] , 
        \zin[0][682] , \zin[0][681] , \zin[0][680] , \zin[0][679] , 
        \zin[0][678] , \zin[0][677] , \zin[0][676] , \zin[0][675] , 
        \zin[0][674] , \zin[0][673] , \zin[0][672] , \zin[0][671] , 
        \zin[0][670] , \zin[0][669] , \zin[0][668] , \zin[0][667] , 
        \zin[0][666] , \zin[0][665] , \zin[0][664] , \zin[0][663] , 
        \zin[0][662] , \zin[0][661] , \zin[0][660] , \zin[0][659] , 
        \zin[0][658] , \zin[0][657] , \zin[0][656] , \zin[0][655] , 
        \zin[0][654] , \zin[0][653] , \zin[0][652] , \zin[0][651] , 
        \zin[0][650] , \zin[0][649] , \zin[0][648] , \zin[0][647] , 
        \zin[0][646] , \zin[0][645] , \zin[0][644] , \zin[0][643] , 
        \zin[0][642] , \zin[0][641] , \zin[0][640] , \zin[0][639] , 
        \zin[0][638] , \zin[0][637] , \zin[0][636] , \zin[0][635] , 
        \zin[0][634] , \zin[0][633] , \zin[0][632] , \zin[0][631] , 
        \zin[0][630] , \zin[0][629] , \zin[0][628] , \zin[0][627] , 
        \zin[0][626] , \zin[0][625] , \zin[0][624] , \zin[0][623] , 
        \zin[0][622] , \zin[0][621] , \zin[0][620] , \zin[0][619] , 
        \zin[0][618] , \zin[0][617] , \zin[0][616] , \zin[0][615] , 
        \zin[0][614] , \zin[0][613] , \zin[0][612] , \zin[0][611] , 
        \zin[0][610] , \zin[0][609] , \zin[0][608] , \zin[0][607] , 
        \zin[0][606] , \zin[0][605] , \zin[0][604] , \zin[0][603] , 
        \zin[0][602] , \zin[0][601] , \zin[0][600] , \zin[0][599] , 
        \zin[0][598] , \zin[0][597] , \zin[0][596] , \zin[0][595] , 
        \zin[0][594] , \zin[0][593] , \zin[0][592] , \zin[0][591] , 
        \zin[0][590] , \zin[0][589] , \zin[0][588] , \zin[0][587] , 
        \zin[0][586] , \zin[0][585] , \zin[0][584] , \zin[0][583] , 
        \zin[0][582] , \zin[0][581] , \zin[0][580] , \zin[0][579] , 
        \zin[0][578] , \zin[0][577] , \zin[0][576] , \zin[0][575] , 
        \zin[0][574] , \zin[0][573] , \zin[0][572] , \zin[0][571] , 
        \zin[0][570] , \zin[0][569] , \zin[0][568] , \zin[0][567] , 
        \zin[0][566] , \zin[0][565] , \zin[0][564] , \zin[0][563] , 
        \zin[0][562] , \zin[0][561] , \zin[0][560] , \zin[0][559] , 
        \zin[0][558] , \zin[0][557] , \zin[0][556] , \zin[0][555] , 
        \zin[0][554] , \zin[0][553] , \zin[0][552] , \zin[0][551] , 
        \zin[0][550] , \zin[0][549] , \zin[0][548] , \zin[0][547] , 
        \zin[0][546] , \zin[0][545] , \zin[0][544] , \zin[0][543] , 
        \zin[0][542] , \zin[0][541] , \zin[0][540] , \zin[0][539] , 
        \zin[0][538] , \zin[0][537] , \zin[0][536] , \zin[0][535] , 
        \zin[0][534] , \zin[0][533] , \zin[0][532] , \zin[0][531] , 
        \zin[0][530] , \zin[0][529] , \zin[0][528] , \zin[0][527] , 
        \zin[0][526] , \zin[0][525] , \zin[0][524] , \zin[0][523] , 
        \zin[0][522] , \zin[0][521] , \zin[0][520] , \zin[0][519] , 
        \zin[0][518] , \zin[0][517] , \zin[0][516] , \zin[0][515] , 
        \zin[0][514] , \zin[0][513] , \zin[0][512] , \zin[0][511] , 
        \zin[0][510] , \zin[0][509] , \zin[0][508] , \zin[0][507] , 
        \zin[0][506] , \zin[0][505] , \zin[0][504] , \zin[0][503] , 
        \zin[0][502] , \zin[0][501] , \zin[0][500] , \zin[0][499] , 
        \zin[0][498] , \zin[0][497] , \zin[0][496] , \zin[0][495] , 
        \zin[0][494] , \zin[0][493] , \zin[0][492] , \zin[0][491] , 
        \zin[0][490] , \zin[0][489] , \zin[0][488] , \zin[0][487] , 
        \zin[0][486] , \zin[0][485] , \zin[0][484] , \zin[0][483] , 
        \zin[0][482] , \zin[0][481] , \zin[0][480] , \zin[0][479] , 
        \zin[0][478] , \zin[0][477] , \zin[0][476] , \zin[0][475] , 
        \zin[0][474] , \zin[0][473] , \zin[0][472] , \zin[0][471] , 
        \zin[0][470] , \zin[0][469] , \zin[0][468] , \zin[0][467] , 
        \zin[0][466] , \zin[0][465] , \zin[0][464] , \zin[0][463] , 
        \zin[0][462] , \zin[0][461] , \zin[0][460] , \zin[0][459] , 
        \zin[0][458] , \zin[0][457] , \zin[0][456] , \zin[0][455] , 
        \zin[0][454] , \zin[0][453] , \zin[0][452] , \zin[0][451] , 
        \zin[0][450] , \zin[0][449] , \zin[0][448] , \zin[0][447] , 
        \zin[0][446] , \zin[0][445] , \zin[0][444] , \zin[0][443] , 
        \zin[0][442] , \zin[0][441] , \zin[0][440] , \zin[0][439] , 
        \zin[0][438] , \zin[0][437] , \zin[0][436] , \zin[0][435] , 
        \zin[0][434] , \zin[0][433] , \zin[0][432] , \zin[0][431] , 
        \zin[0][430] , \zin[0][429] , \zin[0][428] , \zin[0][427] , 
        \zin[0][426] , \zin[0][425] , \zin[0][424] , \zin[0][423] , 
        \zin[0][422] , \zin[0][421] , \zin[0][420] , \zin[0][419] , 
        \zin[0][418] , \zin[0][417] , \zin[0][416] , \zin[0][415] , 
        \zin[0][414] , \zin[0][413] , \zin[0][412] , \zin[0][411] , 
        \zin[0][410] , \zin[0][409] , \zin[0][408] , \zin[0][407] , 
        \zin[0][406] , \zin[0][405] , \zin[0][404] , \zin[0][403] , 
        \zin[0][402] , \zin[0][401] , \zin[0][400] , \zin[0][399] , 
        \zin[0][398] , \zin[0][397] , \zin[0][396] , \zin[0][395] , 
        \zin[0][394] , \zin[0][393] , \zin[0][392] , \zin[0][391] , 
        \zin[0][390] , \zin[0][389] , \zin[0][388] , \zin[0][387] , 
        \zin[0][386] , \zin[0][385] , \zin[0][384] , \zin[0][383] , 
        \zin[0][382] , \zin[0][381] , \zin[0][380] , \zin[0][379] , 
        \zin[0][378] , \zin[0][377] , \zin[0][376] , \zin[0][375] , 
        \zin[0][374] , \zin[0][373] , \zin[0][372] , \zin[0][371] , 
        \zin[0][370] , \zin[0][369] , \zin[0][368] , \zin[0][367] , 
        \zin[0][366] , \zin[0][365] , \zin[0][364] , \zin[0][363] , 
        \zin[0][362] , \zin[0][361] , \zin[0][360] , \zin[0][359] , 
        \zin[0][358] , \zin[0][357] , \zin[0][356] , \zin[0][355] , 
        \zin[0][354] , \zin[0][353] , \zin[0][352] , \zin[0][351] , 
        \zin[0][350] , \zin[0][349] , \zin[0][348] , \zin[0][347] , 
        \zin[0][346] , \zin[0][345] , \zin[0][344] , \zin[0][343] , 
        \zin[0][342] , \zin[0][341] , \zin[0][340] , \zin[0][339] , 
        \zin[0][338] , \zin[0][337] , \zin[0][336] , \zin[0][335] , 
        \zin[0][334] , \zin[0][333] , \zin[0][332] , \zin[0][331] , 
        \zin[0][330] , \zin[0][329] , \zin[0][328] , \zin[0][327] , 
        \zin[0][326] , \zin[0][325] , \zin[0][324] , \zin[0][323] , 
        \zin[0][322] , \zin[0][321] , \zin[0][320] , \zin[0][319] , 
        \zin[0][318] , \zin[0][317] , \zin[0][316] , \zin[0][315] , 
        \zin[0][314] , \zin[0][313] , \zin[0][312] , \zin[0][311] , 
        \zin[0][310] , \zin[0][309] , \zin[0][308] , \zin[0][307] , 
        \zin[0][306] , \zin[0][305] , \zin[0][304] , \zin[0][303] , 
        \zin[0][302] , \zin[0][301] , \zin[0][300] , \zin[0][299] , 
        \zin[0][298] , \zin[0][297] , \zin[0][296] , \zin[0][295] , 
        \zin[0][294] , \zin[0][293] , \zin[0][292] , \zin[0][291] , 
        \zin[0][290] , \zin[0][289] , \zin[0][288] , \zin[0][287] , 
        \zin[0][286] , \zin[0][285] , \zin[0][284] , \zin[0][283] , 
        \zin[0][282] , \zin[0][281] , \zin[0][280] , \zin[0][279] , 
        \zin[0][278] , \zin[0][277] , \zin[0][276] , \zin[0][275] , 
        \zin[0][274] , \zin[0][273] , \zin[0][272] , \zin[0][271] , 
        \zin[0][270] , \zin[0][269] , \zin[0][268] , \zin[0][267] , 
        \zin[0][266] , \zin[0][265] , \zin[0][264] , \zin[0][263] , 
        \zin[0][262] , \zin[0][261] , \zin[0][260] , \zin[0][259] , 
        \zin[0][258] , \zin[0][257] , \zin[0][256] , \zin[0][255] , 
        \zin[0][254] , \zin[0][253] , \zin[0][252] , \zin[0][251] , 
        \zin[0][250] , \zin[0][249] , \zin[0][248] , \zin[0][247] , 
        \zin[0][246] , \zin[0][245] , \zin[0][244] , \zin[0][243] , 
        \zin[0][242] , \zin[0][241] , \zin[0][240] , \zin[0][239] , 
        \zin[0][238] , \zin[0][237] , \zin[0][236] , \zin[0][235] , 
        \zin[0][234] , \zin[0][233] , \zin[0][232] , \zin[0][231] , 
        \zin[0][230] , \zin[0][229] , \zin[0][228] , \zin[0][227] , 
        \zin[0][226] , \zin[0][225] , \zin[0][224] , \zin[0][223] , 
        \zin[0][222] , \zin[0][221] , \zin[0][220] , \zin[0][219] , 
        \zin[0][218] , \zin[0][217] , \zin[0][216] , \zin[0][215] , 
        \zin[0][214] , \zin[0][213] , \zin[0][212] , \zin[0][211] , 
        \zin[0][210] , \zin[0][209] , \zin[0][208] , \zin[0][207] , 
        \zin[0][206] , \zin[0][205] , \zin[0][204] , \zin[0][203] , 
        \zin[0][202] , \zin[0][201] , \zin[0][200] , \zin[0][199] , 
        \zin[0][198] , \zin[0][197] , \zin[0][196] , \zin[0][195] , 
        \zin[0][194] , \zin[0][193] , \zin[0][192] , \zin[0][191] , 
        \zin[0][190] , \zin[0][189] , \zin[0][188] , \zin[0][187] , 
        \zin[0][186] , \zin[0][185] , \zin[0][184] , \zin[0][183] , 
        \zin[0][182] , \zin[0][181] , \zin[0][180] , \zin[0][179] , 
        \zin[0][178] , \zin[0][177] , \zin[0][176] , \zin[0][175] , 
        \zin[0][174] , \zin[0][173] , \zin[0][172] , \zin[0][171] , 
        \zin[0][170] , \zin[0][169] , \zin[0][168] , \zin[0][167] , 
        \zin[0][166] , \zin[0][165] , \zin[0][164] , \zin[0][163] , 
        \zin[0][162] , \zin[0][161] , \zin[0][160] , \zin[0][159] , 
        \zin[0][158] , \zin[0][157] , \zin[0][156] , \zin[0][155] , 
        \zin[0][154] , \zin[0][153] , \zin[0][152] , \zin[0][151] , 
        \zin[0][150] , \zin[0][149] , \zin[0][148] , \zin[0][147] , 
        \zin[0][146] , \zin[0][145] , \zin[0][144] , \zin[0][143] , 
        \zin[0][142] , \zin[0][141] , \zin[0][140] , \zin[0][139] , 
        \zin[0][138] , \zin[0][137] , \zin[0][136] , \zin[0][135] , 
        \zin[0][134] , \zin[0][133] , \zin[0][132] , \zin[0][131] , 
        \zin[0][130] , \zin[0][129] , \zin[0][128] , \zin[0][127] , 
        \zin[0][126] , \zin[0][125] , \zin[0][124] , \zin[0][123] , 
        \zin[0][122] , \zin[0][121] , \zin[0][120] , \zin[0][119] , 
        \zin[0][118] , \zin[0][117] , \zin[0][116] , \zin[0][115] , 
        \zin[0][114] , \zin[0][113] , \zin[0][112] , \zin[0][111] , 
        \zin[0][110] , \zin[0][109] , \zin[0][108] , \zin[0][107] , 
        \zin[0][106] , \zin[0][105] , \zin[0][104] , \zin[0][103] , 
        \zin[0][102] , \zin[0][101] , \zin[0][100] , \zin[0][99] , 
        \zin[0][98] , \zin[0][97] , \zin[0][96] , \zin[0][95] , \zin[0][94] , 
        \zin[0][93] , \zin[0][92] , \zin[0][91] , \zin[0][90] , \zin[0][89] , 
        \zin[0][88] , \zin[0][87] , \zin[0][86] , \zin[0][85] , \zin[0][84] , 
        \zin[0][83] , \zin[0][82] , \zin[0][81] , \zin[0][80] , \zin[0][79] , 
        \zin[0][78] , \zin[0][77] , \zin[0][76] , \zin[0][75] , \zin[0][74] , 
        \zin[0][73] , \zin[0][72] , \zin[0][71] , \zin[0][70] , \zin[0][69] , 
        \zin[0][68] , \zin[0][67] , \zin[0][66] , \zin[0][65] , \zin[0][64] , 
        \zin[0][63] , \zin[0][62] , \zin[0][61] , \zin[0][60] , \zin[0][59] , 
        \zin[0][58] , \zin[0][57] , \zin[0][56] , \zin[0][55] , \zin[0][54] , 
        \zin[0][53] , \zin[0][52] , \zin[0][51] , \zin[0][50] , \zin[0][49] , 
        \zin[0][48] , \zin[0][47] , \zin[0][46] , \zin[0][45] , \zin[0][44] , 
        \zin[0][43] , \zin[0][42] , \zin[0][41] , \zin[0][40] , \zin[0][39] , 
        \zin[0][38] , \zin[0][37] , \zin[0][36] , \zin[0][35] , \zin[0][34] , 
        \zin[0][33] , \zin[0][32] , \zin[0][31] , \zin[0][30] , \zin[0][29] , 
        \zin[0][28] , \zin[0][27] , \zin[0][26] , \zin[0][25] , \zin[0][24] , 
        \zin[0][23] , \zin[0][22] , \zin[0][21] , \zin[0][20] , \zin[0][19] , 
        \zin[0][18] , \zin[0][17] , \zin[0][16] , \zin[0][15] , \zin[0][14] , 
        \zin[0][13] , \zin[0][12] , \zin[0][11] , \zin[0][10] , \zin[0][9] , 
        \zin[0][8] , \zin[0][7] , \zin[0][6] , \zin[0][5] , \zin[0][4] , 
        \zin[0][3] , \zin[0][2] , \zin[0][1] , \zin[0][0] }), .zout({
        SYNOPSYS_UNCONNECTED__0, \zout[0][1024] , o}) );
  DFF \xreg_reg[0]  ( .D(1'b0), .CLK(clk), .RST(start), .I(x[0]), .Q(xin[0])
         );
  DFF \xreg_reg[1]  ( .D(xin[0]), .CLK(clk), .RST(start), .I(x[1]), .Q(xin[1])
         );
  DFF \xreg_reg[2]  ( .D(xin[1]), .CLK(clk), .RST(start), .I(x[2]), .Q(xin[2])
         );
  DFF \xreg_reg[3]  ( .D(xin[2]), .CLK(clk), .RST(start), .I(x[3]), .Q(xin[3])
         );
  DFF \xreg_reg[4]  ( .D(xin[3]), .CLK(clk), .RST(start), .I(x[4]), .Q(xin[4])
         );
  DFF \xreg_reg[5]  ( .D(xin[4]), .CLK(clk), .RST(start), .I(x[5]), .Q(xin[5])
         );
  DFF \xreg_reg[6]  ( .D(xin[5]), .CLK(clk), .RST(start), .I(x[6]), .Q(xin[6])
         );
  DFF \xreg_reg[7]  ( .D(xin[6]), .CLK(clk), .RST(start), .I(x[7]), .Q(xin[7])
         );
  DFF \xreg_reg[8]  ( .D(xin[7]), .CLK(clk), .RST(start), .I(x[8]), .Q(xin[8])
         );
  DFF \xreg_reg[9]  ( .D(xin[8]), .CLK(clk), .RST(start), .I(x[9]), .Q(xin[9])
         );
  DFF \xreg_reg[10]  ( .D(xin[9]), .CLK(clk), .RST(start), .I(x[10]), .Q(
        xin[10]) );
  DFF \xreg_reg[11]  ( .D(xin[10]), .CLK(clk), .RST(start), .I(x[11]), .Q(
        xin[11]) );
  DFF \xreg_reg[12]  ( .D(xin[11]), .CLK(clk), .RST(start), .I(x[12]), .Q(
        xin[12]) );
  DFF \xreg_reg[13]  ( .D(xin[12]), .CLK(clk), .RST(start), .I(x[13]), .Q(
        xin[13]) );
  DFF \xreg_reg[14]  ( .D(xin[13]), .CLK(clk), .RST(start), .I(x[14]), .Q(
        xin[14]) );
  DFF \xreg_reg[15]  ( .D(xin[14]), .CLK(clk), .RST(start), .I(x[15]), .Q(
        xin[15]) );
  DFF \xreg_reg[16]  ( .D(xin[15]), .CLK(clk), .RST(start), .I(x[16]), .Q(
        xin[16]) );
  DFF \xreg_reg[17]  ( .D(xin[16]), .CLK(clk), .RST(start), .I(x[17]), .Q(
        xin[17]) );
  DFF \xreg_reg[18]  ( .D(xin[17]), .CLK(clk), .RST(start), .I(x[18]), .Q(
        xin[18]) );
  DFF \xreg_reg[19]  ( .D(xin[18]), .CLK(clk), .RST(start), .I(x[19]), .Q(
        xin[19]) );
  DFF \xreg_reg[20]  ( .D(xin[19]), .CLK(clk), .RST(start), .I(x[20]), .Q(
        xin[20]) );
  DFF \xreg_reg[21]  ( .D(xin[20]), .CLK(clk), .RST(start), .I(x[21]), .Q(
        xin[21]) );
  DFF \xreg_reg[22]  ( .D(xin[21]), .CLK(clk), .RST(start), .I(x[22]), .Q(
        xin[22]) );
  DFF \xreg_reg[23]  ( .D(xin[22]), .CLK(clk), .RST(start), .I(x[23]), .Q(
        xin[23]) );
  DFF \xreg_reg[24]  ( .D(xin[23]), .CLK(clk), .RST(start), .I(x[24]), .Q(
        xin[24]) );
  DFF \xreg_reg[25]  ( .D(xin[24]), .CLK(clk), .RST(start), .I(x[25]), .Q(
        xin[25]) );
  DFF \xreg_reg[26]  ( .D(xin[25]), .CLK(clk), .RST(start), .I(x[26]), .Q(
        xin[26]) );
  DFF \xreg_reg[27]  ( .D(xin[26]), .CLK(clk), .RST(start), .I(x[27]), .Q(
        xin[27]) );
  DFF \xreg_reg[28]  ( .D(xin[27]), .CLK(clk), .RST(start), .I(x[28]), .Q(
        xin[28]) );
  DFF \xreg_reg[29]  ( .D(xin[28]), .CLK(clk), .RST(start), .I(x[29]), .Q(
        xin[29]) );
  DFF \xreg_reg[30]  ( .D(xin[29]), .CLK(clk), .RST(start), .I(x[30]), .Q(
        xin[30]) );
  DFF \xreg_reg[31]  ( .D(xin[30]), .CLK(clk), .RST(start), .I(x[31]), .Q(
        xin[31]) );
  DFF \xreg_reg[32]  ( .D(xin[31]), .CLK(clk), .RST(start), .I(x[32]), .Q(
        xin[32]) );
  DFF \xreg_reg[33]  ( .D(xin[32]), .CLK(clk), .RST(start), .I(x[33]), .Q(
        xin[33]) );
  DFF \xreg_reg[34]  ( .D(xin[33]), .CLK(clk), .RST(start), .I(x[34]), .Q(
        xin[34]) );
  DFF \xreg_reg[35]  ( .D(xin[34]), .CLK(clk), .RST(start), .I(x[35]), .Q(
        xin[35]) );
  DFF \xreg_reg[36]  ( .D(xin[35]), .CLK(clk), .RST(start), .I(x[36]), .Q(
        xin[36]) );
  DFF \xreg_reg[37]  ( .D(xin[36]), .CLK(clk), .RST(start), .I(x[37]), .Q(
        xin[37]) );
  DFF \xreg_reg[38]  ( .D(xin[37]), .CLK(clk), .RST(start), .I(x[38]), .Q(
        xin[38]) );
  DFF \xreg_reg[39]  ( .D(xin[38]), .CLK(clk), .RST(start), .I(x[39]), .Q(
        xin[39]) );
  DFF \xreg_reg[40]  ( .D(xin[39]), .CLK(clk), .RST(start), .I(x[40]), .Q(
        xin[40]) );
  DFF \xreg_reg[41]  ( .D(xin[40]), .CLK(clk), .RST(start), .I(x[41]), .Q(
        xin[41]) );
  DFF \xreg_reg[42]  ( .D(xin[41]), .CLK(clk), .RST(start), .I(x[42]), .Q(
        xin[42]) );
  DFF \xreg_reg[43]  ( .D(xin[42]), .CLK(clk), .RST(start), .I(x[43]), .Q(
        xin[43]) );
  DFF \xreg_reg[44]  ( .D(xin[43]), .CLK(clk), .RST(start), .I(x[44]), .Q(
        xin[44]) );
  DFF \xreg_reg[45]  ( .D(xin[44]), .CLK(clk), .RST(start), .I(x[45]), .Q(
        xin[45]) );
  DFF \xreg_reg[46]  ( .D(xin[45]), .CLK(clk), .RST(start), .I(x[46]), .Q(
        xin[46]) );
  DFF \xreg_reg[47]  ( .D(xin[46]), .CLK(clk), .RST(start), .I(x[47]), .Q(
        xin[47]) );
  DFF \xreg_reg[48]  ( .D(xin[47]), .CLK(clk), .RST(start), .I(x[48]), .Q(
        xin[48]) );
  DFF \xreg_reg[49]  ( .D(xin[48]), .CLK(clk), .RST(start), .I(x[49]), .Q(
        xin[49]) );
  DFF \xreg_reg[50]  ( .D(xin[49]), .CLK(clk), .RST(start), .I(x[50]), .Q(
        xin[50]) );
  DFF \xreg_reg[51]  ( .D(xin[50]), .CLK(clk), .RST(start), .I(x[51]), .Q(
        xin[51]) );
  DFF \xreg_reg[52]  ( .D(xin[51]), .CLK(clk), .RST(start), .I(x[52]), .Q(
        xin[52]) );
  DFF \xreg_reg[53]  ( .D(xin[52]), .CLK(clk), .RST(start), .I(x[53]), .Q(
        xin[53]) );
  DFF \xreg_reg[54]  ( .D(xin[53]), .CLK(clk), .RST(start), .I(x[54]), .Q(
        xin[54]) );
  DFF \xreg_reg[55]  ( .D(xin[54]), .CLK(clk), .RST(start), .I(x[55]), .Q(
        xin[55]) );
  DFF \xreg_reg[56]  ( .D(xin[55]), .CLK(clk), .RST(start), .I(x[56]), .Q(
        xin[56]) );
  DFF \xreg_reg[57]  ( .D(xin[56]), .CLK(clk), .RST(start), .I(x[57]), .Q(
        xin[57]) );
  DFF \xreg_reg[58]  ( .D(xin[57]), .CLK(clk), .RST(start), .I(x[58]), .Q(
        xin[58]) );
  DFF \xreg_reg[59]  ( .D(xin[58]), .CLK(clk), .RST(start), .I(x[59]), .Q(
        xin[59]) );
  DFF \xreg_reg[60]  ( .D(xin[59]), .CLK(clk), .RST(start), .I(x[60]), .Q(
        xin[60]) );
  DFF \xreg_reg[61]  ( .D(xin[60]), .CLK(clk), .RST(start), .I(x[61]), .Q(
        xin[61]) );
  DFF \xreg_reg[62]  ( .D(xin[61]), .CLK(clk), .RST(start), .I(x[62]), .Q(
        xin[62]) );
  DFF \xreg_reg[63]  ( .D(xin[62]), .CLK(clk), .RST(start), .I(x[63]), .Q(
        xin[63]) );
  DFF \xreg_reg[64]  ( .D(xin[63]), .CLK(clk), .RST(start), .I(x[64]), .Q(
        xin[64]) );
  DFF \xreg_reg[65]  ( .D(xin[64]), .CLK(clk), .RST(start), .I(x[65]), .Q(
        xin[65]) );
  DFF \xreg_reg[66]  ( .D(xin[65]), .CLK(clk), .RST(start), .I(x[66]), .Q(
        xin[66]) );
  DFF \xreg_reg[67]  ( .D(xin[66]), .CLK(clk), .RST(start), .I(x[67]), .Q(
        xin[67]) );
  DFF \xreg_reg[68]  ( .D(xin[67]), .CLK(clk), .RST(start), .I(x[68]), .Q(
        xin[68]) );
  DFF \xreg_reg[69]  ( .D(xin[68]), .CLK(clk), .RST(start), .I(x[69]), .Q(
        xin[69]) );
  DFF \xreg_reg[70]  ( .D(xin[69]), .CLK(clk), .RST(start), .I(x[70]), .Q(
        xin[70]) );
  DFF \xreg_reg[71]  ( .D(xin[70]), .CLK(clk), .RST(start), .I(x[71]), .Q(
        xin[71]) );
  DFF \xreg_reg[72]  ( .D(xin[71]), .CLK(clk), .RST(start), .I(x[72]), .Q(
        xin[72]) );
  DFF \xreg_reg[73]  ( .D(xin[72]), .CLK(clk), .RST(start), .I(x[73]), .Q(
        xin[73]) );
  DFF \xreg_reg[74]  ( .D(xin[73]), .CLK(clk), .RST(start), .I(x[74]), .Q(
        xin[74]) );
  DFF \xreg_reg[75]  ( .D(xin[74]), .CLK(clk), .RST(start), .I(x[75]), .Q(
        xin[75]) );
  DFF \xreg_reg[76]  ( .D(xin[75]), .CLK(clk), .RST(start), .I(x[76]), .Q(
        xin[76]) );
  DFF \xreg_reg[77]  ( .D(xin[76]), .CLK(clk), .RST(start), .I(x[77]), .Q(
        xin[77]) );
  DFF \xreg_reg[78]  ( .D(xin[77]), .CLK(clk), .RST(start), .I(x[78]), .Q(
        xin[78]) );
  DFF \xreg_reg[79]  ( .D(xin[78]), .CLK(clk), .RST(start), .I(x[79]), .Q(
        xin[79]) );
  DFF \xreg_reg[80]  ( .D(xin[79]), .CLK(clk), .RST(start), .I(x[80]), .Q(
        xin[80]) );
  DFF \xreg_reg[81]  ( .D(xin[80]), .CLK(clk), .RST(start), .I(x[81]), .Q(
        xin[81]) );
  DFF \xreg_reg[82]  ( .D(xin[81]), .CLK(clk), .RST(start), .I(x[82]), .Q(
        xin[82]) );
  DFF \xreg_reg[83]  ( .D(xin[82]), .CLK(clk), .RST(start), .I(x[83]), .Q(
        xin[83]) );
  DFF \xreg_reg[84]  ( .D(xin[83]), .CLK(clk), .RST(start), .I(x[84]), .Q(
        xin[84]) );
  DFF \xreg_reg[85]  ( .D(xin[84]), .CLK(clk), .RST(start), .I(x[85]), .Q(
        xin[85]) );
  DFF \xreg_reg[86]  ( .D(xin[85]), .CLK(clk), .RST(start), .I(x[86]), .Q(
        xin[86]) );
  DFF \xreg_reg[87]  ( .D(xin[86]), .CLK(clk), .RST(start), .I(x[87]), .Q(
        xin[87]) );
  DFF \xreg_reg[88]  ( .D(xin[87]), .CLK(clk), .RST(start), .I(x[88]), .Q(
        xin[88]) );
  DFF \xreg_reg[89]  ( .D(xin[88]), .CLK(clk), .RST(start), .I(x[89]), .Q(
        xin[89]) );
  DFF \xreg_reg[90]  ( .D(xin[89]), .CLK(clk), .RST(start), .I(x[90]), .Q(
        xin[90]) );
  DFF \xreg_reg[91]  ( .D(xin[90]), .CLK(clk), .RST(start), .I(x[91]), .Q(
        xin[91]) );
  DFF \xreg_reg[92]  ( .D(xin[91]), .CLK(clk), .RST(start), .I(x[92]), .Q(
        xin[92]) );
  DFF \xreg_reg[93]  ( .D(xin[92]), .CLK(clk), .RST(start), .I(x[93]), .Q(
        xin[93]) );
  DFF \xreg_reg[94]  ( .D(xin[93]), .CLK(clk), .RST(start), .I(x[94]), .Q(
        xin[94]) );
  DFF \xreg_reg[95]  ( .D(xin[94]), .CLK(clk), .RST(start), .I(x[95]), .Q(
        xin[95]) );
  DFF \xreg_reg[96]  ( .D(xin[95]), .CLK(clk), .RST(start), .I(x[96]), .Q(
        xin[96]) );
  DFF \xreg_reg[97]  ( .D(xin[96]), .CLK(clk), .RST(start), .I(x[97]), .Q(
        xin[97]) );
  DFF \xreg_reg[98]  ( .D(xin[97]), .CLK(clk), .RST(start), .I(x[98]), .Q(
        xin[98]) );
  DFF \xreg_reg[99]  ( .D(xin[98]), .CLK(clk), .RST(start), .I(x[99]), .Q(
        xin[99]) );
  DFF \xreg_reg[100]  ( .D(xin[99]), .CLK(clk), .RST(start), .I(x[100]), .Q(
        xin[100]) );
  DFF \xreg_reg[101]  ( .D(xin[100]), .CLK(clk), .RST(start), .I(x[101]), .Q(
        xin[101]) );
  DFF \xreg_reg[102]  ( .D(xin[101]), .CLK(clk), .RST(start), .I(x[102]), .Q(
        xin[102]) );
  DFF \xreg_reg[103]  ( .D(xin[102]), .CLK(clk), .RST(start), .I(x[103]), .Q(
        xin[103]) );
  DFF \xreg_reg[104]  ( .D(xin[103]), .CLK(clk), .RST(start), .I(x[104]), .Q(
        xin[104]) );
  DFF \xreg_reg[105]  ( .D(xin[104]), .CLK(clk), .RST(start), .I(x[105]), .Q(
        xin[105]) );
  DFF \xreg_reg[106]  ( .D(xin[105]), .CLK(clk), .RST(start), .I(x[106]), .Q(
        xin[106]) );
  DFF \xreg_reg[107]  ( .D(xin[106]), .CLK(clk), .RST(start), .I(x[107]), .Q(
        xin[107]) );
  DFF \xreg_reg[108]  ( .D(xin[107]), .CLK(clk), .RST(start), .I(x[108]), .Q(
        xin[108]) );
  DFF \xreg_reg[109]  ( .D(xin[108]), .CLK(clk), .RST(start), .I(x[109]), .Q(
        xin[109]) );
  DFF \xreg_reg[110]  ( .D(xin[109]), .CLK(clk), .RST(start), .I(x[110]), .Q(
        xin[110]) );
  DFF \xreg_reg[111]  ( .D(xin[110]), .CLK(clk), .RST(start), .I(x[111]), .Q(
        xin[111]) );
  DFF \xreg_reg[112]  ( .D(xin[111]), .CLK(clk), .RST(start), .I(x[112]), .Q(
        xin[112]) );
  DFF \xreg_reg[113]  ( .D(xin[112]), .CLK(clk), .RST(start), .I(x[113]), .Q(
        xin[113]) );
  DFF \xreg_reg[114]  ( .D(xin[113]), .CLK(clk), .RST(start), .I(x[114]), .Q(
        xin[114]) );
  DFF \xreg_reg[115]  ( .D(xin[114]), .CLK(clk), .RST(start), .I(x[115]), .Q(
        xin[115]) );
  DFF \xreg_reg[116]  ( .D(xin[115]), .CLK(clk), .RST(start), .I(x[116]), .Q(
        xin[116]) );
  DFF \xreg_reg[117]  ( .D(xin[116]), .CLK(clk), .RST(start), .I(x[117]), .Q(
        xin[117]) );
  DFF \xreg_reg[118]  ( .D(xin[117]), .CLK(clk), .RST(start), .I(x[118]), .Q(
        xin[118]) );
  DFF \xreg_reg[119]  ( .D(xin[118]), .CLK(clk), .RST(start), .I(x[119]), .Q(
        xin[119]) );
  DFF \xreg_reg[120]  ( .D(xin[119]), .CLK(clk), .RST(start), .I(x[120]), .Q(
        xin[120]) );
  DFF \xreg_reg[121]  ( .D(xin[120]), .CLK(clk), .RST(start), .I(x[121]), .Q(
        xin[121]) );
  DFF \xreg_reg[122]  ( .D(xin[121]), .CLK(clk), .RST(start), .I(x[122]), .Q(
        xin[122]) );
  DFF \xreg_reg[123]  ( .D(xin[122]), .CLK(clk), .RST(start), .I(x[123]), .Q(
        xin[123]) );
  DFF \xreg_reg[124]  ( .D(xin[123]), .CLK(clk), .RST(start), .I(x[124]), .Q(
        xin[124]) );
  DFF \xreg_reg[125]  ( .D(xin[124]), .CLK(clk), .RST(start), .I(x[125]), .Q(
        xin[125]) );
  DFF \xreg_reg[126]  ( .D(xin[125]), .CLK(clk), .RST(start), .I(x[126]), .Q(
        xin[126]) );
  DFF \xreg_reg[127]  ( .D(xin[126]), .CLK(clk), .RST(start), .I(x[127]), .Q(
        xin[127]) );
  DFF \xreg_reg[128]  ( .D(xin[127]), .CLK(clk), .RST(start), .I(x[128]), .Q(
        xin[128]) );
  DFF \xreg_reg[129]  ( .D(xin[128]), .CLK(clk), .RST(start), .I(x[129]), .Q(
        xin[129]) );
  DFF \xreg_reg[130]  ( .D(xin[129]), .CLK(clk), .RST(start), .I(x[130]), .Q(
        xin[130]) );
  DFF \xreg_reg[131]  ( .D(xin[130]), .CLK(clk), .RST(start), .I(x[131]), .Q(
        xin[131]) );
  DFF \xreg_reg[132]  ( .D(xin[131]), .CLK(clk), .RST(start), .I(x[132]), .Q(
        xin[132]) );
  DFF \xreg_reg[133]  ( .D(xin[132]), .CLK(clk), .RST(start), .I(x[133]), .Q(
        xin[133]) );
  DFF \xreg_reg[134]  ( .D(xin[133]), .CLK(clk), .RST(start), .I(x[134]), .Q(
        xin[134]) );
  DFF \xreg_reg[135]  ( .D(xin[134]), .CLK(clk), .RST(start), .I(x[135]), .Q(
        xin[135]) );
  DFF \xreg_reg[136]  ( .D(xin[135]), .CLK(clk), .RST(start), .I(x[136]), .Q(
        xin[136]) );
  DFF \xreg_reg[137]  ( .D(xin[136]), .CLK(clk), .RST(start), .I(x[137]), .Q(
        xin[137]) );
  DFF \xreg_reg[138]  ( .D(xin[137]), .CLK(clk), .RST(start), .I(x[138]), .Q(
        xin[138]) );
  DFF \xreg_reg[139]  ( .D(xin[138]), .CLK(clk), .RST(start), .I(x[139]), .Q(
        xin[139]) );
  DFF \xreg_reg[140]  ( .D(xin[139]), .CLK(clk), .RST(start), .I(x[140]), .Q(
        xin[140]) );
  DFF \xreg_reg[141]  ( .D(xin[140]), .CLK(clk), .RST(start), .I(x[141]), .Q(
        xin[141]) );
  DFF \xreg_reg[142]  ( .D(xin[141]), .CLK(clk), .RST(start), .I(x[142]), .Q(
        xin[142]) );
  DFF \xreg_reg[143]  ( .D(xin[142]), .CLK(clk), .RST(start), .I(x[143]), .Q(
        xin[143]) );
  DFF \xreg_reg[144]  ( .D(xin[143]), .CLK(clk), .RST(start), .I(x[144]), .Q(
        xin[144]) );
  DFF \xreg_reg[145]  ( .D(xin[144]), .CLK(clk), .RST(start), .I(x[145]), .Q(
        xin[145]) );
  DFF \xreg_reg[146]  ( .D(xin[145]), .CLK(clk), .RST(start), .I(x[146]), .Q(
        xin[146]) );
  DFF \xreg_reg[147]  ( .D(xin[146]), .CLK(clk), .RST(start), .I(x[147]), .Q(
        xin[147]) );
  DFF \xreg_reg[148]  ( .D(xin[147]), .CLK(clk), .RST(start), .I(x[148]), .Q(
        xin[148]) );
  DFF \xreg_reg[149]  ( .D(xin[148]), .CLK(clk), .RST(start), .I(x[149]), .Q(
        xin[149]) );
  DFF \xreg_reg[150]  ( .D(xin[149]), .CLK(clk), .RST(start), .I(x[150]), .Q(
        xin[150]) );
  DFF \xreg_reg[151]  ( .D(xin[150]), .CLK(clk), .RST(start), .I(x[151]), .Q(
        xin[151]) );
  DFF \xreg_reg[152]  ( .D(xin[151]), .CLK(clk), .RST(start), .I(x[152]), .Q(
        xin[152]) );
  DFF \xreg_reg[153]  ( .D(xin[152]), .CLK(clk), .RST(start), .I(x[153]), .Q(
        xin[153]) );
  DFF \xreg_reg[154]  ( .D(xin[153]), .CLK(clk), .RST(start), .I(x[154]), .Q(
        xin[154]) );
  DFF \xreg_reg[155]  ( .D(xin[154]), .CLK(clk), .RST(start), .I(x[155]), .Q(
        xin[155]) );
  DFF \xreg_reg[156]  ( .D(xin[155]), .CLK(clk), .RST(start), .I(x[156]), .Q(
        xin[156]) );
  DFF \xreg_reg[157]  ( .D(xin[156]), .CLK(clk), .RST(start), .I(x[157]), .Q(
        xin[157]) );
  DFF \xreg_reg[158]  ( .D(xin[157]), .CLK(clk), .RST(start), .I(x[158]), .Q(
        xin[158]) );
  DFF \xreg_reg[159]  ( .D(xin[158]), .CLK(clk), .RST(start), .I(x[159]), .Q(
        xin[159]) );
  DFF \xreg_reg[160]  ( .D(xin[159]), .CLK(clk), .RST(start), .I(x[160]), .Q(
        xin[160]) );
  DFF \xreg_reg[161]  ( .D(xin[160]), .CLK(clk), .RST(start), .I(x[161]), .Q(
        xin[161]) );
  DFF \xreg_reg[162]  ( .D(xin[161]), .CLK(clk), .RST(start), .I(x[162]), .Q(
        xin[162]) );
  DFF \xreg_reg[163]  ( .D(xin[162]), .CLK(clk), .RST(start), .I(x[163]), .Q(
        xin[163]) );
  DFF \xreg_reg[164]  ( .D(xin[163]), .CLK(clk), .RST(start), .I(x[164]), .Q(
        xin[164]) );
  DFF \xreg_reg[165]  ( .D(xin[164]), .CLK(clk), .RST(start), .I(x[165]), .Q(
        xin[165]) );
  DFF \xreg_reg[166]  ( .D(xin[165]), .CLK(clk), .RST(start), .I(x[166]), .Q(
        xin[166]) );
  DFF \xreg_reg[167]  ( .D(xin[166]), .CLK(clk), .RST(start), .I(x[167]), .Q(
        xin[167]) );
  DFF \xreg_reg[168]  ( .D(xin[167]), .CLK(clk), .RST(start), .I(x[168]), .Q(
        xin[168]) );
  DFF \xreg_reg[169]  ( .D(xin[168]), .CLK(clk), .RST(start), .I(x[169]), .Q(
        xin[169]) );
  DFF \xreg_reg[170]  ( .D(xin[169]), .CLK(clk), .RST(start), .I(x[170]), .Q(
        xin[170]) );
  DFF \xreg_reg[171]  ( .D(xin[170]), .CLK(clk), .RST(start), .I(x[171]), .Q(
        xin[171]) );
  DFF \xreg_reg[172]  ( .D(xin[171]), .CLK(clk), .RST(start), .I(x[172]), .Q(
        xin[172]) );
  DFF \xreg_reg[173]  ( .D(xin[172]), .CLK(clk), .RST(start), .I(x[173]), .Q(
        xin[173]) );
  DFF \xreg_reg[174]  ( .D(xin[173]), .CLK(clk), .RST(start), .I(x[174]), .Q(
        xin[174]) );
  DFF \xreg_reg[175]  ( .D(xin[174]), .CLK(clk), .RST(start), .I(x[175]), .Q(
        xin[175]) );
  DFF \xreg_reg[176]  ( .D(xin[175]), .CLK(clk), .RST(start), .I(x[176]), .Q(
        xin[176]) );
  DFF \xreg_reg[177]  ( .D(xin[176]), .CLK(clk), .RST(start), .I(x[177]), .Q(
        xin[177]) );
  DFF \xreg_reg[178]  ( .D(xin[177]), .CLK(clk), .RST(start), .I(x[178]), .Q(
        xin[178]) );
  DFF \xreg_reg[179]  ( .D(xin[178]), .CLK(clk), .RST(start), .I(x[179]), .Q(
        xin[179]) );
  DFF \xreg_reg[180]  ( .D(xin[179]), .CLK(clk), .RST(start), .I(x[180]), .Q(
        xin[180]) );
  DFF \xreg_reg[181]  ( .D(xin[180]), .CLK(clk), .RST(start), .I(x[181]), .Q(
        xin[181]) );
  DFF \xreg_reg[182]  ( .D(xin[181]), .CLK(clk), .RST(start), .I(x[182]), .Q(
        xin[182]) );
  DFF \xreg_reg[183]  ( .D(xin[182]), .CLK(clk), .RST(start), .I(x[183]), .Q(
        xin[183]) );
  DFF \xreg_reg[184]  ( .D(xin[183]), .CLK(clk), .RST(start), .I(x[184]), .Q(
        xin[184]) );
  DFF \xreg_reg[185]  ( .D(xin[184]), .CLK(clk), .RST(start), .I(x[185]), .Q(
        xin[185]) );
  DFF \xreg_reg[186]  ( .D(xin[185]), .CLK(clk), .RST(start), .I(x[186]), .Q(
        xin[186]) );
  DFF \xreg_reg[187]  ( .D(xin[186]), .CLK(clk), .RST(start), .I(x[187]), .Q(
        xin[187]) );
  DFF \xreg_reg[188]  ( .D(xin[187]), .CLK(clk), .RST(start), .I(x[188]), .Q(
        xin[188]) );
  DFF \xreg_reg[189]  ( .D(xin[188]), .CLK(clk), .RST(start), .I(x[189]), .Q(
        xin[189]) );
  DFF \xreg_reg[190]  ( .D(xin[189]), .CLK(clk), .RST(start), .I(x[190]), .Q(
        xin[190]) );
  DFF \xreg_reg[191]  ( .D(xin[190]), .CLK(clk), .RST(start), .I(x[191]), .Q(
        xin[191]) );
  DFF \xreg_reg[192]  ( .D(xin[191]), .CLK(clk), .RST(start), .I(x[192]), .Q(
        xin[192]) );
  DFF \xreg_reg[193]  ( .D(xin[192]), .CLK(clk), .RST(start), .I(x[193]), .Q(
        xin[193]) );
  DFF \xreg_reg[194]  ( .D(xin[193]), .CLK(clk), .RST(start), .I(x[194]), .Q(
        xin[194]) );
  DFF \xreg_reg[195]  ( .D(xin[194]), .CLK(clk), .RST(start), .I(x[195]), .Q(
        xin[195]) );
  DFF \xreg_reg[196]  ( .D(xin[195]), .CLK(clk), .RST(start), .I(x[196]), .Q(
        xin[196]) );
  DFF \xreg_reg[197]  ( .D(xin[196]), .CLK(clk), .RST(start), .I(x[197]), .Q(
        xin[197]) );
  DFF \xreg_reg[198]  ( .D(xin[197]), .CLK(clk), .RST(start), .I(x[198]), .Q(
        xin[198]) );
  DFF \xreg_reg[199]  ( .D(xin[198]), .CLK(clk), .RST(start), .I(x[199]), .Q(
        xin[199]) );
  DFF \xreg_reg[200]  ( .D(xin[199]), .CLK(clk), .RST(start), .I(x[200]), .Q(
        xin[200]) );
  DFF \xreg_reg[201]  ( .D(xin[200]), .CLK(clk), .RST(start), .I(x[201]), .Q(
        xin[201]) );
  DFF \xreg_reg[202]  ( .D(xin[201]), .CLK(clk), .RST(start), .I(x[202]), .Q(
        xin[202]) );
  DFF \xreg_reg[203]  ( .D(xin[202]), .CLK(clk), .RST(start), .I(x[203]), .Q(
        xin[203]) );
  DFF \xreg_reg[204]  ( .D(xin[203]), .CLK(clk), .RST(start), .I(x[204]), .Q(
        xin[204]) );
  DFF \xreg_reg[205]  ( .D(xin[204]), .CLK(clk), .RST(start), .I(x[205]), .Q(
        xin[205]) );
  DFF \xreg_reg[206]  ( .D(xin[205]), .CLK(clk), .RST(start), .I(x[206]), .Q(
        xin[206]) );
  DFF \xreg_reg[207]  ( .D(xin[206]), .CLK(clk), .RST(start), .I(x[207]), .Q(
        xin[207]) );
  DFF \xreg_reg[208]  ( .D(xin[207]), .CLK(clk), .RST(start), .I(x[208]), .Q(
        xin[208]) );
  DFF \xreg_reg[209]  ( .D(xin[208]), .CLK(clk), .RST(start), .I(x[209]), .Q(
        xin[209]) );
  DFF \xreg_reg[210]  ( .D(xin[209]), .CLK(clk), .RST(start), .I(x[210]), .Q(
        xin[210]) );
  DFF \xreg_reg[211]  ( .D(xin[210]), .CLK(clk), .RST(start), .I(x[211]), .Q(
        xin[211]) );
  DFF \xreg_reg[212]  ( .D(xin[211]), .CLK(clk), .RST(start), .I(x[212]), .Q(
        xin[212]) );
  DFF \xreg_reg[213]  ( .D(xin[212]), .CLK(clk), .RST(start), .I(x[213]), .Q(
        xin[213]) );
  DFF \xreg_reg[214]  ( .D(xin[213]), .CLK(clk), .RST(start), .I(x[214]), .Q(
        xin[214]) );
  DFF \xreg_reg[215]  ( .D(xin[214]), .CLK(clk), .RST(start), .I(x[215]), .Q(
        xin[215]) );
  DFF \xreg_reg[216]  ( .D(xin[215]), .CLK(clk), .RST(start), .I(x[216]), .Q(
        xin[216]) );
  DFF \xreg_reg[217]  ( .D(xin[216]), .CLK(clk), .RST(start), .I(x[217]), .Q(
        xin[217]) );
  DFF \xreg_reg[218]  ( .D(xin[217]), .CLK(clk), .RST(start), .I(x[218]), .Q(
        xin[218]) );
  DFF \xreg_reg[219]  ( .D(xin[218]), .CLK(clk), .RST(start), .I(x[219]), .Q(
        xin[219]) );
  DFF \xreg_reg[220]  ( .D(xin[219]), .CLK(clk), .RST(start), .I(x[220]), .Q(
        xin[220]) );
  DFF \xreg_reg[221]  ( .D(xin[220]), .CLK(clk), .RST(start), .I(x[221]), .Q(
        xin[221]) );
  DFF \xreg_reg[222]  ( .D(xin[221]), .CLK(clk), .RST(start), .I(x[222]), .Q(
        xin[222]) );
  DFF \xreg_reg[223]  ( .D(xin[222]), .CLK(clk), .RST(start), .I(x[223]), .Q(
        xin[223]) );
  DFF \xreg_reg[224]  ( .D(xin[223]), .CLK(clk), .RST(start), .I(x[224]), .Q(
        xin[224]) );
  DFF \xreg_reg[225]  ( .D(xin[224]), .CLK(clk), .RST(start), .I(x[225]), .Q(
        xin[225]) );
  DFF \xreg_reg[226]  ( .D(xin[225]), .CLK(clk), .RST(start), .I(x[226]), .Q(
        xin[226]) );
  DFF \xreg_reg[227]  ( .D(xin[226]), .CLK(clk), .RST(start), .I(x[227]), .Q(
        xin[227]) );
  DFF \xreg_reg[228]  ( .D(xin[227]), .CLK(clk), .RST(start), .I(x[228]), .Q(
        xin[228]) );
  DFF \xreg_reg[229]  ( .D(xin[228]), .CLK(clk), .RST(start), .I(x[229]), .Q(
        xin[229]) );
  DFF \xreg_reg[230]  ( .D(xin[229]), .CLK(clk), .RST(start), .I(x[230]), .Q(
        xin[230]) );
  DFF \xreg_reg[231]  ( .D(xin[230]), .CLK(clk), .RST(start), .I(x[231]), .Q(
        xin[231]) );
  DFF \xreg_reg[232]  ( .D(xin[231]), .CLK(clk), .RST(start), .I(x[232]), .Q(
        xin[232]) );
  DFF \xreg_reg[233]  ( .D(xin[232]), .CLK(clk), .RST(start), .I(x[233]), .Q(
        xin[233]) );
  DFF \xreg_reg[234]  ( .D(xin[233]), .CLK(clk), .RST(start), .I(x[234]), .Q(
        xin[234]) );
  DFF \xreg_reg[235]  ( .D(xin[234]), .CLK(clk), .RST(start), .I(x[235]), .Q(
        xin[235]) );
  DFF \xreg_reg[236]  ( .D(xin[235]), .CLK(clk), .RST(start), .I(x[236]), .Q(
        xin[236]) );
  DFF \xreg_reg[237]  ( .D(xin[236]), .CLK(clk), .RST(start), .I(x[237]), .Q(
        xin[237]) );
  DFF \xreg_reg[238]  ( .D(xin[237]), .CLK(clk), .RST(start), .I(x[238]), .Q(
        xin[238]) );
  DFF \xreg_reg[239]  ( .D(xin[238]), .CLK(clk), .RST(start), .I(x[239]), .Q(
        xin[239]) );
  DFF \xreg_reg[240]  ( .D(xin[239]), .CLK(clk), .RST(start), .I(x[240]), .Q(
        xin[240]) );
  DFF \xreg_reg[241]  ( .D(xin[240]), .CLK(clk), .RST(start), .I(x[241]), .Q(
        xin[241]) );
  DFF \xreg_reg[242]  ( .D(xin[241]), .CLK(clk), .RST(start), .I(x[242]), .Q(
        xin[242]) );
  DFF \xreg_reg[243]  ( .D(xin[242]), .CLK(clk), .RST(start), .I(x[243]), .Q(
        xin[243]) );
  DFF \xreg_reg[244]  ( .D(xin[243]), .CLK(clk), .RST(start), .I(x[244]), .Q(
        xin[244]) );
  DFF \xreg_reg[245]  ( .D(xin[244]), .CLK(clk), .RST(start), .I(x[245]), .Q(
        xin[245]) );
  DFF \xreg_reg[246]  ( .D(xin[245]), .CLK(clk), .RST(start), .I(x[246]), .Q(
        xin[246]) );
  DFF \xreg_reg[247]  ( .D(xin[246]), .CLK(clk), .RST(start), .I(x[247]), .Q(
        xin[247]) );
  DFF \xreg_reg[248]  ( .D(xin[247]), .CLK(clk), .RST(start), .I(x[248]), .Q(
        xin[248]) );
  DFF \xreg_reg[249]  ( .D(xin[248]), .CLK(clk), .RST(start), .I(x[249]), .Q(
        xin[249]) );
  DFF \xreg_reg[250]  ( .D(xin[249]), .CLK(clk), .RST(start), .I(x[250]), .Q(
        xin[250]) );
  DFF \xreg_reg[251]  ( .D(xin[250]), .CLK(clk), .RST(start), .I(x[251]), .Q(
        xin[251]) );
  DFF \xreg_reg[252]  ( .D(xin[251]), .CLK(clk), .RST(start), .I(x[252]), .Q(
        xin[252]) );
  DFF \xreg_reg[253]  ( .D(xin[252]), .CLK(clk), .RST(start), .I(x[253]), .Q(
        xin[253]) );
  DFF \xreg_reg[254]  ( .D(xin[253]), .CLK(clk), .RST(start), .I(x[254]), .Q(
        xin[254]) );
  DFF \xreg_reg[255]  ( .D(xin[254]), .CLK(clk), .RST(start), .I(x[255]), .Q(
        xin[255]) );
  DFF \xreg_reg[256]  ( .D(xin[255]), .CLK(clk), .RST(start), .I(x[256]), .Q(
        xin[256]) );
  DFF \xreg_reg[257]  ( .D(xin[256]), .CLK(clk), .RST(start), .I(x[257]), .Q(
        xin[257]) );
  DFF \xreg_reg[258]  ( .D(xin[257]), .CLK(clk), .RST(start), .I(x[258]), .Q(
        xin[258]) );
  DFF \xreg_reg[259]  ( .D(xin[258]), .CLK(clk), .RST(start), .I(x[259]), .Q(
        xin[259]) );
  DFF \xreg_reg[260]  ( .D(xin[259]), .CLK(clk), .RST(start), .I(x[260]), .Q(
        xin[260]) );
  DFF \xreg_reg[261]  ( .D(xin[260]), .CLK(clk), .RST(start), .I(x[261]), .Q(
        xin[261]) );
  DFF \xreg_reg[262]  ( .D(xin[261]), .CLK(clk), .RST(start), .I(x[262]), .Q(
        xin[262]) );
  DFF \xreg_reg[263]  ( .D(xin[262]), .CLK(clk), .RST(start), .I(x[263]), .Q(
        xin[263]) );
  DFF \xreg_reg[264]  ( .D(xin[263]), .CLK(clk), .RST(start), .I(x[264]), .Q(
        xin[264]) );
  DFF \xreg_reg[265]  ( .D(xin[264]), .CLK(clk), .RST(start), .I(x[265]), .Q(
        xin[265]) );
  DFF \xreg_reg[266]  ( .D(xin[265]), .CLK(clk), .RST(start), .I(x[266]), .Q(
        xin[266]) );
  DFF \xreg_reg[267]  ( .D(xin[266]), .CLK(clk), .RST(start), .I(x[267]), .Q(
        xin[267]) );
  DFF \xreg_reg[268]  ( .D(xin[267]), .CLK(clk), .RST(start), .I(x[268]), .Q(
        xin[268]) );
  DFF \xreg_reg[269]  ( .D(xin[268]), .CLK(clk), .RST(start), .I(x[269]), .Q(
        xin[269]) );
  DFF \xreg_reg[270]  ( .D(xin[269]), .CLK(clk), .RST(start), .I(x[270]), .Q(
        xin[270]) );
  DFF \xreg_reg[271]  ( .D(xin[270]), .CLK(clk), .RST(start), .I(x[271]), .Q(
        xin[271]) );
  DFF \xreg_reg[272]  ( .D(xin[271]), .CLK(clk), .RST(start), .I(x[272]), .Q(
        xin[272]) );
  DFF \xreg_reg[273]  ( .D(xin[272]), .CLK(clk), .RST(start), .I(x[273]), .Q(
        xin[273]) );
  DFF \xreg_reg[274]  ( .D(xin[273]), .CLK(clk), .RST(start), .I(x[274]), .Q(
        xin[274]) );
  DFF \xreg_reg[275]  ( .D(xin[274]), .CLK(clk), .RST(start), .I(x[275]), .Q(
        xin[275]) );
  DFF \xreg_reg[276]  ( .D(xin[275]), .CLK(clk), .RST(start), .I(x[276]), .Q(
        xin[276]) );
  DFF \xreg_reg[277]  ( .D(xin[276]), .CLK(clk), .RST(start), .I(x[277]), .Q(
        xin[277]) );
  DFF \xreg_reg[278]  ( .D(xin[277]), .CLK(clk), .RST(start), .I(x[278]), .Q(
        xin[278]) );
  DFF \xreg_reg[279]  ( .D(xin[278]), .CLK(clk), .RST(start), .I(x[279]), .Q(
        xin[279]) );
  DFF \xreg_reg[280]  ( .D(xin[279]), .CLK(clk), .RST(start), .I(x[280]), .Q(
        xin[280]) );
  DFF \xreg_reg[281]  ( .D(xin[280]), .CLK(clk), .RST(start), .I(x[281]), .Q(
        xin[281]) );
  DFF \xreg_reg[282]  ( .D(xin[281]), .CLK(clk), .RST(start), .I(x[282]), .Q(
        xin[282]) );
  DFF \xreg_reg[283]  ( .D(xin[282]), .CLK(clk), .RST(start), .I(x[283]), .Q(
        xin[283]) );
  DFF \xreg_reg[284]  ( .D(xin[283]), .CLK(clk), .RST(start), .I(x[284]), .Q(
        xin[284]) );
  DFF \xreg_reg[285]  ( .D(xin[284]), .CLK(clk), .RST(start), .I(x[285]), .Q(
        xin[285]) );
  DFF \xreg_reg[286]  ( .D(xin[285]), .CLK(clk), .RST(start), .I(x[286]), .Q(
        xin[286]) );
  DFF \xreg_reg[287]  ( .D(xin[286]), .CLK(clk), .RST(start), .I(x[287]), .Q(
        xin[287]) );
  DFF \xreg_reg[288]  ( .D(xin[287]), .CLK(clk), .RST(start), .I(x[288]), .Q(
        xin[288]) );
  DFF \xreg_reg[289]  ( .D(xin[288]), .CLK(clk), .RST(start), .I(x[289]), .Q(
        xin[289]) );
  DFF \xreg_reg[290]  ( .D(xin[289]), .CLK(clk), .RST(start), .I(x[290]), .Q(
        xin[290]) );
  DFF \xreg_reg[291]  ( .D(xin[290]), .CLK(clk), .RST(start), .I(x[291]), .Q(
        xin[291]) );
  DFF \xreg_reg[292]  ( .D(xin[291]), .CLK(clk), .RST(start), .I(x[292]), .Q(
        xin[292]) );
  DFF \xreg_reg[293]  ( .D(xin[292]), .CLK(clk), .RST(start), .I(x[293]), .Q(
        xin[293]) );
  DFF \xreg_reg[294]  ( .D(xin[293]), .CLK(clk), .RST(start), .I(x[294]), .Q(
        xin[294]) );
  DFF \xreg_reg[295]  ( .D(xin[294]), .CLK(clk), .RST(start), .I(x[295]), .Q(
        xin[295]) );
  DFF \xreg_reg[296]  ( .D(xin[295]), .CLK(clk), .RST(start), .I(x[296]), .Q(
        xin[296]) );
  DFF \xreg_reg[297]  ( .D(xin[296]), .CLK(clk), .RST(start), .I(x[297]), .Q(
        xin[297]) );
  DFF \xreg_reg[298]  ( .D(xin[297]), .CLK(clk), .RST(start), .I(x[298]), .Q(
        xin[298]) );
  DFF \xreg_reg[299]  ( .D(xin[298]), .CLK(clk), .RST(start), .I(x[299]), .Q(
        xin[299]) );
  DFF \xreg_reg[300]  ( .D(xin[299]), .CLK(clk), .RST(start), .I(x[300]), .Q(
        xin[300]) );
  DFF \xreg_reg[301]  ( .D(xin[300]), .CLK(clk), .RST(start), .I(x[301]), .Q(
        xin[301]) );
  DFF \xreg_reg[302]  ( .D(xin[301]), .CLK(clk), .RST(start), .I(x[302]), .Q(
        xin[302]) );
  DFF \xreg_reg[303]  ( .D(xin[302]), .CLK(clk), .RST(start), .I(x[303]), .Q(
        xin[303]) );
  DFF \xreg_reg[304]  ( .D(xin[303]), .CLK(clk), .RST(start), .I(x[304]), .Q(
        xin[304]) );
  DFF \xreg_reg[305]  ( .D(xin[304]), .CLK(clk), .RST(start), .I(x[305]), .Q(
        xin[305]) );
  DFF \xreg_reg[306]  ( .D(xin[305]), .CLK(clk), .RST(start), .I(x[306]), .Q(
        xin[306]) );
  DFF \xreg_reg[307]  ( .D(xin[306]), .CLK(clk), .RST(start), .I(x[307]), .Q(
        xin[307]) );
  DFF \xreg_reg[308]  ( .D(xin[307]), .CLK(clk), .RST(start), .I(x[308]), .Q(
        xin[308]) );
  DFF \xreg_reg[309]  ( .D(xin[308]), .CLK(clk), .RST(start), .I(x[309]), .Q(
        xin[309]) );
  DFF \xreg_reg[310]  ( .D(xin[309]), .CLK(clk), .RST(start), .I(x[310]), .Q(
        xin[310]) );
  DFF \xreg_reg[311]  ( .D(xin[310]), .CLK(clk), .RST(start), .I(x[311]), .Q(
        xin[311]) );
  DFF \xreg_reg[312]  ( .D(xin[311]), .CLK(clk), .RST(start), .I(x[312]), .Q(
        xin[312]) );
  DFF \xreg_reg[313]  ( .D(xin[312]), .CLK(clk), .RST(start), .I(x[313]), .Q(
        xin[313]) );
  DFF \xreg_reg[314]  ( .D(xin[313]), .CLK(clk), .RST(start), .I(x[314]), .Q(
        xin[314]) );
  DFF \xreg_reg[315]  ( .D(xin[314]), .CLK(clk), .RST(start), .I(x[315]), .Q(
        xin[315]) );
  DFF \xreg_reg[316]  ( .D(xin[315]), .CLK(clk), .RST(start), .I(x[316]), .Q(
        xin[316]) );
  DFF \xreg_reg[317]  ( .D(xin[316]), .CLK(clk), .RST(start), .I(x[317]), .Q(
        xin[317]) );
  DFF \xreg_reg[318]  ( .D(xin[317]), .CLK(clk), .RST(start), .I(x[318]), .Q(
        xin[318]) );
  DFF \xreg_reg[319]  ( .D(xin[318]), .CLK(clk), .RST(start), .I(x[319]), .Q(
        xin[319]) );
  DFF \xreg_reg[320]  ( .D(xin[319]), .CLK(clk), .RST(start), .I(x[320]), .Q(
        xin[320]) );
  DFF \xreg_reg[321]  ( .D(xin[320]), .CLK(clk), .RST(start), .I(x[321]), .Q(
        xin[321]) );
  DFF \xreg_reg[322]  ( .D(xin[321]), .CLK(clk), .RST(start), .I(x[322]), .Q(
        xin[322]) );
  DFF \xreg_reg[323]  ( .D(xin[322]), .CLK(clk), .RST(start), .I(x[323]), .Q(
        xin[323]) );
  DFF \xreg_reg[324]  ( .D(xin[323]), .CLK(clk), .RST(start), .I(x[324]), .Q(
        xin[324]) );
  DFF \xreg_reg[325]  ( .D(xin[324]), .CLK(clk), .RST(start), .I(x[325]), .Q(
        xin[325]) );
  DFF \xreg_reg[326]  ( .D(xin[325]), .CLK(clk), .RST(start), .I(x[326]), .Q(
        xin[326]) );
  DFF \xreg_reg[327]  ( .D(xin[326]), .CLK(clk), .RST(start), .I(x[327]), .Q(
        xin[327]) );
  DFF \xreg_reg[328]  ( .D(xin[327]), .CLK(clk), .RST(start), .I(x[328]), .Q(
        xin[328]) );
  DFF \xreg_reg[329]  ( .D(xin[328]), .CLK(clk), .RST(start), .I(x[329]), .Q(
        xin[329]) );
  DFF \xreg_reg[330]  ( .D(xin[329]), .CLK(clk), .RST(start), .I(x[330]), .Q(
        xin[330]) );
  DFF \xreg_reg[331]  ( .D(xin[330]), .CLK(clk), .RST(start), .I(x[331]), .Q(
        xin[331]) );
  DFF \xreg_reg[332]  ( .D(xin[331]), .CLK(clk), .RST(start), .I(x[332]), .Q(
        xin[332]) );
  DFF \xreg_reg[333]  ( .D(xin[332]), .CLK(clk), .RST(start), .I(x[333]), .Q(
        xin[333]) );
  DFF \xreg_reg[334]  ( .D(xin[333]), .CLK(clk), .RST(start), .I(x[334]), .Q(
        xin[334]) );
  DFF \xreg_reg[335]  ( .D(xin[334]), .CLK(clk), .RST(start), .I(x[335]), .Q(
        xin[335]) );
  DFF \xreg_reg[336]  ( .D(xin[335]), .CLK(clk), .RST(start), .I(x[336]), .Q(
        xin[336]) );
  DFF \xreg_reg[337]  ( .D(xin[336]), .CLK(clk), .RST(start), .I(x[337]), .Q(
        xin[337]) );
  DFF \xreg_reg[338]  ( .D(xin[337]), .CLK(clk), .RST(start), .I(x[338]), .Q(
        xin[338]) );
  DFF \xreg_reg[339]  ( .D(xin[338]), .CLK(clk), .RST(start), .I(x[339]), .Q(
        xin[339]) );
  DFF \xreg_reg[340]  ( .D(xin[339]), .CLK(clk), .RST(start), .I(x[340]), .Q(
        xin[340]) );
  DFF \xreg_reg[341]  ( .D(xin[340]), .CLK(clk), .RST(start), .I(x[341]), .Q(
        xin[341]) );
  DFF \xreg_reg[342]  ( .D(xin[341]), .CLK(clk), .RST(start), .I(x[342]), .Q(
        xin[342]) );
  DFF \xreg_reg[343]  ( .D(xin[342]), .CLK(clk), .RST(start), .I(x[343]), .Q(
        xin[343]) );
  DFF \xreg_reg[344]  ( .D(xin[343]), .CLK(clk), .RST(start), .I(x[344]), .Q(
        xin[344]) );
  DFF \xreg_reg[345]  ( .D(xin[344]), .CLK(clk), .RST(start), .I(x[345]), .Q(
        xin[345]) );
  DFF \xreg_reg[346]  ( .D(xin[345]), .CLK(clk), .RST(start), .I(x[346]), .Q(
        xin[346]) );
  DFF \xreg_reg[347]  ( .D(xin[346]), .CLK(clk), .RST(start), .I(x[347]), .Q(
        xin[347]) );
  DFF \xreg_reg[348]  ( .D(xin[347]), .CLK(clk), .RST(start), .I(x[348]), .Q(
        xin[348]) );
  DFF \xreg_reg[349]  ( .D(xin[348]), .CLK(clk), .RST(start), .I(x[349]), .Q(
        xin[349]) );
  DFF \xreg_reg[350]  ( .D(xin[349]), .CLK(clk), .RST(start), .I(x[350]), .Q(
        xin[350]) );
  DFF \xreg_reg[351]  ( .D(xin[350]), .CLK(clk), .RST(start), .I(x[351]), .Q(
        xin[351]) );
  DFF \xreg_reg[352]  ( .D(xin[351]), .CLK(clk), .RST(start), .I(x[352]), .Q(
        xin[352]) );
  DFF \xreg_reg[353]  ( .D(xin[352]), .CLK(clk), .RST(start), .I(x[353]), .Q(
        xin[353]) );
  DFF \xreg_reg[354]  ( .D(xin[353]), .CLK(clk), .RST(start), .I(x[354]), .Q(
        xin[354]) );
  DFF \xreg_reg[355]  ( .D(xin[354]), .CLK(clk), .RST(start), .I(x[355]), .Q(
        xin[355]) );
  DFF \xreg_reg[356]  ( .D(xin[355]), .CLK(clk), .RST(start), .I(x[356]), .Q(
        xin[356]) );
  DFF \xreg_reg[357]  ( .D(xin[356]), .CLK(clk), .RST(start), .I(x[357]), .Q(
        xin[357]) );
  DFF \xreg_reg[358]  ( .D(xin[357]), .CLK(clk), .RST(start), .I(x[358]), .Q(
        xin[358]) );
  DFF \xreg_reg[359]  ( .D(xin[358]), .CLK(clk), .RST(start), .I(x[359]), .Q(
        xin[359]) );
  DFF \xreg_reg[360]  ( .D(xin[359]), .CLK(clk), .RST(start), .I(x[360]), .Q(
        xin[360]) );
  DFF \xreg_reg[361]  ( .D(xin[360]), .CLK(clk), .RST(start), .I(x[361]), .Q(
        xin[361]) );
  DFF \xreg_reg[362]  ( .D(xin[361]), .CLK(clk), .RST(start), .I(x[362]), .Q(
        xin[362]) );
  DFF \xreg_reg[363]  ( .D(xin[362]), .CLK(clk), .RST(start), .I(x[363]), .Q(
        xin[363]) );
  DFF \xreg_reg[364]  ( .D(xin[363]), .CLK(clk), .RST(start), .I(x[364]), .Q(
        xin[364]) );
  DFF \xreg_reg[365]  ( .D(xin[364]), .CLK(clk), .RST(start), .I(x[365]), .Q(
        xin[365]) );
  DFF \xreg_reg[366]  ( .D(xin[365]), .CLK(clk), .RST(start), .I(x[366]), .Q(
        xin[366]) );
  DFF \xreg_reg[367]  ( .D(xin[366]), .CLK(clk), .RST(start), .I(x[367]), .Q(
        xin[367]) );
  DFF \xreg_reg[368]  ( .D(xin[367]), .CLK(clk), .RST(start), .I(x[368]), .Q(
        xin[368]) );
  DFF \xreg_reg[369]  ( .D(xin[368]), .CLK(clk), .RST(start), .I(x[369]), .Q(
        xin[369]) );
  DFF \xreg_reg[370]  ( .D(xin[369]), .CLK(clk), .RST(start), .I(x[370]), .Q(
        xin[370]) );
  DFF \xreg_reg[371]  ( .D(xin[370]), .CLK(clk), .RST(start), .I(x[371]), .Q(
        xin[371]) );
  DFF \xreg_reg[372]  ( .D(xin[371]), .CLK(clk), .RST(start), .I(x[372]), .Q(
        xin[372]) );
  DFF \xreg_reg[373]  ( .D(xin[372]), .CLK(clk), .RST(start), .I(x[373]), .Q(
        xin[373]) );
  DFF \xreg_reg[374]  ( .D(xin[373]), .CLK(clk), .RST(start), .I(x[374]), .Q(
        xin[374]) );
  DFF \xreg_reg[375]  ( .D(xin[374]), .CLK(clk), .RST(start), .I(x[375]), .Q(
        xin[375]) );
  DFF \xreg_reg[376]  ( .D(xin[375]), .CLK(clk), .RST(start), .I(x[376]), .Q(
        xin[376]) );
  DFF \xreg_reg[377]  ( .D(xin[376]), .CLK(clk), .RST(start), .I(x[377]), .Q(
        xin[377]) );
  DFF \xreg_reg[378]  ( .D(xin[377]), .CLK(clk), .RST(start), .I(x[378]), .Q(
        xin[378]) );
  DFF \xreg_reg[379]  ( .D(xin[378]), .CLK(clk), .RST(start), .I(x[379]), .Q(
        xin[379]) );
  DFF \xreg_reg[380]  ( .D(xin[379]), .CLK(clk), .RST(start), .I(x[380]), .Q(
        xin[380]) );
  DFF \xreg_reg[381]  ( .D(xin[380]), .CLK(clk), .RST(start), .I(x[381]), .Q(
        xin[381]) );
  DFF \xreg_reg[382]  ( .D(xin[381]), .CLK(clk), .RST(start), .I(x[382]), .Q(
        xin[382]) );
  DFF \xreg_reg[383]  ( .D(xin[382]), .CLK(clk), .RST(start), .I(x[383]), .Q(
        xin[383]) );
  DFF \xreg_reg[384]  ( .D(xin[383]), .CLK(clk), .RST(start), .I(x[384]), .Q(
        xin[384]) );
  DFF \xreg_reg[385]  ( .D(xin[384]), .CLK(clk), .RST(start), .I(x[385]), .Q(
        xin[385]) );
  DFF \xreg_reg[386]  ( .D(xin[385]), .CLK(clk), .RST(start), .I(x[386]), .Q(
        xin[386]) );
  DFF \xreg_reg[387]  ( .D(xin[386]), .CLK(clk), .RST(start), .I(x[387]), .Q(
        xin[387]) );
  DFF \xreg_reg[388]  ( .D(xin[387]), .CLK(clk), .RST(start), .I(x[388]), .Q(
        xin[388]) );
  DFF \xreg_reg[389]  ( .D(xin[388]), .CLK(clk), .RST(start), .I(x[389]), .Q(
        xin[389]) );
  DFF \xreg_reg[390]  ( .D(xin[389]), .CLK(clk), .RST(start), .I(x[390]), .Q(
        xin[390]) );
  DFF \xreg_reg[391]  ( .D(xin[390]), .CLK(clk), .RST(start), .I(x[391]), .Q(
        xin[391]) );
  DFF \xreg_reg[392]  ( .D(xin[391]), .CLK(clk), .RST(start), .I(x[392]), .Q(
        xin[392]) );
  DFF \xreg_reg[393]  ( .D(xin[392]), .CLK(clk), .RST(start), .I(x[393]), .Q(
        xin[393]) );
  DFF \xreg_reg[394]  ( .D(xin[393]), .CLK(clk), .RST(start), .I(x[394]), .Q(
        xin[394]) );
  DFF \xreg_reg[395]  ( .D(xin[394]), .CLK(clk), .RST(start), .I(x[395]), .Q(
        xin[395]) );
  DFF \xreg_reg[396]  ( .D(xin[395]), .CLK(clk), .RST(start), .I(x[396]), .Q(
        xin[396]) );
  DFF \xreg_reg[397]  ( .D(xin[396]), .CLK(clk), .RST(start), .I(x[397]), .Q(
        xin[397]) );
  DFF \xreg_reg[398]  ( .D(xin[397]), .CLK(clk), .RST(start), .I(x[398]), .Q(
        xin[398]) );
  DFF \xreg_reg[399]  ( .D(xin[398]), .CLK(clk), .RST(start), .I(x[399]), .Q(
        xin[399]) );
  DFF \xreg_reg[400]  ( .D(xin[399]), .CLK(clk), .RST(start), .I(x[400]), .Q(
        xin[400]) );
  DFF \xreg_reg[401]  ( .D(xin[400]), .CLK(clk), .RST(start), .I(x[401]), .Q(
        xin[401]) );
  DFF \xreg_reg[402]  ( .D(xin[401]), .CLK(clk), .RST(start), .I(x[402]), .Q(
        xin[402]) );
  DFF \xreg_reg[403]  ( .D(xin[402]), .CLK(clk), .RST(start), .I(x[403]), .Q(
        xin[403]) );
  DFF \xreg_reg[404]  ( .D(xin[403]), .CLK(clk), .RST(start), .I(x[404]), .Q(
        xin[404]) );
  DFF \xreg_reg[405]  ( .D(xin[404]), .CLK(clk), .RST(start), .I(x[405]), .Q(
        xin[405]) );
  DFF \xreg_reg[406]  ( .D(xin[405]), .CLK(clk), .RST(start), .I(x[406]), .Q(
        xin[406]) );
  DFF \xreg_reg[407]  ( .D(xin[406]), .CLK(clk), .RST(start), .I(x[407]), .Q(
        xin[407]) );
  DFF \xreg_reg[408]  ( .D(xin[407]), .CLK(clk), .RST(start), .I(x[408]), .Q(
        xin[408]) );
  DFF \xreg_reg[409]  ( .D(xin[408]), .CLK(clk), .RST(start), .I(x[409]), .Q(
        xin[409]) );
  DFF \xreg_reg[410]  ( .D(xin[409]), .CLK(clk), .RST(start), .I(x[410]), .Q(
        xin[410]) );
  DFF \xreg_reg[411]  ( .D(xin[410]), .CLK(clk), .RST(start), .I(x[411]), .Q(
        xin[411]) );
  DFF \xreg_reg[412]  ( .D(xin[411]), .CLK(clk), .RST(start), .I(x[412]), .Q(
        xin[412]) );
  DFF \xreg_reg[413]  ( .D(xin[412]), .CLK(clk), .RST(start), .I(x[413]), .Q(
        xin[413]) );
  DFF \xreg_reg[414]  ( .D(xin[413]), .CLK(clk), .RST(start), .I(x[414]), .Q(
        xin[414]) );
  DFF \xreg_reg[415]  ( .D(xin[414]), .CLK(clk), .RST(start), .I(x[415]), .Q(
        xin[415]) );
  DFF \xreg_reg[416]  ( .D(xin[415]), .CLK(clk), .RST(start), .I(x[416]), .Q(
        xin[416]) );
  DFF \xreg_reg[417]  ( .D(xin[416]), .CLK(clk), .RST(start), .I(x[417]), .Q(
        xin[417]) );
  DFF \xreg_reg[418]  ( .D(xin[417]), .CLK(clk), .RST(start), .I(x[418]), .Q(
        xin[418]) );
  DFF \xreg_reg[419]  ( .D(xin[418]), .CLK(clk), .RST(start), .I(x[419]), .Q(
        xin[419]) );
  DFF \xreg_reg[420]  ( .D(xin[419]), .CLK(clk), .RST(start), .I(x[420]), .Q(
        xin[420]) );
  DFF \xreg_reg[421]  ( .D(xin[420]), .CLK(clk), .RST(start), .I(x[421]), .Q(
        xin[421]) );
  DFF \xreg_reg[422]  ( .D(xin[421]), .CLK(clk), .RST(start), .I(x[422]), .Q(
        xin[422]) );
  DFF \xreg_reg[423]  ( .D(xin[422]), .CLK(clk), .RST(start), .I(x[423]), .Q(
        xin[423]) );
  DFF \xreg_reg[424]  ( .D(xin[423]), .CLK(clk), .RST(start), .I(x[424]), .Q(
        xin[424]) );
  DFF \xreg_reg[425]  ( .D(xin[424]), .CLK(clk), .RST(start), .I(x[425]), .Q(
        xin[425]) );
  DFF \xreg_reg[426]  ( .D(xin[425]), .CLK(clk), .RST(start), .I(x[426]), .Q(
        xin[426]) );
  DFF \xreg_reg[427]  ( .D(xin[426]), .CLK(clk), .RST(start), .I(x[427]), .Q(
        xin[427]) );
  DFF \xreg_reg[428]  ( .D(xin[427]), .CLK(clk), .RST(start), .I(x[428]), .Q(
        xin[428]) );
  DFF \xreg_reg[429]  ( .D(xin[428]), .CLK(clk), .RST(start), .I(x[429]), .Q(
        xin[429]) );
  DFF \xreg_reg[430]  ( .D(xin[429]), .CLK(clk), .RST(start), .I(x[430]), .Q(
        xin[430]) );
  DFF \xreg_reg[431]  ( .D(xin[430]), .CLK(clk), .RST(start), .I(x[431]), .Q(
        xin[431]) );
  DFF \xreg_reg[432]  ( .D(xin[431]), .CLK(clk), .RST(start), .I(x[432]), .Q(
        xin[432]) );
  DFF \xreg_reg[433]  ( .D(xin[432]), .CLK(clk), .RST(start), .I(x[433]), .Q(
        xin[433]) );
  DFF \xreg_reg[434]  ( .D(xin[433]), .CLK(clk), .RST(start), .I(x[434]), .Q(
        xin[434]) );
  DFF \xreg_reg[435]  ( .D(xin[434]), .CLK(clk), .RST(start), .I(x[435]), .Q(
        xin[435]) );
  DFF \xreg_reg[436]  ( .D(xin[435]), .CLK(clk), .RST(start), .I(x[436]), .Q(
        xin[436]) );
  DFF \xreg_reg[437]  ( .D(xin[436]), .CLK(clk), .RST(start), .I(x[437]), .Q(
        xin[437]) );
  DFF \xreg_reg[438]  ( .D(xin[437]), .CLK(clk), .RST(start), .I(x[438]), .Q(
        xin[438]) );
  DFF \xreg_reg[439]  ( .D(xin[438]), .CLK(clk), .RST(start), .I(x[439]), .Q(
        xin[439]) );
  DFF \xreg_reg[440]  ( .D(xin[439]), .CLK(clk), .RST(start), .I(x[440]), .Q(
        xin[440]) );
  DFF \xreg_reg[441]  ( .D(xin[440]), .CLK(clk), .RST(start), .I(x[441]), .Q(
        xin[441]) );
  DFF \xreg_reg[442]  ( .D(xin[441]), .CLK(clk), .RST(start), .I(x[442]), .Q(
        xin[442]) );
  DFF \xreg_reg[443]  ( .D(xin[442]), .CLK(clk), .RST(start), .I(x[443]), .Q(
        xin[443]) );
  DFF \xreg_reg[444]  ( .D(xin[443]), .CLK(clk), .RST(start), .I(x[444]), .Q(
        xin[444]) );
  DFF \xreg_reg[445]  ( .D(xin[444]), .CLK(clk), .RST(start), .I(x[445]), .Q(
        xin[445]) );
  DFF \xreg_reg[446]  ( .D(xin[445]), .CLK(clk), .RST(start), .I(x[446]), .Q(
        xin[446]) );
  DFF \xreg_reg[447]  ( .D(xin[446]), .CLK(clk), .RST(start), .I(x[447]), .Q(
        xin[447]) );
  DFF \xreg_reg[448]  ( .D(xin[447]), .CLK(clk), .RST(start), .I(x[448]), .Q(
        xin[448]) );
  DFF \xreg_reg[449]  ( .D(xin[448]), .CLK(clk), .RST(start), .I(x[449]), .Q(
        xin[449]) );
  DFF \xreg_reg[450]  ( .D(xin[449]), .CLK(clk), .RST(start), .I(x[450]), .Q(
        xin[450]) );
  DFF \xreg_reg[451]  ( .D(xin[450]), .CLK(clk), .RST(start), .I(x[451]), .Q(
        xin[451]) );
  DFF \xreg_reg[452]  ( .D(xin[451]), .CLK(clk), .RST(start), .I(x[452]), .Q(
        xin[452]) );
  DFF \xreg_reg[453]  ( .D(xin[452]), .CLK(clk), .RST(start), .I(x[453]), .Q(
        xin[453]) );
  DFF \xreg_reg[454]  ( .D(xin[453]), .CLK(clk), .RST(start), .I(x[454]), .Q(
        xin[454]) );
  DFF \xreg_reg[455]  ( .D(xin[454]), .CLK(clk), .RST(start), .I(x[455]), .Q(
        xin[455]) );
  DFF \xreg_reg[456]  ( .D(xin[455]), .CLK(clk), .RST(start), .I(x[456]), .Q(
        xin[456]) );
  DFF \xreg_reg[457]  ( .D(xin[456]), .CLK(clk), .RST(start), .I(x[457]), .Q(
        xin[457]) );
  DFF \xreg_reg[458]  ( .D(xin[457]), .CLK(clk), .RST(start), .I(x[458]), .Q(
        xin[458]) );
  DFF \xreg_reg[459]  ( .D(xin[458]), .CLK(clk), .RST(start), .I(x[459]), .Q(
        xin[459]) );
  DFF \xreg_reg[460]  ( .D(xin[459]), .CLK(clk), .RST(start), .I(x[460]), .Q(
        xin[460]) );
  DFF \xreg_reg[461]  ( .D(xin[460]), .CLK(clk), .RST(start), .I(x[461]), .Q(
        xin[461]) );
  DFF \xreg_reg[462]  ( .D(xin[461]), .CLK(clk), .RST(start), .I(x[462]), .Q(
        xin[462]) );
  DFF \xreg_reg[463]  ( .D(xin[462]), .CLK(clk), .RST(start), .I(x[463]), .Q(
        xin[463]) );
  DFF \xreg_reg[464]  ( .D(xin[463]), .CLK(clk), .RST(start), .I(x[464]), .Q(
        xin[464]) );
  DFF \xreg_reg[465]  ( .D(xin[464]), .CLK(clk), .RST(start), .I(x[465]), .Q(
        xin[465]) );
  DFF \xreg_reg[466]  ( .D(xin[465]), .CLK(clk), .RST(start), .I(x[466]), .Q(
        xin[466]) );
  DFF \xreg_reg[467]  ( .D(xin[466]), .CLK(clk), .RST(start), .I(x[467]), .Q(
        xin[467]) );
  DFF \xreg_reg[468]  ( .D(xin[467]), .CLK(clk), .RST(start), .I(x[468]), .Q(
        xin[468]) );
  DFF \xreg_reg[469]  ( .D(xin[468]), .CLK(clk), .RST(start), .I(x[469]), .Q(
        xin[469]) );
  DFF \xreg_reg[470]  ( .D(xin[469]), .CLK(clk), .RST(start), .I(x[470]), .Q(
        xin[470]) );
  DFF \xreg_reg[471]  ( .D(xin[470]), .CLK(clk), .RST(start), .I(x[471]), .Q(
        xin[471]) );
  DFF \xreg_reg[472]  ( .D(xin[471]), .CLK(clk), .RST(start), .I(x[472]), .Q(
        xin[472]) );
  DFF \xreg_reg[473]  ( .D(xin[472]), .CLK(clk), .RST(start), .I(x[473]), .Q(
        xin[473]) );
  DFF \xreg_reg[474]  ( .D(xin[473]), .CLK(clk), .RST(start), .I(x[474]), .Q(
        xin[474]) );
  DFF \xreg_reg[475]  ( .D(xin[474]), .CLK(clk), .RST(start), .I(x[475]), .Q(
        xin[475]) );
  DFF \xreg_reg[476]  ( .D(xin[475]), .CLK(clk), .RST(start), .I(x[476]), .Q(
        xin[476]) );
  DFF \xreg_reg[477]  ( .D(xin[476]), .CLK(clk), .RST(start), .I(x[477]), .Q(
        xin[477]) );
  DFF \xreg_reg[478]  ( .D(xin[477]), .CLK(clk), .RST(start), .I(x[478]), .Q(
        xin[478]) );
  DFF \xreg_reg[479]  ( .D(xin[478]), .CLK(clk), .RST(start), .I(x[479]), .Q(
        xin[479]) );
  DFF \xreg_reg[480]  ( .D(xin[479]), .CLK(clk), .RST(start), .I(x[480]), .Q(
        xin[480]) );
  DFF \xreg_reg[481]  ( .D(xin[480]), .CLK(clk), .RST(start), .I(x[481]), .Q(
        xin[481]) );
  DFF \xreg_reg[482]  ( .D(xin[481]), .CLK(clk), .RST(start), .I(x[482]), .Q(
        xin[482]) );
  DFF \xreg_reg[483]  ( .D(xin[482]), .CLK(clk), .RST(start), .I(x[483]), .Q(
        xin[483]) );
  DFF \xreg_reg[484]  ( .D(xin[483]), .CLK(clk), .RST(start), .I(x[484]), .Q(
        xin[484]) );
  DFF \xreg_reg[485]  ( .D(xin[484]), .CLK(clk), .RST(start), .I(x[485]), .Q(
        xin[485]) );
  DFF \xreg_reg[486]  ( .D(xin[485]), .CLK(clk), .RST(start), .I(x[486]), .Q(
        xin[486]) );
  DFF \xreg_reg[487]  ( .D(xin[486]), .CLK(clk), .RST(start), .I(x[487]), .Q(
        xin[487]) );
  DFF \xreg_reg[488]  ( .D(xin[487]), .CLK(clk), .RST(start), .I(x[488]), .Q(
        xin[488]) );
  DFF \xreg_reg[489]  ( .D(xin[488]), .CLK(clk), .RST(start), .I(x[489]), .Q(
        xin[489]) );
  DFF \xreg_reg[490]  ( .D(xin[489]), .CLK(clk), .RST(start), .I(x[490]), .Q(
        xin[490]) );
  DFF \xreg_reg[491]  ( .D(xin[490]), .CLK(clk), .RST(start), .I(x[491]), .Q(
        xin[491]) );
  DFF \xreg_reg[492]  ( .D(xin[491]), .CLK(clk), .RST(start), .I(x[492]), .Q(
        xin[492]) );
  DFF \xreg_reg[493]  ( .D(xin[492]), .CLK(clk), .RST(start), .I(x[493]), .Q(
        xin[493]) );
  DFF \xreg_reg[494]  ( .D(xin[493]), .CLK(clk), .RST(start), .I(x[494]), .Q(
        xin[494]) );
  DFF \xreg_reg[495]  ( .D(xin[494]), .CLK(clk), .RST(start), .I(x[495]), .Q(
        xin[495]) );
  DFF \xreg_reg[496]  ( .D(xin[495]), .CLK(clk), .RST(start), .I(x[496]), .Q(
        xin[496]) );
  DFF \xreg_reg[497]  ( .D(xin[496]), .CLK(clk), .RST(start), .I(x[497]), .Q(
        xin[497]) );
  DFF \xreg_reg[498]  ( .D(xin[497]), .CLK(clk), .RST(start), .I(x[498]), .Q(
        xin[498]) );
  DFF \xreg_reg[499]  ( .D(xin[498]), .CLK(clk), .RST(start), .I(x[499]), .Q(
        xin[499]) );
  DFF \xreg_reg[500]  ( .D(xin[499]), .CLK(clk), .RST(start), .I(x[500]), .Q(
        xin[500]) );
  DFF \xreg_reg[501]  ( .D(xin[500]), .CLK(clk), .RST(start), .I(x[501]), .Q(
        xin[501]) );
  DFF \xreg_reg[502]  ( .D(xin[501]), .CLK(clk), .RST(start), .I(x[502]), .Q(
        xin[502]) );
  DFF \xreg_reg[503]  ( .D(xin[502]), .CLK(clk), .RST(start), .I(x[503]), .Q(
        xin[503]) );
  DFF \xreg_reg[504]  ( .D(xin[503]), .CLK(clk), .RST(start), .I(x[504]), .Q(
        xin[504]) );
  DFF \xreg_reg[505]  ( .D(xin[504]), .CLK(clk), .RST(start), .I(x[505]), .Q(
        xin[505]) );
  DFF \xreg_reg[506]  ( .D(xin[505]), .CLK(clk), .RST(start), .I(x[506]), .Q(
        xin[506]) );
  DFF \xreg_reg[507]  ( .D(xin[506]), .CLK(clk), .RST(start), .I(x[507]), .Q(
        xin[507]) );
  DFF \xreg_reg[508]  ( .D(xin[507]), .CLK(clk), .RST(start), .I(x[508]), .Q(
        xin[508]) );
  DFF \xreg_reg[509]  ( .D(xin[508]), .CLK(clk), .RST(start), .I(x[509]), .Q(
        xin[509]) );
  DFF \xreg_reg[510]  ( .D(xin[509]), .CLK(clk), .RST(start), .I(x[510]), .Q(
        xin[510]) );
  DFF \xreg_reg[511]  ( .D(xin[510]), .CLK(clk), .RST(start), .I(x[511]), .Q(
        xin[511]) );
  DFF \xreg_reg[512]  ( .D(xin[511]), .CLK(clk), .RST(start), .I(x[512]), .Q(
        xin[512]) );
  DFF \xreg_reg[513]  ( .D(xin[512]), .CLK(clk), .RST(start), .I(x[513]), .Q(
        xin[513]) );
  DFF \xreg_reg[514]  ( .D(xin[513]), .CLK(clk), .RST(start), .I(x[514]), .Q(
        xin[514]) );
  DFF \xreg_reg[515]  ( .D(xin[514]), .CLK(clk), .RST(start), .I(x[515]), .Q(
        xin[515]) );
  DFF \xreg_reg[516]  ( .D(xin[515]), .CLK(clk), .RST(start), .I(x[516]), .Q(
        xin[516]) );
  DFF \xreg_reg[517]  ( .D(xin[516]), .CLK(clk), .RST(start), .I(x[517]), .Q(
        xin[517]) );
  DFF \xreg_reg[518]  ( .D(xin[517]), .CLK(clk), .RST(start), .I(x[518]), .Q(
        xin[518]) );
  DFF \xreg_reg[519]  ( .D(xin[518]), .CLK(clk), .RST(start), .I(x[519]), .Q(
        xin[519]) );
  DFF \xreg_reg[520]  ( .D(xin[519]), .CLK(clk), .RST(start), .I(x[520]), .Q(
        xin[520]) );
  DFF \xreg_reg[521]  ( .D(xin[520]), .CLK(clk), .RST(start), .I(x[521]), .Q(
        xin[521]) );
  DFF \xreg_reg[522]  ( .D(xin[521]), .CLK(clk), .RST(start), .I(x[522]), .Q(
        xin[522]) );
  DFF \xreg_reg[523]  ( .D(xin[522]), .CLK(clk), .RST(start), .I(x[523]), .Q(
        xin[523]) );
  DFF \xreg_reg[524]  ( .D(xin[523]), .CLK(clk), .RST(start), .I(x[524]), .Q(
        xin[524]) );
  DFF \xreg_reg[525]  ( .D(xin[524]), .CLK(clk), .RST(start), .I(x[525]), .Q(
        xin[525]) );
  DFF \xreg_reg[526]  ( .D(xin[525]), .CLK(clk), .RST(start), .I(x[526]), .Q(
        xin[526]) );
  DFF \xreg_reg[527]  ( .D(xin[526]), .CLK(clk), .RST(start), .I(x[527]), .Q(
        xin[527]) );
  DFF \xreg_reg[528]  ( .D(xin[527]), .CLK(clk), .RST(start), .I(x[528]), .Q(
        xin[528]) );
  DFF \xreg_reg[529]  ( .D(xin[528]), .CLK(clk), .RST(start), .I(x[529]), .Q(
        xin[529]) );
  DFF \xreg_reg[530]  ( .D(xin[529]), .CLK(clk), .RST(start), .I(x[530]), .Q(
        xin[530]) );
  DFF \xreg_reg[531]  ( .D(xin[530]), .CLK(clk), .RST(start), .I(x[531]), .Q(
        xin[531]) );
  DFF \xreg_reg[532]  ( .D(xin[531]), .CLK(clk), .RST(start), .I(x[532]), .Q(
        xin[532]) );
  DFF \xreg_reg[533]  ( .D(xin[532]), .CLK(clk), .RST(start), .I(x[533]), .Q(
        xin[533]) );
  DFF \xreg_reg[534]  ( .D(xin[533]), .CLK(clk), .RST(start), .I(x[534]), .Q(
        xin[534]) );
  DFF \xreg_reg[535]  ( .D(xin[534]), .CLK(clk), .RST(start), .I(x[535]), .Q(
        xin[535]) );
  DFF \xreg_reg[536]  ( .D(xin[535]), .CLK(clk), .RST(start), .I(x[536]), .Q(
        xin[536]) );
  DFF \xreg_reg[537]  ( .D(xin[536]), .CLK(clk), .RST(start), .I(x[537]), .Q(
        xin[537]) );
  DFF \xreg_reg[538]  ( .D(xin[537]), .CLK(clk), .RST(start), .I(x[538]), .Q(
        xin[538]) );
  DFF \xreg_reg[539]  ( .D(xin[538]), .CLK(clk), .RST(start), .I(x[539]), .Q(
        xin[539]) );
  DFF \xreg_reg[540]  ( .D(xin[539]), .CLK(clk), .RST(start), .I(x[540]), .Q(
        xin[540]) );
  DFF \xreg_reg[541]  ( .D(xin[540]), .CLK(clk), .RST(start), .I(x[541]), .Q(
        xin[541]) );
  DFF \xreg_reg[542]  ( .D(xin[541]), .CLK(clk), .RST(start), .I(x[542]), .Q(
        xin[542]) );
  DFF \xreg_reg[543]  ( .D(xin[542]), .CLK(clk), .RST(start), .I(x[543]), .Q(
        xin[543]) );
  DFF \xreg_reg[544]  ( .D(xin[543]), .CLK(clk), .RST(start), .I(x[544]), .Q(
        xin[544]) );
  DFF \xreg_reg[545]  ( .D(xin[544]), .CLK(clk), .RST(start), .I(x[545]), .Q(
        xin[545]) );
  DFF \xreg_reg[546]  ( .D(xin[545]), .CLK(clk), .RST(start), .I(x[546]), .Q(
        xin[546]) );
  DFF \xreg_reg[547]  ( .D(xin[546]), .CLK(clk), .RST(start), .I(x[547]), .Q(
        xin[547]) );
  DFF \xreg_reg[548]  ( .D(xin[547]), .CLK(clk), .RST(start), .I(x[548]), .Q(
        xin[548]) );
  DFF \xreg_reg[549]  ( .D(xin[548]), .CLK(clk), .RST(start), .I(x[549]), .Q(
        xin[549]) );
  DFF \xreg_reg[550]  ( .D(xin[549]), .CLK(clk), .RST(start), .I(x[550]), .Q(
        xin[550]) );
  DFF \xreg_reg[551]  ( .D(xin[550]), .CLK(clk), .RST(start), .I(x[551]), .Q(
        xin[551]) );
  DFF \xreg_reg[552]  ( .D(xin[551]), .CLK(clk), .RST(start), .I(x[552]), .Q(
        xin[552]) );
  DFF \xreg_reg[553]  ( .D(xin[552]), .CLK(clk), .RST(start), .I(x[553]), .Q(
        xin[553]) );
  DFF \xreg_reg[554]  ( .D(xin[553]), .CLK(clk), .RST(start), .I(x[554]), .Q(
        xin[554]) );
  DFF \xreg_reg[555]  ( .D(xin[554]), .CLK(clk), .RST(start), .I(x[555]), .Q(
        xin[555]) );
  DFF \xreg_reg[556]  ( .D(xin[555]), .CLK(clk), .RST(start), .I(x[556]), .Q(
        xin[556]) );
  DFF \xreg_reg[557]  ( .D(xin[556]), .CLK(clk), .RST(start), .I(x[557]), .Q(
        xin[557]) );
  DFF \xreg_reg[558]  ( .D(xin[557]), .CLK(clk), .RST(start), .I(x[558]), .Q(
        xin[558]) );
  DFF \xreg_reg[559]  ( .D(xin[558]), .CLK(clk), .RST(start), .I(x[559]), .Q(
        xin[559]) );
  DFF \xreg_reg[560]  ( .D(xin[559]), .CLK(clk), .RST(start), .I(x[560]), .Q(
        xin[560]) );
  DFF \xreg_reg[561]  ( .D(xin[560]), .CLK(clk), .RST(start), .I(x[561]), .Q(
        xin[561]) );
  DFF \xreg_reg[562]  ( .D(xin[561]), .CLK(clk), .RST(start), .I(x[562]), .Q(
        xin[562]) );
  DFF \xreg_reg[563]  ( .D(xin[562]), .CLK(clk), .RST(start), .I(x[563]), .Q(
        xin[563]) );
  DFF \xreg_reg[564]  ( .D(xin[563]), .CLK(clk), .RST(start), .I(x[564]), .Q(
        xin[564]) );
  DFF \xreg_reg[565]  ( .D(xin[564]), .CLK(clk), .RST(start), .I(x[565]), .Q(
        xin[565]) );
  DFF \xreg_reg[566]  ( .D(xin[565]), .CLK(clk), .RST(start), .I(x[566]), .Q(
        xin[566]) );
  DFF \xreg_reg[567]  ( .D(xin[566]), .CLK(clk), .RST(start), .I(x[567]), .Q(
        xin[567]) );
  DFF \xreg_reg[568]  ( .D(xin[567]), .CLK(clk), .RST(start), .I(x[568]), .Q(
        xin[568]) );
  DFF \xreg_reg[569]  ( .D(xin[568]), .CLK(clk), .RST(start), .I(x[569]), .Q(
        xin[569]) );
  DFF \xreg_reg[570]  ( .D(xin[569]), .CLK(clk), .RST(start), .I(x[570]), .Q(
        xin[570]) );
  DFF \xreg_reg[571]  ( .D(xin[570]), .CLK(clk), .RST(start), .I(x[571]), .Q(
        xin[571]) );
  DFF \xreg_reg[572]  ( .D(xin[571]), .CLK(clk), .RST(start), .I(x[572]), .Q(
        xin[572]) );
  DFF \xreg_reg[573]  ( .D(xin[572]), .CLK(clk), .RST(start), .I(x[573]), .Q(
        xin[573]) );
  DFF \xreg_reg[574]  ( .D(xin[573]), .CLK(clk), .RST(start), .I(x[574]), .Q(
        xin[574]) );
  DFF \xreg_reg[575]  ( .D(xin[574]), .CLK(clk), .RST(start), .I(x[575]), .Q(
        xin[575]) );
  DFF \xreg_reg[576]  ( .D(xin[575]), .CLK(clk), .RST(start), .I(x[576]), .Q(
        xin[576]) );
  DFF \xreg_reg[577]  ( .D(xin[576]), .CLK(clk), .RST(start), .I(x[577]), .Q(
        xin[577]) );
  DFF \xreg_reg[578]  ( .D(xin[577]), .CLK(clk), .RST(start), .I(x[578]), .Q(
        xin[578]) );
  DFF \xreg_reg[579]  ( .D(xin[578]), .CLK(clk), .RST(start), .I(x[579]), .Q(
        xin[579]) );
  DFF \xreg_reg[580]  ( .D(xin[579]), .CLK(clk), .RST(start), .I(x[580]), .Q(
        xin[580]) );
  DFF \xreg_reg[581]  ( .D(xin[580]), .CLK(clk), .RST(start), .I(x[581]), .Q(
        xin[581]) );
  DFF \xreg_reg[582]  ( .D(xin[581]), .CLK(clk), .RST(start), .I(x[582]), .Q(
        xin[582]) );
  DFF \xreg_reg[583]  ( .D(xin[582]), .CLK(clk), .RST(start), .I(x[583]), .Q(
        xin[583]) );
  DFF \xreg_reg[584]  ( .D(xin[583]), .CLK(clk), .RST(start), .I(x[584]), .Q(
        xin[584]) );
  DFF \xreg_reg[585]  ( .D(xin[584]), .CLK(clk), .RST(start), .I(x[585]), .Q(
        xin[585]) );
  DFF \xreg_reg[586]  ( .D(xin[585]), .CLK(clk), .RST(start), .I(x[586]), .Q(
        xin[586]) );
  DFF \xreg_reg[587]  ( .D(xin[586]), .CLK(clk), .RST(start), .I(x[587]), .Q(
        xin[587]) );
  DFF \xreg_reg[588]  ( .D(xin[587]), .CLK(clk), .RST(start), .I(x[588]), .Q(
        xin[588]) );
  DFF \xreg_reg[589]  ( .D(xin[588]), .CLK(clk), .RST(start), .I(x[589]), .Q(
        xin[589]) );
  DFF \xreg_reg[590]  ( .D(xin[589]), .CLK(clk), .RST(start), .I(x[590]), .Q(
        xin[590]) );
  DFF \xreg_reg[591]  ( .D(xin[590]), .CLK(clk), .RST(start), .I(x[591]), .Q(
        xin[591]) );
  DFF \xreg_reg[592]  ( .D(xin[591]), .CLK(clk), .RST(start), .I(x[592]), .Q(
        xin[592]) );
  DFF \xreg_reg[593]  ( .D(xin[592]), .CLK(clk), .RST(start), .I(x[593]), .Q(
        xin[593]) );
  DFF \xreg_reg[594]  ( .D(xin[593]), .CLK(clk), .RST(start), .I(x[594]), .Q(
        xin[594]) );
  DFF \xreg_reg[595]  ( .D(xin[594]), .CLK(clk), .RST(start), .I(x[595]), .Q(
        xin[595]) );
  DFF \xreg_reg[596]  ( .D(xin[595]), .CLK(clk), .RST(start), .I(x[596]), .Q(
        xin[596]) );
  DFF \xreg_reg[597]  ( .D(xin[596]), .CLK(clk), .RST(start), .I(x[597]), .Q(
        xin[597]) );
  DFF \xreg_reg[598]  ( .D(xin[597]), .CLK(clk), .RST(start), .I(x[598]), .Q(
        xin[598]) );
  DFF \xreg_reg[599]  ( .D(xin[598]), .CLK(clk), .RST(start), .I(x[599]), .Q(
        xin[599]) );
  DFF \xreg_reg[600]  ( .D(xin[599]), .CLK(clk), .RST(start), .I(x[600]), .Q(
        xin[600]) );
  DFF \xreg_reg[601]  ( .D(xin[600]), .CLK(clk), .RST(start), .I(x[601]), .Q(
        xin[601]) );
  DFF \xreg_reg[602]  ( .D(xin[601]), .CLK(clk), .RST(start), .I(x[602]), .Q(
        xin[602]) );
  DFF \xreg_reg[603]  ( .D(xin[602]), .CLK(clk), .RST(start), .I(x[603]), .Q(
        xin[603]) );
  DFF \xreg_reg[604]  ( .D(xin[603]), .CLK(clk), .RST(start), .I(x[604]), .Q(
        xin[604]) );
  DFF \xreg_reg[605]  ( .D(xin[604]), .CLK(clk), .RST(start), .I(x[605]), .Q(
        xin[605]) );
  DFF \xreg_reg[606]  ( .D(xin[605]), .CLK(clk), .RST(start), .I(x[606]), .Q(
        xin[606]) );
  DFF \xreg_reg[607]  ( .D(xin[606]), .CLK(clk), .RST(start), .I(x[607]), .Q(
        xin[607]) );
  DFF \xreg_reg[608]  ( .D(xin[607]), .CLK(clk), .RST(start), .I(x[608]), .Q(
        xin[608]) );
  DFF \xreg_reg[609]  ( .D(xin[608]), .CLK(clk), .RST(start), .I(x[609]), .Q(
        xin[609]) );
  DFF \xreg_reg[610]  ( .D(xin[609]), .CLK(clk), .RST(start), .I(x[610]), .Q(
        xin[610]) );
  DFF \xreg_reg[611]  ( .D(xin[610]), .CLK(clk), .RST(start), .I(x[611]), .Q(
        xin[611]) );
  DFF \xreg_reg[612]  ( .D(xin[611]), .CLK(clk), .RST(start), .I(x[612]), .Q(
        xin[612]) );
  DFF \xreg_reg[613]  ( .D(xin[612]), .CLK(clk), .RST(start), .I(x[613]), .Q(
        xin[613]) );
  DFF \xreg_reg[614]  ( .D(xin[613]), .CLK(clk), .RST(start), .I(x[614]), .Q(
        xin[614]) );
  DFF \xreg_reg[615]  ( .D(xin[614]), .CLK(clk), .RST(start), .I(x[615]), .Q(
        xin[615]) );
  DFF \xreg_reg[616]  ( .D(xin[615]), .CLK(clk), .RST(start), .I(x[616]), .Q(
        xin[616]) );
  DFF \xreg_reg[617]  ( .D(xin[616]), .CLK(clk), .RST(start), .I(x[617]), .Q(
        xin[617]) );
  DFF \xreg_reg[618]  ( .D(xin[617]), .CLK(clk), .RST(start), .I(x[618]), .Q(
        xin[618]) );
  DFF \xreg_reg[619]  ( .D(xin[618]), .CLK(clk), .RST(start), .I(x[619]), .Q(
        xin[619]) );
  DFF \xreg_reg[620]  ( .D(xin[619]), .CLK(clk), .RST(start), .I(x[620]), .Q(
        xin[620]) );
  DFF \xreg_reg[621]  ( .D(xin[620]), .CLK(clk), .RST(start), .I(x[621]), .Q(
        xin[621]) );
  DFF \xreg_reg[622]  ( .D(xin[621]), .CLK(clk), .RST(start), .I(x[622]), .Q(
        xin[622]) );
  DFF \xreg_reg[623]  ( .D(xin[622]), .CLK(clk), .RST(start), .I(x[623]), .Q(
        xin[623]) );
  DFF \xreg_reg[624]  ( .D(xin[623]), .CLK(clk), .RST(start), .I(x[624]), .Q(
        xin[624]) );
  DFF \xreg_reg[625]  ( .D(xin[624]), .CLK(clk), .RST(start), .I(x[625]), .Q(
        xin[625]) );
  DFF \xreg_reg[626]  ( .D(xin[625]), .CLK(clk), .RST(start), .I(x[626]), .Q(
        xin[626]) );
  DFF \xreg_reg[627]  ( .D(xin[626]), .CLK(clk), .RST(start), .I(x[627]), .Q(
        xin[627]) );
  DFF \xreg_reg[628]  ( .D(xin[627]), .CLK(clk), .RST(start), .I(x[628]), .Q(
        xin[628]) );
  DFF \xreg_reg[629]  ( .D(xin[628]), .CLK(clk), .RST(start), .I(x[629]), .Q(
        xin[629]) );
  DFF \xreg_reg[630]  ( .D(xin[629]), .CLK(clk), .RST(start), .I(x[630]), .Q(
        xin[630]) );
  DFF \xreg_reg[631]  ( .D(xin[630]), .CLK(clk), .RST(start), .I(x[631]), .Q(
        xin[631]) );
  DFF \xreg_reg[632]  ( .D(xin[631]), .CLK(clk), .RST(start), .I(x[632]), .Q(
        xin[632]) );
  DFF \xreg_reg[633]  ( .D(xin[632]), .CLK(clk), .RST(start), .I(x[633]), .Q(
        xin[633]) );
  DFF \xreg_reg[634]  ( .D(xin[633]), .CLK(clk), .RST(start), .I(x[634]), .Q(
        xin[634]) );
  DFF \xreg_reg[635]  ( .D(xin[634]), .CLK(clk), .RST(start), .I(x[635]), .Q(
        xin[635]) );
  DFF \xreg_reg[636]  ( .D(xin[635]), .CLK(clk), .RST(start), .I(x[636]), .Q(
        xin[636]) );
  DFF \xreg_reg[637]  ( .D(xin[636]), .CLK(clk), .RST(start), .I(x[637]), .Q(
        xin[637]) );
  DFF \xreg_reg[638]  ( .D(xin[637]), .CLK(clk), .RST(start), .I(x[638]), .Q(
        xin[638]) );
  DFF \xreg_reg[639]  ( .D(xin[638]), .CLK(clk), .RST(start), .I(x[639]), .Q(
        xin[639]) );
  DFF \xreg_reg[640]  ( .D(xin[639]), .CLK(clk), .RST(start), .I(x[640]), .Q(
        xin[640]) );
  DFF \xreg_reg[641]  ( .D(xin[640]), .CLK(clk), .RST(start), .I(x[641]), .Q(
        xin[641]) );
  DFF \xreg_reg[642]  ( .D(xin[641]), .CLK(clk), .RST(start), .I(x[642]), .Q(
        xin[642]) );
  DFF \xreg_reg[643]  ( .D(xin[642]), .CLK(clk), .RST(start), .I(x[643]), .Q(
        xin[643]) );
  DFF \xreg_reg[644]  ( .D(xin[643]), .CLK(clk), .RST(start), .I(x[644]), .Q(
        xin[644]) );
  DFF \xreg_reg[645]  ( .D(xin[644]), .CLK(clk), .RST(start), .I(x[645]), .Q(
        xin[645]) );
  DFF \xreg_reg[646]  ( .D(xin[645]), .CLK(clk), .RST(start), .I(x[646]), .Q(
        xin[646]) );
  DFF \xreg_reg[647]  ( .D(xin[646]), .CLK(clk), .RST(start), .I(x[647]), .Q(
        xin[647]) );
  DFF \xreg_reg[648]  ( .D(xin[647]), .CLK(clk), .RST(start), .I(x[648]), .Q(
        xin[648]) );
  DFF \xreg_reg[649]  ( .D(xin[648]), .CLK(clk), .RST(start), .I(x[649]), .Q(
        xin[649]) );
  DFF \xreg_reg[650]  ( .D(xin[649]), .CLK(clk), .RST(start), .I(x[650]), .Q(
        xin[650]) );
  DFF \xreg_reg[651]  ( .D(xin[650]), .CLK(clk), .RST(start), .I(x[651]), .Q(
        xin[651]) );
  DFF \xreg_reg[652]  ( .D(xin[651]), .CLK(clk), .RST(start), .I(x[652]), .Q(
        xin[652]) );
  DFF \xreg_reg[653]  ( .D(xin[652]), .CLK(clk), .RST(start), .I(x[653]), .Q(
        xin[653]) );
  DFF \xreg_reg[654]  ( .D(xin[653]), .CLK(clk), .RST(start), .I(x[654]), .Q(
        xin[654]) );
  DFF \xreg_reg[655]  ( .D(xin[654]), .CLK(clk), .RST(start), .I(x[655]), .Q(
        xin[655]) );
  DFF \xreg_reg[656]  ( .D(xin[655]), .CLK(clk), .RST(start), .I(x[656]), .Q(
        xin[656]) );
  DFF \xreg_reg[657]  ( .D(xin[656]), .CLK(clk), .RST(start), .I(x[657]), .Q(
        xin[657]) );
  DFF \xreg_reg[658]  ( .D(xin[657]), .CLK(clk), .RST(start), .I(x[658]), .Q(
        xin[658]) );
  DFF \xreg_reg[659]  ( .D(xin[658]), .CLK(clk), .RST(start), .I(x[659]), .Q(
        xin[659]) );
  DFF \xreg_reg[660]  ( .D(xin[659]), .CLK(clk), .RST(start), .I(x[660]), .Q(
        xin[660]) );
  DFF \xreg_reg[661]  ( .D(xin[660]), .CLK(clk), .RST(start), .I(x[661]), .Q(
        xin[661]) );
  DFF \xreg_reg[662]  ( .D(xin[661]), .CLK(clk), .RST(start), .I(x[662]), .Q(
        xin[662]) );
  DFF \xreg_reg[663]  ( .D(xin[662]), .CLK(clk), .RST(start), .I(x[663]), .Q(
        xin[663]) );
  DFF \xreg_reg[664]  ( .D(xin[663]), .CLK(clk), .RST(start), .I(x[664]), .Q(
        xin[664]) );
  DFF \xreg_reg[665]  ( .D(xin[664]), .CLK(clk), .RST(start), .I(x[665]), .Q(
        xin[665]) );
  DFF \xreg_reg[666]  ( .D(xin[665]), .CLK(clk), .RST(start), .I(x[666]), .Q(
        xin[666]) );
  DFF \xreg_reg[667]  ( .D(xin[666]), .CLK(clk), .RST(start), .I(x[667]), .Q(
        xin[667]) );
  DFF \xreg_reg[668]  ( .D(xin[667]), .CLK(clk), .RST(start), .I(x[668]), .Q(
        xin[668]) );
  DFF \xreg_reg[669]  ( .D(xin[668]), .CLK(clk), .RST(start), .I(x[669]), .Q(
        xin[669]) );
  DFF \xreg_reg[670]  ( .D(xin[669]), .CLK(clk), .RST(start), .I(x[670]), .Q(
        xin[670]) );
  DFF \xreg_reg[671]  ( .D(xin[670]), .CLK(clk), .RST(start), .I(x[671]), .Q(
        xin[671]) );
  DFF \xreg_reg[672]  ( .D(xin[671]), .CLK(clk), .RST(start), .I(x[672]), .Q(
        xin[672]) );
  DFF \xreg_reg[673]  ( .D(xin[672]), .CLK(clk), .RST(start), .I(x[673]), .Q(
        xin[673]) );
  DFF \xreg_reg[674]  ( .D(xin[673]), .CLK(clk), .RST(start), .I(x[674]), .Q(
        xin[674]) );
  DFF \xreg_reg[675]  ( .D(xin[674]), .CLK(clk), .RST(start), .I(x[675]), .Q(
        xin[675]) );
  DFF \xreg_reg[676]  ( .D(xin[675]), .CLK(clk), .RST(start), .I(x[676]), .Q(
        xin[676]) );
  DFF \xreg_reg[677]  ( .D(xin[676]), .CLK(clk), .RST(start), .I(x[677]), .Q(
        xin[677]) );
  DFF \xreg_reg[678]  ( .D(xin[677]), .CLK(clk), .RST(start), .I(x[678]), .Q(
        xin[678]) );
  DFF \xreg_reg[679]  ( .D(xin[678]), .CLK(clk), .RST(start), .I(x[679]), .Q(
        xin[679]) );
  DFF \xreg_reg[680]  ( .D(xin[679]), .CLK(clk), .RST(start), .I(x[680]), .Q(
        xin[680]) );
  DFF \xreg_reg[681]  ( .D(xin[680]), .CLK(clk), .RST(start), .I(x[681]), .Q(
        xin[681]) );
  DFF \xreg_reg[682]  ( .D(xin[681]), .CLK(clk), .RST(start), .I(x[682]), .Q(
        xin[682]) );
  DFF \xreg_reg[683]  ( .D(xin[682]), .CLK(clk), .RST(start), .I(x[683]), .Q(
        xin[683]) );
  DFF \xreg_reg[684]  ( .D(xin[683]), .CLK(clk), .RST(start), .I(x[684]), .Q(
        xin[684]) );
  DFF \xreg_reg[685]  ( .D(xin[684]), .CLK(clk), .RST(start), .I(x[685]), .Q(
        xin[685]) );
  DFF \xreg_reg[686]  ( .D(xin[685]), .CLK(clk), .RST(start), .I(x[686]), .Q(
        xin[686]) );
  DFF \xreg_reg[687]  ( .D(xin[686]), .CLK(clk), .RST(start), .I(x[687]), .Q(
        xin[687]) );
  DFF \xreg_reg[688]  ( .D(xin[687]), .CLK(clk), .RST(start), .I(x[688]), .Q(
        xin[688]) );
  DFF \xreg_reg[689]  ( .D(xin[688]), .CLK(clk), .RST(start), .I(x[689]), .Q(
        xin[689]) );
  DFF \xreg_reg[690]  ( .D(xin[689]), .CLK(clk), .RST(start), .I(x[690]), .Q(
        xin[690]) );
  DFF \xreg_reg[691]  ( .D(xin[690]), .CLK(clk), .RST(start), .I(x[691]), .Q(
        xin[691]) );
  DFF \xreg_reg[692]  ( .D(xin[691]), .CLK(clk), .RST(start), .I(x[692]), .Q(
        xin[692]) );
  DFF \xreg_reg[693]  ( .D(xin[692]), .CLK(clk), .RST(start), .I(x[693]), .Q(
        xin[693]) );
  DFF \xreg_reg[694]  ( .D(xin[693]), .CLK(clk), .RST(start), .I(x[694]), .Q(
        xin[694]) );
  DFF \xreg_reg[695]  ( .D(xin[694]), .CLK(clk), .RST(start), .I(x[695]), .Q(
        xin[695]) );
  DFF \xreg_reg[696]  ( .D(xin[695]), .CLK(clk), .RST(start), .I(x[696]), .Q(
        xin[696]) );
  DFF \xreg_reg[697]  ( .D(xin[696]), .CLK(clk), .RST(start), .I(x[697]), .Q(
        xin[697]) );
  DFF \xreg_reg[698]  ( .D(xin[697]), .CLK(clk), .RST(start), .I(x[698]), .Q(
        xin[698]) );
  DFF \xreg_reg[699]  ( .D(xin[698]), .CLK(clk), .RST(start), .I(x[699]), .Q(
        xin[699]) );
  DFF \xreg_reg[700]  ( .D(xin[699]), .CLK(clk), .RST(start), .I(x[700]), .Q(
        xin[700]) );
  DFF \xreg_reg[701]  ( .D(xin[700]), .CLK(clk), .RST(start), .I(x[701]), .Q(
        xin[701]) );
  DFF \xreg_reg[702]  ( .D(xin[701]), .CLK(clk), .RST(start), .I(x[702]), .Q(
        xin[702]) );
  DFF \xreg_reg[703]  ( .D(xin[702]), .CLK(clk), .RST(start), .I(x[703]), .Q(
        xin[703]) );
  DFF \xreg_reg[704]  ( .D(xin[703]), .CLK(clk), .RST(start), .I(x[704]), .Q(
        xin[704]) );
  DFF \xreg_reg[705]  ( .D(xin[704]), .CLK(clk), .RST(start), .I(x[705]), .Q(
        xin[705]) );
  DFF \xreg_reg[706]  ( .D(xin[705]), .CLK(clk), .RST(start), .I(x[706]), .Q(
        xin[706]) );
  DFF \xreg_reg[707]  ( .D(xin[706]), .CLK(clk), .RST(start), .I(x[707]), .Q(
        xin[707]) );
  DFF \xreg_reg[708]  ( .D(xin[707]), .CLK(clk), .RST(start), .I(x[708]), .Q(
        xin[708]) );
  DFF \xreg_reg[709]  ( .D(xin[708]), .CLK(clk), .RST(start), .I(x[709]), .Q(
        xin[709]) );
  DFF \xreg_reg[710]  ( .D(xin[709]), .CLK(clk), .RST(start), .I(x[710]), .Q(
        xin[710]) );
  DFF \xreg_reg[711]  ( .D(xin[710]), .CLK(clk), .RST(start), .I(x[711]), .Q(
        xin[711]) );
  DFF \xreg_reg[712]  ( .D(xin[711]), .CLK(clk), .RST(start), .I(x[712]), .Q(
        xin[712]) );
  DFF \xreg_reg[713]  ( .D(xin[712]), .CLK(clk), .RST(start), .I(x[713]), .Q(
        xin[713]) );
  DFF \xreg_reg[714]  ( .D(xin[713]), .CLK(clk), .RST(start), .I(x[714]), .Q(
        xin[714]) );
  DFF \xreg_reg[715]  ( .D(xin[714]), .CLK(clk), .RST(start), .I(x[715]), .Q(
        xin[715]) );
  DFF \xreg_reg[716]  ( .D(xin[715]), .CLK(clk), .RST(start), .I(x[716]), .Q(
        xin[716]) );
  DFF \xreg_reg[717]  ( .D(xin[716]), .CLK(clk), .RST(start), .I(x[717]), .Q(
        xin[717]) );
  DFF \xreg_reg[718]  ( .D(xin[717]), .CLK(clk), .RST(start), .I(x[718]), .Q(
        xin[718]) );
  DFF \xreg_reg[719]  ( .D(xin[718]), .CLK(clk), .RST(start), .I(x[719]), .Q(
        xin[719]) );
  DFF \xreg_reg[720]  ( .D(xin[719]), .CLK(clk), .RST(start), .I(x[720]), .Q(
        xin[720]) );
  DFF \xreg_reg[721]  ( .D(xin[720]), .CLK(clk), .RST(start), .I(x[721]), .Q(
        xin[721]) );
  DFF \xreg_reg[722]  ( .D(xin[721]), .CLK(clk), .RST(start), .I(x[722]), .Q(
        xin[722]) );
  DFF \xreg_reg[723]  ( .D(xin[722]), .CLK(clk), .RST(start), .I(x[723]), .Q(
        xin[723]) );
  DFF \xreg_reg[724]  ( .D(xin[723]), .CLK(clk), .RST(start), .I(x[724]), .Q(
        xin[724]) );
  DFF \xreg_reg[725]  ( .D(xin[724]), .CLK(clk), .RST(start), .I(x[725]), .Q(
        xin[725]) );
  DFF \xreg_reg[726]  ( .D(xin[725]), .CLK(clk), .RST(start), .I(x[726]), .Q(
        xin[726]) );
  DFF \xreg_reg[727]  ( .D(xin[726]), .CLK(clk), .RST(start), .I(x[727]), .Q(
        xin[727]) );
  DFF \xreg_reg[728]  ( .D(xin[727]), .CLK(clk), .RST(start), .I(x[728]), .Q(
        xin[728]) );
  DFF \xreg_reg[729]  ( .D(xin[728]), .CLK(clk), .RST(start), .I(x[729]), .Q(
        xin[729]) );
  DFF \xreg_reg[730]  ( .D(xin[729]), .CLK(clk), .RST(start), .I(x[730]), .Q(
        xin[730]) );
  DFF \xreg_reg[731]  ( .D(xin[730]), .CLK(clk), .RST(start), .I(x[731]), .Q(
        xin[731]) );
  DFF \xreg_reg[732]  ( .D(xin[731]), .CLK(clk), .RST(start), .I(x[732]), .Q(
        xin[732]) );
  DFF \xreg_reg[733]  ( .D(xin[732]), .CLK(clk), .RST(start), .I(x[733]), .Q(
        xin[733]) );
  DFF \xreg_reg[734]  ( .D(xin[733]), .CLK(clk), .RST(start), .I(x[734]), .Q(
        xin[734]) );
  DFF \xreg_reg[735]  ( .D(xin[734]), .CLK(clk), .RST(start), .I(x[735]), .Q(
        xin[735]) );
  DFF \xreg_reg[736]  ( .D(xin[735]), .CLK(clk), .RST(start), .I(x[736]), .Q(
        xin[736]) );
  DFF \xreg_reg[737]  ( .D(xin[736]), .CLK(clk), .RST(start), .I(x[737]), .Q(
        xin[737]) );
  DFF \xreg_reg[738]  ( .D(xin[737]), .CLK(clk), .RST(start), .I(x[738]), .Q(
        xin[738]) );
  DFF \xreg_reg[739]  ( .D(xin[738]), .CLK(clk), .RST(start), .I(x[739]), .Q(
        xin[739]) );
  DFF \xreg_reg[740]  ( .D(xin[739]), .CLK(clk), .RST(start), .I(x[740]), .Q(
        xin[740]) );
  DFF \xreg_reg[741]  ( .D(xin[740]), .CLK(clk), .RST(start), .I(x[741]), .Q(
        xin[741]) );
  DFF \xreg_reg[742]  ( .D(xin[741]), .CLK(clk), .RST(start), .I(x[742]), .Q(
        xin[742]) );
  DFF \xreg_reg[743]  ( .D(xin[742]), .CLK(clk), .RST(start), .I(x[743]), .Q(
        xin[743]) );
  DFF \xreg_reg[744]  ( .D(xin[743]), .CLK(clk), .RST(start), .I(x[744]), .Q(
        xin[744]) );
  DFF \xreg_reg[745]  ( .D(xin[744]), .CLK(clk), .RST(start), .I(x[745]), .Q(
        xin[745]) );
  DFF \xreg_reg[746]  ( .D(xin[745]), .CLK(clk), .RST(start), .I(x[746]), .Q(
        xin[746]) );
  DFF \xreg_reg[747]  ( .D(xin[746]), .CLK(clk), .RST(start), .I(x[747]), .Q(
        xin[747]) );
  DFF \xreg_reg[748]  ( .D(xin[747]), .CLK(clk), .RST(start), .I(x[748]), .Q(
        xin[748]) );
  DFF \xreg_reg[749]  ( .D(xin[748]), .CLK(clk), .RST(start), .I(x[749]), .Q(
        xin[749]) );
  DFF \xreg_reg[750]  ( .D(xin[749]), .CLK(clk), .RST(start), .I(x[750]), .Q(
        xin[750]) );
  DFF \xreg_reg[751]  ( .D(xin[750]), .CLK(clk), .RST(start), .I(x[751]), .Q(
        xin[751]) );
  DFF \xreg_reg[752]  ( .D(xin[751]), .CLK(clk), .RST(start), .I(x[752]), .Q(
        xin[752]) );
  DFF \xreg_reg[753]  ( .D(xin[752]), .CLK(clk), .RST(start), .I(x[753]), .Q(
        xin[753]) );
  DFF \xreg_reg[754]  ( .D(xin[753]), .CLK(clk), .RST(start), .I(x[754]), .Q(
        xin[754]) );
  DFF \xreg_reg[755]  ( .D(xin[754]), .CLK(clk), .RST(start), .I(x[755]), .Q(
        xin[755]) );
  DFF \xreg_reg[756]  ( .D(xin[755]), .CLK(clk), .RST(start), .I(x[756]), .Q(
        xin[756]) );
  DFF \xreg_reg[757]  ( .D(xin[756]), .CLK(clk), .RST(start), .I(x[757]), .Q(
        xin[757]) );
  DFF \xreg_reg[758]  ( .D(xin[757]), .CLK(clk), .RST(start), .I(x[758]), .Q(
        xin[758]) );
  DFF \xreg_reg[759]  ( .D(xin[758]), .CLK(clk), .RST(start), .I(x[759]), .Q(
        xin[759]) );
  DFF \xreg_reg[760]  ( .D(xin[759]), .CLK(clk), .RST(start), .I(x[760]), .Q(
        xin[760]) );
  DFF \xreg_reg[761]  ( .D(xin[760]), .CLK(clk), .RST(start), .I(x[761]), .Q(
        xin[761]) );
  DFF \xreg_reg[762]  ( .D(xin[761]), .CLK(clk), .RST(start), .I(x[762]), .Q(
        xin[762]) );
  DFF \xreg_reg[763]  ( .D(xin[762]), .CLK(clk), .RST(start), .I(x[763]), .Q(
        xin[763]) );
  DFF \xreg_reg[764]  ( .D(xin[763]), .CLK(clk), .RST(start), .I(x[764]), .Q(
        xin[764]) );
  DFF \xreg_reg[765]  ( .D(xin[764]), .CLK(clk), .RST(start), .I(x[765]), .Q(
        xin[765]) );
  DFF \xreg_reg[766]  ( .D(xin[765]), .CLK(clk), .RST(start), .I(x[766]), .Q(
        xin[766]) );
  DFF \xreg_reg[767]  ( .D(xin[766]), .CLK(clk), .RST(start), .I(x[767]), .Q(
        xin[767]) );
  DFF \xreg_reg[768]  ( .D(xin[767]), .CLK(clk), .RST(start), .I(x[768]), .Q(
        xin[768]) );
  DFF \xreg_reg[769]  ( .D(xin[768]), .CLK(clk), .RST(start), .I(x[769]), .Q(
        xin[769]) );
  DFF \xreg_reg[770]  ( .D(xin[769]), .CLK(clk), .RST(start), .I(x[770]), .Q(
        xin[770]) );
  DFF \xreg_reg[771]  ( .D(xin[770]), .CLK(clk), .RST(start), .I(x[771]), .Q(
        xin[771]) );
  DFF \xreg_reg[772]  ( .D(xin[771]), .CLK(clk), .RST(start), .I(x[772]), .Q(
        xin[772]) );
  DFF \xreg_reg[773]  ( .D(xin[772]), .CLK(clk), .RST(start), .I(x[773]), .Q(
        xin[773]) );
  DFF \xreg_reg[774]  ( .D(xin[773]), .CLK(clk), .RST(start), .I(x[774]), .Q(
        xin[774]) );
  DFF \xreg_reg[775]  ( .D(xin[774]), .CLK(clk), .RST(start), .I(x[775]), .Q(
        xin[775]) );
  DFF \xreg_reg[776]  ( .D(xin[775]), .CLK(clk), .RST(start), .I(x[776]), .Q(
        xin[776]) );
  DFF \xreg_reg[777]  ( .D(xin[776]), .CLK(clk), .RST(start), .I(x[777]), .Q(
        xin[777]) );
  DFF \xreg_reg[778]  ( .D(xin[777]), .CLK(clk), .RST(start), .I(x[778]), .Q(
        xin[778]) );
  DFF \xreg_reg[779]  ( .D(xin[778]), .CLK(clk), .RST(start), .I(x[779]), .Q(
        xin[779]) );
  DFF \xreg_reg[780]  ( .D(xin[779]), .CLK(clk), .RST(start), .I(x[780]), .Q(
        xin[780]) );
  DFF \xreg_reg[781]  ( .D(xin[780]), .CLK(clk), .RST(start), .I(x[781]), .Q(
        xin[781]) );
  DFF \xreg_reg[782]  ( .D(xin[781]), .CLK(clk), .RST(start), .I(x[782]), .Q(
        xin[782]) );
  DFF \xreg_reg[783]  ( .D(xin[782]), .CLK(clk), .RST(start), .I(x[783]), .Q(
        xin[783]) );
  DFF \xreg_reg[784]  ( .D(xin[783]), .CLK(clk), .RST(start), .I(x[784]), .Q(
        xin[784]) );
  DFF \xreg_reg[785]  ( .D(xin[784]), .CLK(clk), .RST(start), .I(x[785]), .Q(
        xin[785]) );
  DFF \xreg_reg[786]  ( .D(xin[785]), .CLK(clk), .RST(start), .I(x[786]), .Q(
        xin[786]) );
  DFF \xreg_reg[787]  ( .D(xin[786]), .CLK(clk), .RST(start), .I(x[787]), .Q(
        xin[787]) );
  DFF \xreg_reg[788]  ( .D(xin[787]), .CLK(clk), .RST(start), .I(x[788]), .Q(
        xin[788]) );
  DFF \xreg_reg[789]  ( .D(xin[788]), .CLK(clk), .RST(start), .I(x[789]), .Q(
        xin[789]) );
  DFF \xreg_reg[790]  ( .D(xin[789]), .CLK(clk), .RST(start), .I(x[790]), .Q(
        xin[790]) );
  DFF \xreg_reg[791]  ( .D(xin[790]), .CLK(clk), .RST(start), .I(x[791]), .Q(
        xin[791]) );
  DFF \xreg_reg[792]  ( .D(xin[791]), .CLK(clk), .RST(start), .I(x[792]), .Q(
        xin[792]) );
  DFF \xreg_reg[793]  ( .D(xin[792]), .CLK(clk), .RST(start), .I(x[793]), .Q(
        xin[793]) );
  DFF \xreg_reg[794]  ( .D(xin[793]), .CLK(clk), .RST(start), .I(x[794]), .Q(
        xin[794]) );
  DFF \xreg_reg[795]  ( .D(xin[794]), .CLK(clk), .RST(start), .I(x[795]), .Q(
        xin[795]) );
  DFF \xreg_reg[796]  ( .D(xin[795]), .CLK(clk), .RST(start), .I(x[796]), .Q(
        xin[796]) );
  DFF \xreg_reg[797]  ( .D(xin[796]), .CLK(clk), .RST(start), .I(x[797]), .Q(
        xin[797]) );
  DFF \xreg_reg[798]  ( .D(xin[797]), .CLK(clk), .RST(start), .I(x[798]), .Q(
        xin[798]) );
  DFF \xreg_reg[799]  ( .D(xin[798]), .CLK(clk), .RST(start), .I(x[799]), .Q(
        xin[799]) );
  DFF \xreg_reg[800]  ( .D(xin[799]), .CLK(clk), .RST(start), .I(x[800]), .Q(
        xin[800]) );
  DFF \xreg_reg[801]  ( .D(xin[800]), .CLK(clk), .RST(start), .I(x[801]), .Q(
        xin[801]) );
  DFF \xreg_reg[802]  ( .D(xin[801]), .CLK(clk), .RST(start), .I(x[802]), .Q(
        xin[802]) );
  DFF \xreg_reg[803]  ( .D(xin[802]), .CLK(clk), .RST(start), .I(x[803]), .Q(
        xin[803]) );
  DFF \xreg_reg[804]  ( .D(xin[803]), .CLK(clk), .RST(start), .I(x[804]), .Q(
        xin[804]) );
  DFF \xreg_reg[805]  ( .D(xin[804]), .CLK(clk), .RST(start), .I(x[805]), .Q(
        xin[805]) );
  DFF \xreg_reg[806]  ( .D(xin[805]), .CLK(clk), .RST(start), .I(x[806]), .Q(
        xin[806]) );
  DFF \xreg_reg[807]  ( .D(xin[806]), .CLK(clk), .RST(start), .I(x[807]), .Q(
        xin[807]) );
  DFF \xreg_reg[808]  ( .D(xin[807]), .CLK(clk), .RST(start), .I(x[808]), .Q(
        xin[808]) );
  DFF \xreg_reg[809]  ( .D(xin[808]), .CLK(clk), .RST(start), .I(x[809]), .Q(
        xin[809]) );
  DFF \xreg_reg[810]  ( .D(xin[809]), .CLK(clk), .RST(start), .I(x[810]), .Q(
        xin[810]) );
  DFF \xreg_reg[811]  ( .D(xin[810]), .CLK(clk), .RST(start), .I(x[811]), .Q(
        xin[811]) );
  DFF \xreg_reg[812]  ( .D(xin[811]), .CLK(clk), .RST(start), .I(x[812]), .Q(
        xin[812]) );
  DFF \xreg_reg[813]  ( .D(xin[812]), .CLK(clk), .RST(start), .I(x[813]), .Q(
        xin[813]) );
  DFF \xreg_reg[814]  ( .D(xin[813]), .CLK(clk), .RST(start), .I(x[814]), .Q(
        xin[814]) );
  DFF \xreg_reg[815]  ( .D(xin[814]), .CLK(clk), .RST(start), .I(x[815]), .Q(
        xin[815]) );
  DFF \xreg_reg[816]  ( .D(xin[815]), .CLK(clk), .RST(start), .I(x[816]), .Q(
        xin[816]) );
  DFF \xreg_reg[817]  ( .D(xin[816]), .CLK(clk), .RST(start), .I(x[817]), .Q(
        xin[817]) );
  DFF \xreg_reg[818]  ( .D(xin[817]), .CLK(clk), .RST(start), .I(x[818]), .Q(
        xin[818]) );
  DFF \xreg_reg[819]  ( .D(xin[818]), .CLK(clk), .RST(start), .I(x[819]), .Q(
        xin[819]) );
  DFF \xreg_reg[820]  ( .D(xin[819]), .CLK(clk), .RST(start), .I(x[820]), .Q(
        xin[820]) );
  DFF \xreg_reg[821]  ( .D(xin[820]), .CLK(clk), .RST(start), .I(x[821]), .Q(
        xin[821]) );
  DFF \xreg_reg[822]  ( .D(xin[821]), .CLK(clk), .RST(start), .I(x[822]), .Q(
        xin[822]) );
  DFF \xreg_reg[823]  ( .D(xin[822]), .CLK(clk), .RST(start), .I(x[823]), .Q(
        xin[823]) );
  DFF \xreg_reg[824]  ( .D(xin[823]), .CLK(clk), .RST(start), .I(x[824]), .Q(
        xin[824]) );
  DFF \xreg_reg[825]  ( .D(xin[824]), .CLK(clk), .RST(start), .I(x[825]), .Q(
        xin[825]) );
  DFF \xreg_reg[826]  ( .D(xin[825]), .CLK(clk), .RST(start), .I(x[826]), .Q(
        xin[826]) );
  DFF \xreg_reg[827]  ( .D(xin[826]), .CLK(clk), .RST(start), .I(x[827]), .Q(
        xin[827]) );
  DFF \xreg_reg[828]  ( .D(xin[827]), .CLK(clk), .RST(start), .I(x[828]), .Q(
        xin[828]) );
  DFF \xreg_reg[829]  ( .D(xin[828]), .CLK(clk), .RST(start), .I(x[829]), .Q(
        xin[829]) );
  DFF \xreg_reg[830]  ( .D(xin[829]), .CLK(clk), .RST(start), .I(x[830]), .Q(
        xin[830]) );
  DFF \xreg_reg[831]  ( .D(xin[830]), .CLK(clk), .RST(start), .I(x[831]), .Q(
        xin[831]) );
  DFF \xreg_reg[832]  ( .D(xin[831]), .CLK(clk), .RST(start), .I(x[832]), .Q(
        xin[832]) );
  DFF \xreg_reg[833]  ( .D(xin[832]), .CLK(clk), .RST(start), .I(x[833]), .Q(
        xin[833]) );
  DFF \xreg_reg[834]  ( .D(xin[833]), .CLK(clk), .RST(start), .I(x[834]), .Q(
        xin[834]) );
  DFF \xreg_reg[835]  ( .D(xin[834]), .CLK(clk), .RST(start), .I(x[835]), .Q(
        xin[835]) );
  DFF \xreg_reg[836]  ( .D(xin[835]), .CLK(clk), .RST(start), .I(x[836]), .Q(
        xin[836]) );
  DFF \xreg_reg[837]  ( .D(xin[836]), .CLK(clk), .RST(start), .I(x[837]), .Q(
        xin[837]) );
  DFF \xreg_reg[838]  ( .D(xin[837]), .CLK(clk), .RST(start), .I(x[838]), .Q(
        xin[838]) );
  DFF \xreg_reg[839]  ( .D(xin[838]), .CLK(clk), .RST(start), .I(x[839]), .Q(
        xin[839]) );
  DFF \xreg_reg[840]  ( .D(xin[839]), .CLK(clk), .RST(start), .I(x[840]), .Q(
        xin[840]) );
  DFF \xreg_reg[841]  ( .D(xin[840]), .CLK(clk), .RST(start), .I(x[841]), .Q(
        xin[841]) );
  DFF \xreg_reg[842]  ( .D(xin[841]), .CLK(clk), .RST(start), .I(x[842]), .Q(
        xin[842]) );
  DFF \xreg_reg[843]  ( .D(xin[842]), .CLK(clk), .RST(start), .I(x[843]), .Q(
        xin[843]) );
  DFF \xreg_reg[844]  ( .D(xin[843]), .CLK(clk), .RST(start), .I(x[844]), .Q(
        xin[844]) );
  DFF \xreg_reg[845]  ( .D(xin[844]), .CLK(clk), .RST(start), .I(x[845]), .Q(
        xin[845]) );
  DFF \xreg_reg[846]  ( .D(xin[845]), .CLK(clk), .RST(start), .I(x[846]), .Q(
        xin[846]) );
  DFF \xreg_reg[847]  ( .D(xin[846]), .CLK(clk), .RST(start), .I(x[847]), .Q(
        xin[847]) );
  DFF \xreg_reg[848]  ( .D(xin[847]), .CLK(clk), .RST(start), .I(x[848]), .Q(
        xin[848]) );
  DFF \xreg_reg[849]  ( .D(xin[848]), .CLK(clk), .RST(start), .I(x[849]), .Q(
        xin[849]) );
  DFF \xreg_reg[850]  ( .D(xin[849]), .CLK(clk), .RST(start), .I(x[850]), .Q(
        xin[850]) );
  DFF \xreg_reg[851]  ( .D(xin[850]), .CLK(clk), .RST(start), .I(x[851]), .Q(
        xin[851]) );
  DFF \xreg_reg[852]  ( .D(xin[851]), .CLK(clk), .RST(start), .I(x[852]), .Q(
        xin[852]) );
  DFF \xreg_reg[853]  ( .D(xin[852]), .CLK(clk), .RST(start), .I(x[853]), .Q(
        xin[853]) );
  DFF \xreg_reg[854]  ( .D(xin[853]), .CLK(clk), .RST(start), .I(x[854]), .Q(
        xin[854]) );
  DFF \xreg_reg[855]  ( .D(xin[854]), .CLK(clk), .RST(start), .I(x[855]), .Q(
        xin[855]) );
  DFF \xreg_reg[856]  ( .D(xin[855]), .CLK(clk), .RST(start), .I(x[856]), .Q(
        xin[856]) );
  DFF \xreg_reg[857]  ( .D(xin[856]), .CLK(clk), .RST(start), .I(x[857]), .Q(
        xin[857]) );
  DFF \xreg_reg[858]  ( .D(xin[857]), .CLK(clk), .RST(start), .I(x[858]), .Q(
        xin[858]) );
  DFF \xreg_reg[859]  ( .D(xin[858]), .CLK(clk), .RST(start), .I(x[859]), .Q(
        xin[859]) );
  DFF \xreg_reg[860]  ( .D(xin[859]), .CLK(clk), .RST(start), .I(x[860]), .Q(
        xin[860]) );
  DFF \xreg_reg[861]  ( .D(xin[860]), .CLK(clk), .RST(start), .I(x[861]), .Q(
        xin[861]) );
  DFF \xreg_reg[862]  ( .D(xin[861]), .CLK(clk), .RST(start), .I(x[862]), .Q(
        xin[862]) );
  DFF \xreg_reg[863]  ( .D(xin[862]), .CLK(clk), .RST(start), .I(x[863]), .Q(
        xin[863]) );
  DFF \xreg_reg[864]  ( .D(xin[863]), .CLK(clk), .RST(start), .I(x[864]), .Q(
        xin[864]) );
  DFF \xreg_reg[865]  ( .D(xin[864]), .CLK(clk), .RST(start), .I(x[865]), .Q(
        xin[865]) );
  DFF \xreg_reg[866]  ( .D(xin[865]), .CLK(clk), .RST(start), .I(x[866]), .Q(
        xin[866]) );
  DFF \xreg_reg[867]  ( .D(xin[866]), .CLK(clk), .RST(start), .I(x[867]), .Q(
        xin[867]) );
  DFF \xreg_reg[868]  ( .D(xin[867]), .CLK(clk), .RST(start), .I(x[868]), .Q(
        xin[868]) );
  DFF \xreg_reg[869]  ( .D(xin[868]), .CLK(clk), .RST(start), .I(x[869]), .Q(
        xin[869]) );
  DFF \xreg_reg[870]  ( .D(xin[869]), .CLK(clk), .RST(start), .I(x[870]), .Q(
        xin[870]) );
  DFF \xreg_reg[871]  ( .D(xin[870]), .CLK(clk), .RST(start), .I(x[871]), .Q(
        xin[871]) );
  DFF \xreg_reg[872]  ( .D(xin[871]), .CLK(clk), .RST(start), .I(x[872]), .Q(
        xin[872]) );
  DFF \xreg_reg[873]  ( .D(xin[872]), .CLK(clk), .RST(start), .I(x[873]), .Q(
        xin[873]) );
  DFF \xreg_reg[874]  ( .D(xin[873]), .CLK(clk), .RST(start), .I(x[874]), .Q(
        xin[874]) );
  DFF \xreg_reg[875]  ( .D(xin[874]), .CLK(clk), .RST(start), .I(x[875]), .Q(
        xin[875]) );
  DFF \xreg_reg[876]  ( .D(xin[875]), .CLK(clk), .RST(start), .I(x[876]), .Q(
        xin[876]) );
  DFF \xreg_reg[877]  ( .D(xin[876]), .CLK(clk), .RST(start), .I(x[877]), .Q(
        xin[877]) );
  DFF \xreg_reg[878]  ( .D(xin[877]), .CLK(clk), .RST(start), .I(x[878]), .Q(
        xin[878]) );
  DFF \xreg_reg[879]  ( .D(xin[878]), .CLK(clk), .RST(start), .I(x[879]), .Q(
        xin[879]) );
  DFF \xreg_reg[880]  ( .D(xin[879]), .CLK(clk), .RST(start), .I(x[880]), .Q(
        xin[880]) );
  DFF \xreg_reg[881]  ( .D(xin[880]), .CLK(clk), .RST(start), .I(x[881]), .Q(
        xin[881]) );
  DFF \xreg_reg[882]  ( .D(xin[881]), .CLK(clk), .RST(start), .I(x[882]), .Q(
        xin[882]) );
  DFF \xreg_reg[883]  ( .D(xin[882]), .CLK(clk), .RST(start), .I(x[883]), .Q(
        xin[883]) );
  DFF \xreg_reg[884]  ( .D(xin[883]), .CLK(clk), .RST(start), .I(x[884]), .Q(
        xin[884]) );
  DFF \xreg_reg[885]  ( .D(xin[884]), .CLK(clk), .RST(start), .I(x[885]), .Q(
        xin[885]) );
  DFF \xreg_reg[886]  ( .D(xin[885]), .CLK(clk), .RST(start), .I(x[886]), .Q(
        xin[886]) );
  DFF \xreg_reg[887]  ( .D(xin[886]), .CLK(clk), .RST(start), .I(x[887]), .Q(
        xin[887]) );
  DFF \xreg_reg[888]  ( .D(xin[887]), .CLK(clk), .RST(start), .I(x[888]), .Q(
        xin[888]) );
  DFF \xreg_reg[889]  ( .D(xin[888]), .CLK(clk), .RST(start), .I(x[889]), .Q(
        xin[889]) );
  DFF \xreg_reg[890]  ( .D(xin[889]), .CLK(clk), .RST(start), .I(x[890]), .Q(
        xin[890]) );
  DFF \xreg_reg[891]  ( .D(xin[890]), .CLK(clk), .RST(start), .I(x[891]), .Q(
        xin[891]) );
  DFF \xreg_reg[892]  ( .D(xin[891]), .CLK(clk), .RST(start), .I(x[892]), .Q(
        xin[892]) );
  DFF \xreg_reg[893]  ( .D(xin[892]), .CLK(clk), .RST(start), .I(x[893]), .Q(
        xin[893]) );
  DFF \xreg_reg[894]  ( .D(xin[893]), .CLK(clk), .RST(start), .I(x[894]), .Q(
        xin[894]) );
  DFF \xreg_reg[895]  ( .D(xin[894]), .CLK(clk), .RST(start), .I(x[895]), .Q(
        xin[895]) );
  DFF \xreg_reg[896]  ( .D(xin[895]), .CLK(clk), .RST(start), .I(x[896]), .Q(
        xin[896]) );
  DFF \xreg_reg[897]  ( .D(xin[896]), .CLK(clk), .RST(start), .I(x[897]), .Q(
        xin[897]) );
  DFF \xreg_reg[898]  ( .D(xin[897]), .CLK(clk), .RST(start), .I(x[898]), .Q(
        xin[898]) );
  DFF \xreg_reg[899]  ( .D(xin[898]), .CLK(clk), .RST(start), .I(x[899]), .Q(
        xin[899]) );
  DFF \xreg_reg[900]  ( .D(xin[899]), .CLK(clk), .RST(start), .I(x[900]), .Q(
        xin[900]) );
  DFF \xreg_reg[901]  ( .D(xin[900]), .CLK(clk), .RST(start), .I(x[901]), .Q(
        xin[901]) );
  DFF \xreg_reg[902]  ( .D(xin[901]), .CLK(clk), .RST(start), .I(x[902]), .Q(
        xin[902]) );
  DFF \xreg_reg[903]  ( .D(xin[902]), .CLK(clk), .RST(start), .I(x[903]), .Q(
        xin[903]) );
  DFF \xreg_reg[904]  ( .D(xin[903]), .CLK(clk), .RST(start), .I(x[904]), .Q(
        xin[904]) );
  DFF \xreg_reg[905]  ( .D(xin[904]), .CLK(clk), .RST(start), .I(x[905]), .Q(
        xin[905]) );
  DFF \xreg_reg[906]  ( .D(xin[905]), .CLK(clk), .RST(start), .I(x[906]), .Q(
        xin[906]) );
  DFF \xreg_reg[907]  ( .D(xin[906]), .CLK(clk), .RST(start), .I(x[907]), .Q(
        xin[907]) );
  DFF \xreg_reg[908]  ( .D(xin[907]), .CLK(clk), .RST(start), .I(x[908]), .Q(
        xin[908]) );
  DFF \xreg_reg[909]  ( .D(xin[908]), .CLK(clk), .RST(start), .I(x[909]), .Q(
        xin[909]) );
  DFF \xreg_reg[910]  ( .D(xin[909]), .CLK(clk), .RST(start), .I(x[910]), .Q(
        xin[910]) );
  DFF \xreg_reg[911]  ( .D(xin[910]), .CLK(clk), .RST(start), .I(x[911]), .Q(
        xin[911]) );
  DFF \xreg_reg[912]  ( .D(xin[911]), .CLK(clk), .RST(start), .I(x[912]), .Q(
        xin[912]) );
  DFF \xreg_reg[913]  ( .D(xin[912]), .CLK(clk), .RST(start), .I(x[913]), .Q(
        xin[913]) );
  DFF \xreg_reg[914]  ( .D(xin[913]), .CLK(clk), .RST(start), .I(x[914]), .Q(
        xin[914]) );
  DFF \xreg_reg[915]  ( .D(xin[914]), .CLK(clk), .RST(start), .I(x[915]), .Q(
        xin[915]) );
  DFF \xreg_reg[916]  ( .D(xin[915]), .CLK(clk), .RST(start), .I(x[916]), .Q(
        xin[916]) );
  DFF \xreg_reg[917]  ( .D(xin[916]), .CLK(clk), .RST(start), .I(x[917]), .Q(
        xin[917]) );
  DFF \xreg_reg[918]  ( .D(xin[917]), .CLK(clk), .RST(start), .I(x[918]), .Q(
        xin[918]) );
  DFF \xreg_reg[919]  ( .D(xin[918]), .CLK(clk), .RST(start), .I(x[919]), .Q(
        xin[919]) );
  DFF \xreg_reg[920]  ( .D(xin[919]), .CLK(clk), .RST(start), .I(x[920]), .Q(
        xin[920]) );
  DFF \xreg_reg[921]  ( .D(xin[920]), .CLK(clk), .RST(start), .I(x[921]), .Q(
        xin[921]) );
  DFF \xreg_reg[922]  ( .D(xin[921]), .CLK(clk), .RST(start), .I(x[922]), .Q(
        xin[922]) );
  DFF \xreg_reg[923]  ( .D(xin[922]), .CLK(clk), .RST(start), .I(x[923]), .Q(
        xin[923]) );
  DFF \xreg_reg[924]  ( .D(xin[923]), .CLK(clk), .RST(start), .I(x[924]), .Q(
        xin[924]) );
  DFF \xreg_reg[925]  ( .D(xin[924]), .CLK(clk), .RST(start), .I(x[925]), .Q(
        xin[925]) );
  DFF \xreg_reg[926]  ( .D(xin[925]), .CLK(clk), .RST(start), .I(x[926]), .Q(
        xin[926]) );
  DFF \xreg_reg[927]  ( .D(xin[926]), .CLK(clk), .RST(start), .I(x[927]), .Q(
        xin[927]) );
  DFF \xreg_reg[928]  ( .D(xin[927]), .CLK(clk), .RST(start), .I(x[928]), .Q(
        xin[928]) );
  DFF \xreg_reg[929]  ( .D(xin[928]), .CLK(clk), .RST(start), .I(x[929]), .Q(
        xin[929]) );
  DFF \xreg_reg[930]  ( .D(xin[929]), .CLK(clk), .RST(start), .I(x[930]), .Q(
        xin[930]) );
  DFF \xreg_reg[931]  ( .D(xin[930]), .CLK(clk), .RST(start), .I(x[931]), .Q(
        xin[931]) );
  DFF \xreg_reg[932]  ( .D(xin[931]), .CLK(clk), .RST(start), .I(x[932]), .Q(
        xin[932]) );
  DFF \xreg_reg[933]  ( .D(xin[932]), .CLK(clk), .RST(start), .I(x[933]), .Q(
        xin[933]) );
  DFF \xreg_reg[934]  ( .D(xin[933]), .CLK(clk), .RST(start), .I(x[934]), .Q(
        xin[934]) );
  DFF \xreg_reg[935]  ( .D(xin[934]), .CLK(clk), .RST(start), .I(x[935]), .Q(
        xin[935]) );
  DFF \xreg_reg[936]  ( .D(xin[935]), .CLK(clk), .RST(start), .I(x[936]), .Q(
        xin[936]) );
  DFF \xreg_reg[937]  ( .D(xin[936]), .CLK(clk), .RST(start), .I(x[937]), .Q(
        xin[937]) );
  DFF \xreg_reg[938]  ( .D(xin[937]), .CLK(clk), .RST(start), .I(x[938]), .Q(
        xin[938]) );
  DFF \xreg_reg[939]  ( .D(xin[938]), .CLK(clk), .RST(start), .I(x[939]), .Q(
        xin[939]) );
  DFF \xreg_reg[940]  ( .D(xin[939]), .CLK(clk), .RST(start), .I(x[940]), .Q(
        xin[940]) );
  DFF \xreg_reg[941]  ( .D(xin[940]), .CLK(clk), .RST(start), .I(x[941]), .Q(
        xin[941]) );
  DFF \xreg_reg[942]  ( .D(xin[941]), .CLK(clk), .RST(start), .I(x[942]), .Q(
        xin[942]) );
  DFF \xreg_reg[943]  ( .D(xin[942]), .CLK(clk), .RST(start), .I(x[943]), .Q(
        xin[943]) );
  DFF \xreg_reg[944]  ( .D(xin[943]), .CLK(clk), .RST(start), .I(x[944]), .Q(
        xin[944]) );
  DFF \xreg_reg[945]  ( .D(xin[944]), .CLK(clk), .RST(start), .I(x[945]), .Q(
        xin[945]) );
  DFF \xreg_reg[946]  ( .D(xin[945]), .CLK(clk), .RST(start), .I(x[946]), .Q(
        xin[946]) );
  DFF \xreg_reg[947]  ( .D(xin[946]), .CLK(clk), .RST(start), .I(x[947]), .Q(
        xin[947]) );
  DFF \xreg_reg[948]  ( .D(xin[947]), .CLK(clk), .RST(start), .I(x[948]), .Q(
        xin[948]) );
  DFF \xreg_reg[949]  ( .D(xin[948]), .CLK(clk), .RST(start), .I(x[949]), .Q(
        xin[949]) );
  DFF \xreg_reg[950]  ( .D(xin[949]), .CLK(clk), .RST(start), .I(x[950]), .Q(
        xin[950]) );
  DFF \xreg_reg[951]  ( .D(xin[950]), .CLK(clk), .RST(start), .I(x[951]), .Q(
        xin[951]) );
  DFF \xreg_reg[952]  ( .D(xin[951]), .CLK(clk), .RST(start), .I(x[952]), .Q(
        xin[952]) );
  DFF \xreg_reg[953]  ( .D(xin[952]), .CLK(clk), .RST(start), .I(x[953]), .Q(
        xin[953]) );
  DFF \xreg_reg[954]  ( .D(xin[953]), .CLK(clk), .RST(start), .I(x[954]), .Q(
        xin[954]) );
  DFF \xreg_reg[955]  ( .D(xin[954]), .CLK(clk), .RST(start), .I(x[955]), .Q(
        xin[955]) );
  DFF \xreg_reg[956]  ( .D(xin[955]), .CLK(clk), .RST(start), .I(x[956]), .Q(
        xin[956]) );
  DFF \xreg_reg[957]  ( .D(xin[956]), .CLK(clk), .RST(start), .I(x[957]), .Q(
        xin[957]) );
  DFF \xreg_reg[958]  ( .D(xin[957]), .CLK(clk), .RST(start), .I(x[958]), .Q(
        xin[958]) );
  DFF \xreg_reg[959]  ( .D(xin[958]), .CLK(clk), .RST(start), .I(x[959]), .Q(
        xin[959]) );
  DFF \xreg_reg[960]  ( .D(xin[959]), .CLK(clk), .RST(start), .I(x[960]), .Q(
        xin[960]) );
  DFF \xreg_reg[961]  ( .D(xin[960]), .CLK(clk), .RST(start), .I(x[961]), .Q(
        xin[961]) );
  DFF \xreg_reg[962]  ( .D(xin[961]), .CLK(clk), .RST(start), .I(x[962]), .Q(
        xin[962]) );
  DFF \xreg_reg[963]  ( .D(xin[962]), .CLK(clk), .RST(start), .I(x[963]), .Q(
        xin[963]) );
  DFF \xreg_reg[964]  ( .D(xin[963]), .CLK(clk), .RST(start), .I(x[964]), .Q(
        xin[964]) );
  DFF \xreg_reg[965]  ( .D(xin[964]), .CLK(clk), .RST(start), .I(x[965]), .Q(
        xin[965]) );
  DFF \xreg_reg[966]  ( .D(xin[965]), .CLK(clk), .RST(start), .I(x[966]), .Q(
        xin[966]) );
  DFF \xreg_reg[967]  ( .D(xin[966]), .CLK(clk), .RST(start), .I(x[967]), .Q(
        xin[967]) );
  DFF \xreg_reg[968]  ( .D(xin[967]), .CLK(clk), .RST(start), .I(x[968]), .Q(
        xin[968]) );
  DFF \xreg_reg[969]  ( .D(xin[968]), .CLK(clk), .RST(start), .I(x[969]), .Q(
        xin[969]) );
  DFF \xreg_reg[970]  ( .D(xin[969]), .CLK(clk), .RST(start), .I(x[970]), .Q(
        xin[970]) );
  DFF \xreg_reg[971]  ( .D(xin[970]), .CLK(clk), .RST(start), .I(x[971]), .Q(
        xin[971]) );
  DFF \xreg_reg[972]  ( .D(xin[971]), .CLK(clk), .RST(start), .I(x[972]), .Q(
        xin[972]) );
  DFF \xreg_reg[973]  ( .D(xin[972]), .CLK(clk), .RST(start), .I(x[973]), .Q(
        xin[973]) );
  DFF \xreg_reg[974]  ( .D(xin[973]), .CLK(clk), .RST(start), .I(x[974]), .Q(
        xin[974]) );
  DFF \xreg_reg[975]  ( .D(xin[974]), .CLK(clk), .RST(start), .I(x[975]), .Q(
        xin[975]) );
  DFF \xreg_reg[976]  ( .D(xin[975]), .CLK(clk), .RST(start), .I(x[976]), .Q(
        xin[976]) );
  DFF \xreg_reg[977]  ( .D(xin[976]), .CLK(clk), .RST(start), .I(x[977]), .Q(
        xin[977]) );
  DFF \xreg_reg[978]  ( .D(xin[977]), .CLK(clk), .RST(start), .I(x[978]), .Q(
        xin[978]) );
  DFF \xreg_reg[979]  ( .D(xin[978]), .CLK(clk), .RST(start), .I(x[979]), .Q(
        xin[979]) );
  DFF \xreg_reg[980]  ( .D(xin[979]), .CLK(clk), .RST(start), .I(x[980]), .Q(
        xin[980]) );
  DFF \xreg_reg[981]  ( .D(xin[980]), .CLK(clk), .RST(start), .I(x[981]), .Q(
        xin[981]) );
  DFF \xreg_reg[982]  ( .D(xin[981]), .CLK(clk), .RST(start), .I(x[982]), .Q(
        xin[982]) );
  DFF \xreg_reg[983]  ( .D(xin[982]), .CLK(clk), .RST(start), .I(x[983]), .Q(
        xin[983]) );
  DFF \xreg_reg[984]  ( .D(xin[983]), .CLK(clk), .RST(start), .I(x[984]), .Q(
        xin[984]) );
  DFF \xreg_reg[985]  ( .D(xin[984]), .CLK(clk), .RST(start), .I(x[985]), .Q(
        xin[985]) );
  DFF \xreg_reg[986]  ( .D(xin[985]), .CLK(clk), .RST(start), .I(x[986]), .Q(
        xin[986]) );
  DFF \xreg_reg[987]  ( .D(xin[986]), .CLK(clk), .RST(start), .I(x[987]), .Q(
        xin[987]) );
  DFF \xreg_reg[988]  ( .D(xin[987]), .CLK(clk), .RST(start), .I(x[988]), .Q(
        xin[988]) );
  DFF \xreg_reg[989]  ( .D(xin[988]), .CLK(clk), .RST(start), .I(x[989]), .Q(
        xin[989]) );
  DFF \xreg_reg[990]  ( .D(xin[989]), .CLK(clk), .RST(start), .I(x[990]), .Q(
        xin[990]) );
  DFF \xreg_reg[991]  ( .D(xin[990]), .CLK(clk), .RST(start), .I(x[991]), .Q(
        xin[991]) );
  DFF \xreg_reg[992]  ( .D(xin[991]), .CLK(clk), .RST(start), .I(x[992]), .Q(
        xin[992]) );
  DFF \xreg_reg[993]  ( .D(xin[992]), .CLK(clk), .RST(start), .I(x[993]), .Q(
        xin[993]) );
  DFF \xreg_reg[994]  ( .D(xin[993]), .CLK(clk), .RST(start), .I(x[994]), .Q(
        xin[994]) );
  DFF \xreg_reg[995]  ( .D(xin[994]), .CLK(clk), .RST(start), .I(x[995]), .Q(
        xin[995]) );
  DFF \xreg_reg[996]  ( .D(xin[995]), .CLK(clk), .RST(start), .I(x[996]), .Q(
        xin[996]) );
  DFF \xreg_reg[997]  ( .D(xin[996]), .CLK(clk), .RST(start), .I(x[997]), .Q(
        xin[997]) );
  DFF \xreg_reg[998]  ( .D(xin[997]), .CLK(clk), .RST(start), .I(x[998]), .Q(
        xin[998]) );
  DFF \xreg_reg[999]  ( .D(xin[998]), .CLK(clk), .RST(start), .I(x[999]), .Q(
        xin[999]) );
  DFF \xreg_reg[1000]  ( .D(xin[999]), .CLK(clk), .RST(start), .I(x[1000]), 
        .Q(xin[1000]) );
  DFF \xreg_reg[1001]  ( .D(xin[1000]), .CLK(clk), .RST(start), .I(x[1001]), 
        .Q(xin[1001]) );
  DFF \xreg_reg[1002]  ( .D(xin[1001]), .CLK(clk), .RST(start), .I(x[1002]), 
        .Q(xin[1002]) );
  DFF \xreg_reg[1003]  ( .D(xin[1002]), .CLK(clk), .RST(start), .I(x[1003]), 
        .Q(xin[1003]) );
  DFF \xreg_reg[1004]  ( .D(xin[1003]), .CLK(clk), .RST(start), .I(x[1004]), 
        .Q(xin[1004]) );
  DFF \xreg_reg[1005]  ( .D(xin[1004]), .CLK(clk), .RST(start), .I(x[1005]), 
        .Q(xin[1005]) );
  DFF \xreg_reg[1006]  ( .D(xin[1005]), .CLK(clk), .RST(start), .I(x[1006]), 
        .Q(xin[1006]) );
  DFF \xreg_reg[1007]  ( .D(xin[1006]), .CLK(clk), .RST(start), .I(x[1007]), 
        .Q(xin[1007]) );
  DFF \xreg_reg[1008]  ( .D(xin[1007]), .CLK(clk), .RST(start), .I(x[1008]), 
        .Q(xin[1008]) );
  DFF \xreg_reg[1009]  ( .D(xin[1008]), .CLK(clk), .RST(start), .I(x[1009]), 
        .Q(xin[1009]) );
  DFF \xreg_reg[1010]  ( .D(xin[1009]), .CLK(clk), .RST(start), .I(x[1010]), 
        .Q(xin[1010]) );
  DFF \xreg_reg[1011]  ( .D(xin[1010]), .CLK(clk), .RST(start), .I(x[1011]), 
        .Q(xin[1011]) );
  DFF \xreg_reg[1012]  ( .D(xin[1011]), .CLK(clk), .RST(start), .I(x[1012]), 
        .Q(xin[1012]) );
  DFF \xreg_reg[1013]  ( .D(xin[1012]), .CLK(clk), .RST(start), .I(x[1013]), 
        .Q(xin[1013]) );
  DFF \xreg_reg[1014]  ( .D(xin[1013]), .CLK(clk), .RST(start), .I(x[1014]), 
        .Q(xin[1014]) );
  DFF \xreg_reg[1015]  ( .D(xin[1014]), .CLK(clk), .RST(start), .I(x[1015]), 
        .Q(xin[1015]) );
  DFF \xreg_reg[1016]  ( .D(xin[1015]), .CLK(clk), .RST(start), .I(x[1016]), 
        .Q(xin[1016]) );
  DFF \xreg_reg[1017]  ( .D(xin[1016]), .CLK(clk), .RST(start), .I(x[1017]), 
        .Q(xin[1017]) );
  DFF \xreg_reg[1018]  ( .D(xin[1017]), .CLK(clk), .RST(start), .I(x[1018]), 
        .Q(xin[1018]) );
  DFF \xreg_reg[1019]  ( .D(xin[1018]), .CLK(clk), .RST(start), .I(x[1019]), 
        .Q(xin[1019]) );
  DFF \xreg_reg[1020]  ( .D(xin[1019]), .CLK(clk), .RST(start), .I(x[1020]), 
        .Q(xin[1020]) );
  DFF \xreg_reg[1021]  ( .D(xin[1020]), .CLK(clk), .RST(start), .I(x[1021]), 
        .Q(xin[1021]) );
  DFF \xreg_reg[1022]  ( .D(xin[1021]), .CLK(clk), .RST(start), .I(x[1022]), 
        .Q(xin[1022]) );
  DFF \xreg_reg[1023]  ( .D(xin[1022]), .CLK(clk), .RST(start), .I(x[1023]), 
        .Q(xin[1023]) );
  DFF \zreg_reg[0]  ( .D(o[0]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][0] ) );
  DFF \zreg_reg[1]  ( .D(o[1]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][1] ) );
  DFF \zreg_reg[2]  ( .D(o[2]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][2] ) );
  DFF \zreg_reg[3]  ( .D(o[3]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][3] ) );
  DFF \zreg_reg[4]  ( .D(o[4]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][4] ) );
  DFF \zreg_reg[5]  ( .D(o[5]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][5] ) );
  DFF \zreg_reg[6]  ( .D(o[6]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][6] ) );
  DFF \zreg_reg[7]  ( .D(o[7]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][7] ) );
  DFF \zreg_reg[8]  ( .D(o[8]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][8] ) );
  DFF \zreg_reg[9]  ( .D(o[9]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][9] ) );
  DFF \zreg_reg[10]  ( .D(o[10]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][10] ) );
  DFF \zreg_reg[11]  ( .D(o[11]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][11] ) );
  DFF \zreg_reg[12]  ( .D(o[12]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][12] ) );
  DFF \zreg_reg[13]  ( .D(o[13]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][13] ) );
  DFF \zreg_reg[14]  ( .D(o[14]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][14] ) );
  DFF \zreg_reg[15]  ( .D(o[15]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][15] ) );
  DFF \zreg_reg[16]  ( .D(o[16]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][16] ) );
  DFF \zreg_reg[17]  ( .D(o[17]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][17] ) );
  DFF \zreg_reg[18]  ( .D(o[18]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][18] ) );
  DFF \zreg_reg[19]  ( .D(o[19]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][19] ) );
  DFF \zreg_reg[20]  ( .D(o[20]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][20] ) );
  DFF \zreg_reg[21]  ( .D(o[21]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][21] ) );
  DFF \zreg_reg[22]  ( .D(o[22]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][22] ) );
  DFF \zreg_reg[23]  ( .D(o[23]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][23] ) );
  DFF \zreg_reg[24]  ( .D(o[24]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][24] ) );
  DFF \zreg_reg[25]  ( .D(o[25]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][25] ) );
  DFF \zreg_reg[26]  ( .D(o[26]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][26] ) );
  DFF \zreg_reg[27]  ( .D(o[27]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][27] ) );
  DFF \zreg_reg[28]  ( .D(o[28]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][28] ) );
  DFF \zreg_reg[29]  ( .D(o[29]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][29] ) );
  DFF \zreg_reg[30]  ( .D(o[30]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][30] ) );
  DFF \zreg_reg[31]  ( .D(o[31]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][31] ) );
  DFF \zreg_reg[32]  ( .D(o[32]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][32] ) );
  DFF \zreg_reg[33]  ( .D(o[33]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][33] ) );
  DFF \zreg_reg[34]  ( .D(o[34]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][34] ) );
  DFF \zreg_reg[35]  ( .D(o[35]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][35] ) );
  DFF \zreg_reg[36]  ( .D(o[36]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][36] ) );
  DFF \zreg_reg[37]  ( .D(o[37]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][37] ) );
  DFF \zreg_reg[38]  ( .D(o[38]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][38] ) );
  DFF \zreg_reg[39]  ( .D(o[39]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][39] ) );
  DFF \zreg_reg[40]  ( .D(o[40]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][40] ) );
  DFF \zreg_reg[41]  ( .D(o[41]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][41] ) );
  DFF \zreg_reg[42]  ( .D(o[42]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][42] ) );
  DFF \zreg_reg[43]  ( .D(o[43]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][43] ) );
  DFF \zreg_reg[44]  ( .D(o[44]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][44] ) );
  DFF \zreg_reg[45]  ( .D(o[45]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][45] ) );
  DFF \zreg_reg[46]  ( .D(o[46]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][46] ) );
  DFF \zreg_reg[47]  ( .D(o[47]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][47] ) );
  DFF \zreg_reg[48]  ( .D(o[48]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][48] ) );
  DFF \zreg_reg[49]  ( .D(o[49]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][49] ) );
  DFF \zreg_reg[50]  ( .D(o[50]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][50] ) );
  DFF \zreg_reg[51]  ( .D(o[51]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][51] ) );
  DFF \zreg_reg[52]  ( .D(o[52]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][52] ) );
  DFF \zreg_reg[53]  ( .D(o[53]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][53] ) );
  DFF \zreg_reg[54]  ( .D(o[54]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][54] ) );
  DFF \zreg_reg[55]  ( .D(o[55]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][55] ) );
  DFF \zreg_reg[56]  ( .D(o[56]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][56] ) );
  DFF \zreg_reg[57]  ( .D(o[57]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][57] ) );
  DFF \zreg_reg[58]  ( .D(o[58]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][58] ) );
  DFF \zreg_reg[59]  ( .D(o[59]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][59] ) );
  DFF \zreg_reg[60]  ( .D(o[60]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][60] ) );
  DFF \zreg_reg[61]  ( .D(o[61]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][61] ) );
  DFF \zreg_reg[62]  ( .D(o[62]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][62] ) );
  DFF \zreg_reg[63]  ( .D(o[63]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][63] ) );
  DFF \zreg_reg[64]  ( .D(o[64]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][64] ) );
  DFF \zreg_reg[65]  ( .D(o[65]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][65] ) );
  DFF \zreg_reg[66]  ( .D(o[66]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][66] ) );
  DFF \zreg_reg[67]  ( .D(o[67]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][67] ) );
  DFF \zreg_reg[68]  ( .D(o[68]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][68] ) );
  DFF \zreg_reg[69]  ( .D(o[69]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][69] ) );
  DFF \zreg_reg[70]  ( .D(o[70]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][70] ) );
  DFF \zreg_reg[71]  ( .D(o[71]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][71] ) );
  DFF \zreg_reg[72]  ( .D(o[72]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][72] ) );
  DFF \zreg_reg[73]  ( .D(o[73]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][73] ) );
  DFF \zreg_reg[74]  ( .D(o[74]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][74] ) );
  DFF \zreg_reg[75]  ( .D(o[75]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][75] ) );
  DFF \zreg_reg[76]  ( .D(o[76]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][76] ) );
  DFF \zreg_reg[77]  ( .D(o[77]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][77] ) );
  DFF \zreg_reg[78]  ( .D(o[78]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][78] ) );
  DFF \zreg_reg[79]  ( .D(o[79]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][79] ) );
  DFF \zreg_reg[80]  ( .D(o[80]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][80] ) );
  DFF \zreg_reg[81]  ( .D(o[81]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][81] ) );
  DFF \zreg_reg[82]  ( .D(o[82]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][82] ) );
  DFF \zreg_reg[83]  ( .D(o[83]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][83] ) );
  DFF \zreg_reg[84]  ( .D(o[84]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][84] ) );
  DFF \zreg_reg[85]  ( .D(o[85]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][85] ) );
  DFF \zreg_reg[86]  ( .D(o[86]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][86] ) );
  DFF \zreg_reg[87]  ( .D(o[87]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][87] ) );
  DFF \zreg_reg[88]  ( .D(o[88]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][88] ) );
  DFF \zreg_reg[89]  ( .D(o[89]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][89] ) );
  DFF \zreg_reg[90]  ( .D(o[90]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][90] ) );
  DFF \zreg_reg[91]  ( .D(o[91]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][91] ) );
  DFF \zreg_reg[92]  ( .D(o[92]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][92] ) );
  DFF \zreg_reg[93]  ( .D(o[93]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][93] ) );
  DFF \zreg_reg[94]  ( .D(o[94]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][94] ) );
  DFF \zreg_reg[95]  ( .D(o[95]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][95] ) );
  DFF \zreg_reg[96]  ( .D(o[96]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][96] ) );
  DFF \zreg_reg[97]  ( .D(o[97]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][97] ) );
  DFF \zreg_reg[98]  ( .D(o[98]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][98] ) );
  DFF \zreg_reg[99]  ( .D(o[99]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][99] ) );
  DFF \zreg_reg[100]  ( .D(o[100]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][100] ) );
  DFF \zreg_reg[101]  ( .D(o[101]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][101] ) );
  DFF \zreg_reg[102]  ( .D(o[102]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][102] ) );
  DFF \zreg_reg[103]  ( .D(o[103]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][103] ) );
  DFF \zreg_reg[104]  ( .D(o[104]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][104] ) );
  DFF \zreg_reg[105]  ( .D(o[105]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][105] ) );
  DFF \zreg_reg[106]  ( .D(o[106]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][106] ) );
  DFF \zreg_reg[107]  ( .D(o[107]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][107] ) );
  DFF \zreg_reg[108]  ( .D(o[108]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][108] ) );
  DFF \zreg_reg[109]  ( .D(o[109]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][109] ) );
  DFF \zreg_reg[110]  ( .D(o[110]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][110] ) );
  DFF \zreg_reg[111]  ( .D(o[111]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][111] ) );
  DFF \zreg_reg[112]  ( .D(o[112]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][112] ) );
  DFF \zreg_reg[113]  ( .D(o[113]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][113] ) );
  DFF \zreg_reg[114]  ( .D(o[114]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][114] ) );
  DFF \zreg_reg[115]  ( .D(o[115]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][115] ) );
  DFF \zreg_reg[116]  ( .D(o[116]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][116] ) );
  DFF \zreg_reg[117]  ( .D(o[117]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][117] ) );
  DFF \zreg_reg[118]  ( .D(o[118]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][118] ) );
  DFF \zreg_reg[119]  ( .D(o[119]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][119] ) );
  DFF \zreg_reg[120]  ( .D(o[120]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][120] ) );
  DFF \zreg_reg[121]  ( .D(o[121]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][121] ) );
  DFF \zreg_reg[122]  ( .D(o[122]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][122] ) );
  DFF \zreg_reg[123]  ( .D(o[123]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][123] ) );
  DFF \zreg_reg[124]  ( .D(o[124]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][124] ) );
  DFF \zreg_reg[125]  ( .D(o[125]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][125] ) );
  DFF \zreg_reg[126]  ( .D(o[126]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][126] ) );
  DFF \zreg_reg[127]  ( .D(o[127]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][127] ) );
  DFF \zreg_reg[128]  ( .D(o[128]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][128] ) );
  DFF \zreg_reg[129]  ( .D(o[129]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][129] ) );
  DFF \zreg_reg[130]  ( .D(o[130]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][130] ) );
  DFF \zreg_reg[131]  ( .D(o[131]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][131] ) );
  DFF \zreg_reg[132]  ( .D(o[132]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][132] ) );
  DFF \zreg_reg[133]  ( .D(o[133]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][133] ) );
  DFF \zreg_reg[134]  ( .D(o[134]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][134] ) );
  DFF \zreg_reg[135]  ( .D(o[135]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][135] ) );
  DFF \zreg_reg[136]  ( .D(o[136]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][136] ) );
  DFF \zreg_reg[137]  ( .D(o[137]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][137] ) );
  DFF \zreg_reg[138]  ( .D(o[138]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][138] ) );
  DFF \zreg_reg[139]  ( .D(o[139]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][139] ) );
  DFF \zreg_reg[140]  ( .D(o[140]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][140] ) );
  DFF \zreg_reg[141]  ( .D(o[141]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][141] ) );
  DFF \zreg_reg[142]  ( .D(o[142]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][142] ) );
  DFF \zreg_reg[143]  ( .D(o[143]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][143] ) );
  DFF \zreg_reg[144]  ( .D(o[144]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][144] ) );
  DFF \zreg_reg[145]  ( .D(o[145]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][145] ) );
  DFF \zreg_reg[146]  ( .D(o[146]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][146] ) );
  DFF \zreg_reg[147]  ( .D(o[147]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][147] ) );
  DFF \zreg_reg[148]  ( .D(o[148]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][148] ) );
  DFF \zreg_reg[149]  ( .D(o[149]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][149] ) );
  DFF \zreg_reg[150]  ( .D(o[150]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][150] ) );
  DFF \zreg_reg[151]  ( .D(o[151]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][151] ) );
  DFF \zreg_reg[152]  ( .D(o[152]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][152] ) );
  DFF \zreg_reg[153]  ( .D(o[153]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][153] ) );
  DFF \zreg_reg[154]  ( .D(o[154]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][154] ) );
  DFF \zreg_reg[155]  ( .D(o[155]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][155] ) );
  DFF \zreg_reg[156]  ( .D(o[156]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][156] ) );
  DFF \zreg_reg[157]  ( .D(o[157]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][157] ) );
  DFF \zreg_reg[158]  ( .D(o[158]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][158] ) );
  DFF \zreg_reg[159]  ( .D(o[159]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][159] ) );
  DFF \zreg_reg[160]  ( .D(o[160]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][160] ) );
  DFF \zreg_reg[161]  ( .D(o[161]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][161] ) );
  DFF \zreg_reg[162]  ( .D(o[162]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][162] ) );
  DFF \zreg_reg[163]  ( .D(o[163]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][163] ) );
  DFF \zreg_reg[164]  ( .D(o[164]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][164] ) );
  DFF \zreg_reg[165]  ( .D(o[165]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][165] ) );
  DFF \zreg_reg[166]  ( .D(o[166]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][166] ) );
  DFF \zreg_reg[167]  ( .D(o[167]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][167] ) );
  DFF \zreg_reg[168]  ( .D(o[168]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][168] ) );
  DFF \zreg_reg[169]  ( .D(o[169]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][169] ) );
  DFF \zreg_reg[170]  ( .D(o[170]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][170] ) );
  DFF \zreg_reg[171]  ( .D(o[171]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][171] ) );
  DFF \zreg_reg[172]  ( .D(o[172]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][172] ) );
  DFF \zreg_reg[173]  ( .D(o[173]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][173] ) );
  DFF \zreg_reg[174]  ( .D(o[174]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][174] ) );
  DFF \zreg_reg[175]  ( .D(o[175]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][175] ) );
  DFF \zreg_reg[176]  ( .D(o[176]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][176] ) );
  DFF \zreg_reg[177]  ( .D(o[177]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][177] ) );
  DFF \zreg_reg[178]  ( .D(o[178]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][178] ) );
  DFF \zreg_reg[179]  ( .D(o[179]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][179] ) );
  DFF \zreg_reg[180]  ( .D(o[180]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][180] ) );
  DFF \zreg_reg[181]  ( .D(o[181]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][181] ) );
  DFF \zreg_reg[182]  ( .D(o[182]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][182] ) );
  DFF \zreg_reg[183]  ( .D(o[183]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][183] ) );
  DFF \zreg_reg[184]  ( .D(o[184]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][184] ) );
  DFF \zreg_reg[185]  ( .D(o[185]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][185] ) );
  DFF \zreg_reg[186]  ( .D(o[186]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][186] ) );
  DFF \zreg_reg[187]  ( .D(o[187]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][187] ) );
  DFF \zreg_reg[188]  ( .D(o[188]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][188] ) );
  DFF \zreg_reg[189]  ( .D(o[189]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][189] ) );
  DFF \zreg_reg[190]  ( .D(o[190]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][190] ) );
  DFF \zreg_reg[191]  ( .D(o[191]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][191] ) );
  DFF \zreg_reg[192]  ( .D(o[192]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][192] ) );
  DFF \zreg_reg[193]  ( .D(o[193]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][193] ) );
  DFF \zreg_reg[194]  ( .D(o[194]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][194] ) );
  DFF \zreg_reg[195]  ( .D(o[195]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][195] ) );
  DFF \zreg_reg[196]  ( .D(o[196]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][196] ) );
  DFF \zreg_reg[197]  ( .D(o[197]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][197] ) );
  DFF \zreg_reg[198]  ( .D(o[198]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][198] ) );
  DFF \zreg_reg[199]  ( .D(o[199]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][199] ) );
  DFF \zreg_reg[200]  ( .D(o[200]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][200] ) );
  DFF \zreg_reg[201]  ( .D(o[201]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][201] ) );
  DFF \zreg_reg[202]  ( .D(o[202]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][202] ) );
  DFF \zreg_reg[203]  ( .D(o[203]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][203] ) );
  DFF \zreg_reg[204]  ( .D(o[204]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][204] ) );
  DFF \zreg_reg[205]  ( .D(o[205]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][205] ) );
  DFF \zreg_reg[206]  ( .D(o[206]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][206] ) );
  DFF \zreg_reg[207]  ( .D(o[207]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][207] ) );
  DFF \zreg_reg[208]  ( .D(o[208]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][208] ) );
  DFF \zreg_reg[209]  ( .D(o[209]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][209] ) );
  DFF \zreg_reg[210]  ( .D(o[210]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][210] ) );
  DFF \zreg_reg[211]  ( .D(o[211]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][211] ) );
  DFF \zreg_reg[212]  ( .D(o[212]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][212] ) );
  DFF \zreg_reg[213]  ( .D(o[213]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][213] ) );
  DFF \zreg_reg[214]  ( .D(o[214]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][214] ) );
  DFF \zreg_reg[215]  ( .D(o[215]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][215] ) );
  DFF \zreg_reg[216]  ( .D(o[216]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][216] ) );
  DFF \zreg_reg[217]  ( .D(o[217]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][217] ) );
  DFF \zreg_reg[218]  ( .D(o[218]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][218] ) );
  DFF \zreg_reg[219]  ( .D(o[219]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][219] ) );
  DFF \zreg_reg[220]  ( .D(o[220]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][220] ) );
  DFF \zreg_reg[221]  ( .D(o[221]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][221] ) );
  DFF \zreg_reg[222]  ( .D(o[222]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][222] ) );
  DFF \zreg_reg[223]  ( .D(o[223]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][223] ) );
  DFF \zreg_reg[224]  ( .D(o[224]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][224] ) );
  DFF \zreg_reg[225]  ( .D(o[225]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][225] ) );
  DFF \zreg_reg[226]  ( .D(o[226]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][226] ) );
  DFF \zreg_reg[227]  ( .D(o[227]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][227] ) );
  DFF \zreg_reg[228]  ( .D(o[228]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][228] ) );
  DFF \zreg_reg[229]  ( .D(o[229]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][229] ) );
  DFF \zreg_reg[230]  ( .D(o[230]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][230] ) );
  DFF \zreg_reg[231]  ( .D(o[231]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][231] ) );
  DFF \zreg_reg[232]  ( .D(o[232]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][232] ) );
  DFF \zreg_reg[233]  ( .D(o[233]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][233] ) );
  DFF \zreg_reg[234]  ( .D(o[234]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][234] ) );
  DFF \zreg_reg[235]  ( .D(o[235]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][235] ) );
  DFF \zreg_reg[236]  ( .D(o[236]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][236] ) );
  DFF \zreg_reg[237]  ( .D(o[237]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][237] ) );
  DFF \zreg_reg[238]  ( .D(o[238]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][238] ) );
  DFF \zreg_reg[239]  ( .D(o[239]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][239] ) );
  DFF \zreg_reg[240]  ( .D(o[240]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][240] ) );
  DFF \zreg_reg[241]  ( .D(o[241]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][241] ) );
  DFF \zreg_reg[242]  ( .D(o[242]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][242] ) );
  DFF \zreg_reg[243]  ( .D(o[243]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][243] ) );
  DFF \zreg_reg[244]  ( .D(o[244]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][244] ) );
  DFF \zreg_reg[245]  ( .D(o[245]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][245] ) );
  DFF \zreg_reg[246]  ( .D(o[246]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][246] ) );
  DFF \zreg_reg[247]  ( .D(o[247]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][247] ) );
  DFF \zreg_reg[248]  ( .D(o[248]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][248] ) );
  DFF \zreg_reg[249]  ( .D(o[249]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][249] ) );
  DFF \zreg_reg[250]  ( .D(o[250]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][250] ) );
  DFF \zreg_reg[251]  ( .D(o[251]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][251] ) );
  DFF \zreg_reg[252]  ( .D(o[252]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][252] ) );
  DFF \zreg_reg[253]  ( .D(o[253]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][253] ) );
  DFF \zreg_reg[254]  ( .D(o[254]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][254] ) );
  DFF \zreg_reg[255]  ( .D(o[255]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][255] ) );
  DFF \zreg_reg[256]  ( .D(o[256]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][256] ) );
  DFF \zreg_reg[257]  ( .D(o[257]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][257] ) );
  DFF \zreg_reg[258]  ( .D(o[258]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][258] ) );
  DFF \zreg_reg[259]  ( .D(o[259]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][259] ) );
  DFF \zreg_reg[260]  ( .D(o[260]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][260] ) );
  DFF \zreg_reg[261]  ( .D(o[261]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][261] ) );
  DFF \zreg_reg[262]  ( .D(o[262]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][262] ) );
  DFF \zreg_reg[263]  ( .D(o[263]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][263] ) );
  DFF \zreg_reg[264]  ( .D(o[264]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][264] ) );
  DFF \zreg_reg[265]  ( .D(o[265]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][265] ) );
  DFF \zreg_reg[266]  ( .D(o[266]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][266] ) );
  DFF \zreg_reg[267]  ( .D(o[267]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][267] ) );
  DFF \zreg_reg[268]  ( .D(o[268]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][268] ) );
  DFF \zreg_reg[269]  ( .D(o[269]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][269] ) );
  DFF \zreg_reg[270]  ( .D(o[270]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][270] ) );
  DFF \zreg_reg[271]  ( .D(o[271]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][271] ) );
  DFF \zreg_reg[272]  ( .D(o[272]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][272] ) );
  DFF \zreg_reg[273]  ( .D(o[273]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][273] ) );
  DFF \zreg_reg[274]  ( .D(o[274]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][274] ) );
  DFF \zreg_reg[275]  ( .D(o[275]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][275] ) );
  DFF \zreg_reg[276]  ( .D(o[276]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][276] ) );
  DFF \zreg_reg[277]  ( .D(o[277]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][277] ) );
  DFF \zreg_reg[278]  ( .D(o[278]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][278] ) );
  DFF \zreg_reg[279]  ( .D(o[279]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][279] ) );
  DFF \zreg_reg[280]  ( .D(o[280]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][280] ) );
  DFF \zreg_reg[281]  ( .D(o[281]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][281] ) );
  DFF \zreg_reg[282]  ( .D(o[282]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][282] ) );
  DFF \zreg_reg[283]  ( .D(o[283]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][283] ) );
  DFF \zreg_reg[284]  ( .D(o[284]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][284] ) );
  DFF \zreg_reg[285]  ( .D(o[285]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][285] ) );
  DFF \zreg_reg[286]  ( .D(o[286]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][286] ) );
  DFF \zreg_reg[287]  ( .D(o[287]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][287] ) );
  DFF \zreg_reg[288]  ( .D(o[288]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][288] ) );
  DFF \zreg_reg[289]  ( .D(o[289]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][289] ) );
  DFF \zreg_reg[290]  ( .D(o[290]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][290] ) );
  DFF \zreg_reg[291]  ( .D(o[291]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][291] ) );
  DFF \zreg_reg[292]  ( .D(o[292]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][292] ) );
  DFF \zreg_reg[293]  ( .D(o[293]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][293] ) );
  DFF \zreg_reg[294]  ( .D(o[294]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][294] ) );
  DFF \zreg_reg[295]  ( .D(o[295]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][295] ) );
  DFF \zreg_reg[296]  ( .D(o[296]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][296] ) );
  DFF \zreg_reg[297]  ( .D(o[297]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][297] ) );
  DFF \zreg_reg[298]  ( .D(o[298]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][298] ) );
  DFF \zreg_reg[299]  ( .D(o[299]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][299] ) );
  DFF \zreg_reg[300]  ( .D(o[300]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][300] ) );
  DFF \zreg_reg[301]  ( .D(o[301]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][301] ) );
  DFF \zreg_reg[302]  ( .D(o[302]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][302] ) );
  DFF \zreg_reg[303]  ( .D(o[303]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][303] ) );
  DFF \zreg_reg[304]  ( .D(o[304]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][304] ) );
  DFF \zreg_reg[305]  ( .D(o[305]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][305] ) );
  DFF \zreg_reg[306]  ( .D(o[306]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][306] ) );
  DFF \zreg_reg[307]  ( .D(o[307]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][307] ) );
  DFF \zreg_reg[308]  ( .D(o[308]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][308] ) );
  DFF \zreg_reg[309]  ( .D(o[309]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][309] ) );
  DFF \zreg_reg[310]  ( .D(o[310]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][310] ) );
  DFF \zreg_reg[311]  ( .D(o[311]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][311] ) );
  DFF \zreg_reg[312]  ( .D(o[312]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][312] ) );
  DFF \zreg_reg[313]  ( .D(o[313]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][313] ) );
  DFF \zreg_reg[314]  ( .D(o[314]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][314] ) );
  DFF \zreg_reg[315]  ( .D(o[315]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][315] ) );
  DFF \zreg_reg[316]  ( .D(o[316]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][316] ) );
  DFF \zreg_reg[317]  ( .D(o[317]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][317] ) );
  DFF \zreg_reg[318]  ( .D(o[318]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][318] ) );
  DFF \zreg_reg[319]  ( .D(o[319]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][319] ) );
  DFF \zreg_reg[320]  ( .D(o[320]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][320] ) );
  DFF \zreg_reg[321]  ( .D(o[321]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][321] ) );
  DFF \zreg_reg[322]  ( .D(o[322]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][322] ) );
  DFF \zreg_reg[323]  ( .D(o[323]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][323] ) );
  DFF \zreg_reg[324]  ( .D(o[324]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][324] ) );
  DFF \zreg_reg[325]  ( .D(o[325]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][325] ) );
  DFF \zreg_reg[326]  ( .D(o[326]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][326] ) );
  DFF \zreg_reg[327]  ( .D(o[327]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][327] ) );
  DFF \zreg_reg[328]  ( .D(o[328]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][328] ) );
  DFF \zreg_reg[329]  ( .D(o[329]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][329] ) );
  DFF \zreg_reg[330]  ( .D(o[330]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][330] ) );
  DFF \zreg_reg[331]  ( .D(o[331]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][331] ) );
  DFF \zreg_reg[332]  ( .D(o[332]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][332] ) );
  DFF \zreg_reg[333]  ( .D(o[333]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][333] ) );
  DFF \zreg_reg[334]  ( .D(o[334]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][334] ) );
  DFF \zreg_reg[335]  ( .D(o[335]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][335] ) );
  DFF \zreg_reg[336]  ( .D(o[336]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][336] ) );
  DFF \zreg_reg[337]  ( .D(o[337]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][337] ) );
  DFF \zreg_reg[338]  ( .D(o[338]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][338] ) );
  DFF \zreg_reg[339]  ( .D(o[339]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][339] ) );
  DFF \zreg_reg[340]  ( .D(o[340]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][340] ) );
  DFF \zreg_reg[341]  ( .D(o[341]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][341] ) );
  DFF \zreg_reg[342]  ( .D(o[342]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][342] ) );
  DFF \zreg_reg[343]  ( .D(o[343]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][343] ) );
  DFF \zreg_reg[344]  ( .D(o[344]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][344] ) );
  DFF \zreg_reg[345]  ( .D(o[345]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][345] ) );
  DFF \zreg_reg[346]  ( .D(o[346]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][346] ) );
  DFF \zreg_reg[347]  ( .D(o[347]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][347] ) );
  DFF \zreg_reg[348]  ( .D(o[348]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][348] ) );
  DFF \zreg_reg[349]  ( .D(o[349]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][349] ) );
  DFF \zreg_reg[350]  ( .D(o[350]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][350] ) );
  DFF \zreg_reg[351]  ( .D(o[351]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][351] ) );
  DFF \zreg_reg[352]  ( .D(o[352]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][352] ) );
  DFF \zreg_reg[353]  ( .D(o[353]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][353] ) );
  DFF \zreg_reg[354]  ( .D(o[354]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][354] ) );
  DFF \zreg_reg[355]  ( .D(o[355]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][355] ) );
  DFF \zreg_reg[356]  ( .D(o[356]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][356] ) );
  DFF \zreg_reg[357]  ( .D(o[357]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][357] ) );
  DFF \zreg_reg[358]  ( .D(o[358]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][358] ) );
  DFF \zreg_reg[359]  ( .D(o[359]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][359] ) );
  DFF \zreg_reg[360]  ( .D(o[360]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][360] ) );
  DFF \zreg_reg[361]  ( .D(o[361]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][361] ) );
  DFF \zreg_reg[362]  ( .D(o[362]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][362] ) );
  DFF \zreg_reg[363]  ( .D(o[363]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][363] ) );
  DFF \zreg_reg[364]  ( .D(o[364]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][364] ) );
  DFF \zreg_reg[365]  ( .D(o[365]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][365] ) );
  DFF \zreg_reg[366]  ( .D(o[366]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][366] ) );
  DFF \zreg_reg[367]  ( .D(o[367]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][367] ) );
  DFF \zreg_reg[368]  ( .D(o[368]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][368] ) );
  DFF \zreg_reg[369]  ( .D(o[369]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][369] ) );
  DFF \zreg_reg[370]  ( .D(o[370]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][370] ) );
  DFF \zreg_reg[371]  ( .D(o[371]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][371] ) );
  DFF \zreg_reg[372]  ( .D(o[372]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][372] ) );
  DFF \zreg_reg[373]  ( .D(o[373]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][373] ) );
  DFF \zreg_reg[374]  ( .D(o[374]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][374] ) );
  DFF \zreg_reg[375]  ( .D(o[375]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][375] ) );
  DFF \zreg_reg[376]  ( .D(o[376]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][376] ) );
  DFF \zreg_reg[377]  ( .D(o[377]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][377] ) );
  DFF \zreg_reg[378]  ( .D(o[378]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][378] ) );
  DFF \zreg_reg[379]  ( .D(o[379]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][379] ) );
  DFF \zreg_reg[380]  ( .D(o[380]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][380] ) );
  DFF \zreg_reg[381]  ( .D(o[381]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][381] ) );
  DFF \zreg_reg[382]  ( .D(o[382]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][382] ) );
  DFF \zreg_reg[383]  ( .D(o[383]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][383] ) );
  DFF \zreg_reg[384]  ( .D(o[384]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][384] ) );
  DFF \zreg_reg[385]  ( .D(o[385]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][385] ) );
  DFF \zreg_reg[386]  ( .D(o[386]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][386] ) );
  DFF \zreg_reg[387]  ( .D(o[387]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][387] ) );
  DFF \zreg_reg[388]  ( .D(o[388]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][388] ) );
  DFF \zreg_reg[389]  ( .D(o[389]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][389] ) );
  DFF \zreg_reg[390]  ( .D(o[390]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][390] ) );
  DFF \zreg_reg[391]  ( .D(o[391]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][391] ) );
  DFF \zreg_reg[392]  ( .D(o[392]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][392] ) );
  DFF \zreg_reg[393]  ( .D(o[393]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][393] ) );
  DFF \zreg_reg[394]  ( .D(o[394]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][394] ) );
  DFF \zreg_reg[395]  ( .D(o[395]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][395] ) );
  DFF \zreg_reg[396]  ( .D(o[396]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][396] ) );
  DFF \zreg_reg[397]  ( .D(o[397]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][397] ) );
  DFF \zreg_reg[398]  ( .D(o[398]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][398] ) );
  DFF \zreg_reg[399]  ( .D(o[399]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][399] ) );
  DFF \zreg_reg[400]  ( .D(o[400]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][400] ) );
  DFF \zreg_reg[401]  ( .D(o[401]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][401] ) );
  DFF \zreg_reg[402]  ( .D(o[402]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][402] ) );
  DFF \zreg_reg[403]  ( .D(o[403]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][403] ) );
  DFF \zreg_reg[404]  ( .D(o[404]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][404] ) );
  DFF \zreg_reg[405]  ( .D(o[405]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][405] ) );
  DFF \zreg_reg[406]  ( .D(o[406]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][406] ) );
  DFF \zreg_reg[407]  ( .D(o[407]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][407] ) );
  DFF \zreg_reg[408]  ( .D(o[408]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][408] ) );
  DFF \zreg_reg[409]  ( .D(o[409]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][409] ) );
  DFF \zreg_reg[410]  ( .D(o[410]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][410] ) );
  DFF \zreg_reg[411]  ( .D(o[411]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][411] ) );
  DFF \zreg_reg[412]  ( .D(o[412]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][412] ) );
  DFF \zreg_reg[413]  ( .D(o[413]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][413] ) );
  DFF \zreg_reg[414]  ( .D(o[414]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][414] ) );
  DFF \zreg_reg[415]  ( .D(o[415]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][415] ) );
  DFF \zreg_reg[416]  ( .D(o[416]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][416] ) );
  DFF \zreg_reg[417]  ( .D(o[417]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][417] ) );
  DFF \zreg_reg[418]  ( .D(o[418]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][418] ) );
  DFF \zreg_reg[419]  ( .D(o[419]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][419] ) );
  DFF \zreg_reg[420]  ( .D(o[420]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][420] ) );
  DFF \zreg_reg[421]  ( .D(o[421]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][421] ) );
  DFF \zreg_reg[422]  ( .D(o[422]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][422] ) );
  DFF \zreg_reg[423]  ( .D(o[423]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][423] ) );
  DFF \zreg_reg[424]  ( .D(o[424]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][424] ) );
  DFF \zreg_reg[425]  ( .D(o[425]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][425] ) );
  DFF \zreg_reg[426]  ( .D(o[426]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][426] ) );
  DFF \zreg_reg[427]  ( .D(o[427]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][427] ) );
  DFF \zreg_reg[428]  ( .D(o[428]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][428] ) );
  DFF \zreg_reg[429]  ( .D(o[429]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][429] ) );
  DFF \zreg_reg[430]  ( .D(o[430]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][430] ) );
  DFF \zreg_reg[431]  ( .D(o[431]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][431] ) );
  DFF \zreg_reg[432]  ( .D(o[432]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][432] ) );
  DFF \zreg_reg[433]  ( .D(o[433]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][433] ) );
  DFF \zreg_reg[434]  ( .D(o[434]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][434] ) );
  DFF \zreg_reg[435]  ( .D(o[435]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][435] ) );
  DFF \zreg_reg[436]  ( .D(o[436]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][436] ) );
  DFF \zreg_reg[437]  ( .D(o[437]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][437] ) );
  DFF \zreg_reg[438]  ( .D(o[438]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][438] ) );
  DFF \zreg_reg[439]  ( .D(o[439]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][439] ) );
  DFF \zreg_reg[440]  ( .D(o[440]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][440] ) );
  DFF \zreg_reg[441]  ( .D(o[441]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][441] ) );
  DFF \zreg_reg[442]  ( .D(o[442]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][442] ) );
  DFF \zreg_reg[443]  ( .D(o[443]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][443] ) );
  DFF \zreg_reg[444]  ( .D(o[444]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][444] ) );
  DFF \zreg_reg[445]  ( .D(o[445]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][445] ) );
  DFF \zreg_reg[446]  ( .D(o[446]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][446] ) );
  DFF \zreg_reg[447]  ( .D(o[447]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][447] ) );
  DFF \zreg_reg[448]  ( .D(o[448]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][448] ) );
  DFF \zreg_reg[449]  ( .D(o[449]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][449] ) );
  DFF \zreg_reg[450]  ( .D(o[450]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][450] ) );
  DFF \zreg_reg[451]  ( .D(o[451]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][451] ) );
  DFF \zreg_reg[452]  ( .D(o[452]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][452] ) );
  DFF \zreg_reg[453]  ( .D(o[453]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][453] ) );
  DFF \zreg_reg[454]  ( .D(o[454]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][454] ) );
  DFF \zreg_reg[455]  ( .D(o[455]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][455] ) );
  DFF \zreg_reg[456]  ( .D(o[456]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][456] ) );
  DFF \zreg_reg[457]  ( .D(o[457]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][457] ) );
  DFF \zreg_reg[458]  ( .D(o[458]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][458] ) );
  DFF \zreg_reg[459]  ( .D(o[459]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][459] ) );
  DFF \zreg_reg[460]  ( .D(o[460]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][460] ) );
  DFF \zreg_reg[461]  ( .D(o[461]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][461] ) );
  DFF \zreg_reg[462]  ( .D(o[462]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][462] ) );
  DFF \zreg_reg[463]  ( .D(o[463]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][463] ) );
  DFF \zreg_reg[464]  ( .D(o[464]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][464] ) );
  DFF \zreg_reg[465]  ( .D(o[465]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][465] ) );
  DFF \zreg_reg[466]  ( .D(o[466]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][466] ) );
  DFF \zreg_reg[467]  ( .D(o[467]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][467] ) );
  DFF \zreg_reg[468]  ( .D(o[468]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][468] ) );
  DFF \zreg_reg[469]  ( .D(o[469]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][469] ) );
  DFF \zreg_reg[470]  ( .D(o[470]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][470] ) );
  DFF \zreg_reg[471]  ( .D(o[471]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][471] ) );
  DFF \zreg_reg[472]  ( .D(o[472]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][472] ) );
  DFF \zreg_reg[473]  ( .D(o[473]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][473] ) );
  DFF \zreg_reg[474]  ( .D(o[474]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][474] ) );
  DFF \zreg_reg[475]  ( .D(o[475]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][475] ) );
  DFF \zreg_reg[476]  ( .D(o[476]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][476] ) );
  DFF \zreg_reg[477]  ( .D(o[477]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][477] ) );
  DFF \zreg_reg[478]  ( .D(o[478]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][478] ) );
  DFF \zreg_reg[479]  ( .D(o[479]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][479] ) );
  DFF \zreg_reg[480]  ( .D(o[480]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][480] ) );
  DFF \zreg_reg[481]  ( .D(o[481]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][481] ) );
  DFF \zreg_reg[482]  ( .D(o[482]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][482] ) );
  DFF \zreg_reg[483]  ( .D(o[483]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][483] ) );
  DFF \zreg_reg[484]  ( .D(o[484]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][484] ) );
  DFF \zreg_reg[485]  ( .D(o[485]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][485] ) );
  DFF \zreg_reg[486]  ( .D(o[486]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][486] ) );
  DFF \zreg_reg[487]  ( .D(o[487]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][487] ) );
  DFF \zreg_reg[488]  ( .D(o[488]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][488] ) );
  DFF \zreg_reg[489]  ( .D(o[489]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][489] ) );
  DFF \zreg_reg[490]  ( .D(o[490]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][490] ) );
  DFF \zreg_reg[491]  ( .D(o[491]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][491] ) );
  DFF \zreg_reg[492]  ( .D(o[492]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][492] ) );
  DFF \zreg_reg[493]  ( .D(o[493]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][493] ) );
  DFF \zreg_reg[494]  ( .D(o[494]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][494] ) );
  DFF \zreg_reg[495]  ( .D(o[495]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][495] ) );
  DFF \zreg_reg[496]  ( .D(o[496]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][496] ) );
  DFF \zreg_reg[497]  ( .D(o[497]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][497] ) );
  DFF \zreg_reg[498]  ( .D(o[498]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][498] ) );
  DFF \zreg_reg[499]  ( .D(o[499]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][499] ) );
  DFF \zreg_reg[500]  ( .D(o[500]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][500] ) );
  DFF \zreg_reg[501]  ( .D(o[501]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][501] ) );
  DFF \zreg_reg[502]  ( .D(o[502]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][502] ) );
  DFF \zreg_reg[503]  ( .D(o[503]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][503] ) );
  DFF \zreg_reg[504]  ( .D(o[504]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][504] ) );
  DFF \zreg_reg[505]  ( .D(o[505]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][505] ) );
  DFF \zreg_reg[506]  ( .D(o[506]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][506] ) );
  DFF \zreg_reg[507]  ( .D(o[507]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][507] ) );
  DFF \zreg_reg[508]  ( .D(o[508]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][508] ) );
  DFF \zreg_reg[509]  ( .D(o[509]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][509] ) );
  DFF \zreg_reg[510]  ( .D(o[510]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][510] ) );
  DFF \zreg_reg[511]  ( .D(o[511]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][511] ) );
  DFF \zreg_reg[512]  ( .D(o[512]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][512] ) );
  DFF \zreg_reg[513]  ( .D(o[513]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][513] ) );
  DFF \zreg_reg[514]  ( .D(o[514]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][514] ) );
  DFF \zreg_reg[515]  ( .D(o[515]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][515] ) );
  DFF \zreg_reg[516]  ( .D(o[516]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][516] ) );
  DFF \zreg_reg[517]  ( .D(o[517]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][517] ) );
  DFF \zreg_reg[518]  ( .D(o[518]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][518] ) );
  DFF \zreg_reg[519]  ( .D(o[519]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][519] ) );
  DFF \zreg_reg[520]  ( .D(o[520]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][520] ) );
  DFF \zreg_reg[521]  ( .D(o[521]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][521] ) );
  DFF \zreg_reg[522]  ( .D(o[522]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][522] ) );
  DFF \zreg_reg[523]  ( .D(o[523]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][523] ) );
  DFF \zreg_reg[524]  ( .D(o[524]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][524] ) );
  DFF \zreg_reg[525]  ( .D(o[525]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][525] ) );
  DFF \zreg_reg[526]  ( .D(o[526]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][526] ) );
  DFF \zreg_reg[527]  ( .D(o[527]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][527] ) );
  DFF \zreg_reg[528]  ( .D(o[528]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][528] ) );
  DFF \zreg_reg[529]  ( .D(o[529]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][529] ) );
  DFF \zreg_reg[530]  ( .D(o[530]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][530] ) );
  DFF \zreg_reg[531]  ( .D(o[531]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][531] ) );
  DFF \zreg_reg[532]  ( .D(o[532]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][532] ) );
  DFF \zreg_reg[533]  ( .D(o[533]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][533] ) );
  DFF \zreg_reg[534]  ( .D(o[534]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][534] ) );
  DFF \zreg_reg[535]  ( .D(o[535]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][535] ) );
  DFF \zreg_reg[536]  ( .D(o[536]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][536] ) );
  DFF \zreg_reg[537]  ( .D(o[537]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][537] ) );
  DFF \zreg_reg[538]  ( .D(o[538]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][538] ) );
  DFF \zreg_reg[539]  ( .D(o[539]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][539] ) );
  DFF \zreg_reg[540]  ( .D(o[540]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][540] ) );
  DFF \zreg_reg[541]  ( .D(o[541]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][541] ) );
  DFF \zreg_reg[542]  ( .D(o[542]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][542] ) );
  DFF \zreg_reg[543]  ( .D(o[543]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][543] ) );
  DFF \zreg_reg[544]  ( .D(o[544]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][544] ) );
  DFF \zreg_reg[545]  ( .D(o[545]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][545] ) );
  DFF \zreg_reg[546]  ( .D(o[546]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][546] ) );
  DFF \zreg_reg[547]  ( .D(o[547]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][547] ) );
  DFF \zreg_reg[548]  ( .D(o[548]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][548] ) );
  DFF \zreg_reg[549]  ( .D(o[549]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][549] ) );
  DFF \zreg_reg[550]  ( .D(o[550]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][550] ) );
  DFF \zreg_reg[551]  ( .D(o[551]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][551] ) );
  DFF \zreg_reg[552]  ( .D(o[552]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][552] ) );
  DFF \zreg_reg[553]  ( .D(o[553]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][553] ) );
  DFF \zreg_reg[554]  ( .D(o[554]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][554] ) );
  DFF \zreg_reg[555]  ( .D(o[555]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][555] ) );
  DFF \zreg_reg[556]  ( .D(o[556]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][556] ) );
  DFF \zreg_reg[557]  ( .D(o[557]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][557] ) );
  DFF \zreg_reg[558]  ( .D(o[558]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][558] ) );
  DFF \zreg_reg[559]  ( .D(o[559]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][559] ) );
  DFF \zreg_reg[560]  ( .D(o[560]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][560] ) );
  DFF \zreg_reg[561]  ( .D(o[561]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][561] ) );
  DFF \zreg_reg[562]  ( .D(o[562]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][562] ) );
  DFF \zreg_reg[563]  ( .D(o[563]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][563] ) );
  DFF \zreg_reg[564]  ( .D(o[564]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][564] ) );
  DFF \zreg_reg[565]  ( .D(o[565]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][565] ) );
  DFF \zreg_reg[566]  ( .D(o[566]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][566] ) );
  DFF \zreg_reg[567]  ( .D(o[567]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][567] ) );
  DFF \zreg_reg[568]  ( .D(o[568]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][568] ) );
  DFF \zreg_reg[569]  ( .D(o[569]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][569] ) );
  DFF \zreg_reg[570]  ( .D(o[570]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][570] ) );
  DFF \zreg_reg[571]  ( .D(o[571]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][571] ) );
  DFF \zreg_reg[572]  ( .D(o[572]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][572] ) );
  DFF \zreg_reg[573]  ( .D(o[573]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][573] ) );
  DFF \zreg_reg[574]  ( .D(o[574]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][574] ) );
  DFF \zreg_reg[575]  ( .D(o[575]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][575] ) );
  DFF \zreg_reg[576]  ( .D(o[576]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][576] ) );
  DFF \zreg_reg[577]  ( .D(o[577]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][577] ) );
  DFF \zreg_reg[578]  ( .D(o[578]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][578] ) );
  DFF \zreg_reg[579]  ( .D(o[579]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][579] ) );
  DFF \zreg_reg[580]  ( .D(o[580]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][580] ) );
  DFF \zreg_reg[581]  ( .D(o[581]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][581] ) );
  DFF \zreg_reg[582]  ( .D(o[582]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][582] ) );
  DFF \zreg_reg[583]  ( .D(o[583]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][583] ) );
  DFF \zreg_reg[584]  ( .D(o[584]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][584] ) );
  DFF \zreg_reg[585]  ( .D(o[585]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][585] ) );
  DFF \zreg_reg[586]  ( .D(o[586]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][586] ) );
  DFF \zreg_reg[587]  ( .D(o[587]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][587] ) );
  DFF \zreg_reg[588]  ( .D(o[588]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][588] ) );
  DFF \zreg_reg[589]  ( .D(o[589]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][589] ) );
  DFF \zreg_reg[590]  ( .D(o[590]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][590] ) );
  DFF \zreg_reg[591]  ( .D(o[591]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][591] ) );
  DFF \zreg_reg[592]  ( .D(o[592]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][592] ) );
  DFF \zreg_reg[593]  ( .D(o[593]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][593] ) );
  DFF \zreg_reg[594]  ( .D(o[594]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][594] ) );
  DFF \zreg_reg[595]  ( .D(o[595]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][595] ) );
  DFF \zreg_reg[596]  ( .D(o[596]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][596] ) );
  DFF \zreg_reg[597]  ( .D(o[597]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][597] ) );
  DFF \zreg_reg[598]  ( .D(o[598]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][598] ) );
  DFF \zreg_reg[599]  ( .D(o[599]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][599] ) );
  DFF \zreg_reg[600]  ( .D(o[600]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][600] ) );
  DFF \zreg_reg[601]  ( .D(o[601]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][601] ) );
  DFF \zreg_reg[602]  ( .D(o[602]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][602] ) );
  DFF \zreg_reg[603]  ( .D(o[603]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][603] ) );
  DFF \zreg_reg[604]  ( .D(o[604]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][604] ) );
  DFF \zreg_reg[605]  ( .D(o[605]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][605] ) );
  DFF \zreg_reg[606]  ( .D(o[606]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][606] ) );
  DFF \zreg_reg[607]  ( .D(o[607]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][607] ) );
  DFF \zreg_reg[608]  ( .D(o[608]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][608] ) );
  DFF \zreg_reg[609]  ( .D(o[609]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][609] ) );
  DFF \zreg_reg[610]  ( .D(o[610]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][610] ) );
  DFF \zreg_reg[611]  ( .D(o[611]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][611] ) );
  DFF \zreg_reg[612]  ( .D(o[612]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][612] ) );
  DFF \zreg_reg[613]  ( .D(o[613]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][613] ) );
  DFF \zreg_reg[614]  ( .D(o[614]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][614] ) );
  DFF \zreg_reg[615]  ( .D(o[615]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][615] ) );
  DFF \zreg_reg[616]  ( .D(o[616]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][616] ) );
  DFF \zreg_reg[617]  ( .D(o[617]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][617] ) );
  DFF \zreg_reg[618]  ( .D(o[618]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][618] ) );
  DFF \zreg_reg[619]  ( .D(o[619]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][619] ) );
  DFF \zreg_reg[620]  ( .D(o[620]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][620] ) );
  DFF \zreg_reg[621]  ( .D(o[621]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][621] ) );
  DFF \zreg_reg[622]  ( .D(o[622]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][622] ) );
  DFF \zreg_reg[623]  ( .D(o[623]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][623] ) );
  DFF \zreg_reg[624]  ( .D(o[624]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][624] ) );
  DFF \zreg_reg[625]  ( .D(o[625]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][625] ) );
  DFF \zreg_reg[626]  ( .D(o[626]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][626] ) );
  DFF \zreg_reg[627]  ( .D(o[627]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][627] ) );
  DFF \zreg_reg[628]  ( .D(o[628]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][628] ) );
  DFF \zreg_reg[629]  ( .D(o[629]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][629] ) );
  DFF \zreg_reg[630]  ( .D(o[630]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][630] ) );
  DFF \zreg_reg[631]  ( .D(o[631]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][631] ) );
  DFF \zreg_reg[632]  ( .D(o[632]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][632] ) );
  DFF \zreg_reg[633]  ( .D(o[633]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][633] ) );
  DFF \zreg_reg[634]  ( .D(o[634]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][634] ) );
  DFF \zreg_reg[635]  ( .D(o[635]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][635] ) );
  DFF \zreg_reg[636]  ( .D(o[636]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][636] ) );
  DFF \zreg_reg[637]  ( .D(o[637]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][637] ) );
  DFF \zreg_reg[638]  ( .D(o[638]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][638] ) );
  DFF \zreg_reg[639]  ( .D(o[639]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][639] ) );
  DFF \zreg_reg[640]  ( .D(o[640]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][640] ) );
  DFF \zreg_reg[641]  ( .D(o[641]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][641] ) );
  DFF \zreg_reg[642]  ( .D(o[642]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][642] ) );
  DFF \zreg_reg[643]  ( .D(o[643]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][643] ) );
  DFF \zreg_reg[644]  ( .D(o[644]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][644] ) );
  DFF \zreg_reg[645]  ( .D(o[645]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][645] ) );
  DFF \zreg_reg[646]  ( .D(o[646]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][646] ) );
  DFF \zreg_reg[647]  ( .D(o[647]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][647] ) );
  DFF \zreg_reg[648]  ( .D(o[648]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][648] ) );
  DFF \zreg_reg[649]  ( .D(o[649]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][649] ) );
  DFF \zreg_reg[650]  ( .D(o[650]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][650] ) );
  DFF \zreg_reg[651]  ( .D(o[651]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][651] ) );
  DFF \zreg_reg[652]  ( .D(o[652]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][652] ) );
  DFF \zreg_reg[653]  ( .D(o[653]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][653] ) );
  DFF \zreg_reg[654]  ( .D(o[654]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][654] ) );
  DFF \zreg_reg[655]  ( .D(o[655]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][655] ) );
  DFF \zreg_reg[656]  ( .D(o[656]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][656] ) );
  DFF \zreg_reg[657]  ( .D(o[657]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][657] ) );
  DFF \zreg_reg[658]  ( .D(o[658]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][658] ) );
  DFF \zreg_reg[659]  ( .D(o[659]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][659] ) );
  DFF \zreg_reg[660]  ( .D(o[660]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][660] ) );
  DFF \zreg_reg[661]  ( .D(o[661]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][661] ) );
  DFF \zreg_reg[662]  ( .D(o[662]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][662] ) );
  DFF \zreg_reg[663]  ( .D(o[663]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][663] ) );
  DFF \zreg_reg[664]  ( .D(o[664]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][664] ) );
  DFF \zreg_reg[665]  ( .D(o[665]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][665] ) );
  DFF \zreg_reg[666]  ( .D(o[666]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][666] ) );
  DFF \zreg_reg[667]  ( .D(o[667]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][667] ) );
  DFF \zreg_reg[668]  ( .D(o[668]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][668] ) );
  DFF \zreg_reg[669]  ( .D(o[669]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][669] ) );
  DFF \zreg_reg[670]  ( .D(o[670]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][670] ) );
  DFF \zreg_reg[671]  ( .D(o[671]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][671] ) );
  DFF \zreg_reg[672]  ( .D(o[672]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][672] ) );
  DFF \zreg_reg[673]  ( .D(o[673]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][673] ) );
  DFF \zreg_reg[674]  ( .D(o[674]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][674] ) );
  DFF \zreg_reg[675]  ( .D(o[675]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][675] ) );
  DFF \zreg_reg[676]  ( .D(o[676]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][676] ) );
  DFF \zreg_reg[677]  ( .D(o[677]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][677] ) );
  DFF \zreg_reg[678]  ( .D(o[678]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][678] ) );
  DFF \zreg_reg[679]  ( .D(o[679]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][679] ) );
  DFF \zreg_reg[680]  ( .D(o[680]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][680] ) );
  DFF \zreg_reg[681]  ( .D(o[681]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][681] ) );
  DFF \zreg_reg[682]  ( .D(o[682]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][682] ) );
  DFF \zreg_reg[683]  ( .D(o[683]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][683] ) );
  DFF \zreg_reg[684]  ( .D(o[684]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][684] ) );
  DFF \zreg_reg[685]  ( .D(o[685]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][685] ) );
  DFF \zreg_reg[686]  ( .D(o[686]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][686] ) );
  DFF \zreg_reg[687]  ( .D(o[687]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][687] ) );
  DFF \zreg_reg[688]  ( .D(o[688]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][688] ) );
  DFF \zreg_reg[689]  ( .D(o[689]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][689] ) );
  DFF \zreg_reg[690]  ( .D(o[690]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][690] ) );
  DFF \zreg_reg[691]  ( .D(o[691]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][691] ) );
  DFF \zreg_reg[692]  ( .D(o[692]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][692] ) );
  DFF \zreg_reg[693]  ( .D(o[693]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][693] ) );
  DFF \zreg_reg[694]  ( .D(o[694]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][694] ) );
  DFF \zreg_reg[695]  ( .D(o[695]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][695] ) );
  DFF \zreg_reg[696]  ( .D(o[696]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][696] ) );
  DFF \zreg_reg[697]  ( .D(o[697]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][697] ) );
  DFF \zreg_reg[698]  ( .D(o[698]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][698] ) );
  DFF \zreg_reg[699]  ( .D(o[699]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][699] ) );
  DFF \zreg_reg[700]  ( .D(o[700]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][700] ) );
  DFF \zreg_reg[701]  ( .D(o[701]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][701] ) );
  DFF \zreg_reg[702]  ( .D(o[702]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][702] ) );
  DFF \zreg_reg[703]  ( .D(o[703]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][703] ) );
  DFF \zreg_reg[704]  ( .D(o[704]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][704] ) );
  DFF \zreg_reg[705]  ( .D(o[705]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][705] ) );
  DFF \zreg_reg[706]  ( .D(o[706]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][706] ) );
  DFF \zreg_reg[707]  ( .D(o[707]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][707] ) );
  DFF \zreg_reg[708]  ( .D(o[708]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][708] ) );
  DFF \zreg_reg[709]  ( .D(o[709]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][709] ) );
  DFF \zreg_reg[710]  ( .D(o[710]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][710] ) );
  DFF \zreg_reg[711]  ( .D(o[711]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][711] ) );
  DFF \zreg_reg[712]  ( .D(o[712]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][712] ) );
  DFF \zreg_reg[713]  ( .D(o[713]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][713] ) );
  DFF \zreg_reg[714]  ( .D(o[714]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][714] ) );
  DFF \zreg_reg[715]  ( .D(o[715]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][715] ) );
  DFF \zreg_reg[716]  ( .D(o[716]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][716] ) );
  DFF \zreg_reg[717]  ( .D(o[717]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][717] ) );
  DFF \zreg_reg[718]  ( .D(o[718]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][718] ) );
  DFF \zreg_reg[719]  ( .D(o[719]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][719] ) );
  DFF \zreg_reg[720]  ( .D(o[720]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][720] ) );
  DFF \zreg_reg[721]  ( .D(o[721]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][721] ) );
  DFF \zreg_reg[722]  ( .D(o[722]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][722] ) );
  DFF \zreg_reg[723]  ( .D(o[723]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][723] ) );
  DFF \zreg_reg[724]  ( .D(o[724]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][724] ) );
  DFF \zreg_reg[725]  ( .D(o[725]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][725] ) );
  DFF \zreg_reg[726]  ( .D(o[726]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][726] ) );
  DFF \zreg_reg[727]  ( .D(o[727]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][727] ) );
  DFF \zreg_reg[728]  ( .D(o[728]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][728] ) );
  DFF \zreg_reg[729]  ( .D(o[729]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][729] ) );
  DFF \zreg_reg[730]  ( .D(o[730]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][730] ) );
  DFF \zreg_reg[731]  ( .D(o[731]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][731] ) );
  DFF \zreg_reg[732]  ( .D(o[732]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][732] ) );
  DFF \zreg_reg[733]  ( .D(o[733]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][733] ) );
  DFF \zreg_reg[734]  ( .D(o[734]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][734] ) );
  DFF \zreg_reg[735]  ( .D(o[735]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][735] ) );
  DFF \zreg_reg[736]  ( .D(o[736]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][736] ) );
  DFF \zreg_reg[737]  ( .D(o[737]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][737] ) );
  DFF \zreg_reg[738]  ( .D(o[738]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][738] ) );
  DFF \zreg_reg[739]  ( .D(o[739]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][739] ) );
  DFF \zreg_reg[740]  ( .D(o[740]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][740] ) );
  DFF \zreg_reg[741]  ( .D(o[741]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][741] ) );
  DFF \zreg_reg[742]  ( .D(o[742]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][742] ) );
  DFF \zreg_reg[743]  ( .D(o[743]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][743] ) );
  DFF \zreg_reg[744]  ( .D(o[744]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][744] ) );
  DFF \zreg_reg[745]  ( .D(o[745]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][745] ) );
  DFF \zreg_reg[746]  ( .D(o[746]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][746] ) );
  DFF \zreg_reg[747]  ( .D(o[747]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][747] ) );
  DFF \zreg_reg[748]  ( .D(o[748]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][748] ) );
  DFF \zreg_reg[749]  ( .D(o[749]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][749] ) );
  DFF \zreg_reg[750]  ( .D(o[750]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][750] ) );
  DFF \zreg_reg[751]  ( .D(o[751]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][751] ) );
  DFF \zreg_reg[752]  ( .D(o[752]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][752] ) );
  DFF \zreg_reg[753]  ( .D(o[753]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][753] ) );
  DFF \zreg_reg[754]  ( .D(o[754]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][754] ) );
  DFF \zreg_reg[755]  ( .D(o[755]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][755] ) );
  DFF \zreg_reg[756]  ( .D(o[756]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][756] ) );
  DFF \zreg_reg[757]  ( .D(o[757]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][757] ) );
  DFF \zreg_reg[758]  ( .D(o[758]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][758] ) );
  DFF \zreg_reg[759]  ( .D(o[759]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][759] ) );
  DFF \zreg_reg[760]  ( .D(o[760]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][760] ) );
  DFF \zreg_reg[761]  ( .D(o[761]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][761] ) );
  DFF \zreg_reg[762]  ( .D(o[762]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][762] ) );
  DFF \zreg_reg[763]  ( .D(o[763]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][763] ) );
  DFF \zreg_reg[764]  ( .D(o[764]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][764] ) );
  DFF \zreg_reg[765]  ( .D(o[765]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][765] ) );
  DFF \zreg_reg[766]  ( .D(o[766]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][766] ) );
  DFF \zreg_reg[767]  ( .D(o[767]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][767] ) );
  DFF \zreg_reg[768]  ( .D(o[768]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][768] ) );
  DFF \zreg_reg[769]  ( .D(o[769]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][769] ) );
  DFF \zreg_reg[770]  ( .D(o[770]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][770] ) );
  DFF \zreg_reg[771]  ( .D(o[771]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][771] ) );
  DFF \zreg_reg[772]  ( .D(o[772]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][772] ) );
  DFF \zreg_reg[773]  ( .D(o[773]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][773] ) );
  DFF \zreg_reg[774]  ( .D(o[774]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][774] ) );
  DFF \zreg_reg[775]  ( .D(o[775]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][775] ) );
  DFF \zreg_reg[776]  ( .D(o[776]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][776] ) );
  DFF \zreg_reg[777]  ( .D(o[777]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][777] ) );
  DFF \zreg_reg[778]  ( .D(o[778]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][778] ) );
  DFF \zreg_reg[779]  ( .D(o[779]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][779] ) );
  DFF \zreg_reg[780]  ( .D(o[780]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][780] ) );
  DFF \zreg_reg[781]  ( .D(o[781]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][781] ) );
  DFF \zreg_reg[782]  ( .D(o[782]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][782] ) );
  DFF \zreg_reg[783]  ( .D(o[783]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][783] ) );
  DFF \zreg_reg[784]  ( .D(o[784]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][784] ) );
  DFF \zreg_reg[785]  ( .D(o[785]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][785] ) );
  DFF \zreg_reg[786]  ( .D(o[786]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][786] ) );
  DFF \zreg_reg[787]  ( .D(o[787]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][787] ) );
  DFF \zreg_reg[788]  ( .D(o[788]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][788] ) );
  DFF \zreg_reg[789]  ( .D(o[789]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][789] ) );
  DFF \zreg_reg[790]  ( .D(o[790]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][790] ) );
  DFF \zreg_reg[791]  ( .D(o[791]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][791] ) );
  DFF \zreg_reg[792]  ( .D(o[792]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][792] ) );
  DFF \zreg_reg[793]  ( .D(o[793]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][793] ) );
  DFF \zreg_reg[794]  ( .D(o[794]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][794] ) );
  DFF \zreg_reg[795]  ( .D(o[795]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][795] ) );
  DFF \zreg_reg[796]  ( .D(o[796]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][796] ) );
  DFF \zreg_reg[797]  ( .D(o[797]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][797] ) );
  DFF \zreg_reg[798]  ( .D(o[798]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][798] ) );
  DFF \zreg_reg[799]  ( .D(o[799]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][799] ) );
  DFF \zreg_reg[800]  ( .D(o[800]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][800] ) );
  DFF \zreg_reg[801]  ( .D(o[801]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][801] ) );
  DFF \zreg_reg[802]  ( .D(o[802]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][802] ) );
  DFF \zreg_reg[803]  ( .D(o[803]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][803] ) );
  DFF \zreg_reg[804]  ( .D(o[804]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][804] ) );
  DFF \zreg_reg[805]  ( .D(o[805]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][805] ) );
  DFF \zreg_reg[806]  ( .D(o[806]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][806] ) );
  DFF \zreg_reg[807]  ( .D(o[807]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][807] ) );
  DFF \zreg_reg[808]  ( .D(o[808]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][808] ) );
  DFF \zreg_reg[809]  ( .D(o[809]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][809] ) );
  DFF \zreg_reg[810]  ( .D(o[810]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][810] ) );
  DFF \zreg_reg[811]  ( .D(o[811]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][811] ) );
  DFF \zreg_reg[812]  ( .D(o[812]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][812] ) );
  DFF \zreg_reg[813]  ( .D(o[813]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][813] ) );
  DFF \zreg_reg[814]  ( .D(o[814]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][814] ) );
  DFF \zreg_reg[815]  ( .D(o[815]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][815] ) );
  DFF \zreg_reg[816]  ( .D(o[816]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][816] ) );
  DFF \zreg_reg[817]  ( .D(o[817]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][817] ) );
  DFF \zreg_reg[818]  ( .D(o[818]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][818] ) );
  DFF \zreg_reg[819]  ( .D(o[819]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][819] ) );
  DFF \zreg_reg[820]  ( .D(o[820]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][820] ) );
  DFF \zreg_reg[821]  ( .D(o[821]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][821] ) );
  DFF \zreg_reg[822]  ( .D(o[822]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][822] ) );
  DFF \zreg_reg[823]  ( .D(o[823]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][823] ) );
  DFF \zreg_reg[824]  ( .D(o[824]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][824] ) );
  DFF \zreg_reg[825]  ( .D(o[825]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][825] ) );
  DFF \zreg_reg[826]  ( .D(o[826]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][826] ) );
  DFF \zreg_reg[827]  ( .D(o[827]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][827] ) );
  DFF \zreg_reg[828]  ( .D(o[828]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][828] ) );
  DFF \zreg_reg[829]  ( .D(o[829]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][829] ) );
  DFF \zreg_reg[830]  ( .D(o[830]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][830] ) );
  DFF \zreg_reg[831]  ( .D(o[831]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][831] ) );
  DFF \zreg_reg[832]  ( .D(o[832]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][832] ) );
  DFF \zreg_reg[833]  ( .D(o[833]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][833] ) );
  DFF \zreg_reg[834]  ( .D(o[834]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][834] ) );
  DFF \zreg_reg[835]  ( .D(o[835]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][835] ) );
  DFF \zreg_reg[836]  ( .D(o[836]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][836] ) );
  DFF \zreg_reg[837]  ( .D(o[837]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][837] ) );
  DFF \zreg_reg[838]  ( .D(o[838]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][838] ) );
  DFF \zreg_reg[839]  ( .D(o[839]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][839] ) );
  DFF \zreg_reg[840]  ( .D(o[840]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][840] ) );
  DFF \zreg_reg[841]  ( .D(o[841]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][841] ) );
  DFF \zreg_reg[842]  ( .D(o[842]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][842] ) );
  DFF \zreg_reg[843]  ( .D(o[843]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][843] ) );
  DFF \zreg_reg[844]  ( .D(o[844]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][844] ) );
  DFF \zreg_reg[845]  ( .D(o[845]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][845] ) );
  DFF \zreg_reg[846]  ( .D(o[846]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][846] ) );
  DFF \zreg_reg[847]  ( .D(o[847]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][847] ) );
  DFF \zreg_reg[848]  ( .D(o[848]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][848] ) );
  DFF \zreg_reg[849]  ( .D(o[849]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][849] ) );
  DFF \zreg_reg[850]  ( .D(o[850]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][850] ) );
  DFF \zreg_reg[851]  ( .D(o[851]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][851] ) );
  DFF \zreg_reg[852]  ( .D(o[852]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][852] ) );
  DFF \zreg_reg[853]  ( .D(o[853]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][853] ) );
  DFF \zreg_reg[854]  ( .D(o[854]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][854] ) );
  DFF \zreg_reg[855]  ( .D(o[855]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][855] ) );
  DFF \zreg_reg[856]  ( .D(o[856]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][856] ) );
  DFF \zreg_reg[857]  ( .D(o[857]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][857] ) );
  DFF \zreg_reg[858]  ( .D(o[858]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][858] ) );
  DFF \zreg_reg[859]  ( .D(o[859]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][859] ) );
  DFF \zreg_reg[860]  ( .D(o[860]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][860] ) );
  DFF \zreg_reg[861]  ( .D(o[861]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][861] ) );
  DFF \zreg_reg[862]  ( .D(o[862]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][862] ) );
  DFF \zreg_reg[863]  ( .D(o[863]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][863] ) );
  DFF \zreg_reg[864]  ( .D(o[864]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][864] ) );
  DFF \zreg_reg[865]  ( .D(o[865]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][865] ) );
  DFF \zreg_reg[866]  ( .D(o[866]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][866] ) );
  DFF \zreg_reg[867]  ( .D(o[867]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][867] ) );
  DFF \zreg_reg[868]  ( .D(o[868]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][868] ) );
  DFF \zreg_reg[869]  ( .D(o[869]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][869] ) );
  DFF \zreg_reg[870]  ( .D(o[870]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][870] ) );
  DFF \zreg_reg[871]  ( .D(o[871]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][871] ) );
  DFF \zreg_reg[872]  ( .D(o[872]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][872] ) );
  DFF \zreg_reg[873]  ( .D(o[873]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][873] ) );
  DFF \zreg_reg[874]  ( .D(o[874]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][874] ) );
  DFF \zreg_reg[875]  ( .D(o[875]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][875] ) );
  DFF \zreg_reg[876]  ( .D(o[876]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][876] ) );
  DFF \zreg_reg[877]  ( .D(o[877]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][877] ) );
  DFF \zreg_reg[878]  ( .D(o[878]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][878] ) );
  DFF \zreg_reg[879]  ( .D(o[879]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][879] ) );
  DFF \zreg_reg[880]  ( .D(o[880]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][880] ) );
  DFF \zreg_reg[881]  ( .D(o[881]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][881] ) );
  DFF \zreg_reg[882]  ( .D(o[882]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][882] ) );
  DFF \zreg_reg[883]  ( .D(o[883]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][883] ) );
  DFF \zreg_reg[884]  ( .D(o[884]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][884] ) );
  DFF \zreg_reg[885]  ( .D(o[885]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][885] ) );
  DFF \zreg_reg[886]  ( .D(o[886]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][886] ) );
  DFF \zreg_reg[887]  ( .D(o[887]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][887] ) );
  DFF \zreg_reg[888]  ( .D(o[888]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][888] ) );
  DFF \zreg_reg[889]  ( .D(o[889]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][889] ) );
  DFF \zreg_reg[890]  ( .D(o[890]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][890] ) );
  DFF \zreg_reg[891]  ( .D(o[891]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][891] ) );
  DFF \zreg_reg[892]  ( .D(o[892]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][892] ) );
  DFF \zreg_reg[893]  ( .D(o[893]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][893] ) );
  DFF \zreg_reg[894]  ( .D(o[894]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][894] ) );
  DFF \zreg_reg[895]  ( .D(o[895]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][895] ) );
  DFF \zreg_reg[896]  ( .D(o[896]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][896] ) );
  DFF \zreg_reg[897]  ( .D(o[897]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][897] ) );
  DFF \zreg_reg[898]  ( .D(o[898]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][898] ) );
  DFF \zreg_reg[899]  ( .D(o[899]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][899] ) );
  DFF \zreg_reg[900]  ( .D(o[900]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][900] ) );
  DFF \zreg_reg[901]  ( .D(o[901]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][901] ) );
  DFF \zreg_reg[902]  ( .D(o[902]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][902] ) );
  DFF \zreg_reg[903]  ( .D(o[903]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][903] ) );
  DFF \zreg_reg[904]  ( .D(o[904]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][904] ) );
  DFF \zreg_reg[905]  ( .D(o[905]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][905] ) );
  DFF \zreg_reg[906]  ( .D(o[906]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][906] ) );
  DFF \zreg_reg[907]  ( .D(o[907]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][907] ) );
  DFF \zreg_reg[908]  ( .D(o[908]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][908] ) );
  DFF \zreg_reg[909]  ( .D(o[909]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][909] ) );
  DFF \zreg_reg[910]  ( .D(o[910]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][910] ) );
  DFF \zreg_reg[911]  ( .D(o[911]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][911] ) );
  DFF \zreg_reg[912]  ( .D(o[912]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][912] ) );
  DFF \zreg_reg[913]  ( .D(o[913]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][913] ) );
  DFF \zreg_reg[914]  ( .D(o[914]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][914] ) );
  DFF \zreg_reg[915]  ( .D(o[915]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][915] ) );
  DFF \zreg_reg[916]  ( .D(o[916]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][916] ) );
  DFF \zreg_reg[917]  ( .D(o[917]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][917] ) );
  DFF \zreg_reg[918]  ( .D(o[918]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][918] ) );
  DFF \zreg_reg[919]  ( .D(o[919]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][919] ) );
  DFF \zreg_reg[920]  ( .D(o[920]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][920] ) );
  DFF \zreg_reg[921]  ( .D(o[921]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][921] ) );
  DFF \zreg_reg[922]  ( .D(o[922]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][922] ) );
  DFF \zreg_reg[923]  ( .D(o[923]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][923] ) );
  DFF \zreg_reg[924]  ( .D(o[924]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][924] ) );
  DFF \zreg_reg[925]  ( .D(o[925]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][925] ) );
  DFF \zreg_reg[926]  ( .D(o[926]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][926] ) );
  DFF \zreg_reg[927]  ( .D(o[927]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][927] ) );
  DFF \zreg_reg[928]  ( .D(o[928]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][928] ) );
  DFF \zreg_reg[929]  ( .D(o[929]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][929] ) );
  DFF \zreg_reg[930]  ( .D(o[930]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][930] ) );
  DFF \zreg_reg[931]  ( .D(o[931]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][931] ) );
  DFF \zreg_reg[932]  ( .D(o[932]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][932] ) );
  DFF \zreg_reg[933]  ( .D(o[933]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][933] ) );
  DFF \zreg_reg[934]  ( .D(o[934]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][934] ) );
  DFF \zreg_reg[935]  ( .D(o[935]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][935] ) );
  DFF \zreg_reg[936]  ( .D(o[936]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][936] ) );
  DFF \zreg_reg[937]  ( .D(o[937]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][937] ) );
  DFF \zreg_reg[938]  ( .D(o[938]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][938] ) );
  DFF \zreg_reg[939]  ( .D(o[939]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][939] ) );
  DFF \zreg_reg[940]  ( .D(o[940]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][940] ) );
  DFF \zreg_reg[941]  ( .D(o[941]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][941] ) );
  DFF \zreg_reg[942]  ( .D(o[942]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][942] ) );
  DFF \zreg_reg[943]  ( .D(o[943]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][943] ) );
  DFF \zreg_reg[944]  ( .D(o[944]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][944] ) );
  DFF \zreg_reg[945]  ( .D(o[945]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][945] ) );
  DFF \zreg_reg[946]  ( .D(o[946]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][946] ) );
  DFF \zreg_reg[947]  ( .D(o[947]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][947] ) );
  DFF \zreg_reg[948]  ( .D(o[948]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][948] ) );
  DFF \zreg_reg[949]  ( .D(o[949]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][949] ) );
  DFF \zreg_reg[950]  ( .D(o[950]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][950] ) );
  DFF \zreg_reg[951]  ( .D(o[951]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][951] ) );
  DFF \zreg_reg[952]  ( .D(o[952]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][952] ) );
  DFF \zreg_reg[953]  ( .D(o[953]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][953] ) );
  DFF \zreg_reg[954]  ( .D(o[954]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][954] ) );
  DFF \zreg_reg[955]  ( .D(o[955]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][955] ) );
  DFF \zreg_reg[956]  ( .D(o[956]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][956] ) );
  DFF \zreg_reg[957]  ( .D(o[957]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][957] ) );
  DFF \zreg_reg[958]  ( .D(o[958]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][958] ) );
  DFF \zreg_reg[959]  ( .D(o[959]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][959] ) );
  DFF \zreg_reg[960]  ( .D(o[960]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][960] ) );
  DFF \zreg_reg[961]  ( .D(o[961]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][961] ) );
  DFF \zreg_reg[962]  ( .D(o[962]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][962] ) );
  DFF \zreg_reg[963]  ( .D(o[963]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][963] ) );
  DFF \zreg_reg[964]  ( .D(o[964]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][964] ) );
  DFF \zreg_reg[965]  ( .D(o[965]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][965] ) );
  DFF \zreg_reg[966]  ( .D(o[966]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][966] ) );
  DFF \zreg_reg[967]  ( .D(o[967]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][967] ) );
  DFF \zreg_reg[968]  ( .D(o[968]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][968] ) );
  DFF \zreg_reg[969]  ( .D(o[969]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][969] ) );
  DFF \zreg_reg[970]  ( .D(o[970]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][970] ) );
  DFF \zreg_reg[971]  ( .D(o[971]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][971] ) );
  DFF \zreg_reg[972]  ( .D(o[972]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][972] ) );
  DFF \zreg_reg[973]  ( .D(o[973]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][973] ) );
  DFF \zreg_reg[974]  ( .D(o[974]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][974] ) );
  DFF \zreg_reg[975]  ( .D(o[975]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][975] ) );
  DFF \zreg_reg[976]  ( .D(o[976]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][976] ) );
  DFF \zreg_reg[977]  ( .D(o[977]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][977] ) );
  DFF \zreg_reg[978]  ( .D(o[978]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][978] ) );
  DFF \zreg_reg[979]  ( .D(o[979]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][979] ) );
  DFF \zreg_reg[980]  ( .D(o[980]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][980] ) );
  DFF \zreg_reg[981]  ( .D(o[981]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][981] ) );
  DFF \zreg_reg[982]  ( .D(o[982]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][982] ) );
  DFF \zreg_reg[983]  ( .D(o[983]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][983] ) );
  DFF \zreg_reg[984]  ( .D(o[984]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][984] ) );
  DFF \zreg_reg[985]  ( .D(o[985]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][985] ) );
  DFF \zreg_reg[986]  ( .D(o[986]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][986] ) );
  DFF \zreg_reg[987]  ( .D(o[987]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][987] ) );
  DFF \zreg_reg[988]  ( .D(o[988]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][988] ) );
  DFF \zreg_reg[989]  ( .D(o[989]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][989] ) );
  DFF \zreg_reg[990]  ( .D(o[990]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][990] ) );
  DFF \zreg_reg[991]  ( .D(o[991]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][991] ) );
  DFF \zreg_reg[992]  ( .D(o[992]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][992] ) );
  DFF \zreg_reg[993]  ( .D(o[993]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][993] ) );
  DFF \zreg_reg[994]  ( .D(o[994]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][994] ) );
  DFF \zreg_reg[995]  ( .D(o[995]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][995] ) );
  DFF \zreg_reg[996]  ( .D(o[996]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][996] ) );
  DFF \zreg_reg[997]  ( .D(o[997]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][997] ) );
  DFF \zreg_reg[998]  ( .D(o[998]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][998] ) );
  DFF \zreg_reg[999]  ( .D(o[999]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][999] ) );
  DFF \zreg_reg[1000]  ( .D(o[1000]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][1000] ) );
  DFF \zreg_reg[1001]  ( .D(o[1001]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][1001] ) );
  DFF \zreg_reg[1002]  ( .D(o[1002]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][1002] ) );
  DFF \zreg_reg[1003]  ( .D(o[1003]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][1003] ) );
  DFF \zreg_reg[1004]  ( .D(o[1004]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][1004] ) );
  DFF \zreg_reg[1005]  ( .D(o[1005]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][1005] ) );
  DFF \zreg_reg[1006]  ( .D(o[1006]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][1006] ) );
  DFF \zreg_reg[1007]  ( .D(o[1007]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][1007] ) );
  DFF \zreg_reg[1008]  ( .D(o[1008]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][1008] ) );
  DFF \zreg_reg[1009]  ( .D(o[1009]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][1009] ) );
  DFF \zreg_reg[1010]  ( .D(o[1010]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][1010] ) );
  DFF \zreg_reg[1011]  ( .D(o[1011]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][1011] ) );
  DFF \zreg_reg[1012]  ( .D(o[1012]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][1012] ) );
  DFF \zreg_reg[1013]  ( .D(o[1013]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][1013] ) );
  DFF \zreg_reg[1014]  ( .D(o[1014]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][1014] ) );
  DFF \zreg_reg[1015]  ( .D(o[1015]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][1015] ) );
  DFF \zreg_reg[1016]  ( .D(o[1016]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][1016] ) );
  DFF \zreg_reg[1017]  ( .D(o[1017]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][1017] ) );
  DFF \zreg_reg[1018]  ( .D(o[1018]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][1018] ) );
  DFF \zreg_reg[1019]  ( .D(o[1019]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][1019] ) );
  DFF \zreg_reg[1020]  ( .D(o[1020]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][1020] ) );
  DFF \zreg_reg[1021]  ( .D(o[1021]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][1021] ) );
  DFF \zreg_reg[1022]  ( .D(o[1022]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][1022] ) );
  DFF \zreg_reg[1023]  ( .D(o[1023]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][1023] ) );
  DFF \zreg_reg[1024]  ( .D(\zout[0][1024] ), .CLK(clk), .RST(start), .I(1'b0), 
        .Q(\zin[0][1024] ) );
endmodule


module MUX_N1024_1 ( A, B, S, O );
  input [1023:0] A;
  input [1023:0] B;
  output [1023:0] O;
  input S;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048;

  XOR U1 ( .A(A[9]), .B(n1), .Z(O[9]) );
  AND U2 ( .A(S), .B(n2), .Z(n1) );
  XOR U3 ( .A(B[9]), .B(A[9]), .Z(n2) );
  XOR U4 ( .A(A[99]), .B(n3), .Z(O[99]) );
  AND U5 ( .A(S), .B(n4), .Z(n3) );
  XOR U6 ( .A(B[99]), .B(A[99]), .Z(n4) );
  XOR U7 ( .A(A[999]), .B(n5), .Z(O[999]) );
  AND U8 ( .A(S), .B(n6), .Z(n5) );
  XOR U9 ( .A(B[999]), .B(A[999]), .Z(n6) );
  XOR U10 ( .A(A[998]), .B(n7), .Z(O[998]) );
  AND U11 ( .A(S), .B(n8), .Z(n7) );
  XOR U12 ( .A(B[998]), .B(A[998]), .Z(n8) );
  XOR U13 ( .A(A[997]), .B(n9), .Z(O[997]) );
  AND U14 ( .A(S), .B(n10), .Z(n9) );
  XOR U15 ( .A(B[997]), .B(A[997]), .Z(n10) );
  XOR U16 ( .A(A[996]), .B(n11), .Z(O[996]) );
  AND U17 ( .A(S), .B(n12), .Z(n11) );
  XOR U18 ( .A(B[996]), .B(A[996]), .Z(n12) );
  XOR U19 ( .A(A[995]), .B(n13), .Z(O[995]) );
  AND U20 ( .A(S), .B(n14), .Z(n13) );
  XOR U21 ( .A(B[995]), .B(A[995]), .Z(n14) );
  XOR U22 ( .A(A[994]), .B(n15), .Z(O[994]) );
  AND U23 ( .A(S), .B(n16), .Z(n15) );
  XOR U24 ( .A(B[994]), .B(A[994]), .Z(n16) );
  XOR U25 ( .A(A[993]), .B(n17), .Z(O[993]) );
  AND U26 ( .A(S), .B(n18), .Z(n17) );
  XOR U27 ( .A(B[993]), .B(A[993]), .Z(n18) );
  XOR U28 ( .A(A[992]), .B(n19), .Z(O[992]) );
  AND U29 ( .A(S), .B(n20), .Z(n19) );
  XOR U30 ( .A(B[992]), .B(A[992]), .Z(n20) );
  XOR U31 ( .A(A[991]), .B(n21), .Z(O[991]) );
  AND U32 ( .A(S), .B(n22), .Z(n21) );
  XOR U33 ( .A(B[991]), .B(A[991]), .Z(n22) );
  XOR U34 ( .A(A[990]), .B(n23), .Z(O[990]) );
  AND U35 ( .A(S), .B(n24), .Z(n23) );
  XOR U36 ( .A(B[990]), .B(A[990]), .Z(n24) );
  XOR U37 ( .A(A[98]), .B(n25), .Z(O[98]) );
  AND U38 ( .A(S), .B(n26), .Z(n25) );
  XOR U39 ( .A(B[98]), .B(A[98]), .Z(n26) );
  XOR U40 ( .A(A[989]), .B(n27), .Z(O[989]) );
  AND U41 ( .A(S), .B(n28), .Z(n27) );
  XOR U42 ( .A(B[989]), .B(A[989]), .Z(n28) );
  XOR U43 ( .A(A[988]), .B(n29), .Z(O[988]) );
  AND U44 ( .A(S), .B(n30), .Z(n29) );
  XOR U45 ( .A(B[988]), .B(A[988]), .Z(n30) );
  XOR U46 ( .A(A[987]), .B(n31), .Z(O[987]) );
  AND U47 ( .A(S), .B(n32), .Z(n31) );
  XOR U48 ( .A(B[987]), .B(A[987]), .Z(n32) );
  XOR U49 ( .A(A[986]), .B(n33), .Z(O[986]) );
  AND U50 ( .A(S), .B(n34), .Z(n33) );
  XOR U51 ( .A(B[986]), .B(A[986]), .Z(n34) );
  XOR U52 ( .A(A[985]), .B(n35), .Z(O[985]) );
  AND U53 ( .A(S), .B(n36), .Z(n35) );
  XOR U54 ( .A(B[985]), .B(A[985]), .Z(n36) );
  XOR U55 ( .A(A[984]), .B(n37), .Z(O[984]) );
  AND U56 ( .A(S), .B(n38), .Z(n37) );
  XOR U57 ( .A(B[984]), .B(A[984]), .Z(n38) );
  XOR U58 ( .A(A[983]), .B(n39), .Z(O[983]) );
  AND U59 ( .A(S), .B(n40), .Z(n39) );
  XOR U60 ( .A(B[983]), .B(A[983]), .Z(n40) );
  XOR U61 ( .A(A[982]), .B(n41), .Z(O[982]) );
  AND U62 ( .A(S), .B(n42), .Z(n41) );
  XOR U63 ( .A(B[982]), .B(A[982]), .Z(n42) );
  XOR U64 ( .A(A[981]), .B(n43), .Z(O[981]) );
  AND U65 ( .A(S), .B(n44), .Z(n43) );
  XOR U66 ( .A(B[981]), .B(A[981]), .Z(n44) );
  XOR U67 ( .A(A[980]), .B(n45), .Z(O[980]) );
  AND U68 ( .A(S), .B(n46), .Z(n45) );
  XOR U69 ( .A(B[980]), .B(A[980]), .Z(n46) );
  XOR U70 ( .A(A[97]), .B(n47), .Z(O[97]) );
  AND U71 ( .A(S), .B(n48), .Z(n47) );
  XOR U72 ( .A(B[97]), .B(A[97]), .Z(n48) );
  XOR U73 ( .A(A[979]), .B(n49), .Z(O[979]) );
  AND U74 ( .A(S), .B(n50), .Z(n49) );
  XOR U75 ( .A(B[979]), .B(A[979]), .Z(n50) );
  XOR U76 ( .A(A[978]), .B(n51), .Z(O[978]) );
  AND U77 ( .A(S), .B(n52), .Z(n51) );
  XOR U78 ( .A(B[978]), .B(A[978]), .Z(n52) );
  XOR U79 ( .A(A[977]), .B(n53), .Z(O[977]) );
  AND U80 ( .A(S), .B(n54), .Z(n53) );
  XOR U81 ( .A(B[977]), .B(A[977]), .Z(n54) );
  XOR U82 ( .A(A[976]), .B(n55), .Z(O[976]) );
  AND U83 ( .A(S), .B(n56), .Z(n55) );
  XOR U84 ( .A(B[976]), .B(A[976]), .Z(n56) );
  XOR U85 ( .A(A[975]), .B(n57), .Z(O[975]) );
  AND U86 ( .A(S), .B(n58), .Z(n57) );
  XOR U87 ( .A(B[975]), .B(A[975]), .Z(n58) );
  XOR U88 ( .A(A[974]), .B(n59), .Z(O[974]) );
  AND U89 ( .A(S), .B(n60), .Z(n59) );
  XOR U90 ( .A(B[974]), .B(A[974]), .Z(n60) );
  XOR U91 ( .A(A[973]), .B(n61), .Z(O[973]) );
  AND U92 ( .A(S), .B(n62), .Z(n61) );
  XOR U93 ( .A(B[973]), .B(A[973]), .Z(n62) );
  XOR U94 ( .A(A[972]), .B(n63), .Z(O[972]) );
  AND U95 ( .A(S), .B(n64), .Z(n63) );
  XOR U96 ( .A(B[972]), .B(A[972]), .Z(n64) );
  XOR U97 ( .A(A[971]), .B(n65), .Z(O[971]) );
  AND U98 ( .A(S), .B(n66), .Z(n65) );
  XOR U99 ( .A(B[971]), .B(A[971]), .Z(n66) );
  XOR U100 ( .A(A[970]), .B(n67), .Z(O[970]) );
  AND U101 ( .A(S), .B(n68), .Z(n67) );
  XOR U102 ( .A(B[970]), .B(A[970]), .Z(n68) );
  XOR U103 ( .A(A[96]), .B(n69), .Z(O[96]) );
  AND U104 ( .A(S), .B(n70), .Z(n69) );
  XOR U105 ( .A(B[96]), .B(A[96]), .Z(n70) );
  XOR U106 ( .A(A[969]), .B(n71), .Z(O[969]) );
  AND U107 ( .A(S), .B(n72), .Z(n71) );
  XOR U108 ( .A(B[969]), .B(A[969]), .Z(n72) );
  XOR U109 ( .A(A[968]), .B(n73), .Z(O[968]) );
  AND U110 ( .A(S), .B(n74), .Z(n73) );
  XOR U111 ( .A(B[968]), .B(A[968]), .Z(n74) );
  XOR U112 ( .A(A[967]), .B(n75), .Z(O[967]) );
  AND U113 ( .A(S), .B(n76), .Z(n75) );
  XOR U114 ( .A(B[967]), .B(A[967]), .Z(n76) );
  XOR U115 ( .A(A[966]), .B(n77), .Z(O[966]) );
  AND U116 ( .A(S), .B(n78), .Z(n77) );
  XOR U117 ( .A(B[966]), .B(A[966]), .Z(n78) );
  XOR U118 ( .A(A[965]), .B(n79), .Z(O[965]) );
  AND U119 ( .A(S), .B(n80), .Z(n79) );
  XOR U120 ( .A(B[965]), .B(A[965]), .Z(n80) );
  XOR U121 ( .A(A[964]), .B(n81), .Z(O[964]) );
  AND U122 ( .A(S), .B(n82), .Z(n81) );
  XOR U123 ( .A(B[964]), .B(A[964]), .Z(n82) );
  XOR U124 ( .A(A[963]), .B(n83), .Z(O[963]) );
  AND U125 ( .A(S), .B(n84), .Z(n83) );
  XOR U126 ( .A(B[963]), .B(A[963]), .Z(n84) );
  XOR U127 ( .A(A[962]), .B(n85), .Z(O[962]) );
  AND U128 ( .A(S), .B(n86), .Z(n85) );
  XOR U129 ( .A(B[962]), .B(A[962]), .Z(n86) );
  XOR U130 ( .A(A[961]), .B(n87), .Z(O[961]) );
  AND U131 ( .A(S), .B(n88), .Z(n87) );
  XOR U132 ( .A(B[961]), .B(A[961]), .Z(n88) );
  XOR U133 ( .A(A[960]), .B(n89), .Z(O[960]) );
  AND U134 ( .A(S), .B(n90), .Z(n89) );
  XOR U135 ( .A(B[960]), .B(A[960]), .Z(n90) );
  XOR U136 ( .A(A[95]), .B(n91), .Z(O[95]) );
  AND U137 ( .A(S), .B(n92), .Z(n91) );
  XOR U138 ( .A(B[95]), .B(A[95]), .Z(n92) );
  XOR U139 ( .A(A[959]), .B(n93), .Z(O[959]) );
  AND U140 ( .A(S), .B(n94), .Z(n93) );
  XOR U141 ( .A(B[959]), .B(A[959]), .Z(n94) );
  XOR U142 ( .A(A[958]), .B(n95), .Z(O[958]) );
  AND U143 ( .A(S), .B(n96), .Z(n95) );
  XOR U144 ( .A(B[958]), .B(A[958]), .Z(n96) );
  XOR U145 ( .A(A[957]), .B(n97), .Z(O[957]) );
  AND U146 ( .A(S), .B(n98), .Z(n97) );
  XOR U147 ( .A(B[957]), .B(A[957]), .Z(n98) );
  XOR U148 ( .A(A[956]), .B(n99), .Z(O[956]) );
  AND U149 ( .A(S), .B(n100), .Z(n99) );
  XOR U150 ( .A(B[956]), .B(A[956]), .Z(n100) );
  XOR U151 ( .A(A[955]), .B(n101), .Z(O[955]) );
  AND U152 ( .A(S), .B(n102), .Z(n101) );
  XOR U153 ( .A(B[955]), .B(A[955]), .Z(n102) );
  XOR U154 ( .A(A[954]), .B(n103), .Z(O[954]) );
  AND U155 ( .A(S), .B(n104), .Z(n103) );
  XOR U156 ( .A(B[954]), .B(A[954]), .Z(n104) );
  XOR U157 ( .A(A[953]), .B(n105), .Z(O[953]) );
  AND U158 ( .A(S), .B(n106), .Z(n105) );
  XOR U159 ( .A(B[953]), .B(A[953]), .Z(n106) );
  XOR U160 ( .A(A[952]), .B(n107), .Z(O[952]) );
  AND U161 ( .A(S), .B(n108), .Z(n107) );
  XOR U162 ( .A(B[952]), .B(A[952]), .Z(n108) );
  XOR U163 ( .A(A[951]), .B(n109), .Z(O[951]) );
  AND U164 ( .A(S), .B(n110), .Z(n109) );
  XOR U165 ( .A(B[951]), .B(A[951]), .Z(n110) );
  XOR U166 ( .A(A[950]), .B(n111), .Z(O[950]) );
  AND U167 ( .A(S), .B(n112), .Z(n111) );
  XOR U168 ( .A(B[950]), .B(A[950]), .Z(n112) );
  XOR U169 ( .A(A[94]), .B(n113), .Z(O[94]) );
  AND U170 ( .A(S), .B(n114), .Z(n113) );
  XOR U171 ( .A(B[94]), .B(A[94]), .Z(n114) );
  XOR U172 ( .A(A[949]), .B(n115), .Z(O[949]) );
  AND U173 ( .A(S), .B(n116), .Z(n115) );
  XOR U174 ( .A(B[949]), .B(A[949]), .Z(n116) );
  XOR U175 ( .A(A[948]), .B(n117), .Z(O[948]) );
  AND U176 ( .A(S), .B(n118), .Z(n117) );
  XOR U177 ( .A(B[948]), .B(A[948]), .Z(n118) );
  XOR U178 ( .A(A[947]), .B(n119), .Z(O[947]) );
  AND U179 ( .A(S), .B(n120), .Z(n119) );
  XOR U180 ( .A(B[947]), .B(A[947]), .Z(n120) );
  XOR U181 ( .A(A[946]), .B(n121), .Z(O[946]) );
  AND U182 ( .A(S), .B(n122), .Z(n121) );
  XOR U183 ( .A(B[946]), .B(A[946]), .Z(n122) );
  XOR U184 ( .A(A[945]), .B(n123), .Z(O[945]) );
  AND U185 ( .A(S), .B(n124), .Z(n123) );
  XOR U186 ( .A(B[945]), .B(A[945]), .Z(n124) );
  XOR U187 ( .A(A[944]), .B(n125), .Z(O[944]) );
  AND U188 ( .A(S), .B(n126), .Z(n125) );
  XOR U189 ( .A(B[944]), .B(A[944]), .Z(n126) );
  XOR U190 ( .A(A[943]), .B(n127), .Z(O[943]) );
  AND U191 ( .A(S), .B(n128), .Z(n127) );
  XOR U192 ( .A(B[943]), .B(A[943]), .Z(n128) );
  XOR U193 ( .A(A[942]), .B(n129), .Z(O[942]) );
  AND U194 ( .A(S), .B(n130), .Z(n129) );
  XOR U195 ( .A(B[942]), .B(A[942]), .Z(n130) );
  XOR U196 ( .A(A[941]), .B(n131), .Z(O[941]) );
  AND U197 ( .A(S), .B(n132), .Z(n131) );
  XOR U198 ( .A(B[941]), .B(A[941]), .Z(n132) );
  XOR U199 ( .A(A[940]), .B(n133), .Z(O[940]) );
  AND U200 ( .A(S), .B(n134), .Z(n133) );
  XOR U201 ( .A(B[940]), .B(A[940]), .Z(n134) );
  XOR U202 ( .A(A[93]), .B(n135), .Z(O[93]) );
  AND U203 ( .A(S), .B(n136), .Z(n135) );
  XOR U204 ( .A(B[93]), .B(A[93]), .Z(n136) );
  XOR U205 ( .A(A[939]), .B(n137), .Z(O[939]) );
  AND U206 ( .A(S), .B(n138), .Z(n137) );
  XOR U207 ( .A(B[939]), .B(A[939]), .Z(n138) );
  XOR U208 ( .A(A[938]), .B(n139), .Z(O[938]) );
  AND U209 ( .A(S), .B(n140), .Z(n139) );
  XOR U210 ( .A(B[938]), .B(A[938]), .Z(n140) );
  XOR U211 ( .A(A[937]), .B(n141), .Z(O[937]) );
  AND U212 ( .A(S), .B(n142), .Z(n141) );
  XOR U213 ( .A(B[937]), .B(A[937]), .Z(n142) );
  XOR U214 ( .A(A[936]), .B(n143), .Z(O[936]) );
  AND U215 ( .A(S), .B(n144), .Z(n143) );
  XOR U216 ( .A(B[936]), .B(A[936]), .Z(n144) );
  XOR U217 ( .A(A[935]), .B(n145), .Z(O[935]) );
  AND U218 ( .A(S), .B(n146), .Z(n145) );
  XOR U219 ( .A(B[935]), .B(A[935]), .Z(n146) );
  XOR U220 ( .A(A[934]), .B(n147), .Z(O[934]) );
  AND U221 ( .A(S), .B(n148), .Z(n147) );
  XOR U222 ( .A(B[934]), .B(A[934]), .Z(n148) );
  XOR U223 ( .A(A[933]), .B(n149), .Z(O[933]) );
  AND U224 ( .A(S), .B(n150), .Z(n149) );
  XOR U225 ( .A(B[933]), .B(A[933]), .Z(n150) );
  XOR U226 ( .A(A[932]), .B(n151), .Z(O[932]) );
  AND U227 ( .A(S), .B(n152), .Z(n151) );
  XOR U228 ( .A(B[932]), .B(A[932]), .Z(n152) );
  XOR U229 ( .A(A[931]), .B(n153), .Z(O[931]) );
  AND U230 ( .A(S), .B(n154), .Z(n153) );
  XOR U231 ( .A(B[931]), .B(A[931]), .Z(n154) );
  XOR U232 ( .A(A[930]), .B(n155), .Z(O[930]) );
  AND U233 ( .A(S), .B(n156), .Z(n155) );
  XOR U234 ( .A(B[930]), .B(A[930]), .Z(n156) );
  XOR U235 ( .A(A[92]), .B(n157), .Z(O[92]) );
  AND U236 ( .A(S), .B(n158), .Z(n157) );
  XOR U237 ( .A(B[92]), .B(A[92]), .Z(n158) );
  XOR U238 ( .A(A[929]), .B(n159), .Z(O[929]) );
  AND U239 ( .A(S), .B(n160), .Z(n159) );
  XOR U240 ( .A(B[929]), .B(A[929]), .Z(n160) );
  XOR U241 ( .A(A[928]), .B(n161), .Z(O[928]) );
  AND U242 ( .A(S), .B(n162), .Z(n161) );
  XOR U243 ( .A(B[928]), .B(A[928]), .Z(n162) );
  XOR U244 ( .A(A[927]), .B(n163), .Z(O[927]) );
  AND U245 ( .A(S), .B(n164), .Z(n163) );
  XOR U246 ( .A(B[927]), .B(A[927]), .Z(n164) );
  XOR U247 ( .A(A[926]), .B(n165), .Z(O[926]) );
  AND U248 ( .A(S), .B(n166), .Z(n165) );
  XOR U249 ( .A(B[926]), .B(A[926]), .Z(n166) );
  XOR U250 ( .A(A[925]), .B(n167), .Z(O[925]) );
  AND U251 ( .A(S), .B(n168), .Z(n167) );
  XOR U252 ( .A(B[925]), .B(A[925]), .Z(n168) );
  XOR U253 ( .A(A[924]), .B(n169), .Z(O[924]) );
  AND U254 ( .A(S), .B(n170), .Z(n169) );
  XOR U255 ( .A(B[924]), .B(A[924]), .Z(n170) );
  XOR U256 ( .A(A[923]), .B(n171), .Z(O[923]) );
  AND U257 ( .A(S), .B(n172), .Z(n171) );
  XOR U258 ( .A(B[923]), .B(A[923]), .Z(n172) );
  XOR U259 ( .A(A[922]), .B(n173), .Z(O[922]) );
  AND U260 ( .A(S), .B(n174), .Z(n173) );
  XOR U261 ( .A(B[922]), .B(A[922]), .Z(n174) );
  XOR U262 ( .A(A[921]), .B(n175), .Z(O[921]) );
  AND U263 ( .A(S), .B(n176), .Z(n175) );
  XOR U264 ( .A(B[921]), .B(A[921]), .Z(n176) );
  XOR U265 ( .A(A[920]), .B(n177), .Z(O[920]) );
  AND U266 ( .A(S), .B(n178), .Z(n177) );
  XOR U267 ( .A(B[920]), .B(A[920]), .Z(n178) );
  XOR U268 ( .A(A[91]), .B(n179), .Z(O[91]) );
  AND U269 ( .A(S), .B(n180), .Z(n179) );
  XOR U270 ( .A(B[91]), .B(A[91]), .Z(n180) );
  XOR U271 ( .A(A[919]), .B(n181), .Z(O[919]) );
  AND U272 ( .A(S), .B(n182), .Z(n181) );
  XOR U273 ( .A(B[919]), .B(A[919]), .Z(n182) );
  XOR U274 ( .A(A[918]), .B(n183), .Z(O[918]) );
  AND U275 ( .A(S), .B(n184), .Z(n183) );
  XOR U276 ( .A(B[918]), .B(A[918]), .Z(n184) );
  XOR U277 ( .A(A[917]), .B(n185), .Z(O[917]) );
  AND U278 ( .A(S), .B(n186), .Z(n185) );
  XOR U279 ( .A(B[917]), .B(A[917]), .Z(n186) );
  XOR U280 ( .A(A[916]), .B(n187), .Z(O[916]) );
  AND U281 ( .A(S), .B(n188), .Z(n187) );
  XOR U282 ( .A(B[916]), .B(A[916]), .Z(n188) );
  XOR U283 ( .A(A[915]), .B(n189), .Z(O[915]) );
  AND U284 ( .A(S), .B(n190), .Z(n189) );
  XOR U285 ( .A(B[915]), .B(A[915]), .Z(n190) );
  XOR U286 ( .A(A[914]), .B(n191), .Z(O[914]) );
  AND U287 ( .A(S), .B(n192), .Z(n191) );
  XOR U288 ( .A(B[914]), .B(A[914]), .Z(n192) );
  XOR U289 ( .A(A[913]), .B(n193), .Z(O[913]) );
  AND U290 ( .A(S), .B(n194), .Z(n193) );
  XOR U291 ( .A(B[913]), .B(A[913]), .Z(n194) );
  XOR U292 ( .A(A[912]), .B(n195), .Z(O[912]) );
  AND U293 ( .A(S), .B(n196), .Z(n195) );
  XOR U294 ( .A(B[912]), .B(A[912]), .Z(n196) );
  XOR U295 ( .A(A[911]), .B(n197), .Z(O[911]) );
  AND U296 ( .A(S), .B(n198), .Z(n197) );
  XOR U297 ( .A(B[911]), .B(A[911]), .Z(n198) );
  XOR U298 ( .A(A[910]), .B(n199), .Z(O[910]) );
  AND U299 ( .A(S), .B(n200), .Z(n199) );
  XOR U300 ( .A(B[910]), .B(A[910]), .Z(n200) );
  XOR U301 ( .A(A[90]), .B(n201), .Z(O[90]) );
  AND U302 ( .A(S), .B(n202), .Z(n201) );
  XOR U303 ( .A(B[90]), .B(A[90]), .Z(n202) );
  XOR U304 ( .A(A[909]), .B(n203), .Z(O[909]) );
  AND U305 ( .A(S), .B(n204), .Z(n203) );
  XOR U306 ( .A(B[909]), .B(A[909]), .Z(n204) );
  XOR U307 ( .A(A[908]), .B(n205), .Z(O[908]) );
  AND U308 ( .A(S), .B(n206), .Z(n205) );
  XOR U309 ( .A(B[908]), .B(A[908]), .Z(n206) );
  XOR U310 ( .A(A[907]), .B(n207), .Z(O[907]) );
  AND U311 ( .A(S), .B(n208), .Z(n207) );
  XOR U312 ( .A(B[907]), .B(A[907]), .Z(n208) );
  XOR U313 ( .A(A[906]), .B(n209), .Z(O[906]) );
  AND U314 ( .A(S), .B(n210), .Z(n209) );
  XOR U315 ( .A(B[906]), .B(A[906]), .Z(n210) );
  XOR U316 ( .A(A[905]), .B(n211), .Z(O[905]) );
  AND U317 ( .A(S), .B(n212), .Z(n211) );
  XOR U318 ( .A(B[905]), .B(A[905]), .Z(n212) );
  XOR U319 ( .A(A[904]), .B(n213), .Z(O[904]) );
  AND U320 ( .A(S), .B(n214), .Z(n213) );
  XOR U321 ( .A(B[904]), .B(A[904]), .Z(n214) );
  XOR U322 ( .A(A[903]), .B(n215), .Z(O[903]) );
  AND U323 ( .A(S), .B(n216), .Z(n215) );
  XOR U324 ( .A(B[903]), .B(A[903]), .Z(n216) );
  XOR U325 ( .A(A[902]), .B(n217), .Z(O[902]) );
  AND U326 ( .A(S), .B(n218), .Z(n217) );
  XOR U327 ( .A(B[902]), .B(A[902]), .Z(n218) );
  XOR U328 ( .A(A[901]), .B(n219), .Z(O[901]) );
  AND U329 ( .A(S), .B(n220), .Z(n219) );
  XOR U330 ( .A(B[901]), .B(A[901]), .Z(n220) );
  XOR U331 ( .A(A[900]), .B(n221), .Z(O[900]) );
  AND U332 ( .A(S), .B(n222), .Z(n221) );
  XOR U333 ( .A(B[900]), .B(A[900]), .Z(n222) );
  XOR U334 ( .A(A[8]), .B(n223), .Z(O[8]) );
  AND U335 ( .A(S), .B(n224), .Z(n223) );
  XOR U336 ( .A(B[8]), .B(A[8]), .Z(n224) );
  XOR U337 ( .A(A[89]), .B(n225), .Z(O[89]) );
  AND U338 ( .A(S), .B(n226), .Z(n225) );
  XOR U339 ( .A(B[89]), .B(A[89]), .Z(n226) );
  XOR U340 ( .A(A[899]), .B(n227), .Z(O[899]) );
  AND U341 ( .A(S), .B(n228), .Z(n227) );
  XOR U342 ( .A(B[899]), .B(A[899]), .Z(n228) );
  XOR U343 ( .A(A[898]), .B(n229), .Z(O[898]) );
  AND U344 ( .A(S), .B(n230), .Z(n229) );
  XOR U345 ( .A(B[898]), .B(A[898]), .Z(n230) );
  XOR U346 ( .A(A[897]), .B(n231), .Z(O[897]) );
  AND U347 ( .A(S), .B(n232), .Z(n231) );
  XOR U348 ( .A(B[897]), .B(A[897]), .Z(n232) );
  XOR U349 ( .A(A[896]), .B(n233), .Z(O[896]) );
  AND U350 ( .A(S), .B(n234), .Z(n233) );
  XOR U351 ( .A(B[896]), .B(A[896]), .Z(n234) );
  XOR U352 ( .A(A[895]), .B(n235), .Z(O[895]) );
  AND U353 ( .A(S), .B(n236), .Z(n235) );
  XOR U354 ( .A(B[895]), .B(A[895]), .Z(n236) );
  XOR U355 ( .A(A[894]), .B(n237), .Z(O[894]) );
  AND U356 ( .A(S), .B(n238), .Z(n237) );
  XOR U357 ( .A(B[894]), .B(A[894]), .Z(n238) );
  XOR U358 ( .A(A[893]), .B(n239), .Z(O[893]) );
  AND U359 ( .A(S), .B(n240), .Z(n239) );
  XOR U360 ( .A(B[893]), .B(A[893]), .Z(n240) );
  XOR U361 ( .A(A[892]), .B(n241), .Z(O[892]) );
  AND U362 ( .A(S), .B(n242), .Z(n241) );
  XOR U363 ( .A(B[892]), .B(A[892]), .Z(n242) );
  XOR U364 ( .A(A[891]), .B(n243), .Z(O[891]) );
  AND U365 ( .A(S), .B(n244), .Z(n243) );
  XOR U366 ( .A(B[891]), .B(A[891]), .Z(n244) );
  XOR U367 ( .A(A[890]), .B(n245), .Z(O[890]) );
  AND U368 ( .A(S), .B(n246), .Z(n245) );
  XOR U369 ( .A(B[890]), .B(A[890]), .Z(n246) );
  XOR U370 ( .A(A[88]), .B(n247), .Z(O[88]) );
  AND U371 ( .A(S), .B(n248), .Z(n247) );
  XOR U372 ( .A(B[88]), .B(A[88]), .Z(n248) );
  XOR U373 ( .A(A[889]), .B(n249), .Z(O[889]) );
  AND U374 ( .A(S), .B(n250), .Z(n249) );
  XOR U375 ( .A(B[889]), .B(A[889]), .Z(n250) );
  XOR U376 ( .A(A[888]), .B(n251), .Z(O[888]) );
  AND U377 ( .A(S), .B(n252), .Z(n251) );
  XOR U378 ( .A(B[888]), .B(A[888]), .Z(n252) );
  XOR U379 ( .A(A[887]), .B(n253), .Z(O[887]) );
  AND U380 ( .A(S), .B(n254), .Z(n253) );
  XOR U381 ( .A(B[887]), .B(A[887]), .Z(n254) );
  XOR U382 ( .A(A[886]), .B(n255), .Z(O[886]) );
  AND U383 ( .A(S), .B(n256), .Z(n255) );
  XOR U384 ( .A(B[886]), .B(A[886]), .Z(n256) );
  XOR U385 ( .A(A[885]), .B(n257), .Z(O[885]) );
  AND U386 ( .A(S), .B(n258), .Z(n257) );
  XOR U387 ( .A(B[885]), .B(A[885]), .Z(n258) );
  XOR U388 ( .A(A[884]), .B(n259), .Z(O[884]) );
  AND U389 ( .A(S), .B(n260), .Z(n259) );
  XOR U390 ( .A(B[884]), .B(A[884]), .Z(n260) );
  XOR U391 ( .A(A[883]), .B(n261), .Z(O[883]) );
  AND U392 ( .A(S), .B(n262), .Z(n261) );
  XOR U393 ( .A(B[883]), .B(A[883]), .Z(n262) );
  XOR U394 ( .A(A[882]), .B(n263), .Z(O[882]) );
  AND U395 ( .A(S), .B(n264), .Z(n263) );
  XOR U396 ( .A(B[882]), .B(A[882]), .Z(n264) );
  XOR U397 ( .A(A[881]), .B(n265), .Z(O[881]) );
  AND U398 ( .A(S), .B(n266), .Z(n265) );
  XOR U399 ( .A(B[881]), .B(A[881]), .Z(n266) );
  XOR U400 ( .A(A[880]), .B(n267), .Z(O[880]) );
  AND U401 ( .A(S), .B(n268), .Z(n267) );
  XOR U402 ( .A(B[880]), .B(A[880]), .Z(n268) );
  XOR U403 ( .A(A[87]), .B(n269), .Z(O[87]) );
  AND U404 ( .A(S), .B(n270), .Z(n269) );
  XOR U405 ( .A(B[87]), .B(A[87]), .Z(n270) );
  XOR U406 ( .A(A[879]), .B(n271), .Z(O[879]) );
  AND U407 ( .A(S), .B(n272), .Z(n271) );
  XOR U408 ( .A(B[879]), .B(A[879]), .Z(n272) );
  XOR U409 ( .A(A[878]), .B(n273), .Z(O[878]) );
  AND U410 ( .A(S), .B(n274), .Z(n273) );
  XOR U411 ( .A(B[878]), .B(A[878]), .Z(n274) );
  XOR U412 ( .A(A[877]), .B(n275), .Z(O[877]) );
  AND U413 ( .A(S), .B(n276), .Z(n275) );
  XOR U414 ( .A(B[877]), .B(A[877]), .Z(n276) );
  XOR U415 ( .A(A[876]), .B(n277), .Z(O[876]) );
  AND U416 ( .A(S), .B(n278), .Z(n277) );
  XOR U417 ( .A(B[876]), .B(A[876]), .Z(n278) );
  XOR U418 ( .A(A[875]), .B(n279), .Z(O[875]) );
  AND U419 ( .A(S), .B(n280), .Z(n279) );
  XOR U420 ( .A(B[875]), .B(A[875]), .Z(n280) );
  XOR U421 ( .A(A[874]), .B(n281), .Z(O[874]) );
  AND U422 ( .A(S), .B(n282), .Z(n281) );
  XOR U423 ( .A(B[874]), .B(A[874]), .Z(n282) );
  XOR U424 ( .A(A[873]), .B(n283), .Z(O[873]) );
  AND U425 ( .A(S), .B(n284), .Z(n283) );
  XOR U426 ( .A(B[873]), .B(A[873]), .Z(n284) );
  XOR U427 ( .A(A[872]), .B(n285), .Z(O[872]) );
  AND U428 ( .A(S), .B(n286), .Z(n285) );
  XOR U429 ( .A(B[872]), .B(A[872]), .Z(n286) );
  XOR U430 ( .A(A[871]), .B(n287), .Z(O[871]) );
  AND U431 ( .A(S), .B(n288), .Z(n287) );
  XOR U432 ( .A(B[871]), .B(A[871]), .Z(n288) );
  XOR U433 ( .A(A[870]), .B(n289), .Z(O[870]) );
  AND U434 ( .A(S), .B(n290), .Z(n289) );
  XOR U435 ( .A(B[870]), .B(A[870]), .Z(n290) );
  XOR U436 ( .A(A[86]), .B(n291), .Z(O[86]) );
  AND U437 ( .A(S), .B(n292), .Z(n291) );
  XOR U438 ( .A(B[86]), .B(A[86]), .Z(n292) );
  XOR U439 ( .A(A[869]), .B(n293), .Z(O[869]) );
  AND U440 ( .A(S), .B(n294), .Z(n293) );
  XOR U441 ( .A(B[869]), .B(A[869]), .Z(n294) );
  XOR U442 ( .A(A[868]), .B(n295), .Z(O[868]) );
  AND U443 ( .A(S), .B(n296), .Z(n295) );
  XOR U444 ( .A(B[868]), .B(A[868]), .Z(n296) );
  XOR U445 ( .A(A[867]), .B(n297), .Z(O[867]) );
  AND U446 ( .A(S), .B(n298), .Z(n297) );
  XOR U447 ( .A(B[867]), .B(A[867]), .Z(n298) );
  XOR U448 ( .A(A[866]), .B(n299), .Z(O[866]) );
  AND U449 ( .A(S), .B(n300), .Z(n299) );
  XOR U450 ( .A(B[866]), .B(A[866]), .Z(n300) );
  XOR U451 ( .A(A[865]), .B(n301), .Z(O[865]) );
  AND U452 ( .A(S), .B(n302), .Z(n301) );
  XOR U453 ( .A(B[865]), .B(A[865]), .Z(n302) );
  XOR U454 ( .A(A[864]), .B(n303), .Z(O[864]) );
  AND U455 ( .A(S), .B(n304), .Z(n303) );
  XOR U456 ( .A(B[864]), .B(A[864]), .Z(n304) );
  XOR U457 ( .A(A[863]), .B(n305), .Z(O[863]) );
  AND U458 ( .A(S), .B(n306), .Z(n305) );
  XOR U459 ( .A(B[863]), .B(A[863]), .Z(n306) );
  XOR U460 ( .A(A[862]), .B(n307), .Z(O[862]) );
  AND U461 ( .A(S), .B(n308), .Z(n307) );
  XOR U462 ( .A(B[862]), .B(A[862]), .Z(n308) );
  XOR U463 ( .A(A[861]), .B(n309), .Z(O[861]) );
  AND U464 ( .A(S), .B(n310), .Z(n309) );
  XOR U465 ( .A(B[861]), .B(A[861]), .Z(n310) );
  XOR U466 ( .A(A[860]), .B(n311), .Z(O[860]) );
  AND U467 ( .A(S), .B(n312), .Z(n311) );
  XOR U468 ( .A(B[860]), .B(A[860]), .Z(n312) );
  XOR U469 ( .A(A[85]), .B(n313), .Z(O[85]) );
  AND U470 ( .A(S), .B(n314), .Z(n313) );
  XOR U471 ( .A(B[85]), .B(A[85]), .Z(n314) );
  XOR U472 ( .A(A[859]), .B(n315), .Z(O[859]) );
  AND U473 ( .A(S), .B(n316), .Z(n315) );
  XOR U474 ( .A(B[859]), .B(A[859]), .Z(n316) );
  XOR U475 ( .A(A[858]), .B(n317), .Z(O[858]) );
  AND U476 ( .A(S), .B(n318), .Z(n317) );
  XOR U477 ( .A(B[858]), .B(A[858]), .Z(n318) );
  XOR U478 ( .A(A[857]), .B(n319), .Z(O[857]) );
  AND U479 ( .A(S), .B(n320), .Z(n319) );
  XOR U480 ( .A(B[857]), .B(A[857]), .Z(n320) );
  XOR U481 ( .A(A[856]), .B(n321), .Z(O[856]) );
  AND U482 ( .A(S), .B(n322), .Z(n321) );
  XOR U483 ( .A(B[856]), .B(A[856]), .Z(n322) );
  XOR U484 ( .A(A[855]), .B(n323), .Z(O[855]) );
  AND U485 ( .A(S), .B(n324), .Z(n323) );
  XOR U486 ( .A(B[855]), .B(A[855]), .Z(n324) );
  XOR U487 ( .A(A[854]), .B(n325), .Z(O[854]) );
  AND U488 ( .A(S), .B(n326), .Z(n325) );
  XOR U489 ( .A(B[854]), .B(A[854]), .Z(n326) );
  XOR U490 ( .A(A[853]), .B(n327), .Z(O[853]) );
  AND U491 ( .A(S), .B(n328), .Z(n327) );
  XOR U492 ( .A(B[853]), .B(A[853]), .Z(n328) );
  XOR U493 ( .A(A[852]), .B(n329), .Z(O[852]) );
  AND U494 ( .A(S), .B(n330), .Z(n329) );
  XOR U495 ( .A(B[852]), .B(A[852]), .Z(n330) );
  XOR U496 ( .A(A[851]), .B(n331), .Z(O[851]) );
  AND U497 ( .A(S), .B(n332), .Z(n331) );
  XOR U498 ( .A(B[851]), .B(A[851]), .Z(n332) );
  XOR U499 ( .A(A[850]), .B(n333), .Z(O[850]) );
  AND U500 ( .A(S), .B(n334), .Z(n333) );
  XOR U501 ( .A(B[850]), .B(A[850]), .Z(n334) );
  XOR U502 ( .A(A[84]), .B(n335), .Z(O[84]) );
  AND U503 ( .A(S), .B(n336), .Z(n335) );
  XOR U504 ( .A(B[84]), .B(A[84]), .Z(n336) );
  XOR U505 ( .A(A[849]), .B(n337), .Z(O[849]) );
  AND U506 ( .A(S), .B(n338), .Z(n337) );
  XOR U507 ( .A(B[849]), .B(A[849]), .Z(n338) );
  XOR U508 ( .A(A[848]), .B(n339), .Z(O[848]) );
  AND U509 ( .A(S), .B(n340), .Z(n339) );
  XOR U510 ( .A(B[848]), .B(A[848]), .Z(n340) );
  XOR U511 ( .A(A[847]), .B(n341), .Z(O[847]) );
  AND U512 ( .A(S), .B(n342), .Z(n341) );
  XOR U513 ( .A(B[847]), .B(A[847]), .Z(n342) );
  XOR U514 ( .A(A[846]), .B(n343), .Z(O[846]) );
  AND U515 ( .A(S), .B(n344), .Z(n343) );
  XOR U516 ( .A(B[846]), .B(A[846]), .Z(n344) );
  XOR U517 ( .A(A[845]), .B(n345), .Z(O[845]) );
  AND U518 ( .A(S), .B(n346), .Z(n345) );
  XOR U519 ( .A(B[845]), .B(A[845]), .Z(n346) );
  XOR U520 ( .A(A[844]), .B(n347), .Z(O[844]) );
  AND U521 ( .A(S), .B(n348), .Z(n347) );
  XOR U522 ( .A(B[844]), .B(A[844]), .Z(n348) );
  XOR U523 ( .A(A[843]), .B(n349), .Z(O[843]) );
  AND U524 ( .A(S), .B(n350), .Z(n349) );
  XOR U525 ( .A(B[843]), .B(A[843]), .Z(n350) );
  XOR U526 ( .A(A[842]), .B(n351), .Z(O[842]) );
  AND U527 ( .A(S), .B(n352), .Z(n351) );
  XOR U528 ( .A(B[842]), .B(A[842]), .Z(n352) );
  XOR U529 ( .A(A[841]), .B(n353), .Z(O[841]) );
  AND U530 ( .A(S), .B(n354), .Z(n353) );
  XOR U531 ( .A(B[841]), .B(A[841]), .Z(n354) );
  XOR U532 ( .A(A[840]), .B(n355), .Z(O[840]) );
  AND U533 ( .A(S), .B(n356), .Z(n355) );
  XOR U534 ( .A(B[840]), .B(A[840]), .Z(n356) );
  XOR U535 ( .A(A[83]), .B(n357), .Z(O[83]) );
  AND U536 ( .A(S), .B(n358), .Z(n357) );
  XOR U537 ( .A(B[83]), .B(A[83]), .Z(n358) );
  XOR U538 ( .A(A[839]), .B(n359), .Z(O[839]) );
  AND U539 ( .A(S), .B(n360), .Z(n359) );
  XOR U540 ( .A(B[839]), .B(A[839]), .Z(n360) );
  XOR U541 ( .A(A[838]), .B(n361), .Z(O[838]) );
  AND U542 ( .A(S), .B(n362), .Z(n361) );
  XOR U543 ( .A(B[838]), .B(A[838]), .Z(n362) );
  XOR U544 ( .A(A[837]), .B(n363), .Z(O[837]) );
  AND U545 ( .A(S), .B(n364), .Z(n363) );
  XOR U546 ( .A(B[837]), .B(A[837]), .Z(n364) );
  XOR U547 ( .A(A[836]), .B(n365), .Z(O[836]) );
  AND U548 ( .A(S), .B(n366), .Z(n365) );
  XOR U549 ( .A(B[836]), .B(A[836]), .Z(n366) );
  XOR U550 ( .A(A[835]), .B(n367), .Z(O[835]) );
  AND U551 ( .A(S), .B(n368), .Z(n367) );
  XOR U552 ( .A(B[835]), .B(A[835]), .Z(n368) );
  XOR U553 ( .A(A[834]), .B(n369), .Z(O[834]) );
  AND U554 ( .A(S), .B(n370), .Z(n369) );
  XOR U555 ( .A(B[834]), .B(A[834]), .Z(n370) );
  XOR U556 ( .A(A[833]), .B(n371), .Z(O[833]) );
  AND U557 ( .A(S), .B(n372), .Z(n371) );
  XOR U558 ( .A(B[833]), .B(A[833]), .Z(n372) );
  XOR U559 ( .A(A[832]), .B(n373), .Z(O[832]) );
  AND U560 ( .A(S), .B(n374), .Z(n373) );
  XOR U561 ( .A(B[832]), .B(A[832]), .Z(n374) );
  XOR U562 ( .A(A[831]), .B(n375), .Z(O[831]) );
  AND U563 ( .A(S), .B(n376), .Z(n375) );
  XOR U564 ( .A(B[831]), .B(A[831]), .Z(n376) );
  XOR U565 ( .A(A[830]), .B(n377), .Z(O[830]) );
  AND U566 ( .A(S), .B(n378), .Z(n377) );
  XOR U567 ( .A(B[830]), .B(A[830]), .Z(n378) );
  XOR U568 ( .A(A[82]), .B(n379), .Z(O[82]) );
  AND U569 ( .A(S), .B(n380), .Z(n379) );
  XOR U570 ( .A(B[82]), .B(A[82]), .Z(n380) );
  XOR U571 ( .A(A[829]), .B(n381), .Z(O[829]) );
  AND U572 ( .A(S), .B(n382), .Z(n381) );
  XOR U573 ( .A(B[829]), .B(A[829]), .Z(n382) );
  XOR U574 ( .A(A[828]), .B(n383), .Z(O[828]) );
  AND U575 ( .A(S), .B(n384), .Z(n383) );
  XOR U576 ( .A(B[828]), .B(A[828]), .Z(n384) );
  XOR U577 ( .A(A[827]), .B(n385), .Z(O[827]) );
  AND U578 ( .A(S), .B(n386), .Z(n385) );
  XOR U579 ( .A(B[827]), .B(A[827]), .Z(n386) );
  XOR U580 ( .A(A[826]), .B(n387), .Z(O[826]) );
  AND U581 ( .A(S), .B(n388), .Z(n387) );
  XOR U582 ( .A(B[826]), .B(A[826]), .Z(n388) );
  XOR U583 ( .A(A[825]), .B(n389), .Z(O[825]) );
  AND U584 ( .A(S), .B(n390), .Z(n389) );
  XOR U585 ( .A(B[825]), .B(A[825]), .Z(n390) );
  XOR U586 ( .A(A[824]), .B(n391), .Z(O[824]) );
  AND U587 ( .A(S), .B(n392), .Z(n391) );
  XOR U588 ( .A(B[824]), .B(A[824]), .Z(n392) );
  XOR U589 ( .A(A[823]), .B(n393), .Z(O[823]) );
  AND U590 ( .A(S), .B(n394), .Z(n393) );
  XOR U591 ( .A(B[823]), .B(A[823]), .Z(n394) );
  XOR U592 ( .A(A[822]), .B(n395), .Z(O[822]) );
  AND U593 ( .A(S), .B(n396), .Z(n395) );
  XOR U594 ( .A(B[822]), .B(A[822]), .Z(n396) );
  XOR U595 ( .A(A[821]), .B(n397), .Z(O[821]) );
  AND U596 ( .A(S), .B(n398), .Z(n397) );
  XOR U597 ( .A(B[821]), .B(A[821]), .Z(n398) );
  XOR U598 ( .A(A[820]), .B(n399), .Z(O[820]) );
  AND U599 ( .A(S), .B(n400), .Z(n399) );
  XOR U600 ( .A(B[820]), .B(A[820]), .Z(n400) );
  XOR U601 ( .A(A[81]), .B(n401), .Z(O[81]) );
  AND U602 ( .A(S), .B(n402), .Z(n401) );
  XOR U603 ( .A(B[81]), .B(A[81]), .Z(n402) );
  XOR U604 ( .A(A[819]), .B(n403), .Z(O[819]) );
  AND U605 ( .A(S), .B(n404), .Z(n403) );
  XOR U606 ( .A(B[819]), .B(A[819]), .Z(n404) );
  XOR U607 ( .A(A[818]), .B(n405), .Z(O[818]) );
  AND U608 ( .A(S), .B(n406), .Z(n405) );
  XOR U609 ( .A(B[818]), .B(A[818]), .Z(n406) );
  XOR U610 ( .A(A[817]), .B(n407), .Z(O[817]) );
  AND U611 ( .A(S), .B(n408), .Z(n407) );
  XOR U612 ( .A(B[817]), .B(A[817]), .Z(n408) );
  XOR U613 ( .A(A[816]), .B(n409), .Z(O[816]) );
  AND U614 ( .A(S), .B(n410), .Z(n409) );
  XOR U615 ( .A(B[816]), .B(A[816]), .Z(n410) );
  XOR U616 ( .A(A[815]), .B(n411), .Z(O[815]) );
  AND U617 ( .A(S), .B(n412), .Z(n411) );
  XOR U618 ( .A(B[815]), .B(A[815]), .Z(n412) );
  XOR U619 ( .A(A[814]), .B(n413), .Z(O[814]) );
  AND U620 ( .A(S), .B(n414), .Z(n413) );
  XOR U621 ( .A(B[814]), .B(A[814]), .Z(n414) );
  XOR U622 ( .A(A[813]), .B(n415), .Z(O[813]) );
  AND U623 ( .A(S), .B(n416), .Z(n415) );
  XOR U624 ( .A(B[813]), .B(A[813]), .Z(n416) );
  XOR U625 ( .A(A[812]), .B(n417), .Z(O[812]) );
  AND U626 ( .A(S), .B(n418), .Z(n417) );
  XOR U627 ( .A(B[812]), .B(A[812]), .Z(n418) );
  XOR U628 ( .A(A[811]), .B(n419), .Z(O[811]) );
  AND U629 ( .A(S), .B(n420), .Z(n419) );
  XOR U630 ( .A(B[811]), .B(A[811]), .Z(n420) );
  XOR U631 ( .A(A[810]), .B(n421), .Z(O[810]) );
  AND U632 ( .A(S), .B(n422), .Z(n421) );
  XOR U633 ( .A(B[810]), .B(A[810]), .Z(n422) );
  XOR U634 ( .A(A[80]), .B(n423), .Z(O[80]) );
  AND U635 ( .A(S), .B(n424), .Z(n423) );
  XOR U636 ( .A(B[80]), .B(A[80]), .Z(n424) );
  XOR U637 ( .A(A[809]), .B(n425), .Z(O[809]) );
  AND U638 ( .A(S), .B(n426), .Z(n425) );
  XOR U639 ( .A(B[809]), .B(A[809]), .Z(n426) );
  XOR U640 ( .A(A[808]), .B(n427), .Z(O[808]) );
  AND U641 ( .A(S), .B(n428), .Z(n427) );
  XOR U642 ( .A(B[808]), .B(A[808]), .Z(n428) );
  XOR U643 ( .A(A[807]), .B(n429), .Z(O[807]) );
  AND U644 ( .A(S), .B(n430), .Z(n429) );
  XOR U645 ( .A(B[807]), .B(A[807]), .Z(n430) );
  XOR U646 ( .A(A[806]), .B(n431), .Z(O[806]) );
  AND U647 ( .A(S), .B(n432), .Z(n431) );
  XOR U648 ( .A(B[806]), .B(A[806]), .Z(n432) );
  XOR U649 ( .A(A[805]), .B(n433), .Z(O[805]) );
  AND U650 ( .A(S), .B(n434), .Z(n433) );
  XOR U651 ( .A(B[805]), .B(A[805]), .Z(n434) );
  XOR U652 ( .A(A[804]), .B(n435), .Z(O[804]) );
  AND U653 ( .A(S), .B(n436), .Z(n435) );
  XOR U654 ( .A(B[804]), .B(A[804]), .Z(n436) );
  XOR U655 ( .A(A[803]), .B(n437), .Z(O[803]) );
  AND U656 ( .A(S), .B(n438), .Z(n437) );
  XOR U657 ( .A(B[803]), .B(A[803]), .Z(n438) );
  XOR U658 ( .A(A[802]), .B(n439), .Z(O[802]) );
  AND U659 ( .A(S), .B(n440), .Z(n439) );
  XOR U660 ( .A(B[802]), .B(A[802]), .Z(n440) );
  XOR U661 ( .A(A[801]), .B(n441), .Z(O[801]) );
  AND U662 ( .A(S), .B(n442), .Z(n441) );
  XOR U663 ( .A(B[801]), .B(A[801]), .Z(n442) );
  XOR U664 ( .A(A[800]), .B(n443), .Z(O[800]) );
  AND U665 ( .A(S), .B(n444), .Z(n443) );
  XOR U666 ( .A(B[800]), .B(A[800]), .Z(n444) );
  XOR U667 ( .A(A[7]), .B(n445), .Z(O[7]) );
  AND U668 ( .A(S), .B(n446), .Z(n445) );
  XOR U669 ( .A(B[7]), .B(A[7]), .Z(n446) );
  XOR U670 ( .A(A[79]), .B(n447), .Z(O[79]) );
  AND U671 ( .A(S), .B(n448), .Z(n447) );
  XOR U672 ( .A(B[79]), .B(A[79]), .Z(n448) );
  XOR U673 ( .A(A[799]), .B(n449), .Z(O[799]) );
  AND U674 ( .A(S), .B(n450), .Z(n449) );
  XOR U675 ( .A(B[799]), .B(A[799]), .Z(n450) );
  XOR U676 ( .A(A[798]), .B(n451), .Z(O[798]) );
  AND U677 ( .A(S), .B(n452), .Z(n451) );
  XOR U678 ( .A(B[798]), .B(A[798]), .Z(n452) );
  XOR U679 ( .A(A[797]), .B(n453), .Z(O[797]) );
  AND U680 ( .A(S), .B(n454), .Z(n453) );
  XOR U681 ( .A(B[797]), .B(A[797]), .Z(n454) );
  XOR U682 ( .A(A[796]), .B(n455), .Z(O[796]) );
  AND U683 ( .A(S), .B(n456), .Z(n455) );
  XOR U684 ( .A(B[796]), .B(A[796]), .Z(n456) );
  XOR U685 ( .A(A[795]), .B(n457), .Z(O[795]) );
  AND U686 ( .A(S), .B(n458), .Z(n457) );
  XOR U687 ( .A(B[795]), .B(A[795]), .Z(n458) );
  XOR U688 ( .A(A[794]), .B(n459), .Z(O[794]) );
  AND U689 ( .A(S), .B(n460), .Z(n459) );
  XOR U690 ( .A(B[794]), .B(A[794]), .Z(n460) );
  XOR U691 ( .A(A[793]), .B(n461), .Z(O[793]) );
  AND U692 ( .A(S), .B(n462), .Z(n461) );
  XOR U693 ( .A(B[793]), .B(A[793]), .Z(n462) );
  XOR U694 ( .A(A[792]), .B(n463), .Z(O[792]) );
  AND U695 ( .A(S), .B(n464), .Z(n463) );
  XOR U696 ( .A(B[792]), .B(A[792]), .Z(n464) );
  XOR U697 ( .A(A[791]), .B(n465), .Z(O[791]) );
  AND U698 ( .A(S), .B(n466), .Z(n465) );
  XOR U699 ( .A(B[791]), .B(A[791]), .Z(n466) );
  XOR U700 ( .A(A[790]), .B(n467), .Z(O[790]) );
  AND U701 ( .A(S), .B(n468), .Z(n467) );
  XOR U702 ( .A(B[790]), .B(A[790]), .Z(n468) );
  XOR U703 ( .A(A[78]), .B(n469), .Z(O[78]) );
  AND U704 ( .A(S), .B(n470), .Z(n469) );
  XOR U705 ( .A(B[78]), .B(A[78]), .Z(n470) );
  XOR U706 ( .A(A[789]), .B(n471), .Z(O[789]) );
  AND U707 ( .A(S), .B(n472), .Z(n471) );
  XOR U708 ( .A(B[789]), .B(A[789]), .Z(n472) );
  XOR U709 ( .A(A[788]), .B(n473), .Z(O[788]) );
  AND U710 ( .A(S), .B(n474), .Z(n473) );
  XOR U711 ( .A(B[788]), .B(A[788]), .Z(n474) );
  XOR U712 ( .A(A[787]), .B(n475), .Z(O[787]) );
  AND U713 ( .A(S), .B(n476), .Z(n475) );
  XOR U714 ( .A(B[787]), .B(A[787]), .Z(n476) );
  XOR U715 ( .A(A[786]), .B(n477), .Z(O[786]) );
  AND U716 ( .A(S), .B(n478), .Z(n477) );
  XOR U717 ( .A(B[786]), .B(A[786]), .Z(n478) );
  XOR U718 ( .A(A[785]), .B(n479), .Z(O[785]) );
  AND U719 ( .A(S), .B(n480), .Z(n479) );
  XOR U720 ( .A(B[785]), .B(A[785]), .Z(n480) );
  XOR U721 ( .A(A[784]), .B(n481), .Z(O[784]) );
  AND U722 ( .A(S), .B(n482), .Z(n481) );
  XOR U723 ( .A(B[784]), .B(A[784]), .Z(n482) );
  XOR U724 ( .A(A[783]), .B(n483), .Z(O[783]) );
  AND U725 ( .A(S), .B(n484), .Z(n483) );
  XOR U726 ( .A(B[783]), .B(A[783]), .Z(n484) );
  XOR U727 ( .A(A[782]), .B(n485), .Z(O[782]) );
  AND U728 ( .A(S), .B(n486), .Z(n485) );
  XOR U729 ( .A(B[782]), .B(A[782]), .Z(n486) );
  XOR U730 ( .A(A[781]), .B(n487), .Z(O[781]) );
  AND U731 ( .A(S), .B(n488), .Z(n487) );
  XOR U732 ( .A(B[781]), .B(A[781]), .Z(n488) );
  XOR U733 ( .A(A[780]), .B(n489), .Z(O[780]) );
  AND U734 ( .A(S), .B(n490), .Z(n489) );
  XOR U735 ( .A(B[780]), .B(A[780]), .Z(n490) );
  XOR U736 ( .A(A[77]), .B(n491), .Z(O[77]) );
  AND U737 ( .A(S), .B(n492), .Z(n491) );
  XOR U738 ( .A(B[77]), .B(A[77]), .Z(n492) );
  XOR U739 ( .A(A[779]), .B(n493), .Z(O[779]) );
  AND U740 ( .A(S), .B(n494), .Z(n493) );
  XOR U741 ( .A(B[779]), .B(A[779]), .Z(n494) );
  XOR U742 ( .A(A[778]), .B(n495), .Z(O[778]) );
  AND U743 ( .A(S), .B(n496), .Z(n495) );
  XOR U744 ( .A(B[778]), .B(A[778]), .Z(n496) );
  XOR U745 ( .A(A[777]), .B(n497), .Z(O[777]) );
  AND U746 ( .A(S), .B(n498), .Z(n497) );
  XOR U747 ( .A(B[777]), .B(A[777]), .Z(n498) );
  XOR U748 ( .A(A[776]), .B(n499), .Z(O[776]) );
  AND U749 ( .A(S), .B(n500), .Z(n499) );
  XOR U750 ( .A(B[776]), .B(A[776]), .Z(n500) );
  XOR U751 ( .A(A[775]), .B(n501), .Z(O[775]) );
  AND U752 ( .A(S), .B(n502), .Z(n501) );
  XOR U753 ( .A(B[775]), .B(A[775]), .Z(n502) );
  XOR U754 ( .A(A[774]), .B(n503), .Z(O[774]) );
  AND U755 ( .A(S), .B(n504), .Z(n503) );
  XOR U756 ( .A(B[774]), .B(A[774]), .Z(n504) );
  XOR U757 ( .A(A[773]), .B(n505), .Z(O[773]) );
  AND U758 ( .A(S), .B(n506), .Z(n505) );
  XOR U759 ( .A(B[773]), .B(A[773]), .Z(n506) );
  XOR U760 ( .A(A[772]), .B(n507), .Z(O[772]) );
  AND U761 ( .A(S), .B(n508), .Z(n507) );
  XOR U762 ( .A(B[772]), .B(A[772]), .Z(n508) );
  XOR U763 ( .A(A[771]), .B(n509), .Z(O[771]) );
  AND U764 ( .A(S), .B(n510), .Z(n509) );
  XOR U765 ( .A(B[771]), .B(A[771]), .Z(n510) );
  XOR U766 ( .A(A[770]), .B(n511), .Z(O[770]) );
  AND U767 ( .A(S), .B(n512), .Z(n511) );
  XOR U768 ( .A(B[770]), .B(A[770]), .Z(n512) );
  XOR U769 ( .A(A[76]), .B(n513), .Z(O[76]) );
  AND U770 ( .A(S), .B(n514), .Z(n513) );
  XOR U771 ( .A(B[76]), .B(A[76]), .Z(n514) );
  XOR U772 ( .A(A[769]), .B(n515), .Z(O[769]) );
  AND U773 ( .A(S), .B(n516), .Z(n515) );
  XOR U774 ( .A(B[769]), .B(A[769]), .Z(n516) );
  XOR U775 ( .A(A[768]), .B(n517), .Z(O[768]) );
  AND U776 ( .A(S), .B(n518), .Z(n517) );
  XOR U777 ( .A(B[768]), .B(A[768]), .Z(n518) );
  XOR U778 ( .A(A[767]), .B(n519), .Z(O[767]) );
  AND U779 ( .A(S), .B(n520), .Z(n519) );
  XOR U780 ( .A(B[767]), .B(A[767]), .Z(n520) );
  XOR U781 ( .A(A[766]), .B(n521), .Z(O[766]) );
  AND U782 ( .A(S), .B(n522), .Z(n521) );
  XOR U783 ( .A(B[766]), .B(A[766]), .Z(n522) );
  XOR U784 ( .A(A[765]), .B(n523), .Z(O[765]) );
  AND U785 ( .A(S), .B(n524), .Z(n523) );
  XOR U786 ( .A(B[765]), .B(A[765]), .Z(n524) );
  XOR U787 ( .A(A[764]), .B(n525), .Z(O[764]) );
  AND U788 ( .A(S), .B(n526), .Z(n525) );
  XOR U789 ( .A(B[764]), .B(A[764]), .Z(n526) );
  XOR U790 ( .A(A[763]), .B(n527), .Z(O[763]) );
  AND U791 ( .A(S), .B(n528), .Z(n527) );
  XOR U792 ( .A(B[763]), .B(A[763]), .Z(n528) );
  XOR U793 ( .A(A[762]), .B(n529), .Z(O[762]) );
  AND U794 ( .A(S), .B(n530), .Z(n529) );
  XOR U795 ( .A(B[762]), .B(A[762]), .Z(n530) );
  XOR U796 ( .A(A[761]), .B(n531), .Z(O[761]) );
  AND U797 ( .A(S), .B(n532), .Z(n531) );
  XOR U798 ( .A(B[761]), .B(A[761]), .Z(n532) );
  XOR U799 ( .A(A[760]), .B(n533), .Z(O[760]) );
  AND U800 ( .A(S), .B(n534), .Z(n533) );
  XOR U801 ( .A(B[760]), .B(A[760]), .Z(n534) );
  XOR U802 ( .A(A[75]), .B(n535), .Z(O[75]) );
  AND U803 ( .A(S), .B(n536), .Z(n535) );
  XOR U804 ( .A(B[75]), .B(A[75]), .Z(n536) );
  XOR U805 ( .A(A[759]), .B(n537), .Z(O[759]) );
  AND U806 ( .A(S), .B(n538), .Z(n537) );
  XOR U807 ( .A(B[759]), .B(A[759]), .Z(n538) );
  XOR U808 ( .A(A[758]), .B(n539), .Z(O[758]) );
  AND U809 ( .A(S), .B(n540), .Z(n539) );
  XOR U810 ( .A(B[758]), .B(A[758]), .Z(n540) );
  XOR U811 ( .A(A[757]), .B(n541), .Z(O[757]) );
  AND U812 ( .A(S), .B(n542), .Z(n541) );
  XOR U813 ( .A(B[757]), .B(A[757]), .Z(n542) );
  XOR U814 ( .A(A[756]), .B(n543), .Z(O[756]) );
  AND U815 ( .A(S), .B(n544), .Z(n543) );
  XOR U816 ( .A(B[756]), .B(A[756]), .Z(n544) );
  XOR U817 ( .A(A[755]), .B(n545), .Z(O[755]) );
  AND U818 ( .A(S), .B(n546), .Z(n545) );
  XOR U819 ( .A(B[755]), .B(A[755]), .Z(n546) );
  XOR U820 ( .A(A[754]), .B(n547), .Z(O[754]) );
  AND U821 ( .A(S), .B(n548), .Z(n547) );
  XOR U822 ( .A(B[754]), .B(A[754]), .Z(n548) );
  XOR U823 ( .A(A[753]), .B(n549), .Z(O[753]) );
  AND U824 ( .A(S), .B(n550), .Z(n549) );
  XOR U825 ( .A(B[753]), .B(A[753]), .Z(n550) );
  XOR U826 ( .A(A[752]), .B(n551), .Z(O[752]) );
  AND U827 ( .A(S), .B(n552), .Z(n551) );
  XOR U828 ( .A(B[752]), .B(A[752]), .Z(n552) );
  XOR U829 ( .A(A[751]), .B(n553), .Z(O[751]) );
  AND U830 ( .A(S), .B(n554), .Z(n553) );
  XOR U831 ( .A(B[751]), .B(A[751]), .Z(n554) );
  XOR U832 ( .A(A[750]), .B(n555), .Z(O[750]) );
  AND U833 ( .A(S), .B(n556), .Z(n555) );
  XOR U834 ( .A(B[750]), .B(A[750]), .Z(n556) );
  XOR U835 ( .A(A[74]), .B(n557), .Z(O[74]) );
  AND U836 ( .A(S), .B(n558), .Z(n557) );
  XOR U837 ( .A(B[74]), .B(A[74]), .Z(n558) );
  XOR U838 ( .A(A[749]), .B(n559), .Z(O[749]) );
  AND U839 ( .A(S), .B(n560), .Z(n559) );
  XOR U840 ( .A(B[749]), .B(A[749]), .Z(n560) );
  XOR U841 ( .A(A[748]), .B(n561), .Z(O[748]) );
  AND U842 ( .A(S), .B(n562), .Z(n561) );
  XOR U843 ( .A(B[748]), .B(A[748]), .Z(n562) );
  XOR U844 ( .A(A[747]), .B(n563), .Z(O[747]) );
  AND U845 ( .A(S), .B(n564), .Z(n563) );
  XOR U846 ( .A(B[747]), .B(A[747]), .Z(n564) );
  XOR U847 ( .A(A[746]), .B(n565), .Z(O[746]) );
  AND U848 ( .A(S), .B(n566), .Z(n565) );
  XOR U849 ( .A(B[746]), .B(A[746]), .Z(n566) );
  XOR U850 ( .A(A[745]), .B(n567), .Z(O[745]) );
  AND U851 ( .A(S), .B(n568), .Z(n567) );
  XOR U852 ( .A(B[745]), .B(A[745]), .Z(n568) );
  XOR U853 ( .A(A[744]), .B(n569), .Z(O[744]) );
  AND U854 ( .A(S), .B(n570), .Z(n569) );
  XOR U855 ( .A(B[744]), .B(A[744]), .Z(n570) );
  XOR U856 ( .A(A[743]), .B(n571), .Z(O[743]) );
  AND U857 ( .A(S), .B(n572), .Z(n571) );
  XOR U858 ( .A(B[743]), .B(A[743]), .Z(n572) );
  XOR U859 ( .A(A[742]), .B(n573), .Z(O[742]) );
  AND U860 ( .A(S), .B(n574), .Z(n573) );
  XOR U861 ( .A(B[742]), .B(A[742]), .Z(n574) );
  XOR U862 ( .A(A[741]), .B(n575), .Z(O[741]) );
  AND U863 ( .A(S), .B(n576), .Z(n575) );
  XOR U864 ( .A(B[741]), .B(A[741]), .Z(n576) );
  XOR U865 ( .A(A[740]), .B(n577), .Z(O[740]) );
  AND U866 ( .A(S), .B(n578), .Z(n577) );
  XOR U867 ( .A(B[740]), .B(A[740]), .Z(n578) );
  XOR U868 ( .A(A[73]), .B(n579), .Z(O[73]) );
  AND U869 ( .A(S), .B(n580), .Z(n579) );
  XOR U870 ( .A(B[73]), .B(A[73]), .Z(n580) );
  XOR U871 ( .A(A[739]), .B(n581), .Z(O[739]) );
  AND U872 ( .A(S), .B(n582), .Z(n581) );
  XOR U873 ( .A(B[739]), .B(A[739]), .Z(n582) );
  XOR U874 ( .A(A[738]), .B(n583), .Z(O[738]) );
  AND U875 ( .A(S), .B(n584), .Z(n583) );
  XOR U876 ( .A(B[738]), .B(A[738]), .Z(n584) );
  XOR U877 ( .A(A[737]), .B(n585), .Z(O[737]) );
  AND U878 ( .A(S), .B(n586), .Z(n585) );
  XOR U879 ( .A(B[737]), .B(A[737]), .Z(n586) );
  XOR U880 ( .A(A[736]), .B(n587), .Z(O[736]) );
  AND U881 ( .A(S), .B(n588), .Z(n587) );
  XOR U882 ( .A(B[736]), .B(A[736]), .Z(n588) );
  XOR U883 ( .A(A[735]), .B(n589), .Z(O[735]) );
  AND U884 ( .A(S), .B(n590), .Z(n589) );
  XOR U885 ( .A(B[735]), .B(A[735]), .Z(n590) );
  XOR U886 ( .A(A[734]), .B(n591), .Z(O[734]) );
  AND U887 ( .A(S), .B(n592), .Z(n591) );
  XOR U888 ( .A(B[734]), .B(A[734]), .Z(n592) );
  XOR U889 ( .A(A[733]), .B(n593), .Z(O[733]) );
  AND U890 ( .A(S), .B(n594), .Z(n593) );
  XOR U891 ( .A(B[733]), .B(A[733]), .Z(n594) );
  XOR U892 ( .A(A[732]), .B(n595), .Z(O[732]) );
  AND U893 ( .A(S), .B(n596), .Z(n595) );
  XOR U894 ( .A(B[732]), .B(A[732]), .Z(n596) );
  XOR U895 ( .A(A[731]), .B(n597), .Z(O[731]) );
  AND U896 ( .A(S), .B(n598), .Z(n597) );
  XOR U897 ( .A(B[731]), .B(A[731]), .Z(n598) );
  XOR U898 ( .A(A[730]), .B(n599), .Z(O[730]) );
  AND U899 ( .A(S), .B(n600), .Z(n599) );
  XOR U900 ( .A(B[730]), .B(A[730]), .Z(n600) );
  XOR U901 ( .A(A[72]), .B(n601), .Z(O[72]) );
  AND U902 ( .A(S), .B(n602), .Z(n601) );
  XOR U903 ( .A(B[72]), .B(A[72]), .Z(n602) );
  XOR U904 ( .A(A[729]), .B(n603), .Z(O[729]) );
  AND U905 ( .A(S), .B(n604), .Z(n603) );
  XOR U906 ( .A(B[729]), .B(A[729]), .Z(n604) );
  XOR U907 ( .A(A[728]), .B(n605), .Z(O[728]) );
  AND U908 ( .A(S), .B(n606), .Z(n605) );
  XOR U909 ( .A(B[728]), .B(A[728]), .Z(n606) );
  XOR U910 ( .A(A[727]), .B(n607), .Z(O[727]) );
  AND U911 ( .A(S), .B(n608), .Z(n607) );
  XOR U912 ( .A(B[727]), .B(A[727]), .Z(n608) );
  XOR U913 ( .A(A[726]), .B(n609), .Z(O[726]) );
  AND U914 ( .A(S), .B(n610), .Z(n609) );
  XOR U915 ( .A(B[726]), .B(A[726]), .Z(n610) );
  XOR U916 ( .A(A[725]), .B(n611), .Z(O[725]) );
  AND U917 ( .A(S), .B(n612), .Z(n611) );
  XOR U918 ( .A(B[725]), .B(A[725]), .Z(n612) );
  XOR U919 ( .A(A[724]), .B(n613), .Z(O[724]) );
  AND U920 ( .A(S), .B(n614), .Z(n613) );
  XOR U921 ( .A(B[724]), .B(A[724]), .Z(n614) );
  XOR U922 ( .A(A[723]), .B(n615), .Z(O[723]) );
  AND U923 ( .A(S), .B(n616), .Z(n615) );
  XOR U924 ( .A(B[723]), .B(A[723]), .Z(n616) );
  XOR U925 ( .A(A[722]), .B(n617), .Z(O[722]) );
  AND U926 ( .A(S), .B(n618), .Z(n617) );
  XOR U927 ( .A(B[722]), .B(A[722]), .Z(n618) );
  XOR U928 ( .A(A[721]), .B(n619), .Z(O[721]) );
  AND U929 ( .A(S), .B(n620), .Z(n619) );
  XOR U930 ( .A(B[721]), .B(A[721]), .Z(n620) );
  XOR U931 ( .A(A[720]), .B(n621), .Z(O[720]) );
  AND U932 ( .A(S), .B(n622), .Z(n621) );
  XOR U933 ( .A(B[720]), .B(A[720]), .Z(n622) );
  XOR U934 ( .A(A[71]), .B(n623), .Z(O[71]) );
  AND U935 ( .A(S), .B(n624), .Z(n623) );
  XOR U936 ( .A(B[71]), .B(A[71]), .Z(n624) );
  XOR U937 ( .A(A[719]), .B(n625), .Z(O[719]) );
  AND U938 ( .A(S), .B(n626), .Z(n625) );
  XOR U939 ( .A(B[719]), .B(A[719]), .Z(n626) );
  XOR U940 ( .A(A[718]), .B(n627), .Z(O[718]) );
  AND U941 ( .A(S), .B(n628), .Z(n627) );
  XOR U942 ( .A(B[718]), .B(A[718]), .Z(n628) );
  XOR U943 ( .A(A[717]), .B(n629), .Z(O[717]) );
  AND U944 ( .A(S), .B(n630), .Z(n629) );
  XOR U945 ( .A(B[717]), .B(A[717]), .Z(n630) );
  XOR U946 ( .A(A[716]), .B(n631), .Z(O[716]) );
  AND U947 ( .A(S), .B(n632), .Z(n631) );
  XOR U948 ( .A(B[716]), .B(A[716]), .Z(n632) );
  XOR U949 ( .A(A[715]), .B(n633), .Z(O[715]) );
  AND U950 ( .A(S), .B(n634), .Z(n633) );
  XOR U951 ( .A(B[715]), .B(A[715]), .Z(n634) );
  XOR U952 ( .A(A[714]), .B(n635), .Z(O[714]) );
  AND U953 ( .A(S), .B(n636), .Z(n635) );
  XOR U954 ( .A(B[714]), .B(A[714]), .Z(n636) );
  XOR U955 ( .A(A[713]), .B(n637), .Z(O[713]) );
  AND U956 ( .A(S), .B(n638), .Z(n637) );
  XOR U957 ( .A(B[713]), .B(A[713]), .Z(n638) );
  XOR U958 ( .A(A[712]), .B(n639), .Z(O[712]) );
  AND U959 ( .A(S), .B(n640), .Z(n639) );
  XOR U960 ( .A(B[712]), .B(A[712]), .Z(n640) );
  XOR U961 ( .A(A[711]), .B(n641), .Z(O[711]) );
  AND U962 ( .A(S), .B(n642), .Z(n641) );
  XOR U963 ( .A(B[711]), .B(A[711]), .Z(n642) );
  XOR U964 ( .A(A[710]), .B(n643), .Z(O[710]) );
  AND U965 ( .A(S), .B(n644), .Z(n643) );
  XOR U966 ( .A(B[710]), .B(A[710]), .Z(n644) );
  XOR U967 ( .A(A[70]), .B(n645), .Z(O[70]) );
  AND U968 ( .A(S), .B(n646), .Z(n645) );
  XOR U969 ( .A(B[70]), .B(A[70]), .Z(n646) );
  XOR U970 ( .A(A[709]), .B(n647), .Z(O[709]) );
  AND U971 ( .A(S), .B(n648), .Z(n647) );
  XOR U972 ( .A(B[709]), .B(A[709]), .Z(n648) );
  XOR U973 ( .A(A[708]), .B(n649), .Z(O[708]) );
  AND U974 ( .A(S), .B(n650), .Z(n649) );
  XOR U975 ( .A(B[708]), .B(A[708]), .Z(n650) );
  XOR U976 ( .A(A[707]), .B(n651), .Z(O[707]) );
  AND U977 ( .A(S), .B(n652), .Z(n651) );
  XOR U978 ( .A(B[707]), .B(A[707]), .Z(n652) );
  XOR U979 ( .A(A[706]), .B(n653), .Z(O[706]) );
  AND U980 ( .A(S), .B(n654), .Z(n653) );
  XOR U981 ( .A(B[706]), .B(A[706]), .Z(n654) );
  XOR U982 ( .A(A[705]), .B(n655), .Z(O[705]) );
  AND U983 ( .A(S), .B(n656), .Z(n655) );
  XOR U984 ( .A(B[705]), .B(A[705]), .Z(n656) );
  XOR U985 ( .A(A[704]), .B(n657), .Z(O[704]) );
  AND U986 ( .A(S), .B(n658), .Z(n657) );
  XOR U987 ( .A(B[704]), .B(A[704]), .Z(n658) );
  XOR U988 ( .A(A[703]), .B(n659), .Z(O[703]) );
  AND U989 ( .A(S), .B(n660), .Z(n659) );
  XOR U990 ( .A(B[703]), .B(A[703]), .Z(n660) );
  XOR U991 ( .A(A[702]), .B(n661), .Z(O[702]) );
  AND U992 ( .A(S), .B(n662), .Z(n661) );
  XOR U993 ( .A(B[702]), .B(A[702]), .Z(n662) );
  XOR U994 ( .A(A[701]), .B(n663), .Z(O[701]) );
  AND U995 ( .A(S), .B(n664), .Z(n663) );
  XOR U996 ( .A(B[701]), .B(A[701]), .Z(n664) );
  XOR U997 ( .A(A[700]), .B(n665), .Z(O[700]) );
  AND U998 ( .A(S), .B(n666), .Z(n665) );
  XOR U999 ( .A(B[700]), .B(A[700]), .Z(n666) );
  XOR U1000 ( .A(A[6]), .B(n667), .Z(O[6]) );
  AND U1001 ( .A(S), .B(n668), .Z(n667) );
  XOR U1002 ( .A(B[6]), .B(A[6]), .Z(n668) );
  XOR U1003 ( .A(A[69]), .B(n669), .Z(O[69]) );
  AND U1004 ( .A(S), .B(n670), .Z(n669) );
  XOR U1005 ( .A(B[69]), .B(A[69]), .Z(n670) );
  XOR U1006 ( .A(A[699]), .B(n671), .Z(O[699]) );
  AND U1007 ( .A(S), .B(n672), .Z(n671) );
  XOR U1008 ( .A(B[699]), .B(A[699]), .Z(n672) );
  XOR U1009 ( .A(A[698]), .B(n673), .Z(O[698]) );
  AND U1010 ( .A(S), .B(n674), .Z(n673) );
  XOR U1011 ( .A(B[698]), .B(A[698]), .Z(n674) );
  XOR U1012 ( .A(A[697]), .B(n675), .Z(O[697]) );
  AND U1013 ( .A(S), .B(n676), .Z(n675) );
  XOR U1014 ( .A(B[697]), .B(A[697]), .Z(n676) );
  XOR U1015 ( .A(A[696]), .B(n677), .Z(O[696]) );
  AND U1016 ( .A(S), .B(n678), .Z(n677) );
  XOR U1017 ( .A(B[696]), .B(A[696]), .Z(n678) );
  XOR U1018 ( .A(A[695]), .B(n679), .Z(O[695]) );
  AND U1019 ( .A(S), .B(n680), .Z(n679) );
  XOR U1020 ( .A(B[695]), .B(A[695]), .Z(n680) );
  XOR U1021 ( .A(A[694]), .B(n681), .Z(O[694]) );
  AND U1022 ( .A(S), .B(n682), .Z(n681) );
  XOR U1023 ( .A(B[694]), .B(A[694]), .Z(n682) );
  XOR U1024 ( .A(A[693]), .B(n683), .Z(O[693]) );
  AND U1025 ( .A(S), .B(n684), .Z(n683) );
  XOR U1026 ( .A(B[693]), .B(A[693]), .Z(n684) );
  XOR U1027 ( .A(A[692]), .B(n685), .Z(O[692]) );
  AND U1028 ( .A(S), .B(n686), .Z(n685) );
  XOR U1029 ( .A(B[692]), .B(A[692]), .Z(n686) );
  XOR U1030 ( .A(A[691]), .B(n687), .Z(O[691]) );
  AND U1031 ( .A(S), .B(n688), .Z(n687) );
  XOR U1032 ( .A(B[691]), .B(A[691]), .Z(n688) );
  XOR U1033 ( .A(A[690]), .B(n689), .Z(O[690]) );
  AND U1034 ( .A(S), .B(n690), .Z(n689) );
  XOR U1035 ( .A(B[690]), .B(A[690]), .Z(n690) );
  XOR U1036 ( .A(A[68]), .B(n691), .Z(O[68]) );
  AND U1037 ( .A(S), .B(n692), .Z(n691) );
  XOR U1038 ( .A(B[68]), .B(A[68]), .Z(n692) );
  XOR U1039 ( .A(A[689]), .B(n693), .Z(O[689]) );
  AND U1040 ( .A(S), .B(n694), .Z(n693) );
  XOR U1041 ( .A(B[689]), .B(A[689]), .Z(n694) );
  XOR U1042 ( .A(A[688]), .B(n695), .Z(O[688]) );
  AND U1043 ( .A(S), .B(n696), .Z(n695) );
  XOR U1044 ( .A(B[688]), .B(A[688]), .Z(n696) );
  XOR U1045 ( .A(A[687]), .B(n697), .Z(O[687]) );
  AND U1046 ( .A(S), .B(n698), .Z(n697) );
  XOR U1047 ( .A(B[687]), .B(A[687]), .Z(n698) );
  XOR U1048 ( .A(A[686]), .B(n699), .Z(O[686]) );
  AND U1049 ( .A(S), .B(n700), .Z(n699) );
  XOR U1050 ( .A(B[686]), .B(A[686]), .Z(n700) );
  XOR U1051 ( .A(A[685]), .B(n701), .Z(O[685]) );
  AND U1052 ( .A(S), .B(n702), .Z(n701) );
  XOR U1053 ( .A(B[685]), .B(A[685]), .Z(n702) );
  XOR U1054 ( .A(A[684]), .B(n703), .Z(O[684]) );
  AND U1055 ( .A(S), .B(n704), .Z(n703) );
  XOR U1056 ( .A(B[684]), .B(A[684]), .Z(n704) );
  XOR U1057 ( .A(A[683]), .B(n705), .Z(O[683]) );
  AND U1058 ( .A(S), .B(n706), .Z(n705) );
  XOR U1059 ( .A(B[683]), .B(A[683]), .Z(n706) );
  XOR U1060 ( .A(A[682]), .B(n707), .Z(O[682]) );
  AND U1061 ( .A(S), .B(n708), .Z(n707) );
  XOR U1062 ( .A(B[682]), .B(A[682]), .Z(n708) );
  XOR U1063 ( .A(A[681]), .B(n709), .Z(O[681]) );
  AND U1064 ( .A(S), .B(n710), .Z(n709) );
  XOR U1065 ( .A(B[681]), .B(A[681]), .Z(n710) );
  XOR U1066 ( .A(A[680]), .B(n711), .Z(O[680]) );
  AND U1067 ( .A(S), .B(n712), .Z(n711) );
  XOR U1068 ( .A(B[680]), .B(A[680]), .Z(n712) );
  XOR U1069 ( .A(A[67]), .B(n713), .Z(O[67]) );
  AND U1070 ( .A(S), .B(n714), .Z(n713) );
  XOR U1071 ( .A(B[67]), .B(A[67]), .Z(n714) );
  XOR U1072 ( .A(A[679]), .B(n715), .Z(O[679]) );
  AND U1073 ( .A(S), .B(n716), .Z(n715) );
  XOR U1074 ( .A(B[679]), .B(A[679]), .Z(n716) );
  XOR U1075 ( .A(A[678]), .B(n717), .Z(O[678]) );
  AND U1076 ( .A(S), .B(n718), .Z(n717) );
  XOR U1077 ( .A(B[678]), .B(A[678]), .Z(n718) );
  XOR U1078 ( .A(A[677]), .B(n719), .Z(O[677]) );
  AND U1079 ( .A(S), .B(n720), .Z(n719) );
  XOR U1080 ( .A(B[677]), .B(A[677]), .Z(n720) );
  XOR U1081 ( .A(A[676]), .B(n721), .Z(O[676]) );
  AND U1082 ( .A(S), .B(n722), .Z(n721) );
  XOR U1083 ( .A(B[676]), .B(A[676]), .Z(n722) );
  XOR U1084 ( .A(A[675]), .B(n723), .Z(O[675]) );
  AND U1085 ( .A(S), .B(n724), .Z(n723) );
  XOR U1086 ( .A(B[675]), .B(A[675]), .Z(n724) );
  XOR U1087 ( .A(A[674]), .B(n725), .Z(O[674]) );
  AND U1088 ( .A(S), .B(n726), .Z(n725) );
  XOR U1089 ( .A(B[674]), .B(A[674]), .Z(n726) );
  XOR U1090 ( .A(A[673]), .B(n727), .Z(O[673]) );
  AND U1091 ( .A(S), .B(n728), .Z(n727) );
  XOR U1092 ( .A(B[673]), .B(A[673]), .Z(n728) );
  XOR U1093 ( .A(A[672]), .B(n729), .Z(O[672]) );
  AND U1094 ( .A(S), .B(n730), .Z(n729) );
  XOR U1095 ( .A(B[672]), .B(A[672]), .Z(n730) );
  XOR U1096 ( .A(A[671]), .B(n731), .Z(O[671]) );
  AND U1097 ( .A(S), .B(n732), .Z(n731) );
  XOR U1098 ( .A(B[671]), .B(A[671]), .Z(n732) );
  XOR U1099 ( .A(A[670]), .B(n733), .Z(O[670]) );
  AND U1100 ( .A(S), .B(n734), .Z(n733) );
  XOR U1101 ( .A(B[670]), .B(A[670]), .Z(n734) );
  XOR U1102 ( .A(A[66]), .B(n735), .Z(O[66]) );
  AND U1103 ( .A(S), .B(n736), .Z(n735) );
  XOR U1104 ( .A(B[66]), .B(A[66]), .Z(n736) );
  XOR U1105 ( .A(A[669]), .B(n737), .Z(O[669]) );
  AND U1106 ( .A(S), .B(n738), .Z(n737) );
  XOR U1107 ( .A(B[669]), .B(A[669]), .Z(n738) );
  XOR U1108 ( .A(A[668]), .B(n739), .Z(O[668]) );
  AND U1109 ( .A(S), .B(n740), .Z(n739) );
  XOR U1110 ( .A(B[668]), .B(A[668]), .Z(n740) );
  XOR U1111 ( .A(A[667]), .B(n741), .Z(O[667]) );
  AND U1112 ( .A(S), .B(n742), .Z(n741) );
  XOR U1113 ( .A(B[667]), .B(A[667]), .Z(n742) );
  XOR U1114 ( .A(A[666]), .B(n743), .Z(O[666]) );
  AND U1115 ( .A(S), .B(n744), .Z(n743) );
  XOR U1116 ( .A(B[666]), .B(A[666]), .Z(n744) );
  XOR U1117 ( .A(A[665]), .B(n745), .Z(O[665]) );
  AND U1118 ( .A(S), .B(n746), .Z(n745) );
  XOR U1119 ( .A(B[665]), .B(A[665]), .Z(n746) );
  XOR U1120 ( .A(A[664]), .B(n747), .Z(O[664]) );
  AND U1121 ( .A(S), .B(n748), .Z(n747) );
  XOR U1122 ( .A(B[664]), .B(A[664]), .Z(n748) );
  XOR U1123 ( .A(A[663]), .B(n749), .Z(O[663]) );
  AND U1124 ( .A(S), .B(n750), .Z(n749) );
  XOR U1125 ( .A(B[663]), .B(A[663]), .Z(n750) );
  XOR U1126 ( .A(A[662]), .B(n751), .Z(O[662]) );
  AND U1127 ( .A(S), .B(n752), .Z(n751) );
  XOR U1128 ( .A(B[662]), .B(A[662]), .Z(n752) );
  XOR U1129 ( .A(A[661]), .B(n753), .Z(O[661]) );
  AND U1130 ( .A(S), .B(n754), .Z(n753) );
  XOR U1131 ( .A(B[661]), .B(A[661]), .Z(n754) );
  XOR U1132 ( .A(A[660]), .B(n755), .Z(O[660]) );
  AND U1133 ( .A(S), .B(n756), .Z(n755) );
  XOR U1134 ( .A(B[660]), .B(A[660]), .Z(n756) );
  XOR U1135 ( .A(A[65]), .B(n757), .Z(O[65]) );
  AND U1136 ( .A(S), .B(n758), .Z(n757) );
  XOR U1137 ( .A(B[65]), .B(A[65]), .Z(n758) );
  XOR U1138 ( .A(A[659]), .B(n759), .Z(O[659]) );
  AND U1139 ( .A(S), .B(n760), .Z(n759) );
  XOR U1140 ( .A(B[659]), .B(A[659]), .Z(n760) );
  XOR U1141 ( .A(A[658]), .B(n761), .Z(O[658]) );
  AND U1142 ( .A(S), .B(n762), .Z(n761) );
  XOR U1143 ( .A(B[658]), .B(A[658]), .Z(n762) );
  XOR U1144 ( .A(A[657]), .B(n763), .Z(O[657]) );
  AND U1145 ( .A(S), .B(n764), .Z(n763) );
  XOR U1146 ( .A(B[657]), .B(A[657]), .Z(n764) );
  XOR U1147 ( .A(A[656]), .B(n765), .Z(O[656]) );
  AND U1148 ( .A(S), .B(n766), .Z(n765) );
  XOR U1149 ( .A(B[656]), .B(A[656]), .Z(n766) );
  XOR U1150 ( .A(A[655]), .B(n767), .Z(O[655]) );
  AND U1151 ( .A(S), .B(n768), .Z(n767) );
  XOR U1152 ( .A(B[655]), .B(A[655]), .Z(n768) );
  XOR U1153 ( .A(A[654]), .B(n769), .Z(O[654]) );
  AND U1154 ( .A(S), .B(n770), .Z(n769) );
  XOR U1155 ( .A(B[654]), .B(A[654]), .Z(n770) );
  XOR U1156 ( .A(A[653]), .B(n771), .Z(O[653]) );
  AND U1157 ( .A(S), .B(n772), .Z(n771) );
  XOR U1158 ( .A(B[653]), .B(A[653]), .Z(n772) );
  XOR U1159 ( .A(A[652]), .B(n773), .Z(O[652]) );
  AND U1160 ( .A(S), .B(n774), .Z(n773) );
  XOR U1161 ( .A(B[652]), .B(A[652]), .Z(n774) );
  XOR U1162 ( .A(A[651]), .B(n775), .Z(O[651]) );
  AND U1163 ( .A(S), .B(n776), .Z(n775) );
  XOR U1164 ( .A(B[651]), .B(A[651]), .Z(n776) );
  XOR U1165 ( .A(A[650]), .B(n777), .Z(O[650]) );
  AND U1166 ( .A(S), .B(n778), .Z(n777) );
  XOR U1167 ( .A(B[650]), .B(A[650]), .Z(n778) );
  XOR U1168 ( .A(A[64]), .B(n779), .Z(O[64]) );
  AND U1169 ( .A(S), .B(n780), .Z(n779) );
  XOR U1170 ( .A(B[64]), .B(A[64]), .Z(n780) );
  XOR U1171 ( .A(A[649]), .B(n781), .Z(O[649]) );
  AND U1172 ( .A(S), .B(n782), .Z(n781) );
  XOR U1173 ( .A(B[649]), .B(A[649]), .Z(n782) );
  XOR U1174 ( .A(A[648]), .B(n783), .Z(O[648]) );
  AND U1175 ( .A(S), .B(n784), .Z(n783) );
  XOR U1176 ( .A(B[648]), .B(A[648]), .Z(n784) );
  XOR U1177 ( .A(A[647]), .B(n785), .Z(O[647]) );
  AND U1178 ( .A(S), .B(n786), .Z(n785) );
  XOR U1179 ( .A(B[647]), .B(A[647]), .Z(n786) );
  XOR U1180 ( .A(A[646]), .B(n787), .Z(O[646]) );
  AND U1181 ( .A(S), .B(n788), .Z(n787) );
  XOR U1182 ( .A(B[646]), .B(A[646]), .Z(n788) );
  XOR U1183 ( .A(A[645]), .B(n789), .Z(O[645]) );
  AND U1184 ( .A(S), .B(n790), .Z(n789) );
  XOR U1185 ( .A(B[645]), .B(A[645]), .Z(n790) );
  XOR U1186 ( .A(A[644]), .B(n791), .Z(O[644]) );
  AND U1187 ( .A(S), .B(n792), .Z(n791) );
  XOR U1188 ( .A(B[644]), .B(A[644]), .Z(n792) );
  XOR U1189 ( .A(A[643]), .B(n793), .Z(O[643]) );
  AND U1190 ( .A(S), .B(n794), .Z(n793) );
  XOR U1191 ( .A(B[643]), .B(A[643]), .Z(n794) );
  XOR U1192 ( .A(A[642]), .B(n795), .Z(O[642]) );
  AND U1193 ( .A(S), .B(n796), .Z(n795) );
  XOR U1194 ( .A(B[642]), .B(A[642]), .Z(n796) );
  XOR U1195 ( .A(A[641]), .B(n797), .Z(O[641]) );
  AND U1196 ( .A(S), .B(n798), .Z(n797) );
  XOR U1197 ( .A(B[641]), .B(A[641]), .Z(n798) );
  XOR U1198 ( .A(A[640]), .B(n799), .Z(O[640]) );
  AND U1199 ( .A(S), .B(n800), .Z(n799) );
  XOR U1200 ( .A(B[640]), .B(A[640]), .Z(n800) );
  XOR U1201 ( .A(A[63]), .B(n801), .Z(O[63]) );
  AND U1202 ( .A(S), .B(n802), .Z(n801) );
  XOR U1203 ( .A(B[63]), .B(A[63]), .Z(n802) );
  XOR U1204 ( .A(A[639]), .B(n803), .Z(O[639]) );
  AND U1205 ( .A(S), .B(n804), .Z(n803) );
  XOR U1206 ( .A(B[639]), .B(A[639]), .Z(n804) );
  XOR U1207 ( .A(A[638]), .B(n805), .Z(O[638]) );
  AND U1208 ( .A(S), .B(n806), .Z(n805) );
  XOR U1209 ( .A(B[638]), .B(A[638]), .Z(n806) );
  XOR U1210 ( .A(A[637]), .B(n807), .Z(O[637]) );
  AND U1211 ( .A(S), .B(n808), .Z(n807) );
  XOR U1212 ( .A(B[637]), .B(A[637]), .Z(n808) );
  XOR U1213 ( .A(A[636]), .B(n809), .Z(O[636]) );
  AND U1214 ( .A(S), .B(n810), .Z(n809) );
  XOR U1215 ( .A(B[636]), .B(A[636]), .Z(n810) );
  XOR U1216 ( .A(A[635]), .B(n811), .Z(O[635]) );
  AND U1217 ( .A(S), .B(n812), .Z(n811) );
  XOR U1218 ( .A(B[635]), .B(A[635]), .Z(n812) );
  XOR U1219 ( .A(A[634]), .B(n813), .Z(O[634]) );
  AND U1220 ( .A(S), .B(n814), .Z(n813) );
  XOR U1221 ( .A(B[634]), .B(A[634]), .Z(n814) );
  XOR U1222 ( .A(A[633]), .B(n815), .Z(O[633]) );
  AND U1223 ( .A(S), .B(n816), .Z(n815) );
  XOR U1224 ( .A(B[633]), .B(A[633]), .Z(n816) );
  XOR U1225 ( .A(A[632]), .B(n817), .Z(O[632]) );
  AND U1226 ( .A(S), .B(n818), .Z(n817) );
  XOR U1227 ( .A(B[632]), .B(A[632]), .Z(n818) );
  XOR U1228 ( .A(A[631]), .B(n819), .Z(O[631]) );
  AND U1229 ( .A(S), .B(n820), .Z(n819) );
  XOR U1230 ( .A(B[631]), .B(A[631]), .Z(n820) );
  XOR U1231 ( .A(A[630]), .B(n821), .Z(O[630]) );
  AND U1232 ( .A(S), .B(n822), .Z(n821) );
  XOR U1233 ( .A(B[630]), .B(A[630]), .Z(n822) );
  XOR U1234 ( .A(A[62]), .B(n823), .Z(O[62]) );
  AND U1235 ( .A(S), .B(n824), .Z(n823) );
  XOR U1236 ( .A(B[62]), .B(A[62]), .Z(n824) );
  XOR U1237 ( .A(A[629]), .B(n825), .Z(O[629]) );
  AND U1238 ( .A(S), .B(n826), .Z(n825) );
  XOR U1239 ( .A(B[629]), .B(A[629]), .Z(n826) );
  XOR U1240 ( .A(A[628]), .B(n827), .Z(O[628]) );
  AND U1241 ( .A(S), .B(n828), .Z(n827) );
  XOR U1242 ( .A(B[628]), .B(A[628]), .Z(n828) );
  XOR U1243 ( .A(A[627]), .B(n829), .Z(O[627]) );
  AND U1244 ( .A(S), .B(n830), .Z(n829) );
  XOR U1245 ( .A(B[627]), .B(A[627]), .Z(n830) );
  XOR U1246 ( .A(A[626]), .B(n831), .Z(O[626]) );
  AND U1247 ( .A(S), .B(n832), .Z(n831) );
  XOR U1248 ( .A(B[626]), .B(A[626]), .Z(n832) );
  XOR U1249 ( .A(A[625]), .B(n833), .Z(O[625]) );
  AND U1250 ( .A(S), .B(n834), .Z(n833) );
  XOR U1251 ( .A(B[625]), .B(A[625]), .Z(n834) );
  XOR U1252 ( .A(A[624]), .B(n835), .Z(O[624]) );
  AND U1253 ( .A(S), .B(n836), .Z(n835) );
  XOR U1254 ( .A(B[624]), .B(A[624]), .Z(n836) );
  XOR U1255 ( .A(A[623]), .B(n837), .Z(O[623]) );
  AND U1256 ( .A(S), .B(n838), .Z(n837) );
  XOR U1257 ( .A(B[623]), .B(A[623]), .Z(n838) );
  XOR U1258 ( .A(A[622]), .B(n839), .Z(O[622]) );
  AND U1259 ( .A(S), .B(n840), .Z(n839) );
  XOR U1260 ( .A(B[622]), .B(A[622]), .Z(n840) );
  XOR U1261 ( .A(A[621]), .B(n841), .Z(O[621]) );
  AND U1262 ( .A(S), .B(n842), .Z(n841) );
  XOR U1263 ( .A(B[621]), .B(A[621]), .Z(n842) );
  XOR U1264 ( .A(A[620]), .B(n843), .Z(O[620]) );
  AND U1265 ( .A(S), .B(n844), .Z(n843) );
  XOR U1266 ( .A(B[620]), .B(A[620]), .Z(n844) );
  XOR U1267 ( .A(A[61]), .B(n845), .Z(O[61]) );
  AND U1268 ( .A(S), .B(n846), .Z(n845) );
  XOR U1269 ( .A(B[61]), .B(A[61]), .Z(n846) );
  XOR U1270 ( .A(A[619]), .B(n847), .Z(O[619]) );
  AND U1271 ( .A(S), .B(n848), .Z(n847) );
  XOR U1272 ( .A(B[619]), .B(A[619]), .Z(n848) );
  XOR U1273 ( .A(A[618]), .B(n849), .Z(O[618]) );
  AND U1274 ( .A(S), .B(n850), .Z(n849) );
  XOR U1275 ( .A(B[618]), .B(A[618]), .Z(n850) );
  XOR U1276 ( .A(A[617]), .B(n851), .Z(O[617]) );
  AND U1277 ( .A(S), .B(n852), .Z(n851) );
  XOR U1278 ( .A(B[617]), .B(A[617]), .Z(n852) );
  XOR U1279 ( .A(A[616]), .B(n853), .Z(O[616]) );
  AND U1280 ( .A(S), .B(n854), .Z(n853) );
  XOR U1281 ( .A(B[616]), .B(A[616]), .Z(n854) );
  XOR U1282 ( .A(A[615]), .B(n855), .Z(O[615]) );
  AND U1283 ( .A(S), .B(n856), .Z(n855) );
  XOR U1284 ( .A(B[615]), .B(A[615]), .Z(n856) );
  XOR U1285 ( .A(A[614]), .B(n857), .Z(O[614]) );
  AND U1286 ( .A(S), .B(n858), .Z(n857) );
  XOR U1287 ( .A(B[614]), .B(A[614]), .Z(n858) );
  XOR U1288 ( .A(A[613]), .B(n859), .Z(O[613]) );
  AND U1289 ( .A(S), .B(n860), .Z(n859) );
  XOR U1290 ( .A(B[613]), .B(A[613]), .Z(n860) );
  XOR U1291 ( .A(A[612]), .B(n861), .Z(O[612]) );
  AND U1292 ( .A(S), .B(n862), .Z(n861) );
  XOR U1293 ( .A(B[612]), .B(A[612]), .Z(n862) );
  XOR U1294 ( .A(A[611]), .B(n863), .Z(O[611]) );
  AND U1295 ( .A(S), .B(n864), .Z(n863) );
  XOR U1296 ( .A(B[611]), .B(A[611]), .Z(n864) );
  XOR U1297 ( .A(A[610]), .B(n865), .Z(O[610]) );
  AND U1298 ( .A(S), .B(n866), .Z(n865) );
  XOR U1299 ( .A(B[610]), .B(A[610]), .Z(n866) );
  XOR U1300 ( .A(A[60]), .B(n867), .Z(O[60]) );
  AND U1301 ( .A(S), .B(n868), .Z(n867) );
  XOR U1302 ( .A(B[60]), .B(A[60]), .Z(n868) );
  XOR U1303 ( .A(A[609]), .B(n869), .Z(O[609]) );
  AND U1304 ( .A(S), .B(n870), .Z(n869) );
  XOR U1305 ( .A(B[609]), .B(A[609]), .Z(n870) );
  XOR U1306 ( .A(A[608]), .B(n871), .Z(O[608]) );
  AND U1307 ( .A(S), .B(n872), .Z(n871) );
  XOR U1308 ( .A(B[608]), .B(A[608]), .Z(n872) );
  XOR U1309 ( .A(A[607]), .B(n873), .Z(O[607]) );
  AND U1310 ( .A(S), .B(n874), .Z(n873) );
  XOR U1311 ( .A(B[607]), .B(A[607]), .Z(n874) );
  XOR U1312 ( .A(A[606]), .B(n875), .Z(O[606]) );
  AND U1313 ( .A(S), .B(n876), .Z(n875) );
  XOR U1314 ( .A(B[606]), .B(A[606]), .Z(n876) );
  XOR U1315 ( .A(A[605]), .B(n877), .Z(O[605]) );
  AND U1316 ( .A(S), .B(n878), .Z(n877) );
  XOR U1317 ( .A(B[605]), .B(A[605]), .Z(n878) );
  XOR U1318 ( .A(A[604]), .B(n879), .Z(O[604]) );
  AND U1319 ( .A(S), .B(n880), .Z(n879) );
  XOR U1320 ( .A(B[604]), .B(A[604]), .Z(n880) );
  XOR U1321 ( .A(A[603]), .B(n881), .Z(O[603]) );
  AND U1322 ( .A(S), .B(n882), .Z(n881) );
  XOR U1323 ( .A(B[603]), .B(A[603]), .Z(n882) );
  XOR U1324 ( .A(A[602]), .B(n883), .Z(O[602]) );
  AND U1325 ( .A(S), .B(n884), .Z(n883) );
  XOR U1326 ( .A(B[602]), .B(A[602]), .Z(n884) );
  XOR U1327 ( .A(A[601]), .B(n885), .Z(O[601]) );
  AND U1328 ( .A(S), .B(n886), .Z(n885) );
  XOR U1329 ( .A(B[601]), .B(A[601]), .Z(n886) );
  XOR U1330 ( .A(A[600]), .B(n887), .Z(O[600]) );
  AND U1331 ( .A(S), .B(n888), .Z(n887) );
  XOR U1332 ( .A(B[600]), .B(A[600]), .Z(n888) );
  XOR U1333 ( .A(A[5]), .B(n889), .Z(O[5]) );
  AND U1334 ( .A(S), .B(n890), .Z(n889) );
  XOR U1335 ( .A(B[5]), .B(A[5]), .Z(n890) );
  XOR U1336 ( .A(A[59]), .B(n891), .Z(O[59]) );
  AND U1337 ( .A(S), .B(n892), .Z(n891) );
  XOR U1338 ( .A(B[59]), .B(A[59]), .Z(n892) );
  XOR U1339 ( .A(A[599]), .B(n893), .Z(O[599]) );
  AND U1340 ( .A(S), .B(n894), .Z(n893) );
  XOR U1341 ( .A(B[599]), .B(A[599]), .Z(n894) );
  XOR U1342 ( .A(A[598]), .B(n895), .Z(O[598]) );
  AND U1343 ( .A(S), .B(n896), .Z(n895) );
  XOR U1344 ( .A(B[598]), .B(A[598]), .Z(n896) );
  XOR U1345 ( .A(A[597]), .B(n897), .Z(O[597]) );
  AND U1346 ( .A(S), .B(n898), .Z(n897) );
  XOR U1347 ( .A(B[597]), .B(A[597]), .Z(n898) );
  XOR U1348 ( .A(A[596]), .B(n899), .Z(O[596]) );
  AND U1349 ( .A(S), .B(n900), .Z(n899) );
  XOR U1350 ( .A(B[596]), .B(A[596]), .Z(n900) );
  XOR U1351 ( .A(A[595]), .B(n901), .Z(O[595]) );
  AND U1352 ( .A(S), .B(n902), .Z(n901) );
  XOR U1353 ( .A(B[595]), .B(A[595]), .Z(n902) );
  XOR U1354 ( .A(A[594]), .B(n903), .Z(O[594]) );
  AND U1355 ( .A(S), .B(n904), .Z(n903) );
  XOR U1356 ( .A(B[594]), .B(A[594]), .Z(n904) );
  XOR U1357 ( .A(A[593]), .B(n905), .Z(O[593]) );
  AND U1358 ( .A(S), .B(n906), .Z(n905) );
  XOR U1359 ( .A(B[593]), .B(A[593]), .Z(n906) );
  XOR U1360 ( .A(A[592]), .B(n907), .Z(O[592]) );
  AND U1361 ( .A(S), .B(n908), .Z(n907) );
  XOR U1362 ( .A(B[592]), .B(A[592]), .Z(n908) );
  XOR U1363 ( .A(A[591]), .B(n909), .Z(O[591]) );
  AND U1364 ( .A(S), .B(n910), .Z(n909) );
  XOR U1365 ( .A(B[591]), .B(A[591]), .Z(n910) );
  XOR U1366 ( .A(A[590]), .B(n911), .Z(O[590]) );
  AND U1367 ( .A(S), .B(n912), .Z(n911) );
  XOR U1368 ( .A(B[590]), .B(A[590]), .Z(n912) );
  XOR U1369 ( .A(A[58]), .B(n913), .Z(O[58]) );
  AND U1370 ( .A(S), .B(n914), .Z(n913) );
  XOR U1371 ( .A(B[58]), .B(A[58]), .Z(n914) );
  XOR U1372 ( .A(A[589]), .B(n915), .Z(O[589]) );
  AND U1373 ( .A(S), .B(n916), .Z(n915) );
  XOR U1374 ( .A(B[589]), .B(A[589]), .Z(n916) );
  XOR U1375 ( .A(A[588]), .B(n917), .Z(O[588]) );
  AND U1376 ( .A(S), .B(n918), .Z(n917) );
  XOR U1377 ( .A(B[588]), .B(A[588]), .Z(n918) );
  XOR U1378 ( .A(A[587]), .B(n919), .Z(O[587]) );
  AND U1379 ( .A(S), .B(n920), .Z(n919) );
  XOR U1380 ( .A(B[587]), .B(A[587]), .Z(n920) );
  XOR U1381 ( .A(A[586]), .B(n921), .Z(O[586]) );
  AND U1382 ( .A(S), .B(n922), .Z(n921) );
  XOR U1383 ( .A(B[586]), .B(A[586]), .Z(n922) );
  XOR U1384 ( .A(A[585]), .B(n923), .Z(O[585]) );
  AND U1385 ( .A(S), .B(n924), .Z(n923) );
  XOR U1386 ( .A(B[585]), .B(A[585]), .Z(n924) );
  XOR U1387 ( .A(A[584]), .B(n925), .Z(O[584]) );
  AND U1388 ( .A(S), .B(n926), .Z(n925) );
  XOR U1389 ( .A(B[584]), .B(A[584]), .Z(n926) );
  XOR U1390 ( .A(A[583]), .B(n927), .Z(O[583]) );
  AND U1391 ( .A(S), .B(n928), .Z(n927) );
  XOR U1392 ( .A(B[583]), .B(A[583]), .Z(n928) );
  XOR U1393 ( .A(A[582]), .B(n929), .Z(O[582]) );
  AND U1394 ( .A(S), .B(n930), .Z(n929) );
  XOR U1395 ( .A(B[582]), .B(A[582]), .Z(n930) );
  XOR U1396 ( .A(A[581]), .B(n931), .Z(O[581]) );
  AND U1397 ( .A(S), .B(n932), .Z(n931) );
  XOR U1398 ( .A(B[581]), .B(A[581]), .Z(n932) );
  XOR U1399 ( .A(A[580]), .B(n933), .Z(O[580]) );
  AND U1400 ( .A(S), .B(n934), .Z(n933) );
  XOR U1401 ( .A(B[580]), .B(A[580]), .Z(n934) );
  XOR U1402 ( .A(A[57]), .B(n935), .Z(O[57]) );
  AND U1403 ( .A(S), .B(n936), .Z(n935) );
  XOR U1404 ( .A(B[57]), .B(A[57]), .Z(n936) );
  XOR U1405 ( .A(A[579]), .B(n937), .Z(O[579]) );
  AND U1406 ( .A(S), .B(n938), .Z(n937) );
  XOR U1407 ( .A(B[579]), .B(A[579]), .Z(n938) );
  XOR U1408 ( .A(A[578]), .B(n939), .Z(O[578]) );
  AND U1409 ( .A(S), .B(n940), .Z(n939) );
  XOR U1410 ( .A(B[578]), .B(A[578]), .Z(n940) );
  XOR U1411 ( .A(A[577]), .B(n941), .Z(O[577]) );
  AND U1412 ( .A(S), .B(n942), .Z(n941) );
  XOR U1413 ( .A(B[577]), .B(A[577]), .Z(n942) );
  XOR U1414 ( .A(A[576]), .B(n943), .Z(O[576]) );
  AND U1415 ( .A(S), .B(n944), .Z(n943) );
  XOR U1416 ( .A(B[576]), .B(A[576]), .Z(n944) );
  XOR U1417 ( .A(A[575]), .B(n945), .Z(O[575]) );
  AND U1418 ( .A(S), .B(n946), .Z(n945) );
  XOR U1419 ( .A(B[575]), .B(A[575]), .Z(n946) );
  XOR U1420 ( .A(A[574]), .B(n947), .Z(O[574]) );
  AND U1421 ( .A(S), .B(n948), .Z(n947) );
  XOR U1422 ( .A(B[574]), .B(A[574]), .Z(n948) );
  XOR U1423 ( .A(A[573]), .B(n949), .Z(O[573]) );
  AND U1424 ( .A(S), .B(n950), .Z(n949) );
  XOR U1425 ( .A(B[573]), .B(A[573]), .Z(n950) );
  XOR U1426 ( .A(A[572]), .B(n951), .Z(O[572]) );
  AND U1427 ( .A(S), .B(n952), .Z(n951) );
  XOR U1428 ( .A(B[572]), .B(A[572]), .Z(n952) );
  XOR U1429 ( .A(A[571]), .B(n953), .Z(O[571]) );
  AND U1430 ( .A(S), .B(n954), .Z(n953) );
  XOR U1431 ( .A(B[571]), .B(A[571]), .Z(n954) );
  XOR U1432 ( .A(A[570]), .B(n955), .Z(O[570]) );
  AND U1433 ( .A(S), .B(n956), .Z(n955) );
  XOR U1434 ( .A(B[570]), .B(A[570]), .Z(n956) );
  XOR U1435 ( .A(A[56]), .B(n957), .Z(O[56]) );
  AND U1436 ( .A(S), .B(n958), .Z(n957) );
  XOR U1437 ( .A(B[56]), .B(A[56]), .Z(n958) );
  XOR U1438 ( .A(A[569]), .B(n959), .Z(O[569]) );
  AND U1439 ( .A(S), .B(n960), .Z(n959) );
  XOR U1440 ( .A(B[569]), .B(A[569]), .Z(n960) );
  XOR U1441 ( .A(A[568]), .B(n961), .Z(O[568]) );
  AND U1442 ( .A(S), .B(n962), .Z(n961) );
  XOR U1443 ( .A(B[568]), .B(A[568]), .Z(n962) );
  XOR U1444 ( .A(A[567]), .B(n963), .Z(O[567]) );
  AND U1445 ( .A(S), .B(n964), .Z(n963) );
  XOR U1446 ( .A(B[567]), .B(A[567]), .Z(n964) );
  XOR U1447 ( .A(A[566]), .B(n965), .Z(O[566]) );
  AND U1448 ( .A(S), .B(n966), .Z(n965) );
  XOR U1449 ( .A(B[566]), .B(A[566]), .Z(n966) );
  XOR U1450 ( .A(A[565]), .B(n967), .Z(O[565]) );
  AND U1451 ( .A(S), .B(n968), .Z(n967) );
  XOR U1452 ( .A(B[565]), .B(A[565]), .Z(n968) );
  XOR U1453 ( .A(A[564]), .B(n969), .Z(O[564]) );
  AND U1454 ( .A(S), .B(n970), .Z(n969) );
  XOR U1455 ( .A(B[564]), .B(A[564]), .Z(n970) );
  XOR U1456 ( .A(A[563]), .B(n971), .Z(O[563]) );
  AND U1457 ( .A(S), .B(n972), .Z(n971) );
  XOR U1458 ( .A(B[563]), .B(A[563]), .Z(n972) );
  XOR U1459 ( .A(A[562]), .B(n973), .Z(O[562]) );
  AND U1460 ( .A(S), .B(n974), .Z(n973) );
  XOR U1461 ( .A(B[562]), .B(A[562]), .Z(n974) );
  XOR U1462 ( .A(A[561]), .B(n975), .Z(O[561]) );
  AND U1463 ( .A(S), .B(n976), .Z(n975) );
  XOR U1464 ( .A(B[561]), .B(A[561]), .Z(n976) );
  XOR U1465 ( .A(A[560]), .B(n977), .Z(O[560]) );
  AND U1466 ( .A(S), .B(n978), .Z(n977) );
  XOR U1467 ( .A(B[560]), .B(A[560]), .Z(n978) );
  XOR U1468 ( .A(A[55]), .B(n979), .Z(O[55]) );
  AND U1469 ( .A(S), .B(n980), .Z(n979) );
  XOR U1470 ( .A(B[55]), .B(A[55]), .Z(n980) );
  XOR U1471 ( .A(A[559]), .B(n981), .Z(O[559]) );
  AND U1472 ( .A(S), .B(n982), .Z(n981) );
  XOR U1473 ( .A(B[559]), .B(A[559]), .Z(n982) );
  XOR U1474 ( .A(A[558]), .B(n983), .Z(O[558]) );
  AND U1475 ( .A(S), .B(n984), .Z(n983) );
  XOR U1476 ( .A(B[558]), .B(A[558]), .Z(n984) );
  XOR U1477 ( .A(A[557]), .B(n985), .Z(O[557]) );
  AND U1478 ( .A(S), .B(n986), .Z(n985) );
  XOR U1479 ( .A(B[557]), .B(A[557]), .Z(n986) );
  XOR U1480 ( .A(A[556]), .B(n987), .Z(O[556]) );
  AND U1481 ( .A(S), .B(n988), .Z(n987) );
  XOR U1482 ( .A(B[556]), .B(A[556]), .Z(n988) );
  XOR U1483 ( .A(A[555]), .B(n989), .Z(O[555]) );
  AND U1484 ( .A(S), .B(n990), .Z(n989) );
  XOR U1485 ( .A(B[555]), .B(A[555]), .Z(n990) );
  XOR U1486 ( .A(A[554]), .B(n991), .Z(O[554]) );
  AND U1487 ( .A(S), .B(n992), .Z(n991) );
  XOR U1488 ( .A(B[554]), .B(A[554]), .Z(n992) );
  XOR U1489 ( .A(A[553]), .B(n993), .Z(O[553]) );
  AND U1490 ( .A(S), .B(n994), .Z(n993) );
  XOR U1491 ( .A(B[553]), .B(A[553]), .Z(n994) );
  XOR U1492 ( .A(A[552]), .B(n995), .Z(O[552]) );
  AND U1493 ( .A(S), .B(n996), .Z(n995) );
  XOR U1494 ( .A(B[552]), .B(A[552]), .Z(n996) );
  XOR U1495 ( .A(A[551]), .B(n997), .Z(O[551]) );
  AND U1496 ( .A(S), .B(n998), .Z(n997) );
  XOR U1497 ( .A(B[551]), .B(A[551]), .Z(n998) );
  XOR U1498 ( .A(A[550]), .B(n999), .Z(O[550]) );
  AND U1499 ( .A(S), .B(n1000), .Z(n999) );
  XOR U1500 ( .A(B[550]), .B(A[550]), .Z(n1000) );
  XOR U1501 ( .A(A[54]), .B(n1001), .Z(O[54]) );
  AND U1502 ( .A(S), .B(n1002), .Z(n1001) );
  XOR U1503 ( .A(B[54]), .B(A[54]), .Z(n1002) );
  XOR U1504 ( .A(A[549]), .B(n1003), .Z(O[549]) );
  AND U1505 ( .A(S), .B(n1004), .Z(n1003) );
  XOR U1506 ( .A(B[549]), .B(A[549]), .Z(n1004) );
  XOR U1507 ( .A(A[548]), .B(n1005), .Z(O[548]) );
  AND U1508 ( .A(S), .B(n1006), .Z(n1005) );
  XOR U1509 ( .A(B[548]), .B(A[548]), .Z(n1006) );
  XOR U1510 ( .A(A[547]), .B(n1007), .Z(O[547]) );
  AND U1511 ( .A(S), .B(n1008), .Z(n1007) );
  XOR U1512 ( .A(B[547]), .B(A[547]), .Z(n1008) );
  XOR U1513 ( .A(A[546]), .B(n1009), .Z(O[546]) );
  AND U1514 ( .A(S), .B(n1010), .Z(n1009) );
  XOR U1515 ( .A(B[546]), .B(A[546]), .Z(n1010) );
  XOR U1516 ( .A(A[545]), .B(n1011), .Z(O[545]) );
  AND U1517 ( .A(S), .B(n1012), .Z(n1011) );
  XOR U1518 ( .A(B[545]), .B(A[545]), .Z(n1012) );
  XOR U1519 ( .A(A[544]), .B(n1013), .Z(O[544]) );
  AND U1520 ( .A(S), .B(n1014), .Z(n1013) );
  XOR U1521 ( .A(B[544]), .B(A[544]), .Z(n1014) );
  XOR U1522 ( .A(A[543]), .B(n1015), .Z(O[543]) );
  AND U1523 ( .A(S), .B(n1016), .Z(n1015) );
  XOR U1524 ( .A(B[543]), .B(A[543]), .Z(n1016) );
  XOR U1525 ( .A(A[542]), .B(n1017), .Z(O[542]) );
  AND U1526 ( .A(S), .B(n1018), .Z(n1017) );
  XOR U1527 ( .A(B[542]), .B(A[542]), .Z(n1018) );
  XOR U1528 ( .A(A[541]), .B(n1019), .Z(O[541]) );
  AND U1529 ( .A(S), .B(n1020), .Z(n1019) );
  XOR U1530 ( .A(B[541]), .B(A[541]), .Z(n1020) );
  XOR U1531 ( .A(A[540]), .B(n1021), .Z(O[540]) );
  AND U1532 ( .A(S), .B(n1022), .Z(n1021) );
  XOR U1533 ( .A(B[540]), .B(A[540]), .Z(n1022) );
  XOR U1534 ( .A(A[53]), .B(n1023), .Z(O[53]) );
  AND U1535 ( .A(S), .B(n1024), .Z(n1023) );
  XOR U1536 ( .A(B[53]), .B(A[53]), .Z(n1024) );
  XOR U1537 ( .A(A[539]), .B(n1025), .Z(O[539]) );
  AND U1538 ( .A(S), .B(n1026), .Z(n1025) );
  XOR U1539 ( .A(B[539]), .B(A[539]), .Z(n1026) );
  XOR U1540 ( .A(A[538]), .B(n1027), .Z(O[538]) );
  AND U1541 ( .A(S), .B(n1028), .Z(n1027) );
  XOR U1542 ( .A(B[538]), .B(A[538]), .Z(n1028) );
  XOR U1543 ( .A(A[537]), .B(n1029), .Z(O[537]) );
  AND U1544 ( .A(S), .B(n1030), .Z(n1029) );
  XOR U1545 ( .A(B[537]), .B(A[537]), .Z(n1030) );
  XOR U1546 ( .A(A[536]), .B(n1031), .Z(O[536]) );
  AND U1547 ( .A(S), .B(n1032), .Z(n1031) );
  XOR U1548 ( .A(B[536]), .B(A[536]), .Z(n1032) );
  XOR U1549 ( .A(A[535]), .B(n1033), .Z(O[535]) );
  AND U1550 ( .A(S), .B(n1034), .Z(n1033) );
  XOR U1551 ( .A(B[535]), .B(A[535]), .Z(n1034) );
  XOR U1552 ( .A(A[534]), .B(n1035), .Z(O[534]) );
  AND U1553 ( .A(S), .B(n1036), .Z(n1035) );
  XOR U1554 ( .A(B[534]), .B(A[534]), .Z(n1036) );
  XOR U1555 ( .A(A[533]), .B(n1037), .Z(O[533]) );
  AND U1556 ( .A(S), .B(n1038), .Z(n1037) );
  XOR U1557 ( .A(B[533]), .B(A[533]), .Z(n1038) );
  XOR U1558 ( .A(A[532]), .B(n1039), .Z(O[532]) );
  AND U1559 ( .A(S), .B(n1040), .Z(n1039) );
  XOR U1560 ( .A(B[532]), .B(A[532]), .Z(n1040) );
  XOR U1561 ( .A(A[531]), .B(n1041), .Z(O[531]) );
  AND U1562 ( .A(S), .B(n1042), .Z(n1041) );
  XOR U1563 ( .A(B[531]), .B(A[531]), .Z(n1042) );
  XOR U1564 ( .A(A[530]), .B(n1043), .Z(O[530]) );
  AND U1565 ( .A(S), .B(n1044), .Z(n1043) );
  XOR U1566 ( .A(B[530]), .B(A[530]), .Z(n1044) );
  XOR U1567 ( .A(A[52]), .B(n1045), .Z(O[52]) );
  AND U1568 ( .A(S), .B(n1046), .Z(n1045) );
  XOR U1569 ( .A(B[52]), .B(A[52]), .Z(n1046) );
  XOR U1570 ( .A(A[529]), .B(n1047), .Z(O[529]) );
  AND U1571 ( .A(S), .B(n1048), .Z(n1047) );
  XOR U1572 ( .A(B[529]), .B(A[529]), .Z(n1048) );
  XOR U1573 ( .A(A[528]), .B(n1049), .Z(O[528]) );
  AND U1574 ( .A(S), .B(n1050), .Z(n1049) );
  XOR U1575 ( .A(B[528]), .B(A[528]), .Z(n1050) );
  XOR U1576 ( .A(A[527]), .B(n1051), .Z(O[527]) );
  AND U1577 ( .A(S), .B(n1052), .Z(n1051) );
  XOR U1578 ( .A(B[527]), .B(A[527]), .Z(n1052) );
  XOR U1579 ( .A(A[526]), .B(n1053), .Z(O[526]) );
  AND U1580 ( .A(S), .B(n1054), .Z(n1053) );
  XOR U1581 ( .A(B[526]), .B(A[526]), .Z(n1054) );
  XOR U1582 ( .A(A[525]), .B(n1055), .Z(O[525]) );
  AND U1583 ( .A(S), .B(n1056), .Z(n1055) );
  XOR U1584 ( .A(B[525]), .B(A[525]), .Z(n1056) );
  XOR U1585 ( .A(A[524]), .B(n1057), .Z(O[524]) );
  AND U1586 ( .A(S), .B(n1058), .Z(n1057) );
  XOR U1587 ( .A(B[524]), .B(A[524]), .Z(n1058) );
  XOR U1588 ( .A(A[523]), .B(n1059), .Z(O[523]) );
  AND U1589 ( .A(S), .B(n1060), .Z(n1059) );
  XOR U1590 ( .A(B[523]), .B(A[523]), .Z(n1060) );
  XOR U1591 ( .A(A[522]), .B(n1061), .Z(O[522]) );
  AND U1592 ( .A(S), .B(n1062), .Z(n1061) );
  XOR U1593 ( .A(B[522]), .B(A[522]), .Z(n1062) );
  XOR U1594 ( .A(A[521]), .B(n1063), .Z(O[521]) );
  AND U1595 ( .A(S), .B(n1064), .Z(n1063) );
  XOR U1596 ( .A(B[521]), .B(A[521]), .Z(n1064) );
  XOR U1597 ( .A(A[520]), .B(n1065), .Z(O[520]) );
  AND U1598 ( .A(S), .B(n1066), .Z(n1065) );
  XOR U1599 ( .A(B[520]), .B(A[520]), .Z(n1066) );
  XOR U1600 ( .A(A[51]), .B(n1067), .Z(O[51]) );
  AND U1601 ( .A(S), .B(n1068), .Z(n1067) );
  XOR U1602 ( .A(B[51]), .B(A[51]), .Z(n1068) );
  XOR U1603 ( .A(A[519]), .B(n1069), .Z(O[519]) );
  AND U1604 ( .A(S), .B(n1070), .Z(n1069) );
  XOR U1605 ( .A(B[519]), .B(A[519]), .Z(n1070) );
  XOR U1606 ( .A(A[518]), .B(n1071), .Z(O[518]) );
  AND U1607 ( .A(S), .B(n1072), .Z(n1071) );
  XOR U1608 ( .A(B[518]), .B(A[518]), .Z(n1072) );
  XOR U1609 ( .A(A[517]), .B(n1073), .Z(O[517]) );
  AND U1610 ( .A(S), .B(n1074), .Z(n1073) );
  XOR U1611 ( .A(B[517]), .B(A[517]), .Z(n1074) );
  XOR U1612 ( .A(A[516]), .B(n1075), .Z(O[516]) );
  AND U1613 ( .A(S), .B(n1076), .Z(n1075) );
  XOR U1614 ( .A(B[516]), .B(A[516]), .Z(n1076) );
  XOR U1615 ( .A(A[515]), .B(n1077), .Z(O[515]) );
  AND U1616 ( .A(S), .B(n1078), .Z(n1077) );
  XOR U1617 ( .A(B[515]), .B(A[515]), .Z(n1078) );
  XOR U1618 ( .A(A[514]), .B(n1079), .Z(O[514]) );
  AND U1619 ( .A(S), .B(n1080), .Z(n1079) );
  XOR U1620 ( .A(B[514]), .B(A[514]), .Z(n1080) );
  XOR U1621 ( .A(A[513]), .B(n1081), .Z(O[513]) );
  AND U1622 ( .A(S), .B(n1082), .Z(n1081) );
  XOR U1623 ( .A(B[513]), .B(A[513]), .Z(n1082) );
  XOR U1624 ( .A(A[512]), .B(n1083), .Z(O[512]) );
  AND U1625 ( .A(S), .B(n1084), .Z(n1083) );
  XOR U1626 ( .A(B[512]), .B(A[512]), .Z(n1084) );
  XOR U1627 ( .A(A[511]), .B(n1085), .Z(O[511]) );
  AND U1628 ( .A(S), .B(n1086), .Z(n1085) );
  XOR U1629 ( .A(B[511]), .B(A[511]), .Z(n1086) );
  XOR U1630 ( .A(A[510]), .B(n1087), .Z(O[510]) );
  AND U1631 ( .A(S), .B(n1088), .Z(n1087) );
  XOR U1632 ( .A(B[510]), .B(A[510]), .Z(n1088) );
  XOR U1633 ( .A(A[50]), .B(n1089), .Z(O[50]) );
  AND U1634 ( .A(S), .B(n1090), .Z(n1089) );
  XOR U1635 ( .A(B[50]), .B(A[50]), .Z(n1090) );
  XOR U1636 ( .A(A[509]), .B(n1091), .Z(O[509]) );
  AND U1637 ( .A(S), .B(n1092), .Z(n1091) );
  XOR U1638 ( .A(B[509]), .B(A[509]), .Z(n1092) );
  XOR U1639 ( .A(A[508]), .B(n1093), .Z(O[508]) );
  AND U1640 ( .A(S), .B(n1094), .Z(n1093) );
  XOR U1641 ( .A(B[508]), .B(A[508]), .Z(n1094) );
  XOR U1642 ( .A(A[507]), .B(n1095), .Z(O[507]) );
  AND U1643 ( .A(S), .B(n1096), .Z(n1095) );
  XOR U1644 ( .A(B[507]), .B(A[507]), .Z(n1096) );
  XOR U1645 ( .A(A[506]), .B(n1097), .Z(O[506]) );
  AND U1646 ( .A(S), .B(n1098), .Z(n1097) );
  XOR U1647 ( .A(B[506]), .B(A[506]), .Z(n1098) );
  XOR U1648 ( .A(A[505]), .B(n1099), .Z(O[505]) );
  AND U1649 ( .A(S), .B(n1100), .Z(n1099) );
  XOR U1650 ( .A(B[505]), .B(A[505]), .Z(n1100) );
  XOR U1651 ( .A(A[504]), .B(n1101), .Z(O[504]) );
  AND U1652 ( .A(S), .B(n1102), .Z(n1101) );
  XOR U1653 ( .A(B[504]), .B(A[504]), .Z(n1102) );
  XOR U1654 ( .A(A[503]), .B(n1103), .Z(O[503]) );
  AND U1655 ( .A(S), .B(n1104), .Z(n1103) );
  XOR U1656 ( .A(B[503]), .B(A[503]), .Z(n1104) );
  XOR U1657 ( .A(A[502]), .B(n1105), .Z(O[502]) );
  AND U1658 ( .A(S), .B(n1106), .Z(n1105) );
  XOR U1659 ( .A(B[502]), .B(A[502]), .Z(n1106) );
  XOR U1660 ( .A(A[501]), .B(n1107), .Z(O[501]) );
  AND U1661 ( .A(S), .B(n1108), .Z(n1107) );
  XOR U1662 ( .A(B[501]), .B(A[501]), .Z(n1108) );
  XOR U1663 ( .A(A[500]), .B(n1109), .Z(O[500]) );
  AND U1664 ( .A(S), .B(n1110), .Z(n1109) );
  XOR U1665 ( .A(B[500]), .B(A[500]), .Z(n1110) );
  XOR U1666 ( .A(A[4]), .B(n1111), .Z(O[4]) );
  AND U1667 ( .A(S), .B(n1112), .Z(n1111) );
  XOR U1668 ( .A(B[4]), .B(A[4]), .Z(n1112) );
  XOR U1669 ( .A(A[49]), .B(n1113), .Z(O[49]) );
  AND U1670 ( .A(S), .B(n1114), .Z(n1113) );
  XOR U1671 ( .A(B[49]), .B(A[49]), .Z(n1114) );
  XOR U1672 ( .A(A[499]), .B(n1115), .Z(O[499]) );
  AND U1673 ( .A(S), .B(n1116), .Z(n1115) );
  XOR U1674 ( .A(B[499]), .B(A[499]), .Z(n1116) );
  XOR U1675 ( .A(A[498]), .B(n1117), .Z(O[498]) );
  AND U1676 ( .A(S), .B(n1118), .Z(n1117) );
  XOR U1677 ( .A(B[498]), .B(A[498]), .Z(n1118) );
  XOR U1678 ( .A(A[497]), .B(n1119), .Z(O[497]) );
  AND U1679 ( .A(S), .B(n1120), .Z(n1119) );
  XOR U1680 ( .A(B[497]), .B(A[497]), .Z(n1120) );
  XOR U1681 ( .A(A[496]), .B(n1121), .Z(O[496]) );
  AND U1682 ( .A(S), .B(n1122), .Z(n1121) );
  XOR U1683 ( .A(B[496]), .B(A[496]), .Z(n1122) );
  XOR U1684 ( .A(A[495]), .B(n1123), .Z(O[495]) );
  AND U1685 ( .A(S), .B(n1124), .Z(n1123) );
  XOR U1686 ( .A(B[495]), .B(A[495]), .Z(n1124) );
  XOR U1687 ( .A(A[494]), .B(n1125), .Z(O[494]) );
  AND U1688 ( .A(S), .B(n1126), .Z(n1125) );
  XOR U1689 ( .A(B[494]), .B(A[494]), .Z(n1126) );
  XOR U1690 ( .A(A[493]), .B(n1127), .Z(O[493]) );
  AND U1691 ( .A(S), .B(n1128), .Z(n1127) );
  XOR U1692 ( .A(B[493]), .B(A[493]), .Z(n1128) );
  XOR U1693 ( .A(A[492]), .B(n1129), .Z(O[492]) );
  AND U1694 ( .A(S), .B(n1130), .Z(n1129) );
  XOR U1695 ( .A(B[492]), .B(A[492]), .Z(n1130) );
  XOR U1696 ( .A(A[491]), .B(n1131), .Z(O[491]) );
  AND U1697 ( .A(S), .B(n1132), .Z(n1131) );
  XOR U1698 ( .A(B[491]), .B(A[491]), .Z(n1132) );
  XOR U1699 ( .A(A[490]), .B(n1133), .Z(O[490]) );
  AND U1700 ( .A(S), .B(n1134), .Z(n1133) );
  XOR U1701 ( .A(B[490]), .B(A[490]), .Z(n1134) );
  XOR U1702 ( .A(A[48]), .B(n1135), .Z(O[48]) );
  AND U1703 ( .A(S), .B(n1136), .Z(n1135) );
  XOR U1704 ( .A(B[48]), .B(A[48]), .Z(n1136) );
  XOR U1705 ( .A(A[489]), .B(n1137), .Z(O[489]) );
  AND U1706 ( .A(S), .B(n1138), .Z(n1137) );
  XOR U1707 ( .A(B[489]), .B(A[489]), .Z(n1138) );
  XOR U1708 ( .A(A[488]), .B(n1139), .Z(O[488]) );
  AND U1709 ( .A(S), .B(n1140), .Z(n1139) );
  XOR U1710 ( .A(B[488]), .B(A[488]), .Z(n1140) );
  XOR U1711 ( .A(A[487]), .B(n1141), .Z(O[487]) );
  AND U1712 ( .A(S), .B(n1142), .Z(n1141) );
  XOR U1713 ( .A(B[487]), .B(A[487]), .Z(n1142) );
  XOR U1714 ( .A(A[486]), .B(n1143), .Z(O[486]) );
  AND U1715 ( .A(S), .B(n1144), .Z(n1143) );
  XOR U1716 ( .A(B[486]), .B(A[486]), .Z(n1144) );
  XOR U1717 ( .A(A[485]), .B(n1145), .Z(O[485]) );
  AND U1718 ( .A(S), .B(n1146), .Z(n1145) );
  XOR U1719 ( .A(B[485]), .B(A[485]), .Z(n1146) );
  XOR U1720 ( .A(A[484]), .B(n1147), .Z(O[484]) );
  AND U1721 ( .A(S), .B(n1148), .Z(n1147) );
  XOR U1722 ( .A(B[484]), .B(A[484]), .Z(n1148) );
  XOR U1723 ( .A(A[483]), .B(n1149), .Z(O[483]) );
  AND U1724 ( .A(S), .B(n1150), .Z(n1149) );
  XOR U1725 ( .A(B[483]), .B(A[483]), .Z(n1150) );
  XOR U1726 ( .A(A[482]), .B(n1151), .Z(O[482]) );
  AND U1727 ( .A(S), .B(n1152), .Z(n1151) );
  XOR U1728 ( .A(B[482]), .B(A[482]), .Z(n1152) );
  XOR U1729 ( .A(A[481]), .B(n1153), .Z(O[481]) );
  AND U1730 ( .A(S), .B(n1154), .Z(n1153) );
  XOR U1731 ( .A(B[481]), .B(A[481]), .Z(n1154) );
  XOR U1732 ( .A(A[480]), .B(n1155), .Z(O[480]) );
  AND U1733 ( .A(S), .B(n1156), .Z(n1155) );
  XOR U1734 ( .A(B[480]), .B(A[480]), .Z(n1156) );
  XOR U1735 ( .A(A[47]), .B(n1157), .Z(O[47]) );
  AND U1736 ( .A(S), .B(n1158), .Z(n1157) );
  XOR U1737 ( .A(B[47]), .B(A[47]), .Z(n1158) );
  XOR U1738 ( .A(A[479]), .B(n1159), .Z(O[479]) );
  AND U1739 ( .A(S), .B(n1160), .Z(n1159) );
  XOR U1740 ( .A(B[479]), .B(A[479]), .Z(n1160) );
  XOR U1741 ( .A(A[478]), .B(n1161), .Z(O[478]) );
  AND U1742 ( .A(S), .B(n1162), .Z(n1161) );
  XOR U1743 ( .A(B[478]), .B(A[478]), .Z(n1162) );
  XOR U1744 ( .A(A[477]), .B(n1163), .Z(O[477]) );
  AND U1745 ( .A(S), .B(n1164), .Z(n1163) );
  XOR U1746 ( .A(B[477]), .B(A[477]), .Z(n1164) );
  XOR U1747 ( .A(A[476]), .B(n1165), .Z(O[476]) );
  AND U1748 ( .A(S), .B(n1166), .Z(n1165) );
  XOR U1749 ( .A(B[476]), .B(A[476]), .Z(n1166) );
  XOR U1750 ( .A(A[475]), .B(n1167), .Z(O[475]) );
  AND U1751 ( .A(S), .B(n1168), .Z(n1167) );
  XOR U1752 ( .A(B[475]), .B(A[475]), .Z(n1168) );
  XOR U1753 ( .A(A[474]), .B(n1169), .Z(O[474]) );
  AND U1754 ( .A(S), .B(n1170), .Z(n1169) );
  XOR U1755 ( .A(B[474]), .B(A[474]), .Z(n1170) );
  XOR U1756 ( .A(A[473]), .B(n1171), .Z(O[473]) );
  AND U1757 ( .A(S), .B(n1172), .Z(n1171) );
  XOR U1758 ( .A(B[473]), .B(A[473]), .Z(n1172) );
  XOR U1759 ( .A(A[472]), .B(n1173), .Z(O[472]) );
  AND U1760 ( .A(S), .B(n1174), .Z(n1173) );
  XOR U1761 ( .A(B[472]), .B(A[472]), .Z(n1174) );
  XOR U1762 ( .A(A[471]), .B(n1175), .Z(O[471]) );
  AND U1763 ( .A(S), .B(n1176), .Z(n1175) );
  XOR U1764 ( .A(B[471]), .B(A[471]), .Z(n1176) );
  XOR U1765 ( .A(A[470]), .B(n1177), .Z(O[470]) );
  AND U1766 ( .A(S), .B(n1178), .Z(n1177) );
  XOR U1767 ( .A(B[470]), .B(A[470]), .Z(n1178) );
  XOR U1768 ( .A(A[46]), .B(n1179), .Z(O[46]) );
  AND U1769 ( .A(S), .B(n1180), .Z(n1179) );
  XOR U1770 ( .A(B[46]), .B(A[46]), .Z(n1180) );
  XOR U1771 ( .A(A[469]), .B(n1181), .Z(O[469]) );
  AND U1772 ( .A(S), .B(n1182), .Z(n1181) );
  XOR U1773 ( .A(B[469]), .B(A[469]), .Z(n1182) );
  XOR U1774 ( .A(A[468]), .B(n1183), .Z(O[468]) );
  AND U1775 ( .A(S), .B(n1184), .Z(n1183) );
  XOR U1776 ( .A(B[468]), .B(A[468]), .Z(n1184) );
  XOR U1777 ( .A(A[467]), .B(n1185), .Z(O[467]) );
  AND U1778 ( .A(S), .B(n1186), .Z(n1185) );
  XOR U1779 ( .A(B[467]), .B(A[467]), .Z(n1186) );
  XOR U1780 ( .A(A[466]), .B(n1187), .Z(O[466]) );
  AND U1781 ( .A(S), .B(n1188), .Z(n1187) );
  XOR U1782 ( .A(B[466]), .B(A[466]), .Z(n1188) );
  XOR U1783 ( .A(A[465]), .B(n1189), .Z(O[465]) );
  AND U1784 ( .A(S), .B(n1190), .Z(n1189) );
  XOR U1785 ( .A(B[465]), .B(A[465]), .Z(n1190) );
  XOR U1786 ( .A(A[464]), .B(n1191), .Z(O[464]) );
  AND U1787 ( .A(S), .B(n1192), .Z(n1191) );
  XOR U1788 ( .A(B[464]), .B(A[464]), .Z(n1192) );
  XOR U1789 ( .A(A[463]), .B(n1193), .Z(O[463]) );
  AND U1790 ( .A(S), .B(n1194), .Z(n1193) );
  XOR U1791 ( .A(B[463]), .B(A[463]), .Z(n1194) );
  XOR U1792 ( .A(A[462]), .B(n1195), .Z(O[462]) );
  AND U1793 ( .A(S), .B(n1196), .Z(n1195) );
  XOR U1794 ( .A(B[462]), .B(A[462]), .Z(n1196) );
  XOR U1795 ( .A(A[461]), .B(n1197), .Z(O[461]) );
  AND U1796 ( .A(S), .B(n1198), .Z(n1197) );
  XOR U1797 ( .A(B[461]), .B(A[461]), .Z(n1198) );
  XOR U1798 ( .A(A[460]), .B(n1199), .Z(O[460]) );
  AND U1799 ( .A(S), .B(n1200), .Z(n1199) );
  XOR U1800 ( .A(B[460]), .B(A[460]), .Z(n1200) );
  XOR U1801 ( .A(A[45]), .B(n1201), .Z(O[45]) );
  AND U1802 ( .A(S), .B(n1202), .Z(n1201) );
  XOR U1803 ( .A(B[45]), .B(A[45]), .Z(n1202) );
  XOR U1804 ( .A(A[459]), .B(n1203), .Z(O[459]) );
  AND U1805 ( .A(S), .B(n1204), .Z(n1203) );
  XOR U1806 ( .A(B[459]), .B(A[459]), .Z(n1204) );
  XOR U1807 ( .A(A[458]), .B(n1205), .Z(O[458]) );
  AND U1808 ( .A(S), .B(n1206), .Z(n1205) );
  XOR U1809 ( .A(B[458]), .B(A[458]), .Z(n1206) );
  XOR U1810 ( .A(A[457]), .B(n1207), .Z(O[457]) );
  AND U1811 ( .A(S), .B(n1208), .Z(n1207) );
  XOR U1812 ( .A(B[457]), .B(A[457]), .Z(n1208) );
  XOR U1813 ( .A(A[456]), .B(n1209), .Z(O[456]) );
  AND U1814 ( .A(S), .B(n1210), .Z(n1209) );
  XOR U1815 ( .A(B[456]), .B(A[456]), .Z(n1210) );
  XOR U1816 ( .A(A[455]), .B(n1211), .Z(O[455]) );
  AND U1817 ( .A(S), .B(n1212), .Z(n1211) );
  XOR U1818 ( .A(B[455]), .B(A[455]), .Z(n1212) );
  XOR U1819 ( .A(A[454]), .B(n1213), .Z(O[454]) );
  AND U1820 ( .A(S), .B(n1214), .Z(n1213) );
  XOR U1821 ( .A(B[454]), .B(A[454]), .Z(n1214) );
  XOR U1822 ( .A(A[453]), .B(n1215), .Z(O[453]) );
  AND U1823 ( .A(S), .B(n1216), .Z(n1215) );
  XOR U1824 ( .A(B[453]), .B(A[453]), .Z(n1216) );
  XOR U1825 ( .A(A[452]), .B(n1217), .Z(O[452]) );
  AND U1826 ( .A(S), .B(n1218), .Z(n1217) );
  XOR U1827 ( .A(B[452]), .B(A[452]), .Z(n1218) );
  XOR U1828 ( .A(A[451]), .B(n1219), .Z(O[451]) );
  AND U1829 ( .A(S), .B(n1220), .Z(n1219) );
  XOR U1830 ( .A(B[451]), .B(A[451]), .Z(n1220) );
  XOR U1831 ( .A(A[450]), .B(n1221), .Z(O[450]) );
  AND U1832 ( .A(S), .B(n1222), .Z(n1221) );
  XOR U1833 ( .A(B[450]), .B(A[450]), .Z(n1222) );
  XOR U1834 ( .A(A[44]), .B(n1223), .Z(O[44]) );
  AND U1835 ( .A(S), .B(n1224), .Z(n1223) );
  XOR U1836 ( .A(B[44]), .B(A[44]), .Z(n1224) );
  XOR U1837 ( .A(A[449]), .B(n1225), .Z(O[449]) );
  AND U1838 ( .A(S), .B(n1226), .Z(n1225) );
  XOR U1839 ( .A(B[449]), .B(A[449]), .Z(n1226) );
  XOR U1840 ( .A(A[448]), .B(n1227), .Z(O[448]) );
  AND U1841 ( .A(S), .B(n1228), .Z(n1227) );
  XOR U1842 ( .A(B[448]), .B(A[448]), .Z(n1228) );
  XOR U1843 ( .A(A[447]), .B(n1229), .Z(O[447]) );
  AND U1844 ( .A(S), .B(n1230), .Z(n1229) );
  XOR U1845 ( .A(B[447]), .B(A[447]), .Z(n1230) );
  XOR U1846 ( .A(A[446]), .B(n1231), .Z(O[446]) );
  AND U1847 ( .A(S), .B(n1232), .Z(n1231) );
  XOR U1848 ( .A(B[446]), .B(A[446]), .Z(n1232) );
  XOR U1849 ( .A(A[445]), .B(n1233), .Z(O[445]) );
  AND U1850 ( .A(S), .B(n1234), .Z(n1233) );
  XOR U1851 ( .A(B[445]), .B(A[445]), .Z(n1234) );
  XOR U1852 ( .A(A[444]), .B(n1235), .Z(O[444]) );
  AND U1853 ( .A(S), .B(n1236), .Z(n1235) );
  XOR U1854 ( .A(B[444]), .B(A[444]), .Z(n1236) );
  XOR U1855 ( .A(A[443]), .B(n1237), .Z(O[443]) );
  AND U1856 ( .A(S), .B(n1238), .Z(n1237) );
  XOR U1857 ( .A(B[443]), .B(A[443]), .Z(n1238) );
  XOR U1858 ( .A(A[442]), .B(n1239), .Z(O[442]) );
  AND U1859 ( .A(S), .B(n1240), .Z(n1239) );
  XOR U1860 ( .A(B[442]), .B(A[442]), .Z(n1240) );
  XOR U1861 ( .A(A[441]), .B(n1241), .Z(O[441]) );
  AND U1862 ( .A(S), .B(n1242), .Z(n1241) );
  XOR U1863 ( .A(B[441]), .B(A[441]), .Z(n1242) );
  XOR U1864 ( .A(A[440]), .B(n1243), .Z(O[440]) );
  AND U1865 ( .A(S), .B(n1244), .Z(n1243) );
  XOR U1866 ( .A(B[440]), .B(A[440]), .Z(n1244) );
  XOR U1867 ( .A(A[43]), .B(n1245), .Z(O[43]) );
  AND U1868 ( .A(S), .B(n1246), .Z(n1245) );
  XOR U1869 ( .A(B[43]), .B(A[43]), .Z(n1246) );
  XOR U1870 ( .A(A[439]), .B(n1247), .Z(O[439]) );
  AND U1871 ( .A(S), .B(n1248), .Z(n1247) );
  XOR U1872 ( .A(B[439]), .B(A[439]), .Z(n1248) );
  XOR U1873 ( .A(A[438]), .B(n1249), .Z(O[438]) );
  AND U1874 ( .A(S), .B(n1250), .Z(n1249) );
  XOR U1875 ( .A(B[438]), .B(A[438]), .Z(n1250) );
  XOR U1876 ( .A(A[437]), .B(n1251), .Z(O[437]) );
  AND U1877 ( .A(S), .B(n1252), .Z(n1251) );
  XOR U1878 ( .A(B[437]), .B(A[437]), .Z(n1252) );
  XOR U1879 ( .A(A[436]), .B(n1253), .Z(O[436]) );
  AND U1880 ( .A(S), .B(n1254), .Z(n1253) );
  XOR U1881 ( .A(B[436]), .B(A[436]), .Z(n1254) );
  XOR U1882 ( .A(A[435]), .B(n1255), .Z(O[435]) );
  AND U1883 ( .A(S), .B(n1256), .Z(n1255) );
  XOR U1884 ( .A(B[435]), .B(A[435]), .Z(n1256) );
  XOR U1885 ( .A(A[434]), .B(n1257), .Z(O[434]) );
  AND U1886 ( .A(S), .B(n1258), .Z(n1257) );
  XOR U1887 ( .A(B[434]), .B(A[434]), .Z(n1258) );
  XOR U1888 ( .A(A[433]), .B(n1259), .Z(O[433]) );
  AND U1889 ( .A(S), .B(n1260), .Z(n1259) );
  XOR U1890 ( .A(B[433]), .B(A[433]), .Z(n1260) );
  XOR U1891 ( .A(A[432]), .B(n1261), .Z(O[432]) );
  AND U1892 ( .A(S), .B(n1262), .Z(n1261) );
  XOR U1893 ( .A(B[432]), .B(A[432]), .Z(n1262) );
  XOR U1894 ( .A(A[431]), .B(n1263), .Z(O[431]) );
  AND U1895 ( .A(S), .B(n1264), .Z(n1263) );
  XOR U1896 ( .A(B[431]), .B(A[431]), .Z(n1264) );
  XOR U1897 ( .A(A[430]), .B(n1265), .Z(O[430]) );
  AND U1898 ( .A(S), .B(n1266), .Z(n1265) );
  XOR U1899 ( .A(B[430]), .B(A[430]), .Z(n1266) );
  XOR U1900 ( .A(A[42]), .B(n1267), .Z(O[42]) );
  AND U1901 ( .A(S), .B(n1268), .Z(n1267) );
  XOR U1902 ( .A(B[42]), .B(A[42]), .Z(n1268) );
  XOR U1903 ( .A(A[429]), .B(n1269), .Z(O[429]) );
  AND U1904 ( .A(S), .B(n1270), .Z(n1269) );
  XOR U1905 ( .A(B[429]), .B(A[429]), .Z(n1270) );
  XOR U1906 ( .A(A[428]), .B(n1271), .Z(O[428]) );
  AND U1907 ( .A(S), .B(n1272), .Z(n1271) );
  XOR U1908 ( .A(B[428]), .B(A[428]), .Z(n1272) );
  XOR U1909 ( .A(A[427]), .B(n1273), .Z(O[427]) );
  AND U1910 ( .A(S), .B(n1274), .Z(n1273) );
  XOR U1911 ( .A(B[427]), .B(A[427]), .Z(n1274) );
  XOR U1912 ( .A(A[426]), .B(n1275), .Z(O[426]) );
  AND U1913 ( .A(S), .B(n1276), .Z(n1275) );
  XOR U1914 ( .A(B[426]), .B(A[426]), .Z(n1276) );
  XOR U1915 ( .A(A[425]), .B(n1277), .Z(O[425]) );
  AND U1916 ( .A(S), .B(n1278), .Z(n1277) );
  XOR U1917 ( .A(B[425]), .B(A[425]), .Z(n1278) );
  XOR U1918 ( .A(A[424]), .B(n1279), .Z(O[424]) );
  AND U1919 ( .A(S), .B(n1280), .Z(n1279) );
  XOR U1920 ( .A(B[424]), .B(A[424]), .Z(n1280) );
  XOR U1921 ( .A(A[423]), .B(n1281), .Z(O[423]) );
  AND U1922 ( .A(S), .B(n1282), .Z(n1281) );
  XOR U1923 ( .A(B[423]), .B(A[423]), .Z(n1282) );
  XOR U1924 ( .A(A[422]), .B(n1283), .Z(O[422]) );
  AND U1925 ( .A(S), .B(n1284), .Z(n1283) );
  XOR U1926 ( .A(B[422]), .B(A[422]), .Z(n1284) );
  XOR U1927 ( .A(A[421]), .B(n1285), .Z(O[421]) );
  AND U1928 ( .A(S), .B(n1286), .Z(n1285) );
  XOR U1929 ( .A(B[421]), .B(A[421]), .Z(n1286) );
  XOR U1930 ( .A(A[420]), .B(n1287), .Z(O[420]) );
  AND U1931 ( .A(S), .B(n1288), .Z(n1287) );
  XOR U1932 ( .A(B[420]), .B(A[420]), .Z(n1288) );
  XOR U1933 ( .A(A[41]), .B(n1289), .Z(O[41]) );
  AND U1934 ( .A(S), .B(n1290), .Z(n1289) );
  XOR U1935 ( .A(B[41]), .B(A[41]), .Z(n1290) );
  XOR U1936 ( .A(A[419]), .B(n1291), .Z(O[419]) );
  AND U1937 ( .A(S), .B(n1292), .Z(n1291) );
  XOR U1938 ( .A(B[419]), .B(A[419]), .Z(n1292) );
  XOR U1939 ( .A(A[418]), .B(n1293), .Z(O[418]) );
  AND U1940 ( .A(S), .B(n1294), .Z(n1293) );
  XOR U1941 ( .A(B[418]), .B(A[418]), .Z(n1294) );
  XOR U1942 ( .A(A[417]), .B(n1295), .Z(O[417]) );
  AND U1943 ( .A(S), .B(n1296), .Z(n1295) );
  XOR U1944 ( .A(B[417]), .B(A[417]), .Z(n1296) );
  XOR U1945 ( .A(A[416]), .B(n1297), .Z(O[416]) );
  AND U1946 ( .A(S), .B(n1298), .Z(n1297) );
  XOR U1947 ( .A(B[416]), .B(A[416]), .Z(n1298) );
  XOR U1948 ( .A(A[415]), .B(n1299), .Z(O[415]) );
  AND U1949 ( .A(S), .B(n1300), .Z(n1299) );
  XOR U1950 ( .A(B[415]), .B(A[415]), .Z(n1300) );
  XOR U1951 ( .A(A[414]), .B(n1301), .Z(O[414]) );
  AND U1952 ( .A(S), .B(n1302), .Z(n1301) );
  XOR U1953 ( .A(B[414]), .B(A[414]), .Z(n1302) );
  XOR U1954 ( .A(A[413]), .B(n1303), .Z(O[413]) );
  AND U1955 ( .A(S), .B(n1304), .Z(n1303) );
  XOR U1956 ( .A(B[413]), .B(A[413]), .Z(n1304) );
  XOR U1957 ( .A(A[412]), .B(n1305), .Z(O[412]) );
  AND U1958 ( .A(S), .B(n1306), .Z(n1305) );
  XOR U1959 ( .A(B[412]), .B(A[412]), .Z(n1306) );
  XOR U1960 ( .A(A[411]), .B(n1307), .Z(O[411]) );
  AND U1961 ( .A(S), .B(n1308), .Z(n1307) );
  XOR U1962 ( .A(B[411]), .B(A[411]), .Z(n1308) );
  XOR U1963 ( .A(A[410]), .B(n1309), .Z(O[410]) );
  AND U1964 ( .A(S), .B(n1310), .Z(n1309) );
  XOR U1965 ( .A(B[410]), .B(A[410]), .Z(n1310) );
  XOR U1966 ( .A(A[40]), .B(n1311), .Z(O[40]) );
  AND U1967 ( .A(S), .B(n1312), .Z(n1311) );
  XOR U1968 ( .A(B[40]), .B(A[40]), .Z(n1312) );
  XOR U1969 ( .A(A[409]), .B(n1313), .Z(O[409]) );
  AND U1970 ( .A(S), .B(n1314), .Z(n1313) );
  XOR U1971 ( .A(B[409]), .B(A[409]), .Z(n1314) );
  XOR U1972 ( .A(A[408]), .B(n1315), .Z(O[408]) );
  AND U1973 ( .A(S), .B(n1316), .Z(n1315) );
  XOR U1974 ( .A(B[408]), .B(A[408]), .Z(n1316) );
  XOR U1975 ( .A(A[407]), .B(n1317), .Z(O[407]) );
  AND U1976 ( .A(S), .B(n1318), .Z(n1317) );
  XOR U1977 ( .A(B[407]), .B(A[407]), .Z(n1318) );
  XOR U1978 ( .A(A[406]), .B(n1319), .Z(O[406]) );
  AND U1979 ( .A(S), .B(n1320), .Z(n1319) );
  XOR U1980 ( .A(B[406]), .B(A[406]), .Z(n1320) );
  XOR U1981 ( .A(A[405]), .B(n1321), .Z(O[405]) );
  AND U1982 ( .A(S), .B(n1322), .Z(n1321) );
  XOR U1983 ( .A(B[405]), .B(A[405]), .Z(n1322) );
  XOR U1984 ( .A(A[404]), .B(n1323), .Z(O[404]) );
  AND U1985 ( .A(S), .B(n1324), .Z(n1323) );
  XOR U1986 ( .A(B[404]), .B(A[404]), .Z(n1324) );
  XOR U1987 ( .A(A[403]), .B(n1325), .Z(O[403]) );
  AND U1988 ( .A(S), .B(n1326), .Z(n1325) );
  XOR U1989 ( .A(B[403]), .B(A[403]), .Z(n1326) );
  XOR U1990 ( .A(A[402]), .B(n1327), .Z(O[402]) );
  AND U1991 ( .A(S), .B(n1328), .Z(n1327) );
  XOR U1992 ( .A(B[402]), .B(A[402]), .Z(n1328) );
  XOR U1993 ( .A(A[401]), .B(n1329), .Z(O[401]) );
  AND U1994 ( .A(S), .B(n1330), .Z(n1329) );
  XOR U1995 ( .A(B[401]), .B(A[401]), .Z(n1330) );
  XOR U1996 ( .A(A[400]), .B(n1331), .Z(O[400]) );
  AND U1997 ( .A(S), .B(n1332), .Z(n1331) );
  XOR U1998 ( .A(B[400]), .B(A[400]), .Z(n1332) );
  XOR U1999 ( .A(A[3]), .B(n1333), .Z(O[3]) );
  AND U2000 ( .A(S), .B(n1334), .Z(n1333) );
  XOR U2001 ( .A(B[3]), .B(A[3]), .Z(n1334) );
  XOR U2002 ( .A(A[39]), .B(n1335), .Z(O[39]) );
  AND U2003 ( .A(S), .B(n1336), .Z(n1335) );
  XOR U2004 ( .A(B[39]), .B(A[39]), .Z(n1336) );
  XOR U2005 ( .A(A[399]), .B(n1337), .Z(O[399]) );
  AND U2006 ( .A(S), .B(n1338), .Z(n1337) );
  XOR U2007 ( .A(B[399]), .B(A[399]), .Z(n1338) );
  XOR U2008 ( .A(A[398]), .B(n1339), .Z(O[398]) );
  AND U2009 ( .A(S), .B(n1340), .Z(n1339) );
  XOR U2010 ( .A(B[398]), .B(A[398]), .Z(n1340) );
  XOR U2011 ( .A(A[397]), .B(n1341), .Z(O[397]) );
  AND U2012 ( .A(S), .B(n1342), .Z(n1341) );
  XOR U2013 ( .A(B[397]), .B(A[397]), .Z(n1342) );
  XOR U2014 ( .A(A[396]), .B(n1343), .Z(O[396]) );
  AND U2015 ( .A(S), .B(n1344), .Z(n1343) );
  XOR U2016 ( .A(B[396]), .B(A[396]), .Z(n1344) );
  XOR U2017 ( .A(A[395]), .B(n1345), .Z(O[395]) );
  AND U2018 ( .A(S), .B(n1346), .Z(n1345) );
  XOR U2019 ( .A(B[395]), .B(A[395]), .Z(n1346) );
  XOR U2020 ( .A(A[394]), .B(n1347), .Z(O[394]) );
  AND U2021 ( .A(S), .B(n1348), .Z(n1347) );
  XOR U2022 ( .A(B[394]), .B(A[394]), .Z(n1348) );
  XOR U2023 ( .A(A[393]), .B(n1349), .Z(O[393]) );
  AND U2024 ( .A(S), .B(n1350), .Z(n1349) );
  XOR U2025 ( .A(B[393]), .B(A[393]), .Z(n1350) );
  XOR U2026 ( .A(A[392]), .B(n1351), .Z(O[392]) );
  AND U2027 ( .A(S), .B(n1352), .Z(n1351) );
  XOR U2028 ( .A(B[392]), .B(A[392]), .Z(n1352) );
  XOR U2029 ( .A(A[391]), .B(n1353), .Z(O[391]) );
  AND U2030 ( .A(S), .B(n1354), .Z(n1353) );
  XOR U2031 ( .A(B[391]), .B(A[391]), .Z(n1354) );
  XOR U2032 ( .A(A[390]), .B(n1355), .Z(O[390]) );
  AND U2033 ( .A(S), .B(n1356), .Z(n1355) );
  XOR U2034 ( .A(B[390]), .B(A[390]), .Z(n1356) );
  XOR U2035 ( .A(A[38]), .B(n1357), .Z(O[38]) );
  AND U2036 ( .A(S), .B(n1358), .Z(n1357) );
  XOR U2037 ( .A(B[38]), .B(A[38]), .Z(n1358) );
  XOR U2038 ( .A(A[389]), .B(n1359), .Z(O[389]) );
  AND U2039 ( .A(S), .B(n1360), .Z(n1359) );
  XOR U2040 ( .A(B[389]), .B(A[389]), .Z(n1360) );
  XOR U2041 ( .A(A[388]), .B(n1361), .Z(O[388]) );
  AND U2042 ( .A(S), .B(n1362), .Z(n1361) );
  XOR U2043 ( .A(B[388]), .B(A[388]), .Z(n1362) );
  XOR U2044 ( .A(A[387]), .B(n1363), .Z(O[387]) );
  AND U2045 ( .A(S), .B(n1364), .Z(n1363) );
  XOR U2046 ( .A(B[387]), .B(A[387]), .Z(n1364) );
  XOR U2047 ( .A(A[386]), .B(n1365), .Z(O[386]) );
  AND U2048 ( .A(S), .B(n1366), .Z(n1365) );
  XOR U2049 ( .A(B[386]), .B(A[386]), .Z(n1366) );
  XOR U2050 ( .A(A[385]), .B(n1367), .Z(O[385]) );
  AND U2051 ( .A(S), .B(n1368), .Z(n1367) );
  XOR U2052 ( .A(B[385]), .B(A[385]), .Z(n1368) );
  XOR U2053 ( .A(A[384]), .B(n1369), .Z(O[384]) );
  AND U2054 ( .A(S), .B(n1370), .Z(n1369) );
  XOR U2055 ( .A(B[384]), .B(A[384]), .Z(n1370) );
  XOR U2056 ( .A(A[383]), .B(n1371), .Z(O[383]) );
  AND U2057 ( .A(S), .B(n1372), .Z(n1371) );
  XOR U2058 ( .A(B[383]), .B(A[383]), .Z(n1372) );
  XOR U2059 ( .A(A[382]), .B(n1373), .Z(O[382]) );
  AND U2060 ( .A(S), .B(n1374), .Z(n1373) );
  XOR U2061 ( .A(B[382]), .B(A[382]), .Z(n1374) );
  XOR U2062 ( .A(A[381]), .B(n1375), .Z(O[381]) );
  AND U2063 ( .A(S), .B(n1376), .Z(n1375) );
  XOR U2064 ( .A(B[381]), .B(A[381]), .Z(n1376) );
  XOR U2065 ( .A(A[380]), .B(n1377), .Z(O[380]) );
  AND U2066 ( .A(S), .B(n1378), .Z(n1377) );
  XOR U2067 ( .A(B[380]), .B(A[380]), .Z(n1378) );
  XOR U2068 ( .A(A[37]), .B(n1379), .Z(O[37]) );
  AND U2069 ( .A(S), .B(n1380), .Z(n1379) );
  XOR U2070 ( .A(B[37]), .B(A[37]), .Z(n1380) );
  XOR U2071 ( .A(A[379]), .B(n1381), .Z(O[379]) );
  AND U2072 ( .A(S), .B(n1382), .Z(n1381) );
  XOR U2073 ( .A(B[379]), .B(A[379]), .Z(n1382) );
  XOR U2074 ( .A(A[378]), .B(n1383), .Z(O[378]) );
  AND U2075 ( .A(S), .B(n1384), .Z(n1383) );
  XOR U2076 ( .A(B[378]), .B(A[378]), .Z(n1384) );
  XOR U2077 ( .A(A[377]), .B(n1385), .Z(O[377]) );
  AND U2078 ( .A(S), .B(n1386), .Z(n1385) );
  XOR U2079 ( .A(B[377]), .B(A[377]), .Z(n1386) );
  XOR U2080 ( .A(A[376]), .B(n1387), .Z(O[376]) );
  AND U2081 ( .A(S), .B(n1388), .Z(n1387) );
  XOR U2082 ( .A(B[376]), .B(A[376]), .Z(n1388) );
  XOR U2083 ( .A(A[375]), .B(n1389), .Z(O[375]) );
  AND U2084 ( .A(S), .B(n1390), .Z(n1389) );
  XOR U2085 ( .A(B[375]), .B(A[375]), .Z(n1390) );
  XOR U2086 ( .A(A[374]), .B(n1391), .Z(O[374]) );
  AND U2087 ( .A(S), .B(n1392), .Z(n1391) );
  XOR U2088 ( .A(B[374]), .B(A[374]), .Z(n1392) );
  XOR U2089 ( .A(A[373]), .B(n1393), .Z(O[373]) );
  AND U2090 ( .A(S), .B(n1394), .Z(n1393) );
  XOR U2091 ( .A(B[373]), .B(A[373]), .Z(n1394) );
  XOR U2092 ( .A(A[372]), .B(n1395), .Z(O[372]) );
  AND U2093 ( .A(S), .B(n1396), .Z(n1395) );
  XOR U2094 ( .A(B[372]), .B(A[372]), .Z(n1396) );
  XOR U2095 ( .A(A[371]), .B(n1397), .Z(O[371]) );
  AND U2096 ( .A(S), .B(n1398), .Z(n1397) );
  XOR U2097 ( .A(B[371]), .B(A[371]), .Z(n1398) );
  XOR U2098 ( .A(A[370]), .B(n1399), .Z(O[370]) );
  AND U2099 ( .A(S), .B(n1400), .Z(n1399) );
  XOR U2100 ( .A(B[370]), .B(A[370]), .Z(n1400) );
  XOR U2101 ( .A(A[36]), .B(n1401), .Z(O[36]) );
  AND U2102 ( .A(S), .B(n1402), .Z(n1401) );
  XOR U2103 ( .A(B[36]), .B(A[36]), .Z(n1402) );
  XOR U2104 ( .A(A[369]), .B(n1403), .Z(O[369]) );
  AND U2105 ( .A(S), .B(n1404), .Z(n1403) );
  XOR U2106 ( .A(B[369]), .B(A[369]), .Z(n1404) );
  XOR U2107 ( .A(A[368]), .B(n1405), .Z(O[368]) );
  AND U2108 ( .A(S), .B(n1406), .Z(n1405) );
  XOR U2109 ( .A(B[368]), .B(A[368]), .Z(n1406) );
  XOR U2110 ( .A(A[367]), .B(n1407), .Z(O[367]) );
  AND U2111 ( .A(S), .B(n1408), .Z(n1407) );
  XOR U2112 ( .A(B[367]), .B(A[367]), .Z(n1408) );
  XOR U2113 ( .A(A[366]), .B(n1409), .Z(O[366]) );
  AND U2114 ( .A(S), .B(n1410), .Z(n1409) );
  XOR U2115 ( .A(B[366]), .B(A[366]), .Z(n1410) );
  XOR U2116 ( .A(A[365]), .B(n1411), .Z(O[365]) );
  AND U2117 ( .A(S), .B(n1412), .Z(n1411) );
  XOR U2118 ( .A(B[365]), .B(A[365]), .Z(n1412) );
  XOR U2119 ( .A(A[364]), .B(n1413), .Z(O[364]) );
  AND U2120 ( .A(S), .B(n1414), .Z(n1413) );
  XOR U2121 ( .A(B[364]), .B(A[364]), .Z(n1414) );
  XOR U2122 ( .A(A[363]), .B(n1415), .Z(O[363]) );
  AND U2123 ( .A(S), .B(n1416), .Z(n1415) );
  XOR U2124 ( .A(B[363]), .B(A[363]), .Z(n1416) );
  XOR U2125 ( .A(A[362]), .B(n1417), .Z(O[362]) );
  AND U2126 ( .A(S), .B(n1418), .Z(n1417) );
  XOR U2127 ( .A(B[362]), .B(A[362]), .Z(n1418) );
  XOR U2128 ( .A(A[361]), .B(n1419), .Z(O[361]) );
  AND U2129 ( .A(S), .B(n1420), .Z(n1419) );
  XOR U2130 ( .A(B[361]), .B(A[361]), .Z(n1420) );
  XOR U2131 ( .A(A[360]), .B(n1421), .Z(O[360]) );
  AND U2132 ( .A(S), .B(n1422), .Z(n1421) );
  XOR U2133 ( .A(B[360]), .B(A[360]), .Z(n1422) );
  XOR U2134 ( .A(A[35]), .B(n1423), .Z(O[35]) );
  AND U2135 ( .A(S), .B(n1424), .Z(n1423) );
  XOR U2136 ( .A(B[35]), .B(A[35]), .Z(n1424) );
  XOR U2137 ( .A(A[359]), .B(n1425), .Z(O[359]) );
  AND U2138 ( .A(S), .B(n1426), .Z(n1425) );
  XOR U2139 ( .A(B[359]), .B(A[359]), .Z(n1426) );
  XOR U2140 ( .A(A[358]), .B(n1427), .Z(O[358]) );
  AND U2141 ( .A(S), .B(n1428), .Z(n1427) );
  XOR U2142 ( .A(B[358]), .B(A[358]), .Z(n1428) );
  XOR U2143 ( .A(A[357]), .B(n1429), .Z(O[357]) );
  AND U2144 ( .A(S), .B(n1430), .Z(n1429) );
  XOR U2145 ( .A(B[357]), .B(A[357]), .Z(n1430) );
  XOR U2146 ( .A(A[356]), .B(n1431), .Z(O[356]) );
  AND U2147 ( .A(S), .B(n1432), .Z(n1431) );
  XOR U2148 ( .A(B[356]), .B(A[356]), .Z(n1432) );
  XOR U2149 ( .A(A[355]), .B(n1433), .Z(O[355]) );
  AND U2150 ( .A(S), .B(n1434), .Z(n1433) );
  XOR U2151 ( .A(B[355]), .B(A[355]), .Z(n1434) );
  XOR U2152 ( .A(A[354]), .B(n1435), .Z(O[354]) );
  AND U2153 ( .A(S), .B(n1436), .Z(n1435) );
  XOR U2154 ( .A(B[354]), .B(A[354]), .Z(n1436) );
  XOR U2155 ( .A(A[353]), .B(n1437), .Z(O[353]) );
  AND U2156 ( .A(S), .B(n1438), .Z(n1437) );
  XOR U2157 ( .A(B[353]), .B(A[353]), .Z(n1438) );
  XOR U2158 ( .A(A[352]), .B(n1439), .Z(O[352]) );
  AND U2159 ( .A(S), .B(n1440), .Z(n1439) );
  XOR U2160 ( .A(B[352]), .B(A[352]), .Z(n1440) );
  XOR U2161 ( .A(A[351]), .B(n1441), .Z(O[351]) );
  AND U2162 ( .A(S), .B(n1442), .Z(n1441) );
  XOR U2163 ( .A(B[351]), .B(A[351]), .Z(n1442) );
  XOR U2164 ( .A(A[350]), .B(n1443), .Z(O[350]) );
  AND U2165 ( .A(S), .B(n1444), .Z(n1443) );
  XOR U2166 ( .A(B[350]), .B(A[350]), .Z(n1444) );
  XOR U2167 ( .A(A[34]), .B(n1445), .Z(O[34]) );
  AND U2168 ( .A(S), .B(n1446), .Z(n1445) );
  XOR U2169 ( .A(B[34]), .B(A[34]), .Z(n1446) );
  XOR U2170 ( .A(A[349]), .B(n1447), .Z(O[349]) );
  AND U2171 ( .A(S), .B(n1448), .Z(n1447) );
  XOR U2172 ( .A(B[349]), .B(A[349]), .Z(n1448) );
  XOR U2173 ( .A(A[348]), .B(n1449), .Z(O[348]) );
  AND U2174 ( .A(S), .B(n1450), .Z(n1449) );
  XOR U2175 ( .A(B[348]), .B(A[348]), .Z(n1450) );
  XOR U2176 ( .A(A[347]), .B(n1451), .Z(O[347]) );
  AND U2177 ( .A(S), .B(n1452), .Z(n1451) );
  XOR U2178 ( .A(B[347]), .B(A[347]), .Z(n1452) );
  XOR U2179 ( .A(A[346]), .B(n1453), .Z(O[346]) );
  AND U2180 ( .A(S), .B(n1454), .Z(n1453) );
  XOR U2181 ( .A(B[346]), .B(A[346]), .Z(n1454) );
  XOR U2182 ( .A(A[345]), .B(n1455), .Z(O[345]) );
  AND U2183 ( .A(S), .B(n1456), .Z(n1455) );
  XOR U2184 ( .A(B[345]), .B(A[345]), .Z(n1456) );
  XOR U2185 ( .A(A[344]), .B(n1457), .Z(O[344]) );
  AND U2186 ( .A(S), .B(n1458), .Z(n1457) );
  XOR U2187 ( .A(B[344]), .B(A[344]), .Z(n1458) );
  XOR U2188 ( .A(A[343]), .B(n1459), .Z(O[343]) );
  AND U2189 ( .A(S), .B(n1460), .Z(n1459) );
  XOR U2190 ( .A(B[343]), .B(A[343]), .Z(n1460) );
  XOR U2191 ( .A(A[342]), .B(n1461), .Z(O[342]) );
  AND U2192 ( .A(S), .B(n1462), .Z(n1461) );
  XOR U2193 ( .A(B[342]), .B(A[342]), .Z(n1462) );
  XOR U2194 ( .A(A[341]), .B(n1463), .Z(O[341]) );
  AND U2195 ( .A(S), .B(n1464), .Z(n1463) );
  XOR U2196 ( .A(B[341]), .B(A[341]), .Z(n1464) );
  XOR U2197 ( .A(A[340]), .B(n1465), .Z(O[340]) );
  AND U2198 ( .A(S), .B(n1466), .Z(n1465) );
  XOR U2199 ( .A(B[340]), .B(A[340]), .Z(n1466) );
  XOR U2200 ( .A(A[33]), .B(n1467), .Z(O[33]) );
  AND U2201 ( .A(S), .B(n1468), .Z(n1467) );
  XOR U2202 ( .A(B[33]), .B(A[33]), .Z(n1468) );
  XOR U2203 ( .A(A[339]), .B(n1469), .Z(O[339]) );
  AND U2204 ( .A(S), .B(n1470), .Z(n1469) );
  XOR U2205 ( .A(B[339]), .B(A[339]), .Z(n1470) );
  XOR U2206 ( .A(A[338]), .B(n1471), .Z(O[338]) );
  AND U2207 ( .A(S), .B(n1472), .Z(n1471) );
  XOR U2208 ( .A(B[338]), .B(A[338]), .Z(n1472) );
  XOR U2209 ( .A(A[337]), .B(n1473), .Z(O[337]) );
  AND U2210 ( .A(S), .B(n1474), .Z(n1473) );
  XOR U2211 ( .A(B[337]), .B(A[337]), .Z(n1474) );
  XOR U2212 ( .A(A[336]), .B(n1475), .Z(O[336]) );
  AND U2213 ( .A(S), .B(n1476), .Z(n1475) );
  XOR U2214 ( .A(B[336]), .B(A[336]), .Z(n1476) );
  XOR U2215 ( .A(A[335]), .B(n1477), .Z(O[335]) );
  AND U2216 ( .A(S), .B(n1478), .Z(n1477) );
  XOR U2217 ( .A(B[335]), .B(A[335]), .Z(n1478) );
  XOR U2218 ( .A(A[334]), .B(n1479), .Z(O[334]) );
  AND U2219 ( .A(S), .B(n1480), .Z(n1479) );
  XOR U2220 ( .A(B[334]), .B(A[334]), .Z(n1480) );
  XOR U2221 ( .A(A[333]), .B(n1481), .Z(O[333]) );
  AND U2222 ( .A(S), .B(n1482), .Z(n1481) );
  XOR U2223 ( .A(B[333]), .B(A[333]), .Z(n1482) );
  XOR U2224 ( .A(A[332]), .B(n1483), .Z(O[332]) );
  AND U2225 ( .A(S), .B(n1484), .Z(n1483) );
  XOR U2226 ( .A(B[332]), .B(A[332]), .Z(n1484) );
  XOR U2227 ( .A(A[331]), .B(n1485), .Z(O[331]) );
  AND U2228 ( .A(S), .B(n1486), .Z(n1485) );
  XOR U2229 ( .A(B[331]), .B(A[331]), .Z(n1486) );
  XOR U2230 ( .A(A[330]), .B(n1487), .Z(O[330]) );
  AND U2231 ( .A(S), .B(n1488), .Z(n1487) );
  XOR U2232 ( .A(B[330]), .B(A[330]), .Z(n1488) );
  XOR U2233 ( .A(A[32]), .B(n1489), .Z(O[32]) );
  AND U2234 ( .A(S), .B(n1490), .Z(n1489) );
  XOR U2235 ( .A(B[32]), .B(A[32]), .Z(n1490) );
  XOR U2236 ( .A(A[329]), .B(n1491), .Z(O[329]) );
  AND U2237 ( .A(S), .B(n1492), .Z(n1491) );
  XOR U2238 ( .A(B[329]), .B(A[329]), .Z(n1492) );
  XOR U2239 ( .A(A[328]), .B(n1493), .Z(O[328]) );
  AND U2240 ( .A(S), .B(n1494), .Z(n1493) );
  XOR U2241 ( .A(B[328]), .B(A[328]), .Z(n1494) );
  XOR U2242 ( .A(A[327]), .B(n1495), .Z(O[327]) );
  AND U2243 ( .A(S), .B(n1496), .Z(n1495) );
  XOR U2244 ( .A(B[327]), .B(A[327]), .Z(n1496) );
  XOR U2245 ( .A(A[326]), .B(n1497), .Z(O[326]) );
  AND U2246 ( .A(S), .B(n1498), .Z(n1497) );
  XOR U2247 ( .A(B[326]), .B(A[326]), .Z(n1498) );
  XOR U2248 ( .A(A[325]), .B(n1499), .Z(O[325]) );
  AND U2249 ( .A(S), .B(n1500), .Z(n1499) );
  XOR U2250 ( .A(B[325]), .B(A[325]), .Z(n1500) );
  XOR U2251 ( .A(A[324]), .B(n1501), .Z(O[324]) );
  AND U2252 ( .A(S), .B(n1502), .Z(n1501) );
  XOR U2253 ( .A(B[324]), .B(A[324]), .Z(n1502) );
  XOR U2254 ( .A(A[323]), .B(n1503), .Z(O[323]) );
  AND U2255 ( .A(S), .B(n1504), .Z(n1503) );
  XOR U2256 ( .A(B[323]), .B(A[323]), .Z(n1504) );
  XOR U2257 ( .A(A[322]), .B(n1505), .Z(O[322]) );
  AND U2258 ( .A(S), .B(n1506), .Z(n1505) );
  XOR U2259 ( .A(B[322]), .B(A[322]), .Z(n1506) );
  XOR U2260 ( .A(A[321]), .B(n1507), .Z(O[321]) );
  AND U2261 ( .A(S), .B(n1508), .Z(n1507) );
  XOR U2262 ( .A(B[321]), .B(A[321]), .Z(n1508) );
  XOR U2263 ( .A(A[320]), .B(n1509), .Z(O[320]) );
  AND U2264 ( .A(S), .B(n1510), .Z(n1509) );
  XOR U2265 ( .A(B[320]), .B(A[320]), .Z(n1510) );
  XOR U2266 ( .A(A[31]), .B(n1511), .Z(O[31]) );
  AND U2267 ( .A(S), .B(n1512), .Z(n1511) );
  XOR U2268 ( .A(B[31]), .B(A[31]), .Z(n1512) );
  XOR U2269 ( .A(A[319]), .B(n1513), .Z(O[319]) );
  AND U2270 ( .A(S), .B(n1514), .Z(n1513) );
  XOR U2271 ( .A(B[319]), .B(A[319]), .Z(n1514) );
  XOR U2272 ( .A(A[318]), .B(n1515), .Z(O[318]) );
  AND U2273 ( .A(S), .B(n1516), .Z(n1515) );
  XOR U2274 ( .A(B[318]), .B(A[318]), .Z(n1516) );
  XOR U2275 ( .A(A[317]), .B(n1517), .Z(O[317]) );
  AND U2276 ( .A(S), .B(n1518), .Z(n1517) );
  XOR U2277 ( .A(B[317]), .B(A[317]), .Z(n1518) );
  XOR U2278 ( .A(A[316]), .B(n1519), .Z(O[316]) );
  AND U2279 ( .A(S), .B(n1520), .Z(n1519) );
  XOR U2280 ( .A(B[316]), .B(A[316]), .Z(n1520) );
  XOR U2281 ( .A(A[315]), .B(n1521), .Z(O[315]) );
  AND U2282 ( .A(S), .B(n1522), .Z(n1521) );
  XOR U2283 ( .A(B[315]), .B(A[315]), .Z(n1522) );
  XOR U2284 ( .A(A[314]), .B(n1523), .Z(O[314]) );
  AND U2285 ( .A(S), .B(n1524), .Z(n1523) );
  XOR U2286 ( .A(B[314]), .B(A[314]), .Z(n1524) );
  XOR U2287 ( .A(A[313]), .B(n1525), .Z(O[313]) );
  AND U2288 ( .A(S), .B(n1526), .Z(n1525) );
  XOR U2289 ( .A(B[313]), .B(A[313]), .Z(n1526) );
  XOR U2290 ( .A(A[312]), .B(n1527), .Z(O[312]) );
  AND U2291 ( .A(S), .B(n1528), .Z(n1527) );
  XOR U2292 ( .A(B[312]), .B(A[312]), .Z(n1528) );
  XOR U2293 ( .A(A[311]), .B(n1529), .Z(O[311]) );
  AND U2294 ( .A(S), .B(n1530), .Z(n1529) );
  XOR U2295 ( .A(B[311]), .B(A[311]), .Z(n1530) );
  XOR U2296 ( .A(A[310]), .B(n1531), .Z(O[310]) );
  AND U2297 ( .A(S), .B(n1532), .Z(n1531) );
  XOR U2298 ( .A(B[310]), .B(A[310]), .Z(n1532) );
  XOR U2299 ( .A(A[30]), .B(n1533), .Z(O[30]) );
  AND U2300 ( .A(S), .B(n1534), .Z(n1533) );
  XOR U2301 ( .A(B[30]), .B(A[30]), .Z(n1534) );
  XOR U2302 ( .A(A[309]), .B(n1535), .Z(O[309]) );
  AND U2303 ( .A(S), .B(n1536), .Z(n1535) );
  XOR U2304 ( .A(B[309]), .B(A[309]), .Z(n1536) );
  XOR U2305 ( .A(A[308]), .B(n1537), .Z(O[308]) );
  AND U2306 ( .A(S), .B(n1538), .Z(n1537) );
  XOR U2307 ( .A(B[308]), .B(A[308]), .Z(n1538) );
  XOR U2308 ( .A(A[307]), .B(n1539), .Z(O[307]) );
  AND U2309 ( .A(S), .B(n1540), .Z(n1539) );
  XOR U2310 ( .A(B[307]), .B(A[307]), .Z(n1540) );
  XOR U2311 ( .A(A[306]), .B(n1541), .Z(O[306]) );
  AND U2312 ( .A(S), .B(n1542), .Z(n1541) );
  XOR U2313 ( .A(B[306]), .B(A[306]), .Z(n1542) );
  XOR U2314 ( .A(A[305]), .B(n1543), .Z(O[305]) );
  AND U2315 ( .A(S), .B(n1544), .Z(n1543) );
  XOR U2316 ( .A(B[305]), .B(A[305]), .Z(n1544) );
  XOR U2317 ( .A(A[304]), .B(n1545), .Z(O[304]) );
  AND U2318 ( .A(S), .B(n1546), .Z(n1545) );
  XOR U2319 ( .A(B[304]), .B(A[304]), .Z(n1546) );
  XOR U2320 ( .A(A[303]), .B(n1547), .Z(O[303]) );
  AND U2321 ( .A(S), .B(n1548), .Z(n1547) );
  XOR U2322 ( .A(B[303]), .B(A[303]), .Z(n1548) );
  XOR U2323 ( .A(A[302]), .B(n1549), .Z(O[302]) );
  AND U2324 ( .A(S), .B(n1550), .Z(n1549) );
  XOR U2325 ( .A(B[302]), .B(A[302]), .Z(n1550) );
  XOR U2326 ( .A(A[301]), .B(n1551), .Z(O[301]) );
  AND U2327 ( .A(S), .B(n1552), .Z(n1551) );
  XOR U2328 ( .A(B[301]), .B(A[301]), .Z(n1552) );
  XOR U2329 ( .A(A[300]), .B(n1553), .Z(O[300]) );
  AND U2330 ( .A(S), .B(n1554), .Z(n1553) );
  XOR U2331 ( .A(B[300]), .B(A[300]), .Z(n1554) );
  XOR U2332 ( .A(A[2]), .B(n1555), .Z(O[2]) );
  AND U2333 ( .A(S), .B(n1556), .Z(n1555) );
  XOR U2334 ( .A(B[2]), .B(A[2]), .Z(n1556) );
  XOR U2335 ( .A(A[29]), .B(n1557), .Z(O[29]) );
  AND U2336 ( .A(S), .B(n1558), .Z(n1557) );
  XOR U2337 ( .A(B[29]), .B(A[29]), .Z(n1558) );
  XOR U2338 ( .A(A[299]), .B(n1559), .Z(O[299]) );
  AND U2339 ( .A(S), .B(n1560), .Z(n1559) );
  XOR U2340 ( .A(B[299]), .B(A[299]), .Z(n1560) );
  XOR U2341 ( .A(A[298]), .B(n1561), .Z(O[298]) );
  AND U2342 ( .A(S), .B(n1562), .Z(n1561) );
  XOR U2343 ( .A(B[298]), .B(A[298]), .Z(n1562) );
  XOR U2344 ( .A(A[297]), .B(n1563), .Z(O[297]) );
  AND U2345 ( .A(S), .B(n1564), .Z(n1563) );
  XOR U2346 ( .A(B[297]), .B(A[297]), .Z(n1564) );
  XOR U2347 ( .A(A[296]), .B(n1565), .Z(O[296]) );
  AND U2348 ( .A(S), .B(n1566), .Z(n1565) );
  XOR U2349 ( .A(B[296]), .B(A[296]), .Z(n1566) );
  XOR U2350 ( .A(A[295]), .B(n1567), .Z(O[295]) );
  AND U2351 ( .A(S), .B(n1568), .Z(n1567) );
  XOR U2352 ( .A(B[295]), .B(A[295]), .Z(n1568) );
  XOR U2353 ( .A(A[294]), .B(n1569), .Z(O[294]) );
  AND U2354 ( .A(S), .B(n1570), .Z(n1569) );
  XOR U2355 ( .A(B[294]), .B(A[294]), .Z(n1570) );
  XOR U2356 ( .A(A[293]), .B(n1571), .Z(O[293]) );
  AND U2357 ( .A(S), .B(n1572), .Z(n1571) );
  XOR U2358 ( .A(B[293]), .B(A[293]), .Z(n1572) );
  XOR U2359 ( .A(A[292]), .B(n1573), .Z(O[292]) );
  AND U2360 ( .A(S), .B(n1574), .Z(n1573) );
  XOR U2361 ( .A(B[292]), .B(A[292]), .Z(n1574) );
  XOR U2362 ( .A(A[291]), .B(n1575), .Z(O[291]) );
  AND U2363 ( .A(S), .B(n1576), .Z(n1575) );
  XOR U2364 ( .A(B[291]), .B(A[291]), .Z(n1576) );
  XOR U2365 ( .A(A[290]), .B(n1577), .Z(O[290]) );
  AND U2366 ( .A(S), .B(n1578), .Z(n1577) );
  XOR U2367 ( .A(B[290]), .B(A[290]), .Z(n1578) );
  XOR U2368 ( .A(A[28]), .B(n1579), .Z(O[28]) );
  AND U2369 ( .A(S), .B(n1580), .Z(n1579) );
  XOR U2370 ( .A(B[28]), .B(A[28]), .Z(n1580) );
  XOR U2371 ( .A(A[289]), .B(n1581), .Z(O[289]) );
  AND U2372 ( .A(S), .B(n1582), .Z(n1581) );
  XOR U2373 ( .A(B[289]), .B(A[289]), .Z(n1582) );
  XOR U2374 ( .A(A[288]), .B(n1583), .Z(O[288]) );
  AND U2375 ( .A(S), .B(n1584), .Z(n1583) );
  XOR U2376 ( .A(B[288]), .B(A[288]), .Z(n1584) );
  XOR U2377 ( .A(A[287]), .B(n1585), .Z(O[287]) );
  AND U2378 ( .A(S), .B(n1586), .Z(n1585) );
  XOR U2379 ( .A(B[287]), .B(A[287]), .Z(n1586) );
  XOR U2380 ( .A(A[286]), .B(n1587), .Z(O[286]) );
  AND U2381 ( .A(S), .B(n1588), .Z(n1587) );
  XOR U2382 ( .A(B[286]), .B(A[286]), .Z(n1588) );
  XOR U2383 ( .A(A[285]), .B(n1589), .Z(O[285]) );
  AND U2384 ( .A(S), .B(n1590), .Z(n1589) );
  XOR U2385 ( .A(B[285]), .B(A[285]), .Z(n1590) );
  XOR U2386 ( .A(A[284]), .B(n1591), .Z(O[284]) );
  AND U2387 ( .A(S), .B(n1592), .Z(n1591) );
  XOR U2388 ( .A(B[284]), .B(A[284]), .Z(n1592) );
  XOR U2389 ( .A(A[283]), .B(n1593), .Z(O[283]) );
  AND U2390 ( .A(S), .B(n1594), .Z(n1593) );
  XOR U2391 ( .A(B[283]), .B(A[283]), .Z(n1594) );
  XOR U2392 ( .A(A[282]), .B(n1595), .Z(O[282]) );
  AND U2393 ( .A(S), .B(n1596), .Z(n1595) );
  XOR U2394 ( .A(B[282]), .B(A[282]), .Z(n1596) );
  XOR U2395 ( .A(A[281]), .B(n1597), .Z(O[281]) );
  AND U2396 ( .A(S), .B(n1598), .Z(n1597) );
  XOR U2397 ( .A(B[281]), .B(A[281]), .Z(n1598) );
  XOR U2398 ( .A(A[280]), .B(n1599), .Z(O[280]) );
  AND U2399 ( .A(S), .B(n1600), .Z(n1599) );
  XOR U2400 ( .A(B[280]), .B(A[280]), .Z(n1600) );
  XOR U2401 ( .A(A[27]), .B(n1601), .Z(O[27]) );
  AND U2402 ( .A(S), .B(n1602), .Z(n1601) );
  XOR U2403 ( .A(B[27]), .B(A[27]), .Z(n1602) );
  XOR U2404 ( .A(A[279]), .B(n1603), .Z(O[279]) );
  AND U2405 ( .A(S), .B(n1604), .Z(n1603) );
  XOR U2406 ( .A(B[279]), .B(A[279]), .Z(n1604) );
  XOR U2407 ( .A(A[278]), .B(n1605), .Z(O[278]) );
  AND U2408 ( .A(S), .B(n1606), .Z(n1605) );
  XOR U2409 ( .A(B[278]), .B(A[278]), .Z(n1606) );
  XOR U2410 ( .A(A[277]), .B(n1607), .Z(O[277]) );
  AND U2411 ( .A(S), .B(n1608), .Z(n1607) );
  XOR U2412 ( .A(B[277]), .B(A[277]), .Z(n1608) );
  XOR U2413 ( .A(A[276]), .B(n1609), .Z(O[276]) );
  AND U2414 ( .A(S), .B(n1610), .Z(n1609) );
  XOR U2415 ( .A(B[276]), .B(A[276]), .Z(n1610) );
  XOR U2416 ( .A(A[275]), .B(n1611), .Z(O[275]) );
  AND U2417 ( .A(S), .B(n1612), .Z(n1611) );
  XOR U2418 ( .A(B[275]), .B(A[275]), .Z(n1612) );
  XOR U2419 ( .A(A[274]), .B(n1613), .Z(O[274]) );
  AND U2420 ( .A(S), .B(n1614), .Z(n1613) );
  XOR U2421 ( .A(B[274]), .B(A[274]), .Z(n1614) );
  XOR U2422 ( .A(A[273]), .B(n1615), .Z(O[273]) );
  AND U2423 ( .A(S), .B(n1616), .Z(n1615) );
  XOR U2424 ( .A(B[273]), .B(A[273]), .Z(n1616) );
  XOR U2425 ( .A(A[272]), .B(n1617), .Z(O[272]) );
  AND U2426 ( .A(S), .B(n1618), .Z(n1617) );
  XOR U2427 ( .A(B[272]), .B(A[272]), .Z(n1618) );
  XOR U2428 ( .A(A[271]), .B(n1619), .Z(O[271]) );
  AND U2429 ( .A(S), .B(n1620), .Z(n1619) );
  XOR U2430 ( .A(B[271]), .B(A[271]), .Z(n1620) );
  XOR U2431 ( .A(A[270]), .B(n1621), .Z(O[270]) );
  AND U2432 ( .A(S), .B(n1622), .Z(n1621) );
  XOR U2433 ( .A(B[270]), .B(A[270]), .Z(n1622) );
  XOR U2434 ( .A(A[26]), .B(n1623), .Z(O[26]) );
  AND U2435 ( .A(S), .B(n1624), .Z(n1623) );
  XOR U2436 ( .A(B[26]), .B(A[26]), .Z(n1624) );
  XOR U2437 ( .A(A[269]), .B(n1625), .Z(O[269]) );
  AND U2438 ( .A(S), .B(n1626), .Z(n1625) );
  XOR U2439 ( .A(B[269]), .B(A[269]), .Z(n1626) );
  XOR U2440 ( .A(A[268]), .B(n1627), .Z(O[268]) );
  AND U2441 ( .A(S), .B(n1628), .Z(n1627) );
  XOR U2442 ( .A(B[268]), .B(A[268]), .Z(n1628) );
  XOR U2443 ( .A(A[267]), .B(n1629), .Z(O[267]) );
  AND U2444 ( .A(S), .B(n1630), .Z(n1629) );
  XOR U2445 ( .A(B[267]), .B(A[267]), .Z(n1630) );
  XOR U2446 ( .A(A[266]), .B(n1631), .Z(O[266]) );
  AND U2447 ( .A(S), .B(n1632), .Z(n1631) );
  XOR U2448 ( .A(B[266]), .B(A[266]), .Z(n1632) );
  XOR U2449 ( .A(A[265]), .B(n1633), .Z(O[265]) );
  AND U2450 ( .A(S), .B(n1634), .Z(n1633) );
  XOR U2451 ( .A(B[265]), .B(A[265]), .Z(n1634) );
  XOR U2452 ( .A(A[264]), .B(n1635), .Z(O[264]) );
  AND U2453 ( .A(S), .B(n1636), .Z(n1635) );
  XOR U2454 ( .A(B[264]), .B(A[264]), .Z(n1636) );
  XOR U2455 ( .A(A[263]), .B(n1637), .Z(O[263]) );
  AND U2456 ( .A(S), .B(n1638), .Z(n1637) );
  XOR U2457 ( .A(B[263]), .B(A[263]), .Z(n1638) );
  XOR U2458 ( .A(A[262]), .B(n1639), .Z(O[262]) );
  AND U2459 ( .A(S), .B(n1640), .Z(n1639) );
  XOR U2460 ( .A(B[262]), .B(A[262]), .Z(n1640) );
  XOR U2461 ( .A(A[261]), .B(n1641), .Z(O[261]) );
  AND U2462 ( .A(S), .B(n1642), .Z(n1641) );
  XOR U2463 ( .A(B[261]), .B(A[261]), .Z(n1642) );
  XOR U2464 ( .A(A[260]), .B(n1643), .Z(O[260]) );
  AND U2465 ( .A(S), .B(n1644), .Z(n1643) );
  XOR U2466 ( .A(B[260]), .B(A[260]), .Z(n1644) );
  XOR U2467 ( .A(A[25]), .B(n1645), .Z(O[25]) );
  AND U2468 ( .A(S), .B(n1646), .Z(n1645) );
  XOR U2469 ( .A(B[25]), .B(A[25]), .Z(n1646) );
  XOR U2470 ( .A(A[259]), .B(n1647), .Z(O[259]) );
  AND U2471 ( .A(S), .B(n1648), .Z(n1647) );
  XOR U2472 ( .A(B[259]), .B(A[259]), .Z(n1648) );
  XOR U2473 ( .A(A[258]), .B(n1649), .Z(O[258]) );
  AND U2474 ( .A(S), .B(n1650), .Z(n1649) );
  XOR U2475 ( .A(B[258]), .B(A[258]), .Z(n1650) );
  XOR U2476 ( .A(A[257]), .B(n1651), .Z(O[257]) );
  AND U2477 ( .A(S), .B(n1652), .Z(n1651) );
  XOR U2478 ( .A(B[257]), .B(A[257]), .Z(n1652) );
  XOR U2479 ( .A(A[256]), .B(n1653), .Z(O[256]) );
  AND U2480 ( .A(S), .B(n1654), .Z(n1653) );
  XOR U2481 ( .A(B[256]), .B(A[256]), .Z(n1654) );
  XOR U2482 ( .A(A[255]), .B(n1655), .Z(O[255]) );
  AND U2483 ( .A(S), .B(n1656), .Z(n1655) );
  XOR U2484 ( .A(B[255]), .B(A[255]), .Z(n1656) );
  XOR U2485 ( .A(A[254]), .B(n1657), .Z(O[254]) );
  AND U2486 ( .A(S), .B(n1658), .Z(n1657) );
  XOR U2487 ( .A(B[254]), .B(A[254]), .Z(n1658) );
  XOR U2488 ( .A(A[253]), .B(n1659), .Z(O[253]) );
  AND U2489 ( .A(S), .B(n1660), .Z(n1659) );
  XOR U2490 ( .A(B[253]), .B(A[253]), .Z(n1660) );
  XOR U2491 ( .A(A[252]), .B(n1661), .Z(O[252]) );
  AND U2492 ( .A(S), .B(n1662), .Z(n1661) );
  XOR U2493 ( .A(B[252]), .B(A[252]), .Z(n1662) );
  XOR U2494 ( .A(A[251]), .B(n1663), .Z(O[251]) );
  AND U2495 ( .A(S), .B(n1664), .Z(n1663) );
  XOR U2496 ( .A(B[251]), .B(A[251]), .Z(n1664) );
  XOR U2497 ( .A(A[250]), .B(n1665), .Z(O[250]) );
  AND U2498 ( .A(S), .B(n1666), .Z(n1665) );
  XOR U2499 ( .A(B[250]), .B(A[250]), .Z(n1666) );
  XOR U2500 ( .A(A[24]), .B(n1667), .Z(O[24]) );
  AND U2501 ( .A(S), .B(n1668), .Z(n1667) );
  XOR U2502 ( .A(B[24]), .B(A[24]), .Z(n1668) );
  XOR U2503 ( .A(A[249]), .B(n1669), .Z(O[249]) );
  AND U2504 ( .A(S), .B(n1670), .Z(n1669) );
  XOR U2505 ( .A(B[249]), .B(A[249]), .Z(n1670) );
  XOR U2506 ( .A(A[248]), .B(n1671), .Z(O[248]) );
  AND U2507 ( .A(S), .B(n1672), .Z(n1671) );
  XOR U2508 ( .A(B[248]), .B(A[248]), .Z(n1672) );
  XOR U2509 ( .A(A[247]), .B(n1673), .Z(O[247]) );
  AND U2510 ( .A(S), .B(n1674), .Z(n1673) );
  XOR U2511 ( .A(B[247]), .B(A[247]), .Z(n1674) );
  XOR U2512 ( .A(A[246]), .B(n1675), .Z(O[246]) );
  AND U2513 ( .A(S), .B(n1676), .Z(n1675) );
  XOR U2514 ( .A(B[246]), .B(A[246]), .Z(n1676) );
  XOR U2515 ( .A(A[245]), .B(n1677), .Z(O[245]) );
  AND U2516 ( .A(S), .B(n1678), .Z(n1677) );
  XOR U2517 ( .A(B[245]), .B(A[245]), .Z(n1678) );
  XOR U2518 ( .A(A[244]), .B(n1679), .Z(O[244]) );
  AND U2519 ( .A(S), .B(n1680), .Z(n1679) );
  XOR U2520 ( .A(B[244]), .B(A[244]), .Z(n1680) );
  XOR U2521 ( .A(A[243]), .B(n1681), .Z(O[243]) );
  AND U2522 ( .A(S), .B(n1682), .Z(n1681) );
  XOR U2523 ( .A(B[243]), .B(A[243]), .Z(n1682) );
  XOR U2524 ( .A(A[242]), .B(n1683), .Z(O[242]) );
  AND U2525 ( .A(S), .B(n1684), .Z(n1683) );
  XOR U2526 ( .A(B[242]), .B(A[242]), .Z(n1684) );
  XOR U2527 ( .A(A[241]), .B(n1685), .Z(O[241]) );
  AND U2528 ( .A(S), .B(n1686), .Z(n1685) );
  XOR U2529 ( .A(B[241]), .B(A[241]), .Z(n1686) );
  XOR U2530 ( .A(A[240]), .B(n1687), .Z(O[240]) );
  AND U2531 ( .A(S), .B(n1688), .Z(n1687) );
  XOR U2532 ( .A(B[240]), .B(A[240]), .Z(n1688) );
  XOR U2533 ( .A(A[23]), .B(n1689), .Z(O[23]) );
  AND U2534 ( .A(S), .B(n1690), .Z(n1689) );
  XOR U2535 ( .A(B[23]), .B(A[23]), .Z(n1690) );
  XOR U2536 ( .A(A[239]), .B(n1691), .Z(O[239]) );
  AND U2537 ( .A(S), .B(n1692), .Z(n1691) );
  XOR U2538 ( .A(B[239]), .B(A[239]), .Z(n1692) );
  XOR U2539 ( .A(A[238]), .B(n1693), .Z(O[238]) );
  AND U2540 ( .A(S), .B(n1694), .Z(n1693) );
  XOR U2541 ( .A(B[238]), .B(A[238]), .Z(n1694) );
  XOR U2542 ( .A(A[237]), .B(n1695), .Z(O[237]) );
  AND U2543 ( .A(S), .B(n1696), .Z(n1695) );
  XOR U2544 ( .A(B[237]), .B(A[237]), .Z(n1696) );
  XOR U2545 ( .A(A[236]), .B(n1697), .Z(O[236]) );
  AND U2546 ( .A(S), .B(n1698), .Z(n1697) );
  XOR U2547 ( .A(B[236]), .B(A[236]), .Z(n1698) );
  XOR U2548 ( .A(A[235]), .B(n1699), .Z(O[235]) );
  AND U2549 ( .A(S), .B(n1700), .Z(n1699) );
  XOR U2550 ( .A(B[235]), .B(A[235]), .Z(n1700) );
  XOR U2551 ( .A(A[234]), .B(n1701), .Z(O[234]) );
  AND U2552 ( .A(S), .B(n1702), .Z(n1701) );
  XOR U2553 ( .A(B[234]), .B(A[234]), .Z(n1702) );
  XOR U2554 ( .A(A[233]), .B(n1703), .Z(O[233]) );
  AND U2555 ( .A(S), .B(n1704), .Z(n1703) );
  XOR U2556 ( .A(B[233]), .B(A[233]), .Z(n1704) );
  XOR U2557 ( .A(A[232]), .B(n1705), .Z(O[232]) );
  AND U2558 ( .A(S), .B(n1706), .Z(n1705) );
  XOR U2559 ( .A(B[232]), .B(A[232]), .Z(n1706) );
  XOR U2560 ( .A(A[231]), .B(n1707), .Z(O[231]) );
  AND U2561 ( .A(S), .B(n1708), .Z(n1707) );
  XOR U2562 ( .A(B[231]), .B(A[231]), .Z(n1708) );
  XOR U2563 ( .A(A[230]), .B(n1709), .Z(O[230]) );
  AND U2564 ( .A(S), .B(n1710), .Z(n1709) );
  XOR U2565 ( .A(B[230]), .B(A[230]), .Z(n1710) );
  XOR U2566 ( .A(A[22]), .B(n1711), .Z(O[22]) );
  AND U2567 ( .A(S), .B(n1712), .Z(n1711) );
  XOR U2568 ( .A(B[22]), .B(A[22]), .Z(n1712) );
  XOR U2569 ( .A(A[229]), .B(n1713), .Z(O[229]) );
  AND U2570 ( .A(S), .B(n1714), .Z(n1713) );
  XOR U2571 ( .A(B[229]), .B(A[229]), .Z(n1714) );
  XOR U2572 ( .A(A[228]), .B(n1715), .Z(O[228]) );
  AND U2573 ( .A(S), .B(n1716), .Z(n1715) );
  XOR U2574 ( .A(B[228]), .B(A[228]), .Z(n1716) );
  XOR U2575 ( .A(A[227]), .B(n1717), .Z(O[227]) );
  AND U2576 ( .A(S), .B(n1718), .Z(n1717) );
  XOR U2577 ( .A(B[227]), .B(A[227]), .Z(n1718) );
  XOR U2578 ( .A(A[226]), .B(n1719), .Z(O[226]) );
  AND U2579 ( .A(S), .B(n1720), .Z(n1719) );
  XOR U2580 ( .A(B[226]), .B(A[226]), .Z(n1720) );
  XOR U2581 ( .A(A[225]), .B(n1721), .Z(O[225]) );
  AND U2582 ( .A(S), .B(n1722), .Z(n1721) );
  XOR U2583 ( .A(B[225]), .B(A[225]), .Z(n1722) );
  XOR U2584 ( .A(A[224]), .B(n1723), .Z(O[224]) );
  AND U2585 ( .A(S), .B(n1724), .Z(n1723) );
  XOR U2586 ( .A(B[224]), .B(A[224]), .Z(n1724) );
  XOR U2587 ( .A(A[223]), .B(n1725), .Z(O[223]) );
  AND U2588 ( .A(S), .B(n1726), .Z(n1725) );
  XOR U2589 ( .A(B[223]), .B(A[223]), .Z(n1726) );
  XOR U2590 ( .A(A[222]), .B(n1727), .Z(O[222]) );
  AND U2591 ( .A(S), .B(n1728), .Z(n1727) );
  XOR U2592 ( .A(B[222]), .B(A[222]), .Z(n1728) );
  XOR U2593 ( .A(A[221]), .B(n1729), .Z(O[221]) );
  AND U2594 ( .A(S), .B(n1730), .Z(n1729) );
  XOR U2595 ( .A(B[221]), .B(A[221]), .Z(n1730) );
  XOR U2596 ( .A(A[220]), .B(n1731), .Z(O[220]) );
  AND U2597 ( .A(S), .B(n1732), .Z(n1731) );
  XOR U2598 ( .A(B[220]), .B(A[220]), .Z(n1732) );
  XOR U2599 ( .A(A[21]), .B(n1733), .Z(O[21]) );
  AND U2600 ( .A(S), .B(n1734), .Z(n1733) );
  XOR U2601 ( .A(B[21]), .B(A[21]), .Z(n1734) );
  XOR U2602 ( .A(A[219]), .B(n1735), .Z(O[219]) );
  AND U2603 ( .A(S), .B(n1736), .Z(n1735) );
  XOR U2604 ( .A(B[219]), .B(A[219]), .Z(n1736) );
  XOR U2605 ( .A(A[218]), .B(n1737), .Z(O[218]) );
  AND U2606 ( .A(S), .B(n1738), .Z(n1737) );
  XOR U2607 ( .A(B[218]), .B(A[218]), .Z(n1738) );
  XOR U2608 ( .A(A[217]), .B(n1739), .Z(O[217]) );
  AND U2609 ( .A(S), .B(n1740), .Z(n1739) );
  XOR U2610 ( .A(B[217]), .B(A[217]), .Z(n1740) );
  XOR U2611 ( .A(A[216]), .B(n1741), .Z(O[216]) );
  AND U2612 ( .A(S), .B(n1742), .Z(n1741) );
  XOR U2613 ( .A(B[216]), .B(A[216]), .Z(n1742) );
  XOR U2614 ( .A(A[215]), .B(n1743), .Z(O[215]) );
  AND U2615 ( .A(S), .B(n1744), .Z(n1743) );
  XOR U2616 ( .A(B[215]), .B(A[215]), .Z(n1744) );
  XOR U2617 ( .A(A[214]), .B(n1745), .Z(O[214]) );
  AND U2618 ( .A(S), .B(n1746), .Z(n1745) );
  XOR U2619 ( .A(B[214]), .B(A[214]), .Z(n1746) );
  XOR U2620 ( .A(A[213]), .B(n1747), .Z(O[213]) );
  AND U2621 ( .A(S), .B(n1748), .Z(n1747) );
  XOR U2622 ( .A(B[213]), .B(A[213]), .Z(n1748) );
  XOR U2623 ( .A(A[212]), .B(n1749), .Z(O[212]) );
  AND U2624 ( .A(S), .B(n1750), .Z(n1749) );
  XOR U2625 ( .A(B[212]), .B(A[212]), .Z(n1750) );
  XOR U2626 ( .A(A[211]), .B(n1751), .Z(O[211]) );
  AND U2627 ( .A(S), .B(n1752), .Z(n1751) );
  XOR U2628 ( .A(B[211]), .B(A[211]), .Z(n1752) );
  XOR U2629 ( .A(A[210]), .B(n1753), .Z(O[210]) );
  AND U2630 ( .A(S), .B(n1754), .Z(n1753) );
  XOR U2631 ( .A(B[210]), .B(A[210]), .Z(n1754) );
  XOR U2632 ( .A(A[20]), .B(n1755), .Z(O[20]) );
  AND U2633 ( .A(S), .B(n1756), .Z(n1755) );
  XOR U2634 ( .A(B[20]), .B(A[20]), .Z(n1756) );
  XOR U2635 ( .A(A[209]), .B(n1757), .Z(O[209]) );
  AND U2636 ( .A(S), .B(n1758), .Z(n1757) );
  XOR U2637 ( .A(B[209]), .B(A[209]), .Z(n1758) );
  XOR U2638 ( .A(A[208]), .B(n1759), .Z(O[208]) );
  AND U2639 ( .A(S), .B(n1760), .Z(n1759) );
  XOR U2640 ( .A(B[208]), .B(A[208]), .Z(n1760) );
  XOR U2641 ( .A(A[207]), .B(n1761), .Z(O[207]) );
  AND U2642 ( .A(S), .B(n1762), .Z(n1761) );
  XOR U2643 ( .A(B[207]), .B(A[207]), .Z(n1762) );
  XOR U2644 ( .A(A[206]), .B(n1763), .Z(O[206]) );
  AND U2645 ( .A(S), .B(n1764), .Z(n1763) );
  XOR U2646 ( .A(B[206]), .B(A[206]), .Z(n1764) );
  XOR U2647 ( .A(A[205]), .B(n1765), .Z(O[205]) );
  AND U2648 ( .A(S), .B(n1766), .Z(n1765) );
  XOR U2649 ( .A(B[205]), .B(A[205]), .Z(n1766) );
  XOR U2650 ( .A(A[204]), .B(n1767), .Z(O[204]) );
  AND U2651 ( .A(S), .B(n1768), .Z(n1767) );
  XOR U2652 ( .A(B[204]), .B(A[204]), .Z(n1768) );
  XOR U2653 ( .A(A[203]), .B(n1769), .Z(O[203]) );
  AND U2654 ( .A(S), .B(n1770), .Z(n1769) );
  XOR U2655 ( .A(B[203]), .B(A[203]), .Z(n1770) );
  XOR U2656 ( .A(A[202]), .B(n1771), .Z(O[202]) );
  AND U2657 ( .A(S), .B(n1772), .Z(n1771) );
  XOR U2658 ( .A(B[202]), .B(A[202]), .Z(n1772) );
  XOR U2659 ( .A(A[201]), .B(n1773), .Z(O[201]) );
  AND U2660 ( .A(S), .B(n1774), .Z(n1773) );
  XOR U2661 ( .A(B[201]), .B(A[201]), .Z(n1774) );
  XOR U2662 ( .A(A[200]), .B(n1775), .Z(O[200]) );
  AND U2663 ( .A(S), .B(n1776), .Z(n1775) );
  XOR U2664 ( .A(B[200]), .B(A[200]), .Z(n1776) );
  XOR U2665 ( .A(A[1]), .B(n1777), .Z(O[1]) );
  AND U2666 ( .A(S), .B(n1778), .Z(n1777) );
  XOR U2667 ( .A(B[1]), .B(A[1]), .Z(n1778) );
  XOR U2668 ( .A(A[19]), .B(n1779), .Z(O[19]) );
  AND U2669 ( .A(S), .B(n1780), .Z(n1779) );
  XOR U2670 ( .A(B[19]), .B(A[19]), .Z(n1780) );
  XOR U2671 ( .A(A[199]), .B(n1781), .Z(O[199]) );
  AND U2672 ( .A(S), .B(n1782), .Z(n1781) );
  XOR U2673 ( .A(B[199]), .B(A[199]), .Z(n1782) );
  XOR U2674 ( .A(A[198]), .B(n1783), .Z(O[198]) );
  AND U2675 ( .A(S), .B(n1784), .Z(n1783) );
  XOR U2676 ( .A(B[198]), .B(A[198]), .Z(n1784) );
  XOR U2677 ( .A(A[197]), .B(n1785), .Z(O[197]) );
  AND U2678 ( .A(S), .B(n1786), .Z(n1785) );
  XOR U2679 ( .A(B[197]), .B(A[197]), .Z(n1786) );
  XOR U2680 ( .A(A[196]), .B(n1787), .Z(O[196]) );
  AND U2681 ( .A(S), .B(n1788), .Z(n1787) );
  XOR U2682 ( .A(B[196]), .B(A[196]), .Z(n1788) );
  XOR U2683 ( .A(A[195]), .B(n1789), .Z(O[195]) );
  AND U2684 ( .A(S), .B(n1790), .Z(n1789) );
  XOR U2685 ( .A(B[195]), .B(A[195]), .Z(n1790) );
  XOR U2686 ( .A(A[194]), .B(n1791), .Z(O[194]) );
  AND U2687 ( .A(S), .B(n1792), .Z(n1791) );
  XOR U2688 ( .A(B[194]), .B(A[194]), .Z(n1792) );
  XOR U2689 ( .A(A[193]), .B(n1793), .Z(O[193]) );
  AND U2690 ( .A(S), .B(n1794), .Z(n1793) );
  XOR U2691 ( .A(B[193]), .B(A[193]), .Z(n1794) );
  XOR U2692 ( .A(A[192]), .B(n1795), .Z(O[192]) );
  AND U2693 ( .A(S), .B(n1796), .Z(n1795) );
  XOR U2694 ( .A(B[192]), .B(A[192]), .Z(n1796) );
  XOR U2695 ( .A(A[191]), .B(n1797), .Z(O[191]) );
  AND U2696 ( .A(S), .B(n1798), .Z(n1797) );
  XOR U2697 ( .A(B[191]), .B(A[191]), .Z(n1798) );
  XOR U2698 ( .A(A[190]), .B(n1799), .Z(O[190]) );
  AND U2699 ( .A(S), .B(n1800), .Z(n1799) );
  XOR U2700 ( .A(B[190]), .B(A[190]), .Z(n1800) );
  XOR U2701 ( .A(A[18]), .B(n1801), .Z(O[18]) );
  AND U2702 ( .A(S), .B(n1802), .Z(n1801) );
  XOR U2703 ( .A(B[18]), .B(A[18]), .Z(n1802) );
  XOR U2704 ( .A(A[189]), .B(n1803), .Z(O[189]) );
  AND U2705 ( .A(S), .B(n1804), .Z(n1803) );
  XOR U2706 ( .A(B[189]), .B(A[189]), .Z(n1804) );
  XOR U2707 ( .A(A[188]), .B(n1805), .Z(O[188]) );
  AND U2708 ( .A(S), .B(n1806), .Z(n1805) );
  XOR U2709 ( .A(B[188]), .B(A[188]), .Z(n1806) );
  XOR U2710 ( .A(A[187]), .B(n1807), .Z(O[187]) );
  AND U2711 ( .A(S), .B(n1808), .Z(n1807) );
  XOR U2712 ( .A(B[187]), .B(A[187]), .Z(n1808) );
  XOR U2713 ( .A(A[186]), .B(n1809), .Z(O[186]) );
  AND U2714 ( .A(S), .B(n1810), .Z(n1809) );
  XOR U2715 ( .A(B[186]), .B(A[186]), .Z(n1810) );
  XOR U2716 ( .A(A[185]), .B(n1811), .Z(O[185]) );
  AND U2717 ( .A(S), .B(n1812), .Z(n1811) );
  XOR U2718 ( .A(B[185]), .B(A[185]), .Z(n1812) );
  XOR U2719 ( .A(A[184]), .B(n1813), .Z(O[184]) );
  AND U2720 ( .A(S), .B(n1814), .Z(n1813) );
  XOR U2721 ( .A(B[184]), .B(A[184]), .Z(n1814) );
  XOR U2722 ( .A(A[183]), .B(n1815), .Z(O[183]) );
  AND U2723 ( .A(S), .B(n1816), .Z(n1815) );
  XOR U2724 ( .A(B[183]), .B(A[183]), .Z(n1816) );
  XOR U2725 ( .A(A[182]), .B(n1817), .Z(O[182]) );
  AND U2726 ( .A(S), .B(n1818), .Z(n1817) );
  XOR U2727 ( .A(B[182]), .B(A[182]), .Z(n1818) );
  XOR U2728 ( .A(A[181]), .B(n1819), .Z(O[181]) );
  AND U2729 ( .A(S), .B(n1820), .Z(n1819) );
  XOR U2730 ( .A(B[181]), .B(A[181]), .Z(n1820) );
  XOR U2731 ( .A(A[180]), .B(n1821), .Z(O[180]) );
  AND U2732 ( .A(S), .B(n1822), .Z(n1821) );
  XOR U2733 ( .A(B[180]), .B(A[180]), .Z(n1822) );
  XOR U2734 ( .A(A[17]), .B(n1823), .Z(O[17]) );
  AND U2735 ( .A(S), .B(n1824), .Z(n1823) );
  XOR U2736 ( .A(B[17]), .B(A[17]), .Z(n1824) );
  XOR U2737 ( .A(A[179]), .B(n1825), .Z(O[179]) );
  AND U2738 ( .A(S), .B(n1826), .Z(n1825) );
  XOR U2739 ( .A(B[179]), .B(A[179]), .Z(n1826) );
  XOR U2740 ( .A(A[178]), .B(n1827), .Z(O[178]) );
  AND U2741 ( .A(S), .B(n1828), .Z(n1827) );
  XOR U2742 ( .A(B[178]), .B(A[178]), .Z(n1828) );
  XOR U2743 ( .A(A[177]), .B(n1829), .Z(O[177]) );
  AND U2744 ( .A(S), .B(n1830), .Z(n1829) );
  XOR U2745 ( .A(B[177]), .B(A[177]), .Z(n1830) );
  XOR U2746 ( .A(A[176]), .B(n1831), .Z(O[176]) );
  AND U2747 ( .A(S), .B(n1832), .Z(n1831) );
  XOR U2748 ( .A(B[176]), .B(A[176]), .Z(n1832) );
  XOR U2749 ( .A(A[175]), .B(n1833), .Z(O[175]) );
  AND U2750 ( .A(S), .B(n1834), .Z(n1833) );
  XOR U2751 ( .A(B[175]), .B(A[175]), .Z(n1834) );
  XOR U2752 ( .A(A[174]), .B(n1835), .Z(O[174]) );
  AND U2753 ( .A(S), .B(n1836), .Z(n1835) );
  XOR U2754 ( .A(B[174]), .B(A[174]), .Z(n1836) );
  XOR U2755 ( .A(A[173]), .B(n1837), .Z(O[173]) );
  AND U2756 ( .A(S), .B(n1838), .Z(n1837) );
  XOR U2757 ( .A(B[173]), .B(A[173]), .Z(n1838) );
  XOR U2758 ( .A(A[172]), .B(n1839), .Z(O[172]) );
  AND U2759 ( .A(S), .B(n1840), .Z(n1839) );
  XOR U2760 ( .A(B[172]), .B(A[172]), .Z(n1840) );
  XOR U2761 ( .A(A[171]), .B(n1841), .Z(O[171]) );
  AND U2762 ( .A(S), .B(n1842), .Z(n1841) );
  XOR U2763 ( .A(B[171]), .B(A[171]), .Z(n1842) );
  XOR U2764 ( .A(A[170]), .B(n1843), .Z(O[170]) );
  AND U2765 ( .A(S), .B(n1844), .Z(n1843) );
  XOR U2766 ( .A(B[170]), .B(A[170]), .Z(n1844) );
  XOR U2767 ( .A(A[16]), .B(n1845), .Z(O[16]) );
  AND U2768 ( .A(S), .B(n1846), .Z(n1845) );
  XOR U2769 ( .A(B[16]), .B(A[16]), .Z(n1846) );
  XOR U2770 ( .A(A[169]), .B(n1847), .Z(O[169]) );
  AND U2771 ( .A(S), .B(n1848), .Z(n1847) );
  XOR U2772 ( .A(B[169]), .B(A[169]), .Z(n1848) );
  XOR U2773 ( .A(A[168]), .B(n1849), .Z(O[168]) );
  AND U2774 ( .A(S), .B(n1850), .Z(n1849) );
  XOR U2775 ( .A(B[168]), .B(A[168]), .Z(n1850) );
  XOR U2776 ( .A(A[167]), .B(n1851), .Z(O[167]) );
  AND U2777 ( .A(S), .B(n1852), .Z(n1851) );
  XOR U2778 ( .A(B[167]), .B(A[167]), .Z(n1852) );
  XOR U2779 ( .A(A[166]), .B(n1853), .Z(O[166]) );
  AND U2780 ( .A(S), .B(n1854), .Z(n1853) );
  XOR U2781 ( .A(B[166]), .B(A[166]), .Z(n1854) );
  XOR U2782 ( .A(A[165]), .B(n1855), .Z(O[165]) );
  AND U2783 ( .A(S), .B(n1856), .Z(n1855) );
  XOR U2784 ( .A(B[165]), .B(A[165]), .Z(n1856) );
  XOR U2785 ( .A(A[164]), .B(n1857), .Z(O[164]) );
  AND U2786 ( .A(S), .B(n1858), .Z(n1857) );
  XOR U2787 ( .A(B[164]), .B(A[164]), .Z(n1858) );
  XOR U2788 ( .A(A[163]), .B(n1859), .Z(O[163]) );
  AND U2789 ( .A(S), .B(n1860), .Z(n1859) );
  XOR U2790 ( .A(B[163]), .B(A[163]), .Z(n1860) );
  XOR U2791 ( .A(A[162]), .B(n1861), .Z(O[162]) );
  AND U2792 ( .A(S), .B(n1862), .Z(n1861) );
  XOR U2793 ( .A(B[162]), .B(A[162]), .Z(n1862) );
  XOR U2794 ( .A(A[161]), .B(n1863), .Z(O[161]) );
  AND U2795 ( .A(S), .B(n1864), .Z(n1863) );
  XOR U2796 ( .A(B[161]), .B(A[161]), .Z(n1864) );
  XOR U2797 ( .A(A[160]), .B(n1865), .Z(O[160]) );
  AND U2798 ( .A(S), .B(n1866), .Z(n1865) );
  XOR U2799 ( .A(B[160]), .B(A[160]), .Z(n1866) );
  XOR U2800 ( .A(A[15]), .B(n1867), .Z(O[15]) );
  AND U2801 ( .A(S), .B(n1868), .Z(n1867) );
  XOR U2802 ( .A(B[15]), .B(A[15]), .Z(n1868) );
  XOR U2803 ( .A(A[159]), .B(n1869), .Z(O[159]) );
  AND U2804 ( .A(S), .B(n1870), .Z(n1869) );
  XOR U2805 ( .A(B[159]), .B(A[159]), .Z(n1870) );
  XOR U2806 ( .A(A[158]), .B(n1871), .Z(O[158]) );
  AND U2807 ( .A(S), .B(n1872), .Z(n1871) );
  XOR U2808 ( .A(B[158]), .B(A[158]), .Z(n1872) );
  XOR U2809 ( .A(A[157]), .B(n1873), .Z(O[157]) );
  AND U2810 ( .A(S), .B(n1874), .Z(n1873) );
  XOR U2811 ( .A(B[157]), .B(A[157]), .Z(n1874) );
  XOR U2812 ( .A(A[156]), .B(n1875), .Z(O[156]) );
  AND U2813 ( .A(S), .B(n1876), .Z(n1875) );
  XOR U2814 ( .A(B[156]), .B(A[156]), .Z(n1876) );
  XOR U2815 ( .A(A[155]), .B(n1877), .Z(O[155]) );
  AND U2816 ( .A(S), .B(n1878), .Z(n1877) );
  XOR U2817 ( .A(B[155]), .B(A[155]), .Z(n1878) );
  XOR U2818 ( .A(A[154]), .B(n1879), .Z(O[154]) );
  AND U2819 ( .A(S), .B(n1880), .Z(n1879) );
  XOR U2820 ( .A(B[154]), .B(A[154]), .Z(n1880) );
  XOR U2821 ( .A(A[153]), .B(n1881), .Z(O[153]) );
  AND U2822 ( .A(S), .B(n1882), .Z(n1881) );
  XOR U2823 ( .A(B[153]), .B(A[153]), .Z(n1882) );
  XOR U2824 ( .A(A[152]), .B(n1883), .Z(O[152]) );
  AND U2825 ( .A(S), .B(n1884), .Z(n1883) );
  XOR U2826 ( .A(B[152]), .B(A[152]), .Z(n1884) );
  XOR U2827 ( .A(A[151]), .B(n1885), .Z(O[151]) );
  AND U2828 ( .A(S), .B(n1886), .Z(n1885) );
  XOR U2829 ( .A(B[151]), .B(A[151]), .Z(n1886) );
  XOR U2830 ( .A(A[150]), .B(n1887), .Z(O[150]) );
  AND U2831 ( .A(S), .B(n1888), .Z(n1887) );
  XOR U2832 ( .A(B[150]), .B(A[150]), .Z(n1888) );
  XOR U2833 ( .A(A[14]), .B(n1889), .Z(O[14]) );
  AND U2834 ( .A(S), .B(n1890), .Z(n1889) );
  XOR U2835 ( .A(B[14]), .B(A[14]), .Z(n1890) );
  XOR U2836 ( .A(A[149]), .B(n1891), .Z(O[149]) );
  AND U2837 ( .A(S), .B(n1892), .Z(n1891) );
  XOR U2838 ( .A(B[149]), .B(A[149]), .Z(n1892) );
  XOR U2839 ( .A(A[148]), .B(n1893), .Z(O[148]) );
  AND U2840 ( .A(S), .B(n1894), .Z(n1893) );
  XOR U2841 ( .A(B[148]), .B(A[148]), .Z(n1894) );
  XOR U2842 ( .A(A[147]), .B(n1895), .Z(O[147]) );
  AND U2843 ( .A(S), .B(n1896), .Z(n1895) );
  XOR U2844 ( .A(B[147]), .B(A[147]), .Z(n1896) );
  XOR U2845 ( .A(A[146]), .B(n1897), .Z(O[146]) );
  AND U2846 ( .A(S), .B(n1898), .Z(n1897) );
  XOR U2847 ( .A(B[146]), .B(A[146]), .Z(n1898) );
  XOR U2848 ( .A(A[145]), .B(n1899), .Z(O[145]) );
  AND U2849 ( .A(S), .B(n1900), .Z(n1899) );
  XOR U2850 ( .A(B[145]), .B(A[145]), .Z(n1900) );
  XOR U2851 ( .A(A[144]), .B(n1901), .Z(O[144]) );
  AND U2852 ( .A(S), .B(n1902), .Z(n1901) );
  XOR U2853 ( .A(B[144]), .B(A[144]), .Z(n1902) );
  XOR U2854 ( .A(A[143]), .B(n1903), .Z(O[143]) );
  AND U2855 ( .A(S), .B(n1904), .Z(n1903) );
  XOR U2856 ( .A(B[143]), .B(A[143]), .Z(n1904) );
  XOR U2857 ( .A(A[142]), .B(n1905), .Z(O[142]) );
  AND U2858 ( .A(S), .B(n1906), .Z(n1905) );
  XOR U2859 ( .A(B[142]), .B(A[142]), .Z(n1906) );
  XOR U2860 ( .A(A[141]), .B(n1907), .Z(O[141]) );
  AND U2861 ( .A(S), .B(n1908), .Z(n1907) );
  XOR U2862 ( .A(B[141]), .B(A[141]), .Z(n1908) );
  XOR U2863 ( .A(A[140]), .B(n1909), .Z(O[140]) );
  AND U2864 ( .A(S), .B(n1910), .Z(n1909) );
  XOR U2865 ( .A(B[140]), .B(A[140]), .Z(n1910) );
  XOR U2866 ( .A(A[13]), .B(n1911), .Z(O[13]) );
  AND U2867 ( .A(S), .B(n1912), .Z(n1911) );
  XOR U2868 ( .A(B[13]), .B(A[13]), .Z(n1912) );
  XOR U2869 ( .A(A[139]), .B(n1913), .Z(O[139]) );
  AND U2870 ( .A(S), .B(n1914), .Z(n1913) );
  XOR U2871 ( .A(B[139]), .B(A[139]), .Z(n1914) );
  XOR U2872 ( .A(A[138]), .B(n1915), .Z(O[138]) );
  AND U2873 ( .A(S), .B(n1916), .Z(n1915) );
  XOR U2874 ( .A(B[138]), .B(A[138]), .Z(n1916) );
  XOR U2875 ( .A(A[137]), .B(n1917), .Z(O[137]) );
  AND U2876 ( .A(S), .B(n1918), .Z(n1917) );
  XOR U2877 ( .A(B[137]), .B(A[137]), .Z(n1918) );
  XOR U2878 ( .A(A[136]), .B(n1919), .Z(O[136]) );
  AND U2879 ( .A(S), .B(n1920), .Z(n1919) );
  XOR U2880 ( .A(B[136]), .B(A[136]), .Z(n1920) );
  XOR U2881 ( .A(A[135]), .B(n1921), .Z(O[135]) );
  AND U2882 ( .A(S), .B(n1922), .Z(n1921) );
  XOR U2883 ( .A(B[135]), .B(A[135]), .Z(n1922) );
  XOR U2884 ( .A(A[134]), .B(n1923), .Z(O[134]) );
  AND U2885 ( .A(S), .B(n1924), .Z(n1923) );
  XOR U2886 ( .A(B[134]), .B(A[134]), .Z(n1924) );
  XOR U2887 ( .A(A[133]), .B(n1925), .Z(O[133]) );
  AND U2888 ( .A(S), .B(n1926), .Z(n1925) );
  XOR U2889 ( .A(B[133]), .B(A[133]), .Z(n1926) );
  XOR U2890 ( .A(A[132]), .B(n1927), .Z(O[132]) );
  AND U2891 ( .A(S), .B(n1928), .Z(n1927) );
  XOR U2892 ( .A(B[132]), .B(A[132]), .Z(n1928) );
  XOR U2893 ( .A(A[131]), .B(n1929), .Z(O[131]) );
  AND U2894 ( .A(S), .B(n1930), .Z(n1929) );
  XOR U2895 ( .A(B[131]), .B(A[131]), .Z(n1930) );
  XOR U2896 ( .A(A[130]), .B(n1931), .Z(O[130]) );
  AND U2897 ( .A(S), .B(n1932), .Z(n1931) );
  XOR U2898 ( .A(B[130]), .B(A[130]), .Z(n1932) );
  XOR U2899 ( .A(A[12]), .B(n1933), .Z(O[12]) );
  AND U2900 ( .A(S), .B(n1934), .Z(n1933) );
  XOR U2901 ( .A(B[12]), .B(A[12]), .Z(n1934) );
  XOR U2902 ( .A(A[129]), .B(n1935), .Z(O[129]) );
  AND U2903 ( .A(S), .B(n1936), .Z(n1935) );
  XOR U2904 ( .A(B[129]), .B(A[129]), .Z(n1936) );
  XOR U2905 ( .A(A[128]), .B(n1937), .Z(O[128]) );
  AND U2906 ( .A(S), .B(n1938), .Z(n1937) );
  XOR U2907 ( .A(B[128]), .B(A[128]), .Z(n1938) );
  XOR U2908 ( .A(A[127]), .B(n1939), .Z(O[127]) );
  AND U2909 ( .A(S), .B(n1940), .Z(n1939) );
  XOR U2910 ( .A(B[127]), .B(A[127]), .Z(n1940) );
  XOR U2911 ( .A(A[126]), .B(n1941), .Z(O[126]) );
  AND U2912 ( .A(S), .B(n1942), .Z(n1941) );
  XOR U2913 ( .A(B[126]), .B(A[126]), .Z(n1942) );
  XOR U2914 ( .A(A[125]), .B(n1943), .Z(O[125]) );
  AND U2915 ( .A(S), .B(n1944), .Z(n1943) );
  XOR U2916 ( .A(B[125]), .B(A[125]), .Z(n1944) );
  XOR U2917 ( .A(A[124]), .B(n1945), .Z(O[124]) );
  AND U2918 ( .A(S), .B(n1946), .Z(n1945) );
  XOR U2919 ( .A(B[124]), .B(A[124]), .Z(n1946) );
  XOR U2920 ( .A(A[123]), .B(n1947), .Z(O[123]) );
  AND U2921 ( .A(S), .B(n1948), .Z(n1947) );
  XOR U2922 ( .A(B[123]), .B(A[123]), .Z(n1948) );
  XOR U2923 ( .A(A[122]), .B(n1949), .Z(O[122]) );
  AND U2924 ( .A(S), .B(n1950), .Z(n1949) );
  XOR U2925 ( .A(B[122]), .B(A[122]), .Z(n1950) );
  XOR U2926 ( .A(A[121]), .B(n1951), .Z(O[121]) );
  AND U2927 ( .A(S), .B(n1952), .Z(n1951) );
  XOR U2928 ( .A(B[121]), .B(A[121]), .Z(n1952) );
  XOR U2929 ( .A(A[120]), .B(n1953), .Z(O[120]) );
  AND U2930 ( .A(S), .B(n1954), .Z(n1953) );
  XOR U2931 ( .A(B[120]), .B(A[120]), .Z(n1954) );
  XOR U2932 ( .A(A[11]), .B(n1955), .Z(O[11]) );
  AND U2933 ( .A(S), .B(n1956), .Z(n1955) );
  XOR U2934 ( .A(B[11]), .B(A[11]), .Z(n1956) );
  XOR U2935 ( .A(A[119]), .B(n1957), .Z(O[119]) );
  AND U2936 ( .A(S), .B(n1958), .Z(n1957) );
  XOR U2937 ( .A(B[119]), .B(A[119]), .Z(n1958) );
  XOR U2938 ( .A(A[118]), .B(n1959), .Z(O[118]) );
  AND U2939 ( .A(S), .B(n1960), .Z(n1959) );
  XOR U2940 ( .A(B[118]), .B(A[118]), .Z(n1960) );
  XOR U2941 ( .A(A[117]), .B(n1961), .Z(O[117]) );
  AND U2942 ( .A(S), .B(n1962), .Z(n1961) );
  XOR U2943 ( .A(B[117]), .B(A[117]), .Z(n1962) );
  XOR U2944 ( .A(A[116]), .B(n1963), .Z(O[116]) );
  AND U2945 ( .A(S), .B(n1964), .Z(n1963) );
  XOR U2946 ( .A(B[116]), .B(A[116]), .Z(n1964) );
  XOR U2947 ( .A(A[115]), .B(n1965), .Z(O[115]) );
  AND U2948 ( .A(S), .B(n1966), .Z(n1965) );
  XOR U2949 ( .A(B[115]), .B(A[115]), .Z(n1966) );
  XOR U2950 ( .A(A[114]), .B(n1967), .Z(O[114]) );
  AND U2951 ( .A(S), .B(n1968), .Z(n1967) );
  XOR U2952 ( .A(B[114]), .B(A[114]), .Z(n1968) );
  XOR U2953 ( .A(A[113]), .B(n1969), .Z(O[113]) );
  AND U2954 ( .A(S), .B(n1970), .Z(n1969) );
  XOR U2955 ( .A(B[113]), .B(A[113]), .Z(n1970) );
  XOR U2956 ( .A(A[112]), .B(n1971), .Z(O[112]) );
  AND U2957 ( .A(S), .B(n1972), .Z(n1971) );
  XOR U2958 ( .A(B[112]), .B(A[112]), .Z(n1972) );
  XOR U2959 ( .A(A[111]), .B(n1973), .Z(O[111]) );
  AND U2960 ( .A(S), .B(n1974), .Z(n1973) );
  XOR U2961 ( .A(B[111]), .B(A[111]), .Z(n1974) );
  XOR U2962 ( .A(A[110]), .B(n1975), .Z(O[110]) );
  AND U2963 ( .A(S), .B(n1976), .Z(n1975) );
  XOR U2964 ( .A(B[110]), .B(A[110]), .Z(n1976) );
  XOR U2965 ( .A(A[10]), .B(n1977), .Z(O[10]) );
  AND U2966 ( .A(S), .B(n1978), .Z(n1977) );
  XOR U2967 ( .A(B[10]), .B(A[10]), .Z(n1978) );
  XOR U2968 ( .A(A[109]), .B(n1979), .Z(O[109]) );
  AND U2969 ( .A(S), .B(n1980), .Z(n1979) );
  XOR U2970 ( .A(B[109]), .B(A[109]), .Z(n1980) );
  XOR U2971 ( .A(A[108]), .B(n1981), .Z(O[108]) );
  AND U2972 ( .A(S), .B(n1982), .Z(n1981) );
  XOR U2973 ( .A(B[108]), .B(A[108]), .Z(n1982) );
  XOR U2974 ( .A(A[107]), .B(n1983), .Z(O[107]) );
  AND U2975 ( .A(S), .B(n1984), .Z(n1983) );
  XOR U2976 ( .A(B[107]), .B(A[107]), .Z(n1984) );
  XOR U2977 ( .A(A[106]), .B(n1985), .Z(O[106]) );
  AND U2978 ( .A(S), .B(n1986), .Z(n1985) );
  XOR U2979 ( .A(B[106]), .B(A[106]), .Z(n1986) );
  XOR U2980 ( .A(A[105]), .B(n1987), .Z(O[105]) );
  AND U2981 ( .A(S), .B(n1988), .Z(n1987) );
  XOR U2982 ( .A(B[105]), .B(A[105]), .Z(n1988) );
  XOR U2983 ( .A(A[104]), .B(n1989), .Z(O[104]) );
  AND U2984 ( .A(S), .B(n1990), .Z(n1989) );
  XOR U2985 ( .A(B[104]), .B(A[104]), .Z(n1990) );
  XOR U2986 ( .A(A[103]), .B(n1991), .Z(O[103]) );
  AND U2987 ( .A(S), .B(n1992), .Z(n1991) );
  XOR U2988 ( .A(B[103]), .B(A[103]), .Z(n1992) );
  XOR U2989 ( .A(A[102]), .B(n1993), .Z(O[102]) );
  AND U2990 ( .A(S), .B(n1994), .Z(n1993) );
  XOR U2991 ( .A(B[102]), .B(A[102]), .Z(n1994) );
  XOR U2992 ( .A(A[1023]), .B(n1995), .Z(O[1023]) );
  AND U2993 ( .A(S), .B(n1996), .Z(n1995) );
  XOR U2994 ( .A(B[1023]), .B(A[1023]), .Z(n1996) );
  XOR U2995 ( .A(A[1022]), .B(n1997), .Z(O[1022]) );
  AND U2996 ( .A(S), .B(n1998), .Z(n1997) );
  XOR U2997 ( .A(B[1022]), .B(A[1022]), .Z(n1998) );
  XOR U2998 ( .A(A[1021]), .B(n1999), .Z(O[1021]) );
  AND U2999 ( .A(S), .B(n2000), .Z(n1999) );
  XOR U3000 ( .A(B[1021]), .B(A[1021]), .Z(n2000) );
  XOR U3001 ( .A(A[1020]), .B(n2001), .Z(O[1020]) );
  AND U3002 ( .A(S), .B(n2002), .Z(n2001) );
  XOR U3003 ( .A(B[1020]), .B(A[1020]), .Z(n2002) );
  XOR U3004 ( .A(A[101]), .B(n2003), .Z(O[101]) );
  AND U3005 ( .A(S), .B(n2004), .Z(n2003) );
  XOR U3006 ( .A(B[101]), .B(A[101]), .Z(n2004) );
  XOR U3007 ( .A(A[1019]), .B(n2005), .Z(O[1019]) );
  AND U3008 ( .A(S), .B(n2006), .Z(n2005) );
  XOR U3009 ( .A(B[1019]), .B(A[1019]), .Z(n2006) );
  XOR U3010 ( .A(A[1018]), .B(n2007), .Z(O[1018]) );
  AND U3011 ( .A(S), .B(n2008), .Z(n2007) );
  XOR U3012 ( .A(B[1018]), .B(A[1018]), .Z(n2008) );
  XOR U3013 ( .A(A[1017]), .B(n2009), .Z(O[1017]) );
  AND U3014 ( .A(S), .B(n2010), .Z(n2009) );
  XOR U3015 ( .A(B[1017]), .B(A[1017]), .Z(n2010) );
  XOR U3016 ( .A(A[1016]), .B(n2011), .Z(O[1016]) );
  AND U3017 ( .A(S), .B(n2012), .Z(n2011) );
  XOR U3018 ( .A(B[1016]), .B(A[1016]), .Z(n2012) );
  XOR U3019 ( .A(A[1015]), .B(n2013), .Z(O[1015]) );
  AND U3020 ( .A(S), .B(n2014), .Z(n2013) );
  XOR U3021 ( .A(B[1015]), .B(A[1015]), .Z(n2014) );
  XOR U3022 ( .A(A[1014]), .B(n2015), .Z(O[1014]) );
  AND U3023 ( .A(S), .B(n2016), .Z(n2015) );
  XOR U3024 ( .A(B[1014]), .B(A[1014]), .Z(n2016) );
  XOR U3025 ( .A(A[1013]), .B(n2017), .Z(O[1013]) );
  AND U3026 ( .A(S), .B(n2018), .Z(n2017) );
  XOR U3027 ( .A(B[1013]), .B(A[1013]), .Z(n2018) );
  XOR U3028 ( .A(A[1012]), .B(n2019), .Z(O[1012]) );
  AND U3029 ( .A(S), .B(n2020), .Z(n2019) );
  XOR U3030 ( .A(B[1012]), .B(A[1012]), .Z(n2020) );
  XOR U3031 ( .A(A[1011]), .B(n2021), .Z(O[1011]) );
  AND U3032 ( .A(S), .B(n2022), .Z(n2021) );
  XOR U3033 ( .A(B[1011]), .B(A[1011]), .Z(n2022) );
  XOR U3034 ( .A(A[1010]), .B(n2023), .Z(O[1010]) );
  AND U3035 ( .A(S), .B(n2024), .Z(n2023) );
  XOR U3036 ( .A(B[1010]), .B(A[1010]), .Z(n2024) );
  XOR U3037 ( .A(A[100]), .B(n2025), .Z(O[100]) );
  AND U3038 ( .A(S), .B(n2026), .Z(n2025) );
  XOR U3039 ( .A(B[100]), .B(A[100]), .Z(n2026) );
  XOR U3040 ( .A(A[1009]), .B(n2027), .Z(O[1009]) );
  AND U3041 ( .A(S), .B(n2028), .Z(n2027) );
  XOR U3042 ( .A(B[1009]), .B(A[1009]), .Z(n2028) );
  XOR U3043 ( .A(A[1008]), .B(n2029), .Z(O[1008]) );
  AND U3044 ( .A(S), .B(n2030), .Z(n2029) );
  XOR U3045 ( .A(B[1008]), .B(A[1008]), .Z(n2030) );
  XOR U3046 ( .A(A[1007]), .B(n2031), .Z(O[1007]) );
  AND U3047 ( .A(S), .B(n2032), .Z(n2031) );
  XOR U3048 ( .A(B[1007]), .B(A[1007]), .Z(n2032) );
  XOR U3049 ( .A(A[1006]), .B(n2033), .Z(O[1006]) );
  AND U3050 ( .A(S), .B(n2034), .Z(n2033) );
  XOR U3051 ( .A(B[1006]), .B(A[1006]), .Z(n2034) );
  XOR U3052 ( .A(A[1005]), .B(n2035), .Z(O[1005]) );
  AND U3053 ( .A(S), .B(n2036), .Z(n2035) );
  XOR U3054 ( .A(B[1005]), .B(A[1005]), .Z(n2036) );
  XOR U3055 ( .A(A[1004]), .B(n2037), .Z(O[1004]) );
  AND U3056 ( .A(S), .B(n2038), .Z(n2037) );
  XOR U3057 ( .A(B[1004]), .B(A[1004]), .Z(n2038) );
  XOR U3058 ( .A(A[1003]), .B(n2039), .Z(O[1003]) );
  AND U3059 ( .A(S), .B(n2040), .Z(n2039) );
  XOR U3060 ( .A(B[1003]), .B(A[1003]), .Z(n2040) );
  XOR U3061 ( .A(A[1002]), .B(n2041), .Z(O[1002]) );
  AND U3062 ( .A(S), .B(n2042), .Z(n2041) );
  XOR U3063 ( .A(B[1002]), .B(A[1002]), .Z(n2042) );
  XOR U3064 ( .A(A[1001]), .B(n2043), .Z(O[1001]) );
  AND U3065 ( .A(S), .B(n2044), .Z(n2043) );
  XOR U3066 ( .A(B[1001]), .B(A[1001]), .Z(n2044) );
  XOR U3067 ( .A(A[1000]), .B(n2045), .Z(O[1000]) );
  AND U3068 ( .A(S), .B(n2046), .Z(n2045) );
  XOR U3069 ( .A(B[1000]), .B(A[1000]), .Z(n2046) );
  XOR U3070 ( .A(A[0]), .B(n2047), .Z(O[0]) );
  AND U3071 ( .A(S), .B(n2048), .Z(n2047) );
  XOR U3072 ( .A(B[0]), .B(A[0]), .Z(n2048) );
endmodule


module MUX_N1024_2 ( A, B, S, O );
  input [1023:0] A;
  input [1023:0] B;
  output [1023:0] O;
  input S;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046;

  XOR U1 ( .A(B[8]), .B(n1), .Z(O[9]) );
  AND U2 ( .A(S), .B(n2), .Z(n1) );
  XOR U3 ( .A(B[9]), .B(B[8]), .Z(n2) );
  XOR U4 ( .A(B[98]), .B(n3), .Z(O[99]) );
  AND U5 ( .A(S), .B(n4), .Z(n3) );
  XOR U6 ( .A(B[99]), .B(B[98]), .Z(n4) );
  XOR U7 ( .A(B[998]), .B(n5), .Z(O[999]) );
  AND U8 ( .A(S), .B(n6), .Z(n5) );
  XOR U9 ( .A(B[999]), .B(B[998]), .Z(n6) );
  XOR U10 ( .A(B[997]), .B(n7), .Z(O[998]) );
  AND U11 ( .A(S), .B(n8), .Z(n7) );
  XOR U12 ( .A(B[998]), .B(B[997]), .Z(n8) );
  XOR U13 ( .A(B[996]), .B(n9), .Z(O[997]) );
  AND U14 ( .A(S), .B(n10), .Z(n9) );
  XOR U15 ( .A(B[997]), .B(B[996]), .Z(n10) );
  XOR U16 ( .A(B[995]), .B(n11), .Z(O[996]) );
  AND U17 ( .A(S), .B(n12), .Z(n11) );
  XOR U18 ( .A(B[996]), .B(B[995]), .Z(n12) );
  XOR U19 ( .A(B[994]), .B(n13), .Z(O[995]) );
  AND U20 ( .A(S), .B(n14), .Z(n13) );
  XOR U21 ( .A(B[995]), .B(B[994]), .Z(n14) );
  XOR U22 ( .A(B[993]), .B(n15), .Z(O[994]) );
  AND U23 ( .A(S), .B(n16), .Z(n15) );
  XOR U24 ( .A(B[994]), .B(B[993]), .Z(n16) );
  XOR U25 ( .A(B[992]), .B(n17), .Z(O[993]) );
  AND U26 ( .A(S), .B(n18), .Z(n17) );
  XOR U27 ( .A(B[993]), .B(B[992]), .Z(n18) );
  XOR U28 ( .A(B[991]), .B(n19), .Z(O[992]) );
  AND U29 ( .A(S), .B(n20), .Z(n19) );
  XOR U30 ( .A(B[992]), .B(B[991]), .Z(n20) );
  XOR U31 ( .A(B[990]), .B(n21), .Z(O[991]) );
  AND U32 ( .A(S), .B(n22), .Z(n21) );
  XOR U33 ( .A(B[991]), .B(B[990]), .Z(n22) );
  XOR U34 ( .A(B[989]), .B(n23), .Z(O[990]) );
  AND U35 ( .A(S), .B(n24), .Z(n23) );
  XOR U36 ( .A(B[990]), .B(B[989]), .Z(n24) );
  XOR U37 ( .A(B[97]), .B(n25), .Z(O[98]) );
  AND U38 ( .A(S), .B(n26), .Z(n25) );
  XOR U39 ( .A(B[98]), .B(B[97]), .Z(n26) );
  XOR U40 ( .A(B[988]), .B(n27), .Z(O[989]) );
  AND U41 ( .A(S), .B(n28), .Z(n27) );
  XOR U42 ( .A(B[989]), .B(B[988]), .Z(n28) );
  XOR U43 ( .A(B[987]), .B(n29), .Z(O[988]) );
  AND U44 ( .A(S), .B(n30), .Z(n29) );
  XOR U45 ( .A(B[988]), .B(B[987]), .Z(n30) );
  XOR U46 ( .A(B[986]), .B(n31), .Z(O[987]) );
  AND U47 ( .A(S), .B(n32), .Z(n31) );
  XOR U48 ( .A(B[987]), .B(B[986]), .Z(n32) );
  XOR U49 ( .A(B[985]), .B(n33), .Z(O[986]) );
  AND U50 ( .A(S), .B(n34), .Z(n33) );
  XOR U51 ( .A(B[986]), .B(B[985]), .Z(n34) );
  XOR U52 ( .A(B[984]), .B(n35), .Z(O[985]) );
  AND U53 ( .A(S), .B(n36), .Z(n35) );
  XOR U54 ( .A(B[985]), .B(B[984]), .Z(n36) );
  XOR U55 ( .A(B[983]), .B(n37), .Z(O[984]) );
  AND U56 ( .A(S), .B(n38), .Z(n37) );
  XOR U57 ( .A(B[984]), .B(B[983]), .Z(n38) );
  XOR U58 ( .A(B[982]), .B(n39), .Z(O[983]) );
  AND U59 ( .A(S), .B(n40), .Z(n39) );
  XOR U60 ( .A(B[983]), .B(B[982]), .Z(n40) );
  XOR U61 ( .A(B[981]), .B(n41), .Z(O[982]) );
  AND U62 ( .A(S), .B(n42), .Z(n41) );
  XOR U63 ( .A(B[982]), .B(B[981]), .Z(n42) );
  XOR U64 ( .A(B[980]), .B(n43), .Z(O[981]) );
  AND U65 ( .A(S), .B(n44), .Z(n43) );
  XOR U66 ( .A(B[981]), .B(B[980]), .Z(n44) );
  XOR U67 ( .A(B[979]), .B(n45), .Z(O[980]) );
  AND U68 ( .A(S), .B(n46), .Z(n45) );
  XOR U69 ( .A(B[980]), .B(B[979]), .Z(n46) );
  XOR U70 ( .A(B[96]), .B(n47), .Z(O[97]) );
  AND U71 ( .A(S), .B(n48), .Z(n47) );
  XOR U72 ( .A(B[97]), .B(B[96]), .Z(n48) );
  XOR U73 ( .A(B[978]), .B(n49), .Z(O[979]) );
  AND U74 ( .A(S), .B(n50), .Z(n49) );
  XOR U75 ( .A(B[979]), .B(B[978]), .Z(n50) );
  XOR U76 ( .A(B[977]), .B(n51), .Z(O[978]) );
  AND U77 ( .A(S), .B(n52), .Z(n51) );
  XOR U78 ( .A(B[978]), .B(B[977]), .Z(n52) );
  XOR U79 ( .A(B[976]), .B(n53), .Z(O[977]) );
  AND U80 ( .A(S), .B(n54), .Z(n53) );
  XOR U81 ( .A(B[977]), .B(B[976]), .Z(n54) );
  XOR U82 ( .A(B[975]), .B(n55), .Z(O[976]) );
  AND U83 ( .A(S), .B(n56), .Z(n55) );
  XOR U84 ( .A(B[976]), .B(B[975]), .Z(n56) );
  XOR U85 ( .A(B[974]), .B(n57), .Z(O[975]) );
  AND U86 ( .A(S), .B(n58), .Z(n57) );
  XOR U87 ( .A(B[975]), .B(B[974]), .Z(n58) );
  XOR U88 ( .A(B[973]), .B(n59), .Z(O[974]) );
  AND U89 ( .A(S), .B(n60), .Z(n59) );
  XOR U90 ( .A(B[974]), .B(B[973]), .Z(n60) );
  XOR U91 ( .A(B[972]), .B(n61), .Z(O[973]) );
  AND U92 ( .A(S), .B(n62), .Z(n61) );
  XOR U93 ( .A(B[973]), .B(B[972]), .Z(n62) );
  XOR U94 ( .A(B[971]), .B(n63), .Z(O[972]) );
  AND U95 ( .A(S), .B(n64), .Z(n63) );
  XOR U96 ( .A(B[972]), .B(B[971]), .Z(n64) );
  XOR U97 ( .A(B[970]), .B(n65), .Z(O[971]) );
  AND U98 ( .A(S), .B(n66), .Z(n65) );
  XOR U99 ( .A(B[971]), .B(B[970]), .Z(n66) );
  XOR U100 ( .A(B[969]), .B(n67), .Z(O[970]) );
  AND U101 ( .A(S), .B(n68), .Z(n67) );
  XOR U102 ( .A(B[970]), .B(B[969]), .Z(n68) );
  XOR U103 ( .A(B[95]), .B(n69), .Z(O[96]) );
  AND U104 ( .A(S), .B(n70), .Z(n69) );
  XOR U105 ( .A(B[96]), .B(B[95]), .Z(n70) );
  XOR U106 ( .A(B[968]), .B(n71), .Z(O[969]) );
  AND U107 ( .A(S), .B(n72), .Z(n71) );
  XOR U108 ( .A(B[969]), .B(B[968]), .Z(n72) );
  XOR U109 ( .A(B[967]), .B(n73), .Z(O[968]) );
  AND U110 ( .A(S), .B(n74), .Z(n73) );
  XOR U111 ( .A(B[968]), .B(B[967]), .Z(n74) );
  XOR U112 ( .A(B[966]), .B(n75), .Z(O[967]) );
  AND U113 ( .A(S), .B(n76), .Z(n75) );
  XOR U114 ( .A(B[967]), .B(B[966]), .Z(n76) );
  XOR U115 ( .A(B[965]), .B(n77), .Z(O[966]) );
  AND U116 ( .A(S), .B(n78), .Z(n77) );
  XOR U117 ( .A(B[966]), .B(B[965]), .Z(n78) );
  XOR U118 ( .A(B[964]), .B(n79), .Z(O[965]) );
  AND U119 ( .A(S), .B(n80), .Z(n79) );
  XOR U120 ( .A(B[965]), .B(B[964]), .Z(n80) );
  XOR U121 ( .A(B[963]), .B(n81), .Z(O[964]) );
  AND U122 ( .A(S), .B(n82), .Z(n81) );
  XOR U123 ( .A(B[964]), .B(B[963]), .Z(n82) );
  XOR U124 ( .A(B[962]), .B(n83), .Z(O[963]) );
  AND U125 ( .A(S), .B(n84), .Z(n83) );
  XOR U126 ( .A(B[963]), .B(B[962]), .Z(n84) );
  XOR U127 ( .A(B[961]), .B(n85), .Z(O[962]) );
  AND U128 ( .A(S), .B(n86), .Z(n85) );
  XOR U129 ( .A(B[962]), .B(B[961]), .Z(n86) );
  XOR U130 ( .A(B[960]), .B(n87), .Z(O[961]) );
  AND U131 ( .A(S), .B(n88), .Z(n87) );
  XOR U132 ( .A(B[961]), .B(B[960]), .Z(n88) );
  XOR U133 ( .A(B[959]), .B(n89), .Z(O[960]) );
  AND U134 ( .A(S), .B(n90), .Z(n89) );
  XOR U135 ( .A(B[960]), .B(B[959]), .Z(n90) );
  XOR U136 ( .A(B[94]), .B(n91), .Z(O[95]) );
  AND U137 ( .A(S), .B(n92), .Z(n91) );
  XOR U138 ( .A(B[95]), .B(B[94]), .Z(n92) );
  XOR U139 ( .A(B[958]), .B(n93), .Z(O[959]) );
  AND U140 ( .A(S), .B(n94), .Z(n93) );
  XOR U141 ( .A(B[959]), .B(B[958]), .Z(n94) );
  XOR U142 ( .A(B[957]), .B(n95), .Z(O[958]) );
  AND U143 ( .A(S), .B(n96), .Z(n95) );
  XOR U144 ( .A(B[958]), .B(B[957]), .Z(n96) );
  XOR U145 ( .A(B[956]), .B(n97), .Z(O[957]) );
  AND U146 ( .A(S), .B(n98), .Z(n97) );
  XOR U147 ( .A(B[957]), .B(B[956]), .Z(n98) );
  XOR U148 ( .A(B[955]), .B(n99), .Z(O[956]) );
  AND U149 ( .A(S), .B(n100), .Z(n99) );
  XOR U150 ( .A(B[956]), .B(B[955]), .Z(n100) );
  XOR U151 ( .A(B[954]), .B(n101), .Z(O[955]) );
  AND U152 ( .A(S), .B(n102), .Z(n101) );
  XOR U153 ( .A(B[955]), .B(B[954]), .Z(n102) );
  XOR U154 ( .A(B[953]), .B(n103), .Z(O[954]) );
  AND U155 ( .A(S), .B(n104), .Z(n103) );
  XOR U156 ( .A(B[954]), .B(B[953]), .Z(n104) );
  XOR U157 ( .A(B[952]), .B(n105), .Z(O[953]) );
  AND U158 ( .A(S), .B(n106), .Z(n105) );
  XOR U159 ( .A(B[953]), .B(B[952]), .Z(n106) );
  XOR U160 ( .A(B[951]), .B(n107), .Z(O[952]) );
  AND U161 ( .A(S), .B(n108), .Z(n107) );
  XOR U162 ( .A(B[952]), .B(B[951]), .Z(n108) );
  XOR U163 ( .A(B[950]), .B(n109), .Z(O[951]) );
  AND U164 ( .A(S), .B(n110), .Z(n109) );
  XOR U165 ( .A(B[951]), .B(B[950]), .Z(n110) );
  XOR U166 ( .A(B[949]), .B(n111), .Z(O[950]) );
  AND U167 ( .A(S), .B(n112), .Z(n111) );
  XOR U168 ( .A(B[950]), .B(B[949]), .Z(n112) );
  XOR U169 ( .A(B[93]), .B(n113), .Z(O[94]) );
  AND U170 ( .A(S), .B(n114), .Z(n113) );
  XOR U171 ( .A(B[94]), .B(B[93]), .Z(n114) );
  XOR U172 ( .A(B[948]), .B(n115), .Z(O[949]) );
  AND U173 ( .A(S), .B(n116), .Z(n115) );
  XOR U174 ( .A(B[949]), .B(B[948]), .Z(n116) );
  XOR U175 ( .A(B[947]), .B(n117), .Z(O[948]) );
  AND U176 ( .A(S), .B(n118), .Z(n117) );
  XOR U177 ( .A(B[948]), .B(B[947]), .Z(n118) );
  XOR U178 ( .A(B[946]), .B(n119), .Z(O[947]) );
  AND U179 ( .A(S), .B(n120), .Z(n119) );
  XOR U180 ( .A(B[947]), .B(B[946]), .Z(n120) );
  XOR U181 ( .A(B[945]), .B(n121), .Z(O[946]) );
  AND U182 ( .A(S), .B(n122), .Z(n121) );
  XOR U183 ( .A(B[946]), .B(B[945]), .Z(n122) );
  XOR U184 ( .A(B[944]), .B(n123), .Z(O[945]) );
  AND U185 ( .A(S), .B(n124), .Z(n123) );
  XOR U186 ( .A(B[945]), .B(B[944]), .Z(n124) );
  XOR U187 ( .A(B[943]), .B(n125), .Z(O[944]) );
  AND U188 ( .A(S), .B(n126), .Z(n125) );
  XOR U189 ( .A(B[944]), .B(B[943]), .Z(n126) );
  XOR U190 ( .A(B[942]), .B(n127), .Z(O[943]) );
  AND U191 ( .A(S), .B(n128), .Z(n127) );
  XOR U192 ( .A(B[943]), .B(B[942]), .Z(n128) );
  XOR U193 ( .A(B[941]), .B(n129), .Z(O[942]) );
  AND U194 ( .A(S), .B(n130), .Z(n129) );
  XOR U195 ( .A(B[942]), .B(B[941]), .Z(n130) );
  XOR U196 ( .A(B[940]), .B(n131), .Z(O[941]) );
  AND U197 ( .A(S), .B(n132), .Z(n131) );
  XOR U198 ( .A(B[941]), .B(B[940]), .Z(n132) );
  XOR U199 ( .A(B[939]), .B(n133), .Z(O[940]) );
  AND U200 ( .A(S), .B(n134), .Z(n133) );
  XOR U201 ( .A(B[940]), .B(B[939]), .Z(n134) );
  XOR U202 ( .A(B[92]), .B(n135), .Z(O[93]) );
  AND U203 ( .A(S), .B(n136), .Z(n135) );
  XOR U204 ( .A(B[93]), .B(B[92]), .Z(n136) );
  XOR U205 ( .A(B[938]), .B(n137), .Z(O[939]) );
  AND U206 ( .A(S), .B(n138), .Z(n137) );
  XOR U207 ( .A(B[939]), .B(B[938]), .Z(n138) );
  XOR U208 ( .A(B[937]), .B(n139), .Z(O[938]) );
  AND U209 ( .A(S), .B(n140), .Z(n139) );
  XOR U210 ( .A(B[938]), .B(B[937]), .Z(n140) );
  XOR U211 ( .A(B[936]), .B(n141), .Z(O[937]) );
  AND U212 ( .A(S), .B(n142), .Z(n141) );
  XOR U213 ( .A(B[937]), .B(B[936]), .Z(n142) );
  XOR U214 ( .A(B[935]), .B(n143), .Z(O[936]) );
  AND U215 ( .A(S), .B(n144), .Z(n143) );
  XOR U216 ( .A(B[936]), .B(B[935]), .Z(n144) );
  XOR U217 ( .A(B[934]), .B(n145), .Z(O[935]) );
  AND U218 ( .A(S), .B(n146), .Z(n145) );
  XOR U219 ( .A(B[935]), .B(B[934]), .Z(n146) );
  XOR U220 ( .A(B[933]), .B(n147), .Z(O[934]) );
  AND U221 ( .A(S), .B(n148), .Z(n147) );
  XOR U222 ( .A(B[934]), .B(B[933]), .Z(n148) );
  XOR U223 ( .A(B[932]), .B(n149), .Z(O[933]) );
  AND U224 ( .A(S), .B(n150), .Z(n149) );
  XOR U225 ( .A(B[933]), .B(B[932]), .Z(n150) );
  XOR U226 ( .A(B[931]), .B(n151), .Z(O[932]) );
  AND U227 ( .A(S), .B(n152), .Z(n151) );
  XOR U228 ( .A(B[932]), .B(B[931]), .Z(n152) );
  XOR U229 ( .A(B[930]), .B(n153), .Z(O[931]) );
  AND U230 ( .A(S), .B(n154), .Z(n153) );
  XOR U231 ( .A(B[931]), .B(B[930]), .Z(n154) );
  XOR U232 ( .A(B[929]), .B(n155), .Z(O[930]) );
  AND U233 ( .A(S), .B(n156), .Z(n155) );
  XOR U234 ( .A(B[930]), .B(B[929]), .Z(n156) );
  XOR U235 ( .A(B[91]), .B(n157), .Z(O[92]) );
  AND U236 ( .A(S), .B(n158), .Z(n157) );
  XOR U237 ( .A(B[92]), .B(B[91]), .Z(n158) );
  XOR U238 ( .A(B[928]), .B(n159), .Z(O[929]) );
  AND U239 ( .A(S), .B(n160), .Z(n159) );
  XOR U240 ( .A(B[929]), .B(B[928]), .Z(n160) );
  XOR U241 ( .A(B[927]), .B(n161), .Z(O[928]) );
  AND U242 ( .A(S), .B(n162), .Z(n161) );
  XOR U243 ( .A(B[928]), .B(B[927]), .Z(n162) );
  XOR U244 ( .A(B[926]), .B(n163), .Z(O[927]) );
  AND U245 ( .A(S), .B(n164), .Z(n163) );
  XOR U246 ( .A(B[927]), .B(B[926]), .Z(n164) );
  XOR U247 ( .A(B[925]), .B(n165), .Z(O[926]) );
  AND U248 ( .A(S), .B(n166), .Z(n165) );
  XOR U249 ( .A(B[926]), .B(B[925]), .Z(n166) );
  XOR U250 ( .A(B[924]), .B(n167), .Z(O[925]) );
  AND U251 ( .A(S), .B(n168), .Z(n167) );
  XOR U252 ( .A(B[925]), .B(B[924]), .Z(n168) );
  XOR U253 ( .A(B[923]), .B(n169), .Z(O[924]) );
  AND U254 ( .A(S), .B(n170), .Z(n169) );
  XOR U255 ( .A(B[924]), .B(B[923]), .Z(n170) );
  XOR U256 ( .A(B[922]), .B(n171), .Z(O[923]) );
  AND U257 ( .A(S), .B(n172), .Z(n171) );
  XOR U258 ( .A(B[923]), .B(B[922]), .Z(n172) );
  XOR U259 ( .A(B[921]), .B(n173), .Z(O[922]) );
  AND U260 ( .A(S), .B(n174), .Z(n173) );
  XOR U261 ( .A(B[922]), .B(B[921]), .Z(n174) );
  XOR U262 ( .A(B[920]), .B(n175), .Z(O[921]) );
  AND U263 ( .A(S), .B(n176), .Z(n175) );
  XOR U264 ( .A(B[921]), .B(B[920]), .Z(n176) );
  XOR U265 ( .A(B[919]), .B(n177), .Z(O[920]) );
  AND U266 ( .A(S), .B(n178), .Z(n177) );
  XOR U267 ( .A(B[920]), .B(B[919]), .Z(n178) );
  XOR U268 ( .A(B[90]), .B(n179), .Z(O[91]) );
  AND U269 ( .A(S), .B(n180), .Z(n179) );
  XOR U270 ( .A(B[91]), .B(B[90]), .Z(n180) );
  XOR U271 ( .A(B[918]), .B(n181), .Z(O[919]) );
  AND U272 ( .A(S), .B(n182), .Z(n181) );
  XOR U273 ( .A(B[919]), .B(B[918]), .Z(n182) );
  XOR U274 ( .A(B[917]), .B(n183), .Z(O[918]) );
  AND U275 ( .A(S), .B(n184), .Z(n183) );
  XOR U276 ( .A(B[918]), .B(B[917]), .Z(n184) );
  XOR U277 ( .A(B[916]), .B(n185), .Z(O[917]) );
  AND U278 ( .A(S), .B(n186), .Z(n185) );
  XOR U279 ( .A(B[917]), .B(B[916]), .Z(n186) );
  XOR U280 ( .A(B[915]), .B(n187), .Z(O[916]) );
  AND U281 ( .A(S), .B(n188), .Z(n187) );
  XOR U282 ( .A(B[916]), .B(B[915]), .Z(n188) );
  XOR U283 ( .A(B[914]), .B(n189), .Z(O[915]) );
  AND U284 ( .A(S), .B(n190), .Z(n189) );
  XOR U285 ( .A(B[915]), .B(B[914]), .Z(n190) );
  XOR U286 ( .A(B[913]), .B(n191), .Z(O[914]) );
  AND U287 ( .A(S), .B(n192), .Z(n191) );
  XOR U288 ( .A(B[914]), .B(B[913]), .Z(n192) );
  XOR U289 ( .A(B[912]), .B(n193), .Z(O[913]) );
  AND U290 ( .A(S), .B(n194), .Z(n193) );
  XOR U291 ( .A(B[913]), .B(B[912]), .Z(n194) );
  XOR U292 ( .A(B[911]), .B(n195), .Z(O[912]) );
  AND U293 ( .A(S), .B(n196), .Z(n195) );
  XOR U294 ( .A(B[912]), .B(B[911]), .Z(n196) );
  XOR U295 ( .A(B[910]), .B(n197), .Z(O[911]) );
  AND U296 ( .A(S), .B(n198), .Z(n197) );
  XOR U297 ( .A(B[911]), .B(B[910]), .Z(n198) );
  XOR U298 ( .A(B[909]), .B(n199), .Z(O[910]) );
  AND U299 ( .A(S), .B(n200), .Z(n199) );
  XOR U300 ( .A(B[910]), .B(B[909]), .Z(n200) );
  XOR U301 ( .A(B[89]), .B(n201), .Z(O[90]) );
  AND U302 ( .A(S), .B(n202), .Z(n201) );
  XOR U303 ( .A(B[90]), .B(B[89]), .Z(n202) );
  XOR U304 ( .A(B[908]), .B(n203), .Z(O[909]) );
  AND U305 ( .A(S), .B(n204), .Z(n203) );
  XOR U306 ( .A(B[909]), .B(B[908]), .Z(n204) );
  XOR U307 ( .A(B[907]), .B(n205), .Z(O[908]) );
  AND U308 ( .A(S), .B(n206), .Z(n205) );
  XOR U309 ( .A(B[908]), .B(B[907]), .Z(n206) );
  XOR U310 ( .A(B[906]), .B(n207), .Z(O[907]) );
  AND U311 ( .A(S), .B(n208), .Z(n207) );
  XOR U312 ( .A(B[907]), .B(B[906]), .Z(n208) );
  XOR U313 ( .A(B[905]), .B(n209), .Z(O[906]) );
  AND U314 ( .A(S), .B(n210), .Z(n209) );
  XOR U315 ( .A(B[906]), .B(B[905]), .Z(n210) );
  XOR U316 ( .A(B[904]), .B(n211), .Z(O[905]) );
  AND U317 ( .A(S), .B(n212), .Z(n211) );
  XOR U318 ( .A(B[905]), .B(B[904]), .Z(n212) );
  XOR U319 ( .A(B[903]), .B(n213), .Z(O[904]) );
  AND U320 ( .A(S), .B(n214), .Z(n213) );
  XOR U321 ( .A(B[904]), .B(B[903]), .Z(n214) );
  XOR U322 ( .A(B[902]), .B(n215), .Z(O[903]) );
  AND U323 ( .A(S), .B(n216), .Z(n215) );
  XOR U324 ( .A(B[903]), .B(B[902]), .Z(n216) );
  XOR U325 ( .A(B[901]), .B(n217), .Z(O[902]) );
  AND U326 ( .A(S), .B(n218), .Z(n217) );
  XOR U327 ( .A(B[902]), .B(B[901]), .Z(n218) );
  XOR U328 ( .A(B[900]), .B(n219), .Z(O[901]) );
  AND U329 ( .A(S), .B(n220), .Z(n219) );
  XOR U330 ( .A(B[901]), .B(B[900]), .Z(n220) );
  XOR U331 ( .A(B[899]), .B(n221), .Z(O[900]) );
  AND U332 ( .A(S), .B(n222), .Z(n221) );
  XOR U333 ( .A(B[900]), .B(B[899]), .Z(n222) );
  XOR U334 ( .A(B[7]), .B(n223), .Z(O[8]) );
  AND U335 ( .A(S), .B(n224), .Z(n223) );
  XOR U336 ( .A(B[8]), .B(B[7]), .Z(n224) );
  XOR U337 ( .A(B[88]), .B(n225), .Z(O[89]) );
  AND U338 ( .A(S), .B(n226), .Z(n225) );
  XOR U339 ( .A(B[89]), .B(B[88]), .Z(n226) );
  XOR U340 ( .A(B[898]), .B(n227), .Z(O[899]) );
  AND U341 ( .A(S), .B(n228), .Z(n227) );
  XOR U342 ( .A(B[899]), .B(B[898]), .Z(n228) );
  XOR U343 ( .A(B[897]), .B(n229), .Z(O[898]) );
  AND U344 ( .A(S), .B(n230), .Z(n229) );
  XOR U345 ( .A(B[898]), .B(B[897]), .Z(n230) );
  XOR U346 ( .A(B[896]), .B(n231), .Z(O[897]) );
  AND U347 ( .A(S), .B(n232), .Z(n231) );
  XOR U348 ( .A(B[897]), .B(B[896]), .Z(n232) );
  XOR U349 ( .A(B[895]), .B(n233), .Z(O[896]) );
  AND U350 ( .A(S), .B(n234), .Z(n233) );
  XOR U351 ( .A(B[896]), .B(B[895]), .Z(n234) );
  XOR U352 ( .A(B[894]), .B(n235), .Z(O[895]) );
  AND U353 ( .A(S), .B(n236), .Z(n235) );
  XOR U354 ( .A(B[895]), .B(B[894]), .Z(n236) );
  XOR U355 ( .A(B[893]), .B(n237), .Z(O[894]) );
  AND U356 ( .A(S), .B(n238), .Z(n237) );
  XOR U357 ( .A(B[894]), .B(B[893]), .Z(n238) );
  XOR U358 ( .A(B[892]), .B(n239), .Z(O[893]) );
  AND U359 ( .A(S), .B(n240), .Z(n239) );
  XOR U360 ( .A(B[893]), .B(B[892]), .Z(n240) );
  XOR U361 ( .A(B[891]), .B(n241), .Z(O[892]) );
  AND U362 ( .A(S), .B(n242), .Z(n241) );
  XOR U363 ( .A(B[892]), .B(B[891]), .Z(n242) );
  XOR U364 ( .A(B[890]), .B(n243), .Z(O[891]) );
  AND U365 ( .A(S), .B(n244), .Z(n243) );
  XOR U366 ( .A(B[891]), .B(B[890]), .Z(n244) );
  XOR U367 ( .A(B[889]), .B(n245), .Z(O[890]) );
  AND U368 ( .A(S), .B(n246), .Z(n245) );
  XOR U369 ( .A(B[890]), .B(B[889]), .Z(n246) );
  XOR U370 ( .A(B[87]), .B(n247), .Z(O[88]) );
  AND U371 ( .A(S), .B(n248), .Z(n247) );
  XOR U372 ( .A(B[88]), .B(B[87]), .Z(n248) );
  XOR U373 ( .A(B[888]), .B(n249), .Z(O[889]) );
  AND U374 ( .A(S), .B(n250), .Z(n249) );
  XOR U375 ( .A(B[889]), .B(B[888]), .Z(n250) );
  XOR U376 ( .A(B[887]), .B(n251), .Z(O[888]) );
  AND U377 ( .A(S), .B(n252), .Z(n251) );
  XOR U378 ( .A(B[888]), .B(B[887]), .Z(n252) );
  XOR U379 ( .A(B[886]), .B(n253), .Z(O[887]) );
  AND U380 ( .A(S), .B(n254), .Z(n253) );
  XOR U381 ( .A(B[887]), .B(B[886]), .Z(n254) );
  XOR U382 ( .A(B[885]), .B(n255), .Z(O[886]) );
  AND U383 ( .A(S), .B(n256), .Z(n255) );
  XOR U384 ( .A(B[886]), .B(B[885]), .Z(n256) );
  XOR U385 ( .A(B[884]), .B(n257), .Z(O[885]) );
  AND U386 ( .A(S), .B(n258), .Z(n257) );
  XOR U387 ( .A(B[885]), .B(B[884]), .Z(n258) );
  XOR U388 ( .A(B[883]), .B(n259), .Z(O[884]) );
  AND U389 ( .A(S), .B(n260), .Z(n259) );
  XOR U390 ( .A(B[884]), .B(B[883]), .Z(n260) );
  XOR U391 ( .A(B[882]), .B(n261), .Z(O[883]) );
  AND U392 ( .A(S), .B(n262), .Z(n261) );
  XOR U393 ( .A(B[883]), .B(B[882]), .Z(n262) );
  XOR U394 ( .A(B[881]), .B(n263), .Z(O[882]) );
  AND U395 ( .A(S), .B(n264), .Z(n263) );
  XOR U396 ( .A(B[882]), .B(B[881]), .Z(n264) );
  XOR U397 ( .A(B[880]), .B(n265), .Z(O[881]) );
  AND U398 ( .A(S), .B(n266), .Z(n265) );
  XOR U399 ( .A(B[881]), .B(B[880]), .Z(n266) );
  XOR U400 ( .A(B[879]), .B(n267), .Z(O[880]) );
  AND U401 ( .A(S), .B(n268), .Z(n267) );
  XOR U402 ( .A(B[880]), .B(B[879]), .Z(n268) );
  XOR U403 ( .A(B[86]), .B(n269), .Z(O[87]) );
  AND U404 ( .A(S), .B(n270), .Z(n269) );
  XOR U405 ( .A(B[87]), .B(B[86]), .Z(n270) );
  XOR U406 ( .A(B[878]), .B(n271), .Z(O[879]) );
  AND U407 ( .A(S), .B(n272), .Z(n271) );
  XOR U408 ( .A(B[879]), .B(B[878]), .Z(n272) );
  XOR U409 ( .A(B[877]), .B(n273), .Z(O[878]) );
  AND U410 ( .A(S), .B(n274), .Z(n273) );
  XOR U411 ( .A(B[878]), .B(B[877]), .Z(n274) );
  XOR U412 ( .A(B[876]), .B(n275), .Z(O[877]) );
  AND U413 ( .A(S), .B(n276), .Z(n275) );
  XOR U414 ( .A(B[877]), .B(B[876]), .Z(n276) );
  XOR U415 ( .A(B[875]), .B(n277), .Z(O[876]) );
  AND U416 ( .A(S), .B(n278), .Z(n277) );
  XOR U417 ( .A(B[876]), .B(B[875]), .Z(n278) );
  XOR U418 ( .A(B[874]), .B(n279), .Z(O[875]) );
  AND U419 ( .A(S), .B(n280), .Z(n279) );
  XOR U420 ( .A(B[875]), .B(B[874]), .Z(n280) );
  XOR U421 ( .A(B[873]), .B(n281), .Z(O[874]) );
  AND U422 ( .A(S), .B(n282), .Z(n281) );
  XOR U423 ( .A(B[874]), .B(B[873]), .Z(n282) );
  XOR U424 ( .A(B[872]), .B(n283), .Z(O[873]) );
  AND U425 ( .A(S), .B(n284), .Z(n283) );
  XOR U426 ( .A(B[873]), .B(B[872]), .Z(n284) );
  XOR U427 ( .A(B[871]), .B(n285), .Z(O[872]) );
  AND U428 ( .A(S), .B(n286), .Z(n285) );
  XOR U429 ( .A(B[872]), .B(B[871]), .Z(n286) );
  XOR U430 ( .A(B[870]), .B(n287), .Z(O[871]) );
  AND U431 ( .A(S), .B(n288), .Z(n287) );
  XOR U432 ( .A(B[871]), .B(B[870]), .Z(n288) );
  XOR U433 ( .A(B[869]), .B(n289), .Z(O[870]) );
  AND U434 ( .A(S), .B(n290), .Z(n289) );
  XOR U435 ( .A(B[870]), .B(B[869]), .Z(n290) );
  XOR U436 ( .A(B[85]), .B(n291), .Z(O[86]) );
  AND U437 ( .A(S), .B(n292), .Z(n291) );
  XOR U438 ( .A(B[86]), .B(B[85]), .Z(n292) );
  XOR U439 ( .A(B[868]), .B(n293), .Z(O[869]) );
  AND U440 ( .A(S), .B(n294), .Z(n293) );
  XOR U441 ( .A(B[869]), .B(B[868]), .Z(n294) );
  XOR U442 ( .A(B[867]), .B(n295), .Z(O[868]) );
  AND U443 ( .A(S), .B(n296), .Z(n295) );
  XOR U444 ( .A(B[868]), .B(B[867]), .Z(n296) );
  XOR U445 ( .A(B[866]), .B(n297), .Z(O[867]) );
  AND U446 ( .A(S), .B(n298), .Z(n297) );
  XOR U447 ( .A(B[867]), .B(B[866]), .Z(n298) );
  XOR U448 ( .A(B[865]), .B(n299), .Z(O[866]) );
  AND U449 ( .A(S), .B(n300), .Z(n299) );
  XOR U450 ( .A(B[866]), .B(B[865]), .Z(n300) );
  XOR U451 ( .A(B[864]), .B(n301), .Z(O[865]) );
  AND U452 ( .A(S), .B(n302), .Z(n301) );
  XOR U453 ( .A(B[865]), .B(B[864]), .Z(n302) );
  XOR U454 ( .A(B[863]), .B(n303), .Z(O[864]) );
  AND U455 ( .A(S), .B(n304), .Z(n303) );
  XOR U456 ( .A(B[864]), .B(B[863]), .Z(n304) );
  XOR U457 ( .A(B[862]), .B(n305), .Z(O[863]) );
  AND U458 ( .A(S), .B(n306), .Z(n305) );
  XOR U459 ( .A(B[863]), .B(B[862]), .Z(n306) );
  XOR U460 ( .A(B[861]), .B(n307), .Z(O[862]) );
  AND U461 ( .A(S), .B(n308), .Z(n307) );
  XOR U462 ( .A(B[862]), .B(B[861]), .Z(n308) );
  XOR U463 ( .A(B[860]), .B(n309), .Z(O[861]) );
  AND U464 ( .A(S), .B(n310), .Z(n309) );
  XOR U465 ( .A(B[861]), .B(B[860]), .Z(n310) );
  XOR U466 ( .A(B[859]), .B(n311), .Z(O[860]) );
  AND U467 ( .A(S), .B(n312), .Z(n311) );
  XOR U468 ( .A(B[860]), .B(B[859]), .Z(n312) );
  XOR U469 ( .A(B[84]), .B(n313), .Z(O[85]) );
  AND U470 ( .A(S), .B(n314), .Z(n313) );
  XOR U471 ( .A(B[85]), .B(B[84]), .Z(n314) );
  XOR U472 ( .A(B[858]), .B(n315), .Z(O[859]) );
  AND U473 ( .A(S), .B(n316), .Z(n315) );
  XOR U474 ( .A(B[859]), .B(B[858]), .Z(n316) );
  XOR U475 ( .A(B[857]), .B(n317), .Z(O[858]) );
  AND U476 ( .A(S), .B(n318), .Z(n317) );
  XOR U477 ( .A(B[858]), .B(B[857]), .Z(n318) );
  XOR U478 ( .A(B[856]), .B(n319), .Z(O[857]) );
  AND U479 ( .A(S), .B(n320), .Z(n319) );
  XOR U480 ( .A(B[857]), .B(B[856]), .Z(n320) );
  XOR U481 ( .A(B[855]), .B(n321), .Z(O[856]) );
  AND U482 ( .A(S), .B(n322), .Z(n321) );
  XOR U483 ( .A(B[856]), .B(B[855]), .Z(n322) );
  XOR U484 ( .A(B[854]), .B(n323), .Z(O[855]) );
  AND U485 ( .A(S), .B(n324), .Z(n323) );
  XOR U486 ( .A(B[855]), .B(B[854]), .Z(n324) );
  XOR U487 ( .A(B[853]), .B(n325), .Z(O[854]) );
  AND U488 ( .A(S), .B(n326), .Z(n325) );
  XOR U489 ( .A(B[854]), .B(B[853]), .Z(n326) );
  XOR U490 ( .A(B[852]), .B(n327), .Z(O[853]) );
  AND U491 ( .A(S), .B(n328), .Z(n327) );
  XOR U492 ( .A(B[853]), .B(B[852]), .Z(n328) );
  XOR U493 ( .A(B[851]), .B(n329), .Z(O[852]) );
  AND U494 ( .A(S), .B(n330), .Z(n329) );
  XOR U495 ( .A(B[852]), .B(B[851]), .Z(n330) );
  XOR U496 ( .A(B[850]), .B(n331), .Z(O[851]) );
  AND U497 ( .A(S), .B(n332), .Z(n331) );
  XOR U498 ( .A(B[851]), .B(B[850]), .Z(n332) );
  XOR U499 ( .A(B[849]), .B(n333), .Z(O[850]) );
  AND U500 ( .A(S), .B(n334), .Z(n333) );
  XOR U501 ( .A(B[850]), .B(B[849]), .Z(n334) );
  XOR U502 ( .A(B[83]), .B(n335), .Z(O[84]) );
  AND U503 ( .A(S), .B(n336), .Z(n335) );
  XOR U504 ( .A(B[84]), .B(B[83]), .Z(n336) );
  XOR U505 ( .A(B[848]), .B(n337), .Z(O[849]) );
  AND U506 ( .A(S), .B(n338), .Z(n337) );
  XOR U507 ( .A(B[849]), .B(B[848]), .Z(n338) );
  XOR U508 ( .A(B[847]), .B(n339), .Z(O[848]) );
  AND U509 ( .A(S), .B(n340), .Z(n339) );
  XOR U510 ( .A(B[848]), .B(B[847]), .Z(n340) );
  XOR U511 ( .A(B[846]), .B(n341), .Z(O[847]) );
  AND U512 ( .A(S), .B(n342), .Z(n341) );
  XOR U513 ( .A(B[847]), .B(B[846]), .Z(n342) );
  XOR U514 ( .A(B[845]), .B(n343), .Z(O[846]) );
  AND U515 ( .A(S), .B(n344), .Z(n343) );
  XOR U516 ( .A(B[846]), .B(B[845]), .Z(n344) );
  XOR U517 ( .A(B[844]), .B(n345), .Z(O[845]) );
  AND U518 ( .A(S), .B(n346), .Z(n345) );
  XOR U519 ( .A(B[845]), .B(B[844]), .Z(n346) );
  XOR U520 ( .A(B[843]), .B(n347), .Z(O[844]) );
  AND U521 ( .A(S), .B(n348), .Z(n347) );
  XOR U522 ( .A(B[844]), .B(B[843]), .Z(n348) );
  XOR U523 ( .A(B[842]), .B(n349), .Z(O[843]) );
  AND U524 ( .A(S), .B(n350), .Z(n349) );
  XOR U525 ( .A(B[843]), .B(B[842]), .Z(n350) );
  XOR U526 ( .A(B[841]), .B(n351), .Z(O[842]) );
  AND U527 ( .A(S), .B(n352), .Z(n351) );
  XOR U528 ( .A(B[842]), .B(B[841]), .Z(n352) );
  XOR U529 ( .A(B[840]), .B(n353), .Z(O[841]) );
  AND U530 ( .A(S), .B(n354), .Z(n353) );
  XOR U531 ( .A(B[841]), .B(B[840]), .Z(n354) );
  XOR U532 ( .A(B[839]), .B(n355), .Z(O[840]) );
  AND U533 ( .A(S), .B(n356), .Z(n355) );
  XOR U534 ( .A(B[840]), .B(B[839]), .Z(n356) );
  XOR U535 ( .A(B[82]), .B(n357), .Z(O[83]) );
  AND U536 ( .A(S), .B(n358), .Z(n357) );
  XOR U537 ( .A(B[83]), .B(B[82]), .Z(n358) );
  XOR U538 ( .A(B[838]), .B(n359), .Z(O[839]) );
  AND U539 ( .A(S), .B(n360), .Z(n359) );
  XOR U540 ( .A(B[839]), .B(B[838]), .Z(n360) );
  XOR U541 ( .A(B[837]), .B(n361), .Z(O[838]) );
  AND U542 ( .A(S), .B(n362), .Z(n361) );
  XOR U543 ( .A(B[838]), .B(B[837]), .Z(n362) );
  XOR U544 ( .A(B[836]), .B(n363), .Z(O[837]) );
  AND U545 ( .A(S), .B(n364), .Z(n363) );
  XOR U546 ( .A(B[837]), .B(B[836]), .Z(n364) );
  XOR U547 ( .A(B[835]), .B(n365), .Z(O[836]) );
  AND U548 ( .A(S), .B(n366), .Z(n365) );
  XOR U549 ( .A(B[836]), .B(B[835]), .Z(n366) );
  XOR U550 ( .A(B[834]), .B(n367), .Z(O[835]) );
  AND U551 ( .A(S), .B(n368), .Z(n367) );
  XOR U552 ( .A(B[835]), .B(B[834]), .Z(n368) );
  XOR U553 ( .A(B[833]), .B(n369), .Z(O[834]) );
  AND U554 ( .A(S), .B(n370), .Z(n369) );
  XOR U555 ( .A(B[834]), .B(B[833]), .Z(n370) );
  XOR U556 ( .A(B[832]), .B(n371), .Z(O[833]) );
  AND U557 ( .A(S), .B(n372), .Z(n371) );
  XOR U558 ( .A(B[833]), .B(B[832]), .Z(n372) );
  XOR U559 ( .A(B[831]), .B(n373), .Z(O[832]) );
  AND U560 ( .A(S), .B(n374), .Z(n373) );
  XOR U561 ( .A(B[832]), .B(B[831]), .Z(n374) );
  XOR U562 ( .A(B[830]), .B(n375), .Z(O[831]) );
  AND U563 ( .A(S), .B(n376), .Z(n375) );
  XOR U564 ( .A(B[831]), .B(B[830]), .Z(n376) );
  XOR U565 ( .A(B[829]), .B(n377), .Z(O[830]) );
  AND U566 ( .A(S), .B(n378), .Z(n377) );
  XOR U567 ( .A(B[830]), .B(B[829]), .Z(n378) );
  XOR U568 ( .A(B[81]), .B(n379), .Z(O[82]) );
  AND U569 ( .A(S), .B(n380), .Z(n379) );
  XOR U570 ( .A(B[82]), .B(B[81]), .Z(n380) );
  XOR U571 ( .A(B[828]), .B(n381), .Z(O[829]) );
  AND U572 ( .A(S), .B(n382), .Z(n381) );
  XOR U573 ( .A(B[829]), .B(B[828]), .Z(n382) );
  XOR U574 ( .A(B[827]), .B(n383), .Z(O[828]) );
  AND U575 ( .A(S), .B(n384), .Z(n383) );
  XOR U576 ( .A(B[828]), .B(B[827]), .Z(n384) );
  XOR U577 ( .A(B[826]), .B(n385), .Z(O[827]) );
  AND U578 ( .A(S), .B(n386), .Z(n385) );
  XOR U579 ( .A(B[827]), .B(B[826]), .Z(n386) );
  XOR U580 ( .A(B[825]), .B(n387), .Z(O[826]) );
  AND U581 ( .A(S), .B(n388), .Z(n387) );
  XOR U582 ( .A(B[826]), .B(B[825]), .Z(n388) );
  XOR U583 ( .A(B[824]), .B(n389), .Z(O[825]) );
  AND U584 ( .A(S), .B(n390), .Z(n389) );
  XOR U585 ( .A(B[825]), .B(B[824]), .Z(n390) );
  XOR U586 ( .A(B[823]), .B(n391), .Z(O[824]) );
  AND U587 ( .A(S), .B(n392), .Z(n391) );
  XOR U588 ( .A(B[824]), .B(B[823]), .Z(n392) );
  XOR U589 ( .A(B[822]), .B(n393), .Z(O[823]) );
  AND U590 ( .A(S), .B(n394), .Z(n393) );
  XOR U591 ( .A(B[823]), .B(B[822]), .Z(n394) );
  XOR U592 ( .A(B[821]), .B(n395), .Z(O[822]) );
  AND U593 ( .A(S), .B(n396), .Z(n395) );
  XOR U594 ( .A(B[822]), .B(B[821]), .Z(n396) );
  XOR U595 ( .A(B[820]), .B(n397), .Z(O[821]) );
  AND U596 ( .A(S), .B(n398), .Z(n397) );
  XOR U597 ( .A(B[821]), .B(B[820]), .Z(n398) );
  XOR U598 ( .A(B[819]), .B(n399), .Z(O[820]) );
  AND U599 ( .A(S), .B(n400), .Z(n399) );
  XOR U600 ( .A(B[820]), .B(B[819]), .Z(n400) );
  XOR U601 ( .A(B[80]), .B(n401), .Z(O[81]) );
  AND U602 ( .A(S), .B(n402), .Z(n401) );
  XOR U603 ( .A(B[81]), .B(B[80]), .Z(n402) );
  XOR U604 ( .A(B[818]), .B(n403), .Z(O[819]) );
  AND U605 ( .A(S), .B(n404), .Z(n403) );
  XOR U606 ( .A(B[819]), .B(B[818]), .Z(n404) );
  XOR U607 ( .A(B[817]), .B(n405), .Z(O[818]) );
  AND U608 ( .A(S), .B(n406), .Z(n405) );
  XOR U609 ( .A(B[818]), .B(B[817]), .Z(n406) );
  XOR U610 ( .A(B[816]), .B(n407), .Z(O[817]) );
  AND U611 ( .A(S), .B(n408), .Z(n407) );
  XOR U612 ( .A(B[817]), .B(B[816]), .Z(n408) );
  XOR U613 ( .A(B[815]), .B(n409), .Z(O[816]) );
  AND U614 ( .A(S), .B(n410), .Z(n409) );
  XOR U615 ( .A(B[816]), .B(B[815]), .Z(n410) );
  XOR U616 ( .A(B[814]), .B(n411), .Z(O[815]) );
  AND U617 ( .A(S), .B(n412), .Z(n411) );
  XOR U618 ( .A(B[815]), .B(B[814]), .Z(n412) );
  XOR U619 ( .A(B[813]), .B(n413), .Z(O[814]) );
  AND U620 ( .A(S), .B(n414), .Z(n413) );
  XOR U621 ( .A(B[814]), .B(B[813]), .Z(n414) );
  XOR U622 ( .A(B[812]), .B(n415), .Z(O[813]) );
  AND U623 ( .A(S), .B(n416), .Z(n415) );
  XOR U624 ( .A(B[813]), .B(B[812]), .Z(n416) );
  XOR U625 ( .A(B[811]), .B(n417), .Z(O[812]) );
  AND U626 ( .A(S), .B(n418), .Z(n417) );
  XOR U627 ( .A(B[812]), .B(B[811]), .Z(n418) );
  XOR U628 ( .A(B[810]), .B(n419), .Z(O[811]) );
  AND U629 ( .A(S), .B(n420), .Z(n419) );
  XOR U630 ( .A(B[811]), .B(B[810]), .Z(n420) );
  XOR U631 ( .A(B[809]), .B(n421), .Z(O[810]) );
  AND U632 ( .A(S), .B(n422), .Z(n421) );
  XOR U633 ( .A(B[810]), .B(B[809]), .Z(n422) );
  XOR U634 ( .A(B[79]), .B(n423), .Z(O[80]) );
  AND U635 ( .A(S), .B(n424), .Z(n423) );
  XOR U636 ( .A(B[80]), .B(B[79]), .Z(n424) );
  XOR U637 ( .A(B[808]), .B(n425), .Z(O[809]) );
  AND U638 ( .A(S), .B(n426), .Z(n425) );
  XOR U639 ( .A(B[809]), .B(B[808]), .Z(n426) );
  XOR U640 ( .A(B[807]), .B(n427), .Z(O[808]) );
  AND U641 ( .A(S), .B(n428), .Z(n427) );
  XOR U642 ( .A(B[808]), .B(B[807]), .Z(n428) );
  XOR U643 ( .A(B[806]), .B(n429), .Z(O[807]) );
  AND U644 ( .A(S), .B(n430), .Z(n429) );
  XOR U645 ( .A(B[807]), .B(B[806]), .Z(n430) );
  XOR U646 ( .A(B[805]), .B(n431), .Z(O[806]) );
  AND U647 ( .A(S), .B(n432), .Z(n431) );
  XOR U648 ( .A(B[806]), .B(B[805]), .Z(n432) );
  XOR U649 ( .A(B[804]), .B(n433), .Z(O[805]) );
  AND U650 ( .A(S), .B(n434), .Z(n433) );
  XOR U651 ( .A(B[805]), .B(B[804]), .Z(n434) );
  XOR U652 ( .A(B[803]), .B(n435), .Z(O[804]) );
  AND U653 ( .A(S), .B(n436), .Z(n435) );
  XOR U654 ( .A(B[804]), .B(B[803]), .Z(n436) );
  XOR U655 ( .A(B[802]), .B(n437), .Z(O[803]) );
  AND U656 ( .A(S), .B(n438), .Z(n437) );
  XOR U657 ( .A(B[803]), .B(B[802]), .Z(n438) );
  XOR U658 ( .A(B[801]), .B(n439), .Z(O[802]) );
  AND U659 ( .A(S), .B(n440), .Z(n439) );
  XOR U660 ( .A(B[802]), .B(B[801]), .Z(n440) );
  XOR U661 ( .A(B[800]), .B(n441), .Z(O[801]) );
  AND U662 ( .A(S), .B(n442), .Z(n441) );
  XOR U663 ( .A(B[801]), .B(B[800]), .Z(n442) );
  XOR U664 ( .A(B[799]), .B(n443), .Z(O[800]) );
  AND U665 ( .A(S), .B(n444), .Z(n443) );
  XOR U666 ( .A(B[800]), .B(B[799]), .Z(n444) );
  XOR U667 ( .A(B[6]), .B(n445), .Z(O[7]) );
  AND U668 ( .A(S), .B(n446), .Z(n445) );
  XOR U669 ( .A(B[7]), .B(B[6]), .Z(n446) );
  XOR U670 ( .A(B[78]), .B(n447), .Z(O[79]) );
  AND U671 ( .A(S), .B(n448), .Z(n447) );
  XOR U672 ( .A(B[79]), .B(B[78]), .Z(n448) );
  XOR U673 ( .A(B[798]), .B(n449), .Z(O[799]) );
  AND U674 ( .A(S), .B(n450), .Z(n449) );
  XOR U675 ( .A(B[799]), .B(B[798]), .Z(n450) );
  XOR U676 ( .A(B[797]), .B(n451), .Z(O[798]) );
  AND U677 ( .A(S), .B(n452), .Z(n451) );
  XOR U678 ( .A(B[798]), .B(B[797]), .Z(n452) );
  XOR U679 ( .A(B[796]), .B(n453), .Z(O[797]) );
  AND U680 ( .A(S), .B(n454), .Z(n453) );
  XOR U681 ( .A(B[797]), .B(B[796]), .Z(n454) );
  XOR U682 ( .A(B[795]), .B(n455), .Z(O[796]) );
  AND U683 ( .A(S), .B(n456), .Z(n455) );
  XOR U684 ( .A(B[796]), .B(B[795]), .Z(n456) );
  XOR U685 ( .A(B[794]), .B(n457), .Z(O[795]) );
  AND U686 ( .A(S), .B(n458), .Z(n457) );
  XOR U687 ( .A(B[795]), .B(B[794]), .Z(n458) );
  XOR U688 ( .A(B[793]), .B(n459), .Z(O[794]) );
  AND U689 ( .A(S), .B(n460), .Z(n459) );
  XOR U690 ( .A(B[794]), .B(B[793]), .Z(n460) );
  XOR U691 ( .A(B[792]), .B(n461), .Z(O[793]) );
  AND U692 ( .A(S), .B(n462), .Z(n461) );
  XOR U693 ( .A(B[793]), .B(B[792]), .Z(n462) );
  XOR U694 ( .A(B[791]), .B(n463), .Z(O[792]) );
  AND U695 ( .A(S), .B(n464), .Z(n463) );
  XOR U696 ( .A(B[792]), .B(B[791]), .Z(n464) );
  XOR U697 ( .A(B[790]), .B(n465), .Z(O[791]) );
  AND U698 ( .A(S), .B(n466), .Z(n465) );
  XOR U699 ( .A(B[791]), .B(B[790]), .Z(n466) );
  XOR U700 ( .A(B[789]), .B(n467), .Z(O[790]) );
  AND U701 ( .A(S), .B(n468), .Z(n467) );
  XOR U702 ( .A(B[790]), .B(B[789]), .Z(n468) );
  XOR U703 ( .A(B[77]), .B(n469), .Z(O[78]) );
  AND U704 ( .A(S), .B(n470), .Z(n469) );
  XOR U705 ( .A(B[78]), .B(B[77]), .Z(n470) );
  XOR U706 ( .A(B[788]), .B(n471), .Z(O[789]) );
  AND U707 ( .A(S), .B(n472), .Z(n471) );
  XOR U708 ( .A(B[789]), .B(B[788]), .Z(n472) );
  XOR U709 ( .A(B[787]), .B(n473), .Z(O[788]) );
  AND U710 ( .A(S), .B(n474), .Z(n473) );
  XOR U711 ( .A(B[788]), .B(B[787]), .Z(n474) );
  XOR U712 ( .A(B[786]), .B(n475), .Z(O[787]) );
  AND U713 ( .A(S), .B(n476), .Z(n475) );
  XOR U714 ( .A(B[787]), .B(B[786]), .Z(n476) );
  XOR U715 ( .A(B[785]), .B(n477), .Z(O[786]) );
  AND U716 ( .A(S), .B(n478), .Z(n477) );
  XOR U717 ( .A(B[786]), .B(B[785]), .Z(n478) );
  XOR U718 ( .A(B[784]), .B(n479), .Z(O[785]) );
  AND U719 ( .A(S), .B(n480), .Z(n479) );
  XOR U720 ( .A(B[785]), .B(B[784]), .Z(n480) );
  XOR U721 ( .A(B[783]), .B(n481), .Z(O[784]) );
  AND U722 ( .A(S), .B(n482), .Z(n481) );
  XOR U723 ( .A(B[784]), .B(B[783]), .Z(n482) );
  XOR U724 ( .A(B[782]), .B(n483), .Z(O[783]) );
  AND U725 ( .A(S), .B(n484), .Z(n483) );
  XOR U726 ( .A(B[783]), .B(B[782]), .Z(n484) );
  XOR U727 ( .A(B[781]), .B(n485), .Z(O[782]) );
  AND U728 ( .A(S), .B(n486), .Z(n485) );
  XOR U729 ( .A(B[782]), .B(B[781]), .Z(n486) );
  XOR U730 ( .A(B[780]), .B(n487), .Z(O[781]) );
  AND U731 ( .A(S), .B(n488), .Z(n487) );
  XOR U732 ( .A(B[781]), .B(B[780]), .Z(n488) );
  XOR U733 ( .A(B[779]), .B(n489), .Z(O[780]) );
  AND U734 ( .A(S), .B(n490), .Z(n489) );
  XOR U735 ( .A(B[780]), .B(B[779]), .Z(n490) );
  XOR U736 ( .A(B[76]), .B(n491), .Z(O[77]) );
  AND U737 ( .A(S), .B(n492), .Z(n491) );
  XOR U738 ( .A(B[77]), .B(B[76]), .Z(n492) );
  XOR U739 ( .A(B[778]), .B(n493), .Z(O[779]) );
  AND U740 ( .A(S), .B(n494), .Z(n493) );
  XOR U741 ( .A(B[779]), .B(B[778]), .Z(n494) );
  XOR U742 ( .A(B[777]), .B(n495), .Z(O[778]) );
  AND U743 ( .A(S), .B(n496), .Z(n495) );
  XOR U744 ( .A(B[778]), .B(B[777]), .Z(n496) );
  XOR U745 ( .A(B[776]), .B(n497), .Z(O[777]) );
  AND U746 ( .A(S), .B(n498), .Z(n497) );
  XOR U747 ( .A(B[777]), .B(B[776]), .Z(n498) );
  XOR U748 ( .A(B[775]), .B(n499), .Z(O[776]) );
  AND U749 ( .A(S), .B(n500), .Z(n499) );
  XOR U750 ( .A(B[776]), .B(B[775]), .Z(n500) );
  XOR U751 ( .A(B[774]), .B(n501), .Z(O[775]) );
  AND U752 ( .A(S), .B(n502), .Z(n501) );
  XOR U753 ( .A(B[775]), .B(B[774]), .Z(n502) );
  XOR U754 ( .A(B[773]), .B(n503), .Z(O[774]) );
  AND U755 ( .A(S), .B(n504), .Z(n503) );
  XOR U756 ( .A(B[774]), .B(B[773]), .Z(n504) );
  XOR U757 ( .A(B[772]), .B(n505), .Z(O[773]) );
  AND U758 ( .A(S), .B(n506), .Z(n505) );
  XOR U759 ( .A(B[773]), .B(B[772]), .Z(n506) );
  XOR U760 ( .A(B[771]), .B(n507), .Z(O[772]) );
  AND U761 ( .A(S), .B(n508), .Z(n507) );
  XOR U762 ( .A(B[772]), .B(B[771]), .Z(n508) );
  XOR U763 ( .A(B[770]), .B(n509), .Z(O[771]) );
  AND U764 ( .A(S), .B(n510), .Z(n509) );
  XOR U765 ( .A(B[771]), .B(B[770]), .Z(n510) );
  XOR U766 ( .A(B[769]), .B(n511), .Z(O[770]) );
  AND U767 ( .A(S), .B(n512), .Z(n511) );
  XOR U768 ( .A(B[770]), .B(B[769]), .Z(n512) );
  XOR U769 ( .A(B[75]), .B(n513), .Z(O[76]) );
  AND U770 ( .A(S), .B(n514), .Z(n513) );
  XOR U771 ( .A(B[76]), .B(B[75]), .Z(n514) );
  XOR U772 ( .A(B[768]), .B(n515), .Z(O[769]) );
  AND U773 ( .A(S), .B(n516), .Z(n515) );
  XOR U774 ( .A(B[769]), .B(B[768]), .Z(n516) );
  XOR U775 ( .A(B[767]), .B(n517), .Z(O[768]) );
  AND U776 ( .A(S), .B(n518), .Z(n517) );
  XOR U777 ( .A(B[768]), .B(B[767]), .Z(n518) );
  XOR U778 ( .A(B[766]), .B(n519), .Z(O[767]) );
  AND U779 ( .A(S), .B(n520), .Z(n519) );
  XOR U780 ( .A(B[767]), .B(B[766]), .Z(n520) );
  XOR U781 ( .A(B[765]), .B(n521), .Z(O[766]) );
  AND U782 ( .A(S), .B(n522), .Z(n521) );
  XOR U783 ( .A(B[766]), .B(B[765]), .Z(n522) );
  XOR U784 ( .A(B[764]), .B(n523), .Z(O[765]) );
  AND U785 ( .A(S), .B(n524), .Z(n523) );
  XOR U786 ( .A(B[765]), .B(B[764]), .Z(n524) );
  XOR U787 ( .A(B[763]), .B(n525), .Z(O[764]) );
  AND U788 ( .A(S), .B(n526), .Z(n525) );
  XOR U789 ( .A(B[764]), .B(B[763]), .Z(n526) );
  XOR U790 ( .A(B[762]), .B(n527), .Z(O[763]) );
  AND U791 ( .A(S), .B(n528), .Z(n527) );
  XOR U792 ( .A(B[763]), .B(B[762]), .Z(n528) );
  XOR U793 ( .A(B[761]), .B(n529), .Z(O[762]) );
  AND U794 ( .A(S), .B(n530), .Z(n529) );
  XOR U795 ( .A(B[762]), .B(B[761]), .Z(n530) );
  XOR U796 ( .A(B[760]), .B(n531), .Z(O[761]) );
  AND U797 ( .A(S), .B(n532), .Z(n531) );
  XOR U798 ( .A(B[761]), .B(B[760]), .Z(n532) );
  XOR U799 ( .A(B[759]), .B(n533), .Z(O[760]) );
  AND U800 ( .A(S), .B(n534), .Z(n533) );
  XOR U801 ( .A(B[760]), .B(B[759]), .Z(n534) );
  XOR U802 ( .A(B[74]), .B(n535), .Z(O[75]) );
  AND U803 ( .A(S), .B(n536), .Z(n535) );
  XOR U804 ( .A(B[75]), .B(B[74]), .Z(n536) );
  XOR U805 ( .A(B[758]), .B(n537), .Z(O[759]) );
  AND U806 ( .A(S), .B(n538), .Z(n537) );
  XOR U807 ( .A(B[759]), .B(B[758]), .Z(n538) );
  XOR U808 ( .A(B[757]), .B(n539), .Z(O[758]) );
  AND U809 ( .A(S), .B(n540), .Z(n539) );
  XOR U810 ( .A(B[758]), .B(B[757]), .Z(n540) );
  XOR U811 ( .A(B[756]), .B(n541), .Z(O[757]) );
  AND U812 ( .A(S), .B(n542), .Z(n541) );
  XOR U813 ( .A(B[757]), .B(B[756]), .Z(n542) );
  XOR U814 ( .A(B[755]), .B(n543), .Z(O[756]) );
  AND U815 ( .A(S), .B(n544), .Z(n543) );
  XOR U816 ( .A(B[756]), .B(B[755]), .Z(n544) );
  XOR U817 ( .A(B[754]), .B(n545), .Z(O[755]) );
  AND U818 ( .A(S), .B(n546), .Z(n545) );
  XOR U819 ( .A(B[755]), .B(B[754]), .Z(n546) );
  XOR U820 ( .A(B[753]), .B(n547), .Z(O[754]) );
  AND U821 ( .A(S), .B(n548), .Z(n547) );
  XOR U822 ( .A(B[754]), .B(B[753]), .Z(n548) );
  XOR U823 ( .A(B[752]), .B(n549), .Z(O[753]) );
  AND U824 ( .A(S), .B(n550), .Z(n549) );
  XOR U825 ( .A(B[753]), .B(B[752]), .Z(n550) );
  XOR U826 ( .A(B[751]), .B(n551), .Z(O[752]) );
  AND U827 ( .A(S), .B(n552), .Z(n551) );
  XOR U828 ( .A(B[752]), .B(B[751]), .Z(n552) );
  XOR U829 ( .A(B[750]), .B(n553), .Z(O[751]) );
  AND U830 ( .A(S), .B(n554), .Z(n553) );
  XOR U831 ( .A(B[751]), .B(B[750]), .Z(n554) );
  XOR U832 ( .A(B[749]), .B(n555), .Z(O[750]) );
  AND U833 ( .A(S), .B(n556), .Z(n555) );
  XOR U834 ( .A(B[750]), .B(B[749]), .Z(n556) );
  XOR U835 ( .A(B[73]), .B(n557), .Z(O[74]) );
  AND U836 ( .A(S), .B(n558), .Z(n557) );
  XOR U837 ( .A(B[74]), .B(B[73]), .Z(n558) );
  XOR U838 ( .A(B[748]), .B(n559), .Z(O[749]) );
  AND U839 ( .A(S), .B(n560), .Z(n559) );
  XOR U840 ( .A(B[749]), .B(B[748]), .Z(n560) );
  XOR U841 ( .A(B[747]), .B(n561), .Z(O[748]) );
  AND U842 ( .A(S), .B(n562), .Z(n561) );
  XOR U843 ( .A(B[748]), .B(B[747]), .Z(n562) );
  XOR U844 ( .A(B[746]), .B(n563), .Z(O[747]) );
  AND U845 ( .A(S), .B(n564), .Z(n563) );
  XOR U846 ( .A(B[747]), .B(B[746]), .Z(n564) );
  XOR U847 ( .A(B[745]), .B(n565), .Z(O[746]) );
  AND U848 ( .A(S), .B(n566), .Z(n565) );
  XOR U849 ( .A(B[746]), .B(B[745]), .Z(n566) );
  XOR U850 ( .A(B[744]), .B(n567), .Z(O[745]) );
  AND U851 ( .A(S), .B(n568), .Z(n567) );
  XOR U852 ( .A(B[745]), .B(B[744]), .Z(n568) );
  XOR U853 ( .A(B[743]), .B(n569), .Z(O[744]) );
  AND U854 ( .A(S), .B(n570), .Z(n569) );
  XOR U855 ( .A(B[744]), .B(B[743]), .Z(n570) );
  XOR U856 ( .A(B[742]), .B(n571), .Z(O[743]) );
  AND U857 ( .A(S), .B(n572), .Z(n571) );
  XOR U858 ( .A(B[743]), .B(B[742]), .Z(n572) );
  XOR U859 ( .A(B[741]), .B(n573), .Z(O[742]) );
  AND U860 ( .A(S), .B(n574), .Z(n573) );
  XOR U861 ( .A(B[742]), .B(B[741]), .Z(n574) );
  XOR U862 ( .A(B[740]), .B(n575), .Z(O[741]) );
  AND U863 ( .A(S), .B(n576), .Z(n575) );
  XOR U864 ( .A(B[741]), .B(B[740]), .Z(n576) );
  XOR U865 ( .A(B[739]), .B(n577), .Z(O[740]) );
  AND U866 ( .A(S), .B(n578), .Z(n577) );
  XOR U867 ( .A(B[740]), .B(B[739]), .Z(n578) );
  XOR U868 ( .A(B[72]), .B(n579), .Z(O[73]) );
  AND U869 ( .A(S), .B(n580), .Z(n579) );
  XOR U870 ( .A(B[73]), .B(B[72]), .Z(n580) );
  XOR U871 ( .A(B[738]), .B(n581), .Z(O[739]) );
  AND U872 ( .A(S), .B(n582), .Z(n581) );
  XOR U873 ( .A(B[739]), .B(B[738]), .Z(n582) );
  XOR U874 ( .A(B[737]), .B(n583), .Z(O[738]) );
  AND U875 ( .A(S), .B(n584), .Z(n583) );
  XOR U876 ( .A(B[738]), .B(B[737]), .Z(n584) );
  XOR U877 ( .A(B[736]), .B(n585), .Z(O[737]) );
  AND U878 ( .A(S), .B(n586), .Z(n585) );
  XOR U879 ( .A(B[737]), .B(B[736]), .Z(n586) );
  XOR U880 ( .A(B[735]), .B(n587), .Z(O[736]) );
  AND U881 ( .A(S), .B(n588), .Z(n587) );
  XOR U882 ( .A(B[736]), .B(B[735]), .Z(n588) );
  XOR U883 ( .A(B[734]), .B(n589), .Z(O[735]) );
  AND U884 ( .A(S), .B(n590), .Z(n589) );
  XOR U885 ( .A(B[735]), .B(B[734]), .Z(n590) );
  XOR U886 ( .A(B[733]), .B(n591), .Z(O[734]) );
  AND U887 ( .A(S), .B(n592), .Z(n591) );
  XOR U888 ( .A(B[734]), .B(B[733]), .Z(n592) );
  XOR U889 ( .A(B[732]), .B(n593), .Z(O[733]) );
  AND U890 ( .A(S), .B(n594), .Z(n593) );
  XOR U891 ( .A(B[733]), .B(B[732]), .Z(n594) );
  XOR U892 ( .A(B[731]), .B(n595), .Z(O[732]) );
  AND U893 ( .A(S), .B(n596), .Z(n595) );
  XOR U894 ( .A(B[732]), .B(B[731]), .Z(n596) );
  XOR U895 ( .A(B[730]), .B(n597), .Z(O[731]) );
  AND U896 ( .A(S), .B(n598), .Z(n597) );
  XOR U897 ( .A(B[731]), .B(B[730]), .Z(n598) );
  XOR U898 ( .A(B[729]), .B(n599), .Z(O[730]) );
  AND U899 ( .A(S), .B(n600), .Z(n599) );
  XOR U900 ( .A(B[730]), .B(B[729]), .Z(n600) );
  XOR U901 ( .A(B[71]), .B(n601), .Z(O[72]) );
  AND U902 ( .A(S), .B(n602), .Z(n601) );
  XOR U903 ( .A(B[72]), .B(B[71]), .Z(n602) );
  XOR U904 ( .A(B[728]), .B(n603), .Z(O[729]) );
  AND U905 ( .A(S), .B(n604), .Z(n603) );
  XOR U906 ( .A(B[729]), .B(B[728]), .Z(n604) );
  XOR U907 ( .A(B[727]), .B(n605), .Z(O[728]) );
  AND U908 ( .A(S), .B(n606), .Z(n605) );
  XOR U909 ( .A(B[728]), .B(B[727]), .Z(n606) );
  XOR U910 ( .A(B[726]), .B(n607), .Z(O[727]) );
  AND U911 ( .A(S), .B(n608), .Z(n607) );
  XOR U912 ( .A(B[727]), .B(B[726]), .Z(n608) );
  XOR U913 ( .A(B[725]), .B(n609), .Z(O[726]) );
  AND U914 ( .A(S), .B(n610), .Z(n609) );
  XOR U915 ( .A(B[726]), .B(B[725]), .Z(n610) );
  XOR U916 ( .A(B[724]), .B(n611), .Z(O[725]) );
  AND U917 ( .A(S), .B(n612), .Z(n611) );
  XOR U918 ( .A(B[725]), .B(B[724]), .Z(n612) );
  XOR U919 ( .A(B[723]), .B(n613), .Z(O[724]) );
  AND U920 ( .A(S), .B(n614), .Z(n613) );
  XOR U921 ( .A(B[724]), .B(B[723]), .Z(n614) );
  XOR U922 ( .A(B[722]), .B(n615), .Z(O[723]) );
  AND U923 ( .A(S), .B(n616), .Z(n615) );
  XOR U924 ( .A(B[723]), .B(B[722]), .Z(n616) );
  XOR U925 ( .A(B[721]), .B(n617), .Z(O[722]) );
  AND U926 ( .A(S), .B(n618), .Z(n617) );
  XOR U927 ( .A(B[722]), .B(B[721]), .Z(n618) );
  XOR U928 ( .A(B[720]), .B(n619), .Z(O[721]) );
  AND U929 ( .A(S), .B(n620), .Z(n619) );
  XOR U930 ( .A(B[721]), .B(B[720]), .Z(n620) );
  XOR U931 ( .A(B[719]), .B(n621), .Z(O[720]) );
  AND U932 ( .A(S), .B(n622), .Z(n621) );
  XOR U933 ( .A(B[720]), .B(B[719]), .Z(n622) );
  XOR U934 ( .A(B[70]), .B(n623), .Z(O[71]) );
  AND U935 ( .A(S), .B(n624), .Z(n623) );
  XOR U936 ( .A(B[71]), .B(B[70]), .Z(n624) );
  XOR U937 ( .A(B[718]), .B(n625), .Z(O[719]) );
  AND U938 ( .A(S), .B(n626), .Z(n625) );
  XOR U939 ( .A(B[719]), .B(B[718]), .Z(n626) );
  XOR U940 ( .A(B[717]), .B(n627), .Z(O[718]) );
  AND U941 ( .A(S), .B(n628), .Z(n627) );
  XOR U942 ( .A(B[718]), .B(B[717]), .Z(n628) );
  XOR U943 ( .A(B[716]), .B(n629), .Z(O[717]) );
  AND U944 ( .A(S), .B(n630), .Z(n629) );
  XOR U945 ( .A(B[717]), .B(B[716]), .Z(n630) );
  XOR U946 ( .A(B[715]), .B(n631), .Z(O[716]) );
  AND U947 ( .A(S), .B(n632), .Z(n631) );
  XOR U948 ( .A(B[716]), .B(B[715]), .Z(n632) );
  XOR U949 ( .A(B[714]), .B(n633), .Z(O[715]) );
  AND U950 ( .A(S), .B(n634), .Z(n633) );
  XOR U951 ( .A(B[715]), .B(B[714]), .Z(n634) );
  XOR U952 ( .A(B[713]), .B(n635), .Z(O[714]) );
  AND U953 ( .A(S), .B(n636), .Z(n635) );
  XOR U954 ( .A(B[714]), .B(B[713]), .Z(n636) );
  XOR U955 ( .A(B[712]), .B(n637), .Z(O[713]) );
  AND U956 ( .A(S), .B(n638), .Z(n637) );
  XOR U957 ( .A(B[713]), .B(B[712]), .Z(n638) );
  XOR U958 ( .A(B[711]), .B(n639), .Z(O[712]) );
  AND U959 ( .A(S), .B(n640), .Z(n639) );
  XOR U960 ( .A(B[712]), .B(B[711]), .Z(n640) );
  XOR U961 ( .A(B[710]), .B(n641), .Z(O[711]) );
  AND U962 ( .A(S), .B(n642), .Z(n641) );
  XOR U963 ( .A(B[711]), .B(B[710]), .Z(n642) );
  XOR U964 ( .A(B[709]), .B(n643), .Z(O[710]) );
  AND U965 ( .A(S), .B(n644), .Z(n643) );
  XOR U966 ( .A(B[710]), .B(B[709]), .Z(n644) );
  XOR U967 ( .A(B[69]), .B(n645), .Z(O[70]) );
  AND U968 ( .A(S), .B(n646), .Z(n645) );
  XOR U969 ( .A(B[70]), .B(B[69]), .Z(n646) );
  XOR U970 ( .A(B[708]), .B(n647), .Z(O[709]) );
  AND U971 ( .A(S), .B(n648), .Z(n647) );
  XOR U972 ( .A(B[709]), .B(B[708]), .Z(n648) );
  XOR U973 ( .A(B[707]), .B(n649), .Z(O[708]) );
  AND U974 ( .A(S), .B(n650), .Z(n649) );
  XOR U975 ( .A(B[708]), .B(B[707]), .Z(n650) );
  XOR U976 ( .A(B[706]), .B(n651), .Z(O[707]) );
  AND U977 ( .A(S), .B(n652), .Z(n651) );
  XOR U978 ( .A(B[707]), .B(B[706]), .Z(n652) );
  XOR U979 ( .A(B[705]), .B(n653), .Z(O[706]) );
  AND U980 ( .A(S), .B(n654), .Z(n653) );
  XOR U981 ( .A(B[706]), .B(B[705]), .Z(n654) );
  XOR U982 ( .A(B[704]), .B(n655), .Z(O[705]) );
  AND U983 ( .A(S), .B(n656), .Z(n655) );
  XOR U984 ( .A(B[705]), .B(B[704]), .Z(n656) );
  XOR U985 ( .A(B[703]), .B(n657), .Z(O[704]) );
  AND U986 ( .A(S), .B(n658), .Z(n657) );
  XOR U987 ( .A(B[704]), .B(B[703]), .Z(n658) );
  XOR U988 ( .A(B[702]), .B(n659), .Z(O[703]) );
  AND U989 ( .A(S), .B(n660), .Z(n659) );
  XOR U990 ( .A(B[703]), .B(B[702]), .Z(n660) );
  XOR U991 ( .A(B[701]), .B(n661), .Z(O[702]) );
  AND U992 ( .A(S), .B(n662), .Z(n661) );
  XOR U993 ( .A(B[702]), .B(B[701]), .Z(n662) );
  XOR U994 ( .A(B[700]), .B(n663), .Z(O[701]) );
  AND U995 ( .A(S), .B(n664), .Z(n663) );
  XOR U996 ( .A(B[701]), .B(B[700]), .Z(n664) );
  XOR U997 ( .A(B[699]), .B(n665), .Z(O[700]) );
  AND U998 ( .A(S), .B(n666), .Z(n665) );
  XOR U999 ( .A(B[700]), .B(B[699]), .Z(n666) );
  XOR U1000 ( .A(B[5]), .B(n667), .Z(O[6]) );
  AND U1001 ( .A(S), .B(n668), .Z(n667) );
  XOR U1002 ( .A(B[6]), .B(B[5]), .Z(n668) );
  XOR U1003 ( .A(B[68]), .B(n669), .Z(O[69]) );
  AND U1004 ( .A(S), .B(n670), .Z(n669) );
  XOR U1005 ( .A(B[69]), .B(B[68]), .Z(n670) );
  XOR U1006 ( .A(B[698]), .B(n671), .Z(O[699]) );
  AND U1007 ( .A(S), .B(n672), .Z(n671) );
  XOR U1008 ( .A(B[699]), .B(B[698]), .Z(n672) );
  XOR U1009 ( .A(B[697]), .B(n673), .Z(O[698]) );
  AND U1010 ( .A(S), .B(n674), .Z(n673) );
  XOR U1011 ( .A(B[698]), .B(B[697]), .Z(n674) );
  XOR U1012 ( .A(B[696]), .B(n675), .Z(O[697]) );
  AND U1013 ( .A(S), .B(n676), .Z(n675) );
  XOR U1014 ( .A(B[697]), .B(B[696]), .Z(n676) );
  XOR U1015 ( .A(B[695]), .B(n677), .Z(O[696]) );
  AND U1016 ( .A(S), .B(n678), .Z(n677) );
  XOR U1017 ( .A(B[696]), .B(B[695]), .Z(n678) );
  XOR U1018 ( .A(B[694]), .B(n679), .Z(O[695]) );
  AND U1019 ( .A(S), .B(n680), .Z(n679) );
  XOR U1020 ( .A(B[695]), .B(B[694]), .Z(n680) );
  XOR U1021 ( .A(B[693]), .B(n681), .Z(O[694]) );
  AND U1022 ( .A(S), .B(n682), .Z(n681) );
  XOR U1023 ( .A(B[694]), .B(B[693]), .Z(n682) );
  XOR U1024 ( .A(B[692]), .B(n683), .Z(O[693]) );
  AND U1025 ( .A(S), .B(n684), .Z(n683) );
  XOR U1026 ( .A(B[693]), .B(B[692]), .Z(n684) );
  XOR U1027 ( .A(B[691]), .B(n685), .Z(O[692]) );
  AND U1028 ( .A(S), .B(n686), .Z(n685) );
  XOR U1029 ( .A(B[692]), .B(B[691]), .Z(n686) );
  XOR U1030 ( .A(B[690]), .B(n687), .Z(O[691]) );
  AND U1031 ( .A(S), .B(n688), .Z(n687) );
  XOR U1032 ( .A(B[691]), .B(B[690]), .Z(n688) );
  XOR U1033 ( .A(B[689]), .B(n689), .Z(O[690]) );
  AND U1034 ( .A(S), .B(n690), .Z(n689) );
  XOR U1035 ( .A(B[690]), .B(B[689]), .Z(n690) );
  XOR U1036 ( .A(B[67]), .B(n691), .Z(O[68]) );
  AND U1037 ( .A(S), .B(n692), .Z(n691) );
  XOR U1038 ( .A(B[68]), .B(B[67]), .Z(n692) );
  XOR U1039 ( .A(B[688]), .B(n693), .Z(O[689]) );
  AND U1040 ( .A(S), .B(n694), .Z(n693) );
  XOR U1041 ( .A(B[689]), .B(B[688]), .Z(n694) );
  XOR U1042 ( .A(B[687]), .B(n695), .Z(O[688]) );
  AND U1043 ( .A(S), .B(n696), .Z(n695) );
  XOR U1044 ( .A(B[688]), .B(B[687]), .Z(n696) );
  XOR U1045 ( .A(B[686]), .B(n697), .Z(O[687]) );
  AND U1046 ( .A(S), .B(n698), .Z(n697) );
  XOR U1047 ( .A(B[687]), .B(B[686]), .Z(n698) );
  XOR U1048 ( .A(B[685]), .B(n699), .Z(O[686]) );
  AND U1049 ( .A(S), .B(n700), .Z(n699) );
  XOR U1050 ( .A(B[686]), .B(B[685]), .Z(n700) );
  XOR U1051 ( .A(B[684]), .B(n701), .Z(O[685]) );
  AND U1052 ( .A(S), .B(n702), .Z(n701) );
  XOR U1053 ( .A(B[685]), .B(B[684]), .Z(n702) );
  XOR U1054 ( .A(B[683]), .B(n703), .Z(O[684]) );
  AND U1055 ( .A(S), .B(n704), .Z(n703) );
  XOR U1056 ( .A(B[684]), .B(B[683]), .Z(n704) );
  XOR U1057 ( .A(B[682]), .B(n705), .Z(O[683]) );
  AND U1058 ( .A(S), .B(n706), .Z(n705) );
  XOR U1059 ( .A(B[683]), .B(B[682]), .Z(n706) );
  XOR U1060 ( .A(B[681]), .B(n707), .Z(O[682]) );
  AND U1061 ( .A(S), .B(n708), .Z(n707) );
  XOR U1062 ( .A(B[682]), .B(B[681]), .Z(n708) );
  XOR U1063 ( .A(B[680]), .B(n709), .Z(O[681]) );
  AND U1064 ( .A(S), .B(n710), .Z(n709) );
  XOR U1065 ( .A(B[681]), .B(B[680]), .Z(n710) );
  XOR U1066 ( .A(B[679]), .B(n711), .Z(O[680]) );
  AND U1067 ( .A(S), .B(n712), .Z(n711) );
  XOR U1068 ( .A(B[680]), .B(B[679]), .Z(n712) );
  XOR U1069 ( .A(B[66]), .B(n713), .Z(O[67]) );
  AND U1070 ( .A(S), .B(n714), .Z(n713) );
  XOR U1071 ( .A(B[67]), .B(B[66]), .Z(n714) );
  XOR U1072 ( .A(B[678]), .B(n715), .Z(O[679]) );
  AND U1073 ( .A(S), .B(n716), .Z(n715) );
  XOR U1074 ( .A(B[679]), .B(B[678]), .Z(n716) );
  XOR U1075 ( .A(B[677]), .B(n717), .Z(O[678]) );
  AND U1076 ( .A(S), .B(n718), .Z(n717) );
  XOR U1077 ( .A(B[678]), .B(B[677]), .Z(n718) );
  XOR U1078 ( .A(B[676]), .B(n719), .Z(O[677]) );
  AND U1079 ( .A(S), .B(n720), .Z(n719) );
  XOR U1080 ( .A(B[677]), .B(B[676]), .Z(n720) );
  XOR U1081 ( .A(B[675]), .B(n721), .Z(O[676]) );
  AND U1082 ( .A(S), .B(n722), .Z(n721) );
  XOR U1083 ( .A(B[676]), .B(B[675]), .Z(n722) );
  XOR U1084 ( .A(B[674]), .B(n723), .Z(O[675]) );
  AND U1085 ( .A(S), .B(n724), .Z(n723) );
  XOR U1086 ( .A(B[675]), .B(B[674]), .Z(n724) );
  XOR U1087 ( .A(B[673]), .B(n725), .Z(O[674]) );
  AND U1088 ( .A(S), .B(n726), .Z(n725) );
  XOR U1089 ( .A(B[674]), .B(B[673]), .Z(n726) );
  XOR U1090 ( .A(B[672]), .B(n727), .Z(O[673]) );
  AND U1091 ( .A(S), .B(n728), .Z(n727) );
  XOR U1092 ( .A(B[673]), .B(B[672]), .Z(n728) );
  XOR U1093 ( .A(B[671]), .B(n729), .Z(O[672]) );
  AND U1094 ( .A(S), .B(n730), .Z(n729) );
  XOR U1095 ( .A(B[672]), .B(B[671]), .Z(n730) );
  XOR U1096 ( .A(B[670]), .B(n731), .Z(O[671]) );
  AND U1097 ( .A(S), .B(n732), .Z(n731) );
  XOR U1098 ( .A(B[671]), .B(B[670]), .Z(n732) );
  XOR U1099 ( .A(B[669]), .B(n733), .Z(O[670]) );
  AND U1100 ( .A(S), .B(n734), .Z(n733) );
  XOR U1101 ( .A(B[670]), .B(B[669]), .Z(n734) );
  XOR U1102 ( .A(B[65]), .B(n735), .Z(O[66]) );
  AND U1103 ( .A(S), .B(n736), .Z(n735) );
  XOR U1104 ( .A(B[66]), .B(B[65]), .Z(n736) );
  XOR U1105 ( .A(B[668]), .B(n737), .Z(O[669]) );
  AND U1106 ( .A(S), .B(n738), .Z(n737) );
  XOR U1107 ( .A(B[669]), .B(B[668]), .Z(n738) );
  XOR U1108 ( .A(B[667]), .B(n739), .Z(O[668]) );
  AND U1109 ( .A(S), .B(n740), .Z(n739) );
  XOR U1110 ( .A(B[668]), .B(B[667]), .Z(n740) );
  XOR U1111 ( .A(B[666]), .B(n741), .Z(O[667]) );
  AND U1112 ( .A(S), .B(n742), .Z(n741) );
  XOR U1113 ( .A(B[667]), .B(B[666]), .Z(n742) );
  XOR U1114 ( .A(B[665]), .B(n743), .Z(O[666]) );
  AND U1115 ( .A(S), .B(n744), .Z(n743) );
  XOR U1116 ( .A(B[666]), .B(B[665]), .Z(n744) );
  XOR U1117 ( .A(B[664]), .B(n745), .Z(O[665]) );
  AND U1118 ( .A(S), .B(n746), .Z(n745) );
  XOR U1119 ( .A(B[665]), .B(B[664]), .Z(n746) );
  XOR U1120 ( .A(B[663]), .B(n747), .Z(O[664]) );
  AND U1121 ( .A(S), .B(n748), .Z(n747) );
  XOR U1122 ( .A(B[664]), .B(B[663]), .Z(n748) );
  XOR U1123 ( .A(B[662]), .B(n749), .Z(O[663]) );
  AND U1124 ( .A(S), .B(n750), .Z(n749) );
  XOR U1125 ( .A(B[663]), .B(B[662]), .Z(n750) );
  XOR U1126 ( .A(B[661]), .B(n751), .Z(O[662]) );
  AND U1127 ( .A(S), .B(n752), .Z(n751) );
  XOR U1128 ( .A(B[662]), .B(B[661]), .Z(n752) );
  XOR U1129 ( .A(B[660]), .B(n753), .Z(O[661]) );
  AND U1130 ( .A(S), .B(n754), .Z(n753) );
  XOR U1131 ( .A(B[661]), .B(B[660]), .Z(n754) );
  XOR U1132 ( .A(B[659]), .B(n755), .Z(O[660]) );
  AND U1133 ( .A(S), .B(n756), .Z(n755) );
  XOR U1134 ( .A(B[660]), .B(B[659]), .Z(n756) );
  XOR U1135 ( .A(B[64]), .B(n757), .Z(O[65]) );
  AND U1136 ( .A(S), .B(n758), .Z(n757) );
  XOR U1137 ( .A(B[65]), .B(B[64]), .Z(n758) );
  XOR U1138 ( .A(B[658]), .B(n759), .Z(O[659]) );
  AND U1139 ( .A(S), .B(n760), .Z(n759) );
  XOR U1140 ( .A(B[659]), .B(B[658]), .Z(n760) );
  XOR U1141 ( .A(B[657]), .B(n761), .Z(O[658]) );
  AND U1142 ( .A(S), .B(n762), .Z(n761) );
  XOR U1143 ( .A(B[658]), .B(B[657]), .Z(n762) );
  XOR U1144 ( .A(B[656]), .B(n763), .Z(O[657]) );
  AND U1145 ( .A(S), .B(n764), .Z(n763) );
  XOR U1146 ( .A(B[657]), .B(B[656]), .Z(n764) );
  XOR U1147 ( .A(B[655]), .B(n765), .Z(O[656]) );
  AND U1148 ( .A(S), .B(n766), .Z(n765) );
  XOR U1149 ( .A(B[656]), .B(B[655]), .Z(n766) );
  XOR U1150 ( .A(B[654]), .B(n767), .Z(O[655]) );
  AND U1151 ( .A(S), .B(n768), .Z(n767) );
  XOR U1152 ( .A(B[655]), .B(B[654]), .Z(n768) );
  XOR U1153 ( .A(B[653]), .B(n769), .Z(O[654]) );
  AND U1154 ( .A(S), .B(n770), .Z(n769) );
  XOR U1155 ( .A(B[654]), .B(B[653]), .Z(n770) );
  XOR U1156 ( .A(B[652]), .B(n771), .Z(O[653]) );
  AND U1157 ( .A(S), .B(n772), .Z(n771) );
  XOR U1158 ( .A(B[653]), .B(B[652]), .Z(n772) );
  XOR U1159 ( .A(B[651]), .B(n773), .Z(O[652]) );
  AND U1160 ( .A(S), .B(n774), .Z(n773) );
  XOR U1161 ( .A(B[652]), .B(B[651]), .Z(n774) );
  XOR U1162 ( .A(B[650]), .B(n775), .Z(O[651]) );
  AND U1163 ( .A(S), .B(n776), .Z(n775) );
  XOR U1164 ( .A(B[651]), .B(B[650]), .Z(n776) );
  XOR U1165 ( .A(B[649]), .B(n777), .Z(O[650]) );
  AND U1166 ( .A(S), .B(n778), .Z(n777) );
  XOR U1167 ( .A(B[650]), .B(B[649]), .Z(n778) );
  XOR U1168 ( .A(B[63]), .B(n779), .Z(O[64]) );
  AND U1169 ( .A(S), .B(n780), .Z(n779) );
  XOR U1170 ( .A(B[64]), .B(B[63]), .Z(n780) );
  XOR U1171 ( .A(B[648]), .B(n781), .Z(O[649]) );
  AND U1172 ( .A(S), .B(n782), .Z(n781) );
  XOR U1173 ( .A(B[649]), .B(B[648]), .Z(n782) );
  XOR U1174 ( .A(B[647]), .B(n783), .Z(O[648]) );
  AND U1175 ( .A(S), .B(n784), .Z(n783) );
  XOR U1176 ( .A(B[648]), .B(B[647]), .Z(n784) );
  XOR U1177 ( .A(B[646]), .B(n785), .Z(O[647]) );
  AND U1178 ( .A(S), .B(n786), .Z(n785) );
  XOR U1179 ( .A(B[647]), .B(B[646]), .Z(n786) );
  XOR U1180 ( .A(B[645]), .B(n787), .Z(O[646]) );
  AND U1181 ( .A(S), .B(n788), .Z(n787) );
  XOR U1182 ( .A(B[646]), .B(B[645]), .Z(n788) );
  XOR U1183 ( .A(B[644]), .B(n789), .Z(O[645]) );
  AND U1184 ( .A(S), .B(n790), .Z(n789) );
  XOR U1185 ( .A(B[645]), .B(B[644]), .Z(n790) );
  XOR U1186 ( .A(B[643]), .B(n791), .Z(O[644]) );
  AND U1187 ( .A(S), .B(n792), .Z(n791) );
  XOR U1188 ( .A(B[644]), .B(B[643]), .Z(n792) );
  XOR U1189 ( .A(B[642]), .B(n793), .Z(O[643]) );
  AND U1190 ( .A(S), .B(n794), .Z(n793) );
  XOR U1191 ( .A(B[643]), .B(B[642]), .Z(n794) );
  XOR U1192 ( .A(B[641]), .B(n795), .Z(O[642]) );
  AND U1193 ( .A(S), .B(n796), .Z(n795) );
  XOR U1194 ( .A(B[642]), .B(B[641]), .Z(n796) );
  XOR U1195 ( .A(B[640]), .B(n797), .Z(O[641]) );
  AND U1196 ( .A(S), .B(n798), .Z(n797) );
  XOR U1197 ( .A(B[641]), .B(B[640]), .Z(n798) );
  XOR U1198 ( .A(B[639]), .B(n799), .Z(O[640]) );
  AND U1199 ( .A(S), .B(n800), .Z(n799) );
  XOR U1200 ( .A(B[640]), .B(B[639]), .Z(n800) );
  XOR U1201 ( .A(B[62]), .B(n801), .Z(O[63]) );
  AND U1202 ( .A(S), .B(n802), .Z(n801) );
  XOR U1203 ( .A(B[63]), .B(B[62]), .Z(n802) );
  XOR U1204 ( .A(B[638]), .B(n803), .Z(O[639]) );
  AND U1205 ( .A(S), .B(n804), .Z(n803) );
  XOR U1206 ( .A(B[639]), .B(B[638]), .Z(n804) );
  XOR U1207 ( .A(B[637]), .B(n805), .Z(O[638]) );
  AND U1208 ( .A(S), .B(n806), .Z(n805) );
  XOR U1209 ( .A(B[638]), .B(B[637]), .Z(n806) );
  XOR U1210 ( .A(B[636]), .B(n807), .Z(O[637]) );
  AND U1211 ( .A(S), .B(n808), .Z(n807) );
  XOR U1212 ( .A(B[637]), .B(B[636]), .Z(n808) );
  XOR U1213 ( .A(B[635]), .B(n809), .Z(O[636]) );
  AND U1214 ( .A(S), .B(n810), .Z(n809) );
  XOR U1215 ( .A(B[636]), .B(B[635]), .Z(n810) );
  XOR U1216 ( .A(B[634]), .B(n811), .Z(O[635]) );
  AND U1217 ( .A(S), .B(n812), .Z(n811) );
  XOR U1218 ( .A(B[635]), .B(B[634]), .Z(n812) );
  XOR U1219 ( .A(B[633]), .B(n813), .Z(O[634]) );
  AND U1220 ( .A(S), .B(n814), .Z(n813) );
  XOR U1221 ( .A(B[634]), .B(B[633]), .Z(n814) );
  XOR U1222 ( .A(B[632]), .B(n815), .Z(O[633]) );
  AND U1223 ( .A(S), .B(n816), .Z(n815) );
  XOR U1224 ( .A(B[633]), .B(B[632]), .Z(n816) );
  XOR U1225 ( .A(B[631]), .B(n817), .Z(O[632]) );
  AND U1226 ( .A(S), .B(n818), .Z(n817) );
  XOR U1227 ( .A(B[632]), .B(B[631]), .Z(n818) );
  XOR U1228 ( .A(B[630]), .B(n819), .Z(O[631]) );
  AND U1229 ( .A(S), .B(n820), .Z(n819) );
  XOR U1230 ( .A(B[631]), .B(B[630]), .Z(n820) );
  XOR U1231 ( .A(B[629]), .B(n821), .Z(O[630]) );
  AND U1232 ( .A(S), .B(n822), .Z(n821) );
  XOR U1233 ( .A(B[630]), .B(B[629]), .Z(n822) );
  XOR U1234 ( .A(B[61]), .B(n823), .Z(O[62]) );
  AND U1235 ( .A(S), .B(n824), .Z(n823) );
  XOR U1236 ( .A(B[62]), .B(B[61]), .Z(n824) );
  XOR U1237 ( .A(B[628]), .B(n825), .Z(O[629]) );
  AND U1238 ( .A(S), .B(n826), .Z(n825) );
  XOR U1239 ( .A(B[629]), .B(B[628]), .Z(n826) );
  XOR U1240 ( .A(B[627]), .B(n827), .Z(O[628]) );
  AND U1241 ( .A(S), .B(n828), .Z(n827) );
  XOR U1242 ( .A(B[628]), .B(B[627]), .Z(n828) );
  XOR U1243 ( .A(B[626]), .B(n829), .Z(O[627]) );
  AND U1244 ( .A(S), .B(n830), .Z(n829) );
  XOR U1245 ( .A(B[627]), .B(B[626]), .Z(n830) );
  XOR U1246 ( .A(B[625]), .B(n831), .Z(O[626]) );
  AND U1247 ( .A(S), .B(n832), .Z(n831) );
  XOR U1248 ( .A(B[626]), .B(B[625]), .Z(n832) );
  XOR U1249 ( .A(B[624]), .B(n833), .Z(O[625]) );
  AND U1250 ( .A(S), .B(n834), .Z(n833) );
  XOR U1251 ( .A(B[625]), .B(B[624]), .Z(n834) );
  XOR U1252 ( .A(B[623]), .B(n835), .Z(O[624]) );
  AND U1253 ( .A(S), .B(n836), .Z(n835) );
  XOR U1254 ( .A(B[624]), .B(B[623]), .Z(n836) );
  XOR U1255 ( .A(B[622]), .B(n837), .Z(O[623]) );
  AND U1256 ( .A(S), .B(n838), .Z(n837) );
  XOR U1257 ( .A(B[623]), .B(B[622]), .Z(n838) );
  XOR U1258 ( .A(B[621]), .B(n839), .Z(O[622]) );
  AND U1259 ( .A(S), .B(n840), .Z(n839) );
  XOR U1260 ( .A(B[622]), .B(B[621]), .Z(n840) );
  XOR U1261 ( .A(B[620]), .B(n841), .Z(O[621]) );
  AND U1262 ( .A(S), .B(n842), .Z(n841) );
  XOR U1263 ( .A(B[621]), .B(B[620]), .Z(n842) );
  XOR U1264 ( .A(B[619]), .B(n843), .Z(O[620]) );
  AND U1265 ( .A(S), .B(n844), .Z(n843) );
  XOR U1266 ( .A(B[620]), .B(B[619]), .Z(n844) );
  XOR U1267 ( .A(B[60]), .B(n845), .Z(O[61]) );
  AND U1268 ( .A(S), .B(n846), .Z(n845) );
  XOR U1269 ( .A(B[61]), .B(B[60]), .Z(n846) );
  XOR U1270 ( .A(B[618]), .B(n847), .Z(O[619]) );
  AND U1271 ( .A(S), .B(n848), .Z(n847) );
  XOR U1272 ( .A(B[619]), .B(B[618]), .Z(n848) );
  XOR U1273 ( .A(B[617]), .B(n849), .Z(O[618]) );
  AND U1274 ( .A(S), .B(n850), .Z(n849) );
  XOR U1275 ( .A(B[618]), .B(B[617]), .Z(n850) );
  XOR U1276 ( .A(B[616]), .B(n851), .Z(O[617]) );
  AND U1277 ( .A(S), .B(n852), .Z(n851) );
  XOR U1278 ( .A(B[617]), .B(B[616]), .Z(n852) );
  XOR U1279 ( .A(B[615]), .B(n853), .Z(O[616]) );
  AND U1280 ( .A(S), .B(n854), .Z(n853) );
  XOR U1281 ( .A(B[616]), .B(B[615]), .Z(n854) );
  XOR U1282 ( .A(B[614]), .B(n855), .Z(O[615]) );
  AND U1283 ( .A(S), .B(n856), .Z(n855) );
  XOR U1284 ( .A(B[615]), .B(B[614]), .Z(n856) );
  XOR U1285 ( .A(B[613]), .B(n857), .Z(O[614]) );
  AND U1286 ( .A(S), .B(n858), .Z(n857) );
  XOR U1287 ( .A(B[614]), .B(B[613]), .Z(n858) );
  XOR U1288 ( .A(B[612]), .B(n859), .Z(O[613]) );
  AND U1289 ( .A(S), .B(n860), .Z(n859) );
  XOR U1290 ( .A(B[613]), .B(B[612]), .Z(n860) );
  XOR U1291 ( .A(B[611]), .B(n861), .Z(O[612]) );
  AND U1292 ( .A(S), .B(n862), .Z(n861) );
  XOR U1293 ( .A(B[612]), .B(B[611]), .Z(n862) );
  XOR U1294 ( .A(B[610]), .B(n863), .Z(O[611]) );
  AND U1295 ( .A(S), .B(n864), .Z(n863) );
  XOR U1296 ( .A(B[611]), .B(B[610]), .Z(n864) );
  XOR U1297 ( .A(B[609]), .B(n865), .Z(O[610]) );
  AND U1298 ( .A(S), .B(n866), .Z(n865) );
  XOR U1299 ( .A(B[610]), .B(B[609]), .Z(n866) );
  XOR U1300 ( .A(B[59]), .B(n867), .Z(O[60]) );
  AND U1301 ( .A(S), .B(n868), .Z(n867) );
  XOR U1302 ( .A(B[60]), .B(B[59]), .Z(n868) );
  XOR U1303 ( .A(B[608]), .B(n869), .Z(O[609]) );
  AND U1304 ( .A(S), .B(n870), .Z(n869) );
  XOR U1305 ( .A(B[609]), .B(B[608]), .Z(n870) );
  XOR U1306 ( .A(B[607]), .B(n871), .Z(O[608]) );
  AND U1307 ( .A(S), .B(n872), .Z(n871) );
  XOR U1308 ( .A(B[608]), .B(B[607]), .Z(n872) );
  XOR U1309 ( .A(B[606]), .B(n873), .Z(O[607]) );
  AND U1310 ( .A(S), .B(n874), .Z(n873) );
  XOR U1311 ( .A(B[607]), .B(B[606]), .Z(n874) );
  XOR U1312 ( .A(B[605]), .B(n875), .Z(O[606]) );
  AND U1313 ( .A(S), .B(n876), .Z(n875) );
  XOR U1314 ( .A(B[606]), .B(B[605]), .Z(n876) );
  XOR U1315 ( .A(B[604]), .B(n877), .Z(O[605]) );
  AND U1316 ( .A(S), .B(n878), .Z(n877) );
  XOR U1317 ( .A(B[605]), .B(B[604]), .Z(n878) );
  XOR U1318 ( .A(B[603]), .B(n879), .Z(O[604]) );
  AND U1319 ( .A(S), .B(n880), .Z(n879) );
  XOR U1320 ( .A(B[604]), .B(B[603]), .Z(n880) );
  XOR U1321 ( .A(B[602]), .B(n881), .Z(O[603]) );
  AND U1322 ( .A(S), .B(n882), .Z(n881) );
  XOR U1323 ( .A(B[603]), .B(B[602]), .Z(n882) );
  XOR U1324 ( .A(B[601]), .B(n883), .Z(O[602]) );
  AND U1325 ( .A(S), .B(n884), .Z(n883) );
  XOR U1326 ( .A(B[602]), .B(B[601]), .Z(n884) );
  XOR U1327 ( .A(B[600]), .B(n885), .Z(O[601]) );
  AND U1328 ( .A(S), .B(n886), .Z(n885) );
  XOR U1329 ( .A(B[601]), .B(B[600]), .Z(n886) );
  XOR U1330 ( .A(B[599]), .B(n887), .Z(O[600]) );
  AND U1331 ( .A(S), .B(n888), .Z(n887) );
  XOR U1332 ( .A(B[600]), .B(B[599]), .Z(n888) );
  XOR U1333 ( .A(B[4]), .B(n889), .Z(O[5]) );
  AND U1334 ( .A(S), .B(n890), .Z(n889) );
  XOR U1335 ( .A(B[5]), .B(B[4]), .Z(n890) );
  XOR U1336 ( .A(B[58]), .B(n891), .Z(O[59]) );
  AND U1337 ( .A(S), .B(n892), .Z(n891) );
  XOR U1338 ( .A(B[59]), .B(B[58]), .Z(n892) );
  XOR U1339 ( .A(B[598]), .B(n893), .Z(O[599]) );
  AND U1340 ( .A(S), .B(n894), .Z(n893) );
  XOR U1341 ( .A(B[599]), .B(B[598]), .Z(n894) );
  XOR U1342 ( .A(B[597]), .B(n895), .Z(O[598]) );
  AND U1343 ( .A(S), .B(n896), .Z(n895) );
  XOR U1344 ( .A(B[598]), .B(B[597]), .Z(n896) );
  XOR U1345 ( .A(B[596]), .B(n897), .Z(O[597]) );
  AND U1346 ( .A(S), .B(n898), .Z(n897) );
  XOR U1347 ( .A(B[597]), .B(B[596]), .Z(n898) );
  XOR U1348 ( .A(B[595]), .B(n899), .Z(O[596]) );
  AND U1349 ( .A(S), .B(n900), .Z(n899) );
  XOR U1350 ( .A(B[596]), .B(B[595]), .Z(n900) );
  XOR U1351 ( .A(B[594]), .B(n901), .Z(O[595]) );
  AND U1352 ( .A(S), .B(n902), .Z(n901) );
  XOR U1353 ( .A(B[595]), .B(B[594]), .Z(n902) );
  XOR U1354 ( .A(B[593]), .B(n903), .Z(O[594]) );
  AND U1355 ( .A(S), .B(n904), .Z(n903) );
  XOR U1356 ( .A(B[594]), .B(B[593]), .Z(n904) );
  XOR U1357 ( .A(B[592]), .B(n905), .Z(O[593]) );
  AND U1358 ( .A(S), .B(n906), .Z(n905) );
  XOR U1359 ( .A(B[593]), .B(B[592]), .Z(n906) );
  XOR U1360 ( .A(B[591]), .B(n907), .Z(O[592]) );
  AND U1361 ( .A(S), .B(n908), .Z(n907) );
  XOR U1362 ( .A(B[592]), .B(B[591]), .Z(n908) );
  XOR U1363 ( .A(B[590]), .B(n909), .Z(O[591]) );
  AND U1364 ( .A(S), .B(n910), .Z(n909) );
  XOR U1365 ( .A(B[591]), .B(B[590]), .Z(n910) );
  XOR U1366 ( .A(B[589]), .B(n911), .Z(O[590]) );
  AND U1367 ( .A(S), .B(n912), .Z(n911) );
  XOR U1368 ( .A(B[590]), .B(B[589]), .Z(n912) );
  XOR U1369 ( .A(B[57]), .B(n913), .Z(O[58]) );
  AND U1370 ( .A(S), .B(n914), .Z(n913) );
  XOR U1371 ( .A(B[58]), .B(B[57]), .Z(n914) );
  XOR U1372 ( .A(B[588]), .B(n915), .Z(O[589]) );
  AND U1373 ( .A(S), .B(n916), .Z(n915) );
  XOR U1374 ( .A(B[589]), .B(B[588]), .Z(n916) );
  XOR U1375 ( .A(B[587]), .B(n917), .Z(O[588]) );
  AND U1376 ( .A(S), .B(n918), .Z(n917) );
  XOR U1377 ( .A(B[588]), .B(B[587]), .Z(n918) );
  XOR U1378 ( .A(B[586]), .B(n919), .Z(O[587]) );
  AND U1379 ( .A(S), .B(n920), .Z(n919) );
  XOR U1380 ( .A(B[587]), .B(B[586]), .Z(n920) );
  XOR U1381 ( .A(B[585]), .B(n921), .Z(O[586]) );
  AND U1382 ( .A(S), .B(n922), .Z(n921) );
  XOR U1383 ( .A(B[586]), .B(B[585]), .Z(n922) );
  XOR U1384 ( .A(B[584]), .B(n923), .Z(O[585]) );
  AND U1385 ( .A(S), .B(n924), .Z(n923) );
  XOR U1386 ( .A(B[585]), .B(B[584]), .Z(n924) );
  XOR U1387 ( .A(B[583]), .B(n925), .Z(O[584]) );
  AND U1388 ( .A(S), .B(n926), .Z(n925) );
  XOR U1389 ( .A(B[584]), .B(B[583]), .Z(n926) );
  XOR U1390 ( .A(B[582]), .B(n927), .Z(O[583]) );
  AND U1391 ( .A(S), .B(n928), .Z(n927) );
  XOR U1392 ( .A(B[583]), .B(B[582]), .Z(n928) );
  XOR U1393 ( .A(B[581]), .B(n929), .Z(O[582]) );
  AND U1394 ( .A(S), .B(n930), .Z(n929) );
  XOR U1395 ( .A(B[582]), .B(B[581]), .Z(n930) );
  XOR U1396 ( .A(B[580]), .B(n931), .Z(O[581]) );
  AND U1397 ( .A(S), .B(n932), .Z(n931) );
  XOR U1398 ( .A(B[581]), .B(B[580]), .Z(n932) );
  XOR U1399 ( .A(B[579]), .B(n933), .Z(O[580]) );
  AND U1400 ( .A(S), .B(n934), .Z(n933) );
  XOR U1401 ( .A(B[580]), .B(B[579]), .Z(n934) );
  XOR U1402 ( .A(B[56]), .B(n935), .Z(O[57]) );
  AND U1403 ( .A(S), .B(n936), .Z(n935) );
  XOR U1404 ( .A(B[57]), .B(B[56]), .Z(n936) );
  XOR U1405 ( .A(B[578]), .B(n937), .Z(O[579]) );
  AND U1406 ( .A(S), .B(n938), .Z(n937) );
  XOR U1407 ( .A(B[579]), .B(B[578]), .Z(n938) );
  XOR U1408 ( .A(B[577]), .B(n939), .Z(O[578]) );
  AND U1409 ( .A(S), .B(n940), .Z(n939) );
  XOR U1410 ( .A(B[578]), .B(B[577]), .Z(n940) );
  XOR U1411 ( .A(B[576]), .B(n941), .Z(O[577]) );
  AND U1412 ( .A(S), .B(n942), .Z(n941) );
  XOR U1413 ( .A(B[577]), .B(B[576]), .Z(n942) );
  XOR U1414 ( .A(B[575]), .B(n943), .Z(O[576]) );
  AND U1415 ( .A(S), .B(n944), .Z(n943) );
  XOR U1416 ( .A(B[576]), .B(B[575]), .Z(n944) );
  XOR U1417 ( .A(B[574]), .B(n945), .Z(O[575]) );
  AND U1418 ( .A(S), .B(n946), .Z(n945) );
  XOR U1419 ( .A(B[575]), .B(B[574]), .Z(n946) );
  XOR U1420 ( .A(B[573]), .B(n947), .Z(O[574]) );
  AND U1421 ( .A(S), .B(n948), .Z(n947) );
  XOR U1422 ( .A(B[574]), .B(B[573]), .Z(n948) );
  XOR U1423 ( .A(B[572]), .B(n949), .Z(O[573]) );
  AND U1424 ( .A(S), .B(n950), .Z(n949) );
  XOR U1425 ( .A(B[573]), .B(B[572]), .Z(n950) );
  XOR U1426 ( .A(B[571]), .B(n951), .Z(O[572]) );
  AND U1427 ( .A(S), .B(n952), .Z(n951) );
  XOR U1428 ( .A(B[572]), .B(B[571]), .Z(n952) );
  XOR U1429 ( .A(B[570]), .B(n953), .Z(O[571]) );
  AND U1430 ( .A(S), .B(n954), .Z(n953) );
  XOR U1431 ( .A(B[571]), .B(B[570]), .Z(n954) );
  XOR U1432 ( .A(B[569]), .B(n955), .Z(O[570]) );
  AND U1433 ( .A(S), .B(n956), .Z(n955) );
  XOR U1434 ( .A(B[570]), .B(B[569]), .Z(n956) );
  XOR U1435 ( .A(B[55]), .B(n957), .Z(O[56]) );
  AND U1436 ( .A(S), .B(n958), .Z(n957) );
  XOR U1437 ( .A(B[56]), .B(B[55]), .Z(n958) );
  XOR U1438 ( .A(B[568]), .B(n959), .Z(O[569]) );
  AND U1439 ( .A(S), .B(n960), .Z(n959) );
  XOR U1440 ( .A(B[569]), .B(B[568]), .Z(n960) );
  XOR U1441 ( .A(B[567]), .B(n961), .Z(O[568]) );
  AND U1442 ( .A(S), .B(n962), .Z(n961) );
  XOR U1443 ( .A(B[568]), .B(B[567]), .Z(n962) );
  XOR U1444 ( .A(B[566]), .B(n963), .Z(O[567]) );
  AND U1445 ( .A(S), .B(n964), .Z(n963) );
  XOR U1446 ( .A(B[567]), .B(B[566]), .Z(n964) );
  XOR U1447 ( .A(B[565]), .B(n965), .Z(O[566]) );
  AND U1448 ( .A(S), .B(n966), .Z(n965) );
  XOR U1449 ( .A(B[566]), .B(B[565]), .Z(n966) );
  XOR U1450 ( .A(B[564]), .B(n967), .Z(O[565]) );
  AND U1451 ( .A(S), .B(n968), .Z(n967) );
  XOR U1452 ( .A(B[565]), .B(B[564]), .Z(n968) );
  XOR U1453 ( .A(B[563]), .B(n969), .Z(O[564]) );
  AND U1454 ( .A(S), .B(n970), .Z(n969) );
  XOR U1455 ( .A(B[564]), .B(B[563]), .Z(n970) );
  XOR U1456 ( .A(B[562]), .B(n971), .Z(O[563]) );
  AND U1457 ( .A(S), .B(n972), .Z(n971) );
  XOR U1458 ( .A(B[563]), .B(B[562]), .Z(n972) );
  XOR U1459 ( .A(B[561]), .B(n973), .Z(O[562]) );
  AND U1460 ( .A(S), .B(n974), .Z(n973) );
  XOR U1461 ( .A(B[562]), .B(B[561]), .Z(n974) );
  XOR U1462 ( .A(B[560]), .B(n975), .Z(O[561]) );
  AND U1463 ( .A(S), .B(n976), .Z(n975) );
  XOR U1464 ( .A(B[561]), .B(B[560]), .Z(n976) );
  XOR U1465 ( .A(B[559]), .B(n977), .Z(O[560]) );
  AND U1466 ( .A(S), .B(n978), .Z(n977) );
  XOR U1467 ( .A(B[560]), .B(B[559]), .Z(n978) );
  XOR U1468 ( .A(B[54]), .B(n979), .Z(O[55]) );
  AND U1469 ( .A(S), .B(n980), .Z(n979) );
  XOR U1470 ( .A(B[55]), .B(B[54]), .Z(n980) );
  XOR U1471 ( .A(B[558]), .B(n981), .Z(O[559]) );
  AND U1472 ( .A(S), .B(n982), .Z(n981) );
  XOR U1473 ( .A(B[559]), .B(B[558]), .Z(n982) );
  XOR U1474 ( .A(B[557]), .B(n983), .Z(O[558]) );
  AND U1475 ( .A(S), .B(n984), .Z(n983) );
  XOR U1476 ( .A(B[558]), .B(B[557]), .Z(n984) );
  XOR U1477 ( .A(B[556]), .B(n985), .Z(O[557]) );
  AND U1478 ( .A(S), .B(n986), .Z(n985) );
  XOR U1479 ( .A(B[557]), .B(B[556]), .Z(n986) );
  XOR U1480 ( .A(B[555]), .B(n987), .Z(O[556]) );
  AND U1481 ( .A(S), .B(n988), .Z(n987) );
  XOR U1482 ( .A(B[556]), .B(B[555]), .Z(n988) );
  XOR U1483 ( .A(B[554]), .B(n989), .Z(O[555]) );
  AND U1484 ( .A(S), .B(n990), .Z(n989) );
  XOR U1485 ( .A(B[555]), .B(B[554]), .Z(n990) );
  XOR U1486 ( .A(B[553]), .B(n991), .Z(O[554]) );
  AND U1487 ( .A(S), .B(n992), .Z(n991) );
  XOR U1488 ( .A(B[554]), .B(B[553]), .Z(n992) );
  XOR U1489 ( .A(B[552]), .B(n993), .Z(O[553]) );
  AND U1490 ( .A(S), .B(n994), .Z(n993) );
  XOR U1491 ( .A(B[553]), .B(B[552]), .Z(n994) );
  XOR U1492 ( .A(B[551]), .B(n995), .Z(O[552]) );
  AND U1493 ( .A(S), .B(n996), .Z(n995) );
  XOR U1494 ( .A(B[552]), .B(B[551]), .Z(n996) );
  XOR U1495 ( .A(B[550]), .B(n997), .Z(O[551]) );
  AND U1496 ( .A(S), .B(n998), .Z(n997) );
  XOR U1497 ( .A(B[551]), .B(B[550]), .Z(n998) );
  XOR U1498 ( .A(B[549]), .B(n999), .Z(O[550]) );
  AND U1499 ( .A(S), .B(n1000), .Z(n999) );
  XOR U1500 ( .A(B[550]), .B(B[549]), .Z(n1000) );
  XOR U1501 ( .A(B[53]), .B(n1001), .Z(O[54]) );
  AND U1502 ( .A(S), .B(n1002), .Z(n1001) );
  XOR U1503 ( .A(B[54]), .B(B[53]), .Z(n1002) );
  XOR U1504 ( .A(B[548]), .B(n1003), .Z(O[549]) );
  AND U1505 ( .A(S), .B(n1004), .Z(n1003) );
  XOR U1506 ( .A(B[549]), .B(B[548]), .Z(n1004) );
  XOR U1507 ( .A(B[547]), .B(n1005), .Z(O[548]) );
  AND U1508 ( .A(S), .B(n1006), .Z(n1005) );
  XOR U1509 ( .A(B[548]), .B(B[547]), .Z(n1006) );
  XOR U1510 ( .A(B[546]), .B(n1007), .Z(O[547]) );
  AND U1511 ( .A(S), .B(n1008), .Z(n1007) );
  XOR U1512 ( .A(B[547]), .B(B[546]), .Z(n1008) );
  XOR U1513 ( .A(B[545]), .B(n1009), .Z(O[546]) );
  AND U1514 ( .A(S), .B(n1010), .Z(n1009) );
  XOR U1515 ( .A(B[546]), .B(B[545]), .Z(n1010) );
  XOR U1516 ( .A(B[544]), .B(n1011), .Z(O[545]) );
  AND U1517 ( .A(S), .B(n1012), .Z(n1011) );
  XOR U1518 ( .A(B[545]), .B(B[544]), .Z(n1012) );
  XOR U1519 ( .A(B[543]), .B(n1013), .Z(O[544]) );
  AND U1520 ( .A(S), .B(n1014), .Z(n1013) );
  XOR U1521 ( .A(B[544]), .B(B[543]), .Z(n1014) );
  XOR U1522 ( .A(B[542]), .B(n1015), .Z(O[543]) );
  AND U1523 ( .A(S), .B(n1016), .Z(n1015) );
  XOR U1524 ( .A(B[543]), .B(B[542]), .Z(n1016) );
  XOR U1525 ( .A(B[541]), .B(n1017), .Z(O[542]) );
  AND U1526 ( .A(S), .B(n1018), .Z(n1017) );
  XOR U1527 ( .A(B[542]), .B(B[541]), .Z(n1018) );
  XOR U1528 ( .A(B[540]), .B(n1019), .Z(O[541]) );
  AND U1529 ( .A(S), .B(n1020), .Z(n1019) );
  XOR U1530 ( .A(B[541]), .B(B[540]), .Z(n1020) );
  XOR U1531 ( .A(B[539]), .B(n1021), .Z(O[540]) );
  AND U1532 ( .A(S), .B(n1022), .Z(n1021) );
  XOR U1533 ( .A(B[540]), .B(B[539]), .Z(n1022) );
  XOR U1534 ( .A(B[52]), .B(n1023), .Z(O[53]) );
  AND U1535 ( .A(S), .B(n1024), .Z(n1023) );
  XOR U1536 ( .A(B[53]), .B(B[52]), .Z(n1024) );
  XOR U1537 ( .A(B[538]), .B(n1025), .Z(O[539]) );
  AND U1538 ( .A(S), .B(n1026), .Z(n1025) );
  XOR U1539 ( .A(B[539]), .B(B[538]), .Z(n1026) );
  XOR U1540 ( .A(B[537]), .B(n1027), .Z(O[538]) );
  AND U1541 ( .A(S), .B(n1028), .Z(n1027) );
  XOR U1542 ( .A(B[538]), .B(B[537]), .Z(n1028) );
  XOR U1543 ( .A(B[536]), .B(n1029), .Z(O[537]) );
  AND U1544 ( .A(S), .B(n1030), .Z(n1029) );
  XOR U1545 ( .A(B[537]), .B(B[536]), .Z(n1030) );
  XOR U1546 ( .A(B[535]), .B(n1031), .Z(O[536]) );
  AND U1547 ( .A(S), .B(n1032), .Z(n1031) );
  XOR U1548 ( .A(B[536]), .B(B[535]), .Z(n1032) );
  XOR U1549 ( .A(B[534]), .B(n1033), .Z(O[535]) );
  AND U1550 ( .A(S), .B(n1034), .Z(n1033) );
  XOR U1551 ( .A(B[535]), .B(B[534]), .Z(n1034) );
  XOR U1552 ( .A(B[533]), .B(n1035), .Z(O[534]) );
  AND U1553 ( .A(S), .B(n1036), .Z(n1035) );
  XOR U1554 ( .A(B[534]), .B(B[533]), .Z(n1036) );
  XOR U1555 ( .A(B[532]), .B(n1037), .Z(O[533]) );
  AND U1556 ( .A(S), .B(n1038), .Z(n1037) );
  XOR U1557 ( .A(B[533]), .B(B[532]), .Z(n1038) );
  XOR U1558 ( .A(B[531]), .B(n1039), .Z(O[532]) );
  AND U1559 ( .A(S), .B(n1040), .Z(n1039) );
  XOR U1560 ( .A(B[532]), .B(B[531]), .Z(n1040) );
  XOR U1561 ( .A(B[530]), .B(n1041), .Z(O[531]) );
  AND U1562 ( .A(S), .B(n1042), .Z(n1041) );
  XOR U1563 ( .A(B[531]), .B(B[530]), .Z(n1042) );
  XOR U1564 ( .A(B[529]), .B(n1043), .Z(O[530]) );
  AND U1565 ( .A(S), .B(n1044), .Z(n1043) );
  XOR U1566 ( .A(B[530]), .B(B[529]), .Z(n1044) );
  XOR U1567 ( .A(B[51]), .B(n1045), .Z(O[52]) );
  AND U1568 ( .A(S), .B(n1046), .Z(n1045) );
  XOR U1569 ( .A(B[52]), .B(B[51]), .Z(n1046) );
  XOR U1570 ( .A(B[528]), .B(n1047), .Z(O[529]) );
  AND U1571 ( .A(S), .B(n1048), .Z(n1047) );
  XOR U1572 ( .A(B[529]), .B(B[528]), .Z(n1048) );
  XOR U1573 ( .A(B[527]), .B(n1049), .Z(O[528]) );
  AND U1574 ( .A(S), .B(n1050), .Z(n1049) );
  XOR U1575 ( .A(B[528]), .B(B[527]), .Z(n1050) );
  XOR U1576 ( .A(B[526]), .B(n1051), .Z(O[527]) );
  AND U1577 ( .A(S), .B(n1052), .Z(n1051) );
  XOR U1578 ( .A(B[527]), .B(B[526]), .Z(n1052) );
  XOR U1579 ( .A(B[525]), .B(n1053), .Z(O[526]) );
  AND U1580 ( .A(S), .B(n1054), .Z(n1053) );
  XOR U1581 ( .A(B[526]), .B(B[525]), .Z(n1054) );
  XOR U1582 ( .A(B[524]), .B(n1055), .Z(O[525]) );
  AND U1583 ( .A(S), .B(n1056), .Z(n1055) );
  XOR U1584 ( .A(B[525]), .B(B[524]), .Z(n1056) );
  XOR U1585 ( .A(B[523]), .B(n1057), .Z(O[524]) );
  AND U1586 ( .A(S), .B(n1058), .Z(n1057) );
  XOR U1587 ( .A(B[524]), .B(B[523]), .Z(n1058) );
  XOR U1588 ( .A(B[522]), .B(n1059), .Z(O[523]) );
  AND U1589 ( .A(S), .B(n1060), .Z(n1059) );
  XOR U1590 ( .A(B[523]), .B(B[522]), .Z(n1060) );
  XOR U1591 ( .A(B[521]), .B(n1061), .Z(O[522]) );
  AND U1592 ( .A(S), .B(n1062), .Z(n1061) );
  XOR U1593 ( .A(B[522]), .B(B[521]), .Z(n1062) );
  XOR U1594 ( .A(B[520]), .B(n1063), .Z(O[521]) );
  AND U1595 ( .A(S), .B(n1064), .Z(n1063) );
  XOR U1596 ( .A(B[521]), .B(B[520]), .Z(n1064) );
  XOR U1597 ( .A(B[519]), .B(n1065), .Z(O[520]) );
  AND U1598 ( .A(S), .B(n1066), .Z(n1065) );
  XOR U1599 ( .A(B[520]), .B(B[519]), .Z(n1066) );
  XOR U1600 ( .A(B[50]), .B(n1067), .Z(O[51]) );
  AND U1601 ( .A(S), .B(n1068), .Z(n1067) );
  XOR U1602 ( .A(B[51]), .B(B[50]), .Z(n1068) );
  XOR U1603 ( .A(B[518]), .B(n1069), .Z(O[519]) );
  AND U1604 ( .A(S), .B(n1070), .Z(n1069) );
  XOR U1605 ( .A(B[519]), .B(B[518]), .Z(n1070) );
  XOR U1606 ( .A(B[517]), .B(n1071), .Z(O[518]) );
  AND U1607 ( .A(S), .B(n1072), .Z(n1071) );
  XOR U1608 ( .A(B[518]), .B(B[517]), .Z(n1072) );
  XOR U1609 ( .A(B[516]), .B(n1073), .Z(O[517]) );
  AND U1610 ( .A(S), .B(n1074), .Z(n1073) );
  XOR U1611 ( .A(B[517]), .B(B[516]), .Z(n1074) );
  XOR U1612 ( .A(B[515]), .B(n1075), .Z(O[516]) );
  AND U1613 ( .A(S), .B(n1076), .Z(n1075) );
  XOR U1614 ( .A(B[516]), .B(B[515]), .Z(n1076) );
  XOR U1615 ( .A(B[514]), .B(n1077), .Z(O[515]) );
  AND U1616 ( .A(S), .B(n1078), .Z(n1077) );
  XOR U1617 ( .A(B[515]), .B(B[514]), .Z(n1078) );
  XOR U1618 ( .A(B[513]), .B(n1079), .Z(O[514]) );
  AND U1619 ( .A(S), .B(n1080), .Z(n1079) );
  XOR U1620 ( .A(B[514]), .B(B[513]), .Z(n1080) );
  XOR U1621 ( .A(B[512]), .B(n1081), .Z(O[513]) );
  AND U1622 ( .A(S), .B(n1082), .Z(n1081) );
  XOR U1623 ( .A(B[513]), .B(B[512]), .Z(n1082) );
  XOR U1624 ( .A(B[511]), .B(n1083), .Z(O[512]) );
  AND U1625 ( .A(S), .B(n1084), .Z(n1083) );
  XOR U1626 ( .A(B[512]), .B(B[511]), .Z(n1084) );
  XOR U1627 ( .A(B[510]), .B(n1085), .Z(O[511]) );
  AND U1628 ( .A(S), .B(n1086), .Z(n1085) );
  XOR U1629 ( .A(B[511]), .B(B[510]), .Z(n1086) );
  XOR U1630 ( .A(B[509]), .B(n1087), .Z(O[510]) );
  AND U1631 ( .A(S), .B(n1088), .Z(n1087) );
  XOR U1632 ( .A(B[510]), .B(B[509]), .Z(n1088) );
  XOR U1633 ( .A(B[49]), .B(n1089), .Z(O[50]) );
  AND U1634 ( .A(S), .B(n1090), .Z(n1089) );
  XOR U1635 ( .A(B[50]), .B(B[49]), .Z(n1090) );
  XOR U1636 ( .A(B[508]), .B(n1091), .Z(O[509]) );
  AND U1637 ( .A(S), .B(n1092), .Z(n1091) );
  XOR U1638 ( .A(B[509]), .B(B[508]), .Z(n1092) );
  XOR U1639 ( .A(B[507]), .B(n1093), .Z(O[508]) );
  AND U1640 ( .A(S), .B(n1094), .Z(n1093) );
  XOR U1641 ( .A(B[508]), .B(B[507]), .Z(n1094) );
  XOR U1642 ( .A(B[506]), .B(n1095), .Z(O[507]) );
  AND U1643 ( .A(S), .B(n1096), .Z(n1095) );
  XOR U1644 ( .A(B[507]), .B(B[506]), .Z(n1096) );
  XOR U1645 ( .A(B[505]), .B(n1097), .Z(O[506]) );
  AND U1646 ( .A(S), .B(n1098), .Z(n1097) );
  XOR U1647 ( .A(B[506]), .B(B[505]), .Z(n1098) );
  XOR U1648 ( .A(B[504]), .B(n1099), .Z(O[505]) );
  AND U1649 ( .A(S), .B(n1100), .Z(n1099) );
  XOR U1650 ( .A(B[505]), .B(B[504]), .Z(n1100) );
  XOR U1651 ( .A(B[503]), .B(n1101), .Z(O[504]) );
  AND U1652 ( .A(S), .B(n1102), .Z(n1101) );
  XOR U1653 ( .A(B[504]), .B(B[503]), .Z(n1102) );
  XOR U1654 ( .A(B[502]), .B(n1103), .Z(O[503]) );
  AND U1655 ( .A(S), .B(n1104), .Z(n1103) );
  XOR U1656 ( .A(B[503]), .B(B[502]), .Z(n1104) );
  XOR U1657 ( .A(B[501]), .B(n1105), .Z(O[502]) );
  AND U1658 ( .A(S), .B(n1106), .Z(n1105) );
  XOR U1659 ( .A(B[502]), .B(B[501]), .Z(n1106) );
  XOR U1660 ( .A(B[500]), .B(n1107), .Z(O[501]) );
  AND U1661 ( .A(S), .B(n1108), .Z(n1107) );
  XOR U1662 ( .A(B[501]), .B(B[500]), .Z(n1108) );
  XOR U1663 ( .A(B[499]), .B(n1109), .Z(O[500]) );
  AND U1664 ( .A(S), .B(n1110), .Z(n1109) );
  XOR U1665 ( .A(B[500]), .B(B[499]), .Z(n1110) );
  XOR U1666 ( .A(B[3]), .B(n1111), .Z(O[4]) );
  AND U1667 ( .A(S), .B(n1112), .Z(n1111) );
  XOR U1668 ( .A(B[4]), .B(B[3]), .Z(n1112) );
  XOR U1669 ( .A(B[48]), .B(n1113), .Z(O[49]) );
  AND U1670 ( .A(S), .B(n1114), .Z(n1113) );
  XOR U1671 ( .A(B[49]), .B(B[48]), .Z(n1114) );
  XOR U1672 ( .A(B[498]), .B(n1115), .Z(O[499]) );
  AND U1673 ( .A(S), .B(n1116), .Z(n1115) );
  XOR U1674 ( .A(B[499]), .B(B[498]), .Z(n1116) );
  XOR U1675 ( .A(B[497]), .B(n1117), .Z(O[498]) );
  AND U1676 ( .A(S), .B(n1118), .Z(n1117) );
  XOR U1677 ( .A(B[498]), .B(B[497]), .Z(n1118) );
  XOR U1678 ( .A(B[496]), .B(n1119), .Z(O[497]) );
  AND U1679 ( .A(S), .B(n1120), .Z(n1119) );
  XOR U1680 ( .A(B[497]), .B(B[496]), .Z(n1120) );
  XOR U1681 ( .A(B[495]), .B(n1121), .Z(O[496]) );
  AND U1682 ( .A(S), .B(n1122), .Z(n1121) );
  XOR U1683 ( .A(B[496]), .B(B[495]), .Z(n1122) );
  XOR U1684 ( .A(B[494]), .B(n1123), .Z(O[495]) );
  AND U1685 ( .A(S), .B(n1124), .Z(n1123) );
  XOR U1686 ( .A(B[495]), .B(B[494]), .Z(n1124) );
  XOR U1687 ( .A(B[493]), .B(n1125), .Z(O[494]) );
  AND U1688 ( .A(S), .B(n1126), .Z(n1125) );
  XOR U1689 ( .A(B[494]), .B(B[493]), .Z(n1126) );
  XOR U1690 ( .A(B[492]), .B(n1127), .Z(O[493]) );
  AND U1691 ( .A(S), .B(n1128), .Z(n1127) );
  XOR U1692 ( .A(B[493]), .B(B[492]), .Z(n1128) );
  XOR U1693 ( .A(B[491]), .B(n1129), .Z(O[492]) );
  AND U1694 ( .A(S), .B(n1130), .Z(n1129) );
  XOR U1695 ( .A(B[492]), .B(B[491]), .Z(n1130) );
  XOR U1696 ( .A(B[490]), .B(n1131), .Z(O[491]) );
  AND U1697 ( .A(S), .B(n1132), .Z(n1131) );
  XOR U1698 ( .A(B[491]), .B(B[490]), .Z(n1132) );
  XOR U1699 ( .A(B[489]), .B(n1133), .Z(O[490]) );
  AND U1700 ( .A(S), .B(n1134), .Z(n1133) );
  XOR U1701 ( .A(B[490]), .B(B[489]), .Z(n1134) );
  XOR U1702 ( .A(B[47]), .B(n1135), .Z(O[48]) );
  AND U1703 ( .A(S), .B(n1136), .Z(n1135) );
  XOR U1704 ( .A(B[48]), .B(B[47]), .Z(n1136) );
  XOR U1705 ( .A(B[488]), .B(n1137), .Z(O[489]) );
  AND U1706 ( .A(S), .B(n1138), .Z(n1137) );
  XOR U1707 ( .A(B[489]), .B(B[488]), .Z(n1138) );
  XOR U1708 ( .A(B[487]), .B(n1139), .Z(O[488]) );
  AND U1709 ( .A(S), .B(n1140), .Z(n1139) );
  XOR U1710 ( .A(B[488]), .B(B[487]), .Z(n1140) );
  XOR U1711 ( .A(B[486]), .B(n1141), .Z(O[487]) );
  AND U1712 ( .A(S), .B(n1142), .Z(n1141) );
  XOR U1713 ( .A(B[487]), .B(B[486]), .Z(n1142) );
  XOR U1714 ( .A(B[485]), .B(n1143), .Z(O[486]) );
  AND U1715 ( .A(S), .B(n1144), .Z(n1143) );
  XOR U1716 ( .A(B[486]), .B(B[485]), .Z(n1144) );
  XOR U1717 ( .A(B[484]), .B(n1145), .Z(O[485]) );
  AND U1718 ( .A(S), .B(n1146), .Z(n1145) );
  XOR U1719 ( .A(B[485]), .B(B[484]), .Z(n1146) );
  XOR U1720 ( .A(B[483]), .B(n1147), .Z(O[484]) );
  AND U1721 ( .A(S), .B(n1148), .Z(n1147) );
  XOR U1722 ( .A(B[484]), .B(B[483]), .Z(n1148) );
  XOR U1723 ( .A(B[482]), .B(n1149), .Z(O[483]) );
  AND U1724 ( .A(S), .B(n1150), .Z(n1149) );
  XOR U1725 ( .A(B[483]), .B(B[482]), .Z(n1150) );
  XOR U1726 ( .A(B[481]), .B(n1151), .Z(O[482]) );
  AND U1727 ( .A(S), .B(n1152), .Z(n1151) );
  XOR U1728 ( .A(B[482]), .B(B[481]), .Z(n1152) );
  XOR U1729 ( .A(B[480]), .B(n1153), .Z(O[481]) );
  AND U1730 ( .A(S), .B(n1154), .Z(n1153) );
  XOR U1731 ( .A(B[481]), .B(B[480]), .Z(n1154) );
  XOR U1732 ( .A(B[479]), .B(n1155), .Z(O[480]) );
  AND U1733 ( .A(S), .B(n1156), .Z(n1155) );
  XOR U1734 ( .A(B[480]), .B(B[479]), .Z(n1156) );
  XOR U1735 ( .A(B[46]), .B(n1157), .Z(O[47]) );
  AND U1736 ( .A(S), .B(n1158), .Z(n1157) );
  XOR U1737 ( .A(B[47]), .B(B[46]), .Z(n1158) );
  XOR U1738 ( .A(B[478]), .B(n1159), .Z(O[479]) );
  AND U1739 ( .A(S), .B(n1160), .Z(n1159) );
  XOR U1740 ( .A(B[479]), .B(B[478]), .Z(n1160) );
  XOR U1741 ( .A(B[477]), .B(n1161), .Z(O[478]) );
  AND U1742 ( .A(S), .B(n1162), .Z(n1161) );
  XOR U1743 ( .A(B[478]), .B(B[477]), .Z(n1162) );
  XOR U1744 ( .A(B[476]), .B(n1163), .Z(O[477]) );
  AND U1745 ( .A(S), .B(n1164), .Z(n1163) );
  XOR U1746 ( .A(B[477]), .B(B[476]), .Z(n1164) );
  XOR U1747 ( .A(B[475]), .B(n1165), .Z(O[476]) );
  AND U1748 ( .A(S), .B(n1166), .Z(n1165) );
  XOR U1749 ( .A(B[476]), .B(B[475]), .Z(n1166) );
  XOR U1750 ( .A(B[474]), .B(n1167), .Z(O[475]) );
  AND U1751 ( .A(S), .B(n1168), .Z(n1167) );
  XOR U1752 ( .A(B[475]), .B(B[474]), .Z(n1168) );
  XOR U1753 ( .A(B[473]), .B(n1169), .Z(O[474]) );
  AND U1754 ( .A(S), .B(n1170), .Z(n1169) );
  XOR U1755 ( .A(B[474]), .B(B[473]), .Z(n1170) );
  XOR U1756 ( .A(B[472]), .B(n1171), .Z(O[473]) );
  AND U1757 ( .A(S), .B(n1172), .Z(n1171) );
  XOR U1758 ( .A(B[473]), .B(B[472]), .Z(n1172) );
  XOR U1759 ( .A(B[471]), .B(n1173), .Z(O[472]) );
  AND U1760 ( .A(S), .B(n1174), .Z(n1173) );
  XOR U1761 ( .A(B[472]), .B(B[471]), .Z(n1174) );
  XOR U1762 ( .A(B[470]), .B(n1175), .Z(O[471]) );
  AND U1763 ( .A(S), .B(n1176), .Z(n1175) );
  XOR U1764 ( .A(B[471]), .B(B[470]), .Z(n1176) );
  XOR U1765 ( .A(B[469]), .B(n1177), .Z(O[470]) );
  AND U1766 ( .A(S), .B(n1178), .Z(n1177) );
  XOR U1767 ( .A(B[470]), .B(B[469]), .Z(n1178) );
  XOR U1768 ( .A(B[45]), .B(n1179), .Z(O[46]) );
  AND U1769 ( .A(S), .B(n1180), .Z(n1179) );
  XOR U1770 ( .A(B[46]), .B(B[45]), .Z(n1180) );
  XOR U1771 ( .A(B[468]), .B(n1181), .Z(O[469]) );
  AND U1772 ( .A(S), .B(n1182), .Z(n1181) );
  XOR U1773 ( .A(B[469]), .B(B[468]), .Z(n1182) );
  XOR U1774 ( .A(B[467]), .B(n1183), .Z(O[468]) );
  AND U1775 ( .A(S), .B(n1184), .Z(n1183) );
  XOR U1776 ( .A(B[468]), .B(B[467]), .Z(n1184) );
  XOR U1777 ( .A(B[466]), .B(n1185), .Z(O[467]) );
  AND U1778 ( .A(S), .B(n1186), .Z(n1185) );
  XOR U1779 ( .A(B[467]), .B(B[466]), .Z(n1186) );
  XOR U1780 ( .A(B[465]), .B(n1187), .Z(O[466]) );
  AND U1781 ( .A(S), .B(n1188), .Z(n1187) );
  XOR U1782 ( .A(B[466]), .B(B[465]), .Z(n1188) );
  XOR U1783 ( .A(B[464]), .B(n1189), .Z(O[465]) );
  AND U1784 ( .A(S), .B(n1190), .Z(n1189) );
  XOR U1785 ( .A(B[465]), .B(B[464]), .Z(n1190) );
  XOR U1786 ( .A(B[463]), .B(n1191), .Z(O[464]) );
  AND U1787 ( .A(S), .B(n1192), .Z(n1191) );
  XOR U1788 ( .A(B[464]), .B(B[463]), .Z(n1192) );
  XOR U1789 ( .A(B[462]), .B(n1193), .Z(O[463]) );
  AND U1790 ( .A(S), .B(n1194), .Z(n1193) );
  XOR U1791 ( .A(B[463]), .B(B[462]), .Z(n1194) );
  XOR U1792 ( .A(B[461]), .B(n1195), .Z(O[462]) );
  AND U1793 ( .A(S), .B(n1196), .Z(n1195) );
  XOR U1794 ( .A(B[462]), .B(B[461]), .Z(n1196) );
  XOR U1795 ( .A(B[460]), .B(n1197), .Z(O[461]) );
  AND U1796 ( .A(S), .B(n1198), .Z(n1197) );
  XOR U1797 ( .A(B[461]), .B(B[460]), .Z(n1198) );
  XOR U1798 ( .A(B[459]), .B(n1199), .Z(O[460]) );
  AND U1799 ( .A(S), .B(n1200), .Z(n1199) );
  XOR U1800 ( .A(B[460]), .B(B[459]), .Z(n1200) );
  XOR U1801 ( .A(B[44]), .B(n1201), .Z(O[45]) );
  AND U1802 ( .A(S), .B(n1202), .Z(n1201) );
  XOR U1803 ( .A(B[45]), .B(B[44]), .Z(n1202) );
  XOR U1804 ( .A(B[458]), .B(n1203), .Z(O[459]) );
  AND U1805 ( .A(S), .B(n1204), .Z(n1203) );
  XOR U1806 ( .A(B[459]), .B(B[458]), .Z(n1204) );
  XOR U1807 ( .A(B[457]), .B(n1205), .Z(O[458]) );
  AND U1808 ( .A(S), .B(n1206), .Z(n1205) );
  XOR U1809 ( .A(B[458]), .B(B[457]), .Z(n1206) );
  XOR U1810 ( .A(B[456]), .B(n1207), .Z(O[457]) );
  AND U1811 ( .A(S), .B(n1208), .Z(n1207) );
  XOR U1812 ( .A(B[457]), .B(B[456]), .Z(n1208) );
  XOR U1813 ( .A(B[455]), .B(n1209), .Z(O[456]) );
  AND U1814 ( .A(S), .B(n1210), .Z(n1209) );
  XOR U1815 ( .A(B[456]), .B(B[455]), .Z(n1210) );
  XOR U1816 ( .A(B[454]), .B(n1211), .Z(O[455]) );
  AND U1817 ( .A(S), .B(n1212), .Z(n1211) );
  XOR U1818 ( .A(B[455]), .B(B[454]), .Z(n1212) );
  XOR U1819 ( .A(B[453]), .B(n1213), .Z(O[454]) );
  AND U1820 ( .A(S), .B(n1214), .Z(n1213) );
  XOR U1821 ( .A(B[454]), .B(B[453]), .Z(n1214) );
  XOR U1822 ( .A(B[452]), .B(n1215), .Z(O[453]) );
  AND U1823 ( .A(S), .B(n1216), .Z(n1215) );
  XOR U1824 ( .A(B[453]), .B(B[452]), .Z(n1216) );
  XOR U1825 ( .A(B[451]), .B(n1217), .Z(O[452]) );
  AND U1826 ( .A(S), .B(n1218), .Z(n1217) );
  XOR U1827 ( .A(B[452]), .B(B[451]), .Z(n1218) );
  XOR U1828 ( .A(B[450]), .B(n1219), .Z(O[451]) );
  AND U1829 ( .A(S), .B(n1220), .Z(n1219) );
  XOR U1830 ( .A(B[451]), .B(B[450]), .Z(n1220) );
  XOR U1831 ( .A(B[449]), .B(n1221), .Z(O[450]) );
  AND U1832 ( .A(S), .B(n1222), .Z(n1221) );
  XOR U1833 ( .A(B[450]), .B(B[449]), .Z(n1222) );
  XOR U1834 ( .A(B[43]), .B(n1223), .Z(O[44]) );
  AND U1835 ( .A(S), .B(n1224), .Z(n1223) );
  XOR U1836 ( .A(B[44]), .B(B[43]), .Z(n1224) );
  XOR U1837 ( .A(B[448]), .B(n1225), .Z(O[449]) );
  AND U1838 ( .A(S), .B(n1226), .Z(n1225) );
  XOR U1839 ( .A(B[449]), .B(B[448]), .Z(n1226) );
  XOR U1840 ( .A(B[447]), .B(n1227), .Z(O[448]) );
  AND U1841 ( .A(S), .B(n1228), .Z(n1227) );
  XOR U1842 ( .A(B[448]), .B(B[447]), .Z(n1228) );
  XOR U1843 ( .A(B[446]), .B(n1229), .Z(O[447]) );
  AND U1844 ( .A(S), .B(n1230), .Z(n1229) );
  XOR U1845 ( .A(B[447]), .B(B[446]), .Z(n1230) );
  XOR U1846 ( .A(B[445]), .B(n1231), .Z(O[446]) );
  AND U1847 ( .A(S), .B(n1232), .Z(n1231) );
  XOR U1848 ( .A(B[446]), .B(B[445]), .Z(n1232) );
  XOR U1849 ( .A(B[444]), .B(n1233), .Z(O[445]) );
  AND U1850 ( .A(S), .B(n1234), .Z(n1233) );
  XOR U1851 ( .A(B[445]), .B(B[444]), .Z(n1234) );
  XOR U1852 ( .A(B[443]), .B(n1235), .Z(O[444]) );
  AND U1853 ( .A(S), .B(n1236), .Z(n1235) );
  XOR U1854 ( .A(B[444]), .B(B[443]), .Z(n1236) );
  XOR U1855 ( .A(B[442]), .B(n1237), .Z(O[443]) );
  AND U1856 ( .A(S), .B(n1238), .Z(n1237) );
  XOR U1857 ( .A(B[443]), .B(B[442]), .Z(n1238) );
  XOR U1858 ( .A(B[441]), .B(n1239), .Z(O[442]) );
  AND U1859 ( .A(S), .B(n1240), .Z(n1239) );
  XOR U1860 ( .A(B[442]), .B(B[441]), .Z(n1240) );
  XOR U1861 ( .A(B[440]), .B(n1241), .Z(O[441]) );
  AND U1862 ( .A(S), .B(n1242), .Z(n1241) );
  XOR U1863 ( .A(B[441]), .B(B[440]), .Z(n1242) );
  XOR U1864 ( .A(B[439]), .B(n1243), .Z(O[440]) );
  AND U1865 ( .A(S), .B(n1244), .Z(n1243) );
  XOR U1866 ( .A(B[440]), .B(B[439]), .Z(n1244) );
  XOR U1867 ( .A(B[42]), .B(n1245), .Z(O[43]) );
  AND U1868 ( .A(S), .B(n1246), .Z(n1245) );
  XOR U1869 ( .A(B[43]), .B(B[42]), .Z(n1246) );
  XOR U1870 ( .A(B[438]), .B(n1247), .Z(O[439]) );
  AND U1871 ( .A(S), .B(n1248), .Z(n1247) );
  XOR U1872 ( .A(B[439]), .B(B[438]), .Z(n1248) );
  XOR U1873 ( .A(B[437]), .B(n1249), .Z(O[438]) );
  AND U1874 ( .A(S), .B(n1250), .Z(n1249) );
  XOR U1875 ( .A(B[438]), .B(B[437]), .Z(n1250) );
  XOR U1876 ( .A(B[436]), .B(n1251), .Z(O[437]) );
  AND U1877 ( .A(S), .B(n1252), .Z(n1251) );
  XOR U1878 ( .A(B[437]), .B(B[436]), .Z(n1252) );
  XOR U1879 ( .A(B[435]), .B(n1253), .Z(O[436]) );
  AND U1880 ( .A(S), .B(n1254), .Z(n1253) );
  XOR U1881 ( .A(B[436]), .B(B[435]), .Z(n1254) );
  XOR U1882 ( .A(B[434]), .B(n1255), .Z(O[435]) );
  AND U1883 ( .A(S), .B(n1256), .Z(n1255) );
  XOR U1884 ( .A(B[435]), .B(B[434]), .Z(n1256) );
  XOR U1885 ( .A(B[433]), .B(n1257), .Z(O[434]) );
  AND U1886 ( .A(S), .B(n1258), .Z(n1257) );
  XOR U1887 ( .A(B[434]), .B(B[433]), .Z(n1258) );
  XOR U1888 ( .A(B[432]), .B(n1259), .Z(O[433]) );
  AND U1889 ( .A(S), .B(n1260), .Z(n1259) );
  XOR U1890 ( .A(B[433]), .B(B[432]), .Z(n1260) );
  XOR U1891 ( .A(B[431]), .B(n1261), .Z(O[432]) );
  AND U1892 ( .A(S), .B(n1262), .Z(n1261) );
  XOR U1893 ( .A(B[432]), .B(B[431]), .Z(n1262) );
  XOR U1894 ( .A(B[430]), .B(n1263), .Z(O[431]) );
  AND U1895 ( .A(S), .B(n1264), .Z(n1263) );
  XOR U1896 ( .A(B[431]), .B(B[430]), .Z(n1264) );
  XOR U1897 ( .A(B[429]), .B(n1265), .Z(O[430]) );
  AND U1898 ( .A(S), .B(n1266), .Z(n1265) );
  XOR U1899 ( .A(B[430]), .B(B[429]), .Z(n1266) );
  XOR U1900 ( .A(B[41]), .B(n1267), .Z(O[42]) );
  AND U1901 ( .A(S), .B(n1268), .Z(n1267) );
  XOR U1902 ( .A(B[42]), .B(B[41]), .Z(n1268) );
  XOR U1903 ( .A(B[428]), .B(n1269), .Z(O[429]) );
  AND U1904 ( .A(S), .B(n1270), .Z(n1269) );
  XOR U1905 ( .A(B[429]), .B(B[428]), .Z(n1270) );
  XOR U1906 ( .A(B[427]), .B(n1271), .Z(O[428]) );
  AND U1907 ( .A(S), .B(n1272), .Z(n1271) );
  XOR U1908 ( .A(B[428]), .B(B[427]), .Z(n1272) );
  XOR U1909 ( .A(B[426]), .B(n1273), .Z(O[427]) );
  AND U1910 ( .A(S), .B(n1274), .Z(n1273) );
  XOR U1911 ( .A(B[427]), .B(B[426]), .Z(n1274) );
  XOR U1912 ( .A(B[425]), .B(n1275), .Z(O[426]) );
  AND U1913 ( .A(S), .B(n1276), .Z(n1275) );
  XOR U1914 ( .A(B[426]), .B(B[425]), .Z(n1276) );
  XOR U1915 ( .A(B[424]), .B(n1277), .Z(O[425]) );
  AND U1916 ( .A(S), .B(n1278), .Z(n1277) );
  XOR U1917 ( .A(B[425]), .B(B[424]), .Z(n1278) );
  XOR U1918 ( .A(B[423]), .B(n1279), .Z(O[424]) );
  AND U1919 ( .A(S), .B(n1280), .Z(n1279) );
  XOR U1920 ( .A(B[424]), .B(B[423]), .Z(n1280) );
  XOR U1921 ( .A(B[422]), .B(n1281), .Z(O[423]) );
  AND U1922 ( .A(S), .B(n1282), .Z(n1281) );
  XOR U1923 ( .A(B[423]), .B(B[422]), .Z(n1282) );
  XOR U1924 ( .A(B[421]), .B(n1283), .Z(O[422]) );
  AND U1925 ( .A(S), .B(n1284), .Z(n1283) );
  XOR U1926 ( .A(B[422]), .B(B[421]), .Z(n1284) );
  XOR U1927 ( .A(B[420]), .B(n1285), .Z(O[421]) );
  AND U1928 ( .A(S), .B(n1286), .Z(n1285) );
  XOR U1929 ( .A(B[421]), .B(B[420]), .Z(n1286) );
  XOR U1930 ( .A(B[419]), .B(n1287), .Z(O[420]) );
  AND U1931 ( .A(S), .B(n1288), .Z(n1287) );
  XOR U1932 ( .A(B[420]), .B(B[419]), .Z(n1288) );
  XOR U1933 ( .A(B[40]), .B(n1289), .Z(O[41]) );
  AND U1934 ( .A(S), .B(n1290), .Z(n1289) );
  XOR U1935 ( .A(B[41]), .B(B[40]), .Z(n1290) );
  XOR U1936 ( .A(B[418]), .B(n1291), .Z(O[419]) );
  AND U1937 ( .A(S), .B(n1292), .Z(n1291) );
  XOR U1938 ( .A(B[419]), .B(B[418]), .Z(n1292) );
  XOR U1939 ( .A(B[417]), .B(n1293), .Z(O[418]) );
  AND U1940 ( .A(S), .B(n1294), .Z(n1293) );
  XOR U1941 ( .A(B[418]), .B(B[417]), .Z(n1294) );
  XOR U1942 ( .A(B[416]), .B(n1295), .Z(O[417]) );
  AND U1943 ( .A(S), .B(n1296), .Z(n1295) );
  XOR U1944 ( .A(B[417]), .B(B[416]), .Z(n1296) );
  XOR U1945 ( .A(B[415]), .B(n1297), .Z(O[416]) );
  AND U1946 ( .A(S), .B(n1298), .Z(n1297) );
  XOR U1947 ( .A(B[416]), .B(B[415]), .Z(n1298) );
  XOR U1948 ( .A(B[414]), .B(n1299), .Z(O[415]) );
  AND U1949 ( .A(S), .B(n1300), .Z(n1299) );
  XOR U1950 ( .A(B[415]), .B(B[414]), .Z(n1300) );
  XOR U1951 ( .A(B[413]), .B(n1301), .Z(O[414]) );
  AND U1952 ( .A(S), .B(n1302), .Z(n1301) );
  XOR U1953 ( .A(B[414]), .B(B[413]), .Z(n1302) );
  XOR U1954 ( .A(B[412]), .B(n1303), .Z(O[413]) );
  AND U1955 ( .A(S), .B(n1304), .Z(n1303) );
  XOR U1956 ( .A(B[413]), .B(B[412]), .Z(n1304) );
  XOR U1957 ( .A(B[411]), .B(n1305), .Z(O[412]) );
  AND U1958 ( .A(S), .B(n1306), .Z(n1305) );
  XOR U1959 ( .A(B[412]), .B(B[411]), .Z(n1306) );
  XOR U1960 ( .A(B[410]), .B(n1307), .Z(O[411]) );
  AND U1961 ( .A(S), .B(n1308), .Z(n1307) );
  XOR U1962 ( .A(B[411]), .B(B[410]), .Z(n1308) );
  XOR U1963 ( .A(B[409]), .B(n1309), .Z(O[410]) );
  AND U1964 ( .A(S), .B(n1310), .Z(n1309) );
  XOR U1965 ( .A(B[410]), .B(B[409]), .Z(n1310) );
  XOR U1966 ( .A(B[39]), .B(n1311), .Z(O[40]) );
  AND U1967 ( .A(S), .B(n1312), .Z(n1311) );
  XOR U1968 ( .A(B[40]), .B(B[39]), .Z(n1312) );
  XOR U1969 ( .A(B[408]), .B(n1313), .Z(O[409]) );
  AND U1970 ( .A(S), .B(n1314), .Z(n1313) );
  XOR U1971 ( .A(B[409]), .B(B[408]), .Z(n1314) );
  XOR U1972 ( .A(B[407]), .B(n1315), .Z(O[408]) );
  AND U1973 ( .A(S), .B(n1316), .Z(n1315) );
  XOR U1974 ( .A(B[408]), .B(B[407]), .Z(n1316) );
  XOR U1975 ( .A(B[406]), .B(n1317), .Z(O[407]) );
  AND U1976 ( .A(S), .B(n1318), .Z(n1317) );
  XOR U1977 ( .A(B[407]), .B(B[406]), .Z(n1318) );
  XOR U1978 ( .A(B[405]), .B(n1319), .Z(O[406]) );
  AND U1979 ( .A(S), .B(n1320), .Z(n1319) );
  XOR U1980 ( .A(B[406]), .B(B[405]), .Z(n1320) );
  XOR U1981 ( .A(B[404]), .B(n1321), .Z(O[405]) );
  AND U1982 ( .A(S), .B(n1322), .Z(n1321) );
  XOR U1983 ( .A(B[405]), .B(B[404]), .Z(n1322) );
  XOR U1984 ( .A(B[403]), .B(n1323), .Z(O[404]) );
  AND U1985 ( .A(S), .B(n1324), .Z(n1323) );
  XOR U1986 ( .A(B[404]), .B(B[403]), .Z(n1324) );
  XOR U1987 ( .A(B[402]), .B(n1325), .Z(O[403]) );
  AND U1988 ( .A(S), .B(n1326), .Z(n1325) );
  XOR U1989 ( .A(B[403]), .B(B[402]), .Z(n1326) );
  XOR U1990 ( .A(B[401]), .B(n1327), .Z(O[402]) );
  AND U1991 ( .A(S), .B(n1328), .Z(n1327) );
  XOR U1992 ( .A(B[402]), .B(B[401]), .Z(n1328) );
  XOR U1993 ( .A(B[400]), .B(n1329), .Z(O[401]) );
  AND U1994 ( .A(S), .B(n1330), .Z(n1329) );
  XOR U1995 ( .A(B[401]), .B(B[400]), .Z(n1330) );
  XOR U1996 ( .A(B[399]), .B(n1331), .Z(O[400]) );
  AND U1997 ( .A(S), .B(n1332), .Z(n1331) );
  XOR U1998 ( .A(B[400]), .B(B[399]), .Z(n1332) );
  XOR U1999 ( .A(B[2]), .B(n1333), .Z(O[3]) );
  AND U2000 ( .A(S), .B(n1334), .Z(n1333) );
  XOR U2001 ( .A(B[3]), .B(B[2]), .Z(n1334) );
  XOR U2002 ( .A(B[38]), .B(n1335), .Z(O[39]) );
  AND U2003 ( .A(S), .B(n1336), .Z(n1335) );
  XOR U2004 ( .A(B[39]), .B(B[38]), .Z(n1336) );
  XOR U2005 ( .A(B[398]), .B(n1337), .Z(O[399]) );
  AND U2006 ( .A(S), .B(n1338), .Z(n1337) );
  XOR U2007 ( .A(B[399]), .B(B[398]), .Z(n1338) );
  XOR U2008 ( .A(B[397]), .B(n1339), .Z(O[398]) );
  AND U2009 ( .A(S), .B(n1340), .Z(n1339) );
  XOR U2010 ( .A(B[398]), .B(B[397]), .Z(n1340) );
  XOR U2011 ( .A(B[396]), .B(n1341), .Z(O[397]) );
  AND U2012 ( .A(S), .B(n1342), .Z(n1341) );
  XOR U2013 ( .A(B[397]), .B(B[396]), .Z(n1342) );
  XOR U2014 ( .A(B[395]), .B(n1343), .Z(O[396]) );
  AND U2015 ( .A(S), .B(n1344), .Z(n1343) );
  XOR U2016 ( .A(B[396]), .B(B[395]), .Z(n1344) );
  XOR U2017 ( .A(B[394]), .B(n1345), .Z(O[395]) );
  AND U2018 ( .A(S), .B(n1346), .Z(n1345) );
  XOR U2019 ( .A(B[395]), .B(B[394]), .Z(n1346) );
  XOR U2020 ( .A(B[393]), .B(n1347), .Z(O[394]) );
  AND U2021 ( .A(S), .B(n1348), .Z(n1347) );
  XOR U2022 ( .A(B[394]), .B(B[393]), .Z(n1348) );
  XOR U2023 ( .A(B[392]), .B(n1349), .Z(O[393]) );
  AND U2024 ( .A(S), .B(n1350), .Z(n1349) );
  XOR U2025 ( .A(B[393]), .B(B[392]), .Z(n1350) );
  XOR U2026 ( .A(B[391]), .B(n1351), .Z(O[392]) );
  AND U2027 ( .A(S), .B(n1352), .Z(n1351) );
  XOR U2028 ( .A(B[392]), .B(B[391]), .Z(n1352) );
  XOR U2029 ( .A(B[390]), .B(n1353), .Z(O[391]) );
  AND U2030 ( .A(S), .B(n1354), .Z(n1353) );
  XOR U2031 ( .A(B[391]), .B(B[390]), .Z(n1354) );
  XOR U2032 ( .A(B[389]), .B(n1355), .Z(O[390]) );
  AND U2033 ( .A(S), .B(n1356), .Z(n1355) );
  XOR U2034 ( .A(B[390]), .B(B[389]), .Z(n1356) );
  XOR U2035 ( .A(B[37]), .B(n1357), .Z(O[38]) );
  AND U2036 ( .A(S), .B(n1358), .Z(n1357) );
  XOR U2037 ( .A(B[38]), .B(B[37]), .Z(n1358) );
  XOR U2038 ( .A(B[388]), .B(n1359), .Z(O[389]) );
  AND U2039 ( .A(S), .B(n1360), .Z(n1359) );
  XOR U2040 ( .A(B[389]), .B(B[388]), .Z(n1360) );
  XOR U2041 ( .A(B[387]), .B(n1361), .Z(O[388]) );
  AND U2042 ( .A(S), .B(n1362), .Z(n1361) );
  XOR U2043 ( .A(B[388]), .B(B[387]), .Z(n1362) );
  XOR U2044 ( .A(B[386]), .B(n1363), .Z(O[387]) );
  AND U2045 ( .A(S), .B(n1364), .Z(n1363) );
  XOR U2046 ( .A(B[387]), .B(B[386]), .Z(n1364) );
  XOR U2047 ( .A(B[385]), .B(n1365), .Z(O[386]) );
  AND U2048 ( .A(S), .B(n1366), .Z(n1365) );
  XOR U2049 ( .A(B[386]), .B(B[385]), .Z(n1366) );
  XOR U2050 ( .A(B[384]), .B(n1367), .Z(O[385]) );
  AND U2051 ( .A(S), .B(n1368), .Z(n1367) );
  XOR U2052 ( .A(B[385]), .B(B[384]), .Z(n1368) );
  XOR U2053 ( .A(B[383]), .B(n1369), .Z(O[384]) );
  AND U2054 ( .A(S), .B(n1370), .Z(n1369) );
  XOR U2055 ( .A(B[384]), .B(B[383]), .Z(n1370) );
  XOR U2056 ( .A(B[382]), .B(n1371), .Z(O[383]) );
  AND U2057 ( .A(S), .B(n1372), .Z(n1371) );
  XOR U2058 ( .A(B[383]), .B(B[382]), .Z(n1372) );
  XOR U2059 ( .A(B[381]), .B(n1373), .Z(O[382]) );
  AND U2060 ( .A(S), .B(n1374), .Z(n1373) );
  XOR U2061 ( .A(B[382]), .B(B[381]), .Z(n1374) );
  XOR U2062 ( .A(B[380]), .B(n1375), .Z(O[381]) );
  AND U2063 ( .A(S), .B(n1376), .Z(n1375) );
  XOR U2064 ( .A(B[381]), .B(B[380]), .Z(n1376) );
  XOR U2065 ( .A(B[379]), .B(n1377), .Z(O[380]) );
  AND U2066 ( .A(S), .B(n1378), .Z(n1377) );
  XOR U2067 ( .A(B[380]), .B(B[379]), .Z(n1378) );
  XOR U2068 ( .A(B[36]), .B(n1379), .Z(O[37]) );
  AND U2069 ( .A(S), .B(n1380), .Z(n1379) );
  XOR U2070 ( .A(B[37]), .B(B[36]), .Z(n1380) );
  XOR U2071 ( .A(B[378]), .B(n1381), .Z(O[379]) );
  AND U2072 ( .A(S), .B(n1382), .Z(n1381) );
  XOR U2073 ( .A(B[379]), .B(B[378]), .Z(n1382) );
  XOR U2074 ( .A(B[377]), .B(n1383), .Z(O[378]) );
  AND U2075 ( .A(S), .B(n1384), .Z(n1383) );
  XOR U2076 ( .A(B[378]), .B(B[377]), .Z(n1384) );
  XOR U2077 ( .A(B[376]), .B(n1385), .Z(O[377]) );
  AND U2078 ( .A(S), .B(n1386), .Z(n1385) );
  XOR U2079 ( .A(B[377]), .B(B[376]), .Z(n1386) );
  XOR U2080 ( .A(B[375]), .B(n1387), .Z(O[376]) );
  AND U2081 ( .A(S), .B(n1388), .Z(n1387) );
  XOR U2082 ( .A(B[376]), .B(B[375]), .Z(n1388) );
  XOR U2083 ( .A(B[374]), .B(n1389), .Z(O[375]) );
  AND U2084 ( .A(S), .B(n1390), .Z(n1389) );
  XOR U2085 ( .A(B[375]), .B(B[374]), .Z(n1390) );
  XOR U2086 ( .A(B[373]), .B(n1391), .Z(O[374]) );
  AND U2087 ( .A(S), .B(n1392), .Z(n1391) );
  XOR U2088 ( .A(B[374]), .B(B[373]), .Z(n1392) );
  XOR U2089 ( .A(B[372]), .B(n1393), .Z(O[373]) );
  AND U2090 ( .A(S), .B(n1394), .Z(n1393) );
  XOR U2091 ( .A(B[373]), .B(B[372]), .Z(n1394) );
  XOR U2092 ( .A(B[371]), .B(n1395), .Z(O[372]) );
  AND U2093 ( .A(S), .B(n1396), .Z(n1395) );
  XOR U2094 ( .A(B[372]), .B(B[371]), .Z(n1396) );
  XOR U2095 ( .A(B[370]), .B(n1397), .Z(O[371]) );
  AND U2096 ( .A(S), .B(n1398), .Z(n1397) );
  XOR U2097 ( .A(B[371]), .B(B[370]), .Z(n1398) );
  XOR U2098 ( .A(B[369]), .B(n1399), .Z(O[370]) );
  AND U2099 ( .A(S), .B(n1400), .Z(n1399) );
  XOR U2100 ( .A(B[370]), .B(B[369]), .Z(n1400) );
  XOR U2101 ( .A(B[35]), .B(n1401), .Z(O[36]) );
  AND U2102 ( .A(S), .B(n1402), .Z(n1401) );
  XOR U2103 ( .A(B[36]), .B(B[35]), .Z(n1402) );
  XOR U2104 ( .A(B[368]), .B(n1403), .Z(O[369]) );
  AND U2105 ( .A(S), .B(n1404), .Z(n1403) );
  XOR U2106 ( .A(B[369]), .B(B[368]), .Z(n1404) );
  XOR U2107 ( .A(B[367]), .B(n1405), .Z(O[368]) );
  AND U2108 ( .A(S), .B(n1406), .Z(n1405) );
  XOR U2109 ( .A(B[368]), .B(B[367]), .Z(n1406) );
  XOR U2110 ( .A(B[366]), .B(n1407), .Z(O[367]) );
  AND U2111 ( .A(S), .B(n1408), .Z(n1407) );
  XOR U2112 ( .A(B[367]), .B(B[366]), .Z(n1408) );
  XOR U2113 ( .A(B[365]), .B(n1409), .Z(O[366]) );
  AND U2114 ( .A(S), .B(n1410), .Z(n1409) );
  XOR U2115 ( .A(B[366]), .B(B[365]), .Z(n1410) );
  XOR U2116 ( .A(B[364]), .B(n1411), .Z(O[365]) );
  AND U2117 ( .A(S), .B(n1412), .Z(n1411) );
  XOR U2118 ( .A(B[365]), .B(B[364]), .Z(n1412) );
  XOR U2119 ( .A(B[363]), .B(n1413), .Z(O[364]) );
  AND U2120 ( .A(S), .B(n1414), .Z(n1413) );
  XOR U2121 ( .A(B[364]), .B(B[363]), .Z(n1414) );
  XOR U2122 ( .A(B[362]), .B(n1415), .Z(O[363]) );
  AND U2123 ( .A(S), .B(n1416), .Z(n1415) );
  XOR U2124 ( .A(B[363]), .B(B[362]), .Z(n1416) );
  XOR U2125 ( .A(B[361]), .B(n1417), .Z(O[362]) );
  AND U2126 ( .A(S), .B(n1418), .Z(n1417) );
  XOR U2127 ( .A(B[362]), .B(B[361]), .Z(n1418) );
  XOR U2128 ( .A(B[360]), .B(n1419), .Z(O[361]) );
  AND U2129 ( .A(S), .B(n1420), .Z(n1419) );
  XOR U2130 ( .A(B[361]), .B(B[360]), .Z(n1420) );
  XOR U2131 ( .A(B[359]), .B(n1421), .Z(O[360]) );
  AND U2132 ( .A(S), .B(n1422), .Z(n1421) );
  XOR U2133 ( .A(B[360]), .B(B[359]), .Z(n1422) );
  XOR U2134 ( .A(B[34]), .B(n1423), .Z(O[35]) );
  AND U2135 ( .A(S), .B(n1424), .Z(n1423) );
  XOR U2136 ( .A(B[35]), .B(B[34]), .Z(n1424) );
  XOR U2137 ( .A(B[358]), .B(n1425), .Z(O[359]) );
  AND U2138 ( .A(S), .B(n1426), .Z(n1425) );
  XOR U2139 ( .A(B[359]), .B(B[358]), .Z(n1426) );
  XOR U2140 ( .A(B[357]), .B(n1427), .Z(O[358]) );
  AND U2141 ( .A(S), .B(n1428), .Z(n1427) );
  XOR U2142 ( .A(B[358]), .B(B[357]), .Z(n1428) );
  XOR U2143 ( .A(B[356]), .B(n1429), .Z(O[357]) );
  AND U2144 ( .A(S), .B(n1430), .Z(n1429) );
  XOR U2145 ( .A(B[357]), .B(B[356]), .Z(n1430) );
  XOR U2146 ( .A(B[355]), .B(n1431), .Z(O[356]) );
  AND U2147 ( .A(S), .B(n1432), .Z(n1431) );
  XOR U2148 ( .A(B[356]), .B(B[355]), .Z(n1432) );
  XOR U2149 ( .A(B[354]), .B(n1433), .Z(O[355]) );
  AND U2150 ( .A(S), .B(n1434), .Z(n1433) );
  XOR U2151 ( .A(B[355]), .B(B[354]), .Z(n1434) );
  XOR U2152 ( .A(B[353]), .B(n1435), .Z(O[354]) );
  AND U2153 ( .A(S), .B(n1436), .Z(n1435) );
  XOR U2154 ( .A(B[354]), .B(B[353]), .Z(n1436) );
  XOR U2155 ( .A(B[352]), .B(n1437), .Z(O[353]) );
  AND U2156 ( .A(S), .B(n1438), .Z(n1437) );
  XOR U2157 ( .A(B[353]), .B(B[352]), .Z(n1438) );
  XOR U2158 ( .A(B[351]), .B(n1439), .Z(O[352]) );
  AND U2159 ( .A(S), .B(n1440), .Z(n1439) );
  XOR U2160 ( .A(B[352]), .B(B[351]), .Z(n1440) );
  XOR U2161 ( .A(B[350]), .B(n1441), .Z(O[351]) );
  AND U2162 ( .A(S), .B(n1442), .Z(n1441) );
  XOR U2163 ( .A(B[351]), .B(B[350]), .Z(n1442) );
  XOR U2164 ( .A(B[349]), .B(n1443), .Z(O[350]) );
  AND U2165 ( .A(S), .B(n1444), .Z(n1443) );
  XOR U2166 ( .A(B[350]), .B(B[349]), .Z(n1444) );
  XOR U2167 ( .A(B[33]), .B(n1445), .Z(O[34]) );
  AND U2168 ( .A(S), .B(n1446), .Z(n1445) );
  XOR U2169 ( .A(B[34]), .B(B[33]), .Z(n1446) );
  XOR U2170 ( .A(B[348]), .B(n1447), .Z(O[349]) );
  AND U2171 ( .A(S), .B(n1448), .Z(n1447) );
  XOR U2172 ( .A(B[349]), .B(B[348]), .Z(n1448) );
  XOR U2173 ( .A(B[347]), .B(n1449), .Z(O[348]) );
  AND U2174 ( .A(S), .B(n1450), .Z(n1449) );
  XOR U2175 ( .A(B[348]), .B(B[347]), .Z(n1450) );
  XOR U2176 ( .A(B[346]), .B(n1451), .Z(O[347]) );
  AND U2177 ( .A(S), .B(n1452), .Z(n1451) );
  XOR U2178 ( .A(B[347]), .B(B[346]), .Z(n1452) );
  XOR U2179 ( .A(B[345]), .B(n1453), .Z(O[346]) );
  AND U2180 ( .A(S), .B(n1454), .Z(n1453) );
  XOR U2181 ( .A(B[346]), .B(B[345]), .Z(n1454) );
  XOR U2182 ( .A(B[344]), .B(n1455), .Z(O[345]) );
  AND U2183 ( .A(S), .B(n1456), .Z(n1455) );
  XOR U2184 ( .A(B[345]), .B(B[344]), .Z(n1456) );
  XOR U2185 ( .A(B[343]), .B(n1457), .Z(O[344]) );
  AND U2186 ( .A(S), .B(n1458), .Z(n1457) );
  XOR U2187 ( .A(B[344]), .B(B[343]), .Z(n1458) );
  XOR U2188 ( .A(B[342]), .B(n1459), .Z(O[343]) );
  AND U2189 ( .A(S), .B(n1460), .Z(n1459) );
  XOR U2190 ( .A(B[343]), .B(B[342]), .Z(n1460) );
  XOR U2191 ( .A(B[341]), .B(n1461), .Z(O[342]) );
  AND U2192 ( .A(S), .B(n1462), .Z(n1461) );
  XOR U2193 ( .A(B[342]), .B(B[341]), .Z(n1462) );
  XOR U2194 ( .A(B[340]), .B(n1463), .Z(O[341]) );
  AND U2195 ( .A(S), .B(n1464), .Z(n1463) );
  XOR U2196 ( .A(B[341]), .B(B[340]), .Z(n1464) );
  XOR U2197 ( .A(B[339]), .B(n1465), .Z(O[340]) );
  AND U2198 ( .A(S), .B(n1466), .Z(n1465) );
  XOR U2199 ( .A(B[340]), .B(B[339]), .Z(n1466) );
  XOR U2200 ( .A(B[32]), .B(n1467), .Z(O[33]) );
  AND U2201 ( .A(S), .B(n1468), .Z(n1467) );
  XOR U2202 ( .A(B[33]), .B(B[32]), .Z(n1468) );
  XOR U2203 ( .A(B[338]), .B(n1469), .Z(O[339]) );
  AND U2204 ( .A(S), .B(n1470), .Z(n1469) );
  XOR U2205 ( .A(B[339]), .B(B[338]), .Z(n1470) );
  XOR U2206 ( .A(B[337]), .B(n1471), .Z(O[338]) );
  AND U2207 ( .A(S), .B(n1472), .Z(n1471) );
  XOR U2208 ( .A(B[338]), .B(B[337]), .Z(n1472) );
  XOR U2209 ( .A(B[336]), .B(n1473), .Z(O[337]) );
  AND U2210 ( .A(S), .B(n1474), .Z(n1473) );
  XOR U2211 ( .A(B[337]), .B(B[336]), .Z(n1474) );
  XOR U2212 ( .A(B[335]), .B(n1475), .Z(O[336]) );
  AND U2213 ( .A(S), .B(n1476), .Z(n1475) );
  XOR U2214 ( .A(B[336]), .B(B[335]), .Z(n1476) );
  XOR U2215 ( .A(B[334]), .B(n1477), .Z(O[335]) );
  AND U2216 ( .A(S), .B(n1478), .Z(n1477) );
  XOR U2217 ( .A(B[335]), .B(B[334]), .Z(n1478) );
  XOR U2218 ( .A(B[333]), .B(n1479), .Z(O[334]) );
  AND U2219 ( .A(S), .B(n1480), .Z(n1479) );
  XOR U2220 ( .A(B[334]), .B(B[333]), .Z(n1480) );
  XOR U2221 ( .A(B[332]), .B(n1481), .Z(O[333]) );
  AND U2222 ( .A(S), .B(n1482), .Z(n1481) );
  XOR U2223 ( .A(B[333]), .B(B[332]), .Z(n1482) );
  XOR U2224 ( .A(B[331]), .B(n1483), .Z(O[332]) );
  AND U2225 ( .A(S), .B(n1484), .Z(n1483) );
  XOR U2226 ( .A(B[332]), .B(B[331]), .Z(n1484) );
  XOR U2227 ( .A(B[330]), .B(n1485), .Z(O[331]) );
  AND U2228 ( .A(S), .B(n1486), .Z(n1485) );
  XOR U2229 ( .A(B[331]), .B(B[330]), .Z(n1486) );
  XOR U2230 ( .A(B[329]), .B(n1487), .Z(O[330]) );
  AND U2231 ( .A(S), .B(n1488), .Z(n1487) );
  XOR U2232 ( .A(B[330]), .B(B[329]), .Z(n1488) );
  XOR U2233 ( .A(B[31]), .B(n1489), .Z(O[32]) );
  AND U2234 ( .A(S), .B(n1490), .Z(n1489) );
  XOR U2235 ( .A(B[32]), .B(B[31]), .Z(n1490) );
  XOR U2236 ( .A(B[328]), .B(n1491), .Z(O[329]) );
  AND U2237 ( .A(S), .B(n1492), .Z(n1491) );
  XOR U2238 ( .A(B[329]), .B(B[328]), .Z(n1492) );
  XOR U2239 ( .A(B[327]), .B(n1493), .Z(O[328]) );
  AND U2240 ( .A(S), .B(n1494), .Z(n1493) );
  XOR U2241 ( .A(B[328]), .B(B[327]), .Z(n1494) );
  XOR U2242 ( .A(B[326]), .B(n1495), .Z(O[327]) );
  AND U2243 ( .A(S), .B(n1496), .Z(n1495) );
  XOR U2244 ( .A(B[327]), .B(B[326]), .Z(n1496) );
  XOR U2245 ( .A(B[325]), .B(n1497), .Z(O[326]) );
  AND U2246 ( .A(S), .B(n1498), .Z(n1497) );
  XOR U2247 ( .A(B[326]), .B(B[325]), .Z(n1498) );
  XOR U2248 ( .A(B[324]), .B(n1499), .Z(O[325]) );
  AND U2249 ( .A(S), .B(n1500), .Z(n1499) );
  XOR U2250 ( .A(B[325]), .B(B[324]), .Z(n1500) );
  XOR U2251 ( .A(B[323]), .B(n1501), .Z(O[324]) );
  AND U2252 ( .A(S), .B(n1502), .Z(n1501) );
  XOR U2253 ( .A(B[324]), .B(B[323]), .Z(n1502) );
  XOR U2254 ( .A(B[322]), .B(n1503), .Z(O[323]) );
  AND U2255 ( .A(S), .B(n1504), .Z(n1503) );
  XOR U2256 ( .A(B[323]), .B(B[322]), .Z(n1504) );
  XOR U2257 ( .A(B[321]), .B(n1505), .Z(O[322]) );
  AND U2258 ( .A(S), .B(n1506), .Z(n1505) );
  XOR U2259 ( .A(B[322]), .B(B[321]), .Z(n1506) );
  XOR U2260 ( .A(B[320]), .B(n1507), .Z(O[321]) );
  AND U2261 ( .A(S), .B(n1508), .Z(n1507) );
  XOR U2262 ( .A(B[321]), .B(B[320]), .Z(n1508) );
  XOR U2263 ( .A(B[319]), .B(n1509), .Z(O[320]) );
  AND U2264 ( .A(S), .B(n1510), .Z(n1509) );
  XOR U2265 ( .A(B[320]), .B(B[319]), .Z(n1510) );
  XOR U2266 ( .A(B[30]), .B(n1511), .Z(O[31]) );
  AND U2267 ( .A(S), .B(n1512), .Z(n1511) );
  XOR U2268 ( .A(B[31]), .B(B[30]), .Z(n1512) );
  XOR U2269 ( .A(B[318]), .B(n1513), .Z(O[319]) );
  AND U2270 ( .A(S), .B(n1514), .Z(n1513) );
  XOR U2271 ( .A(B[319]), .B(B[318]), .Z(n1514) );
  XOR U2272 ( .A(B[317]), .B(n1515), .Z(O[318]) );
  AND U2273 ( .A(S), .B(n1516), .Z(n1515) );
  XOR U2274 ( .A(B[318]), .B(B[317]), .Z(n1516) );
  XOR U2275 ( .A(B[316]), .B(n1517), .Z(O[317]) );
  AND U2276 ( .A(S), .B(n1518), .Z(n1517) );
  XOR U2277 ( .A(B[317]), .B(B[316]), .Z(n1518) );
  XOR U2278 ( .A(B[315]), .B(n1519), .Z(O[316]) );
  AND U2279 ( .A(S), .B(n1520), .Z(n1519) );
  XOR U2280 ( .A(B[316]), .B(B[315]), .Z(n1520) );
  XOR U2281 ( .A(B[314]), .B(n1521), .Z(O[315]) );
  AND U2282 ( .A(S), .B(n1522), .Z(n1521) );
  XOR U2283 ( .A(B[315]), .B(B[314]), .Z(n1522) );
  XOR U2284 ( .A(B[313]), .B(n1523), .Z(O[314]) );
  AND U2285 ( .A(S), .B(n1524), .Z(n1523) );
  XOR U2286 ( .A(B[314]), .B(B[313]), .Z(n1524) );
  XOR U2287 ( .A(B[312]), .B(n1525), .Z(O[313]) );
  AND U2288 ( .A(S), .B(n1526), .Z(n1525) );
  XOR U2289 ( .A(B[313]), .B(B[312]), .Z(n1526) );
  XOR U2290 ( .A(B[311]), .B(n1527), .Z(O[312]) );
  AND U2291 ( .A(S), .B(n1528), .Z(n1527) );
  XOR U2292 ( .A(B[312]), .B(B[311]), .Z(n1528) );
  XOR U2293 ( .A(B[310]), .B(n1529), .Z(O[311]) );
  AND U2294 ( .A(S), .B(n1530), .Z(n1529) );
  XOR U2295 ( .A(B[311]), .B(B[310]), .Z(n1530) );
  XOR U2296 ( .A(B[309]), .B(n1531), .Z(O[310]) );
  AND U2297 ( .A(S), .B(n1532), .Z(n1531) );
  XOR U2298 ( .A(B[310]), .B(B[309]), .Z(n1532) );
  XOR U2299 ( .A(B[29]), .B(n1533), .Z(O[30]) );
  AND U2300 ( .A(S), .B(n1534), .Z(n1533) );
  XOR U2301 ( .A(B[30]), .B(B[29]), .Z(n1534) );
  XOR U2302 ( .A(B[308]), .B(n1535), .Z(O[309]) );
  AND U2303 ( .A(S), .B(n1536), .Z(n1535) );
  XOR U2304 ( .A(B[309]), .B(B[308]), .Z(n1536) );
  XOR U2305 ( .A(B[307]), .B(n1537), .Z(O[308]) );
  AND U2306 ( .A(S), .B(n1538), .Z(n1537) );
  XOR U2307 ( .A(B[308]), .B(B[307]), .Z(n1538) );
  XOR U2308 ( .A(B[306]), .B(n1539), .Z(O[307]) );
  AND U2309 ( .A(S), .B(n1540), .Z(n1539) );
  XOR U2310 ( .A(B[307]), .B(B[306]), .Z(n1540) );
  XOR U2311 ( .A(B[305]), .B(n1541), .Z(O[306]) );
  AND U2312 ( .A(S), .B(n1542), .Z(n1541) );
  XOR U2313 ( .A(B[306]), .B(B[305]), .Z(n1542) );
  XOR U2314 ( .A(B[304]), .B(n1543), .Z(O[305]) );
  AND U2315 ( .A(S), .B(n1544), .Z(n1543) );
  XOR U2316 ( .A(B[305]), .B(B[304]), .Z(n1544) );
  XOR U2317 ( .A(B[303]), .B(n1545), .Z(O[304]) );
  AND U2318 ( .A(S), .B(n1546), .Z(n1545) );
  XOR U2319 ( .A(B[304]), .B(B[303]), .Z(n1546) );
  XOR U2320 ( .A(B[302]), .B(n1547), .Z(O[303]) );
  AND U2321 ( .A(S), .B(n1548), .Z(n1547) );
  XOR U2322 ( .A(B[303]), .B(B[302]), .Z(n1548) );
  XOR U2323 ( .A(B[301]), .B(n1549), .Z(O[302]) );
  AND U2324 ( .A(S), .B(n1550), .Z(n1549) );
  XOR U2325 ( .A(B[302]), .B(B[301]), .Z(n1550) );
  XOR U2326 ( .A(B[300]), .B(n1551), .Z(O[301]) );
  AND U2327 ( .A(S), .B(n1552), .Z(n1551) );
  XOR U2328 ( .A(B[301]), .B(B[300]), .Z(n1552) );
  XOR U2329 ( .A(B[299]), .B(n1553), .Z(O[300]) );
  AND U2330 ( .A(S), .B(n1554), .Z(n1553) );
  XOR U2331 ( .A(B[300]), .B(B[299]), .Z(n1554) );
  XOR U2332 ( .A(B[1]), .B(n1555), .Z(O[2]) );
  AND U2333 ( .A(S), .B(n1556), .Z(n1555) );
  XOR U2334 ( .A(B[2]), .B(B[1]), .Z(n1556) );
  XOR U2335 ( .A(B[28]), .B(n1557), .Z(O[29]) );
  AND U2336 ( .A(S), .B(n1558), .Z(n1557) );
  XOR U2337 ( .A(B[29]), .B(B[28]), .Z(n1558) );
  XOR U2338 ( .A(B[298]), .B(n1559), .Z(O[299]) );
  AND U2339 ( .A(S), .B(n1560), .Z(n1559) );
  XOR U2340 ( .A(B[299]), .B(B[298]), .Z(n1560) );
  XOR U2341 ( .A(B[297]), .B(n1561), .Z(O[298]) );
  AND U2342 ( .A(S), .B(n1562), .Z(n1561) );
  XOR U2343 ( .A(B[298]), .B(B[297]), .Z(n1562) );
  XOR U2344 ( .A(B[296]), .B(n1563), .Z(O[297]) );
  AND U2345 ( .A(S), .B(n1564), .Z(n1563) );
  XOR U2346 ( .A(B[297]), .B(B[296]), .Z(n1564) );
  XOR U2347 ( .A(B[295]), .B(n1565), .Z(O[296]) );
  AND U2348 ( .A(S), .B(n1566), .Z(n1565) );
  XOR U2349 ( .A(B[296]), .B(B[295]), .Z(n1566) );
  XOR U2350 ( .A(B[294]), .B(n1567), .Z(O[295]) );
  AND U2351 ( .A(S), .B(n1568), .Z(n1567) );
  XOR U2352 ( .A(B[295]), .B(B[294]), .Z(n1568) );
  XOR U2353 ( .A(B[293]), .B(n1569), .Z(O[294]) );
  AND U2354 ( .A(S), .B(n1570), .Z(n1569) );
  XOR U2355 ( .A(B[294]), .B(B[293]), .Z(n1570) );
  XOR U2356 ( .A(B[292]), .B(n1571), .Z(O[293]) );
  AND U2357 ( .A(S), .B(n1572), .Z(n1571) );
  XOR U2358 ( .A(B[293]), .B(B[292]), .Z(n1572) );
  XOR U2359 ( .A(B[291]), .B(n1573), .Z(O[292]) );
  AND U2360 ( .A(S), .B(n1574), .Z(n1573) );
  XOR U2361 ( .A(B[292]), .B(B[291]), .Z(n1574) );
  XOR U2362 ( .A(B[290]), .B(n1575), .Z(O[291]) );
  AND U2363 ( .A(S), .B(n1576), .Z(n1575) );
  XOR U2364 ( .A(B[291]), .B(B[290]), .Z(n1576) );
  XOR U2365 ( .A(B[289]), .B(n1577), .Z(O[290]) );
  AND U2366 ( .A(S), .B(n1578), .Z(n1577) );
  XOR U2367 ( .A(B[290]), .B(B[289]), .Z(n1578) );
  XOR U2368 ( .A(B[27]), .B(n1579), .Z(O[28]) );
  AND U2369 ( .A(S), .B(n1580), .Z(n1579) );
  XOR U2370 ( .A(B[28]), .B(B[27]), .Z(n1580) );
  XOR U2371 ( .A(B[288]), .B(n1581), .Z(O[289]) );
  AND U2372 ( .A(S), .B(n1582), .Z(n1581) );
  XOR U2373 ( .A(B[289]), .B(B[288]), .Z(n1582) );
  XOR U2374 ( .A(B[287]), .B(n1583), .Z(O[288]) );
  AND U2375 ( .A(S), .B(n1584), .Z(n1583) );
  XOR U2376 ( .A(B[288]), .B(B[287]), .Z(n1584) );
  XOR U2377 ( .A(B[286]), .B(n1585), .Z(O[287]) );
  AND U2378 ( .A(S), .B(n1586), .Z(n1585) );
  XOR U2379 ( .A(B[287]), .B(B[286]), .Z(n1586) );
  XOR U2380 ( .A(B[285]), .B(n1587), .Z(O[286]) );
  AND U2381 ( .A(S), .B(n1588), .Z(n1587) );
  XOR U2382 ( .A(B[286]), .B(B[285]), .Z(n1588) );
  XOR U2383 ( .A(B[284]), .B(n1589), .Z(O[285]) );
  AND U2384 ( .A(S), .B(n1590), .Z(n1589) );
  XOR U2385 ( .A(B[285]), .B(B[284]), .Z(n1590) );
  XOR U2386 ( .A(B[283]), .B(n1591), .Z(O[284]) );
  AND U2387 ( .A(S), .B(n1592), .Z(n1591) );
  XOR U2388 ( .A(B[284]), .B(B[283]), .Z(n1592) );
  XOR U2389 ( .A(B[282]), .B(n1593), .Z(O[283]) );
  AND U2390 ( .A(S), .B(n1594), .Z(n1593) );
  XOR U2391 ( .A(B[283]), .B(B[282]), .Z(n1594) );
  XOR U2392 ( .A(B[281]), .B(n1595), .Z(O[282]) );
  AND U2393 ( .A(S), .B(n1596), .Z(n1595) );
  XOR U2394 ( .A(B[282]), .B(B[281]), .Z(n1596) );
  XOR U2395 ( .A(B[280]), .B(n1597), .Z(O[281]) );
  AND U2396 ( .A(S), .B(n1598), .Z(n1597) );
  XOR U2397 ( .A(B[281]), .B(B[280]), .Z(n1598) );
  XOR U2398 ( .A(B[279]), .B(n1599), .Z(O[280]) );
  AND U2399 ( .A(S), .B(n1600), .Z(n1599) );
  XOR U2400 ( .A(B[280]), .B(B[279]), .Z(n1600) );
  XOR U2401 ( .A(B[26]), .B(n1601), .Z(O[27]) );
  AND U2402 ( .A(S), .B(n1602), .Z(n1601) );
  XOR U2403 ( .A(B[27]), .B(B[26]), .Z(n1602) );
  XOR U2404 ( .A(B[278]), .B(n1603), .Z(O[279]) );
  AND U2405 ( .A(S), .B(n1604), .Z(n1603) );
  XOR U2406 ( .A(B[279]), .B(B[278]), .Z(n1604) );
  XOR U2407 ( .A(B[277]), .B(n1605), .Z(O[278]) );
  AND U2408 ( .A(S), .B(n1606), .Z(n1605) );
  XOR U2409 ( .A(B[278]), .B(B[277]), .Z(n1606) );
  XOR U2410 ( .A(B[276]), .B(n1607), .Z(O[277]) );
  AND U2411 ( .A(S), .B(n1608), .Z(n1607) );
  XOR U2412 ( .A(B[277]), .B(B[276]), .Z(n1608) );
  XOR U2413 ( .A(B[275]), .B(n1609), .Z(O[276]) );
  AND U2414 ( .A(S), .B(n1610), .Z(n1609) );
  XOR U2415 ( .A(B[276]), .B(B[275]), .Z(n1610) );
  XOR U2416 ( .A(B[274]), .B(n1611), .Z(O[275]) );
  AND U2417 ( .A(S), .B(n1612), .Z(n1611) );
  XOR U2418 ( .A(B[275]), .B(B[274]), .Z(n1612) );
  XOR U2419 ( .A(B[273]), .B(n1613), .Z(O[274]) );
  AND U2420 ( .A(S), .B(n1614), .Z(n1613) );
  XOR U2421 ( .A(B[274]), .B(B[273]), .Z(n1614) );
  XOR U2422 ( .A(B[272]), .B(n1615), .Z(O[273]) );
  AND U2423 ( .A(S), .B(n1616), .Z(n1615) );
  XOR U2424 ( .A(B[273]), .B(B[272]), .Z(n1616) );
  XOR U2425 ( .A(B[271]), .B(n1617), .Z(O[272]) );
  AND U2426 ( .A(S), .B(n1618), .Z(n1617) );
  XOR U2427 ( .A(B[272]), .B(B[271]), .Z(n1618) );
  XOR U2428 ( .A(B[270]), .B(n1619), .Z(O[271]) );
  AND U2429 ( .A(S), .B(n1620), .Z(n1619) );
  XOR U2430 ( .A(B[271]), .B(B[270]), .Z(n1620) );
  XOR U2431 ( .A(B[269]), .B(n1621), .Z(O[270]) );
  AND U2432 ( .A(S), .B(n1622), .Z(n1621) );
  XOR U2433 ( .A(B[270]), .B(B[269]), .Z(n1622) );
  XOR U2434 ( .A(B[25]), .B(n1623), .Z(O[26]) );
  AND U2435 ( .A(S), .B(n1624), .Z(n1623) );
  XOR U2436 ( .A(B[26]), .B(B[25]), .Z(n1624) );
  XOR U2437 ( .A(B[268]), .B(n1625), .Z(O[269]) );
  AND U2438 ( .A(S), .B(n1626), .Z(n1625) );
  XOR U2439 ( .A(B[269]), .B(B[268]), .Z(n1626) );
  XOR U2440 ( .A(B[267]), .B(n1627), .Z(O[268]) );
  AND U2441 ( .A(S), .B(n1628), .Z(n1627) );
  XOR U2442 ( .A(B[268]), .B(B[267]), .Z(n1628) );
  XOR U2443 ( .A(B[266]), .B(n1629), .Z(O[267]) );
  AND U2444 ( .A(S), .B(n1630), .Z(n1629) );
  XOR U2445 ( .A(B[267]), .B(B[266]), .Z(n1630) );
  XOR U2446 ( .A(B[265]), .B(n1631), .Z(O[266]) );
  AND U2447 ( .A(S), .B(n1632), .Z(n1631) );
  XOR U2448 ( .A(B[266]), .B(B[265]), .Z(n1632) );
  XOR U2449 ( .A(B[264]), .B(n1633), .Z(O[265]) );
  AND U2450 ( .A(S), .B(n1634), .Z(n1633) );
  XOR U2451 ( .A(B[265]), .B(B[264]), .Z(n1634) );
  XOR U2452 ( .A(B[263]), .B(n1635), .Z(O[264]) );
  AND U2453 ( .A(S), .B(n1636), .Z(n1635) );
  XOR U2454 ( .A(B[264]), .B(B[263]), .Z(n1636) );
  XOR U2455 ( .A(B[262]), .B(n1637), .Z(O[263]) );
  AND U2456 ( .A(S), .B(n1638), .Z(n1637) );
  XOR U2457 ( .A(B[263]), .B(B[262]), .Z(n1638) );
  XOR U2458 ( .A(B[261]), .B(n1639), .Z(O[262]) );
  AND U2459 ( .A(S), .B(n1640), .Z(n1639) );
  XOR U2460 ( .A(B[262]), .B(B[261]), .Z(n1640) );
  XOR U2461 ( .A(B[260]), .B(n1641), .Z(O[261]) );
  AND U2462 ( .A(S), .B(n1642), .Z(n1641) );
  XOR U2463 ( .A(B[261]), .B(B[260]), .Z(n1642) );
  XOR U2464 ( .A(B[259]), .B(n1643), .Z(O[260]) );
  AND U2465 ( .A(S), .B(n1644), .Z(n1643) );
  XOR U2466 ( .A(B[260]), .B(B[259]), .Z(n1644) );
  XOR U2467 ( .A(B[24]), .B(n1645), .Z(O[25]) );
  AND U2468 ( .A(S), .B(n1646), .Z(n1645) );
  XOR U2469 ( .A(B[25]), .B(B[24]), .Z(n1646) );
  XOR U2470 ( .A(B[258]), .B(n1647), .Z(O[259]) );
  AND U2471 ( .A(S), .B(n1648), .Z(n1647) );
  XOR U2472 ( .A(B[259]), .B(B[258]), .Z(n1648) );
  XOR U2473 ( .A(B[257]), .B(n1649), .Z(O[258]) );
  AND U2474 ( .A(S), .B(n1650), .Z(n1649) );
  XOR U2475 ( .A(B[258]), .B(B[257]), .Z(n1650) );
  XOR U2476 ( .A(B[256]), .B(n1651), .Z(O[257]) );
  AND U2477 ( .A(S), .B(n1652), .Z(n1651) );
  XOR U2478 ( .A(B[257]), .B(B[256]), .Z(n1652) );
  XOR U2479 ( .A(B[255]), .B(n1653), .Z(O[256]) );
  AND U2480 ( .A(S), .B(n1654), .Z(n1653) );
  XOR U2481 ( .A(B[256]), .B(B[255]), .Z(n1654) );
  XOR U2482 ( .A(B[254]), .B(n1655), .Z(O[255]) );
  AND U2483 ( .A(S), .B(n1656), .Z(n1655) );
  XOR U2484 ( .A(B[255]), .B(B[254]), .Z(n1656) );
  XOR U2485 ( .A(B[253]), .B(n1657), .Z(O[254]) );
  AND U2486 ( .A(S), .B(n1658), .Z(n1657) );
  XOR U2487 ( .A(B[254]), .B(B[253]), .Z(n1658) );
  XOR U2488 ( .A(B[252]), .B(n1659), .Z(O[253]) );
  AND U2489 ( .A(S), .B(n1660), .Z(n1659) );
  XOR U2490 ( .A(B[253]), .B(B[252]), .Z(n1660) );
  XOR U2491 ( .A(B[251]), .B(n1661), .Z(O[252]) );
  AND U2492 ( .A(S), .B(n1662), .Z(n1661) );
  XOR U2493 ( .A(B[252]), .B(B[251]), .Z(n1662) );
  XOR U2494 ( .A(B[250]), .B(n1663), .Z(O[251]) );
  AND U2495 ( .A(S), .B(n1664), .Z(n1663) );
  XOR U2496 ( .A(B[251]), .B(B[250]), .Z(n1664) );
  XOR U2497 ( .A(B[249]), .B(n1665), .Z(O[250]) );
  AND U2498 ( .A(S), .B(n1666), .Z(n1665) );
  XOR U2499 ( .A(B[250]), .B(B[249]), .Z(n1666) );
  XOR U2500 ( .A(B[23]), .B(n1667), .Z(O[24]) );
  AND U2501 ( .A(S), .B(n1668), .Z(n1667) );
  XOR U2502 ( .A(B[24]), .B(B[23]), .Z(n1668) );
  XOR U2503 ( .A(B[248]), .B(n1669), .Z(O[249]) );
  AND U2504 ( .A(S), .B(n1670), .Z(n1669) );
  XOR U2505 ( .A(B[249]), .B(B[248]), .Z(n1670) );
  XOR U2506 ( .A(B[247]), .B(n1671), .Z(O[248]) );
  AND U2507 ( .A(S), .B(n1672), .Z(n1671) );
  XOR U2508 ( .A(B[248]), .B(B[247]), .Z(n1672) );
  XOR U2509 ( .A(B[246]), .B(n1673), .Z(O[247]) );
  AND U2510 ( .A(S), .B(n1674), .Z(n1673) );
  XOR U2511 ( .A(B[247]), .B(B[246]), .Z(n1674) );
  XOR U2512 ( .A(B[245]), .B(n1675), .Z(O[246]) );
  AND U2513 ( .A(S), .B(n1676), .Z(n1675) );
  XOR U2514 ( .A(B[246]), .B(B[245]), .Z(n1676) );
  XOR U2515 ( .A(B[244]), .B(n1677), .Z(O[245]) );
  AND U2516 ( .A(S), .B(n1678), .Z(n1677) );
  XOR U2517 ( .A(B[245]), .B(B[244]), .Z(n1678) );
  XOR U2518 ( .A(B[243]), .B(n1679), .Z(O[244]) );
  AND U2519 ( .A(S), .B(n1680), .Z(n1679) );
  XOR U2520 ( .A(B[244]), .B(B[243]), .Z(n1680) );
  XOR U2521 ( .A(B[242]), .B(n1681), .Z(O[243]) );
  AND U2522 ( .A(S), .B(n1682), .Z(n1681) );
  XOR U2523 ( .A(B[243]), .B(B[242]), .Z(n1682) );
  XOR U2524 ( .A(B[241]), .B(n1683), .Z(O[242]) );
  AND U2525 ( .A(S), .B(n1684), .Z(n1683) );
  XOR U2526 ( .A(B[242]), .B(B[241]), .Z(n1684) );
  XOR U2527 ( .A(B[240]), .B(n1685), .Z(O[241]) );
  AND U2528 ( .A(S), .B(n1686), .Z(n1685) );
  XOR U2529 ( .A(B[241]), .B(B[240]), .Z(n1686) );
  XOR U2530 ( .A(B[239]), .B(n1687), .Z(O[240]) );
  AND U2531 ( .A(S), .B(n1688), .Z(n1687) );
  XOR U2532 ( .A(B[240]), .B(B[239]), .Z(n1688) );
  XOR U2533 ( .A(B[22]), .B(n1689), .Z(O[23]) );
  AND U2534 ( .A(S), .B(n1690), .Z(n1689) );
  XOR U2535 ( .A(B[23]), .B(B[22]), .Z(n1690) );
  XOR U2536 ( .A(B[238]), .B(n1691), .Z(O[239]) );
  AND U2537 ( .A(S), .B(n1692), .Z(n1691) );
  XOR U2538 ( .A(B[239]), .B(B[238]), .Z(n1692) );
  XOR U2539 ( .A(B[237]), .B(n1693), .Z(O[238]) );
  AND U2540 ( .A(S), .B(n1694), .Z(n1693) );
  XOR U2541 ( .A(B[238]), .B(B[237]), .Z(n1694) );
  XOR U2542 ( .A(B[236]), .B(n1695), .Z(O[237]) );
  AND U2543 ( .A(S), .B(n1696), .Z(n1695) );
  XOR U2544 ( .A(B[237]), .B(B[236]), .Z(n1696) );
  XOR U2545 ( .A(B[235]), .B(n1697), .Z(O[236]) );
  AND U2546 ( .A(S), .B(n1698), .Z(n1697) );
  XOR U2547 ( .A(B[236]), .B(B[235]), .Z(n1698) );
  XOR U2548 ( .A(B[234]), .B(n1699), .Z(O[235]) );
  AND U2549 ( .A(S), .B(n1700), .Z(n1699) );
  XOR U2550 ( .A(B[235]), .B(B[234]), .Z(n1700) );
  XOR U2551 ( .A(B[233]), .B(n1701), .Z(O[234]) );
  AND U2552 ( .A(S), .B(n1702), .Z(n1701) );
  XOR U2553 ( .A(B[234]), .B(B[233]), .Z(n1702) );
  XOR U2554 ( .A(B[232]), .B(n1703), .Z(O[233]) );
  AND U2555 ( .A(S), .B(n1704), .Z(n1703) );
  XOR U2556 ( .A(B[233]), .B(B[232]), .Z(n1704) );
  XOR U2557 ( .A(B[231]), .B(n1705), .Z(O[232]) );
  AND U2558 ( .A(S), .B(n1706), .Z(n1705) );
  XOR U2559 ( .A(B[232]), .B(B[231]), .Z(n1706) );
  XOR U2560 ( .A(B[230]), .B(n1707), .Z(O[231]) );
  AND U2561 ( .A(S), .B(n1708), .Z(n1707) );
  XOR U2562 ( .A(B[231]), .B(B[230]), .Z(n1708) );
  XOR U2563 ( .A(B[229]), .B(n1709), .Z(O[230]) );
  AND U2564 ( .A(S), .B(n1710), .Z(n1709) );
  XOR U2565 ( .A(B[230]), .B(B[229]), .Z(n1710) );
  XOR U2566 ( .A(B[21]), .B(n1711), .Z(O[22]) );
  AND U2567 ( .A(S), .B(n1712), .Z(n1711) );
  XOR U2568 ( .A(B[22]), .B(B[21]), .Z(n1712) );
  XOR U2569 ( .A(B[228]), .B(n1713), .Z(O[229]) );
  AND U2570 ( .A(S), .B(n1714), .Z(n1713) );
  XOR U2571 ( .A(B[229]), .B(B[228]), .Z(n1714) );
  XOR U2572 ( .A(B[227]), .B(n1715), .Z(O[228]) );
  AND U2573 ( .A(S), .B(n1716), .Z(n1715) );
  XOR U2574 ( .A(B[228]), .B(B[227]), .Z(n1716) );
  XOR U2575 ( .A(B[226]), .B(n1717), .Z(O[227]) );
  AND U2576 ( .A(S), .B(n1718), .Z(n1717) );
  XOR U2577 ( .A(B[227]), .B(B[226]), .Z(n1718) );
  XOR U2578 ( .A(B[225]), .B(n1719), .Z(O[226]) );
  AND U2579 ( .A(S), .B(n1720), .Z(n1719) );
  XOR U2580 ( .A(B[226]), .B(B[225]), .Z(n1720) );
  XOR U2581 ( .A(B[224]), .B(n1721), .Z(O[225]) );
  AND U2582 ( .A(S), .B(n1722), .Z(n1721) );
  XOR U2583 ( .A(B[225]), .B(B[224]), .Z(n1722) );
  XOR U2584 ( .A(B[223]), .B(n1723), .Z(O[224]) );
  AND U2585 ( .A(S), .B(n1724), .Z(n1723) );
  XOR U2586 ( .A(B[224]), .B(B[223]), .Z(n1724) );
  XOR U2587 ( .A(B[222]), .B(n1725), .Z(O[223]) );
  AND U2588 ( .A(S), .B(n1726), .Z(n1725) );
  XOR U2589 ( .A(B[223]), .B(B[222]), .Z(n1726) );
  XOR U2590 ( .A(B[221]), .B(n1727), .Z(O[222]) );
  AND U2591 ( .A(S), .B(n1728), .Z(n1727) );
  XOR U2592 ( .A(B[222]), .B(B[221]), .Z(n1728) );
  XOR U2593 ( .A(B[220]), .B(n1729), .Z(O[221]) );
  AND U2594 ( .A(S), .B(n1730), .Z(n1729) );
  XOR U2595 ( .A(B[221]), .B(B[220]), .Z(n1730) );
  XOR U2596 ( .A(B[219]), .B(n1731), .Z(O[220]) );
  AND U2597 ( .A(S), .B(n1732), .Z(n1731) );
  XOR U2598 ( .A(B[220]), .B(B[219]), .Z(n1732) );
  XOR U2599 ( .A(B[20]), .B(n1733), .Z(O[21]) );
  AND U2600 ( .A(S), .B(n1734), .Z(n1733) );
  XOR U2601 ( .A(B[21]), .B(B[20]), .Z(n1734) );
  XOR U2602 ( .A(B[218]), .B(n1735), .Z(O[219]) );
  AND U2603 ( .A(S), .B(n1736), .Z(n1735) );
  XOR U2604 ( .A(B[219]), .B(B[218]), .Z(n1736) );
  XOR U2605 ( .A(B[217]), .B(n1737), .Z(O[218]) );
  AND U2606 ( .A(S), .B(n1738), .Z(n1737) );
  XOR U2607 ( .A(B[218]), .B(B[217]), .Z(n1738) );
  XOR U2608 ( .A(B[216]), .B(n1739), .Z(O[217]) );
  AND U2609 ( .A(S), .B(n1740), .Z(n1739) );
  XOR U2610 ( .A(B[217]), .B(B[216]), .Z(n1740) );
  XOR U2611 ( .A(B[215]), .B(n1741), .Z(O[216]) );
  AND U2612 ( .A(S), .B(n1742), .Z(n1741) );
  XOR U2613 ( .A(B[216]), .B(B[215]), .Z(n1742) );
  XOR U2614 ( .A(B[214]), .B(n1743), .Z(O[215]) );
  AND U2615 ( .A(S), .B(n1744), .Z(n1743) );
  XOR U2616 ( .A(B[215]), .B(B[214]), .Z(n1744) );
  XOR U2617 ( .A(B[213]), .B(n1745), .Z(O[214]) );
  AND U2618 ( .A(S), .B(n1746), .Z(n1745) );
  XOR U2619 ( .A(B[214]), .B(B[213]), .Z(n1746) );
  XOR U2620 ( .A(B[212]), .B(n1747), .Z(O[213]) );
  AND U2621 ( .A(S), .B(n1748), .Z(n1747) );
  XOR U2622 ( .A(B[213]), .B(B[212]), .Z(n1748) );
  XOR U2623 ( .A(B[211]), .B(n1749), .Z(O[212]) );
  AND U2624 ( .A(S), .B(n1750), .Z(n1749) );
  XOR U2625 ( .A(B[212]), .B(B[211]), .Z(n1750) );
  XOR U2626 ( .A(B[210]), .B(n1751), .Z(O[211]) );
  AND U2627 ( .A(S), .B(n1752), .Z(n1751) );
  XOR U2628 ( .A(B[211]), .B(B[210]), .Z(n1752) );
  XOR U2629 ( .A(B[209]), .B(n1753), .Z(O[210]) );
  AND U2630 ( .A(S), .B(n1754), .Z(n1753) );
  XOR U2631 ( .A(B[210]), .B(B[209]), .Z(n1754) );
  XOR U2632 ( .A(B[19]), .B(n1755), .Z(O[20]) );
  AND U2633 ( .A(S), .B(n1756), .Z(n1755) );
  XOR U2634 ( .A(B[20]), .B(B[19]), .Z(n1756) );
  XOR U2635 ( .A(B[208]), .B(n1757), .Z(O[209]) );
  AND U2636 ( .A(S), .B(n1758), .Z(n1757) );
  XOR U2637 ( .A(B[209]), .B(B[208]), .Z(n1758) );
  XOR U2638 ( .A(B[207]), .B(n1759), .Z(O[208]) );
  AND U2639 ( .A(S), .B(n1760), .Z(n1759) );
  XOR U2640 ( .A(B[208]), .B(B[207]), .Z(n1760) );
  XOR U2641 ( .A(B[206]), .B(n1761), .Z(O[207]) );
  AND U2642 ( .A(S), .B(n1762), .Z(n1761) );
  XOR U2643 ( .A(B[207]), .B(B[206]), .Z(n1762) );
  XOR U2644 ( .A(B[205]), .B(n1763), .Z(O[206]) );
  AND U2645 ( .A(S), .B(n1764), .Z(n1763) );
  XOR U2646 ( .A(B[206]), .B(B[205]), .Z(n1764) );
  XOR U2647 ( .A(B[204]), .B(n1765), .Z(O[205]) );
  AND U2648 ( .A(S), .B(n1766), .Z(n1765) );
  XOR U2649 ( .A(B[205]), .B(B[204]), .Z(n1766) );
  XOR U2650 ( .A(B[203]), .B(n1767), .Z(O[204]) );
  AND U2651 ( .A(S), .B(n1768), .Z(n1767) );
  XOR U2652 ( .A(B[204]), .B(B[203]), .Z(n1768) );
  XOR U2653 ( .A(B[202]), .B(n1769), .Z(O[203]) );
  AND U2654 ( .A(S), .B(n1770), .Z(n1769) );
  XOR U2655 ( .A(B[203]), .B(B[202]), .Z(n1770) );
  XOR U2656 ( .A(B[201]), .B(n1771), .Z(O[202]) );
  AND U2657 ( .A(S), .B(n1772), .Z(n1771) );
  XOR U2658 ( .A(B[202]), .B(B[201]), .Z(n1772) );
  XOR U2659 ( .A(B[200]), .B(n1773), .Z(O[201]) );
  AND U2660 ( .A(S), .B(n1774), .Z(n1773) );
  XOR U2661 ( .A(B[201]), .B(B[200]), .Z(n1774) );
  XOR U2662 ( .A(B[199]), .B(n1775), .Z(O[200]) );
  AND U2663 ( .A(S), .B(n1776), .Z(n1775) );
  XOR U2664 ( .A(B[200]), .B(B[199]), .Z(n1776) );
  XOR U2665 ( .A(B[0]), .B(n1777), .Z(O[1]) );
  AND U2666 ( .A(S), .B(n1778), .Z(n1777) );
  XOR U2667 ( .A(B[1]), .B(B[0]), .Z(n1778) );
  XOR U2668 ( .A(B[18]), .B(n1779), .Z(O[19]) );
  AND U2669 ( .A(S), .B(n1780), .Z(n1779) );
  XOR U2670 ( .A(B[19]), .B(B[18]), .Z(n1780) );
  XOR U2671 ( .A(B[198]), .B(n1781), .Z(O[199]) );
  AND U2672 ( .A(S), .B(n1782), .Z(n1781) );
  XOR U2673 ( .A(B[199]), .B(B[198]), .Z(n1782) );
  XOR U2674 ( .A(B[197]), .B(n1783), .Z(O[198]) );
  AND U2675 ( .A(S), .B(n1784), .Z(n1783) );
  XOR U2676 ( .A(B[198]), .B(B[197]), .Z(n1784) );
  XOR U2677 ( .A(B[196]), .B(n1785), .Z(O[197]) );
  AND U2678 ( .A(S), .B(n1786), .Z(n1785) );
  XOR U2679 ( .A(B[197]), .B(B[196]), .Z(n1786) );
  XOR U2680 ( .A(B[195]), .B(n1787), .Z(O[196]) );
  AND U2681 ( .A(S), .B(n1788), .Z(n1787) );
  XOR U2682 ( .A(B[196]), .B(B[195]), .Z(n1788) );
  XOR U2683 ( .A(B[194]), .B(n1789), .Z(O[195]) );
  AND U2684 ( .A(S), .B(n1790), .Z(n1789) );
  XOR U2685 ( .A(B[195]), .B(B[194]), .Z(n1790) );
  XOR U2686 ( .A(B[193]), .B(n1791), .Z(O[194]) );
  AND U2687 ( .A(S), .B(n1792), .Z(n1791) );
  XOR U2688 ( .A(B[194]), .B(B[193]), .Z(n1792) );
  XOR U2689 ( .A(B[192]), .B(n1793), .Z(O[193]) );
  AND U2690 ( .A(S), .B(n1794), .Z(n1793) );
  XOR U2691 ( .A(B[193]), .B(B[192]), .Z(n1794) );
  XOR U2692 ( .A(B[191]), .B(n1795), .Z(O[192]) );
  AND U2693 ( .A(S), .B(n1796), .Z(n1795) );
  XOR U2694 ( .A(B[192]), .B(B[191]), .Z(n1796) );
  XOR U2695 ( .A(B[190]), .B(n1797), .Z(O[191]) );
  AND U2696 ( .A(S), .B(n1798), .Z(n1797) );
  XOR U2697 ( .A(B[191]), .B(B[190]), .Z(n1798) );
  XOR U2698 ( .A(B[189]), .B(n1799), .Z(O[190]) );
  AND U2699 ( .A(S), .B(n1800), .Z(n1799) );
  XOR U2700 ( .A(B[190]), .B(B[189]), .Z(n1800) );
  XOR U2701 ( .A(B[17]), .B(n1801), .Z(O[18]) );
  AND U2702 ( .A(S), .B(n1802), .Z(n1801) );
  XOR U2703 ( .A(B[18]), .B(B[17]), .Z(n1802) );
  XOR U2704 ( .A(B[188]), .B(n1803), .Z(O[189]) );
  AND U2705 ( .A(S), .B(n1804), .Z(n1803) );
  XOR U2706 ( .A(B[189]), .B(B[188]), .Z(n1804) );
  XOR U2707 ( .A(B[187]), .B(n1805), .Z(O[188]) );
  AND U2708 ( .A(S), .B(n1806), .Z(n1805) );
  XOR U2709 ( .A(B[188]), .B(B[187]), .Z(n1806) );
  XOR U2710 ( .A(B[186]), .B(n1807), .Z(O[187]) );
  AND U2711 ( .A(S), .B(n1808), .Z(n1807) );
  XOR U2712 ( .A(B[187]), .B(B[186]), .Z(n1808) );
  XOR U2713 ( .A(B[185]), .B(n1809), .Z(O[186]) );
  AND U2714 ( .A(S), .B(n1810), .Z(n1809) );
  XOR U2715 ( .A(B[186]), .B(B[185]), .Z(n1810) );
  XOR U2716 ( .A(B[184]), .B(n1811), .Z(O[185]) );
  AND U2717 ( .A(S), .B(n1812), .Z(n1811) );
  XOR U2718 ( .A(B[185]), .B(B[184]), .Z(n1812) );
  XOR U2719 ( .A(B[183]), .B(n1813), .Z(O[184]) );
  AND U2720 ( .A(S), .B(n1814), .Z(n1813) );
  XOR U2721 ( .A(B[184]), .B(B[183]), .Z(n1814) );
  XOR U2722 ( .A(B[182]), .B(n1815), .Z(O[183]) );
  AND U2723 ( .A(S), .B(n1816), .Z(n1815) );
  XOR U2724 ( .A(B[183]), .B(B[182]), .Z(n1816) );
  XOR U2725 ( .A(B[181]), .B(n1817), .Z(O[182]) );
  AND U2726 ( .A(S), .B(n1818), .Z(n1817) );
  XOR U2727 ( .A(B[182]), .B(B[181]), .Z(n1818) );
  XOR U2728 ( .A(B[180]), .B(n1819), .Z(O[181]) );
  AND U2729 ( .A(S), .B(n1820), .Z(n1819) );
  XOR U2730 ( .A(B[181]), .B(B[180]), .Z(n1820) );
  XOR U2731 ( .A(B[179]), .B(n1821), .Z(O[180]) );
  AND U2732 ( .A(S), .B(n1822), .Z(n1821) );
  XOR U2733 ( .A(B[180]), .B(B[179]), .Z(n1822) );
  XOR U2734 ( .A(B[16]), .B(n1823), .Z(O[17]) );
  AND U2735 ( .A(S), .B(n1824), .Z(n1823) );
  XOR U2736 ( .A(B[17]), .B(B[16]), .Z(n1824) );
  XOR U2737 ( .A(B[178]), .B(n1825), .Z(O[179]) );
  AND U2738 ( .A(S), .B(n1826), .Z(n1825) );
  XOR U2739 ( .A(B[179]), .B(B[178]), .Z(n1826) );
  XOR U2740 ( .A(B[177]), .B(n1827), .Z(O[178]) );
  AND U2741 ( .A(S), .B(n1828), .Z(n1827) );
  XOR U2742 ( .A(B[178]), .B(B[177]), .Z(n1828) );
  XOR U2743 ( .A(B[176]), .B(n1829), .Z(O[177]) );
  AND U2744 ( .A(S), .B(n1830), .Z(n1829) );
  XOR U2745 ( .A(B[177]), .B(B[176]), .Z(n1830) );
  XOR U2746 ( .A(B[175]), .B(n1831), .Z(O[176]) );
  AND U2747 ( .A(S), .B(n1832), .Z(n1831) );
  XOR U2748 ( .A(B[176]), .B(B[175]), .Z(n1832) );
  XOR U2749 ( .A(B[174]), .B(n1833), .Z(O[175]) );
  AND U2750 ( .A(S), .B(n1834), .Z(n1833) );
  XOR U2751 ( .A(B[175]), .B(B[174]), .Z(n1834) );
  XOR U2752 ( .A(B[173]), .B(n1835), .Z(O[174]) );
  AND U2753 ( .A(S), .B(n1836), .Z(n1835) );
  XOR U2754 ( .A(B[174]), .B(B[173]), .Z(n1836) );
  XOR U2755 ( .A(B[172]), .B(n1837), .Z(O[173]) );
  AND U2756 ( .A(S), .B(n1838), .Z(n1837) );
  XOR U2757 ( .A(B[173]), .B(B[172]), .Z(n1838) );
  XOR U2758 ( .A(B[171]), .B(n1839), .Z(O[172]) );
  AND U2759 ( .A(S), .B(n1840), .Z(n1839) );
  XOR U2760 ( .A(B[172]), .B(B[171]), .Z(n1840) );
  XOR U2761 ( .A(B[170]), .B(n1841), .Z(O[171]) );
  AND U2762 ( .A(S), .B(n1842), .Z(n1841) );
  XOR U2763 ( .A(B[171]), .B(B[170]), .Z(n1842) );
  XOR U2764 ( .A(B[169]), .B(n1843), .Z(O[170]) );
  AND U2765 ( .A(S), .B(n1844), .Z(n1843) );
  XOR U2766 ( .A(B[170]), .B(B[169]), .Z(n1844) );
  XOR U2767 ( .A(B[15]), .B(n1845), .Z(O[16]) );
  AND U2768 ( .A(S), .B(n1846), .Z(n1845) );
  XOR U2769 ( .A(B[16]), .B(B[15]), .Z(n1846) );
  XOR U2770 ( .A(B[168]), .B(n1847), .Z(O[169]) );
  AND U2771 ( .A(S), .B(n1848), .Z(n1847) );
  XOR U2772 ( .A(B[169]), .B(B[168]), .Z(n1848) );
  XOR U2773 ( .A(B[167]), .B(n1849), .Z(O[168]) );
  AND U2774 ( .A(S), .B(n1850), .Z(n1849) );
  XOR U2775 ( .A(B[168]), .B(B[167]), .Z(n1850) );
  XOR U2776 ( .A(B[166]), .B(n1851), .Z(O[167]) );
  AND U2777 ( .A(S), .B(n1852), .Z(n1851) );
  XOR U2778 ( .A(B[167]), .B(B[166]), .Z(n1852) );
  XOR U2779 ( .A(B[165]), .B(n1853), .Z(O[166]) );
  AND U2780 ( .A(S), .B(n1854), .Z(n1853) );
  XOR U2781 ( .A(B[166]), .B(B[165]), .Z(n1854) );
  XOR U2782 ( .A(B[164]), .B(n1855), .Z(O[165]) );
  AND U2783 ( .A(S), .B(n1856), .Z(n1855) );
  XOR U2784 ( .A(B[165]), .B(B[164]), .Z(n1856) );
  XOR U2785 ( .A(B[163]), .B(n1857), .Z(O[164]) );
  AND U2786 ( .A(S), .B(n1858), .Z(n1857) );
  XOR U2787 ( .A(B[164]), .B(B[163]), .Z(n1858) );
  XOR U2788 ( .A(B[162]), .B(n1859), .Z(O[163]) );
  AND U2789 ( .A(S), .B(n1860), .Z(n1859) );
  XOR U2790 ( .A(B[163]), .B(B[162]), .Z(n1860) );
  XOR U2791 ( .A(B[161]), .B(n1861), .Z(O[162]) );
  AND U2792 ( .A(S), .B(n1862), .Z(n1861) );
  XOR U2793 ( .A(B[162]), .B(B[161]), .Z(n1862) );
  XOR U2794 ( .A(B[160]), .B(n1863), .Z(O[161]) );
  AND U2795 ( .A(S), .B(n1864), .Z(n1863) );
  XOR U2796 ( .A(B[161]), .B(B[160]), .Z(n1864) );
  XOR U2797 ( .A(B[159]), .B(n1865), .Z(O[160]) );
  AND U2798 ( .A(S), .B(n1866), .Z(n1865) );
  XOR U2799 ( .A(B[160]), .B(B[159]), .Z(n1866) );
  XOR U2800 ( .A(B[14]), .B(n1867), .Z(O[15]) );
  AND U2801 ( .A(S), .B(n1868), .Z(n1867) );
  XOR U2802 ( .A(B[15]), .B(B[14]), .Z(n1868) );
  XOR U2803 ( .A(B[158]), .B(n1869), .Z(O[159]) );
  AND U2804 ( .A(S), .B(n1870), .Z(n1869) );
  XOR U2805 ( .A(B[159]), .B(B[158]), .Z(n1870) );
  XOR U2806 ( .A(B[157]), .B(n1871), .Z(O[158]) );
  AND U2807 ( .A(S), .B(n1872), .Z(n1871) );
  XOR U2808 ( .A(B[158]), .B(B[157]), .Z(n1872) );
  XOR U2809 ( .A(B[156]), .B(n1873), .Z(O[157]) );
  AND U2810 ( .A(S), .B(n1874), .Z(n1873) );
  XOR U2811 ( .A(B[157]), .B(B[156]), .Z(n1874) );
  XOR U2812 ( .A(B[155]), .B(n1875), .Z(O[156]) );
  AND U2813 ( .A(S), .B(n1876), .Z(n1875) );
  XOR U2814 ( .A(B[156]), .B(B[155]), .Z(n1876) );
  XOR U2815 ( .A(B[154]), .B(n1877), .Z(O[155]) );
  AND U2816 ( .A(S), .B(n1878), .Z(n1877) );
  XOR U2817 ( .A(B[155]), .B(B[154]), .Z(n1878) );
  XOR U2818 ( .A(B[153]), .B(n1879), .Z(O[154]) );
  AND U2819 ( .A(S), .B(n1880), .Z(n1879) );
  XOR U2820 ( .A(B[154]), .B(B[153]), .Z(n1880) );
  XOR U2821 ( .A(B[152]), .B(n1881), .Z(O[153]) );
  AND U2822 ( .A(S), .B(n1882), .Z(n1881) );
  XOR U2823 ( .A(B[153]), .B(B[152]), .Z(n1882) );
  XOR U2824 ( .A(B[151]), .B(n1883), .Z(O[152]) );
  AND U2825 ( .A(S), .B(n1884), .Z(n1883) );
  XOR U2826 ( .A(B[152]), .B(B[151]), .Z(n1884) );
  XOR U2827 ( .A(B[150]), .B(n1885), .Z(O[151]) );
  AND U2828 ( .A(S), .B(n1886), .Z(n1885) );
  XOR U2829 ( .A(B[151]), .B(B[150]), .Z(n1886) );
  XOR U2830 ( .A(B[149]), .B(n1887), .Z(O[150]) );
  AND U2831 ( .A(S), .B(n1888), .Z(n1887) );
  XOR U2832 ( .A(B[150]), .B(B[149]), .Z(n1888) );
  XOR U2833 ( .A(B[13]), .B(n1889), .Z(O[14]) );
  AND U2834 ( .A(S), .B(n1890), .Z(n1889) );
  XOR U2835 ( .A(B[14]), .B(B[13]), .Z(n1890) );
  XOR U2836 ( .A(B[148]), .B(n1891), .Z(O[149]) );
  AND U2837 ( .A(S), .B(n1892), .Z(n1891) );
  XOR U2838 ( .A(B[149]), .B(B[148]), .Z(n1892) );
  XOR U2839 ( .A(B[147]), .B(n1893), .Z(O[148]) );
  AND U2840 ( .A(S), .B(n1894), .Z(n1893) );
  XOR U2841 ( .A(B[148]), .B(B[147]), .Z(n1894) );
  XOR U2842 ( .A(B[146]), .B(n1895), .Z(O[147]) );
  AND U2843 ( .A(S), .B(n1896), .Z(n1895) );
  XOR U2844 ( .A(B[147]), .B(B[146]), .Z(n1896) );
  XOR U2845 ( .A(B[145]), .B(n1897), .Z(O[146]) );
  AND U2846 ( .A(S), .B(n1898), .Z(n1897) );
  XOR U2847 ( .A(B[146]), .B(B[145]), .Z(n1898) );
  XOR U2848 ( .A(B[144]), .B(n1899), .Z(O[145]) );
  AND U2849 ( .A(S), .B(n1900), .Z(n1899) );
  XOR U2850 ( .A(B[145]), .B(B[144]), .Z(n1900) );
  XOR U2851 ( .A(B[143]), .B(n1901), .Z(O[144]) );
  AND U2852 ( .A(S), .B(n1902), .Z(n1901) );
  XOR U2853 ( .A(B[144]), .B(B[143]), .Z(n1902) );
  XOR U2854 ( .A(B[142]), .B(n1903), .Z(O[143]) );
  AND U2855 ( .A(S), .B(n1904), .Z(n1903) );
  XOR U2856 ( .A(B[143]), .B(B[142]), .Z(n1904) );
  XOR U2857 ( .A(B[141]), .B(n1905), .Z(O[142]) );
  AND U2858 ( .A(S), .B(n1906), .Z(n1905) );
  XOR U2859 ( .A(B[142]), .B(B[141]), .Z(n1906) );
  XOR U2860 ( .A(B[140]), .B(n1907), .Z(O[141]) );
  AND U2861 ( .A(S), .B(n1908), .Z(n1907) );
  XOR U2862 ( .A(B[141]), .B(B[140]), .Z(n1908) );
  XOR U2863 ( .A(B[139]), .B(n1909), .Z(O[140]) );
  AND U2864 ( .A(S), .B(n1910), .Z(n1909) );
  XOR U2865 ( .A(B[140]), .B(B[139]), .Z(n1910) );
  XOR U2866 ( .A(B[12]), .B(n1911), .Z(O[13]) );
  AND U2867 ( .A(S), .B(n1912), .Z(n1911) );
  XOR U2868 ( .A(B[13]), .B(B[12]), .Z(n1912) );
  XOR U2869 ( .A(B[138]), .B(n1913), .Z(O[139]) );
  AND U2870 ( .A(S), .B(n1914), .Z(n1913) );
  XOR U2871 ( .A(B[139]), .B(B[138]), .Z(n1914) );
  XOR U2872 ( .A(B[137]), .B(n1915), .Z(O[138]) );
  AND U2873 ( .A(S), .B(n1916), .Z(n1915) );
  XOR U2874 ( .A(B[138]), .B(B[137]), .Z(n1916) );
  XOR U2875 ( .A(B[136]), .B(n1917), .Z(O[137]) );
  AND U2876 ( .A(S), .B(n1918), .Z(n1917) );
  XOR U2877 ( .A(B[137]), .B(B[136]), .Z(n1918) );
  XOR U2878 ( .A(B[135]), .B(n1919), .Z(O[136]) );
  AND U2879 ( .A(S), .B(n1920), .Z(n1919) );
  XOR U2880 ( .A(B[136]), .B(B[135]), .Z(n1920) );
  XOR U2881 ( .A(B[134]), .B(n1921), .Z(O[135]) );
  AND U2882 ( .A(S), .B(n1922), .Z(n1921) );
  XOR U2883 ( .A(B[135]), .B(B[134]), .Z(n1922) );
  XOR U2884 ( .A(B[133]), .B(n1923), .Z(O[134]) );
  AND U2885 ( .A(S), .B(n1924), .Z(n1923) );
  XOR U2886 ( .A(B[134]), .B(B[133]), .Z(n1924) );
  XOR U2887 ( .A(B[132]), .B(n1925), .Z(O[133]) );
  AND U2888 ( .A(S), .B(n1926), .Z(n1925) );
  XOR U2889 ( .A(B[133]), .B(B[132]), .Z(n1926) );
  XOR U2890 ( .A(B[131]), .B(n1927), .Z(O[132]) );
  AND U2891 ( .A(S), .B(n1928), .Z(n1927) );
  XOR U2892 ( .A(B[132]), .B(B[131]), .Z(n1928) );
  XOR U2893 ( .A(B[130]), .B(n1929), .Z(O[131]) );
  AND U2894 ( .A(S), .B(n1930), .Z(n1929) );
  XOR U2895 ( .A(B[131]), .B(B[130]), .Z(n1930) );
  XOR U2896 ( .A(B[129]), .B(n1931), .Z(O[130]) );
  AND U2897 ( .A(S), .B(n1932), .Z(n1931) );
  XOR U2898 ( .A(B[130]), .B(B[129]), .Z(n1932) );
  XOR U2899 ( .A(B[11]), .B(n1933), .Z(O[12]) );
  AND U2900 ( .A(S), .B(n1934), .Z(n1933) );
  XOR U2901 ( .A(B[12]), .B(B[11]), .Z(n1934) );
  XOR U2902 ( .A(B[128]), .B(n1935), .Z(O[129]) );
  AND U2903 ( .A(S), .B(n1936), .Z(n1935) );
  XOR U2904 ( .A(B[129]), .B(B[128]), .Z(n1936) );
  XOR U2905 ( .A(B[127]), .B(n1937), .Z(O[128]) );
  AND U2906 ( .A(S), .B(n1938), .Z(n1937) );
  XOR U2907 ( .A(B[128]), .B(B[127]), .Z(n1938) );
  XOR U2908 ( .A(B[126]), .B(n1939), .Z(O[127]) );
  AND U2909 ( .A(S), .B(n1940), .Z(n1939) );
  XOR U2910 ( .A(B[127]), .B(B[126]), .Z(n1940) );
  XOR U2911 ( .A(B[125]), .B(n1941), .Z(O[126]) );
  AND U2912 ( .A(S), .B(n1942), .Z(n1941) );
  XOR U2913 ( .A(B[126]), .B(B[125]), .Z(n1942) );
  XOR U2914 ( .A(B[124]), .B(n1943), .Z(O[125]) );
  AND U2915 ( .A(S), .B(n1944), .Z(n1943) );
  XOR U2916 ( .A(B[125]), .B(B[124]), .Z(n1944) );
  XOR U2917 ( .A(B[123]), .B(n1945), .Z(O[124]) );
  AND U2918 ( .A(S), .B(n1946), .Z(n1945) );
  XOR U2919 ( .A(B[124]), .B(B[123]), .Z(n1946) );
  XOR U2920 ( .A(B[122]), .B(n1947), .Z(O[123]) );
  AND U2921 ( .A(S), .B(n1948), .Z(n1947) );
  XOR U2922 ( .A(B[123]), .B(B[122]), .Z(n1948) );
  XOR U2923 ( .A(B[121]), .B(n1949), .Z(O[122]) );
  AND U2924 ( .A(S), .B(n1950), .Z(n1949) );
  XOR U2925 ( .A(B[122]), .B(B[121]), .Z(n1950) );
  XOR U2926 ( .A(B[120]), .B(n1951), .Z(O[121]) );
  AND U2927 ( .A(S), .B(n1952), .Z(n1951) );
  XOR U2928 ( .A(B[121]), .B(B[120]), .Z(n1952) );
  XOR U2929 ( .A(B[119]), .B(n1953), .Z(O[120]) );
  AND U2930 ( .A(S), .B(n1954), .Z(n1953) );
  XOR U2931 ( .A(B[120]), .B(B[119]), .Z(n1954) );
  XOR U2932 ( .A(B[10]), .B(n1955), .Z(O[11]) );
  AND U2933 ( .A(S), .B(n1956), .Z(n1955) );
  XOR U2934 ( .A(B[11]), .B(B[10]), .Z(n1956) );
  XOR U2935 ( .A(B[118]), .B(n1957), .Z(O[119]) );
  AND U2936 ( .A(S), .B(n1958), .Z(n1957) );
  XOR U2937 ( .A(B[119]), .B(B[118]), .Z(n1958) );
  XOR U2938 ( .A(B[117]), .B(n1959), .Z(O[118]) );
  AND U2939 ( .A(S), .B(n1960), .Z(n1959) );
  XOR U2940 ( .A(B[118]), .B(B[117]), .Z(n1960) );
  XOR U2941 ( .A(B[116]), .B(n1961), .Z(O[117]) );
  AND U2942 ( .A(S), .B(n1962), .Z(n1961) );
  XOR U2943 ( .A(B[117]), .B(B[116]), .Z(n1962) );
  XOR U2944 ( .A(B[115]), .B(n1963), .Z(O[116]) );
  AND U2945 ( .A(S), .B(n1964), .Z(n1963) );
  XOR U2946 ( .A(B[116]), .B(B[115]), .Z(n1964) );
  XOR U2947 ( .A(B[114]), .B(n1965), .Z(O[115]) );
  AND U2948 ( .A(S), .B(n1966), .Z(n1965) );
  XOR U2949 ( .A(B[115]), .B(B[114]), .Z(n1966) );
  XOR U2950 ( .A(B[113]), .B(n1967), .Z(O[114]) );
  AND U2951 ( .A(S), .B(n1968), .Z(n1967) );
  XOR U2952 ( .A(B[114]), .B(B[113]), .Z(n1968) );
  XOR U2953 ( .A(B[112]), .B(n1969), .Z(O[113]) );
  AND U2954 ( .A(S), .B(n1970), .Z(n1969) );
  XOR U2955 ( .A(B[113]), .B(B[112]), .Z(n1970) );
  XOR U2956 ( .A(B[111]), .B(n1971), .Z(O[112]) );
  AND U2957 ( .A(S), .B(n1972), .Z(n1971) );
  XOR U2958 ( .A(B[112]), .B(B[111]), .Z(n1972) );
  XOR U2959 ( .A(B[110]), .B(n1973), .Z(O[111]) );
  AND U2960 ( .A(S), .B(n1974), .Z(n1973) );
  XOR U2961 ( .A(B[111]), .B(B[110]), .Z(n1974) );
  XOR U2962 ( .A(B[109]), .B(n1975), .Z(O[110]) );
  AND U2963 ( .A(S), .B(n1976), .Z(n1975) );
  XOR U2964 ( .A(B[110]), .B(B[109]), .Z(n1976) );
  XOR U2965 ( .A(B[9]), .B(n1977), .Z(O[10]) );
  AND U2966 ( .A(S), .B(n1978), .Z(n1977) );
  XOR U2967 ( .A(B[9]), .B(B[10]), .Z(n1978) );
  XOR U2968 ( .A(B[108]), .B(n1979), .Z(O[109]) );
  AND U2969 ( .A(S), .B(n1980), .Z(n1979) );
  XOR U2970 ( .A(B[109]), .B(B[108]), .Z(n1980) );
  XOR U2971 ( .A(B[107]), .B(n1981), .Z(O[108]) );
  AND U2972 ( .A(S), .B(n1982), .Z(n1981) );
  XOR U2973 ( .A(B[108]), .B(B[107]), .Z(n1982) );
  XOR U2974 ( .A(B[106]), .B(n1983), .Z(O[107]) );
  AND U2975 ( .A(S), .B(n1984), .Z(n1983) );
  XOR U2976 ( .A(B[107]), .B(B[106]), .Z(n1984) );
  XOR U2977 ( .A(B[105]), .B(n1985), .Z(O[106]) );
  AND U2978 ( .A(S), .B(n1986), .Z(n1985) );
  XOR U2979 ( .A(B[106]), .B(B[105]), .Z(n1986) );
  XOR U2980 ( .A(B[104]), .B(n1987), .Z(O[105]) );
  AND U2981 ( .A(S), .B(n1988), .Z(n1987) );
  XOR U2982 ( .A(B[105]), .B(B[104]), .Z(n1988) );
  XOR U2983 ( .A(B[103]), .B(n1989), .Z(O[104]) );
  AND U2984 ( .A(S), .B(n1990), .Z(n1989) );
  XOR U2985 ( .A(B[104]), .B(B[103]), .Z(n1990) );
  XOR U2986 ( .A(B[102]), .B(n1991), .Z(O[103]) );
  AND U2987 ( .A(S), .B(n1992), .Z(n1991) );
  XOR U2988 ( .A(B[103]), .B(B[102]), .Z(n1992) );
  XOR U2989 ( .A(B[101]), .B(n1993), .Z(O[102]) );
  AND U2990 ( .A(S), .B(n1994), .Z(n1993) );
  XOR U2991 ( .A(B[102]), .B(B[101]), .Z(n1994) );
  XOR U2992 ( .A(B[1022]), .B(n1995), .Z(O[1023]) );
  AND U2993 ( .A(S), .B(n1996), .Z(n1995) );
  XOR U2994 ( .A(B[1023]), .B(B[1022]), .Z(n1996) );
  XOR U2995 ( .A(B[1021]), .B(n1997), .Z(O[1022]) );
  AND U2996 ( .A(S), .B(n1998), .Z(n1997) );
  XOR U2997 ( .A(B[1022]), .B(B[1021]), .Z(n1998) );
  XOR U2998 ( .A(B[1020]), .B(n1999), .Z(O[1021]) );
  AND U2999 ( .A(S), .B(n2000), .Z(n1999) );
  XOR U3000 ( .A(B[1021]), .B(B[1020]), .Z(n2000) );
  XOR U3001 ( .A(B[1019]), .B(n2001), .Z(O[1020]) );
  AND U3002 ( .A(S), .B(n2002), .Z(n2001) );
  XOR U3003 ( .A(B[1020]), .B(B[1019]), .Z(n2002) );
  XOR U3004 ( .A(B[100]), .B(n2003), .Z(O[101]) );
  AND U3005 ( .A(S), .B(n2004), .Z(n2003) );
  XOR U3006 ( .A(B[101]), .B(B[100]), .Z(n2004) );
  XOR U3007 ( .A(B[1018]), .B(n2005), .Z(O[1019]) );
  AND U3008 ( .A(S), .B(n2006), .Z(n2005) );
  XOR U3009 ( .A(B[1019]), .B(B[1018]), .Z(n2006) );
  XOR U3010 ( .A(B[1017]), .B(n2007), .Z(O[1018]) );
  AND U3011 ( .A(S), .B(n2008), .Z(n2007) );
  XOR U3012 ( .A(B[1018]), .B(B[1017]), .Z(n2008) );
  XOR U3013 ( .A(B[1016]), .B(n2009), .Z(O[1017]) );
  AND U3014 ( .A(S), .B(n2010), .Z(n2009) );
  XOR U3015 ( .A(B[1017]), .B(B[1016]), .Z(n2010) );
  XOR U3016 ( .A(B[1015]), .B(n2011), .Z(O[1016]) );
  AND U3017 ( .A(S), .B(n2012), .Z(n2011) );
  XOR U3018 ( .A(B[1016]), .B(B[1015]), .Z(n2012) );
  XOR U3019 ( .A(B[1014]), .B(n2013), .Z(O[1015]) );
  AND U3020 ( .A(S), .B(n2014), .Z(n2013) );
  XOR U3021 ( .A(B[1015]), .B(B[1014]), .Z(n2014) );
  XOR U3022 ( .A(B[1013]), .B(n2015), .Z(O[1014]) );
  AND U3023 ( .A(S), .B(n2016), .Z(n2015) );
  XOR U3024 ( .A(B[1014]), .B(B[1013]), .Z(n2016) );
  XOR U3025 ( .A(B[1012]), .B(n2017), .Z(O[1013]) );
  AND U3026 ( .A(S), .B(n2018), .Z(n2017) );
  XOR U3027 ( .A(B[1013]), .B(B[1012]), .Z(n2018) );
  XOR U3028 ( .A(B[1011]), .B(n2019), .Z(O[1012]) );
  AND U3029 ( .A(S), .B(n2020), .Z(n2019) );
  XOR U3030 ( .A(B[1012]), .B(B[1011]), .Z(n2020) );
  XOR U3031 ( .A(B[1010]), .B(n2021), .Z(O[1011]) );
  AND U3032 ( .A(S), .B(n2022), .Z(n2021) );
  XOR U3033 ( .A(B[1011]), .B(B[1010]), .Z(n2022) );
  XOR U3034 ( .A(B[1009]), .B(n2023), .Z(O[1010]) );
  AND U3035 ( .A(S), .B(n2024), .Z(n2023) );
  XOR U3036 ( .A(B[1010]), .B(B[1009]), .Z(n2024) );
  XOR U3037 ( .A(B[99]), .B(n2025), .Z(O[100]) );
  AND U3038 ( .A(S), .B(n2026), .Z(n2025) );
  XOR U3039 ( .A(B[99]), .B(B[100]), .Z(n2026) );
  XOR U3040 ( .A(B[1008]), .B(n2027), .Z(O[1009]) );
  AND U3041 ( .A(S), .B(n2028), .Z(n2027) );
  XOR U3042 ( .A(B[1009]), .B(B[1008]), .Z(n2028) );
  XOR U3043 ( .A(B[1007]), .B(n2029), .Z(O[1008]) );
  AND U3044 ( .A(S), .B(n2030), .Z(n2029) );
  XOR U3045 ( .A(B[1008]), .B(B[1007]), .Z(n2030) );
  XOR U3046 ( .A(B[1006]), .B(n2031), .Z(O[1007]) );
  AND U3047 ( .A(S), .B(n2032), .Z(n2031) );
  XOR U3048 ( .A(B[1007]), .B(B[1006]), .Z(n2032) );
  XOR U3049 ( .A(B[1005]), .B(n2033), .Z(O[1006]) );
  AND U3050 ( .A(S), .B(n2034), .Z(n2033) );
  XOR U3051 ( .A(B[1006]), .B(B[1005]), .Z(n2034) );
  XOR U3052 ( .A(B[1004]), .B(n2035), .Z(O[1005]) );
  AND U3053 ( .A(S), .B(n2036), .Z(n2035) );
  XOR U3054 ( .A(B[1005]), .B(B[1004]), .Z(n2036) );
  XOR U3055 ( .A(B[1003]), .B(n2037), .Z(O[1004]) );
  AND U3056 ( .A(S), .B(n2038), .Z(n2037) );
  XOR U3057 ( .A(B[1004]), .B(B[1003]), .Z(n2038) );
  XOR U3058 ( .A(B[1002]), .B(n2039), .Z(O[1003]) );
  AND U3059 ( .A(S), .B(n2040), .Z(n2039) );
  XOR U3060 ( .A(B[1003]), .B(B[1002]), .Z(n2040) );
  XOR U3061 ( .A(B[1001]), .B(n2041), .Z(O[1002]) );
  AND U3062 ( .A(S), .B(n2042), .Z(n2041) );
  XOR U3063 ( .A(B[1002]), .B(B[1001]), .Z(n2042) );
  XOR U3064 ( .A(B[1000]), .B(n2043), .Z(O[1001]) );
  AND U3065 ( .A(S), .B(n2044), .Z(n2043) );
  XOR U3066 ( .A(B[1001]), .B(B[1000]), .Z(n2044) );
  XOR U3067 ( .A(B[999]), .B(n2045), .Z(O[1000]) );
  AND U3068 ( .A(S), .B(n2046), .Z(n2045) );
  XOR U3069 ( .A(B[999]), .B(B[1000]), .Z(n2046) );
  AND U3070 ( .A(B[0]), .B(S), .Z(O[0]) );
endmodule


module modexp_2N_NN_N1024_CC2097152 ( clk, rst, m, e, n, c );
  input [1023:0] m;
  input [1023:0] e;
  input [1023:0] n;
  output [1023:0] c;
  input clk, rst;
  wire   _0_net_, first_one, mul_pow, n6, n8, n1033, n1034, n1035, n1036;
  wire   [1023:0] start_in;
  wire   [1023:0] ein;
  wire   [1023:0] creg_next;
  wire   [1023:0] o;
  wire   [1023:0] ereg_next;
  wire   [1023:0] y;

  MUX_N1024_0 MUX_4 ( .A(o), .B(c), .S(_0_net_), .O(creg_next) );
  MUX_N1024_2 MUX_6 ( .A({ein[1022:0], 1'b0}), .B(ein), .S(mul_pow), .O(
        ereg_next) );
  MUX_N1024_1 MUX_9 ( .A(m), .B(c), .S(mul_pow), .O(y) );
  modmult_N1024_CC1024 modmult_1 ( .clk(clk), .rst(1'b0), .start(start_in[0]), 
        .x(c), .y(y), .n(n), .o(o) );
  DFF \start_reg_reg[0]  ( .D(start_in[1023]), .CLK(clk), .RST(rst), .I(1'b1), 
        .Q(start_in[0]) );
  DFF \start_reg_reg[1]  ( .D(start_in[0]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[1]) );
  DFF \start_reg_reg[2]  ( .D(start_in[1]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[2]) );
  DFF \start_reg_reg[3]  ( .D(start_in[2]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[3]) );
  DFF \start_reg_reg[4]  ( .D(start_in[3]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[4]) );
  DFF \start_reg_reg[5]  ( .D(start_in[4]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[5]) );
  DFF \start_reg_reg[6]  ( .D(start_in[5]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[6]) );
  DFF \start_reg_reg[7]  ( .D(start_in[6]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[7]) );
  DFF \start_reg_reg[8]  ( .D(start_in[7]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[8]) );
  DFF \start_reg_reg[9]  ( .D(start_in[8]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[9]) );
  DFF \start_reg_reg[10]  ( .D(start_in[9]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[10]) );
  DFF \start_reg_reg[11]  ( .D(start_in[10]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[11]) );
  DFF \start_reg_reg[12]  ( .D(start_in[11]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[12]) );
  DFF \start_reg_reg[13]  ( .D(start_in[12]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[13]) );
  DFF \start_reg_reg[14]  ( .D(start_in[13]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[14]) );
  DFF \start_reg_reg[15]  ( .D(start_in[14]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[15]) );
  DFF \start_reg_reg[16]  ( .D(start_in[15]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[16]) );
  DFF \start_reg_reg[17]  ( .D(start_in[16]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[17]) );
  DFF \start_reg_reg[18]  ( .D(start_in[17]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[18]) );
  DFF \start_reg_reg[19]  ( .D(start_in[18]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[19]) );
  DFF \start_reg_reg[20]  ( .D(start_in[19]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[20]) );
  DFF \start_reg_reg[21]  ( .D(start_in[20]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[21]) );
  DFF \start_reg_reg[22]  ( .D(start_in[21]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[22]) );
  DFF \start_reg_reg[23]  ( .D(start_in[22]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[23]) );
  DFF \start_reg_reg[24]  ( .D(start_in[23]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[24]) );
  DFF \start_reg_reg[25]  ( .D(start_in[24]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[25]) );
  DFF \start_reg_reg[26]  ( .D(start_in[25]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[26]) );
  DFF \start_reg_reg[27]  ( .D(start_in[26]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[27]) );
  DFF \start_reg_reg[28]  ( .D(start_in[27]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[28]) );
  DFF \start_reg_reg[29]  ( .D(start_in[28]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[29]) );
  DFF \start_reg_reg[30]  ( .D(start_in[29]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[30]) );
  DFF \start_reg_reg[31]  ( .D(start_in[30]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[31]) );
  DFF \start_reg_reg[32]  ( .D(start_in[31]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[32]) );
  DFF \start_reg_reg[33]  ( .D(start_in[32]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[33]) );
  DFF \start_reg_reg[34]  ( .D(start_in[33]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[34]) );
  DFF \start_reg_reg[35]  ( .D(start_in[34]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[35]) );
  DFF \start_reg_reg[36]  ( .D(start_in[35]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[36]) );
  DFF \start_reg_reg[37]  ( .D(start_in[36]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[37]) );
  DFF \start_reg_reg[38]  ( .D(start_in[37]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[38]) );
  DFF \start_reg_reg[39]  ( .D(start_in[38]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[39]) );
  DFF \start_reg_reg[40]  ( .D(start_in[39]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[40]) );
  DFF \start_reg_reg[41]  ( .D(start_in[40]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[41]) );
  DFF \start_reg_reg[42]  ( .D(start_in[41]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[42]) );
  DFF \start_reg_reg[43]  ( .D(start_in[42]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[43]) );
  DFF \start_reg_reg[44]  ( .D(start_in[43]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[44]) );
  DFF \start_reg_reg[45]  ( .D(start_in[44]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[45]) );
  DFF \start_reg_reg[46]  ( .D(start_in[45]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[46]) );
  DFF \start_reg_reg[47]  ( .D(start_in[46]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[47]) );
  DFF \start_reg_reg[48]  ( .D(start_in[47]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[48]) );
  DFF \start_reg_reg[49]  ( .D(start_in[48]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[49]) );
  DFF \start_reg_reg[50]  ( .D(start_in[49]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[50]) );
  DFF \start_reg_reg[51]  ( .D(start_in[50]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[51]) );
  DFF \start_reg_reg[52]  ( .D(start_in[51]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[52]) );
  DFF \start_reg_reg[53]  ( .D(start_in[52]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[53]) );
  DFF \start_reg_reg[54]  ( .D(start_in[53]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[54]) );
  DFF \start_reg_reg[55]  ( .D(start_in[54]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[55]) );
  DFF \start_reg_reg[56]  ( .D(start_in[55]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[56]) );
  DFF \start_reg_reg[57]  ( .D(start_in[56]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[57]) );
  DFF \start_reg_reg[58]  ( .D(start_in[57]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[58]) );
  DFF \start_reg_reg[59]  ( .D(start_in[58]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[59]) );
  DFF \start_reg_reg[60]  ( .D(start_in[59]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[60]) );
  DFF \start_reg_reg[61]  ( .D(start_in[60]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[61]) );
  DFF \start_reg_reg[62]  ( .D(start_in[61]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[62]) );
  DFF \start_reg_reg[63]  ( .D(start_in[62]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[63]) );
  DFF \start_reg_reg[64]  ( .D(start_in[63]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[64]) );
  DFF \start_reg_reg[65]  ( .D(start_in[64]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[65]) );
  DFF \start_reg_reg[66]  ( .D(start_in[65]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[66]) );
  DFF \start_reg_reg[67]  ( .D(start_in[66]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[67]) );
  DFF \start_reg_reg[68]  ( .D(start_in[67]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[68]) );
  DFF \start_reg_reg[69]  ( .D(start_in[68]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[69]) );
  DFF \start_reg_reg[70]  ( .D(start_in[69]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[70]) );
  DFF \start_reg_reg[71]  ( .D(start_in[70]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[71]) );
  DFF \start_reg_reg[72]  ( .D(start_in[71]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[72]) );
  DFF \start_reg_reg[73]  ( .D(start_in[72]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[73]) );
  DFF \start_reg_reg[74]  ( .D(start_in[73]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[74]) );
  DFF \start_reg_reg[75]  ( .D(start_in[74]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[75]) );
  DFF \start_reg_reg[76]  ( .D(start_in[75]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[76]) );
  DFF \start_reg_reg[77]  ( .D(start_in[76]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[77]) );
  DFF \start_reg_reg[78]  ( .D(start_in[77]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[78]) );
  DFF \start_reg_reg[79]  ( .D(start_in[78]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[79]) );
  DFF \start_reg_reg[80]  ( .D(start_in[79]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[80]) );
  DFF \start_reg_reg[81]  ( .D(start_in[80]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[81]) );
  DFF \start_reg_reg[82]  ( .D(start_in[81]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[82]) );
  DFF \start_reg_reg[83]  ( .D(start_in[82]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[83]) );
  DFF \start_reg_reg[84]  ( .D(start_in[83]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[84]) );
  DFF \start_reg_reg[85]  ( .D(start_in[84]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[85]) );
  DFF \start_reg_reg[86]  ( .D(start_in[85]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[86]) );
  DFF \start_reg_reg[87]  ( .D(start_in[86]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[87]) );
  DFF \start_reg_reg[88]  ( .D(start_in[87]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[88]) );
  DFF \start_reg_reg[89]  ( .D(start_in[88]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[89]) );
  DFF \start_reg_reg[90]  ( .D(start_in[89]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[90]) );
  DFF \start_reg_reg[91]  ( .D(start_in[90]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[91]) );
  DFF \start_reg_reg[92]  ( .D(start_in[91]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[92]) );
  DFF \start_reg_reg[93]  ( .D(start_in[92]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[93]) );
  DFF \start_reg_reg[94]  ( .D(start_in[93]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[94]) );
  DFF \start_reg_reg[95]  ( .D(start_in[94]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[95]) );
  DFF \start_reg_reg[96]  ( .D(start_in[95]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[96]) );
  DFF \start_reg_reg[97]  ( .D(start_in[96]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[97]) );
  DFF \start_reg_reg[98]  ( .D(start_in[97]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[98]) );
  DFF \start_reg_reg[99]  ( .D(start_in[98]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[99]) );
  DFF \start_reg_reg[100]  ( .D(start_in[99]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[100]) );
  DFF \start_reg_reg[101]  ( .D(start_in[100]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[101]) );
  DFF \start_reg_reg[102]  ( .D(start_in[101]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[102]) );
  DFF \start_reg_reg[103]  ( .D(start_in[102]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[103]) );
  DFF \start_reg_reg[104]  ( .D(start_in[103]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[104]) );
  DFF \start_reg_reg[105]  ( .D(start_in[104]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[105]) );
  DFF \start_reg_reg[106]  ( .D(start_in[105]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[106]) );
  DFF \start_reg_reg[107]  ( .D(start_in[106]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[107]) );
  DFF \start_reg_reg[108]  ( .D(start_in[107]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[108]) );
  DFF \start_reg_reg[109]  ( .D(start_in[108]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[109]) );
  DFF \start_reg_reg[110]  ( .D(start_in[109]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[110]) );
  DFF \start_reg_reg[111]  ( .D(start_in[110]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[111]) );
  DFF \start_reg_reg[112]  ( .D(start_in[111]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[112]) );
  DFF \start_reg_reg[113]  ( .D(start_in[112]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[113]) );
  DFF \start_reg_reg[114]  ( .D(start_in[113]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[114]) );
  DFF \start_reg_reg[115]  ( .D(start_in[114]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[115]) );
  DFF \start_reg_reg[116]  ( .D(start_in[115]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[116]) );
  DFF \start_reg_reg[117]  ( .D(start_in[116]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[117]) );
  DFF \start_reg_reg[118]  ( .D(start_in[117]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[118]) );
  DFF \start_reg_reg[119]  ( .D(start_in[118]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[119]) );
  DFF \start_reg_reg[120]  ( .D(start_in[119]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[120]) );
  DFF \start_reg_reg[121]  ( .D(start_in[120]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[121]) );
  DFF \start_reg_reg[122]  ( .D(start_in[121]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[122]) );
  DFF \start_reg_reg[123]  ( .D(start_in[122]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[123]) );
  DFF \start_reg_reg[124]  ( .D(start_in[123]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[124]) );
  DFF \start_reg_reg[125]  ( .D(start_in[124]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[125]) );
  DFF \start_reg_reg[126]  ( .D(start_in[125]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[126]) );
  DFF \start_reg_reg[127]  ( .D(start_in[126]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[127]) );
  DFF \start_reg_reg[128]  ( .D(start_in[127]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[128]) );
  DFF \start_reg_reg[129]  ( .D(start_in[128]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[129]) );
  DFF \start_reg_reg[130]  ( .D(start_in[129]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[130]) );
  DFF \start_reg_reg[131]  ( .D(start_in[130]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[131]) );
  DFF \start_reg_reg[132]  ( .D(start_in[131]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[132]) );
  DFF \start_reg_reg[133]  ( .D(start_in[132]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[133]) );
  DFF \start_reg_reg[134]  ( .D(start_in[133]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[134]) );
  DFF \start_reg_reg[135]  ( .D(start_in[134]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[135]) );
  DFF \start_reg_reg[136]  ( .D(start_in[135]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[136]) );
  DFF \start_reg_reg[137]  ( .D(start_in[136]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[137]) );
  DFF \start_reg_reg[138]  ( .D(start_in[137]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[138]) );
  DFF \start_reg_reg[139]  ( .D(start_in[138]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[139]) );
  DFF \start_reg_reg[140]  ( .D(start_in[139]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[140]) );
  DFF \start_reg_reg[141]  ( .D(start_in[140]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[141]) );
  DFF \start_reg_reg[142]  ( .D(start_in[141]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[142]) );
  DFF \start_reg_reg[143]  ( .D(start_in[142]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[143]) );
  DFF \start_reg_reg[144]  ( .D(start_in[143]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[144]) );
  DFF \start_reg_reg[145]  ( .D(start_in[144]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[145]) );
  DFF \start_reg_reg[146]  ( .D(start_in[145]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[146]) );
  DFF \start_reg_reg[147]  ( .D(start_in[146]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[147]) );
  DFF \start_reg_reg[148]  ( .D(start_in[147]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[148]) );
  DFF \start_reg_reg[149]  ( .D(start_in[148]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[149]) );
  DFF \start_reg_reg[150]  ( .D(start_in[149]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[150]) );
  DFF \start_reg_reg[151]  ( .D(start_in[150]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[151]) );
  DFF \start_reg_reg[152]  ( .D(start_in[151]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[152]) );
  DFF \start_reg_reg[153]  ( .D(start_in[152]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[153]) );
  DFF \start_reg_reg[154]  ( .D(start_in[153]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[154]) );
  DFF \start_reg_reg[155]  ( .D(start_in[154]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[155]) );
  DFF \start_reg_reg[156]  ( .D(start_in[155]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[156]) );
  DFF \start_reg_reg[157]  ( .D(start_in[156]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[157]) );
  DFF \start_reg_reg[158]  ( .D(start_in[157]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[158]) );
  DFF \start_reg_reg[159]  ( .D(start_in[158]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[159]) );
  DFF \start_reg_reg[160]  ( .D(start_in[159]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[160]) );
  DFF \start_reg_reg[161]  ( .D(start_in[160]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[161]) );
  DFF \start_reg_reg[162]  ( .D(start_in[161]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[162]) );
  DFF \start_reg_reg[163]  ( .D(start_in[162]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[163]) );
  DFF \start_reg_reg[164]  ( .D(start_in[163]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[164]) );
  DFF \start_reg_reg[165]  ( .D(start_in[164]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[165]) );
  DFF \start_reg_reg[166]  ( .D(start_in[165]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[166]) );
  DFF \start_reg_reg[167]  ( .D(start_in[166]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[167]) );
  DFF \start_reg_reg[168]  ( .D(start_in[167]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[168]) );
  DFF \start_reg_reg[169]  ( .D(start_in[168]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[169]) );
  DFF \start_reg_reg[170]  ( .D(start_in[169]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[170]) );
  DFF \start_reg_reg[171]  ( .D(start_in[170]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[171]) );
  DFF \start_reg_reg[172]  ( .D(start_in[171]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[172]) );
  DFF \start_reg_reg[173]  ( .D(start_in[172]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[173]) );
  DFF \start_reg_reg[174]  ( .D(start_in[173]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[174]) );
  DFF \start_reg_reg[175]  ( .D(start_in[174]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[175]) );
  DFF \start_reg_reg[176]  ( .D(start_in[175]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[176]) );
  DFF \start_reg_reg[177]  ( .D(start_in[176]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[177]) );
  DFF \start_reg_reg[178]  ( .D(start_in[177]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[178]) );
  DFF \start_reg_reg[179]  ( .D(start_in[178]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[179]) );
  DFF \start_reg_reg[180]  ( .D(start_in[179]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[180]) );
  DFF \start_reg_reg[181]  ( .D(start_in[180]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[181]) );
  DFF \start_reg_reg[182]  ( .D(start_in[181]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[182]) );
  DFF \start_reg_reg[183]  ( .D(start_in[182]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[183]) );
  DFF \start_reg_reg[184]  ( .D(start_in[183]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[184]) );
  DFF \start_reg_reg[185]  ( .D(start_in[184]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[185]) );
  DFF \start_reg_reg[186]  ( .D(start_in[185]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[186]) );
  DFF \start_reg_reg[187]  ( .D(start_in[186]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[187]) );
  DFF \start_reg_reg[188]  ( .D(start_in[187]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[188]) );
  DFF \start_reg_reg[189]  ( .D(start_in[188]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[189]) );
  DFF \start_reg_reg[190]  ( .D(start_in[189]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[190]) );
  DFF \start_reg_reg[191]  ( .D(start_in[190]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[191]) );
  DFF \start_reg_reg[192]  ( .D(start_in[191]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[192]) );
  DFF \start_reg_reg[193]  ( .D(start_in[192]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[193]) );
  DFF \start_reg_reg[194]  ( .D(start_in[193]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[194]) );
  DFF \start_reg_reg[195]  ( .D(start_in[194]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[195]) );
  DFF \start_reg_reg[196]  ( .D(start_in[195]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[196]) );
  DFF \start_reg_reg[197]  ( .D(start_in[196]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[197]) );
  DFF \start_reg_reg[198]  ( .D(start_in[197]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[198]) );
  DFF \start_reg_reg[199]  ( .D(start_in[198]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[199]) );
  DFF \start_reg_reg[200]  ( .D(start_in[199]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[200]) );
  DFF \start_reg_reg[201]  ( .D(start_in[200]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[201]) );
  DFF \start_reg_reg[202]  ( .D(start_in[201]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[202]) );
  DFF \start_reg_reg[203]  ( .D(start_in[202]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[203]) );
  DFF \start_reg_reg[204]  ( .D(start_in[203]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[204]) );
  DFF \start_reg_reg[205]  ( .D(start_in[204]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[205]) );
  DFF \start_reg_reg[206]  ( .D(start_in[205]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[206]) );
  DFF \start_reg_reg[207]  ( .D(start_in[206]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[207]) );
  DFF \start_reg_reg[208]  ( .D(start_in[207]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[208]) );
  DFF \start_reg_reg[209]  ( .D(start_in[208]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[209]) );
  DFF \start_reg_reg[210]  ( .D(start_in[209]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[210]) );
  DFF \start_reg_reg[211]  ( .D(start_in[210]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[211]) );
  DFF \start_reg_reg[212]  ( .D(start_in[211]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[212]) );
  DFF \start_reg_reg[213]  ( .D(start_in[212]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[213]) );
  DFF \start_reg_reg[214]  ( .D(start_in[213]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[214]) );
  DFF \start_reg_reg[215]  ( .D(start_in[214]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[215]) );
  DFF \start_reg_reg[216]  ( .D(start_in[215]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[216]) );
  DFF \start_reg_reg[217]  ( .D(start_in[216]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[217]) );
  DFF \start_reg_reg[218]  ( .D(start_in[217]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[218]) );
  DFF \start_reg_reg[219]  ( .D(start_in[218]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[219]) );
  DFF \start_reg_reg[220]  ( .D(start_in[219]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[220]) );
  DFF \start_reg_reg[221]  ( .D(start_in[220]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[221]) );
  DFF \start_reg_reg[222]  ( .D(start_in[221]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[222]) );
  DFF \start_reg_reg[223]  ( .D(start_in[222]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[223]) );
  DFF \start_reg_reg[224]  ( .D(start_in[223]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[224]) );
  DFF \start_reg_reg[225]  ( .D(start_in[224]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[225]) );
  DFF \start_reg_reg[226]  ( .D(start_in[225]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[226]) );
  DFF \start_reg_reg[227]  ( .D(start_in[226]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[227]) );
  DFF \start_reg_reg[228]  ( .D(start_in[227]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[228]) );
  DFF \start_reg_reg[229]  ( .D(start_in[228]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[229]) );
  DFF \start_reg_reg[230]  ( .D(start_in[229]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[230]) );
  DFF \start_reg_reg[231]  ( .D(start_in[230]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[231]) );
  DFF \start_reg_reg[232]  ( .D(start_in[231]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[232]) );
  DFF \start_reg_reg[233]  ( .D(start_in[232]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[233]) );
  DFF \start_reg_reg[234]  ( .D(start_in[233]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[234]) );
  DFF \start_reg_reg[235]  ( .D(start_in[234]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[235]) );
  DFF \start_reg_reg[236]  ( .D(start_in[235]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[236]) );
  DFF \start_reg_reg[237]  ( .D(start_in[236]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[237]) );
  DFF \start_reg_reg[238]  ( .D(start_in[237]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[238]) );
  DFF \start_reg_reg[239]  ( .D(start_in[238]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[239]) );
  DFF \start_reg_reg[240]  ( .D(start_in[239]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[240]) );
  DFF \start_reg_reg[241]  ( .D(start_in[240]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[241]) );
  DFF \start_reg_reg[242]  ( .D(start_in[241]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[242]) );
  DFF \start_reg_reg[243]  ( .D(start_in[242]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[243]) );
  DFF \start_reg_reg[244]  ( .D(start_in[243]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[244]) );
  DFF \start_reg_reg[245]  ( .D(start_in[244]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[245]) );
  DFF \start_reg_reg[246]  ( .D(start_in[245]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[246]) );
  DFF \start_reg_reg[247]  ( .D(start_in[246]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[247]) );
  DFF \start_reg_reg[248]  ( .D(start_in[247]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[248]) );
  DFF \start_reg_reg[249]  ( .D(start_in[248]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[249]) );
  DFF \start_reg_reg[250]  ( .D(start_in[249]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[250]) );
  DFF \start_reg_reg[251]  ( .D(start_in[250]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[251]) );
  DFF \start_reg_reg[252]  ( .D(start_in[251]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[252]) );
  DFF \start_reg_reg[253]  ( .D(start_in[252]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[253]) );
  DFF \start_reg_reg[254]  ( .D(start_in[253]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[254]) );
  DFF \start_reg_reg[255]  ( .D(start_in[254]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[255]) );
  DFF \start_reg_reg[256]  ( .D(start_in[255]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[256]) );
  DFF \start_reg_reg[257]  ( .D(start_in[256]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[257]) );
  DFF \start_reg_reg[258]  ( .D(start_in[257]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[258]) );
  DFF \start_reg_reg[259]  ( .D(start_in[258]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[259]) );
  DFF \start_reg_reg[260]  ( .D(start_in[259]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[260]) );
  DFF \start_reg_reg[261]  ( .D(start_in[260]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[261]) );
  DFF \start_reg_reg[262]  ( .D(start_in[261]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[262]) );
  DFF \start_reg_reg[263]  ( .D(start_in[262]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[263]) );
  DFF \start_reg_reg[264]  ( .D(start_in[263]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[264]) );
  DFF \start_reg_reg[265]  ( .D(start_in[264]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[265]) );
  DFF \start_reg_reg[266]  ( .D(start_in[265]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[266]) );
  DFF \start_reg_reg[267]  ( .D(start_in[266]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[267]) );
  DFF \start_reg_reg[268]  ( .D(start_in[267]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[268]) );
  DFF \start_reg_reg[269]  ( .D(start_in[268]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[269]) );
  DFF \start_reg_reg[270]  ( .D(start_in[269]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[270]) );
  DFF \start_reg_reg[271]  ( .D(start_in[270]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[271]) );
  DFF \start_reg_reg[272]  ( .D(start_in[271]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[272]) );
  DFF \start_reg_reg[273]  ( .D(start_in[272]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[273]) );
  DFF \start_reg_reg[274]  ( .D(start_in[273]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[274]) );
  DFF \start_reg_reg[275]  ( .D(start_in[274]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[275]) );
  DFF \start_reg_reg[276]  ( .D(start_in[275]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[276]) );
  DFF \start_reg_reg[277]  ( .D(start_in[276]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[277]) );
  DFF \start_reg_reg[278]  ( .D(start_in[277]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[278]) );
  DFF \start_reg_reg[279]  ( .D(start_in[278]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[279]) );
  DFF \start_reg_reg[280]  ( .D(start_in[279]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[280]) );
  DFF \start_reg_reg[281]  ( .D(start_in[280]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[281]) );
  DFF \start_reg_reg[282]  ( .D(start_in[281]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[282]) );
  DFF \start_reg_reg[283]  ( .D(start_in[282]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[283]) );
  DFF \start_reg_reg[284]  ( .D(start_in[283]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[284]) );
  DFF \start_reg_reg[285]  ( .D(start_in[284]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[285]) );
  DFF \start_reg_reg[286]  ( .D(start_in[285]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[286]) );
  DFF \start_reg_reg[287]  ( .D(start_in[286]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[287]) );
  DFF \start_reg_reg[288]  ( .D(start_in[287]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[288]) );
  DFF \start_reg_reg[289]  ( .D(start_in[288]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[289]) );
  DFF \start_reg_reg[290]  ( .D(start_in[289]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[290]) );
  DFF \start_reg_reg[291]  ( .D(start_in[290]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[291]) );
  DFF \start_reg_reg[292]  ( .D(start_in[291]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[292]) );
  DFF \start_reg_reg[293]  ( .D(start_in[292]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[293]) );
  DFF \start_reg_reg[294]  ( .D(start_in[293]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[294]) );
  DFF \start_reg_reg[295]  ( .D(start_in[294]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[295]) );
  DFF \start_reg_reg[296]  ( .D(start_in[295]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[296]) );
  DFF \start_reg_reg[297]  ( .D(start_in[296]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[297]) );
  DFF \start_reg_reg[298]  ( .D(start_in[297]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[298]) );
  DFF \start_reg_reg[299]  ( .D(start_in[298]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[299]) );
  DFF \start_reg_reg[300]  ( .D(start_in[299]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[300]) );
  DFF \start_reg_reg[301]  ( .D(start_in[300]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[301]) );
  DFF \start_reg_reg[302]  ( .D(start_in[301]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[302]) );
  DFF \start_reg_reg[303]  ( .D(start_in[302]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[303]) );
  DFF \start_reg_reg[304]  ( .D(start_in[303]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[304]) );
  DFF \start_reg_reg[305]  ( .D(start_in[304]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[305]) );
  DFF \start_reg_reg[306]  ( .D(start_in[305]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[306]) );
  DFF \start_reg_reg[307]  ( .D(start_in[306]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[307]) );
  DFF \start_reg_reg[308]  ( .D(start_in[307]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[308]) );
  DFF \start_reg_reg[309]  ( .D(start_in[308]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[309]) );
  DFF \start_reg_reg[310]  ( .D(start_in[309]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[310]) );
  DFF \start_reg_reg[311]  ( .D(start_in[310]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[311]) );
  DFF \start_reg_reg[312]  ( .D(start_in[311]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[312]) );
  DFF \start_reg_reg[313]  ( .D(start_in[312]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[313]) );
  DFF \start_reg_reg[314]  ( .D(start_in[313]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[314]) );
  DFF \start_reg_reg[315]  ( .D(start_in[314]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[315]) );
  DFF \start_reg_reg[316]  ( .D(start_in[315]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[316]) );
  DFF \start_reg_reg[317]  ( .D(start_in[316]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[317]) );
  DFF \start_reg_reg[318]  ( .D(start_in[317]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[318]) );
  DFF \start_reg_reg[319]  ( .D(start_in[318]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[319]) );
  DFF \start_reg_reg[320]  ( .D(start_in[319]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[320]) );
  DFF \start_reg_reg[321]  ( .D(start_in[320]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[321]) );
  DFF \start_reg_reg[322]  ( .D(start_in[321]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[322]) );
  DFF \start_reg_reg[323]  ( .D(start_in[322]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[323]) );
  DFF \start_reg_reg[324]  ( .D(start_in[323]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[324]) );
  DFF \start_reg_reg[325]  ( .D(start_in[324]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[325]) );
  DFF \start_reg_reg[326]  ( .D(start_in[325]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[326]) );
  DFF \start_reg_reg[327]  ( .D(start_in[326]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[327]) );
  DFF \start_reg_reg[328]  ( .D(start_in[327]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[328]) );
  DFF \start_reg_reg[329]  ( .D(start_in[328]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[329]) );
  DFF \start_reg_reg[330]  ( .D(start_in[329]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[330]) );
  DFF \start_reg_reg[331]  ( .D(start_in[330]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[331]) );
  DFF \start_reg_reg[332]  ( .D(start_in[331]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[332]) );
  DFF \start_reg_reg[333]  ( .D(start_in[332]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[333]) );
  DFF \start_reg_reg[334]  ( .D(start_in[333]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[334]) );
  DFF \start_reg_reg[335]  ( .D(start_in[334]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[335]) );
  DFF \start_reg_reg[336]  ( .D(start_in[335]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[336]) );
  DFF \start_reg_reg[337]  ( .D(start_in[336]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[337]) );
  DFF \start_reg_reg[338]  ( .D(start_in[337]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[338]) );
  DFF \start_reg_reg[339]  ( .D(start_in[338]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[339]) );
  DFF \start_reg_reg[340]  ( .D(start_in[339]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[340]) );
  DFF \start_reg_reg[341]  ( .D(start_in[340]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[341]) );
  DFF \start_reg_reg[342]  ( .D(start_in[341]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[342]) );
  DFF \start_reg_reg[343]  ( .D(start_in[342]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[343]) );
  DFF \start_reg_reg[344]  ( .D(start_in[343]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[344]) );
  DFF \start_reg_reg[345]  ( .D(start_in[344]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[345]) );
  DFF \start_reg_reg[346]  ( .D(start_in[345]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[346]) );
  DFF \start_reg_reg[347]  ( .D(start_in[346]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[347]) );
  DFF \start_reg_reg[348]  ( .D(start_in[347]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[348]) );
  DFF \start_reg_reg[349]  ( .D(start_in[348]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[349]) );
  DFF \start_reg_reg[350]  ( .D(start_in[349]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[350]) );
  DFF \start_reg_reg[351]  ( .D(start_in[350]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[351]) );
  DFF \start_reg_reg[352]  ( .D(start_in[351]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[352]) );
  DFF \start_reg_reg[353]  ( .D(start_in[352]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[353]) );
  DFF \start_reg_reg[354]  ( .D(start_in[353]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[354]) );
  DFF \start_reg_reg[355]  ( .D(start_in[354]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[355]) );
  DFF \start_reg_reg[356]  ( .D(start_in[355]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[356]) );
  DFF \start_reg_reg[357]  ( .D(start_in[356]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[357]) );
  DFF \start_reg_reg[358]  ( .D(start_in[357]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[358]) );
  DFF \start_reg_reg[359]  ( .D(start_in[358]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[359]) );
  DFF \start_reg_reg[360]  ( .D(start_in[359]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[360]) );
  DFF \start_reg_reg[361]  ( .D(start_in[360]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[361]) );
  DFF \start_reg_reg[362]  ( .D(start_in[361]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[362]) );
  DFF \start_reg_reg[363]  ( .D(start_in[362]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[363]) );
  DFF \start_reg_reg[364]  ( .D(start_in[363]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[364]) );
  DFF \start_reg_reg[365]  ( .D(start_in[364]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[365]) );
  DFF \start_reg_reg[366]  ( .D(start_in[365]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[366]) );
  DFF \start_reg_reg[367]  ( .D(start_in[366]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[367]) );
  DFF \start_reg_reg[368]  ( .D(start_in[367]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[368]) );
  DFF \start_reg_reg[369]  ( .D(start_in[368]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[369]) );
  DFF \start_reg_reg[370]  ( .D(start_in[369]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[370]) );
  DFF \start_reg_reg[371]  ( .D(start_in[370]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[371]) );
  DFF \start_reg_reg[372]  ( .D(start_in[371]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[372]) );
  DFF \start_reg_reg[373]  ( .D(start_in[372]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[373]) );
  DFF \start_reg_reg[374]  ( .D(start_in[373]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[374]) );
  DFF \start_reg_reg[375]  ( .D(start_in[374]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[375]) );
  DFF \start_reg_reg[376]  ( .D(start_in[375]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[376]) );
  DFF \start_reg_reg[377]  ( .D(start_in[376]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[377]) );
  DFF \start_reg_reg[378]  ( .D(start_in[377]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[378]) );
  DFF \start_reg_reg[379]  ( .D(start_in[378]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[379]) );
  DFF \start_reg_reg[380]  ( .D(start_in[379]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[380]) );
  DFF \start_reg_reg[381]  ( .D(start_in[380]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[381]) );
  DFF \start_reg_reg[382]  ( .D(start_in[381]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[382]) );
  DFF \start_reg_reg[383]  ( .D(start_in[382]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[383]) );
  DFF \start_reg_reg[384]  ( .D(start_in[383]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[384]) );
  DFF \start_reg_reg[385]  ( .D(start_in[384]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[385]) );
  DFF \start_reg_reg[386]  ( .D(start_in[385]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[386]) );
  DFF \start_reg_reg[387]  ( .D(start_in[386]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[387]) );
  DFF \start_reg_reg[388]  ( .D(start_in[387]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[388]) );
  DFF \start_reg_reg[389]  ( .D(start_in[388]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[389]) );
  DFF \start_reg_reg[390]  ( .D(start_in[389]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[390]) );
  DFF \start_reg_reg[391]  ( .D(start_in[390]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[391]) );
  DFF \start_reg_reg[392]  ( .D(start_in[391]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[392]) );
  DFF \start_reg_reg[393]  ( .D(start_in[392]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[393]) );
  DFF \start_reg_reg[394]  ( .D(start_in[393]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[394]) );
  DFF \start_reg_reg[395]  ( .D(start_in[394]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[395]) );
  DFF \start_reg_reg[396]  ( .D(start_in[395]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[396]) );
  DFF \start_reg_reg[397]  ( .D(start_in[396]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[397]) );
  DFF \start_reg_reg[398]  ( .D(start_in[397]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[398]) );
  DFF \start_reg_reg[399]  ( .D(start_in[398]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[399]) );
  DFF \start_reg_reg[400]  ( .D(start_in[399]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[400]) );
  DFF \start_reg_reg[401]  ( .D(start_in[400]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[401]) );
  DFF \start_reg_reg[402]  ( .D(start_in[401]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[402]) );
  DFF \start_reg_reg[403]  ( .D(start_in[402]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[403]) );
  DFF \start_reg_reg[404]  ( .D(start_in[403]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[404]) );
  DFF \start_reg_reg[405]  ( .D(start_in[404]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[405]) );
  DFF \start_reg_reg[406]  ( .D(start_in[405]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[406]) );
  DFF \start_reg_reg[407]  ( .D(start_in[406]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[407]) );
  DFF \start_reg_reg[408]  ( .D(start_in[407]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[408]) );
  DFF \start_reg_reg[409]  ( .D(start_in[408]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[409]) );
  DFF \start_reg_reg[410]  ( .D(start_in[409]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[410]) );
  DFF \start_reg_reg[411]  ( .D(start_in[410]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[411]) );
  DFF \start_reg_reg[412]  ( .D(start_in[411]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[412]) );
  DFF \start_reg_reg[413]  ( .D(start_in[412]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[413]) );
  DFF \start_reg_reg[414]  ( .D(start_in[413]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[414]) );
  DFF \start_reg_reg[415]  ( .D(start_in[414]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[415]) );
  DFF \start_reg_reg[416]  ( .D(start_in[415]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[416]) );
  DFF \start_reg_reg[417]  ( .D(start_in[416]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[417]) );
  DFF \start_reg_reg[418]  ( .D(start_in[417]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[418]) );
  DFF \start_reg_reg[419]  ( .D(start_in[418]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[419]) );
  DFF \start_reg_reg[420]  ( .D(start_in[419]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[420]) );
  DFF \start_reg_reg[421]  ( .D(start_in[420]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[421]) );
  DFF \start_reg_reg[422]  ( .D(start_in[421]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[422]) );
  DFF \start_reg_reg[423]  ( .D(start_in[422]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[423]) );
  DFF \start_reg_reg[424]  ( .D(start_in[423]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[424]) );
  DFF \start_reg_reg[425]  ( .D(start_in[424]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[425]) );
  DFF \start_reg_reg[426]  ( .D(start_in[425]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[426]) );
  DFF \start_reg_reg[427]  ( .D(start_in[426]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[427]) );
  DFF \start_reg_reg[428]  ( .D(start_in[427]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[428]) );
  DFF \start_reg_reg[429]  ( .D(start_in[428]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[429]) );
  DFF \start_reg_reg[430]  ( .D(start_in[429]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[430]) );
  DFF \start_reg_reg[431]  ( .D(start_in[430]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[431]) );
  DFF \start_reg_reg[432]  ( .D(start_in[431]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[432]) );
  DFF \start_reg_reg[433]  ( .D(start_in[432]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[433]) );
  DFF \start_reg_reg[434]  ( .D(start_in[433]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[434]) );
  DFF \start_reg_reg[435]  ( .D(start_in[434]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[435]) );
  DFF \start_reg_reg[436]  ( .D(start_in[435]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[436]) );
  DFF \start_reg_reg[437]  ( .D(start_in[436]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[437]) );
  DFF \start_reg_reg[438]  ( .D(start_in[437]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[438]) );
  DFF \start_reg_reg[439]  ( .D(start_in[438]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[439]) );
  DFF \start_reg_reg[440]  ( .D(start_in[439]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[440]) );
  DFF \start_reg_reg[441]  ( .D(start_in[440]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[441]) );
  DFF \start_reg_reg[442]  ( .D(start_in[441]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[442]) );
  DFF \start_reg_reg[443]  ( .D(start_in[442]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[443]) );
  DFF \start_reg_reg[444]  ( .D(start_in[443]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[444]) );
  DFF \start_reg_reg[445]  ( .D(start_in[444]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[445]) );
  DFF \start_reg_reg[446]  ( .D(start_in[445]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[446]) );
  DFF \start_reg_reg[447]  ( .D(start_in[446]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[447]) );
  DFF \start_reg_reg[448]  ( .D(start_in[447]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[448]) );
  DFF \start_reg_reg[449]  ( .D(start_in[448]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[449]) );
  DFF \start_reg_reg[450]  ( .D(start_in[449]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[450]) );
  DFF \start_reg_reg[451]  ( .D(start_in[450]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[451]) );
  DFF \start_reg_reg[452]  ( .D(start_in[451]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[452]) );
  DFF \start_reg_reg[453]  ( .D(start_in[452]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[453]) );
  DFF \start_reg_reg[454]  ( .D(start_in[453]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[454]) );
  DFF \start_reg_reg[455]  ( .D(start_in[454]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[455]) );
  DFF \start_reg_reg[456]  ( .D(start_in[455]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[456]) );
  DFF \start_reg_reg[457]  ( .D(start_in[456]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[457]) );
  DFF \start_reg_reg[458]  ( .D(start_in[457]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[458]) );
  DFF \start_reg_reg[459]  ( .D(start_in[458]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[459]) );
  DFF \start_reg_reg[460]  ( .D(start_in[459]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[460]) );
  DFF \start_reg_reg[461]  ( .D(start_in[460]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[461]) );
  DFF \start_reg_reg[462]  ( .D(start_in[461]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[462]) );
  DFF \start_reg_reg[463]  ( .D(start_in[462]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[463]) );
  DFF \start_reg_reg[464]  ( .D(start_in[463]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[464]) );
  DFF \start_reg_reg[465]  ( .D(start_in[464]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[465]) );
  DFF \start_reg_reg[466]  ( .D(start_in[465]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[466]) );
  DFF \start_reg_reg[467]  ( .D(start_in[466]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[467]) );
  DFF \start_reg_reg[468]  ( .D(start_in[467]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[468]) );
  DFF \start_reg_reg[469]  ( .D(start_in[468]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[469]) );
  DFF \start_reg_reg[470]  ( .D(start_in[469]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[470]) );
  DFF \start_reg_reg[471]  ( .D(start_in[470]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[471]) );
  DFF \start_reg_reg[472]  ( .D(start_in[471]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[472]) );
  DFF \start_reg_reg[473]  ( .D(start_in[472]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[473]) );
  DFF \start_reg_reg[474]  ( .D(start_in[473]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[474]) );
  DFF \start_reg_reg[475]  ( .D(start_in[474]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[475]) );
  DFF \start_reg_reg[476]  ( .D(start_in[475]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[476]) );
  DFF \start_reg_reg[477]  ( .D(start_in[476]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[477]) );
  DFF \start_reg_reg[478]  ( .D(start_in[477]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[478]) );
  DFF \start_reg_reg[479]  ( .D(start_in[478]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[479]) );
  DFF \start_reg_reg[480]  ( .D(start_in[479]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[480]) );
  DFF \start_reg_reg[481]  ( .D(start_in[480]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[481]) );
  DFF \start_reg_reg[482]  ( .D(start_in[481]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[482]) );
  DFF \start_reg_reg[483]  ( .D(start_in[482]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[483]) );
  DFF \start_reg_reg[484]  ( .D(start_in[483]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[484]) );
  DFF \start_reg_reg[485]  ( .D(start_in[484]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[485]) );
  DFF \start_reg_reg[486]  ( .D(start_in[485]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[486]) );
  DFF \start_reg_reg[487]  ( .D(start_in[486]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[487]) );
  DFF \start_reg_reg[488]  ( .D(start_in[487]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[488]) );
  DFF \start_reg_reg[489]  ( .D(start_in[488]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[489]) );
  DFF \start_reg_reg[490]  ( .D(start_in[489]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[490]) );
  DFF \start_reg_reg[491]  ( .D(start_in[490]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[491]) );
  DFF \start_reg_reg[492]  ( .D(start_in[491]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[492]) );
  DFF \start_reg_reg[493]  ( .D(start_in[492]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[493]) );
  DFF \start_reg_reg[494]  ( .D(start_in[493]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[494]) );
  DFF \start_reg_reg[495]  ( .D(start_in[494]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[495]) );
  DFF \start_reg_reg[496]  ( .D(start_in[495]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[496]) );
  DFF \start_reg_reg[497]  ( .D(start_in[496]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[497]) );
  DFF \start_reg_reg[498]  ( .D(start_in[497]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[498]) );
  DFF \start_reg_reg[499]  ( .D(start_in[498]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[499]) );
  DFF \start_reg_reg[500]  ( .D(start_in[499]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[500]) );
  DFF \start_reg_reg[501]  ( .D(start_in[500]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[501]) );
  DFF \start_reg_reg[502]  ( .D(start_in[501]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[502]) );
  DFF \start_reg_reg[503]  ( .D(start_in[502]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[503]) );
  DFF \start_reg_reg[504]  ( .D(start_in[503]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[504]) );
  DFF \start_reg_reg[505]  ( .D(start_in[504]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[505]) );
  DFF \start_reg_reg[506]  ( .D(start_in[505]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[506]) );
  DFF \start_reg_reg[507]  ( .D(start_in[506]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[507]) );
  DFF \start_reg_reg[508]  ( .D(start_in[507]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[508]) );
  DFF \start_reg_reg[509]  ( .D(start_in[508]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[509]) );
  DFF \start_reg_reg[510]  ( .D(start_in[509]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[510]) );
  DFF \start_reg_reg[511]  ( .D(start_in[510]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[511]) );
  DFF \start_reg_reg[512]  ( .D(start_in[511]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[512]) );
  DFF \start_reg_reg[513]  ( .D(start_in[512]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[513]) );
  DFF \start_reg_reg[514]  ( .D(start_in[513]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[514]) );
  DFF \start_reg_reg[515]  ( .D(start_in[514]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[515]) );
  DFF \start_reg_reg[516]  ( .D(start_in[515]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[516]) );
  DFF \start_reg_reg[517]  ( .D(start_in[516]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[517]) );
  DFF \start_reg_reg[518]  ( .D(start_in[517]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[518]) );
  DFF \start_reg_reg[519]  ( .D(start_in[518]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[519]) );
  DFF \start_reg_reg[520]  ( .D(start_in[519]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[520]) );
  DFF \start_reg_reg[521]  ( .D(start_in[520]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[521]) );
  DFF \start_reg_reg[522]  ( .D(start_in[521]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[522]) );
  DFF \start_reg_reg[523]  ( .D(start_in[522]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[523]) );
  DFF \start_reg_reg[524]  ( .D(start_in[523]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[524]) );
  DFF \start_reg_reg[525]  ( .D(start_in[524]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[525]) );
  DFF \start_reg_reg[526]  ( .D(start_in[525]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[526]) );
  DFF \start_reg_reg[527]  ( .D(start_in[526]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[527]) );
  DFF \start_reg_reg[528]  ( .D(start_in[527]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[528]) );
  DFF \start_reg_reg[529]  ( .D(start_in[528]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[529]) );
  DFF \start_reg_reg[530]  ( .D(start_in[529]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[530]) );
  DFF \start_reg_reg[531]  ( .D(start_in[530]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[531]) );
  DFF \start_reg_reg[532]  ( .D(start_in[531]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[532]) );
  DFF \start_reg_reg[533]  ( .D(start_in[532]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[533]) );
  DFF \start_reg_reg[534]  ( .D(start_in[533]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[534]) );
  DFF \start_reg_reg[535]  ( .D(start_in[534]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[535]) );
  DFF \start_reg_reg[536]  ( .D(start_in[535]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[536]) );
  DFF \start_reg_reg[537]  ( .D(start_in[536]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[537]) );
  DFF \start_reg_reg[538]  ( .D(start_in[537]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[538]) );
  DFF \start_reg_reg[539]  ( .D(start_in[538]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[539]) );
  DFF \start_reg_reg[540]  ( .D(start_in[539]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[540]) );
  DFF \start_reg_reg[541]  ( .D(start_in[540]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[541]) );
  DFF \start_reg_reg[542]  ( .D(start_in[541]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[542]) );
  DFF \start_reg_reg[543]  ( .D(start_in[542]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[543]) );
  DFF \start_reg_reg[544]  ( .D(start_in[543]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[544]) );
  DFF \start_reg_reg[545]  ( .D(start_in[544]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[545]) );
  DFF \start_reg_reg[546]  ( .D(start_in[545]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[546]) );
  DFF \start_reg_reg[547]  ( .D(start_in[546]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[547]) );
  DFF \start_reg_reg[548]  ( .D(start_in[547]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[548]) );
  DFF \start_reg_reg[549]  ( .D(start_in[548]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[549]) );
  DFF \start_reg_reg[550]  ( .D(start_in[549]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[550]) );
  DFF \start_reg_reg[551]  ( .D(start_in[550]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[551]) );
  DFF \start_reg_reg[552]  ( .D(start_in[551]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[552]) );
  DFF \start_reg_reg[553]  ( .D(start_in[552]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[553]) );
  DFF \start_reg_reg[554]  ( .D(start_in[553]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[554]) );
  DFF \start_reg_reg[555]  ( .D(start_in[554]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[555]) );
  DFF \start_reg_reg[556]  ( .D(start_in[555]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[556]) );
  DFF \start_reg_reg[557]  ( .D(start_in[556]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[557]) );
  DFF \start_reg_reg[558]  ( .D(start_in[557]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[558]) );
  DFF \start_reg_reg[559]  ( .D(start_in[558]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[559]) );
  DFF \start_reg_reg[560]  ( .D(start_in[559]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[560]) );
  DFF \start_reg_reg[561]  ( .D(start_in[560]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[561]) );
  DFF \start_reg_reg[562]  ( .D(start_in[561]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[562]) );
  DFF \start_reg_reg[563]  ( .D(start_in[562]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[563]) );
  DFF \start_reg_reg[564]  ( .D(start_in[563]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[564]) );
  DFF \start_reg_reg[565]  ( .D(start_in[564]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[565]) );
  DFF \start_reg_reg[566]  ( .D(start_in[565]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[566]) );
  DFF \start_reg_reg[567]  ( .D(start_in[566]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[567]) );
  DFF \start_reg_reg[568]  ( .D(start_in[567]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[568]) );
  DFF \start_reg_reg[569]  ( .D(start_in[568]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[569]) );
  DFF \start_reg_reg[570]  ( .D(start_in[569]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[570]) );
  DFF \start_reg_reg[571]  ( .D(start_in[570]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[571]) );
  DFF \start_reg_reg[572]  ( .D(start_in[571]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[572]) );
  DFF \start_reg_reg[573]  ( .D(start_in[572]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[573]) );
  DFF \start_reg_reg[574]  ( .D(start_in[573]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[574]) );
  DFF \start_reg_reg[575]  ( .D(start_in[574]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[575]) );
  DFF \start_reg_reg[576]  ( .D(start_in[575]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[576]) );
  DFF \start_reg_reg[577]  ( .D(start_in[576]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[577]) );
  DFF \start_reg_reg[578]  ( .D(start_in[577]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[578]) );
  DFF \start_reg_reg[579]  ( .D(start_in[578]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[579]) );
  DFF \start_reg_reg[580]  ( .D(start_in[579]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[580]) );
  DFF \start_reg_reg[581]  ( .D(start_in[580]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[581]) );
  DFF \start_reg_reg[582]  ( .D(start_in[581]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[582]) );
  DFF \start_reg_reg[583]  ( .D(start_in[582]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[583]) );
  DFF \start_reg_reg[584]  ( .D(start_in[583]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[584]) );
  DFF \start_reg_reg[585]  ( .D(start_in[584]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[585]) );
  DFF \start_reg_reg[586]  ( .D(start_in[585]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[586]) );
  DFF \start_reg_reg[587]  ( .D(start_in[586]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[587]) );
  DFF \start_reg_reg[588]  ( .D(start_in[587]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[588]) );
  DFF \start_reg_reg[589]  ( .D(start_in[588]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[589]) );
  DFF \start_reg_reg[590]  ( .D(start_in[589]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[590]) );
  DFF \start_reg_reg[591]  ( .D(start_in[590]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[591]) );
  DFF \start_reg_reg[592]  ( .D(start_in[591]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[592]) );
  DFF \start_reg_reg[593]  ( .D(start_in[592]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[593]) );
  DFF \start_reg_reg[594]  ( .D(start_in[593]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[594]) );
  DFF \start_reg_reg[595]  ( .D(start_in[594]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[595]) );
  DFF \start_reg_reg[596]  ( .D(start_in[595]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[596]) );
  DFF \start_reg_reg[597]  ( .D(start_in[596]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[597]) );
  DFF \start_reg_reg[598]  ( .D(start_in[597]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[598]) );
  DFF \start_reg_reg[599]  ( .D(start_in[598]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[599]) );
  DFF \start_reg_reg[600]  ( .D(start_in[599]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[600]) );
  DFF \start_reg_reg[601]  ( .D(start_in[600]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[601]) );
  DFF \start_reg_reg[602]  ( .D(start_in[601]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[602]) );
  DFF \start_reg_reg[603]  ( .D(start_in[602]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[603]) );
  DFF \start_reg_reg[604]  ( .D(start_in[603]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[604]) );
  DFF \start_reg_reg[605]  ( .D(start_in[604]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[605]) );
  DFF \start_reg_reg[606]  ( .D(start_in[605]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[606]) );
  DFF \start_reg_reg[607]  ( .D(start_in[606]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[607]) );
  DFF \start_reg_reg[608]  ( .D(start_in[607]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[608]) );
  DFF \start_reg_reg[609]  ( .D(start_in[608]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[609]) );
  DFF \start_reg_reg[610]  ( .D(start_in[609]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[610]) );
  DFF \start_reg_reg[611]  ( .D(start_in[610]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[611]) );
  DFF \start_reg_reg[612]  ( .D(start_in[611]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[612]) );
  DFF \start_reg_reg[613]  ( .D(start_in[612]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[613]) );
  DFF \start_reg_reg[614]  ( .D(start_in[613]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[614]) );
  DFF \start_reg_reg[615]  ( .D(start_in[614]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[615]) );
  DFF \start_reg_reg[616]  ( .D(start_in[615]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[616]) );
  DFF \start_reg_reg[617]  ( .D(start_in[616]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[617]) );
  DFF \start_reg_reg[618]  ( .D(start_in[617]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[618]) );
  DFF \start_reg_reg[619]  ( .D(start_in[618]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[619]) );
  DFF \start_reg_reg[620]  ( .D(start_in[619]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[620]) );
  DFF \start_reg_reg[621]  ( .D(start_in[620]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[621]) );
  DFF \start_reg_reg[622]  ( .D(start_in[621]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[622]) );
  DFF \start_reg_reg[623]  ( .D(start_in[622]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[623]) );
  DFF \start_reg_reg[624]  ( .D(start_in[623]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[624]) );
  DFF \start_reg_reg[625]  ( .D(start_in[624]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[625]) );
  DFF \start_reg_reg[626]  ( .D(start_in[625]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[626]) );
  DFF \start_reg_reg[627]  ( .D(start_in[626]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[627]) );
  DFF \start_reg_reg[628]  ( .D(start_in[627]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[628]) );
  DFF \start_reg_reg[629]  ( .D(start_in[628]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[629]) );
  DFF \start_reg_reg[630]  ( .D(start_in[629]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[630]) );
  DFF \start_reg_reg[631]  ( .D(start_in[630]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[631]) );
  DFF \start_reg_reg[632]  ( .D(start_in[631]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[632]) );
  DFF \start_reg_reg[633]  ( .D(start_in[632]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[633]) );
  DFF \start_reg_reg[634]  ( .D(start_in[633]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[634]) );
  DFF \start_reg_reg[635]  ( .D(start_in[634]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[635]) );
  DFF \start_reg_reg[636]  ( .D(start_in[635]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[636]) );
  DFF \start_reg_reg[637]  ( .D(start_in[636]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[637]) );
  DFF \start_reg_reg[638]  ( .D(start_in[637]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[638]) );
  DFF \start_reg_reg[639]  ( .D(start_in[638]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[639]) );
  DFF \start_reg_reg[640]  ( .D(start_in[639]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[640]) );
  DFF \start_reg_reg[641]  ( .D(start_in[640]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[641]) );
  DFF \start_reg_reg[642]  ( .D(start_in[641]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[642]) );
  DFF \start_reg_reg[643]  ( .D(start_in[642]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[643]) );
  DFF \start_reg_reg[644]  ( .D(start_in[643]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[644]) );
  DFF \start_reg_reg[645]  ( .D(start_in[644]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[645]) );
  DFF \start_reg_reg[646]  ( .D(start_in[645]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[646]) );
  DFF \start_reg_reg[647]  ( .D(start_in[646]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[647]) );
  DFF \start_reg_reg[648]  ( .D(start_in[647]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[648]) );
  DFF \start_reg_reg[649]  ( .D(start_in[648]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[649]) );
  DFF \start_reg_reg[650]  ( .D(start_in[649]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[650]) );
  DFF \start_reg_reg[651]  ( .D(start_in[650]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[651]) );
  DFF \start_reg_reg[652]  ( .D(start_in[651]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[652]) );
  DFF \start_reg_reg[653]  ( .D(start_in[652]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[653]) );
  DFF \start_reg_reg[654]  ( .D(start_in[653]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[654]) );
  DFF \start_reg_reg[655]  ( .D(start_in[654]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[655]) );
  DFF \start_reg_reg[656]  ( .D(start_in[655]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[656]) );
  DFF \start_reg_reg[657]  ( .D(start_in[656]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[657]) );
  DFF \start_reg_reg[658]  ( .D(start_in[657]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[658]) );
  DFF \start_reg_reg[659]  ( .D(start_in[658]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[659]) );
  DFF \start_reg_reg[660]  ( .D(start_in[659]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[660]) );
  DFF \start_reg_reg[661]  ( .D(start_in[660]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[661]) );
  DFF \start_reg_reg[662]  ( .D(start_in[661]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[662]) );
  DFF \start_reg_reg[663]  ( .D(start_in[662]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[663]) );
  DFF \start_reg_reg[664]  ( .D(start_in[663]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[664]) );
  DFF \start_reg_reg[665]  ( .D(start_in[664]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[665]) );
  DFF \start_reg_reg[666]  ( .D(start_in[665]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[666]) );
  DFF \start_reg_reg[667]  ( .D(start_in[666]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[667]) );
  DFF \start_reg_reg[668]  ( .D(start_in[667]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[668]) );
  DFF \start_reg_reg[669]  ( .D(start_in[668]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[669]) );
  DFF \start_reg_reg[670]  ( .D(start_in[669]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[670]) );
  DFF \start_reg_reg[671]  ( .D(start_in[670]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[671]) );
  DFF \start_reg_reg[672]  ( .D(start_in[671]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[672]) );
  DFF \start_reg_reg[673]  ( .D(start_in[672]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[673]) );
  DFF \start_reg_reg[674]  ( .D(start_in[673]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[674]) );
  DFF \start_reg_reg[675]  ( .D(start_in[674]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[675]) );
  DFF \start_reg_reg[676]  ( .D(start_in[675]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[676]) );
  DFF \start_reg_reg[677]  ( .D(start_in[676]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[677]) );
  DFF \start_reg_reg[678]  ( .D(start_in[677]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[678]) );
  DFF \start_reg_reg[679]  ( .D(start_in[678]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[679]) );
  DFF \start_reg_reg[680]  ( .D(start_in[679]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[680]) );
  DFF \start_reg_reg[681]  ( .D(start_in[680]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[681]) );
  DFF \start_reg_reg[682]  ( .D(start_in[681]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[682]) );
  DFF \start_reg_reg[683]  ( .D(start_in[682]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[683]) );
  DFF \start_reg_reg[684]  ( .D(start_in[683]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[684]) );
  DFF \start_reg_reg[685]  ( .D(start_in[684]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[685]) );
  DFF \start_reg_reg[686]  ( .D(start_in[685]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[686]) );
  DFF \start_reg_reg[687]  ( .D(start_in[686]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[687]) );
  DFF \start_reg_reg[688]  ( .D(start_in[687]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[688]) );
  DFF \start_reg_reg[689]  ( .D(start_in[688]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[689]) );
  DFF \start_reg_reg[690]  ( .D(start_in[689]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[690]) );
  DFF \start_reg_reg[691]  ( .D(start_in[690]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[691]) );
  DFF \start_reg_reg[692]  ( .D(start_in[691]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[692]) );
  DFF \start_reg_reg[693]  ( .D(start_in[692]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[693]) );
  DFF \start_reg_reg[694]  ( .D(start_in[693]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[694]) );
  DFF \start_reg_reg[695]  ( .D(start_in[694]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[695]) );
  DFF \start_reg_reg[696]  ( .D(start_in[695]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[696]) );
  DFF \start_reg_reg[697]  ( .D(start_in[696]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[697]) );
  DFF \start_reg_reg[698]  ( .D(start_in[697]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[698]) );
  DFF \start_reg_reg[699]  ( .D(start_in[698]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[699]) );
  DFF \start_reg_reg[700]  ( .D(start_in[699]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[700]) );
  DFF \start_reg_reg[701]  ( .D(start_in[700]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[701]) );
  DFF \start_reg_reg[702]  ( .D(start_in[701]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[702]) );
  DFF \start_reg_reg[703]  ( .D(start_in[702]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[703]) );
  DFF \start_reg_reg[704]  ( .D(start_in[703]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[704]) );
  DFF \start_reg_reg[705]  ( .D(start_in[704]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[705]) );
  DFF \start_reg_reg[706]  ( .D(start_in[705]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[706]) );
  DFF \start_reg_reg[707]  ( .D(start_in[706]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[707]) );
  DFF \start_reg_reg[708]  ( .D(start_in[707]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[708]) );
  DFF \start_reg_reg[709]  ( .D(start_in[708]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[709]) );
  DFF \start_reg_reg[710]  ( .D(start_in[709]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[710]) );
  DFF \start_reg_reg[711]  ( .D(start_in[710]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[711]) );
  DFF \start_reg_reg[712]  ( .D(start_in[711]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[712]) );
  DFF \start_reg_reg[713]  ( .D(start_in[712]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[713]) );
  DFF \start_reg_reg[714]  ( .D(start_in[713]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[714]) );
  DFF \start_reg_reg[715]  ( .D(start_in[714]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[715]) );
  DFF \start_reg_reg[716]  ( .D(start_in[715]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[716]) );
  DFF \start_reg_reg[717]  ( .D(start_in[716]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[717]) );
  DFF \start_reg_reg[718]  ( .D(start_in[717]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[718]) );
  DFF \start_reg_reg[719]  ( .D(start_in[718]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[719]) );
  DFF \start_reg_reg[720]  ( .D(start_in[719]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[720]) );
  DFF \start_reg_reg[721]  ( .D(start_in[720]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[721]) );
  DFF \start_reg_reg[722]  ( .D(start_in[721]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[722]) );
  DFF \start_reg_reg[723]  ( .D(start_in[722]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[723]) );
  DFF \start_reg_reg[724]  ( .D(start_in[723]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[724]) );
  DFF \start_reg_reg[725]  ( .D(start_in[724]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[725]) );
  DFF \start_reg_reg[726]  ( .D(start_in[725]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[726]) );
  DFF \start_reg_reg[727]  ( .D(start_in[726]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[727]) );
  DFF \start_reg_reg[728]  ( .D(start_in[727]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[728]) );
  DFF \start_reg_reg[729]  ( .D(start_in[728]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[729]) );
  DFF \start_reg_reg[730]  ( .D(start_in[729]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[730]) );
  DFF \start_reg_reg[731]  ( .D(start_in[730]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[731]) );
  DFF \start_reg_reg[732]  ( .D(start_in[731]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[732]) );
  DFF \start_reg_reg[733]  ( .D(start_in[732]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[733]) );
  DFF \start_reg_reg[734]  ( .D(start_in[733]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[734]) );
  DFF \start_reg_reg[735]  ( .D(start_in[734]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[735]) );
  DFF \start_reg_reg[736]  ( .D(start_in[735]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[736]) );
  DFF \start_reg_reg[737]  ( .D(start_in[736]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[737]) );
  DFF \start_reg_reg[738]  ( .D(start_in[737]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[738]) );
  DFF \start_reg_reg[739]  ( .D(start_in[738]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[739]) );
  DFF \start_reg_reg[740]  ( .D(start_in[739]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[740]) );
  DFF \start_reg_reg[741]  ( .D(start_in[740]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[741]) );
  DFF \start_reg_reg[742]  ( .D(start_in[741]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[742]) );
  DFF \start_reg_reg[743]  ( .D(start_in[742]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[743]) );
  DFF \start_reg_reg[744]  ( .D(start_in[743]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[744]) );
  DFF \start_reg_reg[745]  ( .D(start_in[744]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[745]) );
  DFF \start_reg_reg[746]  ( .D(start_in[745]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[746]) );
  DFF \start_reg_reg[747]  ( .D(start_in[746]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[747]) );
  DFF \start_reg_reg[748]  ( .D(start_in[747]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[748]) );
  DFF \start_reg_reg[749]  ( .D(start_in[748]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[749]) );
  DFF \start_reg_reg[750]  ( .D(start_in[749]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[750]) );
  DFF \start_reg_reg[751]  ( .D(start_in[750]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[751]) );
  DFF \start_reg_reg[752]  ( .D(start_in[751]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[752]) );
  DFF \start_reg_reg[753]  ( .D(start_in[752]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[753]) );
  DFF \start_reg_reg[754]  ( .D(start_in[753]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[754]) );
  DFF \start_reg_reg[755]  ( .D(start_in[754]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[755]) );
  DFF \start_reg_reg[756]  ( .D(start_in[755]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[756]) );
  DFF \start_reg_reg[757]  ( .D(start_in[756]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[757]) );
  DFF \start_reg_reg[758]  ( .D(start_in[757]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[758]) );
  DFF \start_reg_reg[759]  ( .D(start_in[758]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[759]) );
  DFF \start_reg_reg[760]  ( .D(start_in[759]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[760]) );
  DFF \start_reg_reg[761]  ( .D(start_in[760]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[761]) );
  DFF \start_reg_reg[762]  ( .D(start_in[761]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[762]) );
  DFF \start_reg_reg[763]  ( .D(start_in[762]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[763]) );
  DFF \start_reg_reg[764]  ( .D(start_in[763]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[764]) );
  DFF \start_reg_reg[765]  ( .D(start_in[764]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[765]) );
  DFF \start_reg_reg[766]  ( .D(start_in[765]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[766]) );
  DFF \start_reg_reg[767]  ( .D(start_in[766]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[767]) );
  DFF \start_reg_reg[768]  ( .D(start_in[767]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[768]) );
  DFF \start_reg_reg[769]  ( .D(start_in[768]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[769]) );
  DFF \start_reg_reg[770]  ( .D(start_in[769]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[770]) );
  DFF \start_reg_reg[771]  ( .D(start_in[770]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[771]) );
  DFF \start_reg_reg[772]  ( .D(start_in[771]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[772]) );
  DFF \start_reg_reg[773]  ( .D(start_in[772]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[773]) );
  DFF \start_reg_reg[774]  ( .D(start_in[773]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[774]) );
  DFF \start_reg_reg[775]  ( .D(start_in[774]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[775]) );
  DFF \start_reg_reg[776]  ( .D(start_in[775]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[776]) );
  DFF \start_reg_reg[777]  ( .D(start_in[776]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[777]) );
  DFF \start_reg_reg[778]  ( .D(start_in[777]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[778]) );
  DFF \start_reg_reg[779]  ( .D(start_in[778]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[779]) );
  DFF \start_reg_reg[780]  ( .D(start_in[779]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[780]) );
  DFF \start_reg_reg[781]  ( .D(start_in[780]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[781]) );
  DFF \start_reg_reg[782]  ( .D(start_in[781]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[782]) );
  DFF \start_reg_reg[783]  ( .D(start_in[782]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[783]) );
  DFF \start_reg_reg[784]  ( .D(start_in[783]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[784]) );
  DFF \start_reg_reg[785]  ( .D(start_in[784]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[785]) );
  DFF \start_reg_reg[786]  ( .D(start_in[785]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[786]) );
  DFF \start_reg_reg[787]  ( .D(start_in[786]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[787]) );
  DFF \start_reg_reg[788]  ( .D(start_in[787]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[788]) );
  DFF \start_reg_reg[789]  ( .D(start_in[788]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[789]) );
  DFF \start_reg_reg[790]  ( .D(start_in[789]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[790]) );
  DFF \start_reg_reg[791]  ( .D(start_in[790]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[791]) );
  DFF \start_reg_reg[792]  ( .D(start_in[791]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[792]) );
  DFF \start_reg_reg[793]  ( .D(start_in[792]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[793]) );
  DFF \start_reg_reg[794]  ( .D(start_in[793]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[794]) );
  DFF \start_reg_reg[795]  ( .D(start_in[794]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[795]) );
  DFF \start_reg_reg[796]  ( .D(start_in[795]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[796]) );
  DFF \start_reg_reg[797]  ( .D(start_in[796]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[797]) );
  DFF \start_reg_reg[798]  ( .D(start_in[797]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[798]) );
  DFF \start_reg_reg[799]  ( .D(start_in[798]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[799]) );
  DFF \start_reg_reg[800]  ( .D(start_in[799]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[800]) );
  DFF \start_reg_reg[801]  ( .D(start_in[800]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[801]) );
  DFF \start_reg_reg[802]  ( .D(start_in[801]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[802]) );
  DFF \start_reg_reg[803]  ( .D(start_in[802]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[803]) );
  DFF \start_reg_reg[804]  ( .D(start_in[803]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[804]) );
  DFF \start_reg_reg[805]  ( .D(start_in[804]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[805]) );
  DFF \start_reg_reg[806]  ( .D(start_in[805]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[806]) );
  DFF \start_reg_reg[807]  ( .D(start_in[806]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[807]) );
  DFF \start_reg_reg[808]  ( .D(start_in[807]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[808]) );
  DFF \start_reg_reg[809]  ( .D(start_in[808]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[809]) );
  DFF \start_reg_reg[810]  ( .D(start_in[809]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[810]) );
  DFF \start_reg_reg[811]  ( .D(start_in[810]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[811]) );
  DFF \start_reg_reg[812]  ( .D(start_in[811]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[812]) );
  DFF \start_reg_reg[813]  ( .D(start_in[812]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[813]) );
  DFF \start_reg_reg[814]  ( .D(start_in[813]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[814]) );
  DFF \start_reg_reg[815]  ( .D(start_in[814]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[815]) );
  DFF \start_reg_reg[816]  ( .D(start_in[815]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[816]) );
  DFF \start_reg_reg[817]  ( .D(start_in[816]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[817]) );
  DFF \start_reg_reg[818]  ( .D(start_in[817]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[818]) );
  DFF \start_reg_reg[819]  ( .D(start_in[818]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[819]) );
  DFF \start_reg_reg[820]  ( .D(start_in[819]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[820]) );
  DFF \start_reg_reg[821]  ( .D(start_in[820]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[821]) );
  DFF \start_reg_reg[822]  ( .D(start_in[821]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[822]) );
  DFF \start_reg_reg[823]  ( .D(start_in[822]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[823]) );
  DFF \start_reg_reg[824]  ( .D(start_in[823]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[824]) );
  DFF \start_reg_reg[825]  ( .D(start_in[824]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[825]) );
  DFF \start_reg_reg[826]  ( .D(start_in[825]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[826]) );
  DFF \start_reg_reg[827]  ( .D(start_in[826]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[827]) );
  DFF \start_reg_reg[828]  ( .D(start_in[827]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[828]) );
  DFF \start_reg_reg[829]  ( .D(start_in[828]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[829]) );
  DFF \start_reg_reg[830]  ( .D(start_in[829]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[830]) );
  DFF \start_reg_reg[831]  ( .D(start_in[830]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[831]) );
  DFF \start_reg_reg[832]  ( .D(start_in[831]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[832]) );
  DFF \start_reg_reg[833]  ( .D(start_in[832]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[833]) );
  DFF \start_reg_reg[834]  ( .D(start_in[833]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[834]) );
  DFF \start_reg_reg[835]  ( .D(start_in[834]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[835]) );
  DFF \start_reg_reg[836]  ( .D(start_in[835]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[836]) );
  DFF \start_reg_reg[837]  ( .D(start_in[836]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[837]) );
  DFF \start_reg_reg[838]  ( .D(start_in[837]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[838]) );
  DFF \start_reg_reg[839]  ( .D(start_in[838]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[839]) );
  DFF \start_reg_reg[840]  ( .D(start_in[839]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[840]) );
  DFF \start_reg_reg[841]  ( .D(start_in[840]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[841]) );
  DFF \start_reg_reg[842]  ( .D(start_in[841]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[842]) );
  DFF \start_reg_reg[843]  ( .D(start_in[842]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[843]) );
  DFF \start_reg_reg[844]  ( .D(start_in[843]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[844]) );
  DFF \start_reg_reg[845]  ( .D(start_in[844]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[845]) );
  DFF \start_reg_reg[846]  ( .D(start_in[845]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[846]) );
  DFF \start_reg_reg[847]  ( .D(start_in[846]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[847]) );
  DFF \start_reg_reg[848]  ( .D(start_in[847]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[848]) );
  DFF \start_reg_reg[849]  ( .D(start_in[848]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[849]) );
  DFF \start_reg_reg[850]  ( .D(start_in[849]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[850]) );
  DFF \start_reg_reg[851]  ( .D(start_in[850]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[851]) );
  DFF \start_reg_reg[852]  ( .D(start_in[851]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[852]) );
  DFF \start_reg_reg[853]  ( .D(start_in[852]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[853]) );
  DFF \start_reg_reg[854]  ( .D(start_in[853]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[854]) );
  DFF \start_reg_reg[855]  ( .D(start_in[854]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[855]) );
  DFF \start_reg_reg[856]  ( .D(start_in[855]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[856]) );
  DFF \start_reg_reg[857]  ( .D(start_in[856]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[857]) );
  DFF \start_reg_reg[858]  ( .D(start_in[857]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[858]) );
  DFF \start_reg_reg[859]  ( .D(start_in[858]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[859]) );
  DFF \start_reg_reg[860]  ( .D(start_in[859]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[860]) );
  DFF \start_reg_reg[861]  ( .D(start_in[860]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[861]) );
  DFF \start_reg_reg[862]  ( .D(start_in[861]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[862]) );
  DFF \start_reg_reg[863]  ( .D(start_in[862]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[863]) );
  DFF \start_reg_reg[864]  ( .D(start_in[863]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[864]) );
  DFF \start_reg_reg[865]  ( .D(start_in[864]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[865]) );
  DFF \start_reg_reg[866]  ( .D(start_in[865]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[866]) );
  DFF \start_reg_reg[867]  ( .D(start_in[866]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[867]) );
  DFF \start_reg_reg[868]  ( .D(start_in[867]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[868]) );
  DFF \start_reg_reg[869]  ( .D(start_in[868]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[869]) );
  DFF \start_reg_reg[870]  ( .D(start_in[869]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[870]) );
  DFF \start_reg_reg[871]  ( .D(start_in[870]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[871]) );
  DFF \start_reg_reg[872]  ( .D(start_in[871]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[872]) );
  DFF \start_reg_reg[873]  ( .D(start_in[872]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[873]) );
  DFF \start_reg_reg[874]  ( .D(start_in[873]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[874]) );
  DFF \start_reg_reg[875]  ( .D(start_in[874]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[875]) );
  DFF \start_reg_reg[876]  ( .D(start_in[875]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[876]) );
  DFF \start_reg_reg[877]  ( .D(start_in[876]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[877]) );
  DFF \start_reg_reg[878]  ( .D(start_in[877]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[878]) );
  DFF \start_reg_reg[879]  ( .D(start_in[878]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[879]) );
  DFF \start_reg_reg[880]  ( .D(start_in[879]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[880]) );
  DFF \start_reg_reg[881]  ( .D(start_in[880]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[881]) );
  DFF \start_reg_reg[882]  ( .D(start_in[881]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[882]) );
  DFF \start_reg_reg[883]  ( .D(start_in[882]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[883]) );
  DFF \start_reg_reg[884]  ( .D(start_in[883]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[884]) );
  DFF \start_reg_reg[885]  ( .D(start_in[884]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[885]) );
  DFF \start_reg_reg[886]  ( .D(start_in[885]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[886]) );
  DFF \start_reg_reg[887]  ( .D(start_in[886]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[887]) );
  DFF \start_reg_reg[888]  ( .D(start_in[887]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[888]) );
  DFF \start_reg_reg[889]  ( .D(start_in[888]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[889]) );
  DFF \start_reg_reg[890]  ( .D(start_in[889]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[890]) );
  DFF \start_reg_reg[891]  ( .D(start_in[890]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[891]) );
  DFF \start_reg_reg[892]  ( .D(start_in[891]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[892]) );
  DFF \start_reg_reg[893]  ( .D(start_in[892]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[893]) );
  DFF \start_reg_reg[894]  ( .D(start_in[893]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[894]) );
  DFF \start_reg_reg[895]  ( .D(start_in[894]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[895]) );
  DFF \start_reg_reg[896]  ( .D(start_in[895]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[896]) );
  DFF \start_reg_reg[897]  ( .D(start_in[896]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[897]) );
  DFF \start_reg_reg[898]  ( .D(start_in[897]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[898]) );
  DFF \start_reg_reg[899]  ( .D(start_in[898]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[899]) );
  DFF \start_reg_reg[900]  ( .D(start_in[899]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[900]) );
  DFF \start_reg_reg[901]  ( .D(start_in[900]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[901]) );
  DFF \start_reg_reg[902]  ( .D(start_in[901]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[902]) );
  DFF \start_reg_reg[903]  ( .D(start_in[902]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[903]) );
  DFF \start_reg_reg[904]  ( .D(start_in[903]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[904]) );
  DFF \start_reg_reg[905]  ( .D(start_in[904]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[905]) );
  DFF \start_reg_reg[906]  ( .D(start_in[905]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[906]) );
  DFF \start_reg_reg[907]  ( .D(start_in[906]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[907]) );
  DFF \start_reg_reg[908]  ( .D(start_in[907]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[908]) );
  DFF \start_reg_reg[909]  ( .D(start_in[908]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[909]) );
  DFF \start_reg_reg[910]  ( .D(start_in[909]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[910]) );
  DFF \start_reg_reg[911]  ( .D(start_in[910]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[911]) );
  DFF \start_reg_reg[912]  ( .D(start_in[911]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[912]) );
  DFF \start_reg_reg[913]  ( .D(start_in[912]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[913]) );
  DFF \start_reg_reg[914]  ( .D(start_in[913]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[914]) );
  DFF \start_reg_reg[915]  ( .D(start_in[914]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[915]) );
  DFF \start_reg_reg[916]  ( .D(start_in[915]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[916]) );
  DFF \start_reg_reg[917]  ( .D(start_in[916]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[917]) );
  DFF \start_reg_reg[918]  ( .D(start_in[917]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[918]) );
  DFF \start_reg_reg[919]  ( .D(start_in[918]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[919]) );
  DFF \start_reg_reg[920]  ( .D(start_in[919]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[920]) );
  DFF \start_reg_reg[921]  ( .D(start_in[920]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[921]) );
  DFF \start_reg_reg[922]  ( .D(start_in[921]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[922]) );
  DFF \start_reg_reg[923]  ( .D(start_in[922]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[923]) );
  DFF \start_reg_reg[924]  ( .D(start_in[923]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[924]) );
  DFF \start_reg_reg[925]  ( .D(start_in[924]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[925]) );
  DFF \start_reg_reg[926]  ( .D(start_in[925]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[926]) );
  DFF \start_reg_reg[927]  ( .D(start_in[926]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[927]) );
  DFF \start_reg_reg[928]  ( .D(start_in[927]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[928]) );
  DFF \start_reg_reg[929]  ( .D(start_in[928]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[929]) );
  DFF \start_reg_reg[930]  ( .D(start_in[929]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[930]) );
  DFF \start_reg_reg[931]  ( .D(start_in[930]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[931]) );
  DFF \start_reg_reg[932]  ( .D(start_in[931]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[932]) );
  DFF \start_reg_reg[933]  ( .D(start_in[932]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[933]) );
  DFF \start_reg_reg[934]  ( .D(start_in[933]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[934]) );
  DFF \start_reg_reg[935]  ( .D(start_in[934]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[935]) );
  DFF \start_reg_reg[936]  ( .D(start_in[935]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[936]) );
  DFF \start_reg_reg[937]  ( .D(start_in[936]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[937]) );
  DFF \start_reg_reg[938]  ( .D(start_in[937]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[938]) );
  DFF \start_reg_reg[939]  ( .D(start_in[938]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[939]) );
  DFF \start_reg_reg[940]  ( .D(start_in[939]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[940]) );
  DFF \start_reg_reg[941]  ( .D(start_in[940]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[941]) );
  DFF \start_reg_reg[942]  ( .D(start_in[941]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[942]) );
  DFF \start_reg_reg[943]  ( .D(start_in[942]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[943]) );
  DFF \start_reg_reg[944]  ( .D(start_in[943]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[944]) );
  DFF \start_reg_reg[945]  ( .D(start_in[944]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[945]) );
  DFF \start_reg_reg[946]  ( .D(start_in[945]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[946]) );
  DFF \start_reg_reg[947]  ( .D(start_in[946]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[947]) );
  DFF \start_reg_reg[948]  ( .D(start_in[947]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[948]) );
  DFF \start_reg_reg[949]  ( .D(start_in[948]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[949]) );
  DFF \start_reg_reg[950]  ( .D(start_in[949]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[950]) );
  DFF \start_reg_reg[951]  ( .D(start_in[950]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[951]) );
  DFF \start_reg_reg[952]  ( .D(start_in[951]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[952]) );
  DFF \start_reg_reg[953]  ( .D(start_in[952]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[953]) );
  DFF \start_reg_reg[954]  ( .D(start_in[953]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[954]) );
  DFF \start_reg_reg[955]  ( .D(start_in[954]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[955]) );
  DFF \start_reg_reg[956]  ( .D(start_in[955]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[956]) );
  DFF \start_reg_reg[957]  ( .D(start_in[956]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[957]) );
  DFF \start_reg_reg[958]  ( .D(start_in[957]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[958]) );
  DFF \start_reg_reg[959]  ( .D(start_in[958]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[959]) );
  DFF \start_reg_reg[960]  ( .D(start_in[959]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[960]) );
  DFF \start_reg_reg[961]  ( .D(start_in[960]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[961]) );
  DFF \start_reg_reg[962]  ( .D(start_in[961]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[962]) );
  DFF \start_reg_reg[963]  ( .D(start_in[962]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[963]) );
  DFF \start_reg_reg[964]  ( .D(start_in[963]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[964]) );
  DFF \start_reg_reg[965]  ( .D(start_in[964]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[965]) );
  DFF \start_reg_reg[966]  ( .D(start_in[965]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[966]) );
  DFF \start_reg_reg[967]  ( .D(start_in[966]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[967]) );
  DFF \start_reg_reg[968]  ( .D(start_in[967]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[968]) );
  DFF \start_reg_reg[969]  ( .D(start_in[968]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[969]) );
  DFF \start_reg_reg[970]  ( .D(start_in[969]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[970]) );
  DFF \start_reg_reg[971]  ( .D(start_in[970]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[971]) );
  DFF \start_reg_reg[972]  ( .D(start_in[971]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[972]) );
  DFF \start_reg_reg[973]  ( .D(start_in[972]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[973]) );
  DFF \start_reg_reg[974]  ( .D(start_in[973]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[974]) );
  DFF \start_reg_reg[975]  ( .D(start_in[974]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[975]) );
  DFF \start_reg_reg[976]  ( .D(start_in[975]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[976]) );
  DFF \start_reg_reg[977]  ( .D(start_in[976]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[977]) );
  DFF \start_reg_reg[978]  ( .D(start_in[977]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[978]) );
  DFF \start_reg_reg[979]  ( .D(start_in[978]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[979]) );
  DFF \start_reg_reg[980]  ( .D(start_in[979]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[980]) );
  DFF \start_reg_reg[981]  ( .D(start_in[980]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[981]) );
  DFF \start_reg_reg[982]  ( .D(start_in[981]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[982]) );
  DFF \start_reg_reg[983]  ( .D(start_in[982]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[983]) );
  DFF \start_reg_reg[984]  ( .D(start_in[983]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[984]) );
  DFF \start_reg_reg[985]  ( .D(start_in[984]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[985]) );
  DFF \start_reg_reg[986]  ( .D(start_in[985]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[986]) );
  DFF \start_reg_reg[987]  ( .D(start_in[986]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[987]) );
  DFF \start_reg_reg[988]  ( .D(start_in[987]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[988]) );
  DFF \start_reg_reg[989]  ( .D(start_in[988]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[989]) );
  DFF \start_reg_reg[990]  ( .D(start_in[989]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[990]) );
  DFF \start_reg_reg[991]  ( .D(start_in[990]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[991]) );
  DFF \start_reg_reg[992]  ( .D(start_in[991]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[992]) );
  DFF \start_reg_reg[993]  ( .D(start_in[992]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[993]) );
  DFF \start_reg_reg[994]  ( .D(start_in[993]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[994]) );
  DFF \start_reg_reg[995]  ( .D(start_in[994]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[995]) );
  DFF \start_reg_reg[996]  ( .D(start_in[995]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[996]) );
  DFF \start_reg_reg[997]  ( .D(start_in[996]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[997]) );
  DFF \start_reg_reg[998]  ( .D(start_in[997]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[998]) );
  DFF \start_reg_reg[999]  ( .D(start_in[998]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[999]) );
  DFF \start_reg_reg[1000]  ( .D(start_in[999]), .CLK(clk), .RST(rst), .I(1'b0), .Q(start_in[1000]) );
  DFF \start_reg_reg[1001]  ( .D(start_in[1000]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1001]) );
  DFF \start_reg_reg[1002]  ( .D(start_in[1001]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1002]) );
  DFF \start_reg_reg[1003]  ( .D(start_in[1002]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1003]) );
  DFF \start_reg_reg[1004]  ( .D(start_in[1003]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1004]) );
  DFF \start_reg_reg[1005]  ( .D(start_in[1004]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1005]) );
  DFF \start_reg_reg[1006]  ( .D(start_in[1005]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1006]) );
  DFF \start_reg_reg[1007]  ( .D(start_in[1006]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1007]) );
  DFF \start_reg_reg[1008]  ( .D(start_in[1007]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1008]) );
  DFF \start_reg_reg[1009]  ( .D(start_in[1008]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1009]) );
  DFF \start_reg_reg[1010]  ( .D(start_in[1009]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1010]) );
  DFF \start_reg_reg[1011]  ( .D(start_in[1010]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1011]) );
  DFF \start_reg_reg[1012]  ( .D(start_in[1011]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1012]) );
  DFF \start_reg_reg[1013]  ( .D(start_in[1012]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1013]) );
  DFF \start_reg_reg[1014]  ( .D(start_in[1013]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1014]) );
  DFF \start_reg_reg[1015]  ( .D(start_in[1014]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1015]) );
  DFF \start_reg_reg[1016]  ( .D(start_in[1015]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1016]) );
  DFF \start_reg_reg[1017]  ( .D(start_in[1016]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1017]) );
  DFF \start_reg_reg[1018]  ( .D(start_in[1017]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1018]) );
  DFF \start_reg_reg[1019]  ( .D(start_in[1018]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1019]) );
  DFF \start_reg_reg[1020]  ( .D(start_in[1019]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1020]) );
  DFF \start_reg_reg[1021]  ( .D(start_in[1020]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1021]) );
  DFF \start_reg_reg[1022]  ( .D(start_in[1021]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1022]) );
  DFF \start_reg_reg[1023]  ( .D(start_in[1022]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1023]) );
  DFF mul_pow_reg ( .D(n8), .CLK(clk), .RST(rst), .I(1'b0), .Q(mul_pow) );
  DFF \ereg_reg[0]  ( .D(ereg_next[0]), .CLK(clk), .RST(rst), .I(e[0]), .Q(
        ein[0]) );
  DFF \ereg_reg[1]  ( .D(ereg_next[1]), .CLK(clk), .RST(rst), .I(e[1]), .Q(
        ein[1]) );
  DFF \ereg_reg[2]  ( .D(ereg_next[2]), .CLK(clk), .RST(rst), .I(e[2]), .Q(
        ein[2]) );
  DFF \ereg_reg[3]  ( .D(ereg_next[3]), .CLK(clk), .RST(rst), .I(e[3]), .Q(
        ein[3]) );
  DFF \ereg_reg[4]  ( .D(ereg_next[4]), .CLK(clk), .RST(rst), .I(e[4]), .Q(
        ein[4]) );
  DFF \ereg_reg[5]  ( .D(ereg_next[5]), .CLK(clk), .RST(rst), .I(e[5]), .Q(
        ein[5]) );
  DFF \ereg_reg[6]  ( .D(ereg_next[6]), .CLK(clk), .RST(rst), .I(e[6]), .Q(
        ein[6]) );
  DFF \ereg_reg[7]  ( .D(ereg_next[7]), .CLK(clk), .RST(rst), .I(e[7]), .Q(
        ein[7]) );
  DFF \ereg_reg[8]  ( .D(ereg_next[8]), .CLK(clk), .RST(rst), .I(e[8]), .Q(
        ein[8]) );
  DFF \ereg_reg[9]  ( .D(ereg_next[9]), .CLK(clk), .RST(rst), .I(e[9]), .Q(
        ein[9]) );
  DFF \ereg_reg[10]  ( .D(ereg_next[10]), .CLK(clk), .RST(rst), .I(e[10]), .Q(
        ein[10]) );
  DFF \ereg_reg[11]  ( .D(ereg_next[11]), .CLK(clk), .RST(rst), .I(e[11]), .Q(
        ein[11]) );
  DFF \ereg_reg[12]  ( .D(ereg_next[12]), .CLK(clk), .RST(rst), .I(e[12]), .Q(
        ein[12]) );
  DFF \ereg_reg[13]  ( .D(ereg_next[13]), .CLK(clk), .RST(rst), .I(e[13]), .Q(
        ein[13]) );
  DFF \ereg_reg[14]  ( .D(ereg_next[14]), .CLK(clk), .RST(rst), .I(e[14]), .Q(
        ein[14]) );
  DFF \ereg_reg[15]  ( .D(ereg_next[15]), .CLK(clk), .RST(rst), .I(e[15]), .Q(
        ein[15]) );
  DFF \ereg_reg[16]  ( .D(ereg_next[16]), .CLK(clk), .RST(rst), .I(e[16]), .Q(
        ein[16]) );
  DFF \ereg_reg[17]  ( .D(ereg_next[17]), .CLK(clk), .RST(rst), .I(e[17]), .Q(
        ein[17]) );
  DFF \ereg_reg[18]  ( .D(ereg_next[18]), .CLK(clk), .RST(rst), .I(e[18]), .Q(
        ein[18]) );
  DFF \ereg_reg[19]  ( .D(ereg_next[19]), .CLK(clk), .RST(rst), .I(e[19]), .Q(
        ein[19]) );
  DFF \ereg_reg[20]  ( .D(ereg_next[20]), .CLK(clk), .RST(rst), .I(e[20]), .Q(
        ein[20]) );
  DFF \ereg_reg[21]  ( .D(ereg_next[21]), .CLK(clk), .RST(rst), .I(e[21]), .Q(
        ein[21]) );
  DFF \ereg_reg[22]  ( .D(ereg_next[22]), .CLK(clk), .RST(rst), .I(e[22]), .Q(
        ein[22]) );
  DFF \ereg_reg[23]  ( .D(ereg_next[23]), .CLK(clk), .RST(rst), .I(e[23]), .Q(
        ein[23]) );
  DFF \ereg_reg[24]  ( .D(ereg_next[24]), .CLK(clk), .RST(rst), .I(e[24]), .Q(
        ein[24]) );
  DFF \ereg_reg[25]  ( .D(ereg_next[25]), .CLK(clk), .RST(rst), .I(e[25]), .Q(
        ein[25]) );
  DFF \ereg_reg[26]  ( .D(ereg_next[26]), .CLK(clk), .RST(rst), .I(e[26]), .Q(
        ein[26]) );
  DFF \ereg_reg[27]  ( .D(ereg_next[27]), .CLK(clk), .RST(rst), .I(e[27]), .Q(
        ein[27]) );
  DFF \ereg_reg[28]  ( .D(ereg_next[28]), .CLK(clk), .RST(rst), .I(e[28]), .Q(
        ein[28]) );
  DFF \ereg_reg[29]  ( .D(ereg_next[29]), .CLK(clk), .RST(rst), .I(e[29]), .Q(
        ein[29]) );
  DFF \ereg_reg[30]  ( .D(ereg_next[30]), .CLK(clk), .RST(rst), .I(e[30]), .Q(
        ein[30]) );
  DFF \ereg_reg[31]  ( .D(ereg_next[31]), .CLK(clk), .RST(rst), .I(e[31]), .Q(
        ein[31]) );
  DFF \ereg_reg[32]  ( .D(ereg_next[32]), .CLK(clk), .RST(rst), .I(e[32]), .Q(
        ein[32]) );
  DFF \ereg_reg[33]  ( .D(ereg_next[33]), .CLK(clk), .RST(rst), .I(e[33]), .Q(
        ein[33]) );
  DFF \ereg_reg[34]  ( .D(ereg_next[34]), .CLK(clk), .RST(rst), .I(e[34]), .Q(
        ein[34]) );
  DFF \ereg_reg[35]  ( .D(ereg_next[35]), .CLK(clk), .RST(rst), .I(e[35]), .Q(
        ein[35]) );
  DFF \ereg_reg[36]  ( .D(ereg_next[36]), .CLK(clk), .RST(rst), .I(e[36]), .Q(
        ein[36]) );
  DFF \ereg_reg[37]  ( .D(ereg_next[37]), .CLK(clk), .RST(rst), .I(e[37]), .Q(
        ein[37]) );
  DFF \ereg_reg[38]  ( .D(ereg_next[38]), .CLK(clk), .RST(rst), .I(e[38]), .Q(
        ein[38]) );
  DFF \ereg_reg[39]  ( .D(ereg_next[39]), .CLK(clk), .RST(rst), .I(e[39]), .Q(
        ein[39]) );
  DFF \ereg_reg[40]  ( .D(ereg_next[40]), .CLK(clk), .RST(rst), .I(e[40]), .Q(
        ein[40]) );
  DFF \ereg_reg[41]  ( .D(ereg_next[41]), .CLK(clk), .RST(rst), .I(e[41]), .Q(
        ein[41]) );
  DFF \ereg_reg[42]  ( .D(ereg_next[42]), .CLK(clk), .RST(rst), .I(e[42]), .Q(
        ein[42]) );
  DFF \ereg_reg[43]  ( .D(ereg_next[43]), .CLK(clk), .RST(rst), .I(e[43]), .Q(
        ein[43]) );
  DFF \ereg_reg[44]  ( .D(ereg_next[44]), .CLK(clk), .RST(rst), .I(e[44]), .Q(
        ein[44]) );
  DFF \ereg_reg[45]  ( .D(ereg_next[45]), .CLK(clk), .RST(rst), .I(e[45]), .Q(
        ein[45]) );
  DFF \ereg_reg[46]  ( .D(ereg_next[46]), .CLK(clk), .RST(rst), .I(e[46]), .Q(
        ein[46]) );
  DFF \ereg_reg[47]  ( .D(ereg_next[47]), .CLK(clk), .RST(rst), .I(e[47]), .Q(
        ein[47]) );
  DFF \ereg_reg[48]  ( .D(ereg_next[48]), .CLK(clk), .RST(rst), .I(e[48]), .Q(
        ein[48]) );
  DFF \ereg_reg[49]  ( .D(ereg_next[49]), .CLK(clk), .RST(rst), .I(e[49]), .Q(
        ein[49]) );
  DFF \ereg_reg[50]  ( .D(ereg_next[50]), .CLK(clk), .RST(rst), .I(e[50]), .Q(
        ein[50]) );
  DFF \ereg_reg[51]  ( .D(ereg_next[51]), .CLK(clk), .RST(rst), .I(e[51]), .Q(
        ein[51]) );
  DFF \ereg_reg[52]  ( .D(ereg_next[52]), .CLK(clk), .RST(rst), .I(e[52]), .Q(
        ein[52]) );
  DFF \ereg_reg[53]  ( .D(ereg_next[53]), .CLK(clk), .RST(rst), .I(e[53]), .Q(
        ein[53]) );
  DFF \ereg_reg[54]  ( .D(ereg_next[54]), .CLK(clk), .RST(rst), .I(e[54]), .Q(
        ein[54]) );
  DFF \ereg_reg[55]  ( .D(ereg_next[55]), .CLK(clk), .RST(rst), .I(e[55]), .Q(
        ein[55]) );
  DFF \ereg_reg[56]  ( .D(ereg_next[56]), .CLK(clk), .RST(rst), .I(e[56]), .Q(
        ein[56]) );
  DFF \ereg_reg[57]  ( .D(ereg_next[57]), .CLK(clk), .RST(rst), .I(e[57]), .Q(
        ein[57]) );
  DFF \ereg_reg[58]  ( .D(ereg_next[58]), .CLK(clk), .RST(rst), .I(e[58]), .Q(
        ein[58]) );
  DFF \ereg_reg[59]  ( .D(ereg_next[59]), .CLK(clk), .RST(rst), .I(e[59]), .Q(
        ein[59]) );
  DFF \ereg_reg[60]  ( .D(ereg_next[60]), .CLK(clk), .RST(rst), .I(e[60]), .Q(
        ein[60]) );
  DFF \ereg_reg[61]  ( .D(ereg_next[61]), .CLK(clk), .RST(rst), .I(e[61]), .Q(
        ein[61]) );
  DFF \ereg_reg[62]  ( .D(ereg_next[62]), .CLK(clk), .RST(rst), .I(e[62]), .Q(
        ein[62]) );
  DFF \ereg_reg[63]  ( .D(ereg_next[63]), .CLK(clk), .RST(rst), .I(e[63]), .Q(
        ein[63]) );
  DFF \ereg_reg[64]  ( .D(ereg_next[64]), .CLK(clk), .RST(rst), .I(e[64]), .Q(
        ein[64]) );
  DFF \ereg_reg[65]  ( .D(ereg_next[65]), .CLK(clk), .RST(rst), .I(e[65]), .Q(
        ein[65]) );
  DFF \ereg_reg[66]  ( .D(ereg_next[66]), .CLK(clk), .RST(rst), .I(e[66]), .Q(
        ein[66]) );
  DFF \ereg_reg[67]  ( .D(ereg_next[67]), .CLK(clk), .RST(rst), .I(e[67]), .Q(
        ein[67]) );
  DFF \ereg_reg[68]  ( .D(ereg_next[68]), .CLK(clk), .RST(rst), .I(e[68]), .Q(
        ein[68]) );
  DFF \ereg_reg[69]  ( .D(ereg_next[69]), .CLK(clk), .RST(rst), .I(e[69]), .Q(
        ein[69]) );
  DFF \ereg_reg[70]  ( .D(ereg_next[70]), .CLK(clk), .RST(rst), .I(e[70]), .Q(
        ein[70]) );
  DFF \ereg_reg[71]  ( .D(ereg_next[71]), .CLK(clk), .RST(rst), .I(e[71]), .Q(
        ein[71]) );
  DFF \ereg_reg[72]  ( .D(ereg_next[72]), .CLK(clk), .RST(rst), .I(e[72]), .Q(
        ein[72]) );
  DFF \ereg_reg[73]  ( .D(ereg_next[73]), .CLK(clk), .RST(rst), .I(e[73]), .Q(
        ein[73]) );
  DFF \ereg_reg[74]  ( .D(ereg_next[74]), .CLK(clk), .RST(rst), .I(e[74]), .Q(
        ein[74]) );
  DFF \ereg_reg[75]  ( .D(ereg_next[75]), .CLK(clk), .RST(rst), .I(e[75]), .Q(
        ein[75]) );
  DFF \ereg_reg[76]  ( .D(ereg_next[76]), .CLK(clk), .RST(rst), .I(e[76]), .Q(
        ein[76]) );
  DFF \ereg_reg[77]  ( .D(ereg_next[77]), .CLK(clk), .RST(rst), .I(e[77]), .Q(
        ein[77]) );
  DFF \ereg_reg[78]  ( .D(ereg_next[78]), .CLK(clk), .RST(rst), .I(e[78]), .Q(
        ein[78]) );
  DFF \ereg_reg[79]  ( .D(ereg_next[79]), .CLK(clk), .RST(rst), .I(e[79]), .Q(
        ein[79]) );
  DFF \ereg_reg[80]  ( .D(ereg_next[80]), .CLK(clk), .RST(rst), .I(e[80]), .Q(
        ein[80]) );
  DFF \ereg_reg[81]  ( .D(ereg_next[81]), .CLK(clk), .RST(rst), .I(e[81]), .Q(
        ein[81]) );
  DFF \ereg_reg[82]  ( .D(ereg_next[82]), .CLK(clk), .RST(rst), .I(e[82]), .Q(
        ein[82]) );
  DFF \ereg_reg[83]  ( .D(ereg_next[83]), .CLK(clk), .RST(rst), .I(e[83]), .Q(
        ein[83]) );
  DFF \ereg_reg[84]  ( .D(ereg_next[84]), .CLK(clk), .RST(rst), .I(e[84]), .Q(
        ein[84]) );
  DFF \ereg_reg[85]  ( .D(ereg_next[85]), .CLK(clk), .RST(rst), .I(e[85]), .Q(
        ein[85]) );
  DFF \ereg_reg[86]  ( .D(ereg_next[86]), .CLK(clk), .RST(rst), .I(e[86]), .Q(
        ein[86]) );
  DFF \ereg_reg[87]  ( .D(ereg_next[87]), .CLK(clk), .RST(rst), .I(e[87]), .Q(
        ein[87]) );
  DFF \ereg_reg[88]  ( .D(ereg_next[88]), .CLK(clk), .RST(rst), .I(e[88]), .Q(
        ein[88]) );
  DFF \ereg_reg[89]  ( .D(ereg_next[89]), .CLK(clk), .RST(rst), .I(e[89]), .Q(
        ein[89]) );
  DFF \ereg_reg[90]  ( .D(ereg_next[90]), .CLK(clk), .RST(rst), .I(e[90]), .Q(
        ein[90]) );
  DFF \ereg_reg[91]  ( .D(ereg_next[91]), .CLK(clk), .RST(rst), .I(e[91]), .Q(
        ein[91]) );
  DFF \ereg_reg[92]  ( .D(ereg_next[92]), .CLK(clk), .RST(rst), .I(e[92]), .Q(
        ein[92]) );
  DFF \ereg_reg[93]  ( .D(ereg_next[93]), .CLK(clk), .RST(rst), .I(e[93]), .Q(
        ein[93]) );
  DFF \ereg_reg[94]  ( .D(ereg_next[94]), .CLK(clk), .RST(rst), .I(e[94]), .Q(
        ein[94]) );
  DFF \ereg_reg[95]  ( .D(ereg_next[95]), .CLK(clk), .RST(rst), .I(e[95]), .Q(
        ein[95]) );
  DFF \ereg_reg[96]  ( .D(ereg_next[96]), .CLK(clk), .RST(rst), .I(e[96]), .Q(
        ein[96]) );
  DFF \ereg_reg[97]  ( .D(ereg_next[97]), .CLK(clk), .RST(rst), .I(e[97]), .Q(
        ein[97]) );
  DFF \ereg_reg[98]  ( .D(ereg_next[98]), .CLK(clk), .RST(rst), .I(e[98]), .Q(
        ein[98]) );
  DFF \ereg_reg[99]  ( .D(ereg_next[99]), .CLK(clk), .RST(rst), .I(e[99]), .Q(
        ein[99]) );
  DFF \ereg_reg[100]  ( .D(ereg_next[100]), .CLK(clk), .RST(rst), .I(e[100]), 
        .Q(ein[100]) );
  DFF \ereg_reg[101]  ( .D(ereg_next[101]), .CLK(clk), .RST(rst), .I(e[101]), 
        .Q(ein[101]) );
  DFF \ereg_reg[102]  ( .D(ereg_next[102]), .CLK(clk), .RST(rst), .I(e[102]), 
        .Q(ein[102]) );
  DFF \ereg_reg[103]  ( .D(ereg_next[103]), .CLK(clk), .RST(rst), .I(e[103]), 
        .Q(ein[103]) );
  DFF \ereg_reg[104]  ( .D(ereg_next[104]), .CLK(clk), .RST(rst), .I(e[104]), 
        .Q(ein[104]) );
  DFF \ereg_reg[105]  ( .D(ereg_next[105]), .CLK(clk), .RST(rst), .I(e[105]), 
        .Q(ein[105]) );
  DFF \ereg_reg[106]  ( .D(ereg_next[106]), .CLK(clk), .RST(rst), .I(e[106]), 
        .Q(ein[106]) );
  DFF \ereg_reg[107]  ( .D(ereg_next[107]), .CLK(clk), .RST(rst), .I(e[107]), 
        .Q(ein[107]) );
  DFF \ereg_reg[108]  ( .D(ereg_next[108]), .CLK(clk), .RST(rst), .I(e[108]), 
        .Q(ein[108]) );
  DFF \ereg_reg[109]  ( .D(ereg_next[109]), .CLK(clk), .RST(rst), .I(e[109]), 
        .Q(ein[109]) );
  DFF \ereg_reg[110]  ( .D(ereg_next[110]), .CLK(clk), .RST(rst), .I(e[110]), 
        .Q(ein[110]) );
  DFF \ereg_reg[111]  ( .D(ereg_next[111]), .CLK(clk), .RST(rst), .I(e[111]), 
        .Q(ein[111]) );
  DFF \ereg_reg[112]  ( .D(ereg_next[112]), .CLK(clk), .RST(rst), .I(e[112]), 
        .Q(ein[112]) );
  DFF \ereg_reg[113]  ( .D(ereg_next[113]), .CLK(clk), .RST(rst), .I(e[113]), 
        .Q(ein[113]) );
  DFF \ereg_reg[114]  ( .D(ereg_next[114]), .CLK(clk), .RST(rst), .I(e[114]), 
        .Q(ein[114]) );
  DFF \ereg_reg[115]  ( .D(ereg_next[115]), .CLK(clk), .RST(rst), .I(e[115]), 
        .Q(ein[115]) );
  DFF \ereg_reg[116]  ( .D(ereg_next[116]), .CLK(clk), .RST(rst), .I(e[116]), 
        .Q(ein[116]) );
  DFF \ereg_reg[117]  ( .D(ereg_next[117]), .CLK(clk), .RST(rst), .I(e[117]), 
        .Q(ein[117]) );
  DFF \ereg_reg[118]  ( .D(ereg_next[118]), .CLK(clk), .RST(rst), .I(e[118]), 
        .Q(ein[118]) );
  DFF \ereg_reg[119]  ( .D(ereg_next[119]), .CLK(clk), .RST(rst), .I(e[119]), 
        .Q(ein[119]) );
  DFF \ereg_reg[120]  ( .D(ereg_next[120]), .CLK(clk), .RST(rst), .I(e[120]), 
        .Q(ein[120]) );
  DFF \ereg_reg[121]  ( .D(ereg_next[121]), .CLK(clk), .RST(rst), .I(e[121]), 
        .Q(ein[121]) );
  DFF \ereg_reg[122]  ( .D(ereg_next[122]), .CLK(clk), .RST(rst), .I(e[122]), 
        .Q(ein[122]) );
  DFF \ereg_reg[123]  ( .D(ereg_next[123]), .CLK(clk), .RST(rst), .I(e[123]), 
        .Q(ein[123]) );
  DFF \ereg_reg[124]  ( .D(ereg_next[124]), .CLK(clk), .RST(rst), .I(e[124]), 
        .Q(ein[124]) );
  DFF \ereg_reg[125]  ( .D(ereg_next[125]), .CLK(clk), .RST(rst), .I(e[125]), 
        .Q(ein[125]) );
  DFF \ereg_reg[126]  ( .D(ereg_next[126]), .CLK(clk), .RST(rst), .I(e[126]), 
        .Q(ein[126]) );
  DFF \ereg_reg[127]  ( .D(ereg_next[127]), .CLK(clk), .RST(rst), .I(e[127]), 
        .Q(ein[127]) );
  DFF \ereg_reg[128]  ( .D(ereg_next[128]), .CLK(clk), .RST(rst), .I(e[128]), 
        .Q(ein[128]) );
  DFF \ereg_reg[129]  ( .D(ereg_next[129]), .CLK(clk), .RST(rst), .I(e[129]), 
        .Q(ein[129]) );
  DFF \ereg_reg[130]  ( .D(ereg_next[130]), .CLK(clk), .RST(rst), .I(e[130]), 
        .Q(ein[130]) );
  DFF \ereg_reg[131]  ( .D(ereg_next[131]), .CLK(clk), .RST(rst), .I(e[131]), 
        .Q(ein[131]) );
  DFF \ereg_reg[132]  ( .D(ereg_next[132]), .CLK(clk), .RST(rst), .I(e[132]), 
        .Q(ein[132]) );
  DFF \ereg_reg[133]  ( .D(ereg_next[133]), .CLK(clk), .RST(rst), .I(e[133]), 
        .Q(ein[133]) );
  DFF \ereg_reg[134]  ( .D(ereg_next[134]), .CLK(clk), .RST(rst), .I(e[134]), 
        .Q(ein[134]) );
  DFF \ereg_reg[135]  ( .D(ereg_next[135]), .CLK(clk), .RST(rst), .I(e[135]), 
        .Q(ein[135]) );
  DFF \ereg_reg[136]  ( .D(ereg_next[136]), .CLK(clk), .RST(rst), .I(e[136]), 
        .Q(ein[136]) );
  DFF \ereg_reg[137]  ( .D(ereg_next[137]), .CLK(clk), .RST(rst), .I(e[137]), 
        .Q(ein[137]) );
  DFF \ereg_reg[138]  ( .D(ereg_next[138]), .CLK(clk), .RST(rst), .I(e[138]), 
        .Q(ein[138]) );
  DFF \ereg_reg[139]  ( .D(ereg_next[139]), .CLK(clk), .RST(rst), .I(e[139]), 
        .Q(ein[139]) );
  DFF \ereg_reg[140]  ( .D(ereg_next[140]), .CLK(clk), .RST(rst), .I(e[140]), 
        .Q(ein[140]) );
  DFF \ereg_reg[141]  ( .D(ereg_next[141]), .CLK(clk), .RST(rst), .I(e[141]), 
        .Q(ein[141]) );
  DFF \ereg_reg[142]  ( .D(ereg_next[142]), .CLK(clk), .RST(rst), .I(e[142]), 
        .Q(ein[142]) );
  DFF \ereg_reg[143]  ( .D(ereg_next[143]), .CLK(clk), .RST(rst), .I(e[143]), 
        .Q(ein[143]) );
  DFF \ereg_reg[144]  ( .D(ereg_next[144]), .CLK(clk), .RST(rst), .I(e[144]), 
        .Q(ein[144]) );
  DFF \ereg_reg[145]  ( .D(ereg_next[145]), .CLK(clk), .RST(rst), .I(e[145]), 
        .Q(ein[145]) );
  DFF \ereg_reg[146]  ( .D(ereg_next[146]), .CLK(clk), .RST(rst), .I(e[146]), 
        .Q(ein[146]) );
  DFF \ereg_reg[147]  ( .D(ereg_next[147]), .CLK(clk), .RST(rst), .I(e[147]), 
        .Q(ein[147]) );
  DFF \ereg_reg[148]  ( .D(ereg_next[148]), .CLK(clk), .RST(rst), .I(e[148]), 
        .Q(ein[148]) );
  DFF \ereg_reg[149]  ( .D(ereg_next[149]), .CLK(clk), .RST(rst), .I(e[149]), 
        .Q(ein[149]) );
  DFF \ereg_reg[150]  ( .D(ereg_next[150]), .CLK(clk), .RST(rst), .I(e[150]), 
        .Q(ein[150]) );
  DFF \ereg_reg[151]  ( .D(ereg_next[151]), .CLK(clk), .RST(rst), .I(e[151]), 
        .Q(ein[151]) );
  DFF \ereg_reg[152]  ( .D(ereg_next[152]), .CLK(clk), .RST(rst), .I(e[152]), 
        .Q(ein[152]) );
  DFF \ereg_reg[153]  ( .D(ereg_next[153]), .CLK(clk), .RST(rst), .I(e[153]), 
        .Q(ein[153]) );
  DFF \ereg_reg[154]  ( .D(ereg_next[154]), .CLK(clk), .RST(rst), .I(e[154]), 
        .Q(ein[154]) );
  DFF \ereg_reg[155]  ( .D(ereg_next[155]), .CLK(clk), .RST(rst), .I(e[155]), 
        .Q(ein[155]) );
  DFF \ereg_reg[156]  ( .D(ereg_next[156]), .CLK(clk), .RST(rst), .I(e[156]), 
        .Q(ein[156]) );
  DFF \ereg_reg[157]  ( .D(ereg_next[157]), .CLK(clk), .RST(rst), .I(e[157]), 
        .Q(ein[157]) );
  DFF \ereg_reg[158]  ( .D(ereg_next[158]), .CLK(clk), .RST(rst), .I(e[158]), 
        .Q(ein[158]) );
  DFF \ereg_reg[159]  ( .D(ereg_next[159]), .CLK(clk), .RST(rst), .I(e[159]), 
        .Q(ein[159]) );
  DFF \ereg_reg[160]  ( .D(ereg_next[160]), .CLK(clk), .RST(rst), .I(e[160]), 
        .Q(ein[160]) );
  DFF \ereg_reg[161]  ( .D(ereg_next[161]), .CLK(clk), .RST(rst), .I(e[161]), 
        .Q(ein[161]) );
  DFF \ereg_reg[162]  ( .D(ereg_next[162]), .CLK(clk), .RST(rst), .I(e[162]), 
        .Q(ein[162]) );
  DFF \ereg_reg[163]  ( .D(ereg_next[163]), .CLK(clk), .RST(rst), .I(e[163]), 
        .Q(ein[163]) );
  DFF \ereg_reg[164]  ( .D(ereg_next[164]), .CLK(clk), .RST(rst), .I(e[164]), 
        .Q(ein[164]) );
  DFF \ereg_reg[165]  ( .D(ereg_next[165]), .CLK(clk), .RST(rst), .I(e[165]), 
        .Q(ein[165]) );
  DFF \ereg_reg[166]  ( .D(ereg_next[166]), .CLK(clk), .RST(rst), .I(e[166]), 
        .Q(ein[166]) );
  DFF \ereg_reg[167]  ( .D(ereg_next[167]), .CLK(clk), .RST(rst), .I(e[167]), 
        .Q(ein[167]) );
  DFF \ereg_reg[168]  ( .D(ereg_next[168]), .CLK(clk), .RST(rst), .I(e[168]), 
        .Q(ein[168]) );
  DFF \ereg_reg[169]  ( .D(ereg_next[169]), .CLK(clk), .RST(rst), .I(e[169]), 
        .Q(ein[169]) );
  DFF \ereg_reg[170]  ( .D(ereg_next[170]), .CLK(clk), .RST(rst), .I(e[170]), 
        .Q(ein[170]) );
  DFF \ereg_reg[171]  ( .D(ereg_next[171]), .CLK(clk), .RST(rst), .I(e[171]), 
        .Q(ein[171]) );
  DFF \ereg_reg[172]  ( .D(ereg_next[172]), .CLK(clk), .RST(rst), .I(e[172]), 
        .Q(ein[172]) );
  DFF \ereg_reg[173]  ( .D(ereg_next[173]), .CLK(clk), .RST(rst), .I(e[173]), 
        .Q(ein[173]) );
  DFF \ereg_reg[174]  ( .D(ereg_next[174]), .CLK(clk), .RST(rst), .I(e[174]), 
        .Q(ein[174]) );
  DFF \ereg_reg[175]  ( .D(ereg_next[175]), .CLK(clk), .RST(rst), .I(e[175]), 
        .Q(ein[175]) );
  DFF \ereg_reg[176]  ( .D(ereg_next[176]), .CLK(clk), .RST(rst), .I(e[176]), 
        .Q(ein[176]) );
  DFF \ereg_reg[177]  ( .D(ereg_next[177]), .CLK(clk), .RST(rst), .I(e[177]), 
        .Q(ein[177]) );
  DFF \ereg_reg[178]  ( .D(ereg_next[178]), .CLK(clk), .RST(rst), .I(e[178]), 
        .Q(ein[178]) );
  DFF \ereg_reg[179]  ( .D(ereg_next[179]), .CLK(clk), .RST(rst), .I(e[179]), 
        .Q(ein[179]) );
  DFF \ereg_reg[180]  ( .D(ereg_next[180]), .CLK(clk), .RST(rst), .I(e[180]), 
        .Q(ein[180]) );
  DFF \ereg_reg[181]  ( .D(ereg_next[181]), .CLK(clk), .RST(rst), .I(e[181]), 
        .Q(ein[181]) );
  DFF \ereg_reg[182]  ( .D(ereg_next[182]), .CLK(clk), .RST(rst), .I(e[182]), 
        .Q(ein[182]) );
  DFF \ereg_reg[183]  ( .D(ereg_next[183]), .CLK(clk), .RST(rst), .I(e[183]), 
        .Q(ein[183]) );
  DFF \ereg_reg[184]  ( .D(ereg_next[184]), .CLK(clk), .RST(rst), .I(e[184]), 
        .Q(ein[184]) );
  DFF \ereg_reg[185]  ( .D(ereg_next[185]), .CLK(clk), .RST(rst), .I(e[185]), 
        .Q(ein[185]) );
  DFF \ereg_reg[186]  ( .D(ereg_next[186]), .CLK(clk), .RST(rst), .I(e[186]), 
        .Q(ein[186]) );
  DFF \ereg_reg[187]  ( .D(ereg_next[187]), .CLK(clk), .RST(rst), .I(e[187]), 
        .Q(ein[187]) );
  DFF \ereg_reg[188]  ( .D(ereg_next[188]), .CLK(clk), .RST(rst), .I(e[188]), 
        .Q(ein[188]) );
  DFF \ereg_reg[189]  ( .D(ereg_next[189]), .CLK(clk), .RST(rst), .I(e[189]), 
        .Q(ein[189]) );
  DFF \ereg_reg[190]  ( .D(ereg_next[190]), .CLK(clk), .RST(rst), .I(e[190]), 
        .Q(ein[190]) );
  DFF \ereg_reg[191]  ( .D(ereg_next[191]), .CLK(clk), .RST(rst), .I(e[191]), 
        .Q(ein[191]) );
  DFF \ereg_reg[192]  ( .D(ereg_next[192]), .CLK(clk), .RST(rst), .I(e[192]), 
        .Q(ein[192]) );
  DFF \ereg_reg[193]  ( .D(ereg_next[193]), .CLK(clk), .RST(rst), .I(e[193]), 
        .Q(ein[193]) );
  DFF \ereg_reg[194]  ( .D(ereg_next[194]), .CLK(clk), .RST(rst), .I(e[194]), 
        .Q(ein[194]) );
  DFF \ereg_reg[195]  ( .D(ereg_next[195]), .CLK(clk), .RST(rst), .I(e[195]), 
        .Q(ein[195]) );
  DFF \ereg_reg[196]  ( .D(ereg_next[196]), .CLK(clk), .RST(rst), .I(e[196]), 
        .Q(ein[196]) );
  DFF \ereg_reg[197]  ( .D(ereg_next[197]), .CLK(clk), .RST(rst), .I(e[197]), 
        .Q(ein[197]) );
  DFF \ereg_reg[198]  ( .D(ereg_next[198]), .CLK(clk), .RST(rst), .I(e[198]), 
        .Q(ein[198]) );
  DFF \ereg_reg[199]  ( .D(ereg_next[199]), .CLK(clk), .RST(rst), .I(e[199]), 
        .Q(ein[199]) );
  DFF \ereg_reg[200]  ( .D(ereg_next[200]), .CLK(clk), .RST(rst), .I(e[200]), 
        .Q(ein[200]) );
  DFF \ereg_reg[201]  ( .D(ereg_next[201]), .CLK(clk), .RST(rst), .I(e[201]), 
        .Q(ein[201]) );
  DFF \ereg_reg[202]  ( .D(ereg_next[202]), .CLK(clk), .RST(rst), .I(e[202]), 
        .Q(ein[202]) );
  DFF \ereg_reg[203]  ( .D(ereg_next[203]), .CLK(clk), .RST(rst), .I(e[203]), 
        .Q(ein[203]) );
  DFF \ereg_reg[204]  ( .D(ereg_next[204]), .CLK(clk), .RST(rst), .I(e[204]), 
        .Q(ein[204]) );
  DFF \ereg_reg[205]  ( .D(ereg_next[205]), .CLK(clk), .RST(rst), .I(e[205]), 
        .Q(ein[205]) );
  DFF \ereg_reg[206]  ( .D(ereg_next[206]), .CLK(clk), .RST(rst), .I(e[206]), 
        .Q(ein[206]) );
  DFF \ereg_reg[207]  ( .D(ereg_next[207]), .CLK(clk), .RST(rst), .I(e[207]), 
        .Q(ein[207]) );
  DFF \ereg_reg[208]  ( .D(ereg_next[208]), .CLK(clk), .RST(rst), .I(e[208]), 
        .Q(ein[208]) );
  DFF \ereg_reg[209]  ( .D(ereg_next[209]), .CLK(clk), .RST(rst), .I(e[209]), 
        .Q(ein[209]) );
  DFF \ereg_reg[210]  ( .D(ereg_next[210]), .CLK(clk), .RST(rst), .I(e[210]), 
        .Q(ein[210]) );
  DFF \ereg_reg[211]  ( .D(ereg_next[211]), .CLK(clk), .RST(rst), .I(e[211]), 
        .Q(ein[211]) );
  DFF \ereg_reg[212]  ( .D(ereg_next[212]), .CLK(clk), .RST(rst), .I(e[212]), 
        .Q(ein[212]) );
  DFF \ereg_reg[213]  ( .D(ereg_next[213]), .CLK(clk), .RST(rst), .I(e[213]), 
        .Q(ein[213]) );
  DFF \ereg_reg[214]  ( .D(ereg_next[214]), .CLK(clk), .RST(rst), .I(e[214]), 
        .Q(ein[214]) );
  DFF \ereg_reg[215]  ( .D(ereg_next[215]), .CLK(clk), .RST(rst), .I(e[215]), 
        .Q(ein[215]) );
  DFF \ereg_reg[216]  ( .D(ereg_next[216]), .CLK(clk), .RST(rst), .I(e[216]), 
        .Q(ein[216]) );
  DFF \ereg_reg[217]  ( .D(ereg_next[217]), .CLK(clk), .RST(rst), .I(e[217]), 
        .Q(ein[217]) );
  DFF \ereg_reg[218]  ( .D(ereg_next[218]), .CLK(clk), .RST(rst), .I(e[218]), 
        .Q(ein[218]) );
  DFF \ereg_reg[219]  ( .D(ereg_next[219]), .CLK(clk), .RST(rst), .I(e[219]), 
        .Q(ein[219]) );
  DFF \ereg_reg[220]  ( .D(ereg_next[220]), .CLK(clk), .RST(rst), .I(e[220]), 
        .Q(ein[220]) );
  DFF \ereg_reg[221]  ( .D(ereg_next[221]), .CLK(clk), .RST(rst), .I(e[221]), 
        .Q(ein[221]) );
  DFF \ereg_reg[222]  ( .D(ereg_next[222]), .CLK(clk), .RST(rst), .I(e[222]), 
        .Q(ein[222]) );
  DFF \ereg_reg[223]  ( .D(ereg_next[223]), .CLK(clk), .RST(rst), .I(e[223]), 
        .Q(ein[223]) );
  DFF \ereg_reg[224]  ( .D(ereg_next[224]), .CLK(clk), .RST(rst), .I(e[224]), 
        .Q(ein[224]) );
  DFF \ereg_reg[225]  ( .D(ereg_next[225]), .CLK(clk), .RST(rst), .I(e[225]), 
        .Q(ein[225]) );
  DFF \ereg_reg[226]  ( .D(ereg_next[226]), .CLK(clk), .RST(rst), .I(e[226]), 
        .Q(ein[226]) );
  DFF \ereg_reg[227]  ( .D(ereg_next[227]), .CLK(clk), .RST(rst), .I(e[227]), 
        .Q(ein[227]) );
  DFF \ereg_reg[228]  ( .D(ereg_next[228]), .CLK(clk), .RST(rst), .I(e[228]), 
        .Q(ein[228]) );
  DFF \ereg_reg[229]  ( .D(ereg_next[229]), .CLK(clk), .RST(rst), .I(e[229]), 
        .Q(ein[229]) );
  DFF \ereg_reg[230]  ( .D(ereg_next[230]), .CLK(clk), .RST(rst), .I(e[230]), 
        .Q(ein[230]) );
  DFF \ereg_reg[231]  ( .D(ereg_next[231]), .CLK(clk), .RST(rst), .I(e[231]), 
        .Q(ein[231]) );
  DFF \ereg_reg[232]  ( .D(ereg_next[232]), .CLK(clk), .RST(rst), .I(e[232]), 
        .Q(ein[232]) );
  DFF \ereg_reg[233]  ( .D(ereg_next[233]), .CLK(clk), .RST(rst), .I(e[233]), 
        .Q(ein[233]) );
  DFF \ereg_reg[234]  ( .D(ereg_next[234]), .CLK(clk), .RST(rst), .I(e[234]), 
        .Q(ein[234]) );
  DFF \ereg_reg[235]  ( .D(ereg_next[235]), .CLK(clk), .RST(rst), .I(e[235]), 
        .Q(ein[235]) );
  DFF \ereg_reg[236]  ( .D(ereg_next[236]), .CLK(clk), .RST(rst), .I(e[236]), 
        .Q(ein[236]) );
  DFF \ereg_reg[237]  ( .D(ereg_next[237]), .CLK(clk), .RST(rst), .I(e[237]), 
        .Q(ein[237]) );
  DFF \ereg_reg[238]  ( .D(ereg_next[238]), .CLK(clk), .RST(rst), .I(e[238]), 
        .Q(ein[238]) );
  DFF \ereg_reg[239]  ( .D(ereg_next[239]), .CLK(clk), .RST(rst), .I(e[239]), 
        .Q(ein[239]) );
  DFF \ereg_reg[240]  ( .D(ereg_next[240]), .CLK(clk), .RST(rst), .I(e[240]), 
        .Q(ein[240]) );
  DFF \ereg_reg[241]  ( .D(ereg_next[241]), .CLK(clk), .RST(rst), .I(e[241]), 
        .Q(ein[241]) );
  DFF \ereg_reg[242]  ( .D(ereg_next[242]), .CLK(clk), .RST(rst), .I(e[242]), 
        .Q(ein[242]) );
  DFF \ereg_reg[243]  ( .D(ereg_next[243]), .CLK(clk), .RST(rst), .I(e[243]), 
        .Q(ein[243]) );
  DFF \ereg_reg[244]  ( .D(ereg_next[244]), .CLK(clk), .RST(rst), .I(e[244]), 
        .Q(ein[244]) );
  DFF \ereg_reg[245]  ( .D(ereg_next[245]), .CLK(clk), .RST(rst), .I(e[245]), 
        .Q(ein[245]) );
  DFF \ereg_reg[246]  ( .D(ereg_next[246]), .CLK(clk), .RST(rst), .I(e[246]), 
        .Q(ein[246]) );
  DFF \ereg_reg[247]  ( .D(ereg_next[247]), .CLK(clk), .RST(rst), .I(e[247]), 
        .Q(ein[247]) );
  DFF \ereg_reg[248]  ( .D(ereg_next[248]), .CLK(clk), .RST(rst), .I(e[248]), 
        .Q(ein[248]) );
  DFF \ereg_reg[249]  ( .D(ereg_next[249]), .CLK(clk), .RST(rst), .I(e[249]), 
        .Q(ein[249]) );
  DFF \ereg_reg[250]  ( .D(ereg_next[250]), .CLK(clk), .RST(rst), .I(e[250]), 
        .Q(ein[250]) );
  DFF \ereg_reg[251]  ( .D(ereg_next[251]), .CLK(clk), .RST(rst), .I(e[251]), 
        .Q(ein[251]) );
  DFF \ereg_reg[252]  ( .D(ereg_next[252]), .CLK(clk), .RST(rst), .I(e[252]), 
        .Q(ein[252]) );
  DFF \ereg_reg[253]  ( .D(ereg_next[253]), .CLK(clk), .RST(rst), .I(e[253]), 
        .Q(ein[253]) );
  DFF \ereg_reg[254]  ( .D(ereg_next[254]), .CLK(clk), .RST(rst), .I(e[254]), 
        .Q(ein[254]) );
  DFF \ereg_reg[255]  ( .D(ereg_next[255]), .CLK(clk), .RST(rst), .I(e[255]), 
        .Q(ein[255]) );
  DFF \ereg_reg[256]  ( .D(ereg_next[256]), .CLK(clk), .RST(rst), .I(e[256]), 
        .Q(ein[256]) );
  DFF \ereg_reg[257]  ( .D(ereg_next[257]), .CLK(clk), .RST(rst), .I(e[257]), 
        .Q(ein[257]) );
  DFF \ereg_reg[258]  ( .D(ereg_next[258]), .CLK(clk), .RST(rst), .I(e[258]), 
        .Q(ein[258]) );
  DFF \ereg_reg[259]  ( .D(ereg_next[259]), .CLK(clk), .RST(rst), .I(e[259]), 
        .Q(ein[259]) );
  DFF \ereg_reg[260]  ( .D(ereg_next[260]), .CLK(clk), .RST(rst), .I(e[260]), 
        .Q(ein[260]) );
  DFF \ereg_reg[261]  ( .D(ereg_next[261]), .CLK(clk), .RST(rst), .I(e[261]), 
        .Q(ein[261]) );
  DFF \ereg_reg[262]  ( .D(ereg_next[262]), .CLK(clk), .RST(rst), .I(e[262]), 
        .Q(ein[262]) );
  DFF \ereg_reg[263]  ( .D(ereg_next[263]), .CLK(clk), .RST(rst), .I(e[263]), 
        .Q(ein[263]) );
  DFF \ereg_reg[264]  ( .D(ereg_next[264]), .CLK(clk), .RST(rst), .I(e[264]), 
        .Q(ein[264]) );
  DFF \ereg_reg[265]  ( .D(ereg_next[265]), .CLK(clk), .RST(rst), .I(e[265]), 
        .Q(ein[265]) );
  DFF \ereg_reg[266]  ( .D(ereg_next[266]), .CLK(clk), .RST(rst), .I(e[266]), 
        .Q(ein[266]) );
  DFF \ereg_reg[267]  ( .D(ereg_next[267]), .CLK(clk), .RST(rst), .I(e[267]), 
        .Q(ein[267]) );
  DFF \ereg_reg[268]  ( .D(ereg_next[268]), .CLK(clk), .RST(rst), .I(e[268]), 
        .Q(ein[268]) );
  DFF \ereg_reg[269]  ( .D(ereg_next[269]), .CLK(clk), .RST(rst), .I(e[269]), 
        .Q(ein[269]) );
  DFF \ereg_reg[270]  ( .D(ereg_next[270]), .CLK(clk), .RST(rst), .I(e[270]), 
        .Q(ein[270]) );
  DFF \ereg_reg[271]  ( .D(ereg_next[271]), .CLK(clk), .RST(rst), .I(e[271]), 
        .Q(ein[271]) );
  DFF \ereg_reg[272]  ( .D(ereg_next[272]), .CLK(clk), .RST(rst), .I(e[272]), 
        .Q(ein[272]) );
  DFF \ereg_reg[273]  ( .D(ereg_next[273]), .CLK(clk), .RST(rst), .I(e[273]), 
        .Q(ein[273]) );
  DFF \ereg_reg[274]  ( .D(ereg_next[274]), .CLK(clk), .RST(rst), .I(e[274]), 
        .Q(ein[274]) );
  DFF \ereg_reg[275]  ( .D(ereg_next[275]), .CLK(clk), .RST(rst), .I(e[275]), 
        .Q(ein[275]) );
  DFF \ereg_reg[276]  ( .D(ereg_next[276]), .CLK(clk), .RST(rst), .I(e[276]), 
        .Q(ein[276]) );
  DFF \ereg_reg[277]  ( .D(ereg_next[277]), .CLK(clk), .RST(rst), .I(e[277]), 
        .Q(ein[277]) );
  DFF \ereg_reg[278]  ( .D(ereg_next[278]), .CLK(clk), .RST(rst), .I(e[278]), 
        .Q(ein[278]) );
  DFF \ereg_reg[279]  ( .D(ereg_next[279]), .CLK(clk), .RST(rst), .I(e[279]), 
        .Q(ein[279]) );
  DFF \ereg_reg[280]  ( .D(ereg_next[280]), .CLK(clk), .RST(rst), .I(e[280]), 
        .Q(ein[280]) );
  DFF \ereg_reg[281]  ( .D(ereg_next[281]), .CLK(clk), .RST(rst), .I(e[281]), 
        .Q(ein[281]) );
  DFF \ereg_reg[282]  ( .D(ereg_next[282]), .CLK(clk), .RST(rst), .I(e[282]), 
        .Q(ein[282]) );
  DFF \ereg_reg[283]  ( .D(ereg_next[283]), .CLK(clk), .RST(rst), .I(e[283]), 
        .Q(ein[283]) );
  DFF \ereg_reg[284]  ( .D(ereg_next[284]), .CLK(clk), .RST(rst), .I(e[284]), 
        .Q(ein[284]) );
  DFF \ereg_reg[285]  ( .D(ereg_next[285]), .CLK(clk), .RST(rst), .I(e[285]), 
        .Q(ein[285]) );
  DFF \ereg_reg[286]  ( .D(ereg_next[286]), .CLK(clk), .RST(rst), .I(e[286]), 
        .Q(ein[286]) );
  DFF \ereg_reg[287]  ( .D(ereg_next[287]), .CLK(clk), .RST(rst), .I(e[287]), 
        .Q(ein[287]) );
  DFF \ereg_reg[288]  ( .D(ereg_next[288]), .CLK(clk), .RST(rst), .I(e[288]), 
        .Q(ein[288]) );
  DFF \ereg_reg[289]  ( .D(ereg_next[289]), .CLK(clk), .RST(rst), .I(e[289]), 
        .Q(ein[289]) );
  DFF \ereg_reg[290]  ( .D(ereg_next[290]), .CLK(clk), .RST(rst), .I(e[290]), 
        .Q(ein[290]) );
  DFF \ereg_reg[291]  ( .D(ereg_next[291]), .CLK(clk), .RST(rst), .I(e[291]), 
        .Q(ein[291]) );
  DFF \ereg_reg[292]  ( .D(ereg_next[292]), .CLK(clk), .RST(rst), .I(e[292]), 
        .Q(ein[292]) );
  DFF \ereg_reg[293]  ( .D(ereg_next[293]), .CLK(clk), .RST(rst), .I(e[293]), 
        .Q(ein[293]) );
  DFF \ereg_reg[294]  ( .D(ereg_next[294]), .CLK(clk), .RST(rst), .I(e[294]), 
        .Q(ein[294]) );
  DFF \ereg_reg[295]  ( .D(ereg_next[295]), .CLK(clk), .RST(rst), .I(e[295]), 
        .Q(ein[295]) );
  DFF \ereg_reg[296]  ( .D(ereg_next[296]), .CLK(clk), .RST(rst), .I(e[296]), 
        .Q(ein[296]) );
  DFF \ereg_reg[297]  ( .D(ereg_next[297]), .CLK(clk), .RST(rst), .I(e[297]), 
        .Q(ein[297]) );
  DFF \ereg_reg[298]  ( .D(ereg_next[298]), .CLK(clk), .RST(rst), .I(e[298]), 
        .Q(ein[298]) );
  DFF \ereg_reg[299]  ( .D(ereg_next[299]), .CLK(clk), .RST(rst), .I(e[299]), 
        .Q(ein[299]) );
  DFF \ereg_reg[300]  ( .D(ereg_next[300]), .CLK(clk), .RST(rst), .I(e[300]), 
        .Q(ein[300]) );
  DFF \ereg_reg[301]  ( .D(ereg_next[301]), .CLK(clk), .RST(rst), .I(e[301]), 
        .Q(ein[301]) );
  DFF \ereg_reg[302]  ( .D(ereg_next[302]), .CLK(clk), .RST(rst), .I(e[302]), 
        .Q(ein[302]) );
  DFF \ereg_reg[303]  ( .D(ereg_next[303]), .CLK(clk), .RST(rst), .I(e[303]), 
        .Q(ein[303]) );
  DFF \ereg_reg[304]  ( .D(ereg_next[304]), .CLK(clk), .RST(rst), .I(e[304]), 
        .Q(ein[304]) );
  DFF \ereg_reg[305]  ( .D(ereg_next[305]), .CLK(clk), .RST(rst), .I(e[305]), 
        .Q(ein[305]) );
  DFF \ereg_reg[306]  ( .D(ereg_next[306]), .CLK(clk), .RST(rst), .I(e[306]), 
        .Q(ein[306]) );
  DFF \ereg_reg[307]  ( .D(ereg_next[307]), .CLK(clk), .RST(rst), .I(e[307]), 
        .Q(ein[307]) );
  DFF \ereg_reg[308]  ( .D(ereg_next[308]), .CLK(clk), .RST(rst), .I(e[308]), 
        .Q(ein[308]) );
  DFF \ereg_reg[309]  ( .D(ereg_next[309]), .CLK(clk), .RST(rst), .I(e[309]), 
        .Q(ein[309]) );
  DFF \ereg_reg[310]  ( .D(ereg_next[310]), .CLK(clk), .RST(rst), .I(e[310]), 
        .Q(ein[310]) );
  DFF \ereg_reg[311]  ( .D(ereg_next[311]), .CLK(clk), .RST(rst), .I(e[311]), 
        .Q(ein[311]) );
  DFF \ereg_reg[312]  ( .D(ereg_next[312]), .CLK(clk), .RST(rst), .I(e[312]), 
        .Q(ein[312]) );
  DFF \ereg_reg[313]  ( .D(ereg_next[313]), .CLK(clk), .RST(rst), .I(e[313]), 
        .Q(ein[313]) );
  DFF \ereg_reg[314]  ( .D(ereg_next[314]), .CLK(clk), .RST(rst), .I(e[314]), 
        .Q(ein[314]) );
  DFF \ereg_reg[315]  ( .D(ereg_next[315]), .CLK(clk), .RST(rst), .I(e[315]), 
        .Q(ein[315]) );
  DFF \ereg_reg[316]  ( .D(ereg_next[316]), .CLK(clk), .RST(rst), .I(e[316]), 
        .Q(ein[316]) );
  DFF \ereg_reg[317]  ( .D(ereg_next[317]), .CLK(clk), .RST(rst), .I(e[317]), 
        .Q(ein[317]) );
  DFF \ereg_reg[318]  ( .D(ereg_next[318]), .CLK(clk), .RST(rst), .I(e[318]), 
        .Q(ein[318]) );
  DFF \ereg_reg[319]  ( .D(ereg_next[319]), .CLK(clk), .RST(rst), .I(e[319]), 
        .Q(ein[319]) );
  DFF \ereg_reg[320]  ( .D(ereg_next[320]), .CLK(clk), .RST(rst), .I(e[320]), 
        .Q(ein[320]) );
  DFF \ereg_reg[321]  ( .D(ereg_next[321]), .CLK(clk), .RST(rst), .I(e[321]), 
        .Q(ein[321]) );
  DFF \ereg_reg[322]  ( .D(ereg_next[322]), .CLK(clk), .RST(rst), .I(e[322]), 
        .Q(ein[322]) );
  DFF \ereg_reg[323]  ( .D(ereg_next[323]), .CLK(clk), .RST(rst), .I(e[323]), 
        .Q(ein[323]) );
  DFF \ereg_reg[324]  ( .D(ereg_next[324]), .CLK(clk), .RST(rst), .I(e[324]), 
        .Q(ein[324]) );
  DFF \ereg_reg[325]  ( .D(ereg_next[325]), .CLK(clk), .RST(rst), .I(e[325]), 
        .Q(ein[325]) );
  DFF \ereg_reg[326]  ( .D(ereg_next[326]), .CLK(clk), .RST(rst), .I(e[326]), 
        .Q(ein[326]) );
  DFF \ereg_reg[327]  ( .D(ereg_next[327]), .CLK(clk), .RST(rst), .I(e[327]), 
        .Q(ein[327]) );
  DFF \ereg_reg[328]  ( .D(ereg_next[328]), .CLK(clk), .RST(rst), .I(e[328]), 
        .Q(ein[328]) );
  DFF \ereg_reg[329]  ( .D(ereg_next[329]), .CLK(clk), .RST(rst), .I(e[329]), 
        .Q(ein[329]) );
  DFF \ereg_reg[330]  ( .D(ereg_next[330]), .CLK(clk), .RST(rst), .I(e[330]), 
        .Q(ein[330]) );
  DFF \ereg_reg[331]  ( .D(ereg_next[331]), .CLK(clk), .RST(rst), .I(e[331]), 
        .Q(ein[331]) );
  DFF \ereg_reg[332]  ( .D(ereg_next[332]), .CLK(clk), .RST(rst), .I(e[332]), 
        .Q(ein[332]) );
  DFF \ereg_reg[333]  ( .D(ereg_next[333]), .CLK(clk), .RST(rst), .I(e[333]), 
        .Q(ein[333]) );
  DFF \ereg_reg[334]  ( .D(ereg_next[334]), .CLK(clk), .RST(rst), .I(e[334]), 
        .Q(ein[334]) );
  DFF \ereg_reg[335]  ( .D(ereg_next[335]), .CLK(clk), .RST(rst), .I(e[335]), 
        .Q(ein[335]) );
  DFF \ereg_reg[336]  ( .D(ereg_next[336]), .CLK(clk), .RST(rst), .I(e[336]), 
        .Q(ein[336]) );
  DFF \ereg_reg[337]  ( .D(ereg_next[337]), .CLK(clk), .RST(rst), .I(e[337]), 
        .Q(ein[337]) );
  DFF \ereg_reg[338]  ( .D(ereg_next[338]), .CLK(clk), .RST(rst), .I(e[338]), 
        .Q(ein[338]) );
  DFF \ereg_reg[339]  ( .D(ereg_next[339]), .CLK(clk), .RST(rst), .I(e[339]), 
        .Q(ein[339]) );
  DFF \ereg_reg[340]  ( .D(ereg_next[340]), .CLK(clk), .RST(rst), .I(e[340]), 
        .Q(ein[340]) );
  DFF \ereg_reg[341]  ( .D(ereg_next[341]), .CLK(clk), .RST(rst), .I(e[341]), 
        .Q(ein[341]) );
  DFF \ereg_reg[342]  ( .D(ereg_next[342]), .CLK(clk), .RST(rst), .I(e[342]), 
        .Q(ein[342]) );
  DFF \ereg_reg[343]  ( .D(ereg_next[343]), .CLK(clk), .RST(rst), .I(e[343]), 
        .Q(ein[343]) );
  DFF \ereg_reg[344]  ( .D(ereg_next[344]), .CLK(clk), .RST(rst), .I(e[344]), 
        .Q(ein[344]) );
  DFF \ereg_reg[345]  ( .D(ereg_next[345]), .CLK(clk), .RST(rst), .I(e[345]), 
        .Q(ein[345]) );
  DFF \ereg_reg[346]  ( .D(ereg_next[346]), .CLK(clk), .RST(rst), .I(e[346]), 
        .Q(ein[346]) );
  DFF \ereg_reg[347]  ( .D(ereg_next[347]), .CLK(clk), .RST(rst), .I(e[347]), 
        .Q(ein[347]) );
  DFF \ereg_reg[348]  ( .D(ereg_next[348]), .CLK(clk), .RST(rst), .I(e[348]), 
        .Q(ein[348]) );
  DFF \ereg_reg[349]  ( .D(ereg_next[349]), .CLK(clk), .RST(rst), .I(e[349]), 
        .Q(ein[349]) );
  DFF \ereg_reg[350]  ( .D(ereg_next[350]), .CLK(clk), .RST(rst), .I(e[350]), 
        .Q(ein[350]) );
  DFF \ereg_reg[351]  ( .D(ereg_next[351]), .CLK(clk), .RST(rst), .I(e[351]), 
        .Q(ein[351]) );
  DFF \ereg_reg[352]  ( .D(ereg_next[352]), .CLK(clk), .RST(rst), .I(e[352]), 
        .Q(ein[352]) );
  DFF \ereg_reg[353]  ( .D(ereg_next[353]), .CLK(clk), .RST(rst), .I(e[353]), 
        .Q(ein[353]) );
  DFF \ereg_reg[354]  ( .D(ereg_next[354]), .CLK(clk), .RST(rst), .I(e[354]), 
        .Q(ein[354]) );
  DFF \ereg_reg[355]  ( .D(ereg_next[355]), .CLK(clk), .RST(rst), .I(e[355]), 
        .Q(ein[355]) );
  DFF \ereg_reg[356]  ( .D(ereg_next[356]), .CLK(clk), .RST(rst), .I(e[356]), 
        .Q(ein[356]) );
  DFF \ereg_reg[357]  ( .D(ereg_next[357]), .CLK(clk), .RST(rst), .I(e[357]), 
        .Q(ein[357]) );
  DFF \ereg_reg[358]  ( .D(ereg_next[358]), .CLK(clk), .RST(rst), .I(e[358]), 
        .Q(ein[358]) );
  DFF \ereg_reg[359]  ( .D(ereg_next[359]), .CLK(clk), .RST(rst), .I(e[359]), 
        .Q(ein[359]) );
  DFF \ereg_reg[360]  ( .D(ereg_next[360]), .CLK(clk), .RST(rst), .I(e[360]), 
        .Q(ein[360]) );
  DFF \ereg_reg[361]  ( .D(ereg_next[361]), .CLK(clk), .RST(rst), .I(e[361]), 
        .Q(ein[361]) );
  DFF \ereg_reg[362]  ( .D(ereg_next[362]), .CLK(clk), .RST(rst), .I(e[362]), 
        .Q(ein[362]) );
  DFF \ereg_reg[363]  ( .D(ereg_next[363]), .CLK(clk), .RST(rst), .I(e[363]), 
        .Q(ein[363]) );
  DFF \ereg_reg[364]  ( .D(ereg_next[364]), .CLK(clk), .RST(rst), .I(e[364]), 
        .Q(ein[364]) );
  DFF \ereg_reg[365]  ( .D(ereg_next[365]), .CLK(clk), .RST(rst), .I(e[365]), 
        .Q(ein[365]) );
  DFF \ereg_reg[366]  ( .D(ereg_next[366]), .CLK(clk), .RST(rst), .I(e[366]), 
        .Q(ein[366]) );
  DFF \ereg_reg[367]  ( .D(ereg_next[367]), .CLK(clk), .RST(rst), .I(e[367]), 
        .Q(ein[367]) );
  DFF \ereg_reg[368]  ( .D(ereg_next[368]), .CLK(clk), .RST(rst), .I(e[368]), 
        .Q(ein[368]) );
  DFF \ereg_reg[369]  ( .D(ereg_next[369]), .CLK(clk), .RST(rst), .I(e[369]), 
        .Q(ein[369]) );
  DFF \ereg_reg[370]  ( .D(ereg_next[370]), .CLK(clk), .RST(rst), .I(e[370]), 
        .Q(ein[370]) );
  DFF \ereg_reg[371]  ( .D(ereg_next[371]), .CLK(clk), .RST(rst), .I(e[371]), 
        .Q(ein[371]) );
  DFF \ereg_reg[372]  ( .D(ereg_next[372]), .CLK(clk), .RST(rst), .I(e[372]), 
        .Q(ein[372]) );
  DFF \ereg_reg[373]  ( .D(ereg_next[373]), .CLK(clk), .RST(rst), .I(e[373]), 
        .Q(ein[373]) );
  DFF \ereg_reg[374]  ( .D(ereg_next[374]), .CLK(clk), .RST(rst), .I(e[374]), 
        .Q(ein[374]) );
  DFF \ereg_reg[375]  ( .D(ereg_next[375]), .CLK(clk), .RST(rst), .I(e[375]), 
        .Q(ein[375]) );
  DFF \ereg_reg[376]  ( .D(ereg_next[376]), .CLK(clk), .RST(rst), .I(e[376]), 
        .Q(ein[376]) );
  DFF \ereg_reg[377]  ( .D(ereg_next[377]), .CLK(clk), .RST(rst), .I(e[377]), 
        .Q(ein[377]) );
  DFF \ereg_reg[378]  ( .D(ereg_next[378]), .CLK(clk), .RST(rst), .I(e[378]), 
        .Q(ein[378]) );
  DFF \ereg_reg[379]  ( .D(ereg_next[379]), .CLK(clk), .RST(rst), .I(e[379]), 
        .Q(ein[379]) );
  DFF \ereg_reg[380]  ( .D(ereg_next[380]), .CLK(clk), .RST(rst), .I(e[380]), 
        .Q(ein[380]) );
  DFF \ereg_reg[381]  ( .D(ereg_next[381]), .CLK(clk), .RST(rst), .I(e[381]), 
        .Q(ein[381]) );
  DFF \ereg_reg[382]  ( .D(ereg_next[382]), .CLK(clk), .RST(rst), .I(e[382]), 
        .Q(ein[382]) );
  DFF \ereg_reg[383]  ( .D(ereg_next[383]), .CLK(clk), .RST(rst), .I(e[383]), 
        .Q(ein[383]) );
  DFF \ereg_reg[384]  ( .D(ereg_next[384]), .CLK(clk), .RST(rst), .I(e[384]), 
        .Q(ein[384]) );
  DFF \ereg_reg[385]  ( .D(ereg_next[385]), .CLK(clk), .RST(rst), .I(e[385]), 
        .Q(ein[385]) );
  DFF \ereg_reg[386]  ( .D(ereg_next[386]), .CLK(clk), .RST(rst), .I(e[386]), 
        .Q(ein[386]) );
  DFF \ereg_reg[387]  ( .D(ereg_next[387]), .CLK(clk), .RST(rst), .I(e[387]), 
        .Q(ein[387]) );
  DFF \ereg_reg[388]  ( .D(ereg_next[388]), .CLK(clk), .RST(rst), .I(e[388]), 
        .Q(ein[388]) );
  DFF \ereg_reg[389]  ( .D(ereg_next[389]), .CLK(clk), .RST(rst), .I(e[389]), 
        .Q(ein[389]) );
  DFF \ereg_reg[390]  ( .D(ereg_next[390]), .CLK(clk), .RST(rst), .I(e[390]), 
        .Q(ein[390]) );
  DFF \ereg_reg[391]  ( .D(ereg_next[391]), .CLK(clk), .RST(rst), .I(e[391]), 
        .Q(ein[391]) );
  DFF \ereg_reg[392]  ( .D(ereg_next[392]), .CLK(clk), .RST(rst), .I(e[392]), 
        .Q(ein[392]) );
  DFF \ereg_reg[393]  ( .D(ereg_next[393]), .CLK(clk), .RST(rst), .I(e[393]), 
        .Q(ein[393]) );
  DFF \ereg_reg[394]  ( .D(ereg_next[394]), .CLK(clk), .RST(rst), .I(e[394]), 
        .Q(ein[394]) );
  DFF \ereg_reg[395]  ( .D(ereg_next[395]), .CLK(clk), .RST(rst), .I(e[395]), 
        .Q(ein[395]) );
  DFF \ereg_reg[396]  ( .D(ereg_next[396]), .CLK(clk), .RST(rst), .I(e[396]), 
        .Q(ein[396]) );
  DFF \ereg_reg[397]  ( .D(ereg_next[397]), .CLK(clk), .RST(rst), .I(e[397]), 
        .Q(ein[397]) );
  DFF \ereg_reg[398]  ( .D(ereg_next[398]), .CLK(clk), .RST(rst), .I(e[398]), 
        .Q(ein[398]) );
  DFF \ereg_reg[399]  ( .D(ereg_next[399]), .CLK(clk), .RST(rst), .I(e[399]), 
        .Q(ein[399]) );
  DFF \ereg_reg[400]  ( .D(ereg_next[400]), .CLK(clk), .RST(rst), .I(e[400]), 
        .Q(ein[400]) );
  DFF \ereg_reg[401]  ( .D(ereg_next[401]), .CLK(clk), .RST(rst), .I(e[401]), 
        .Q(ein[401]) );
  DFF \ereg_reg[402]  ( .D(ereg_next[402]), .CLK(clk), .RST(rst), .I(e[402]), 
        .Q(ein[402]) );
  DFF \ereg_reg[403]  ( .D(ereg_next[403]), .CLK(clk), .RST(rst), .I(e[403]), 
        .Q(ein[403]) );
  DFF \ereg_reg[404]  ( .D(ereg_next[404]), .CLK(clk), .RST(rst), .I(e[404]), 
        .Q(ein[404]) );
  DFF \ereg_reg[405]  ( .D(ereg_next[405]), .CLK(clk), .RST(rst), .I(e[405]), 
        .Q(ein[405]) );
  DFF \ereg_reg[406]  ( .D(ereg_next[406]), .CLK(clk), .RST(rst), .I(e[406]), 
        .Q(ein[406]) );
  DFF \ereg_reg[407]  ( .D(ereg_next[407]), .CLK(clk), .RST(rst), .I(e[407]), 
        .Q(ein[407]) );
  DFF \ereg_reg[408]  ( .D(ereg_next[408]), .CLK(clk), .RST(rst), .I(e[408]), 
        .Q(ein[408]) );
  DFF \ereg_reg[409]  ( .D(ereg_next[409]), .CLK(clk), .RST(rst), .I(e[409]), 
        .Q(ein[409]) );
  DFF \ereg_reg[410]  ( .D(ereg_next[410]), .CLK(clk), .RST(rst), .I(e[410]), 
        .Q(ein[410]) );
  DFF \ereg_reg[411]  ( .D(ereg_next[411]), .CLK(clk), .RST(rst), .I(e[411]), 
        .Q(ein[411]) );
  DFF \ereg_reg[412]  ( .D(ereg_next[412]), .CLK(clk), .RST(rst), .I(e[412]), 
        .Q(ein[412]) );
  DFF \ereg_reg[413]  ( .D(ereg_next[413]), .CLK(clk), .RST(rst), .I(e[413]), 
        .Q(ein[413]) );
  DFF \ereg_reg[414]  ( .D(ereg_next[414]), .CLK(clk), .RST(rst), .I(e[414]), 
        .Q(ein[414]) );
  DFF \ereg_reg[415]  ( .D(ereg_next[415]), .CLK(clk), .RST(rst), .I(e[415]), 
        .Q(ein[415]) );
  DFF \ereg_reg[416]  ( .D(ereg_next[416]), .CLK(clk), .RST(rst), .I(e[416]), 
        .Q(ein[416]) );
  DFF \ereg_reg[417]  ( .D(ereg_next[417]), .CLK(clk), .RST(rst), .I(e[417]), 
        .Q(ein[417]) );
  DFF \ereg_reg[418]  ( .D(ereg_next[418]), .CLK(clk), .RST(rst), .I(e[418]), 
        .Q(ein[418]) );
  DFF \ereg_reg[419]  ( .D(ereg_next[419]), .CLK(clk), .RST(rst), .I(e[419]), 
        .Q(ein[419]) );
  DFF \ereg_reg[420]  ( .D(ereg_next[420]), .CLK(clk), .RST(rst), .I(e[420]), 
        .Q(ein[420]) );
  DFF \ereg_reg[421]  ( .D(ereg_next[421]), .CLK(clk), .RST(rst), .I(e[421]), 
        .Q(ein[421]) );
  DFF \ereg_reg[422]  ( .D(ereg_next[422]), .CLK(clk), .RST(rst), .I(e[422]), 
        .Q(ein[422]) );
  DFF \ereg_reg[423]  ( .D(ereg_next[423]), .CLK(clk), .RST(rst), .I(e[423]), 
        .Q(ein[423]) );
  DFF \ereg_reg[424]  ( .D(ereg_next[424]), .CLK(clk), .RST(rst), .I(e[424]), 
        .Q(ein[424]) );
  DFF \ereg_reg[425]  ( .D(ereg_next[425]), .CLK(clk), .RST(rst), .I(e[425]), 
        .Q(ein[425]) );
  DFF \ereg_reg[426]  ( .D(ereg_next[426]), .CLK(clk), .RST(rst), .I(e[426]), 
        .Q(ein[426]) );
  DFF \ereg_reg[427]  ( .D(ereg_next[427]), .CLK(clk), .RST(rst), .I(e[427]), 
        .Q(ein[427]) );
  DFF \ereg_reg[428]  ( .D(ereg_next[428]), .CLK(clk), .RST(rst), .I(e[428]), 
        .Q(ein[428]) );
  DFF \ereg_reg[429]  ( .D(ereg_next[429]), .CLK(clk), .RST(rst), .I(e[429]), 
        .Q(ein[429]) );
  DFF \ereg_reg[430]  ( .D(ereg_next[430]), .CLK(clk), .RST(rst), .I(e[430]), 
        .Q(ein[430]) );
  DFF \ereg_reg[431]  ( .D(ereg_next[431]), .CLK(clk), .RST(rst), .I(e[431]), 
        .Q(ein[431]) );
  DFF \ereg_reg[432]  ( .D(ereg_next[432]), .CLK(clk), .RST(rst), .I(e[432]), 
        .Q(ein[432]) );
  DFF \ereg_reg[433]  ( .D(ereg_next[433]), .CLK(clk), .RST(rst), .I(e[433]), 
        .Q(ein[433]) );
  DFF \ereg_reg[434]  ( .D(ereg_next[434]), .CLK(clk), .RST(rst), .I(e[434]), 
        .Q(ein[434]) );
  DFF \ereg_reg[435]  ( .D(ereg_next[435]), .CLK(clk), .RST(rst), .I(e[435]), 
        .Q(ein[435]) );
  DFF \ereg_reg[436]  ( .D(ereg_next[436]), .CLK(clk), .RST(rst), .I(e[436]), 
        .Q(ein[436]) );
  DFF \ereg_reg[437]  ( .D(ereg_next[437]), .CLK(clk), .RST(rst), .I(e[437]), 
        .Q(ein[437]) );
  DFF \ereg_reg[438]  ( .D(ereg_next[438]), .CLK(clk), .RST(rst), .I(e[438]), 
        .Q(ein[438]) );
  DFF \ereg_reg[439]  ( .D(ereg_next[439]), .CLK(clk), .RST(rst), .I(e[439]), 
        .Q(ein[439]) );
  DFF \ereg_reg[440]  ( .D(ereg_next[440]), .CLK(clk), .RST(rst), .I(e[440]), 
        .Q(ein[440]) );
  DFF \ereg_reg[441]  ( .D(ereg_next[441]), .CLK(clk), .RST(rst), .I(e[441]), 
        .Q(ein[441]) );
  DFF \ereg_reg[442]  ( .D(ereg_next[442]), .CLK(clk), .RST(rst), .I(e[442]), 
        .Q(ein[442]) );
  DFF \ereg_reg[443]  ( .D(ereg_next[443]), .CLK(clk), .RST(rst), .I(e[443]), 
        .Q(ein[443]) );
  DFF \ereg_reg[444]  ( .D(ereg_next[444]), .CLK(clk), .RST(rst), .I(e[444]), 
        .Q(ein[444]) );
  DFF \ereg_reg[445]  ( .D(ereg_next[445]), .CLK(clk), .RST(rst), .I(e[445]), 
        .Q(ein[445]) );
  DFF \ereg_reg[446]  ( .D(ereg_next[446]), .CLK(clk), .RST(rst), .I(e[446]), 
        .Q(ein[446]) );
  DFF \ereg_reg[447]  ( .D(ereg_next[447]), .CLK(clk), .RST(rst), .I(e[447]), 
        .Q(ein[447]) );
  DFF \ereg_reg[448]  ( .D(ereg_next[448]), .CLK(clk), .RST(rst), .I(e[448]), 
        .Q(ein[448]) );
  DFF \ereg_reg[449]  ( .D(ereg_next[449]), .CLK(clk), .RST(rst), .I(e[449]), 
        .Q(ein[449]) );
  DFF \ereg_reg[450]  ( .D(ereg_next[450]), .CLK(clk), .RST(rst), .I(e[450]), 
        .Q(ein[450]) );
  DFF \ereg_reg[451]  ( .D(ereg_next[451]), .CLK(clk), .RST(rst), .I(e[451]), 
        .Q(ein[451]) );
  DFF \ereg_reg[452]  ( .D(ereg_next[452]), .CLK(clk), .RST(rst), .I(e[452]), 
        .Q(ein[452]) );
  DFF \ereg_reg[453]  ( .D(ereg_next[453]), .CLK(clk), .RST(rst), .I(e[453]), 
        .Q(ein[453]) );
  DFF \ereg_reg[454]  ( .D(ereg_next[454]), .CLK(clk), .RST(rst), .I(e[454]), 
        .Q(ein[454]) );
  DFF \ereg_reg[455]  ( .D(ereg_next[455]), .CLK(clk), .RST(rst), .I(e[455]), 
        .Q(ein[455]) );
  DFF \ereg_reg[456]  ( .D(ereg_next[456]), .CLK(clk), .RST(rst), .I(e[456]), 
        .Q(ein[456]) );
  DFF \ereg_reg[457]  ( .D(ereg_next[457]), .CLK(clk), .RST(rst), .I(e[457]), 
        .Q(ein[457]) );
  DFF \ereg_reg[458]  ( .D(ereg_next[458]), .CLK(clk), .RST(rst), .I(e[458]), 
        .Q(ein[458]) );
  DFF \ereg_reg[459]  ( .D(ereg_next[459]), .CLK(clk), .RST(rst), .I(e[459]), 
        .Q(ein[459]) );
  DFF \ereg_reg[460]  ( .D(ereg_next[460]), .CLK(clk), .RST(rst), .I(e[460]), 
        .Q(ein[460]) );
  DFF \ereg_reg[461]  ( .D(ereg_next[461]), .CLK(clk), .RST(rst), .I(e[461]), 
        .Q(ein[461]) );
  DFF \ereg_reg[462]  ( .D(ereg_next[462]), .CLK(clk), .RST(rst), .I(e[462]), 
        .Q(ein[462]) );
  DFF \ereg_reg[463]  ( .D(ereg_next[463]), .CLK(clk), .RST(rst), .I(e[463]), 
        .Q(ein[463]) );
  DFF \ereg_reg[464]  ( .D(ereg_next[464]), .CLK(clk), .RST(rst), .I(e[464]), 
        .Q(ein[464]) );
  DFF \ereg_reg[465]  ( .D(ereg_next[465]), .CLK(clk), .RST(rst), .I(e[465]), 
        .Q(ein[465]) );
  DFF \ereg_reg[466]  ( .D(ereg_next[466]), .CLK(clk), .RST(rst), .I(e[466]), 
        .Q(ein[466]) );
  DFF \ereg_reg[467]  ( .D(ereg_next[467]), .CLK(clk), .RST(rst), .I(e[467]), 
        .Q(ein[467]) );
  DFF \ereg_reg[468]  ( .D(ereg_next[468]), .CLK(clk), .RST(rst), .I(e[468]), 
        .Q(ein[468]) );
  DFF \ereg_reg[469]  ( .D(ereg_next[469]), .CLK(clk), .RST(rst), .I(e[469]), 
        .Q(ein[469]) );
  DFF \ereg_reg[470]  ( .D(ereg_next[470]), .CLK(clk), .RST(rst), .I(e[470]), 
        .Q(ein[470]) );
  DFF \ereg_reg[471]  ( .D(ereg_next[471]), .CLK(clk), .RST(rst), .I(e[471]), 
        .Q(ein[471]) );
  DFF \ereg_reg[472]  ( .D(ereg_next[472]), .CLK(clk), .RST(rst), .I(e[472]), 
        .Q(ein[472]) );
  DFF \ereg_reg[473]  ( .D(ereg_next[473]), .CLK(clk), .RST(rst), .I(e[473]), 
        .Q(ein[473]) );
  DFF \ereg_reg[474]  ( .D(ereg_next[474]), .CLK(clk), .RST(rst), .I(e[474]), 
        .Q(ein[474]) );
  DFF \ereg_reg[475]  ( .D(ereg_next[475]), .CLK(clk), .RST(rst), .I(e[475]), 
        .Q(ein[475]) );
  DFF \ereg_reg[476]  ( .D(ereg_next[476]), .CLK(clk), .RST(rst), .I(e[476]), 
        .Q(ein[476]) );
  DFF \ereg_reg[477]  ( .D(ereg_next[477]), .CLK(clk), .RST(rst), .I(e[477]), 
        .Q(ein[477]) );
  DFF \ereg_reg[478]  ( .D(ereg_next[478]), .CLK(clk), .RST(rst), .I(e[478]), 
        .Q(ein[478]) );
  DFF \ereg_reg[479]  ( .D(ereg_next[479]), .CLK(clk), .RST(rst), .I(e[479]), 
        .Q(ein[479]) );
  DFF \ereg_reg[480]  ( .D(ereg_next[480]), .CLK(clk), .RST(rst), .I(e[480]), 
        .Q(ein[480]) );
  DFF \ereg_reg[481]  ( .D(ereg_next[481]), .CLK(clk), .RST(rst), .I(e[481]), 
        .Q(ein[481]) );
  DFF \ereg_reg[482]  ( .D(ereg_next[482]), .CLK(clk), .RST(rst), .I(e[482]), 
        .Q(ein[482]) );
  DFF \ereg_reg[483]  ( .D(ereg_next[483]), .CLK(clk), .RST(rst), .I(e[483]), 
        .Q(ein[483]) );
  DFF \ereg_reg[484]  ( .D(ereg_next[484]), .CLK(clk), .RST(rst), .I(e[484]), 
        .Q(ein[484]) );
  DFF \ereg_reg[485]  ( .D(ereg_next[485]), .CLK(clk), .RST(rst), .I(e[485]), 
        .Q(ein[485]) );
  DFF \ereg_reg[486]  ( .D(ereg_next[486]), .CLK(clk), .RST(rst), .I(e[486]), 
        .Q(ein[486]) );
  DFF \ereg_reg[487]  ( .D(ereg_next[487]), .CLK(clk), .RST(rst), .I(e[487]), 
        .Q(ein[487]) );
  DFF \ereg_reg[488]  ( .D(ereg_next[488]), .CLK(clk), .RST(rst), .I(e[488]), 
        .Q(ein[488]) );
  DFF \ereg_reg[489]  ( .D(ereg_next[489]), .CLK(clk), .RST(rst), .I(e[489]), 
        .Q(ein[489]) );
  DFF \ereg_reg[490]  ( .D(ereg_next[490]), .CLK(clk), .RST(rst), .I(e[490]), 
        .Q(ein[490]) );
  DFF \ereg_reg[491]  ( .D(ereg_next[491]), .CLK(clk), .RST(rst), .I(e[491]), 
        .Q(ein[491]) );
  DFF \ereg_reg[492]  ( .D(ereg_next[492]), .CLK(clk), .RST(rst), .I(e[492]), 
        .Q(ein[492]) );
  DFF \ereg_reg[493]  ( .D(ereg_next[493]), .CLK(clk), .RST(rst), .I(e[493]), 
        .Q(ein[493]) );
  DFF \ereg_reg[494]  ( .D(ereg_next[494]), .CLK(clk), .RST(rst), .I(e[494]), 
        .Q(ein[494]) );
  DFF \ereg_reg[495]  ( .D(ereg_next[495]), .CLK(clk), .RST(rst), .I(e[495]), 
        .Q(ein[495]) );
  DFF \ereg_reg[496]  ( .D(ereg_next[496]), .CLK(clk), .RST(rst), .I(e[496]), 
        .Q(ein[496]) );
  DFF \ereg_reg[497]  ( .D(ereg_next[497]), .CLK(clk), .RST(rst), .I(e[497]), 
        .Q(ein[497]) );
  DFF \ereg_reg[498]  ( .D(ereg_next[498]), .CLK(clk), .RST(rst), .I(e[498]), 
        .Q(ein[498]) );
  DFF \ereg_reg[499]  ( .D(ereg_next[499]), .CLK(clk), .RST(rst), .I(e[499]), 
        .Q(ein[499]) );
  DFF \ereg_reg[500]  ( .D(ereg_next[500]), .CLK(clk), .RST(rst), .I(e[500]), 
        .Q(ein[500]) );
  DFF \ereg_reg[501]  ( .D(ereg_next[501]), .CLK(clk), .RST(rst), .I(e[501]), 
        .Q(ein[501]) );
  DFF \ereg_reg[502]  ( .D(ereg_next[502]), .CLK(clk), .RST(rst), .I(e[502]), 
        .Q(ein[502]) );
  DFF \ereg_reg[503]  ( .D(ereg_next[503]), .CLK(clk), .RST(rst), .I(e[503]), 
        .Q(ein[503]) );
  DFF \ereg_reg[504]  ( .D(ereg_next[504]), .CLK(clk), .RST(rst), .I(e[504]), 
        .Q(ein[504]) );
  DFF \ereg_reg[505]  ( .D(ereg_next[505]), .CLK(clk), .RST(rst), .I(e[505]), 
        .Q(ein[505]) );
  DFF \ereg_reg[506]  ( .D(ereg_next[506]), .CLK(clk), .RST(rst), .I(e[506]), 
        .Q(ein[506]) );
  DFF \ereg_reg[507]  ( .D(ereg_next[507]), .CLK(clk), .RST(rst), .I(e[507]), 
        .Q(ein[507]) );
  DFF \ereg_reg[508]  ( .D(ereg_next[508]), .CLK(clk), .RST(rst), .I(e[508]), 
        .Q(ein[508]) );
  DFF \ereg_reg[509]  ( .D(ereg_next[509]), .CLK(clk), .RST(rst), .I(e[509]), 
        .Q(ein[509]) );
  DFF \ereg_reg[510]  ( .D(ereg_next[510]), .CLK(clk), .RST(rst), .I(e[510]), 
        .Q(ein[510]) );
  DFF \ereg_reg[511]  ( .D(ereg_next[511]), .CLK(clk), .RST(rst), .I(e[511]), 
        .Q(ein[511]) );
  DFF \ereg_reg[512]  ( .D(ereg_next[512]), .CLK(clk), .RST(rst), .I(e[512]), 
        .Q(ein[512]) );
  DFF \ereg_reg[513]  ( .D(ereg_next[513]), .CLK(clk), .RST(rst), .I(e[513]), 
        .Q(ein[513]) );
  DFF \ereg_reg[514]  ( .D(ereg_next[514]), .CLK(clk), .RST(rst), .I(e[514]), 
        .Q(ein[514]) );
  DFF \ereg_reg[515]  ( .D(ereg_next[515]), .CLK(clk), .RST(rst), .I(e[515]), 
        .Q(ein[515]) );
  DFF \ereg_reg[516]  ( .D(ereg_next[516]), .CLK(clk), .RST(rst), .I(e[516]), 
        .Q(ein[516]) );
  DFF \ereg_reg[517]  ( .D(ereg_next[517]), .CLK(clk), .RST(rst), .I(e[517]), 
        .Q(ein[517]) );
  DFF \ereg_reg[518]  ( .D(ereg_next[518]), .CLK(clk), .RST(rst), .I(e[518]), 
        .Q(ein[518]) );
  DFF \ereg_reg[519]  ( .D(ereg_next[519]), .CLK(clk), .RST(rst), .I(e[519]), 
        .Q(ein[519]) );
  DFF \ereg_reg[520]  ( .D(ereg_next[520]), .CLK(clk), .RST(rst), .I(e[520]), 
        .Q(ein[520]) );
  DFF \ereg_reg[521]  ( .D(ereg_next[521]), .CLK(clk), .RST(rst), .I(e[521]), 
        .Q(ein[521]) );
  DFF \ereg_reg[522]  ( .D(ereg_next[522]), .CLK(clk), .RST(rst), .I(e[522]), 
        .Q(ein[522]) );
  DFF \ereg_reg[523]  ( .D(ereg_next[523]), .CLK(clk), .RST(rst), .I(e[523]), 
        .Q(ein[523]) );
  DFF \ereg_reg[524]  ( .D(ereg_next[524]), .CLK(clk), .RST(rst), .I(e[524]), 
        .Q(ein[524]) );
  DFF \ereg_reg[525]  ( .D(ereg_next[525]), .CLK(clk), .RST(rst), .I(e[525]), 
        .Q(ein[525]) );
  DFF \ereg_reg[526]  ( .D(ereg_next[526]), .CLK(clk), .RST(rst), .I(e[526]), 
        .Q(ein[526]) );
  DFF \ereg_reg[527]  ( .D(ereg_next[527]), .CLK(clk), .RST(rst), .I(e[527]), 
        .Q(ein[527]) );
  DFF \ereg_reg[528]  ( .D(ereg_next[528]), .CLK(clk), .RST(rst), .I(e[528]), 
        .Q(ein[528]) );
  DFF \ereg_reg[529]  ( .D(ereg_next[529]), .CLK(clk), .RST(rst), .I(e[529]), 
        .Q(ein[529]) );
  DFF \ereg_reg[530]  ( .D(ereg_next[530]), .CLK(clk), .RST(rst), .I(e[530]), 
        .Q(ein[530]) );
  DFF \ereg_reg[531]  ( .D(ereg_next[531]), .CLK(clk), .RST(rst), .I(e[531]), 
        .Q(ein[531]) );
  DFF \ereg_reg[532]  ( .D(ereg_next[532]), .CLK(clk), .RST(rst), .I(e[532]), 
        .Q(ein[532]) );
  DFF \ereg_reg[533]  ( .D(ereg_next[533]), .CLK(clk), .RST(rst), .I(e[533]), 
        .Q(ein[533]) );
  DFF \ereg_reg[534]  ( .D(ereg_next[534]), .CLK(clk), .RST(rst), .I(e[534]), 
        .Q(ein[534]) );
  DFF \ereg_reg[535]  ( .D(ereg_next[535]), .CLK(clk), .RST(rst), .I(e[535]), 
        .Q(ein[535]) );
  DFF \ereg_reg[536]  ( .D(ereg_next[536]), .CLK(clk), .RST(rst), .I(e[536]), 
        .Q(ein[536]) );
  DFF \ereg_reg[537]  ( .D(ereg_next[537]), .CLK(clk), .RST(rst), .I(e[537]), 
        .Q(ein[537]) );
  DFF \ereg_reg[538]  ( .D(ereg_next[538]), .CLK(clk), .RST(rst), .I(e[538]), 
        .Q(ein[538]) );
  DFF \ereg_reg[539]  ( .D(ereg_next[539]), .CLK(clk), .RST(rst), .I(e[539]), 
        .Q(ein[539]) );
  DFF \ereg_reg[540]  ( .D(ereg_next[540]), .CLK(clk), .RST(rst), .I(e[540]), 
        .Q(ein[540]) );
  DFF \ereg_reg[541]  ( .D(ereg_next[541]), .CLK(clk), .RST(rst), .I(e[541]), 
        .Q(ein[541]) );
  DFF \ereg_reg[542]  ( .D(ereg_next[542]), .CLK(clk), .RST(rst), .I(e[542]), 
        .Q(ein[542]) );
  DFF \ereg_reg[543]  ( .D(ereg_next[543]), .CLK(clk), .RST(rst), .I(e[543]), 
        .Q(ein[543]) );
  DFF \ereg_reg[544]  ( .D(ereg_next[544]), .CLK(clk), .RST(rst), .I(e[544]), 
        .Q(ein[544]) );
  DFF \ereg_reg[545]  ( .D(ereg_next[545]), .CLK(clk), .RST(rst), .I(e[545]), 
        .Q(ein[545]) );
  DFF \ereg_reg[546]  ( .D(ereg_next[546]), .CLK(clk), .RST(rst), .I(e[546]), 
        .Q(ein[546]) );
  DFF \ereg_reg[547]  ( .D(ereg_next[547]), .CLK(clk), .RST(rst), .I(e[547]), 
        .Q(ein[547]) );
  DFF \ereg_reg[548]  ( .D(ereg_next[548]), .CLK(clk), .RST(rst), .I(e[548]), 
        .Q(ein[548]) );
  DFF \ereg_reg[549]  ( .D(ereg_next[549]), .CLK(clk), .RST(rst), .I(e[549]), 
        .Q(ein[549]) );
  DFF \ereg_reg[550]  ( .D(ereg_next[550]), .CLK(clk), .RST(rst), .I(e[550]), 
        .Q(ein[550]) );
  DFF \ereg_reg[551]  ( .D(ereg_next[551]), .CLK(clk), .RST(rst), .I(e[551]), 
        .Q(ein[551]) );
  DFF \ereg_reg[552]  ( .D(ereg_next[552]), .CLK(clk), .RST(rst), .I(e[552]), 
        .Q(ein[552]) );
  DFF \ereg_reg[553]  ( .D(ereg_next[553]), .CLK(clk), .RST(rst), .I(e[553]), 
        .Q(ein[553]) );
  DFF \ereg_reg[554]  ( .D(ereg_next[554]), .CLK(clk), .RST(rst), .I(e[554]), 
        .Q(ein[554]) );
  DFF \ereg_reg[555]  ( .D(ereg_next[555]), .CLK(clk), .RST(rst), .I(e[555]), 
        .Q(ein[555]) );
  DFF \ereg_reg[556]  ( .D(ereg_next[556]), .CLK(clk), .RST(rst), .I(e[556]), 
        .Q(ein[556]) );
  DFF \ereg_reg[557]  ( .D(ereg_next[557]), .CLK(clk), .RST(rst), .I(e[557]), 
        .Q(ein[557]) );
  DFF \ereg_reg[558]  ( .D(ereg_next[558]), .CLK(clk), .RST(rst), .I(e[558]), 
        .Q(ein[558]) );
  DFF \ereg_reg[559]  ( .D(ereg_next[559]), .CLK(clk), .RST(rst), .I(e[559]), 
        .Q(ein[559]) );
  DFF \ereg_reg[560]  ( .D(ereg_next[560]), .CLK(clk), .RST(rst), .I(e[560]), 
        .Q(ein[560]) );
  DFF \ereg_reg[561]  ( .D(ereg_next[561]), .CLK(clk), .RST(rst), .I(e[561]), 
        .Q(ein[561]) );
  DFF \ereg_reg[562]  ( .D(ereg_next[562]), .CLK(clk), .RST(rst), .I(e[562]), 
        .Q(ein[562]) );
  DFF \ereg_reg[563]  ( .D(ereg_next[563]), .CLK(clk), .RST(rst), .I(e[563]), 
        .Q(ein[563]) );
  DFF \ereg_reg[564]  ( .D(ereg_next[564]), .CLK(clk), .RST(rst), .I(e[564]), 
        .Q(ein[564]) );
  DFF \ereg_reg[565]  ( .D(ereg_next[565]), .CLK(clk), .RST(rst), .I(e[565]), 
        .Q(ein[565]) );
  DFF \ereg_reg[566]  ( .D(ereg_next[566]), .CLK(clk), .RST(rst), .I(e[566]), 
        .Q(ein[566]) );
  DFF \ereg_reg[567]  ( .D(ereg_next[567]), .CLK(clk), .RST(rst), .I(e[567]), 
        .Q(ein[567]) );
  DFF \ereg_reg[568]  ( .D(ereg_next[568]), .CLK(clk), .RST(rst), .I(e[568]), 
        .Q(ein[568]) );
  DFF \ereg_reg[569]  ( .D(ereg_next[569]), .CLK(clk), .RST(rst), .I(e[569]), 
        .Q(ein[569]) );
  DFF \ereg_reg[570]  ( .D(ereg_next[570]), .CLK(clk), .RST(rst), .I(e[570]), 
        .Q(ein[570]) );
  DFF \ereg_reg[571]  ( .D(ereg_next[571]), .CLK(clk), .RST(rst), .I(e[571]), 
        .Q(ein[571]) );
  DFF \ereg_reg[572]  ( .D(ereg_next[572]), .CLK(clk), .RST(rst), .I(e[572]), 
        .Q(ein[572]) );
  DFF \ereg_reg[573]  ( .D(ereg_next[573]), .CLK(clk), .RST(rst), .I(e[573]), 
        .Q(ein[573]) );
  DFF \ereg_reg[574]  ( .D(ereg_next[574]), .CLK(clk), .RST(rst), .I(e[574]), 
        .Q(ein[574]) );
  DFF \ereg_reg[575]  ( .D(ereg_next[575]), .CLK(clk), .RST(rst), .I(e[575]), 
        .Q(ein[575]) );
  DFF \ereg_reg[576]  ( .D(ereg_next[576]), .CLK(clk), .RST(rst), .I(e[576]), 
        .Q(ein[576]) );
  DFF \ereg_reg[577]  ( .D(ereg_next[577]), .CLK(clk), .RST(rst), .I(e[577]), 
        .Q(ein[577]) );
  DFF \ereg_reg[578]  ( .D(ereg_next[578]), .CLK(clk), .RST(rst), .I(e[578]), 
        .Q(ein[578]) );
  DFF \ereg_reg[579]  ( .D(ereg_next[579]), .CLK(clk), .RST(rst), .I(e[579]), 
        .Q(ein[579]) );
  DFF \ereg_reg[580]  ( .D(ereg_next[580]), .CLK(clk), .RST(rst), .I(e[580]), 
        .Q(ein[580]) );
  DFF \ereg_reg[581]  ( .D(ereg_next[581]), .CLK(clk), .RST(rst), .I(e[581]), 
        .Q(ein[581]) );
  DFF \ereg_reg[582]  ( .D(ereg_next[582]), .CLK(clk), .RST(rst), .I(e[582]), 
        .Q(ein[582]) );
  DFF \ereg_reg[583]  ( .D(ereg_next[583]), .CLK(clk), .RST(rst), .I(e[583]), 
        .Q(ein[583]) );
  DFF \ereg_reg[584]  ( .D(ereg_next[584]), .CLK(clk), .RST(rst), .I(e[584]), 
        .Q(ein[584]) );
  DFF \ereg_reg[585]  ( .D(ereg_next[585]), .CLK(clk), .RST(rst), .I(e[585]), 
        .Q(ein[585]) );
  DFF \ereg_reg[586]  ( .D(ereg_next[586]), .CLK(clk), .RST(rst), .I(e[586]), 
        .Q(ein[586]) );
  DFF \ereg_reg[587]  ( .D(ereg_next[587]), .CLK(clk), .RST(rst), .I(e[587]), 
        .Q(ein[587]) );
  DFF \ereg_reg[588]  ( .D(ereg_next[588]), .CLK(clk), .RST(rst), .I(e[588]), 
        .Q(ein[588]) );
  DFF \ereg_reg[589]  ( .D(ereg_next[589]), .CLK(clk), .RST(rst), .I(e[589]), 
        .Q(ein[589]) );
  DFF \ereg_reg[590]  ( .D(ereg_next[590]), .CLK(clk), .RST(rst), .I(e[590]), 
        .Q(ein[590]) );
  DFF \ereg_reg[591]  ( .D(ereg_next[591]), .CLK(clk), .RST(rst), .I(e[591]), 
        .Q(ein[591]) );
  DFF \ereg_reg[592]  ( .D(ereg_next[592]), .CLK(clk), .RST(rst), .I(e[592]), 
        .Q(ein[592]) );
  DFF \ereg_reg[593]  ( .D(ereg_next[593]), .CLK(clk), .RST(rst), .I(e[593]), 
        .Q(ein[593]) );
  DFF \ereg_reg[594]  ( .D(ereg_next[594]), .CLK(clk), .RST(rst), .I(e[594]), 
        .Q(ein[594]) );
  DFF \ereg_reg[595]  ( .D(ereg_next[595]), .CLK(clk), .RST(rst), .I(e[595]), 
        .Q(ein[595]) );
  DFF \ereg_reg[596]  ( .D(ereg_next[596]), .CLK(clk), .RST(rst), .I(e[596]), 
        .Q(ein[596]) );
  DFF \ereg_reg[597]  ( .D(ereg_next[597]), .CLK(clk), .RST(rst), .I(e[597]), 
        .Q(ein[597]) );
  DFF \ereg_reg[598]  ( .D(ereg_next[598]), .CLK(clk), .RST(rst), .I(e[598]), 
        .Q(ein[598]) );
  DFF \ereg_reg[599]  ( .D(ereg_next[599]), .CLK(clk), .RST(rst), .I(e[599]), 
        .Q(ein[599]) );
  DFF \ereg_reg[600]  ( .D(ereg_next[600]), .CLK(clk), .RST(rst), .I(e[600]), 
        .Q(ein[600]) );
  DFF \ereg_reg[601]  ( .D(ereg_next[601]), .CLK(clk), .RST(rst), .I(e[601]), 
        .Q(ein[601]) );
  DFF \ereg_reg[602]  ( .D(ereg_next[602]), .CLK(clk), .RST(rst), .I(e[602]), 
        .Q(ein[602]) );
  DFF \ereg_reg[603]  ( .D(ereg_next[603]), .CLK(clk), .RST(rst), .I(e[603]), 
        .Q(ein[603]) );
  DFF \ereg_reg[604]  ( .D(ereg_next[604]), .CLK(clk), .RST(rst), .I(e[604]), 
        .Q(ein[604]) );
  DFF \ereg_reg[605]  ( .D(ereg_next[605]), .CLK(clk), .RST(rst), .I(e[605]), 
        .Q(ein[605]) );
  DFF \ereg_reg[606]  ( .D(ereg_next[606]), .CLK(clk), .RST(rst), .I(e[606]), 
        .Q(ein[606]) );
  DFF \ereg_reg[607]  ( .D(ereg_next[607]), .CLK(clk), .RST(rst), .I(e[607]), 
        .Q(ein[607]) );
  DFF \ereg_reg[608]  ( .D(ereg_next[608]), .CLK(clk), .RST(rst), .I(e[608]), 
        .Q(ein[608]) );
  DFF \ereg_reg[609]  ( .D(ereg_next[609]), .CLK(clk), .RST(rst), .I(e[609]), 
        .Q(ein[609]) );
  DFF \ereg_reg[610]  ( .D(ereg_next[610]), .CLK(clk), .RST(rst), .I(e[610]), 
        .Q(ein[610]) );
  DFF \ereg_reg[611]  ( .D(ereg_next[611]), .CLK(clk), .RST(rst), .I(e[611]), 
        .Q(ein[611]) );
  DFF \ereg_reg[612]  ( .D(ereg_next[612]), .CLK(clk), .RST(rst), .I(e[612]), 
        .Q(ein[612]) );
  DFF \ereg_reg[613]  ( .D(ereg_next[613]), .CLK(clk), .RST(rst), .I(e[613]), 
        .Q(ein[613]) );
  DFF \ereg_reg[614]  ( .D(ereg_next[614]), .CLK(clk), .RST(rst), .I(e[614]), 
        .Q(ein[614]) );
  DFF \ereg_reg[615]  ( .D(ereg_next[615]), .CLK(clk), .RST(rst), .I(e[615]), 
        .Q(ein[615]) );
  DFF \ereg_reg[616]  ( .D(ereg_next[616]), .CLK(clk), .RST(rst), .I(e[616]), 
        .Q(ein[616]) );
  DFF \ereg_reg[617]  ( .D(ereg_next[617]), .CLK(clk), .RST(rst), .I(e[617]), 
        .Q(ein[617]) );
  DFF \ereg_reg[618]  ( .D(ereg_next[618]), .CLK(clk), .RST(rst), .I(e[618]), 
        .Q(ein[618]) );
  DFF \ereg_reg[619]  ( .D(ereg_next[619]), .CLK(clk), .RST(rst), .I(e[619]), 
        .Q(ein[619]) );
  DFF \ereg_reg[620]  ( .D(ereg_next[620]), .CLK(clk), .RST(rst), .I(e[620]), 
        .Q(ein[620]) );
  DFF \ereg_reg[621]  ( .D(ereg_next[621]), .CLK(clk), .RST(rst), .I(e[621]), 
        .Q(ein[621]) );
  DFF \ereg_reg[622]  ( .D(ereg_next[622]), .CLK(clk), .RST(rst), .I(e[622]), 
        .Q(ein[622]) );
  DFF \ereg_reg[623]  ( .D(ereg_next[623]), .CLK(clk), .RST(rst), .I(e[623]), 
        .Q(ein[623]) );
  DFF \ereg_reg[624]  ( .D(ereg_next[624]), .CLK(clk), .RST(rst), .I(e[624]), 
        .Q(ein[624]) );
  DFF \ereg_reg[625]  ( .D(ereg_next[625]), .CLK(clk), .RST(rst), .I(e[625]), 
        .Q(ein[625]) );
  DFF \ereg_reg[626]  ( .D(ereg_next[626]), .CLK(clk), .RST(rst), .I(e[626]), 
        .Q(ein[626]) );
  DFF \ereg_reg[627]  ( .D(ereg_next[627]), .CLK(clk), .RST(rst), .I(e[627]), 
        .Q(ein[627]) );
  DFF \ereg_reg[628]  ( .D(ereg_next[628]), .CLK(clk), .RST(rst), .I(e[628]), 
        .Q(ein[628]) );
  DFF \ereg_reg[629]  ( .D(ereg_next[629]), .CLK(clk), .RST(rst), .I(e[629]), 
        .Q(ein[629]) );
  DFF \ereg_reg[630]  ( .D(ereg_next[630]), .CLK(clk), .RST(rst), .I(e[630]), 
        .Q(ein[630]) );
  DFF \ereg_reg[631]  ( .D(ereg_next[631]), .CLK(clk), .RST(rst), .I(e[631]), 
        .Q(ein[631]) );
  DFF \ereg_reg[632]  ( .D(ereg_next[632]), .CLK(clk), .RST(rst), .I(e[632]), 
        .Q(ein[632]) );
  DFF \ereg_reg[633]  ( .D(ereg_next[633]), .CLK(clk), .RST(rst), .I(e[633]), 
        .Q(ein[633]) );
  DFF \ereg_reg[634]  ( .D(ereg_next[634]), .CLK(clk), .RST(rst), .I(e[634]), 
        .Q(ein[634]) );
  DFF \ereg_reg[635]  ( .D(ereg_next[635]), .CLK(clk), .RST(rst), .I(e[635]), 
        .Q(ein[635]) );
  DFF \ereg_reg[636]  ( .D(ereg_next[636]), .CLK(clk), .RST(rst), .I(e[636]), 
        .Q(ein[636]) );
  DFF \ereg_reg[637]  ( .D(ereg_next[637]), .CLK(clk), .RST(rst), .I(e[637]), 
        .Q(ein[637]) );
  DFF \ereg_reg[638]  ( .D(ereg_next[638]), .CLK(clk), .RST(rst), .I(e[638]), 
        .Q(ein[638]) );
  DFF \ereg_reg[639]  ( .D(ereg_next[639]), .CLK(clk), .RST(rst), .I(e[639]), 
        .Q(ein[639]) );
  DFF \ereg_reg[640]  ( .D(ereg_next[640]), .CLK(clk), .RST(rst), .I(e[640]), 
        .Q(ein[640]) );
  DFF \ereg_reg[641]  ( .D(ereg_next[641]), .CLK(clk), .RST(rst), .I(e[641]), 
        .Q(ein[641]) );
  DFF \ereg_reg[642]  ( .D(ereg_next[642]), .CLK(clk), .RST(rst), .I(e[642]), 
        .Q(ein[642]) );
  DFF \ereg_reg[643]  ( .D(ereg_next[643]), .CLK(clk), .RST(rst), .I(e[643]), 
        .Q(ein[643]) );
  DFF \ereg_reg[644]  ( .D(ereg_next[644]), .CLK(clk), .RST(rst), .I(e[644]), 
        .Q(ein[644]) );
  DFF \ereg_reg[645]  ( .D(ereg_next[645]), .CLK(clk), .RST(rst), .I(e[645]), 
        .Q(ein[645]) );
  DFF \ereg_reg[646]  ( .D(ereg_next[646]), .CLK(clk), .RST(rst), .I(e[646]), 
        .Q(ein[646]) );
  DFF \ereg_reg[647]  ( .D(ereg_next[647]), .CLK(clk), .RST(rst), .I(e[647]), 
        .Q(ein[647]) );
  DFF \ereg_reg[648]  ( .D(ereg_next[648]), .CLK(clk), .RST(rst), .I(e[648]), 
        .Q(ein[648]) );
  DFF \ereg_reg[649]  ( .D(ereg_next[649]), .CLK(clk), .RST(rst), .I(e[649]), 
        .Q(ein[649]) );
  DFF \ereg_reg[650]  ( .D(ereg_next[650]), .CLK(clk), .RST(rst), .I(e[650]), 
        .Q(ein[650]) );
  DFF \ereg_reg[651]  ( .D(ereg_next[651]), .CLK(clk), .RST(rst), .I(e[651]), 
        .Q(ein[651]) );
  DFF \ereg_reg[652]  ( .D(ereg_next[652]), .CLK(clk), .RST(rst), .I(e[652]), 
        .Q(ein[652]) );
  DFF \ereg_reg[653]  ( .D(ereg_next[653]), .CLK(clk), .RST(rst), .I(e[653]), 
        .Q(ein[653]) );
  DFF \ereg_reg[654]  ( .D(ereg_next[654]), .CLK(clk), .RST(rst), .I(e[654]), 
        .Q(ein[654]) );
  DFF \ereg_reg[655]  ( .D(ereg_next[655]), .CLK(clk), .RST(rst), .I(e[655]), 
        .Q(ein[655]) );
  DFF \ereg_reg[656]  ( .D(ereg_next[656]), .CLK(clk), .RST(rst), .I(e[656]), 
        .Q(ein[656]) );
  DFF \ereg_reg[657]  ( .D(ereg_next[657]), .CLK(clk), .RST(rst), .I(e[657]), 
        .Q(ein[657]) );
  DFF \ereg_reg[658]  ( .D(ereg_next[658]), .CLK(clk), .RST(rst), .I(e[658]), 
        .Q(ein[658]) );
  DFF \ereg_reg[659]  ( .D(ereg_next[659]), .CLK(clk), .RST(rst), .I(e[659]), 
        .Q(ein[659]) );
  DFF \ereg_reg[660]  ( .D(ereg_next[660]), .CLK(clk), .RST(rst), .I(e[660]), 
        .Q(ein[660]) );
  DFF \ereg_reg[661]  ( .D(ereg_next[661]), .CLK(clk), .RST(rst), .I(e[661]), 
        .Q(ein[661]) );
  DFF \ereg_reg[662]  ( .D(ereg_next[662]), .CLK(clk), .RST(rst), .I(e[662]), 
        .Q(ein[662]) );
  DFF \ereg_reg[663]  ( .D(ereg_next[663]), .CLK(clk), .RST(rst), .I(e[663]), 
        .Q(ein[663]) );
  DFF \ereg_reg[664]  ( .D(ereg_next[664]), .CLK(clk), .RST(rst), .I(e[664]), 
        .Q(ein[664]) );
  DFF \ereg_reg[665]  ( .D(ereg_next[665]), .CLK(clk), .RST(rst), .I(e[665]), 
        .Q(ein[665]) );
  DFF \ereg_reg[666]  ( .D(ereg_next[666]), .CLK(clk), .RST(rst), .I(e[666]), 
        .Q(ein[666]) );
  DFF \ereg_reg[667]  ( .D(ereg_next[667]), .CLK(clk), .RST(rst), .I(e[667]), 
        .Q(ein[667]) );
  DFF \ereg_reg[668]  ( .D(ereg_next[668]), .CLK(clk), .RST(rst), .I(e[668]), 
        .Q(ein[668]) );
  DFF \ereg_reg[669]  ( .D(ereg_next[669]), .CLK(clk), .RST(rst), .I(e[669]), 
        .Q(ein[669]) );
  DFF \ereg_reg[670]  ( .D(ereg_next[670]), .CLK(clk), .RST(rst), .I(e[670]), 
        .Q(ein[670]) );
  DFF \ereg_reg[671]  ( .D(ereg_next[671]), .CLK(clk), .RST(rst), .I(e[671]), 
        .Q(ein[671]) );
  DFF \ereg_reg[672]  ( .D(ereg_next[672]), .CLK(clk), .RST(rst), .I(e[672]), 
        .Q(ein[672]) );
  DFF \ereg_reg[673]  ( .D(ereg_next[673]), .CLK(clk), .RST(rst), .I(e[673]), 
        .Q(ein[673]) );
  DFF \ereg_reg[674]  ( .D(ereg_next[674]), .CLK(clk), .RST(rst), .I(e[674]), 
        .Q(ein[674]) );
  DFF \ereg_reg[675]  ( .D(ereg_next[675]), .CLK(clk), .RST(rst), .I(e[675]), 
        .Q(ein[675]) );
  DFF \ereg_reg[676]  ( .D(ereg_next[676]), .CLK(clk), .RST(rst), .I(e[676]), 
        .Q(ein[676]) );
  DFF \ereg_reg[677]  ( .D(ereg_next[677]), .CLK(clk), .RST(rst), .I(e[677]), 
        .Q(ein[677]) );
  DFF \ereg_reg[678]  ( .D(ereg_next[678]), .CLK(clk), .RST(rst), .I(e[678]), 
        .Q(ein[678]) );
  DFF \ereg_reg[679]  ( .D(ereg_next[679]), .CLK(clk), .RST(rst), .I(e[679]), 
        .Q(ein[679]) );
  DFF \ereg_reg[680]  ( .D(ereg_next[680]), .CLK(clk), .RST(rst), .I(e[680]), 
        .Q(ein[680]) );
  DFF \ereg_reg[681]  ( .D(ereg_next[681]), .CLK(clk), .RST(rst), .I(e[681]), 
        .Q(ein[681]) );
  DFF \ereg_reg[682]  ( .D(ereg_next[682]), .CLK(clk), .RST(rst), .I(e[682]), 
        .Q(ein[682]) );
  DFF \ereg_reg[683]  ( .D(ereg_next[683]), .CLK(clk), .RST(rst), .I(e[683]), 
        .Q(ein[683]) );
  DFF \ereg_reg[684]  ( .D(ereg_next[684]), .CLK(clk), .RST(rst), .I(e[684]), 
        .Q(ein[684]) );
  DFF \ereg_reg[685]  ( .D(ereg_next[685]), .CLK(clk), .RST(rst), .I(e[685]), 
        .Q(ein[685]) );
  DFF \ereg_reg[686]  ( .D(ereg_next[686]), .CLK(clk), .RST(rst), .I(e[686]), 
        .Q(ein[686]) );
  DFF \ereg_reg[687]  ( .D(ereg_next[687]), .CLK(clk), .RST(rst), .I(e[687]), 
        .Q(ein[687]) );
  DFF \ereg_reg[688]  ( .D(ereg_next[688]), .CLK(clk), .RST(rst), .I(e[688]), 
        .Q(ein[688]) );
  DFF \ereg_reg[689]  ( .D(ereg_next[689]), .CLK(clk), .RST(rst), .I(e[689]), 
        .Q(ein[689]) );
  DFF \ereg_reg[690]  ( .D(ereg_next[690]), .CLK(clk), .RST(rst), .I(e[690]), 
        .Q(ein[690]) );
  DFF \ereg_reg[691]  ( .D(ereg_next[691]), .CLK(clk), .RST(rst), .I(e[691]), 
        .Q(ein[691]) );
  DFF \ereg_reg[692]  ( .D(ereg_next[692]), .CLK(clk), .RST(rst), .I(e[692]), 
        .Q(ein[692]) );
  DFF \ereg_reg[693]  ( .D(ereg_next[693]), .CLK(clk), .RST(rst), .I(e[693]), 
        .Q(ein[693]) );
  DFF \ereg_reg[694]  ( .D(ereg_next[694]), .CLK(clk), .RST(rst), .I(e[694]), 
        .Q(ein[694]) );
  DFF \ereg_reg[695]  ( .D(ereg_next[695]), .CLK(clk), .RST(rst), .I(e[695]), 
        .Q(ein[695]) );
  DFF \ereg_reg[696]  ( .D(ereg_next[696]), .CLK(clk), .RST(rst), .I(e[696]), 
        .Q(ein[696]) );
  DFF \ereg_reg[697]  ( .D(ereg_next[697]), .CLK(clk), .RST(rst), .I(e[697]), 
        .Q(ein[697]) );
  DFF \ereg_reg[698]  ( .D(ereg_next[698]), .CLK(clk), .RST(rst), .I(e[698]), 
        .Q(ein[698]) );
  DFF \ereg_reg[699]  ( .D(ereg_next[699]), .CLK(clk), .RST(rst), .I(e[699]), 
        .Q(ein[699]) );
  DFF \ereg_reg[700]  ( .D(ereg_next[700]), .CLK(clk), .RST(rst), .I(e[700]), 
        .Q(ein[700]) );
  DFF \ereg_reg[701]  ( .D(ereg_next[701]), .CLK(clk), .RST(rst), .I(e[701]), 
        .Q(ein[701]) );
  DFF \ereg_reg[702]  ( .D(ereg_next[702]), .CLK(clk), .RST(rst), .I(e[702]), 
        .Q(ein[702]) );
  DFF \ereg_reg[703]  ( .D(ereg_next[703]), .CLK(clk), .RST(rst), .I(e[703]), 
        .Q(ein[703]) );
  DFF \ereg_reg[704]  ( .D(ereg_next[704]), .CLK(clk), .RST(rst), .I(e[704]), 
        .Q(ein[704]) );
  DFF \ereg_reg[705]  ( .D(ereg_next[705]), .CLK(clk), .RST(rst), .I(e[705]), 
        .Q(ein[705]) );
  DFF \ereg_reg[706]  ( .D(ereg_next[706]), .CLK(clk), .RST(rst), .I(e[706]), 
        .Q(ein[706]) );
  DFF \ereg_reg[707]  ( .D(ereg_next[707]), .CLK(clk), .RST(rst), .I(e[707]), 
        .Q(ein[707]) );
  DFF \ereg_reg[708]  ( .D(ereg_next[708]), .CLK(clk), .RST(rst), .I(e[708]), 
        .Q(ein[708]) );
  DFF \ereg_reg[709]  ( .D(ereg_next[709]), .CLK(clk), .RST(rst), .I(e[709]), 
        .Q(ein[709]) );
  DFF \ereg_reg[710]  ( .D(ereg_next[710]), .CLK(clk), .RST(rst), .I(e[710]), 
        .Q(ein[710]) );
  DFF \ereg_reg[711]  ( .D(ereg_next[711]), .CLK(clk), .RST(rst), .I(e[711]), 
        .Q(ein[711]) );
  DFF \ereg_reg[712]  ( .D(ereg_next[712]), .CLK(clk), .RST(rst), .I(e[712]), 
        .Q(ein[712]) );
  DFF \ereg_reg[713]  ( .D(ereg_next[713]), .CLK(clk), .RST(rst), .I(e[713]), 
        .Q(ein[713]) );
  DFF \ereg_reg[714]  ( .D(ereg_next[714]), .CLK(clk), .RST(rst), .I(e[714]), 
        .Q(ein[714]) );
  DFF \ereg_reg[715]  ( .D(ereg_next[715]), .CLK(clk), .RST(rst), .I(e[715]), 
        .Q(ein[715]) );
  DFF \ereg_reg[716]  ( .D(ereg_next[716]), .CLK(clk), .RST(rst), .I(e[716]), 
        .Q(ein[716]) );
  DFF \ereg_reg[717]  ( .D(ereg_next[717]), .CLK(clk), .RST(rst), .I(e[717]), 
        .Q(ein[717]) );
  DFF \ereg_reg[718]  ( .D(ereg_next[718]), .CLK(clk), .RST(rst), .I(e[718]), 
        .Q(ein[718]) );
  DFF \ereg_reg[719]  ( .D(ereg_next[719]), .CLK(clk), .RST(rst), .I(e[719]), 
        .Q(ein[719]) );
  DFF \ereg_reg[720]  ( .D(ereg_next[720]), .CLK(clk), .RST(rst), .I(e[720]), 
        .Q(ein[720]) );
  DFF \ereg_reg[721]  ( .D(ereg_next[721]), .CLK(clk), .RST(rst), .I(e[721]), 
        .Q(ein[721]) );
  DFF \ereg_reg[722]  ( .D(ereg_next[722]), .CLK(clk), .RST(rst), .I(e[722]), 
        .Q(ein[722]) );
  DFF \ereg_reg[723]  ( .D(ereg_next[723]), .CLK(clk), .RST(rst), .I(e[723]), 
        .Q(ein[723]) );
  DFF \ereg_reg[724]  ( .D(ereg_next[724]), .CLK(clk), .RST(rst), .I(e[724]), 
        .Q(ein[724]) );
  DFF \ereg_reg[725]  ( .D(ereg_next[725]), .CLK(clk), .RST(rst), .I(e[725]), 
        .Q(ein[725]) );
  DFF \ereg_reg[726]  ( .D(ereg_next[726]), .CLK(clk), .RST(rst), .I(e[726]), 
        .Q(ein[726]) );
  DFF \ereg_reg[727]  ( .D(ereg_next[727]), .CLK(clk), .RST(rst), .I(e[727]), 
        .Q(ein[727]) );
  DFF \ereg_reg[728]  ( .D(ereg_next[728]), .CLK(clk), .RST(rst), .I(e[728]), 
        .Q(ein[728]) );
  DFF \ereg_reg[729]  ( .D(ereg_next[729]), .CLK(clk), .RST(rst), .I(e[729]), 
        .Q(ein[729]) );
  DFF \ereg_reg[730]  ( .D(ereg_next[730]), .CLK(clk), .RST(rst), .I(e[730]), 
        .Q(ein[730]) );
  DFF \ereg_reg[731]  ( .D(ereg_next[731]), .CLK(clk), .RST(rst), .I(e[731]), 
        .Q(ein[731]) );
  DFF \ereg_reg[732]  ( .D(ereg_next[732]), .CLK(clk), .RST(rst), .I(e[732]), 
        .Q(ein[732]) );
  DFF \ereg_reg[733]  ( .D(ereg_next[733]), .CLK(clk), .RST(rst), .I(e[733]), 
        .Q(ein[733]) );
  DFF \ereg_reg[734]  ( .D(ereg_next[734]), .CLK(clk), .RST(rst), .I(e[734]), 
        .Q(ein[734]) );
  DFF \ereg_reg[735]  ( .D(ereg_next[735]), .CLK(clk), .RST(rst), .I(e[735]), 
        .Q(ein[735]) );
  DFF \ereg_reg[736]  ( .D(ereg_next[736]), .CLK(clk), .RST(rst), .I(e[736]), 
        .Q(ein[736]) );
  DFF \ereg_reg[737]  ( .D(ereg_next[737]), .CLK(clk), .RST(rst), .I(e[737]), 
        .Q(ein[737]) );
  DFF \ereg_reg[738]  ( .D(ereg_next[738]), .CLK(clk), .RST(rst), .I(e[738]), 
        .Q(ein[738]) );
  DFF \ereg_reg[739]  ( .D(ereg_next[739]), .CLK(clk), .RST(rst), .I(e[739]), 
        .Q(ein[739]) );
  DFF \ereg_reg[740]  ( .D(ereg_next[740]), .CLK(clk), .RST(rst), .I(e[740]), 
        .Q(ein[740]) );
  DFF \ereg_reg[741]  ( .D(ereg_next[741]), .CLK(clk), .RST(rst), .I(e[741]), 
        .Q(ein[741]) );
  DFF \ereg_reg[742]  ( .D(ereg_next[742]), .CLK(clk), .RST(rst), .I(e[742]), 
        .Q(ein[742]) );
  DFF \ereg_reg[743]  ( .D(ereg_next[743]), .CLK(clk), .RST(rst), .I(e[743]), 
        .Q(ein[743]) );
  DFF \ereg_reg[744]  ( .D(ereg_next[744]), .CLK(clk), .RST(rst), .I(e[744]), 
        .Q(ein[744]) );
  DFF \ereg_reg[745]  ( .D(ereg_next[745]), .CLK(clk), .RST(rst), .I(e[745]), 
        .Q(ein[745]) );
  DFF \ereg_reg[746]  ( .D(ereg_next[746]), .CLK(clk), .RST(rst), .I(e[746]), 
        .Q(ein[746]) );
  DFF \ereg_reg[747]  ( .D(ereg_next[747]), .CLK(clk), .RST(rst), .I(e[747]), 
        .Q(ein[747]) );
  DFF \ereg_reg[748]  ( .D(ereg_next[748]), .CLK(clk), .RST(rst), .I(e[748]), 
        .Q(ein[748]) );
  DFF \ereg_reg[749]  ( .D(ereg_next[749]), .CLK(clk), .RST(rst), .I(e[749]), 
        .Q(ein[749]) );
  DFF \ereg_reg[750]  ( .D(ereg_next[750]), .CLK(clk), .RST(rst), .I(e[750]), 
        .Q(ein[750]) );
  DFF \ereg_reg[751]  ( .D(ereg_next[751]), .CLK(clk), .RST(rst), .I(e[751]), 
        .Q(ein[751]) );
  DFF \ereg_reg[752]  ( .D(ereg_next[752]), .CLK(clk), .RST(rst), .I(e[752]), 
        .Q(ein[752]) );
  DFF \ereg_reg[753]  ( .D(ereg_next[753]), .CLK(clk), .RST(rst), .I(e[753]), 
        .Q(ein[753]) );
  DFF \ereg_reg[754]  ( .D(ereg_next[754]), .CLK(clk), .RST(rst), .I(e[754]), 
        .Q(ein[754]) );
  DFF \ereg_reg[755]  ( .D(ereg_next[755]), .CLK(clk), .RST(rst), .I(e[755]), 
        .Q(ein[755]) );
  DFF \ereg_reg[756]  ( .D(ereg_next[756]), .CLK(clk), .RST(rst), .I(e[756]), 
        .Q(ein[756]) );
  DFF \ereg_reg[757]  ( .D(ereg_next[757]), .CLK(clk), .RST(rst), .I(e[757]), 
        .Q(ein[757]) );
  DFF \ereg_reg[758]  ( .D(ereg_next[758]), .CLK(clk), .RST(rst), .I(e[758]), 
        .Q(ein[758]) );
  DFF \ereg_reg[759]  ( .D(ereg_next[759]), .CLK(clk), .RST(rst), .I(e[759]), 
        .Q(ein[759]) );
  DFF \ereg_reg[760]  ( .D(ereg_next[760]), .CLK(clk), .RST(rst), .I(e[760]), 
        .Q(ein[760]) );
  DFF \ereg_reg[761]  ( .D(ereg_next[761]), .CLK(clk), .RST(rst), .I(e[761]), 
        .Q(ein[761]) );
  DFF \ereg_reg[762]  ( .D(ereg_next[762]), .CLK(clk), .RST(rst), .I(e[762]), 
        .Q(ein[762]) );
  DFF \ereg_reg[763]  ( .D(ereg_next[763]), .CLK(clk), .RST(rst), .I(e[763]), 
        .Q(ein[763]) );
  DFF \ereg_reg[764]  ( .D(ereg_next[764]), .CLK(clk), .RST(rst), .I(e[764]), 
        .Q(ein[764]) );
  DFF \ereg_reg[765]  ( .D(ereg_next[765]), .CLK(clk), .RST(rst), .I(e[765]), 
        .Q(ein[765]) );
  DFF \ereg_reg[766]  ( .D(ereg_next[766]), .CLK(clk), .RST(rst), .I(e[766]), 
        .Q(ein[766]) );
  DFF \ereg_reg[767]  ( .D(ereg_next[767]), .CLK(clk), .RST(rst), .I(e[767]), 
        .Q(ein[767]) );
  DFF \ereg_reg[768]  ( .D(ereg_next[768]), .CLK(clk), .RST(rst), .I(e[768]), 
        .Q(ein[768]) );
  DFF \ereg_reg[769]  ( .D(ereg_next[769]), .CLK(clk), .RST(rst), .I(e[769]), 
        .Q(ein[769]) );
  DFF \ereg_reg[770]  ( .D(ereg_next[770]), .CLK(clk), .RST(rst), .I(e[770]), 
        .Q(ein[770]) );
  DFF \ereg_reg[771]  ( .D(ereg_next[771]), .CLK(clk), .RST(rst), .I(e[771]), 
        .Q(ein[771]) );
  DFF \ereg_reg[772]  ( .D(ereg_next[772]), .CLK(clk), .RST(rst), .I(e[772]), 
        .Q(ein[772]) );
  DFF \ereg_reg[773]  ( .D(ereg_next[773]), .CLK(clk), .RST(rst), .I(e[773]), 
        .Q(ein[773]) );
  DFF \ereg_reg[774]  ( .D(ereg_next[774]), .CLK(clk), .RST(rst), .I(e[774]), 
        .Q(ein[774]) );
  DFF \ereg_reg[775]  ( .D(ereg_next[775]), .CLK(clk), .RST(rst), .I(e[775]), 
        .Q(ein[775]) );
  DFF \ereg_reg[776]  ( .D(ereg_next[776]), .CLK(clk), .RST(rst), .I(e[776]), 
        .Q(ein[776]) );
  DFF \ereg_reg[777]  ( .D(ereg_next[777]), .CLK(clk), .RST(rst), .I(e[777]), 
        .Q(ein[777]) );
  DFF \ereg_reg[778]  ( .D(ereg_next[778]), .CLK(clk), .RST(rst), .I(e[778]), 
        .Q(ein[778]) );
  DFF \ereg_reg[779]  ( .D(ereg_next[779]), .CLK(clk), .RST(rst), .I(e[779]), 
        .Q(ein[779]) );
  DFF \ereg_reg[780]  ( .D(ereg_next[780]), .CLK(clk), .RST(rst), .I(e[780]), 
        .Q(ein[780]) );
  DFF \ereg_reg[781]  ( .D(ereg_next[781]), .CLK(clk), .RST(rst), .I(e[781]), 
        .Q(ein[781]) );
  DFF \ereg_reg[782]  ( .D(ereg_next[782]), .CLK(clk), .RST(rst), .I(e[782]), 
        .Q(ein[782]) );
  DFF \ereg_reg[783]  ( .D(ereg_next[783]), .CLK(clk), .RST(rst), .I(e[783]), 
        .Q(ein[783]) );
  DFF \ereg_reg[784]  ( .D(ereg_next[784]), .CLK(clk), .RST(rst), .I(e[784]), 
        .Q(ein[784]) );
  DFF \ereg_reg[785]  ( .D(ereg_next[785]), .CLK(clk), .RST(rst), .I(e[785]), 
        .Q(ein[785]) );
  DFF \ereg_reg[786]  ( .D(ereg_next[786]), .CLK(clk), .RST(rst), .I(e[786]), 
        .Q(ein[786]) );
  DFF \ereg_reg[787]  ( .D(ereg_next[787]), .CLK(clk), .RST(rst), .I(e[787]), 
        .Q(ein[787]) );
  DFF \ereg_reg[788]  ( .D(ereg_next[788]), .CLK(clk), .RST(rst), .I(e[788]), 
        .Q(ein[788]) );
  DFF \ereg_reg[789]  ( .D(ereg_next[789]), .CLK(clk), .RST(rst), .I(e[789]), 
        .Q(ein[789]) );
  DFF \ereg_reg[790]  ( .D(ereg_next[790]), .CLK(clk), .RST(rst), .I(e[790]), 
        .Q(ein[790]) );
  DFF \ereg_reg[791]  ( .D(ereg_next[791]), .CLK(clk), .RST(rst), .I(e[791]), 
        .Q(ein[791]) );
  DFF \ereg_reg[792]  ( .D(ereg_next[792]), .CLK(clk), .RST(rst), .I(e[792]), 
        .Q(ein[792]) );
  DFF \ereg_reg[793]  ( .D(ereg_next[793]), .CLK(clk), .RST(rst), .I(e[793]), 
        .Q(ein[793]) );
  DFF \ereg_reg[794]  ( .D(ereg_next[794]), .CLK(clk), .RST(rst), .I(e[794]), 
        .Q(ein[794]) );
  DFF \ereg_reg[795]  ( .D(ereg_next[795]), .CLK(clk), .RST(rst), .I(e[795]), 
        .Q(ein[795]) );
  DFF \ereg_reg[796]  ( .D(ereg_next[796]), .CLK(clk), .RST(rst), .I(e[796]), 
        .Q(ein[796]) );
  DFF \ereg_reg[797]  ( .D(ereg_next[797]), .CLK(clk), .RST(rst), .I(e[797]), 
        .Q(ein[797]) );
  DFF \ereg_reg[798]  ( .D(ereg_next[798]), .CLK(clk), .RST(rst), .I(e[798]), 
        .Q(ein[798]) );
  DFF \ereg_reg[799]  ( .D(ereg_next[799]), .CLK(clk), .RST(rst), .I(e[799]), 
        .Q(ein[799]) );
  DFF \ereg_reg[800]  ( .D(ereg_next[800]), .CLK(clk), .RST(rst), .I(e[800]), 
        .Q(ein[800]) );
  DFF \ereg_reg[801]  ( .D(ereg_next[801]), .CLK(clk), .RST(rst), .I(e[801]), 
        .Q(ein[801]) );
  DFF \ereg_reg[802]  ( .D(ereg_next[802]), .CLK(clk), .RST(rst), .I(e[802]), 
        .Q(ein[802]) );
  DFF \ereg_reg[803]  ( .D(ereg_next[803]), .CLK(clk), .RST(rst), .I(e[803]), 
        .Q(ein[803]) );
  DFF \ereg_reg[804]  ( .D(ereg_next[804]), .CLK(clk), .RST(rst), .I(e[804]), 
        .Q(ein[804]) );
  DFF \ereg_reg[805]  ( .D(ereg_next[805]), .CLK(clk), .RST(rst), .I(e[805]), 
        .Q(ein[805]) );
  DFF \ereg_reg[806]  ( .D(ereg_next[806]), .CLK(clk), .RST(rst), .I(e[806]), 
        .Q(ein[806]) );
  DFF \ereg_reg[807]  ( .D(ereg_next[807]), .CLK(clk), .RST(rst), .I(e[807]), 
        .Q(ein[807]) );
  DFF \ereg_reg[808]  ( .D(ereg_next[808]), .CLK(clk), .RST(rst), .I(e[808]), 
        .Q(ein[808]) );
  DFF \ereg_reg[809]  ( .D(ereg_next[809]), .CLK(clk), .RST(rst), .I(e[809]), 
        .Q(ein[809]) );
  DFF \ereg_reg[810]  ( .D(ereg_next[810]), .CLK(clk), .RST(rst), .I(e[810]), 
        .Q(ein[810]) );
  DFF \ereg_reg[811]  ( .D(ereg_next[811]), .CLK(clk), .RST(rst), .I(e[811]), 
        .Q(ein[811]) );
  DFF \ereg_reg[812]  ( .D(ereg_next[812]), .CLK(clk), .RST(rst), .I(e[812]), 
        .Q(ein[812]) );
  DFF \ereg_reg[813]  ( .D(ereg_next[813]), .CLK(clk), .RST(rst), .I(e[813]), 
        .Q(ein[813]) );
  DFF \ereg_reg[814]  ( .D(ereg_next[814]), .CLK(clk), .RST(rst), .I(e[814]), 
        .Q(ein[814]) );
  DFF \ereg_reg[815]  ( .D(ereg_next[815]), .CLK(clk), .RST(rst), .I(e[815]), 
        .Q(ein[815]) );
  DFF \ereg_reg[816]  ( .D(ereg_next[816]), .CLK(clk), .RST(rst), .I(e[816]), 
        .Q(ein[816]) );
  DFF \ereg_reg[817]  ( .D(ereg_next[817]), .CLK(clk), .RST(rst), .I(e[817]), 
        .Q(ein[817]) );
  DFF \ereg_reg[818]  ( .D(ereg_next[818]), .CLK(clk), .RST(rst), .I(e[818]), 
        .Q(ein[818]) );
  DFF \ereg_reg[819]  ( .D(ereg_next[819]), .CLK(clk), .RST(rst), .I(e[819]), 
        .Q(ein[819]) );
  DFF \ereg_reg[820]  ( .D(ereg_next[820]), .CLK(clk), .RST(rst), .I(e[820]), 
        .Q(ein[820]) );
  DFF \ereg_reg[821]  ( .D(ereg_next[821]), .CLK(clk), .RST(rst), .I(e[821]), 
        .Q(ein[821]) );
  DFF \ereg_reg[822]  ( .D(ereg_next[822]), .CLK(clk), .RST(rst), .I(e[822]), 
        .Q(ein[822]) );
  DFF \ereg_reg[823]  ( .D(ereg_next[823]), .CLK(clk), .RST(rst), .I(e[823]), 
        .Q(ein[823]) );
  DFF \ereg_reg[824]  ( .D(ereg_next[824]), .CLK(clk), .RST(rst), .I(e[824]), 
        .Q(ein[824]) );
  DFF \ereg_reg[825]  ( .D(ereg_next[825]), .CLK(clk), .RST(rst), .I(e[825]), 
        .Q(ein[825]) );
  DFF \ereg_reg[826]  ( .D(ereg_next[826]), .CLK(clk), .RST(rst), .I(e[826]), 
        .Q(ein[826]) );
  DFF \ereg_reg[827]  ( .D(ereg_next[827]), .CLK(clk), .RST(rst), .I(e[827]), 
        .Q(ein[827]) );
  DFF \ereg_reg[828]  ( .D(ereg_next[828]), .CLK(clk), .RST(rst), .I(e[828]), 
        .Q(ein[828]) );
  DFF \ereg_reg[829]  ( .D(ereg_next[829]), .CLK(clk), .RST(rst), .I(e[829]), 
        .Q(ein[829]) );
  DFF \ereg_reg[830]  ( .D(ereg_next[830]), .CLK(clk), .RST(rst), .I(e[830]), 
        .Q(ein[830]) );
  DFF \ereg_reg[831]  ( .D(ereg_next[831]), .CLK(clk), .RST(rst), .I(e[831]), 
        .Q(ein[831]) );
  DFF \ereg_reg[832]  ( .D(ereg_next[832]), .CLK(clk), .RST(rst), .I(e[832]), 
        .Q(ein[832]) );
  DFF \ereg_reg[833]  ( .D(ereg_next[833]), .CLK(clk), .RST(rst), .I(e[833]), 
        .Q(ein[833]) );
  DFF \ereg_reg[834]  ( .D(ereg_next[834]), .CLK(clk), .RST(rst), .I(e[834]), 
        .Q(ein[834]) );
  DFF \ereg_reg[835]  ( .D(ereg_next[835]), .CLK(clk), .RST(rst), .I(e[835]), 
        .Q(ein[835]) );
  DFF \ereg_reg[836]  ( .D(ereg_next[836]), .CLK(clk), .RST(rst), .I(e[836]), 
        .Q(ein[836]) );
  DFF \ereg_reg[837]  ( .D(ereg_next[837]), .CLK(clk), .RST(rst), .I(e[837]), 
        .Q(ein[837]) );
  DFF \ereg_reg[838]  ( .D(ereg_next[838]), .CLK(clk), .RST(rst), .I(e[838]), 
        .Q(ein[838]) );
  DFF \ereg_reg[839]  ( .D(ereg_next[839]), .CLK(clk), .RST(rst), .I(e[839]), 
        .Q(ein[839]) );
  DFF \ereg_reg[840]  ( .D(ereg_next[840]), .CLK(clk), .RST(rst), .I(e[840]), 
        .Q(ein[840]) );
  DFF \ereg_reg[841]  ( .D(ereg_next[841]), .CLK(clk), .RST(rst), .I(e[841]), 
        .Q(ein[841]) );
  DFF \ereg_reg[842]  ( .D(ereg_next[842]), .CLK(clk), .RST(rst), .I(e[842]), 
        .Q(ein[842]) );
  DFF \ereg_reg[843]  ( .D(ereg_next[843]), .CLK(clk), .RST(rst), .I(e[843]), 
        .Q(ein[843]) );
  DFF \ereg_reg[844]  ( .D(ereg_next[844]), .CLK(clk), .RST(rst), .I(e[844]), 
        .Q(ein[844]) );
  DFF \ereg_reg[845]  ( .D(ereg_next[845]), .CLK(clk), .RST(rst), .I(e[845]), 
        .Q(ein[845]) );
  DFF \ereg_reg[846]  ( .D(ereg_next[846]), .CLK(clk), .RST(rst), .I(e[846]), 
        .Q(ein[846]) );
  DFF \ereg_reg[847]  ( .D(ereg_next[847]), .CLK(clk), .RST(rst), .I(e[847]), 
        .Q(ein[847]) );
  DFF \ereg_reg[848]  ( .D(ereg_next[848]), .CLK(clk), .RST(rst), .I(e[848]), 
        .Q(ein[848]) );
  DFF \ereg_reg[849]  ( .D(ereg_next[849]), .CLK(clk), .RST(rst), .I(e[849]), 
        .Q(ein[849]) );
  DFF \ereg_reg[850]  ( .D(ereg_next[850]), .CLK(clk), .RST(rst), .I(e[850]), 
        .Q(ein[850]) );
  DFF \ereg_reg[851]  ( .D(ereg_next[851]), .CLK(clk), .RST(rst), .I(e[851]), 
        .Q(ein[851]) );
  DFF \ereg_reg[852]  ( .D(ereg_next[852]), .CLK(clk), .RST(rst), .I(e[852]), 
        .Q(ein[852]) );
  DFF \ereg_reg[853]  ( .D(ereg_next[853]), .CLK(clk), .RST(rst), .I(e[853]), 
        .Q(ein[853]) );
  DFF \ereg_reg[854]  ( .D(ereg_next[854]), .CLK(clk), .RST(rst), .I(e[854]), 
        .Q(ein[854]) );
  DFF \ereg_reg[855]  ( .D(ereg_next[855]), .CLK(clk), .RST(rst), .I(e[855]), 
        .Q(ein[855]) );
  DFF \ereg_reg[856]  ( .D(ereg_next[856]), .CLK(clk), .RST(rst), .I(e[856]), 
        .Q(ein[856]) );
  DFF \ereg_reg[857]  ( .D(ereg_next[857]), .CLK(clk), .RST(rst), .I(e[857]), 
        .Q(ein[857]) );
  DFF \ereg_reg[858]  ( .D(ereg_next[858]), .CLK(clk), .RST(rst), .I(e[858]), 
        .Q(ein[858]) );
  DFF \ereg_reg[859]  ( .D(ereg_next[859]), .CLK(clk), .RST(rst), .I(e[859]), 
        .Q(ein[859]) );
  DFF \ereg_reg[860]  ( .D(ereg_next[860]), .CLK(clk), .RST(rst), .I(e[860]), 
        .Q(ein[860]) );
  DFF \ereg_reg[861]  ( .D(ereg_next[861]), .CLK(clk), .RST(rst), .I(e[861]), 
        .Q(ein[861]) );
  DFF \ereg_reg[862]  ( .D(ereg_next[862]), .CLK(clk), .RST(rst), .I(e[862]), 
        .Q(ein[862]) );
  DFF \ereg_reg[863]  ( .D(ereg_next[863]), .CLK(clk), .RST(rst), .I(e[863]), 
        .Q(ein[863]) );
  DFF \ereg_reg[864]  ( .D(ereg_next[864]), .CLK(clk), .RST(rst), .I(e[864]), 
        .Q(ein[864]) );
  DFF \ereg_reg[865]  ( .D(ereg_next[865]), .CLK(clk), .RST(rst), .I(e[865]), 
        .Q(ein[865]) );
  DFF \ereg_reg[866]  ( .D(ereg_next[866]), .CLK(clk), .RST(rst), .I(e[866]), 
        .Q(ein[866]) );
  DFF \ereg_reg[867]  ( .D(ereg_next[867]), .CLK(clk), .RST(rst), .I(e[867]), 
        .Q(ein[867]) );
  DFF \ereg_reg[868]  ( .D(ereg_next[868]), .CLK(clk), .RST(rst), .I(e[868]), 
        .Q(ein[868]) );
  DFF \ereg_reg[869]  ( .D(ereg_next[869]), .CLK(clk), .RST(rst), .I(e[869]), 
        .Q(ein[869]) );
  DFF \ereg_reg[870]  ( .D(ereg_next[870]), .CLK(clk), .RST(rst), .I(e[870]), 
        .Q(ein[870]) );
  DFF \ereg_reg[871]  ( .D(ereg_next[871]), .CLK(clk), .RST(rst), .I(e[871]), 
        .Q(ein[871]) );
  DFF \ereg_reg[872]  ( .D(ereg_next[872]), .CLK(clk), .RST(rst), .I(e[872]), 
        .Q(ein[872]) );
  DFF \ereg_reg[873]  ( .D(ereg_next[873]), .CLK(clk), .RST(rst), .I(e[873]), 
        .Q(ein[873]) );
  DFF \ereg_reg[874]  ( .D(ereg_next[874]), .CLK(clk), .RST(rst), .I(e[874]), 
        .Q(ein[874]) );
  DFF \ereg_reg[875]  ( .D(ereg_next[875]), .CLK(clk), .RST(rst), .I(e[875]), 
        .Q(ein[875]) );
  DFF \ereg_reg[876]  ( .D(ereg_next[876]), .CLK(clk), .RST(rst), .I(e[876]), 
        .Q(ein[876]) );
  DFF \ereg_reg[877]  ( .D(ereg_next[877]), .CLK(clk), .RST(rst), .I(e[877]), 
        .Q(ein[877]) );
  DFF \ereg_reg[878]  ( .D(ereg_next[878]), .CLK(clk), .RST(rst), .I(e[878]), 
        .Q(ein[878]) );
  DFF \ereg_reg[879]  ( .D(ereg_next[879]), .CLK(clk), .RST(rst), .I(e[879]), 
        .Q(ein[879]) );
  DFF \ereg_reg[880]  ( .D(ereg_next[880]), .CLK(clk), .RST(rst), .I(e[880]), 
        .Q(ein[880]) );
  DFF \ereg_reg[881]  ( .D(ereg_next[881]), .CLK(clk), .RST(rst), .I(e[881]), 
        .Q(ein[881]) );
  DFF \ereg_reg[882]  ( .D(ereg_next[882]), .CLK(clk), .RST(rst), .I(e[882]), 
        .Q(ein[882]) );
  DFF \ereg_reg[883]  ( .D(ereg_next[883]), .CLK(clk), .RST(rst), .I(e[883]), 
        .Q(ein[883]) );
  DFF \ereg_reg[884]  ( .D(ereg_next[884]), .CLK(clk), .RST(rst), .I(e[884]), 
        .Q(ein[884]) );
  DFF \ereg_reg[885]  ( .D(ereg_next[885]), .CLK(clk), .RST(rst), .I(e[885]), 
        .Q(ein[885]) );
  DFF \ereg_reg[886]  ( .D(ereg_next[886]), .CLK(clk), .RST(rst), .I(e[886]), 
        .Q(ein[886]) );
  DFF \ereg_reg[887]  ( .D(ereg_next[887]), .CLK(clk), .RST(rst), .I(e[887]), 
        .Q(ein[887]) );
  DFF \ereg_reg[888]  ( .D(ereg_next[888]), .CLK(clk), .RST(rst), .I(e[888]), 
        .Q(ein[888]) );
  DFF \ereg_reg[889]  ( .D(ereg_next[889]), .CLK(clk), .RST(rst), .I(e[889]), 
        .Q(ein[889]) );
  DFF \ereg_reg[890]  ( .D(ereg_next[890]), .CLK(clk), .RST(rst), .I(e[890]), 
        .Q(ein[890]) );
  DFF \ereg_reg[891]  ( .D(ereg_next[891]), .CLK(clk), .RST(rst), .I(e[891]), 
        .Q(ein[891]) );
  DFF \ereg_reg[892]  ( .D(ereg_next[892]), .CLK(clk), .RST(rst), .I(e[892]), 
        .Q(ein[892]) );
  DFF \ereg_reg[893]  ( .D(ereg_next[893]), .CLK(clk), .RST(rst), .I(e[893]), 
        .Q(ein[893]) );
  DFF \ereg_reg[894]  ( .D(ereg_next[894]), .CLK(clk), .RST(rst), .I(e[894]), 
        .Q(ein[894]) );
  DFF \ereg_reg[895]  ( .D(ereg_next[895]), .CLK(clk), .RST(rst), .I(e[895]), 
        .Q(ein[895]) );
  DFF \ereg_reg[896]  ( .D(ereg_next[896]), .CLK(clk), .RST(rst), .I(e[896]), 
        .Q(ein[896]) );
  DFF \ereg_reg[897]  ( .D(ereg_next[897]), .CLK(clk), .RST(rst), .I(e[897]), 
        .Q(ein[897]) );
  DFF \ereg_reg[898]  ( .D(ereg_next[898]), .CLK(clk), .RST(rst), .I(e[898]), 
        .Q(ein[898]) );
  DFF \ereg_reg[899]  ( .D(ereg_next[899]), .CLK(clk), .RST(rst), .I(e[899]), 
        .Q(ein[899]) );
  DFF \ereg_reg[900]  ( .D(ereg_next[900]), .CLK(clk), .RST(rst), .I(e[900]), 
        .Q(ein[900]) );
  DFF \ereg_reg[901]  ( .D(ereg_next[901]), .CLK(clk), .RST(rst), .I(e[901]), 
        .Q(ein[901]) );
  DFF \ereg_reg[902]  ( .D(ereg_next[902]), .CLK(clk), .RST(rst), .I(e[902]), 
        .Q(ein[902]) );
  DFF \ereg_reg[903]  ( .D(ereg_next[903]), .CLK(clk), .RST(rst), .I(e[903]), 
        .Q(ein[903]) );
  DFF \ereg_reg[904]  ( .D(ereg_next[904]), .CLK(clk), .RST(rst), .I(e[904]), 
        .Q(ein[904]) );
  DFF \ereg_reg[905]  ( .D(ereg_next[905]), .CLK(clk), .RST(rst), .I(e[905]), 
        .Q(ein[905]) );
  DFF \ereg_reg[906]  ( .D(ereg_next[906]), .CLK(clk), .RST(rst), .I(e[906]), 
        .Q(ein[906]) );
  DFF \ereg_reg[907]  ( .D(ereg_next[907]), .CLK(clk), .RST(rst), .I(e[907]), 
        .Q(ein[907]) );
  DFF \ereg_reg[908]  ( .D(ereg_next[908]), .CLK(clk), .RST(rst), .I(e[908]), 
        .Q(ein[908]) );
  DFF \ereg_reg[909]  ( .D(ereg_next[909]), .CLK(clk), .RST(rst), .I(e[909]), 
        .Q(ein[909]) );
  DFF \ereg_reg[910]  ( .D(ereg_next[910]), .CLK(clk), .RST(rst), .I(e[910]), 
        .Q(ein[910]) );
  DFF \ereg_reg[911]  ( .D(ereg_next[911]), .CLK(clk), .RST(rst), .I(e[911]), 
        .Q(ein[911]) );
  DFF \ereg_reg[912]  ( .D(ereg_next[912]), .CLK(clk), .RST(rst), .I(e[912]), 
        .Q(ein[912]) );
  DFF \ereg_reg[913]  ( .D(ereg_next[913]), .CLK(clk), .RST(rst), .I(e[913]), 
        .Q(ein[913]) );
  DFF \ereg_reg[914]  ( .D(ereg_next[914]), .CLK(clk), .RST(rst), .I(e[914]), 
        .Q(ein[914]) );
  DFF \ereg_reg[915]  ( .D(ereg_next[915]), .CLK(clk), .RST(rst), .I(e[915]), 
        .Q(ein[915]) );
  DFF \ereg_reg[916]  ( .D(ereg_next[916]), .CLK(clk), .RST(rst), .I(e[916]), 
        .Q(ein[916]) );
  DFF \ereg_reg[917]  ( .D(ereg_next[917]), .CLK(clk), .RST(rst), .I(e[917]), 
        .Q(ein[917]) );
  DFF \ereg_reg[918]  ( .D(ereg_next[918]), .CLK(clk), .RST(rst), .I(e[918]), 
        .Q(ein[918]) );
  DFF \ereg_reg[919]  ( .D(ereg_next[919]), .CLK(clk), .RST(rst), .I(e[919]), 
        .Q(ein[919]) );
  DFF \ereg_reg[920]  ( .D(ereg_next[920]), .CLK(clk), .RST(rst), .I(e[920]), 
        .Q(ein[920]) );
  DFF \ereg_reg[921]  ( .D(ereg_next[921]), .CLK(clk), .RST(rst), .I(e[921]), 
        .Q(ein[921]) );
  DFF \ereg_reg[922]  ( .D(ereg_next[922]), .CLK(clk), .RST(rst), .I(e[922]), 
        .Q(ein[922]) );
  DFF \ereg_reg[923]  ( .D(ereg_next[923]), .CLK(clk), .RST(rst), .I(e[923]), 
        .Q(ein[923]) );
  DFF \ereg_reg[924]  ( .D(ereg_next[924]), .CLK(clk), .RST(rst), .I(e[924]), 
        .Q(ein[924]) );
  DFF \ereg_reg[925]  ( .D(ereg_next[925]), .CLK(clk), .RST(rst), .I(e[925]), 
        .Q(ein[925]) );
  DFF \ereg_reg[926]  ( .D(ereg_next[926]), .CLK(clk), .RST(rst), .I(e[926]), 
        .Q(ein[926]) );
  DFF \ereg_reg[927]  ( .D(ereg_next[927]), .CLK(clk), .RST(rst), .I(e[927]), 
        .Q(ein[927]) );
  DFF \ereg_reg[928]  ( .D(ereg_next[928]), .CLK(clk), .RST(rst), .I(e[928]), 
        .Q(ein[928]) );
  DFF \ereg_reg[929]  ( .D(ereg_next[929]), .CLK(clk), .RST(rst), .I(e[929]), 
        .Q(ein[929]) );
  DFF \ereg_reg[930]  ( .D(ereg_next[930]), .CLK(clk), .RST(rst), .I(e[930]), 
        .Q(ein[930]) );
  DFF \ereg_reg[931]  ( .D(ereg_next[931]), .CLK(clk), .RST(rst), .I(e[931]), 
        .Q(ein[931]) );
  DFF \ereg_reg[932]  ( .D(ereg_next[932]), .CLK(clk), .RST(rst), .I(e[932]), 
        .Q(ein[932]) );
  DFF \ereg_reg[933]  ( .D(ereg_next[933]), .CLK(clk), .RST(rst), .I(e[933]), 
        .Q(ein[933]) );
  DFF \ereg_reg[934]  ( .D(ereg_next[934]), .CLK(clk), .RST(rst), .I(e[934]), 
        .Q(ein[934]) );
  DFF \ereg_reg[935]  ( .D(ereg_next[935]), .CLK(clk), .RST(rst), .I(e[935]), 
        .Q(ein[935]) );
  DFF \ereg_reg[936]  ( .D(ereg_next[936]), .CLK(clk), .RST(rst), .I(e[936]), 
        .Q(ein[936]) );
  DFF \ereg_reg[937]  ( .D(ereg_next[937]), .CLK(clk), .RST(rst), .I(e[937]), 
        .Q(ein[937]) );
  DFF \ereg_reg[938]  ( .D(ereg_next[938]), .CLK(clk), .RST(rst), .I(e[938]), 
        .Q(ein[938]) );
  DFF \ereg_reg[939]  ( .D(ereg_next[939]), .CLK(clk), .RST(rst), .I(e[939]), 
        .Q(ein[939]) );
  DFF \ereg_reg[940]  ( .D(ereg_next[940]), .CLK(clk), .RST(rst), .I(e[940]), 
        .Q(ein[940]) );
  DFF \ereg_reg[941]  ( .D(ereg_next[941]), .CLK(clk), .RST(rst), .I(e[941]), 
        .Q(ein[941]) );
  DFF \ereg_reg[942]  ( .D(ereg_next[942]), .CLK(clk), .RST(rst), .I(e[942]), 
        .Q(ein[942]) );
  DFF \ereg_reg[943]  ( .D(ereg_next[943]), .CLK(clk), .RST(rst), .I(e[943]), 
        .Q(ein[943]) );
  DFF \ereg_reg[944]  ( .D(ereg_next[944]), .CLK(clk), .RST(rst), .I(e[944]), 
        .Q(ein[944]) );
  DFF \ereg_reg[945]  ( .D(ereg_next[945]), .CLK(clk), .RST(rst), .I(e[945]), 
        .Q(ein[945]) );
  DFF \ereg_reg[946]  ( .D(ereg_next[946]), .CLK(clk), .RST(rst), .I(e[946]), 
        .Q(ein[946]) );
  DFF \ereg_reg[947]  ( .D(ereg_next[947]), .CLK(clk), .RST(rst), .I(e[947]), 
        .Q(ein[947]) );
  DFF \ereg_reg[948]  ( .D(ereg_next[948]), .CLK(clk), .RST(rst), .I(e[948]), 
        .Q(ein[948]) );
  DFF \ereg_reg[949]  ( .D(ereg_next[949]), .CLK(clk), .RST(rst), .I(e[949]), 
        .Q(ein[949]) );
  DFF \ereg_reg[950]  ( .D(ereg_next[950]), .CLK(clk), .RST(rst), .I(e[950]), 
        .Q(ein[950]) );
  DFF \ereg_reg[951]  ( .D(ereg_next[951]), .CLK(clk), .RST(rst), .I(e[951]), 
        .Q(ein[951]) );
  DFF \ereg_reg[952]  ( .D(ereg_next[952]), .CLK(clk), .RST(rst), .I(e[952]), 
        .Q(ein[952]) );
  DFF \ereg_reg[953]  ( .D(ereg_next[953]), .CLK(clk), .RST(rst), .I(e[953]), 
        .Q(ein[953]) );
  DFF \ereg_reg[954]  ( .D(ereg_next[954]), .CLK(clk), .RST(rst), .I(e[954]), 
        .Q(ein[954]) );
  DFF \ereg_reg[955]  ( .D(ereg_next[955]), .CLK(clk), .RST(rst), .I(e[955]), 
        .Q(ein[955]) );
  DFF \ereg_reg[956]  ( .D(ereg_next[956]), .CLK(clk), .RST(rst), .I(e[956]), 
        .Q(ein[956]) );
  DFF \ereg_reg[957]  ( .D(ereg_next[957]), .CLK(clk), .RST(rst), .I(e[957]), 
        .Q(ein[957]) );
  DFF \ereg_reg[958]  ( .D(ereg_next[958]), .CLK(clk), .RST(rst), .I(e[958]), 
        .Q(ein[958]) );
  DFF \ereg_reg[959]  ( .D(ereg_next[959]), .CLK(clk), .RST(rst), .I(e[959]), 
        .Q(ein[959]) );
  DFF \ereg_reg[960]  ( .D(ereg_next[960]), .CLK(clk), .RST(rst), .I(e[960]), 
        .Q(ein[960]) );
  DFF \ereg_reg[961]  ( .D(ereg_next[961]), .CLK(clk), .RST(rst), .I(e[961]), 
        .Q(ein[961]) );
  DFF \ereg_reg[962]  ( .D(ereg_next[962]), .CLK(clk), .RST(rst), .I(e[962]), 
        .Q(ein[962]) );
  DFF \ereg_reg[963]  ( .D(ereg_next[963]), .CLK(clk), .RST(rst), .I(e[963]), 
        .Q(ein[963]) );
  DFF \ereg_reg[964]  ( .D(ereg_next[964]), .CLK(clk), .RST(rst), .I(e[964]), 
        .Q(ein[964]) );
  DFF \ereg_reg[965]  ( .D(ereg_next[965]), .CLK(clk), .RST(rst), .I(e[965]), 
        .Q(ein[965]) );
  DFF \ereg_reg[966]  ( .D(ereg_next[966]), .CLK(clk), .RST(rst), .I(e[966]), 
        .Q(ein[966]) );
  DFF \ereg_reg[967]  ( .D(ereg_next[967]), .CLK(clk), .RST(rst), .I(e[967]), 
        .Q(ein[967]) );
  DFF \ereg_reg[968]  ( .D(ereg_next[968]), .CLK(clk), .RST(rst), .I(e[968]), 
        .Q(ein[968]) );
  DFF \ereg_reg[969]  ( .D(ereg_next[969]), .CLK(clk), .RST(rst), .I(e[969]), 
        .Q(ein[969]) );
  DFF \ereg_reg[970]  ( .D(ereg_next[970]), .CLK(clk), .RST(rst), .I(e[970]), 
        .Q(ein[970]) );
  DFF \ereg_reg[971]  ( .D(ereg_next[971]), .CLK(clk), .RST(rst), .I(e[971]), 
        .Q(ein[971]) );
  DFF \ereg_reg[972]  ( .D(ereg_next[972]), .CLK(clk), .RST(rst), .I(e[972]), 
        .Q(ein[972]) );
  DFF \ereg_reg[973]  ( .D(ereg_next[973]), .CLK(clk), .RST(rst), .I(e[973]), 
        .Q(ein[973]) );
  DFF \ereg_reg[974]  ( .D(ereg_next[974]), .CLK(clk), .RST(rst), .I(e[974]), 
        .Q(ein[974]) );
  DFF \ereg_reg[975]  ( .D(ereg_next[975]), .CLK(clk), .RST(rst), .I(e[975]), 
        .Q(ein[975]) );
  DFF \ereg_reg[976]  ( .D(ereg_next[976]), .CLK(clk), .RST(rst), .I(e[976]), 
        .Q(ein[976]) );
  DFF \ereg_reg[977]  ( .D(ereg_next[977]), .CLK(clk), .RST(rst), .I(e[977]), 
        .Q(ein[977]) );
  DFF \ereg_reg[978]  ( .D(ereg_next[978]), .CLK(clk), .RST(rst), .I(e[978]), 
        .Q(ein[978]) );
  DFF \ereg_reg[979]  ( .D(ereg_next[979]), .CLK(clk), .RST(rst), .I(e[979]), 
        .Q(ein[979]) );
  DFF \ereg_reg[980]  ( .D(ereg_next[980]), .CLK(clk), .RST(rst), .I(e[980]), 
        .Q(ein[980]) );
  DFF \ereg_reg[981]  ( .D(ereg_next[981]), .CLK(clk), .RST(rst), .I(e[981]), 
        .Q(ein[981]) );
  DFF \ereg_reg[982]  ( .D(ereg_next[982]), .CLK(clk), .RST(rst), .I(e[982]), 
        .Q(ein[982]) );
  DFF \ereg_reg[983]  ( .D(ereg_next[983]), .CLK(clk), .RST(rst), .I(e[983]), 
        .Q(ein[983]) );
  DFF \ereg_reg[984]  ( .D(ereg_next[984]), .CLK(clk), .RST(rst), .I(e[984]), 
        .Q(ein[984]) );
  DFF \ereg_reg[985]  ( .D(ereg_next[985]), .CLK(clk), .RST(rst), .I(e[985]), 
        .Q(ein[985]) );
  DFF \ereg_reg[986]  ( .D(ereg_next[986]), .CLK(clk), .RST(rst), .I(e[986]), 
        .Q(ein[986]) );
  DFF \ereg_reg[987]  ( .D(ereg_next[987]), .CLK(clk), .RST(rst), .I(e[987]), 
        .Q(ein[987]) );
  DFF \ereg_reg[988]  ( .D(ereg_next[988]), .CLK(clk), .RST(rst), .I(e[988]), 
        .Q(ein[988]) );
  DFF \ereg_reg[989]  ( .D(ereg_next[989]), .CLK(clk), .RST(rst), .I(e[989]), 
        .Q(ein[989]) );
  DFF \ereg_reg[990]  ( .D(ereg_next[990]), .CLK(clk), .RST(rst), .I(e[990]), 
        .Q(ein[990]) );
  DFF \ereg_reg[991]  ( .D(ereg_next[991]), .CLK(clk), .RST(rst), .I(e[991]), 
        .Q(ein[991]) );
  DFF \ereg_reg[992]  ( .D(ereg_next[992]), .CLK(clk), .RST(rst), .I(e[992]), 
        .Q(ein[992]) );
  DFF \ereg_reg[993]  ( .D(ereg_next[993]), .CLK(clk), .RST(rst), .I(e[993]), 
        .Q(ein[993]) );
  DFF \ereg_reg[994]  ( .D(ereg_next[994]), .CLK(clk), .RST(rst), .I(e[994]), 
        .Q(ein[994]) );
  DFF \ereg_reg[995]  ( .D(ereg_next[995]), .CLK(clk), .RST(rst), .I(e[995]), 
        .Q(ein[995]) );
  DFF \ereg_reg[996]  ( .D(ereg_next[996]), .CLK(clk), .RST(rst), .I(e[996]), 
        .Q(ein[996]) );
  DFF \ereg_reg[997]  ( .D(ereg_next[997]), .CLK(clk), .RST(rst), .I(e[997]), 
        .Q(ein[997]) );
  DFF \ereg_reg[998]  ( .D(ereg_next[998]), .CLK(clk), .RST(rst), .I(e[998]), 
        .Q(ein[998]) );
  DFF \ereg_reg[999]  ( .D(ereg_next[999]), .CLK(clk), .RST(rst), .I(e[999]), 
        .Q(ein[999]) );
  DFF \ereg_reg[1000]  ( .D(ereg_next[1000]), .CLK(clk), .RST(rst), .I(e[1000]), .Q(ein[1000]) );
  DFF \ereg_reg[1001]  ( .D(ereg_next[1001]), .CLK(clk), .RST(rst), .I(e[1001]), .Q(ein[1001]) );
  DFF \ereg_reg[1002]  ( .D(ereg_next[1002]), .CLK(clk), .RST(rst), .I(e[1002]), .Q(ein[1002]) );
  DFF \ereg_reg[1003]  ( .D(ereg_next[1003]), .CLK(clk), .RST(rst), .I(e[1003]), .Q(ein[1003]) );
  DFF \ereg_reg[1004]  ( .D(ereg_next[1004]), .CLK(clk), .RST(rst), .I(e[1004]), .Q(ein[1004]) );
  DFF \ereg_reg[1005]  ( .D(ereg_next[1005]), .CLK(clk), .RST(rst), .I(e[1005]), .Q(ein[1005]) );
  DFF \ereg_reg[1006]  ( .D(ereg_next[1006]), .CLK(clk), .RST(rst), .I(e[1006]), .Q(ein[1006]) );
  DFF \ereg_reg[1007]  ( .D(ereg_next[1007]), .CLK(clk), .RST(rst), .I(e[1007]), .Q(ein[1007]) );
  DFF \ereg_reg[1008]  ( .D(ereg_next[1008]), .CLK(clk), .RST(rst), .I(e[1008]), .Q(ein[1008]) );
  DFF \ereg_reg[1009]  ( .D(ereg_next[1009]), .CLK(clk), .RST(rst), .I(e[1009]), .Q(ein[1009]) );
  DFF \ereg_reg[1010]  ( .D(ereg_next[1010]), .CLK(clk), .RST(rst), .I(e[1010]), .Q(ein[1010]) );
  DFF \ereg_reg[1011]  ( .D(ereg_next[1011]), .CLK(clk), .RST(rst), .I(e[1011]), .Q(ein[1011]) );
  DFF \ereg_reg[1012]  ( .D(ereg_next[1012]), .CLK(clk), .RST(rst), .I(e[1012]), .Q(ein[1012]) );
  DFF \ereg_reg[1013]  ( .D(ereg_next[1013]), .CLK(clk), .RST(rst), .I(e[1013]), .Q(ein[1013]) );
  DFF \ereg_reg[1014]  ( .D(ereg_next[1014]), .CLK(clk), .RST(rst), .I(e[1014]), .Q(ein[1014]) );
  DFF \ereg_reg[1015]  ( .D(ereg_next[1015]), .CLK(clk), .RST(rst), .I(e[1015]), .Q(ein[1015]) );
  DFF \ereg_reg[1016]  ( .D(ereg_next[1016]), .CLK(clk), .RST(rst), .I(e[1016]), .Q(ein[1016]) );
  DFF \ereg_reg[1017]  ( .D(ereg_next[1017]), .CLK(clk), .RST(rst), .I(e[1017]), .Q(ein[1017]) );
  DFF \ereg_reg[1018]  ( .D(ereg_next[1018]), .CLK(clk), .RST(rst), .I(e[1018]), .Q(ein[1018]) );
  DFF \ereg_reg[1019]  ( .D(ereg_next[1019]), .CLK(clk), .RST(rst), .I(e[1019]), .Q(ein[1019]) );
  DFF \ereg_reg[1020]  ( .D(ereg_next[1020]), .CLK(clk), .RST(rst), .I(e[1020]), .Q(ein[1020]) );
  DFF \ereg_reg[1021]  ( .D(ereg_next[1021]), .CLK(clk), .RST(rst), .I(e[1021]), .Q(ein[1021]) );
  DFF \ereg_reg[1022]  ( .D(ereg_next[1022]), .CLK(clk), .RST(rst), .I(e[1022]), .Q(ein[1022]) );
  DFF \ereg_reg[1023]  ( .D(ereg_next[1023]), .CLK(clk), .RST(rst), .I(e[1023]), .Q(ein[1023]) );
  DFF first_one_reg ( .D(n6), .CLK(clk), .RST(rst), .I(1'b0), .Q(first_one) );
  DFF \creg_reg[0]  ( .D(creg_next[0]), .CLK(clk), .RST(rst), .I(m[0]), .Q(
        c[0]) );
  DFF \creg_reg[1]  ( .D(creg_next[1]), .CLK(clk), .RST(rst), .I(m[1]), .Q(
        c[1]) );
  DFF \creg_reg[2]  ( .D(creg_next[2]), .CLK(clk), .RST(rst), .I(m[2]), .Q(
        c[2]) );
  DFF \creg_reg[3]  ( .D(creg_next[3]), .CLK(clk), .RST(rst), .I(m[3]), .Q(
        c[3]) );
  DFF \creg_reg[4]  ( .D(creg_next[4]), .CLK(clk), .RST(rst), .I(m[4]), .Q(
        c[4]) );
  DFF \creg_reg[5]  ( .D(creg_next[5]), .CLK(clk), .RST(rst), .I(m[5]), .Q(
        c[5]) );
  DFF \creg_reg[6]  ( .D(creg_next[6]), .CLK(clk), .RST(rst), .I(m[6]), .Q(
        c[6]) );
  DFF \creg_reg[7]  ( .D(creg_next[7]), .CLK(clk), .RST(rst), .I(m[7]), .Q(
        c[7]) );
  DFF \creg_reg[8]  ( .D(creg_next[8]), .CLK(clk), .RST(rst), .I(m[8]), .Q(
        c[8]) );
  DFF \creg_reg[9]  ( .D(creg_next[9]), .CLK(clk), .RST(rst), .I(m[9]), .Q(
        c[9]) );
  DFF \creg_reg[10]  ( .D(creg_next[10]), .CLK(clk), .RST(rst), .I(m[10]), .Q(
        c[10]) );
  DFF \creg_reg[11]  ( .D(creg_next[11]), .CLK(clk), .RST(rst), .I(m[11]), .Q(
        c[11]) );
  DFF \creg_reg[12]  ( .D(creg_next[12]), .CLK(clk), .RST(rst), .I(m[12]), .Q(
        c[12]) );
  DFF \creg_reg[13]  ( .D(creg_next[13]), .CLK(clk), .RST(rst), .I(m[13]), .Q(
        c[13]) );
  DFF \creg_reg[14]  ( .D(creg_next[14]), .CLK(clk), .RST(rst), .I(m[14]), .Q(
        c[14]) );
  DFF \creg_reg[15]  ( .D(creg_next[15]), .CLK(clk), .RST(rst), .I(m[15]), .Q(
        c[15]) );
  DFF \creg_reg[16]  ( .D(creg_next[16]), .CLK(clk), .RST(rst), .I(m[16]), .Q(
        c[16]) );
  DFF \creg_reg[17]  ( .D(creg_next[17]), .CLK(clk), .RST(rst), .I(m[17]), .Q(
        c[17]) );
  DFF \creg_reg[18]  ( .D(creg_next[18]), .CLK(clk), .RST(rst), .I(m[18]), .Q(
        c[18]) );
  DFF \creg_reg[19]  ( .D(creg_next[19]), .CLK(clk), .RST(rst), .I(m[19]), .Q(
        c[19]) );
  DFF \creg_reg[20]  ( .D(creg_next[20]), .CLK(clk), .RST(rst), .I(m[20]), .Q(
        c[20]) );
  DFF \creg_reg[21]  ( .D(creg_next[21]), .CLK(clk), .RST(rst), .I(m[21]), .Q(
        c[21]) );
  DFF \creg_reg[22]  ( .D(creg_next[22]), .CLK(clk), .RST(rst), .I(m[22]), .Q(
        c[22]) );
  DFF \creg_reg[23]  ( .D(creg_next[23]), .CLK(clk), .RST(rst), .I(m[23]), .Q(
        c[23]) );
  DFF \creg_reg[24]  ( .D(creg_next[24]), .CLK(clk), .RST(rst), .I(m[24]), .Q(
        c[24]) );
  DFF \creg_reg[25]  ( .D(creg_next[25]), .CLK(clk), .RST(rst), .I(m[25]), .Q(
        c[25]) );
  DFF \creg_reg[26]  ( .D(creg_next[26]), .CLK(clk), .RST(rst), .I(m[26]), .Q(
        c[26]) );
  DFF \creg_reg[27]  ( .D(creg_next[27]), .CLK(clk), .RST(rst), .I(m[27]), .Q(
        c[27]) );
  DFF \creg_reg[28]  ( .D(creg_next[28]), .CLK(clk), .RST(rst), .I(m[28]), .Q(
        c[28]) );
  DFF \creg_reg[29]  ( .D(creg_next[29]), .CLK(clk), .RST(rst), .I(m[29]), .Q(
        c[29]) );
  DFF \creg_reg[30]  ( .D(creg_next[30]), .CLK(clk), .RST(rst), .I(m[30]), .Q(
        c[30]) );
  DFF \creg_reg[31]  ( .D(creg_next[31]), .CLK(clk), .RST(rst), .I(m[31]), .Q(
        c[31]) );
  DFF \creg_reg[32]  ( .D(creg_next[32]), .CLK(clk), .RST(rst), .I(m[32]), .Q(
        c[32]) );
  DFF \creg_reg[33]  ( .D(creg_next[33]), .CLK(clk), .RST(rst), .I(m[33]), .Q(
        c[33]) );
  DFF \creg_reg[34]  ( .D(creg_next[34]), .CLK(clk), .RST(rst), .I(m[34]), .Q(
        c[34]) );
  DFF \creg_reg[35]  ( .D(creg_next[35]), .CLK(clk), .RST(rst), .I(m[35]), .Q(
        c[35]) );
  DFF \creg_reg[36]  ( .D(creg_next[36]), .CLK(clk), .RST(rst), .I(m[36]), .Q(
        c[36]) );
  DFF \creg_reg[37]  ( .D(creg_next[37]), .CLK(clk), .RST(rst), .I(m[37]), .Q(
        c[37]) );
  DFF \creg_reg[38]  ( .D(creg_next[38]), .CLK(clk), .RST(rst), .I(m[38]), .Q(
        c[38]) );
  DFF \creg_reg[39]  ( .D(creg_next[39]), .CLK(clk), .RST(rst), .I(m[39]), .Q(
        c[39]) );
  DFF \creg_reg[40]  ( .D(creg_next[40]), .CLK(clk), .RST(rst), .I(m[40]), .Q(
        c[40]) );
  DFF \creg_reg[41]  ( .D(creg_next[41]), .CLK(clk), .RST(rst), .I(m[41]), .Q(
        c[41]) );
  DFF \creg_reg[42]  ( .D(creg_next[42]), .CLK(clk), .RST(rst), .I(m[42]), .Q(
        c[42]) );
  DFF \creg_reg[43]  ( .D(creg_next[43]), .CLK(clk), .RST(rst), .I(m[43]), .Q(
        c[43]) );
  DFF \creg_reg[44]  ( .D(creg_next[44]), .CLK(clk), .RST(rst), .I(m[44]), .Q(
        c[44]) );
  DFF \creg_reg[45]  ( .D(creg_next[45]), .CLK(clk), .RST(rst), .I(m[45]), .Q(
        c[45]) );
  DFF \creg_reg[46]  ( .D(creg_next[46]), .CLK(clk), .RST(rst), .I(m[46]), .Q(
        c[46]) );
  DFF \creg_reg[47]  ( .D(creg_next[47]), .CLK(clk), .RST(rst), .I(m[47]), .Q(
        c[47]) );
  DFF \creg_reg[48]  ( .D(creg_next[48]), .CLK(clk), .RST(rst), .I(m[48]), .Q(
        c[48]) );
  DFF \creg_reg[49]  ( .D(creg_next[49]), .CLK(clk), .RST(rst), .I(m[49]), .Q(
        c[49]) );
  DFF \creg_reg[50]  ( .D(creg_next[50]), .CLK(clk), .RST(rst), .I(m[50]), .Q(
        c[50]) );
  DFF \creg_reg[51]  ( .D(creg_next[51]), .CLK(clk), .RST(rst), .I(m[51]), .Q(
        c[51]) );
  DFF \creg_reg[52]  ( .D(creg_next[52]), .CLK(clk), .RST(rst), .I(m[52]), .Q(
        c[52]) );
  DFF \creg_reg[53]  ( .D(creg_next[53]), .CLK(clk), .RST(rst), .I(m[53]), .Q(
        c[53]) );
  DFF \creg_reg[54]  ( .D(creg_next[54]), .CLK(clk), .RST(rst), .I(m[54]), .Q(
        c[54]) );
  DFF \creg_reg[55]  ( .D(creg_next[55]), .CLK(clk), .RST(rst), .I(m[55]), .Q(
        c[55]) );
  DFF \creg_reg[56]  ( .D(creg_next[56]), .CLK(clk), .RST(rst), .I(m[56]), .Q(
        c[56]) );
  DFF \creg_reg[57]  ( .D(creg_next[57]), .CLK(clk), .RST(rst), .I(m[57]), .Q(
        c[57]) );
  DFF \creg_reg[58]  ( .D(creg_next[58]), .CLK(clk), .RST(rst), .I(m[58]), .Q(
        c[58]) );
  DFF \creg_reg[59]  ( .D(creg_next[59]), .CLK(clk), .RST(rst), .I(m[59]), .Q(
        c[59]) );
  DFF \creg_reg[60]  ( .D(creg_next[60]), .CLK(clk), .RST(rst), .I(m[60]), .Q(
        c[60]) );
  DFF \creg_reg[61]  ( .D(creg_next[61]), .CLK(clk), .RST(rst), .I(m[61]), .Q(
        c[61]) );
  DFF \creg_reg[62]  ( .D(creg_next[62]), .CLK(clk), .RST(rst), .I(m[62]), .Q(
        c[62]) );
  DFF \creg_reg[63]  ( .D(creg_next[63]), .CLK(clk), .RST(rst), .I(m[63]), .Q(
        c[63]) );
  DFF \creg_reg[64]  ( .D(creg_next[64]), .CLK(clk), .RST(rst), .I(m[64]), .Q(
        c[64]) );
  DFF \creg_reg[65]  ( .D(creg_next[65]), .CLK(clk), .RST(rst), .I(m[65]), .Q(
        c[65]) );
  DFF \creg_reg[66]  ( .D(creg_next[66]), .CLK(clk), .RST(rst), .I(m[66]), .Q(
        c[66]) );
  DFF \creg_reg[67]  ( .D(creg_next[67]), .CLK(clk), .RST(rst), .I(m[67]), .Q(
        c[67]) );
  DFF \creg_reg[68]  ( .D(creg_next[68]), .CLK(clk), .RST(rst), .I(m[68]), .Q(
        c[68]) );
  DFF \creg_reg[69]  ( .D(creg_next[69]), .CLK(clk), .RST(rst), .I(m[69]), .Q(
        c[69]) );
  DFF \creg_reg[70]  ( .D(creg_next[70]), .CLK(clk), .RST(rst), .I(m[70]), .Q(
        c[70]) );
  DFF \creg_reg[71]  ( .D(creg_next[71]), .CLK(clk), .RST(rst), .I(m[71]), .Q(
        c[71]) );
  DFF \creg_reg[72]  ( .D(creg_next[72]), .CLK(clk), .RST(rst), .I(m[72]), .Q(
        c[72]) );
  DFF \creg_reg[73]  ( .D(creg_next[73]), .CLK(clk), .RST(rst), .I(m[73]), .Q(
        c[73]) );
  DFF \creg_reg[74]  ( .D(creg_next[74]), .CLK(clk), .RST(rst), .I(m[74]), .Q(
        c[74]) );
  DFF \creg_reg[75]  ( .D(creg_next[75]), .CLK(clk), .RST(rst), .I(m[75]), .Q(
        c[75]) );
  DFF \creg_reg[76]  ( .D(creg_next[76]), .CLK(clk), .RST(rst), .I(m[76]), .Q(
        c[76]) );
  DFF \creg_reg[77]  ( .D(creg_next[77]), .CLK(clk), .RST(rst), .I(m[77]), .Q(
        c[77]) );
  DFF \creg_reg[78]  ( .D(creg_next[78]), .CLK(clk), .RST(rst), .I(m[78]), .Q(
        c[78]) );
  DFF \creg_reg[79]  ( .D(creg_next[79]), .CLK(clk), .RST(rst), .I(m[79]), .Q(
        c[79]) );
  DFF \creg_reg[80]  ( .D(creg_next[80]), .CLK(clk), .RST(rst), .I(m[80]), .Q(
        c[80]) );
  DFF \creg_reg[81]  ( .D(creg_next[81]), .CLK(clk), .RST(rst), .I(m[81]), .Q(
        c[81]) );
  DFF \creg_reg[82]  ( .D(creg_next[82]), .CLK(clk), .RST(rst), .I(m[82]), .Q(
        c[82]) );
  DFF \creg_reg[83]  ( .D(creg_next[83]), .CLK(clk), .RST(rst), .I(m[83]), .Q(
        c[83]) );
  DFF \creg_reg[84]  ( .D(creg_next[84]), .CLK(clk), .RST(rst), .I(m[84]), .Q(
        c[84]) );
  DFF \creg_reg[85]  ( .D(creg_next[85]), .CLK(clk), .RST(rst), .I(m[85]), .Q(
        c[85]) );
  DFF \creg_reg[86]  ( .D(creg_next[86]), .CLK(clk), .RST(rst), .I(m[86]), .Q(
        c[86]) );
  DFF \creg_reg[87]  ( .D(creg_next[87]), .CLK(clk), .RST(rst), .I(m[87]), .Q(
        c[87]) );
  DFF \creg_reg[88]  ( .D(creg_next[88]), .CLK(clk), .RST(rst), .I(m[88]), .Q(
        c[88]) );
  DFF \creg_reg[89]  ( .D(creg_next[89]), .CLK(clk), .RST(rst), .I(m[89]), .Q(
        c[89]) );
  DFF \creg_reg[90]  ( .D(creg_next[90]), .CLK(clk), .RST(rst), .I(m[90]), .Q(
        c[90]) );
  DFF \creg_reg[91]  ( .D(creg_next[91]), .CLK(clk), .RST(rst), .I(m[91]), .Q(
        c[91]) );
  DFF \creg_reg[92]  ( .D(creg_next[92]), .CLK(clk), .RST(rst), .I(m[92]), .Q(
        c[92]) );
  DFF \creg_reg[93]  ( .D(creg_next[93]), .CLK(clk), .RST(rst), .I(m[93]), .Q(
        c[93]) );
  DFF \creg_reg[94]  ( .D(creg_next[94]), .CLK(clk), .RST(rst), .I(m[94]), .Q(
        c[94]) );
  DFF \creg_reg[95]  ( .D(creg_next[95]), .CLK(clk), .RST(rst), .I(m[95]), .Q(
        c[95]) );
  DFF \creg_reg[96]  ( .D(creg_next[96]), .CLK(clk), .RST(rst), .I(m[96]), .Q(
        c[96]) );
  DFF \creg_reg[97]  ( .D(creg_next[97]), .CLK(clk), .RST(rst), .I(m[97]), .Q(
        c[97]) );
  DFF \creg_reg[98]  ( .D(creg_next[98]), .CLK(clk), .RST(rst), .I(m[98]), .Q(
        c[98]) );
  DFF \creg_reg[99]  ( .D(creg_next[99]), .CLK(clk), .RST(rst), .I(m[99]), .Q(
        c[99]) );
  DFF \creg_reg[100]  ( .D(creg_next[100]), .CLK(clk), .RST(rst), .I(m[100]), 
        .Q(c[100]) );
  DFF \creg_reg[101]  ( .D(creg_next[101]), .CLK(clk), .RST(rst), .I(m[101]), 
        .Q(c[101]) );
  DFF \creg_reg[102]  ( .D(creg_next[102]), .CLK(clk), .RST(rst), .I(m[102]), 
        .Q(c[102]) );
  DFF \creg_reg[103]  ( .D(creg_next[103]), .CLK(clk), .RST(rst), .I(m[103]), 
        .Q(c[103]) );
  DFF \creg_reg[104]  ( .D(creg_next[104]), .CLK(clk), .RST(rst), .I(m[104]), 
        .Q(c[104]) );
  DFF \creg_reg[105]  ( .D(creg_next[105]), .CLK(clk), .RST(rst), .I(m[105]), 
        .Q(c[105]) );
  DFF \creg_reg[106]  ( .D(creg_next[106]), .CLK(clk), .RST(rst), .I(m[106]), 
        .Q(c[106]) );
  DFF \creg_reg[107]  ( .D(creg_next[107]), .CLK(clk), .RST(rst), .I(m[107]), 
        .Q(c[107]) );
  DFF \creg_reg[108]  ( .D(creg_next[108]), .CLK(clk), .RST(rst), .I(m[108]), 
        .Q(c[108]) );
  DFF \creg_reg[109]  ( .D(creg_next[109]), .CLK(clk), .RST(rst), .I(m[109]), 
        .Q(c[109]) );
  DFF \creg_reg[110]  ( .D(creg_next[110]), .CLK(clk), .RST(rst), .I(m[110]), 
        .Q(c[110]) );
  DFF \creg_reg[111]  ( .D(creg_next[111]), .CLK(clk), .RST(rst), .I(m[111]), 
        .Q(c[111]) );
  DFF \creg_reg[112]  ( .D(creg_next[112]), .CLK(clk), .RST(rst), .I(m[112]), 
        .Q(c[112]) );
  DFF \creg_reg[113]  ( .D(creg_next[113]), .CLK(clk), .RST(rst), .I(m[113]), 
        .Q(c[113]) );
  DFF \creg_reg[114]  ( .D(creg_next[114]), .CLK(clk), .RST(rst), .I(m[114]), 
        .Q(c[114]) );
  DFF \creg_reg[115]  ( .D(creg_next[115]), .CLK(clk), .RST(rst), .I(m[115]), 
        .Q(c[115]) );
  DFF \creg_reg[116]  ( .D(creg_next[116]), .CLK(clk), .RST(rst), .I(m[116]), 
        .Q(c[116]) );
  DFF \creg_reg[117]  ( .D(creg_next[117]), .CLK(clk), .RST(rst), .I(m[117]), 
        .Q(c[117]) );
  DFF \creg_reg[118]  ( .D(creg_next[118]), .CLK(clk), .RST(rst), .I(m[118]), 
        .Q(c[118]) );
  DFF \creg_reg[119]  ( .D(creg_next[119]), .CLK(clk), .RST(rst), .I(m[119]), 
        .Q(c[119]) );
  DFF \creg_reg[120]  ( .D(creg_next[120]), .CLK(clk), .RST(rst), .I(m[120]), 
        .Q(c[120]) );
  DFF \creg_reg[121]  ( .D(creg_next[121]), .CLK(clk), .RST(rst), .I(m[121]), 
        .Q(c[121]) );
  DFF \creg_reg[122]  ( .D(creg_next[122]), .CLK(clk), .RST(rst), .I(m[122]), 
        .Q(c[122]) );
  DFF \creg_reg[123]  ( .D(creg_next[123]), .CLK(clk), .RST(rst), .I(m[123]), 
        .Q(c[123]) );
  DFF \creg_reg[124]  ( .D(creg_next[124]), .CLK(clk), .RST(rst), .I(m[124]), 
        .Q(c[124]) );
  DFF \creg_reg[125]  ( .D(creg_next[125]), .CLK(clk), .RST(rst), .I(m[125]), 
        .Q(c[125]) );
  DFF \creg_reg[126]  ( .D(creg_next[126]), .CLK(clk), .RST(rst), .I(m[126]), 
        .Q(c[126]) );
  DFF \creg_reg[127]  ( .D(creg_next[127]), .CLK(clk), .RST(rst), .I(m[127]), 
        .Q(c[127]) );
  DFF \creg_reg[128]  ( .D(creg_next[128]), .CLK(clk), .RST(rst), .I(m[128]), 
        .Q(c[128]) );
  DFF \creg_reg[129]  ( .D(creg_next[129]), .CLK(clk), .RST(rst), .I(m[129]), 
        .Q(c[129]) );
  DFF \creg_reg[130]  ( .D(creg_next[130]), .CLK(clk), .RST(rst), .I(m[130]), 
        .Q(c[130]) );
  DFF \creg_reg[131]  ( .D(creg_next[131]), .CLK(clk), .RST(rst), .I(m[131]), 
        .Q(c[131]) );
  DFF \creg_reg[132]  ( .D(creg_next[132]), .CLK(clk), .RST(rst), .I(m[132]), 
        .Q(c[132]) );
  DFF \creg_reg[133]  ( .D(creg_next[133]), .CLK(clk), .RST(rst), .I(m[133]), 
        .Q(c[133]) );
  DFF \creg_reg[134]  ( .D(creg_next[134]), .CLK(clk), .RST(rst), .I(m[134]), 
        .Q(c[134]) );
  DFF \creg_reg[135]  ( .D(creg_next[135]), .CLK(clk), .RST(rst), .I(m[135]), 
        .Q(c[135]) );
  DFF \creg_reg[136]  ( .D(creg_next[136]), .CLK(clk), .RST(rst), .I(m[136]), 
        .Q(c[136]) );
  DFF \creg_reg[137]  ( .D(creg_next[137]), .CLK(clk), .RST(rst), .I(m[137]), 
        .Q(c[137]) );
  DFF \creg_reg[138]  ( .D(creg_next[138]), .CLK(clk), .RST(rst), .I(m[138]), 
        .Q(c[138]) );
  DFF \creg_reg[139]  ( .D(creg_next[139]), .CLK(clk), .RST(rst), .I(m[139]), 
        .Q(c[139]) );
  DFF \creg_reg[140]  ( .D(creg_next[140]), .CLK(clk), .RST(rst), .I(m[140]), 
        .Q(c[140]) );
  DFF \creg_reg[141]  ( .D(creg_next[141]), .CLK(clk), .RST(rst), .I(m[141]), 
        .Q(c[141]) );
  DFF \creg_reg[142]  ( .D(creg_next[142]), .CLK(clk), .RST(rst), .I(m[142]), 
        .Q(c[142]) );
  DFF \creg_reg[143]  ( .D(creg_next[143]), .CLK(clk), .RST(rst), .I(m[143]), 
        .Q(c[143]) );
  DFF \creg_reg[144]  ( .D(creg_next[144]), .CLK(clk), .RST(rst), .I(m[144]), 
        .Q(c[144]) );
  DFF \creg_reg[145]  ( .D(creg_next[145]), .CLK(clk), .RST(rst), .I(m[145]), 
        .Q(c[145]) );
  DFF \creg_reg[146]  ( .D(creg_next[146]), .CLK(clk), .RST(rst), .I(m[146]), 
        .Q(c[146]) );
  DFF \creg_reg[147]  ( .D(creg_next[147]), .CLK(clk), .RST(rst), .I(m[147]), 
        .Q(c[147]) );
  DFF \creg_reg[148]  ( .D(creg_next[148]), .CLK(clk), .RST(rst), .I(m[148]), 
        .Q(c[148]) );
  DFF \creg_reg[149]  ( .D(creg_next[149]), .CLK(clk), .RST(rst), .I(m[149]), 
        .Q(c[149]) );
  DFF \creg_reg[150]  ( .D(creg_next[150]), .CLK(clk), .RST(rst), .I(m[150]), 
        .Q(c[150]) );
  DFF \creg_reg[151]  ( .D(creg_next[151]), .CLK(clk), .RST(rst), .I(m[151]), 
        .Q(c[151]) );
  DFF \creg_reg[152]  ( .D(creg_next[152]), .CLK(clk), .RST(rst), .I(m[152]), 
        .Q(c[152]) );
  DFF \creg_reg[153]  ( .D(creg_next[153]), .CLK(clk), .RST(rst), .I(m[153]), 
        .Q(c[153]) );
  DFF \creg_reg[154]  ( .D(creg_next[154]), .CLK(clk), .RST(rst), .I(m[154]), 
        .Q(c[154]) );
  DFF \creg_reg[155]  ( .D(creg_next[155]), .CLK(clk), .RST(rst), .I(m[155]), 
        .Q(c[155]) );
  DFF \creg_reg[156]  ( .D(creg_next[156]), .CLK(clk), .RST(rst), .I(m[156]), 
        .Q(c[156]) );
  DFF \creg_reg[157]  ( .D(creg_next[157]), .CLK(clk), .RST(rst), .I(m[157]), 
        .Q(c[157]) );
  DFF \creg_reg[158]  ( .D(creg_next[158]), .CLK(clk), .RST(rst), .I(m[158]), 
        .Q(c[158]) );
  DFF \creg_reg[159]  ( .D(creg_next[159]), .CLK(clk), .RST(rst), .I(m[159]), 
        .Q(c[159]) );
  DFF \creg_reg[160]  ( .D(creg_next[160]), .CLK(clk), .RST(rst), .I(m[160]), 
        .Q(c[160]) );
  DFF \creg_reg[161]  ( .D(creg_next[161]), .CLK(clk), .RST(rst), .I(m[161]), 
        .Q(c[161]) );
  DFF \creg_reg[162]  ( .D(creg_next[162]), .CLK(clk), .RST(rst), .I(m[162]), 
        .Q(c[162]) );
  DFF \creg_reg[163]  ( .D(creg_next[163]), .CLK(clk), .RST(rst), .I(m[163]), 
        .Q(c[163]) );
  DFF \creg_reg[164]  ( .D(creg_next[164]), .CLK(clk), .RST(rst), .I(m[164]), 
        .Q(c[164]) );
  DFF \creg_reg[165]  ( .D(creg_next[165]), .CLK(clk), .RST(rst), .I(m[165]), 
        .Q(c[165]) );
  DFF \creg_reg[166]  ( .D(creg_next[166]), .CLK(clk), .RST(rst), .I(m[166]), 
        .Q(c[166]) );
  DFF \creg_reg[167]  ( .D(creg_next[167]), .CLK(clk), .RST(rst), .I(m[167]), 
        .Q(c[167]) );
  DFF \creg_reg[168]  ( .D(creg_next[168]), .CLK(clk), .RST(rst), .I(m[168]), 
        .Q(c[168]) );
  DFF \creg_reg[169]  ( .D(creg_next[169]), .CLK(clk), .RST(rst), .I(m[169]), 
        .Q(c[169]) );
  DFF \creg_reg[170]  ( .D(creg_next[170]), .CLK(clk), .RST(rst), .I(m[170]), 
        .Q(c[170]) );
  DFF \creg_reg[171]  ( .D(creg_next[171]), .CLK(clk), .RST(rst), .I(m[171]), 
        .Q(c[171]) );
  DFF \creg_reg[172]  ( .D(creg_next[172]), .CLK(clk), .RST(rst), .I(m[172]), 
        .Q(c[172]) );
  DFF \creg_reg[173]  ( .D(creg_next[173]), .CLK(clk), .RST(rst), .I(m[173]), 
        .Q(c[173]) );
  DFF \creg_reg[174]  ( .D(creg_next[174]), .CLK(clk), .RST(rst), .I(m[174]), 
        .Q(c[174]) );
  DFF \creg_reg[175]  ( .D(creg_next[175]), .CLK(clk), .RST(rst), .I(m[175]), 
        .Q(c[175]) );
  DFF \creg_reg[176]  ( .D(creg_next[176]), .CLK(clk), .RST(rst), .I(m[176]), 
        .Q(c[176]) );
  DFF \creg_reg[177]  ( .D(creg_next[177]), .CLK(clk), .RST(rst), .I(m[177]), 
        .Q(c[177]) );
  DFF \creg_reg[178]  ( .D(creg_next[178]), .CLK(clk), .RST(rst), .I(m[178]), 
        .Q(c[178]) );
  DFF \creg_reg[179]  ( .D(creg_next[179]), .CLK(clk), .RST(rst), .I(m[179]), 
        .Q(c[179]) );
  DFF \creg_reg[180]  ( .D(creg_next[180]), .CLK(clk), .RST(rst), .I(m[180]), 
        .Q(c[180]) );
  DFF \creg_reg[181]  ( .D(creg_next[181]), .CLK(clk), .RST(rst), .I(m[181]), 
        .Q(c[181]) );
  DFF \creg_reg[182]  ( .D(creg_next[182]), .CLK(clk), .RST(rst), .I(m[182]), 
        .Q(c[182]) );
  DFF \creg_reg[183]  ( .D(creg_next[183]), .CLK(clk), .RST(rst), .I(m[183]), 
        .Q(c[183]) );
  DFF \creg_reg[184]  ( .D(creg_next[184]), .CLK(clk), .RST(rst), .I(m[184]), 
        .Q(c[184]) );
  DFF \creg_reg[185]  ( .D(creg_next[185]), .CLK(clk), .RST(rst), .I(m[185]), 
        .Q(c[185]) );
  DFF \creg_reg[186]  ( .D(creg_next[186]), .CLK(clk), .RST(rst), .I(m[186]), 
        .Q(c[186]) );
  DFF \creg_reg[187]  ( .D(creg_next[187]), .CLK(clk), .RST(rst), .I(m[187]), 
        .Q(c[187]) );
  DFF \creg_reg[188]  ( .D(creg_next[188]), .CLK(clk), .RST(rst), .I(m[188]), 
        .Q(c[188]) );
  DFF \creg_reg[189]  ( .D(creg_next[189]), .CLK(clk), .RST(rst), .I(m[189]), 
        .Q(c[189]) );
  DFF \creg_reg[190]  ( .D(creg_next[190]), .CLK(clk), .RST(rst), .I(m[190]), 
        .Q(c[190]) );
  DFF \creg_reg[191]  ( .D(creg_next[191]), .CLK(clk), .RST(rst), .I(m[191]), 
        .Q(c[191]) );
  DFF \creg_reg[192]  ( .D(creg_next[192]), .CLK(clk), .RST(rst), .I(m[192]), 
        .Q(c[192]) );
  DFF \creg_reg[193]  ( .D(creg_next[193]), .CLK(clk), .RST(rst), .I(m[193]), 
        .Q(c[193]) );
  DFF \creg_reg[194]  ( .D(creg_next[194]), .CLK(clk), .RST(rst), .I(m[194]), 
        .Q(c[194]) );
  DFF \creg_reg[195]  ( .D(creg_next[195]), .CLK(clk), .RST(rst), .I(m[195]), 
        .Q(c[195]) );
  DFF \creg_reg[196]  ( .D(creg_next[196]), .CLK(clk), .RST(rst), .I(m[196]), 
        .Q(c[196]) );
  DFF \creg_reg[197]  ( .D(creg_next[197]), .CLK(clk), .RST(rst), .I(m[197]), 
        .Q(c[197]) );
  DFF \creg_reg[198]  ( .D(creg_next[198]), .CLK(clk), .RST(rst), .I(m[198]), 
        .Q(c[198]) );
  DFF \creg_reg[199]  ( .D(creg_next[199]), .CLK(clk), .RST(rst), .I(m[199]), 
        .Q(c[199]) );
  DFF \creg_reg[200]  ( .D(creg_next[200]), .CLK(clk), .RST(rst), .I(m[200]), 
        .Q(c[200]) );
  DFF \creg_reg[201]  ( .D(creg_next[201]), .CLK(clk), .RST(rst), .I(m[201]), 
        .Q(c[201]) );
  DFF \creg_reg[202]  ( .D(creg_next[202]), .CLK(clk), .RST(rst), .I(m[202]), 
        .Q(c[202]) );
  DFF \creg_reg[203]  ( .D(creg_next[203]), .CLK(clk), .RST(rst), .I(m[203]), 
        .Q(c[203]) );
  DFF \creg_reg[204]  ( .D(creg_next[204]), .CLK(clk), .RST(rst), .I(m[204]), 
        .Q(c[204]) );
  DFF \creg_reg[205]  ( .D(creg_next[205]), .CLK(clk), .RST(rst), .I(m[205]), 
        .Q(c[205]) );
  DFF \creg_reg[206]  ( .D(creg_next[206]), .CLK(clk), .RST(rst), .I(m[206]), 
        .Q(c[206]) );
  DFF \creg_reg[207]  ( .D(creg_next[207]), .CLK(clk), .RST(rst), .I(m[207]), 
        .Q(c[207]) );
  DFF \creg_reg[208]  ( .D(creg_next[208]), .CLK(clk), .RST(rst), .I(m[208]), 
        .Q(c[208]) );
  DFF \creg_reg[209]  ( .D(creg_next[209]), .CLK(clk), .RST(rst), .I(m[209]), 
        .Q(c[209]) );
  DFF \creg_reg[210]  ( .D(creg_next[210]), .CLK(clk), .RST(rst), .I(m[210]), 
        .Q(c[210]) );
  DFF \creg_reg[211]  ( .D(creg_next[211]), .CLK(clk), .RST(rst), .I(m[211]), 
        .Q(c[211]) );
  DFF \creg_reg[212]  ( .D(creg_next[212]), .CLK(clk), .RST(rst), .I(m[212]), 
        .Q(c[212]) );
  DFF \creg_reg[213]  ( .D(creg_next[213]), .CLK(clk), .RST(rst), .I(m[213]), 
        .Q(c[213]) );
  DFF \creg_reg[214]  ( .D(creg_next[214]), .CLK(clk), .RST(rst), .I(m[214]), 
        .Q(c[214]) );
  DFF \creg_reg[215]  ( .D(creg_next[215]), .CLK(clk), .RST(rst), .I(m[215]), 
        .Q(c[215]) );
  DFF \creg_reg[216]  ( .D(creg_next[216]), .CLK(clk), .RST(rst), .I(m[216]), 
        .Q(c[216]) );
  DFF \creg_reg[217]  ( .D(creg_next[217]), .CLK(clk), .RST(rst), .I(m[217]), 
        .Q(c[217]) );
  DFF \creg_reg[218]  ( .D(creg_next[218]), .CLK(clk), .RST(rst), .I(m[218]), 
        .Q(c[218]) );
  DFF \creg_reg[219]  ( .D(creg_next[219]), .CLK(clk), .RST(rst), .I(m[219]), 
        .Q(c[219]) );
  DFF \creg_reg[220]  ( .D(creg_next[220]), .CLK(clk), .RST(rst), .I(m[220]), 
        .Q(c[220]) );
  DFF \creg_reg[221]  ( .D(creg_next[221]), .CLK(clk), .RST(rst), .I(m[221]), 
        .Q(c[221]) );
  DFF \creg_reg[222]  ( .D(creg_next[222]), .CLK(clk), .RST(rst), .I(m[222]), 
        .Q(c[222]) );
  DFF \creg_reg[223]  ( .D(creg_next[223]), .CLK(clk), .RST(rst), .I(m[223]), 
        .Q(c[223]) );
  DFF \creg_reg[224]  ( .D(creg_next[224]), .CLK(clk), .RST(rst), .I(m[224]), 
        .Q(c[224]) );
  DFF \creg_reg[225]  ( .D(creg_next[225]), .CLK(clk), .RST(rst), .I(m[225]), 
        .Q(c[225]) );
  DFF \creg_reg[226]  ( .D(creg_next[226]), .CLK(clk), .RST(rst), .I(m[226]), 
        .Q(c[226]) );
  DFF \creg_reg[227]  ( .D(creg_next[227]), .CLK(clk), .RST(rst), .I(m[227]), 
        .Q(c[227]) );
  DFF \creg_reg[228]  ( .D(creg_next[228]), .CLK(clk), .RST(rst), .I(m[228]), 
        .Q(c[228]) );
  DFF \creg_reg[229]  ( .D(creg_next[229]), .CLK(clk), .RST(rst), .I(m[229]), 
        .Q(c[229]) );
  DFF \creg_reg[230]  ( .D(creg_next[230]), .CLK(clk), .RST(rst), .I(m[230]), 
        .Q(c[230]) );
  DFF \creg_reg[231]  ( .D(creg_next[231]), .CLK(clk), .RST(rst), .I(m[231]), 
        .Q(c[231]) );
  DFF \creg_reg[232]  ( .D(creg_next[232]), .CLK(clk), .RST(rst), .I(m[232]), 
        .Q(c[232]) );
  DFF \creg_reg[233]  ( .D(creg_next[233]), .CLK(clk), .RST(rst), .I(m[233]), 
        .Q(c[233]) );
  DFF \creg_reg[234]  ( .D(creg_next[234]), .CLK(clk), .RST(rst), .I(m[234]), 
        .Q(c[234]) );
  DFF \creg_reg[235]  ( .D(creg_next[235]), .CLK(clk), .RST(rst), .I(m[235]), 
        .Q(c[235]) );
  DFF \creg_reg[236]  ( .D(creg_next[236]), .CLK(clk), .RST(rst), .I(m[236]), 
        .Q(c[236]) );
  DFF \creg_reg[237]  ( .D(creg_next[237]), .CLK(clk), .RST(rst), .I(m[237]), 
        .Q(c[237]) );
  DFF \creg_reg[238]  ( .D(creg_next[238]), .CLK(clk), .RST(rst), .I(m[238]), 
        .Q(c[238]) );
  DFF \creg_reg[239]  ( .D(creg_next[239]), .CLK(clk), .RST(rst), .I(m[239]), 
        .Q(c[239]) );
  DFF \creg_reg[240]  ( .D(creg_next[240]), .CLK(clk), .RST(rst), .I(m[240]), 
        .Q(c[240]) );
  DFF \creg_reg[241]  ( .D(creg_next[241]), .CLK(clk), .RST(rst), .I(m[241]), 
        .Q(c[241]) );
  DFF \creg_reg[242]  ( .D(creg_next[242]), .CLK(clk), .RST(rst), .I(m[242]), 
        .Q(c[242]) );
  DFF \creg_reg[243]  ( .D(creg_next[243]), .CLK(clk), .RST(rst), .I(m[243]), 
        .Q(c[243]) );
  DFF \creg_reg[244]  ( .D(creg_next[244]), .CLK(clk), .RST(rst), .I(m[244]), 
        .Q(c[244]) );
  DFF \creg_reg[245]  ( .D(creg_next[245]), .CLK(clk), .RST(rst), .I(m[245]), 
        .Q(c[245]) );
  DFF \creg_reg[246]  ( .D(creg_next[246]), .CLK(clk), .RST(rst), .I(m[246]), 
        .Q(c[246]) );
  DFF \creg_reg[247]  ( .D(creg_next[247]), .CLK(clk), .RST(rst), .I(m[247]), 
        .Q(c[247]) );
  DFF \creg_reg[248]  ( .D(creg_next[248]), .CLK(clk), .RST(rst), .I(m[248]), 
        .Q(c[248]) );
  DFF \creg_reg[249]  ( .D(creg_next[249]), .CLK(clk), .RST(rst), .I(m[249]), 
        .Q(c[249]) );
  DFF \creg_reg[250]  ( .D(creg_next[250]), .CLK(clk), .RST(rst), .I(m[250]), 
        .Q(c[250]) );
  DFF \creg_reg[251]  ( .D(creg_next[251]), .CLK(clk), .RST(rst), .I(m[251]), 
        .Q(c[251]) );
  DFF \creg_reg[252]  ( .D(creg_next[252]), .CLK(clk), .RST(rst), .I(m[252]), 
        .Q(c[252]) );
  DFF \creg_reg[253]  ( .D(creg_next[253]), .CLK(clk), .RST(rst), .I(m[253]), 
        .Q(c[253]) );
  DFF \creg_reg[254]  ( .D(creg_next[254]), .CLK(clk), .RST(rst), .I(m[254]), 
        .Q(c[254]) );
  DFF \creg_reg[255]  ( .D(creg_next[255]), .CLK(clk), .RST(rst), .I(m[255]), 
        .Q(c[255]) );
  DFF \creg_reg[256]  ( .D(creg_next[256]), .CLK(clk), .RST(rst), .I(m[256]), 
        .Q(c[256]) );
  DFF \creg_reg[257]  ( .D(creg_next[257]), .CLK(clk), .RST(rst), .I(m[257]), 
        .Q(c[257]) );
  DFF \creg_reg[258]  ( .D(creg_next[258]), .CLK(clk), .RST(rst), .I(m[258]), 
        .Q(c[258]) );
  DFF \creg_reg[259]  ( .D(creg_next[259]), .CLK(clk), .RST(rst), .I(m[259]), 
        .Q(c[259]) );
  DFF \creg_reg[260]  ( .D(creg_next[260]), .CLK(clk), .RST(rst), .I(m[260]), 
        .Q(c[260]) );
  DFF \creg_reg[261]  ( .D(creg_next[261]), .CLK(clk), .RST(rst), .I(m[261]), 
        .Q(c[261]) );
  DFF \creg_reg[262]  ( .D(creg_next[262]), .CLK(clk), .RST(rst), .I(m[262]), 
        .Q(c[262]) );
  DFF \creg_reg[263]  ( .D(creg_next[263]), .CLK(clk), .RST(rst), .I(m[263]), 
        .Q(c[263]) );
  DFF \creg_reg[264]  ( .D(creg_next[264]), .CLK(clk), .RST(rst), .I(m[264]), 
        .Q(c[264]) );
  DFF \creg_reg[265]  ( .D(creg_next[265]), .CLK(clk), .RST(rst), .I(m[265]), 
        .Q(c[265]) );
  DFF \creg_reg[266]  ( .D(creg_next[266]), .CLK(clk), .RST(rst), .I(m[266]), 
        .Q(c[266]) );
  DFF \creg_reg[267]  ( .D(creg_next[267]), .CLK(clk), .RST(rst), .I(m[267]), 
        .Q(c[267]) );
  DFF \creg_reg[268]  ( .D(creg_next[268]), .CLK(clk), .RST(rst), .I(m[268]), 
        .Q(c[268]) );
  DFF \creg_reg[269]  ( .D(creg_next[269]), .CLK(clk), .RST(rst), .I(m[269]), 
        .Q(c[269]) );
  DFF \creg_reg[270]  ( .D(creg_next[270]), .CLK(clk), .RST(rst), .I(m[270]), 
        .Q(c[270]) );
  DFF \creg_reg[271]  ( .D(creg_next[271]), .CLK(clk), .RST(rst), .I(m[271]), 
        .Q(c[271]) );
  DFF \creg_reg[272]  ( .D(creg_next[272]), .CLK(clk), .RST(rst), .I(m[272]), 
        .Q(c[272]) );
  DFF \creg_reg[273]  ( .D(creg_next[273]), .CLK(clk), .RST(rst), .I(m[273]), 
        .Q(c[273]) );
  DFF \creg_reg[274]  ( .D(creg_next[274]), .CLK(clk), .RST(rst), .I(m[274]), 
        .Q(c[274]) );
  DFF \creg_reg[275]  ( .D(creg_next[275]), .CLK(clk), .RST(rst), .I(m[275]), 
        .Q(c[275]) );
  DFF \creg_reg[276]  ( .D(creg_next[276]), .CLK(clk), .RST(rst), .I(m[276]), 
        .Q(c[276]) );
  DFF \creg_reg[277]  ( .D(creg_next[277]), .CLK(clk), .RST(rst), .I(m[277]), 
        .Q(c[277]) );
  DFF \creg_reg[278]  ( .D(creg_next[278]), .CLK(clk), .RST(rst), .I(m[278]), 
        .Q(c[278]) );
  DFF \creg_reg[279]  ( .D(creg_next[279]), .CLK(clk), .RST(rst), .I(m[279]), 
        .Q(c[279]) );
  DFF \creg_reg[280]  ( .D(creg_next[280]), .CLK(clk), .RST(rst), .I(m[280]), 
        .Q(c[280]) );
  DFF \creg_reg[281]  ( .D(creg_next[281]), .CLK(clk), .RST(rst), .I(m[281]), 
        .Q(c[281]) );
  DFF \creg_reg[282]  ( .D(creg_next[282]), .CLK(clk), .RST(rst), .I(m[282]), 
        .Q(c[282]) );
  DFF \creg_reg[283]  ( .D(creg_next[283]), .CLK(clk), .RST(rst), .I(m[283]), 
        .Q(c[283]) );
  DFF \creg_reg[284]  ( .D(creg_next[284]), .CLK(clk), .RST(rst), .I(m[284]), 
        .Q(c[284]) );
  DFF \creg_reg[285]  ( .D(creg_next[285]), .CLK(clk), .RST(rst), .I(m[285]), 
        .Q(c[285]) );
  DFF \creg_reg[286]  ( .D(creg_next[286]), .CLK(clk), .RST(rst), .I(m[286]), 
        .Q(c[286]) );
  DFF \creg_reg[287]  ( .D(creg_next[287]), .CLK(clk), .RST(rst), .I(m[287]), 
        .Q(c[287]) );
  DFF \creg_reg[288]  ( .D(creg_next[288]), .CLK(clk), .RST(rst), .I(m[288]), 
        .Q(c[288]) );
  DFF \creg_reg[289]  ( .D(creg_next[289]), .CLK(clk), .RST(rst), .I(m[289]), 
        .Q(c[289]) );
  DFF \creg_reg[290]  ( .D(creg_next[290]), .CLK(clk), .RST(rst), .I(m[290]), 
        .Q(c[290]) );
  DFF \creg_reg[291]  ( .D(creg_next[291]), .CLK(clk), .RST(rst), .I(m[291]), 
        .Q(c[291]) );
  DFF \creg_reg[292]  ( .D(creg_next[292]), .CLK(clk), .RST(rst), .I(m[292]), 
        .Q(c[292]) );
  DFF \creg_reg[293]  ( .D(creg_next[293]), .CLK(clk), .RST(rst), .I(m[293]), 
        .Q(c[293]) );
  DFF \creg_reg[294]  ( .D(creg_next[294]), .CLK(clk), .RST(rst), .I(m[294]), 
        .Q(c[294]) );
  DFF \creg_reg[295]  ( .D(creg_next[295]), .CLK(clk), .RST(rst), .I(m[295]), 
        .Q(c[295]) );
  DFF \creg_reg[296]  ( .D(creg_next[296]), .CLK(clk), .RST(rst), .I(m[296]), 
        .Q(c[296]) );
  DFF \creg_reg[297]  ( .D(creg_next[297]), .CLK(clk), .RST(rst), .I(m[297]), 
        .Q(c[297]) );
  DFF \creg_reg[298]  ( .D(creg_next[298]), .CLK(clk), .RST(rst), .I(m[298]), 
        .Q(c[298]) );
  DFF \creg_reg[299]  ( .D(creg_next[299]), .CLK(clk), .RST(rst), .I(m[299]), 
        .Q(c[299]) );
  DFF \creg_reg[300]  ( .D(creg_next[300]), .CLK(clk), .RST(rst), .I(m[300]), 
        .Q(c[300]) );
  DFF \creg_reg[301]  ( .D(creg_next[301]), .CLK(clk), .RST(rst), .I(m[301]), 
        .Q(c[301]) );
  DFF \creg_reg[302]  ( .D(creg_next[302]), .CLK(clk), .RST(rst), .I(m[302]), 
        .Q(c[302]) );
  DFF \creg_reg[303]  ( .D(creg_next[303]), .CLK(clk), .RST(rst), .I(m[303]), 
        .Q(c[303]) );
  DFF \creg_reg[304]  ( .D(creg_next[304]), .CLK(clk), .RST(rst), .I(m[304]), 
        .Q(c[304]) );
  DFF \creg_reg[305]  ( .D(creg_next[305]), .CLK(clk), .RST(rst), .I(m[305]), 
        .Q(c[305]) );
  DFF \creg_reg[306]  ( .D(creg_next[306]), .CLK(clk), .RST(rst), .I(m[306]), 
        .Q(c[306]) );
  DFF \creg_reg[307]  ( .D(creg_next[307]), .CLK(clk), .RST(rst), .I(m[307]), 
        .Q(c[307]) );
  DFF \creg_reg[308]  ( .D(creg_next[308]), .CLK(clk), .RST(rst), .I(m[308]), 
        .Q(c[308]) );
  DFF \creg_reg[309]  ( .D(creg_next[309]), .CLK(clk), .RST(rst), .I(m[309]), 
        .Q(c[309]) );
  DFF \creg_reg[310]  ( .D(creg_next[310]), .CLK(clk), .RST(rst), .I(m[310]), 
        .Q(c[310]) );
  DFF \creg_reg[311]  ( .D(creg_next[311]), .CLK(clk), .RST(rst), .I(m[311]), 
        .Q(c[311]) );
  DFF \creg_reg[312]  ( .D(creg_next[312]), .CLK(clk), .RST(rst), .I(m[312]), 
        .Q(c[312]) );
  DFF \creg_reg[313]  ( .D(creg_next[313]), .CLK(clk), .RST(rst), .I(m[313]), 
        .Q(c[313]) );
  DFF \creg_reg[314]  ( .D(creg_next[314]), .CLK(clk), .RST(rst), .I(m[314]), 
        .Q(c[314]) );
  DFF \creg_reg[315]  ( .D(creg_next[315]), .CLK(clk), .RST(rst), .I(m[315]), 
        .Q(c[315]) );
  DFF \creg_reg[316]  ( .D(creg_next[316]), .CLK(clk), .RST(rst), .I(m[316]), 
        .Q(c[316]) );
  DFF \creg_reg[317]  ( .D(creg_next[317]), .CLK(clk), .RST(rst), .I(m[317]), 
        .Q(c[317]) );
  DFF \creg_reg[318]  ( .D(creg_next[318]), .CLK(clk), .RST(rst), .I(m[318]), 
        .Q(c[318]) );
  DFF \creg_reg[319]  ( .D(creg_next[319]), .CLK(clk), .RST(rst), .I(m[319]), 
        .Q(c[319]) );
  DFF \creg_reg[320]  ( .D(creg_next[320]), .CLK(clk), .RST(rst), .I(m[320]), 
        .Q(c[320]) );
  DFF \creg_reg[321]  ( .D(creg_next[321]), .CLK(clk), .RST(rst), .I(m[321]), 
        .Q(c[321]) );
  DFF \creg_reg[322]  ( .D(creg_next[322]), .CLK(clk), .RST(rst), .I(m[322]), 
        .Q(c[322]) );
  DFF \creg_reg[323]  ( .D(creg_next[323]), .CLK(clk), .RST(rst), .I(m[323]), 
        .Q(c[323]) );
  DFF \creg_reg[324]  ( .D(creg_next[324]), .CLK(clk), .RST(rst), .I(m[324]), 
        .Q(c[324]) );
  DFF \creg_reg[325]  ( .D(creg_next[325]), .CLK(clk), .RST(rst), .I(m[325]), 
        .Q(c[325]) );
  DFF \creg_reg[326]  ( .D(creg_next[326]), .CLK(clk), .RST(rst), .I(m[326]), 
        .Q(c[326]) );
  DFF \creg_reg[327]  ( .D(creg_next[327]), .CLK(clk), .RST(rst), .I(m[327]), 
        .Q(c[327]) );
  DFF \creg_reg[328]  ( .D(creg_next[328]), .CLK(clk), .RST(rst), .I(m[328]), 
        .Q(c[328]) );
  DFF \creg_reg[329]  ( .D(creg_next[329]), .CLK(clk), .RST(rst), .I(m[329]), 
        .Q(c[329]) );
  DFF \creg_reg[330]  ( .D(creg_next[330]), .CLK(clk), .RST(rst), .I(m[330]), 
        .Q(c[330]) );
  DFF \creg_reg[331]  ( .D(creg_next[331]), .CLK(clk), .RST(rst), .I(m[331]), 
        .Q(c[331]) );
  DFF \creg_reg[332]  ( .D(creg_next[332]), .CLK(clk), .RST(rst), .I(m[332]), 
        .Q(c[332]) );
  DFF \creg_reg[333]  ( .D(creg_next[333]), .CLK(clk), .RST(rst), .I(m[333]), 
        .Q(c[333]) );
  DFF \creg_reg[334]  ( .D(creg_next[334]), .CLK(clk), .RST(rst), .I(m[334]), 
        .Q(c[334]) );
  DFF \creg_reg[335]  ( .D(creg_next[335]), .CLK(clk), .RST(rst), .I(m[335]), 
        .Q(c[335]) );
  DFF \creg_reg[336]  ( .D(creg_next[336]), .CLK(clk), .RST(rst), .I(m[336]), 
        .Q(c[336]) );
  DFF \creg_reg[337]  ( .D(creg_next[337]), .CLK(clk), .RST(rst), .I(m[337]), 
        .Q(c[337]) );
  DFF \creg_reg[338]  ( .D(creg_next[338]), .CLK(clk), .RST(rst), .I(m[338]), 
        .Q(c[338]) );
  DFF \creg_reg[339]  ( .D(creg_next[339]), .CLK(clk), .RST(rst), .I(m[339]), 
        .Q(c[339]) );
  DFF \creg_reg[340]  ( .D(creg_next[340]), .CLK(clk), .RST(rst), .I(m[340]), 
        .Q(c[340]) );
  DFF \creg_reg[341]  ( .D(creg_next[341]), .CLK(clk), .RST(rst), .I(m[341]), 
        .Q(c[341]) );
  DFF \creg_reg[342]  ( .D(creg_next[342]), .CLK(clk), .RST(rst), .I(m[342]), 
        .Q(c[342]) );
  DFF \creg_reg[343]  ( .D(creg_next[343]), .CLK(clk), .RST(rst), .I(m[343]), 
        .Q(c[343]) );
  DFF \creg_reg[344]  ( .D(creg_next[344]), .CLK(clk), .RST(rst), .I(m[344]), 
        .Q(c[344]) );
  DFF \creg_reg[345]  ( .D(creg_next[345]), .CLK(clk), .RST(rst), .I(m[345]), 
        .Q(c[345]) );
  DFF \creg_reg[346]  ( .D(creg_next[346]), .CLK(clk), .RST(rst), .I(m[346]), 
        .Q(c[346]) );
  DFF \creg_reg[347]  ( .D(creg_next[347]), .CLK(clk), .RST(rst), .I(m[347]), 
        .Q(c[347]) );
  DFF \creg_reg[348]  ( .D(creg_next[348]), .CLK(clk), .RST(rst), .I(m[348]), 
        .Q(c[348]) );
  DFF \creg_reg[349]  ( .D(creg_next[349]), .CLK(clk), .RST(rst), .I(m[349]), 
        .Q(c[349]) );
  DFF \creg_reg[350]  ( .D(creg_next[350]), .CLK(clk), .RST(rst), .I(m[350]), 
        .Q(c[350]) );
  DFF \creg_reg[351]  ( .D(creg_next[351]), .CLK(clk), .RST(rst), .I(m[351]), 
        .Q(c[351]) );
  DFF \creg_reg[352]  ( .D(creg_next[352]), .CLK(clk), .RST(rst), .I(m[352]), 
        .Q(c[352]) );
  DFF \creg_reg[353]  ( .D(creg_next[353]), .CLK(clk), .RST(rst), .I(m[353]), 
        .Q(c[353]) );
  DFF \creg_reg[354]  ( .D(creg_next[354]), .CLK(clk), .RST(rst), .I(m[354]), 
        .Q(c[354]) );
  DFF \creg_reg[355]  ( .D(creg_next[355]), .CLK(clk), .RST(rst), .I(m[355]), 
        .Q(c[355]) );
  DFF \creg_reg[356]  ( .D(creg_next[356]), .CLK(clk), .RST(rst), .I(m[356]), 
        .Q(c[356]) );
  DFF \creg_reg[357]  ( .D(creg_next[357]), .CLK(clk), .RST(rst), .I(m[357]), 
        .Q(c[357]) );
  DFF \creg_reg[358]  ( .D(creg_next[358]), .CLK(clk), .RST(rst), .I(m[358]), 
        .Q(c[358]) );
  DFF \creg_reg[359]  ( .D(creg_next[359]), .CLK(clk), .RST(rst), .I(m[359]), 
        .Q(c[359]) );
  DFF \creg_reg[360]  ( .D(creg_next[360]), .CLK(clk), .RST(rst), .I(m[360]), 
        .Q(c[360]) );
  DFF \creg_reg[361]  ( .D(creg_next[361]), .CLK(clk), .RST(rst), .I(m[361]), 
        .Q(c[361]) );
  DFF \creg_reg[362]  ( .D(creg_next[362]), .CLK(clk), .RST(rst), .I(m[362]), 
        .Q(c[362]) );
  DFF \creg_reg[363]  ( .D(creg_next[363]), .CLK(clk), .RST(rst), .I(m[363]), 
        .Q(c[363]) );
  DFF \creg_reg[364]  ( .D(creg_next[364]), .CLK(clk), .RST(rst), .I(m[364]), 
        .Q(c[364]) );
  DFF \creg_reg[365]  ( .D(creg_next[365]), .CLK(clk), .RST(rst), .I(m[365]), 
        .Q(c[365]) );
  DFF \creg_reg[366]  ( .D(creg_next[366]), .CLK(clk), .RST(rst), .I(m[366]), 
        .Q(c[366]) );
  DFF \creg_reg[367]  ( .D(creg_next[367]), .CLK(clk), .RST(rst), .I(m[367]), 
        .Q(c[367]) );
  DFF \creg_reg[368]  ( .D(creg_next[368]), .CLK(clk), .RST(rst), .I(m[368]), 
        .Q(c[368]) );
  DFF \creg_reg[369]  ( .D(creg_next[369]), .CLK(clk), .RST(rst), .I(m[369]), 
        .Q(c[369]) );
  DFF \creg_reg[370]  ( .D(creg_next[370]), .CLK(clk), .RST(rst), .I(m[370]), 
        .Q(c[370]) );
  DFF \creg_reg[371]  ( .D(creg_next[371]), .CLK(clk), .RST(rst), .I(m[371]), 
        .Q(c[371]) );
  DFF \creg_reg[372]  ( .D(creg_next[372]), .CLK(clk), .RST(rst), .I(m[372]), 
        .Q(c[372]) );
  DFF \creg_reg[373]  ( .D(creg_next[373]), .CLK(clk), .RST(rst), .I(m[373]), 
        .Q(c[373]) );
  DFF \creg_reg[374]  ( .D(creg_next[374]), .CLK(clk), .RST(rst), .I(m[374]), 
        .Q(c[374]) );
  DFF \creg_reg[375]  ( .D(creg_next[375]), .CLK(clk), .RST(rst), .I(m[375]), 
        .Q(c[375]) );
  DFF \creg_reg[376]  ( .D(creg_next[376]), .CLK(clk), .RST(rst), .I(m[376]), 
        .Q(c[376]) );
  DFF \creg_reg[377]  ( .D(creg_next[377]), .CLK(clk), .RST(rst), .I(m[377]), 
        .Q(c[377]) );
  DFF \creg_reg[378]  ( .D(creg_next[378]), .CLK(clk), .RST(rst), .I(m[378]), 
        .Q(c[378]) );
  DFF \creg_reg[379]  ( .D(creg_next[379]), .CLK(clk), .RST(rst), .I(m[379]), 
        .Q(c[379]) );
  DFF \creg_reg[380]  ( .D(creg_next[380]), .CLK(clk), .RST(rst), .I(m[380]), 
        .Q(c[380]) );
  DFF \creg_reg[381]  ( .D(creg_next[381]), .CLK(clk), .RST(rst), .I(m[381]), 
        .Q(c[381]) );
  DFF \creg_reg[382]  ( .D(creg_next[382]), .CLK(clk), .RST(rst), .I(m[382]), 
        .Q(c[382]) );
  DFF \creg_reg[383]  ( .D(creg_next[383]), .CLK(clk), .RST(rst), .I(m[383]), 
        .Q(c[383]) );
  DFF \creg_reg[384]  ( .D(creg_next[384]), .CLK(clk), .RST(rst), .I(m[384]), 
        .Q(c[384]) );
  DFF \creg_reg[385]  ( .D(creg_next[385]), .CLK(clk), .RST(rst), .I(m[385]), 
        .Q(c[385]) );
  DFF \creg_reg[386]  ( .D(creg_next[386]), .CLK(clk), .RST(rst), .I(m[386]), 
        .Q(c[386]) );
  DFF \creg_reg[387]  ( .D(creg_next[387]), .CLK(clk), .RST(rst), .I(m[387]), 
        .Q(c[387]) );
  DFF \creg_reg[388]  ( .D(creg_next[388]), .CLK(clk), .RST(rst), .I(m[388]), 
        .Q(c[388]) );
  DFF \creg_reg[389]  ( .D(creg_next[389]), .CLK(clk), .RST(rst), .I(m[389]), 
        .Q(c[389]) );
  DFF \creg_reg[390]  ( .D(creg_next[390]), .CLK(clk), .RST(rst), .I(m[390]), 
        .Q(c[390]) );
  DFF \creg_reg[391]  ( .D(creg_next[391]), .CLK(clk), .RST(rst), .I(m[391]), 
        .Q(c[391]) );
  DFF \creg_reg[392]  ( .D(creg_next[392]), .CLK(clk), .RST(rst), .I(m[392]), 
        .Q(c[392]) );
  DFF \creg_reg[393]  ( .D(creg_next[393]), .CLK(clk), .RST(rst), .I(m[393]), 
        .Q(c[393]) );
  DFF \creg_reg[394]  ( .D(creg_next[394]), .CLK(clk), .RST(rst), .I(m[394]), 
        .Q(c[394]) );
  DFF \creg_reg[395]  ( .D(creg_next[395]), .CLK(clk), .RST(rst), .I(m[395]), 
        .Q(c[395]) );
  DFF \creg_reg[396]  ( .D(creg_next[396]), .CLK(clk), .RST(rst), .I(m[396]), 
        .Q(c[396]) );
  DFF \creg_reg[397]  ( .D(creg_next[397]), .CLK(clk), .RST(rst), .I(m[397]), 
        .Q(c[397]) );
  DFF \creg_reg[398]  ( .D(creg_next[398]), .CLK(clk), .RST(rst), .I(m[398]), 
        .Q(c[398]) );
  DFF \creg_reg[399]  ( .D(creg_next[399]), .CLK(clk), .RST(rst), .I(m[399]), 
        .Q(c[399]) );
  DFF \creg_reg[400]  ( .D(creg_next[400]), .CLK(clk), .RST(rst), .I(m[400]), 
        .Q(c[400]) );
  DFF \creg_reg[401]  ( .D(creg_next[401]), .CLK(clk), .RST(rst), .I(m[401]), 
        .Q(c[401]) );
  DFF \creg_reg[402]  ( .D(creg_next[402]), .CLK(clk), .RST(rst), .I(m[402]), 
        .Q(c[402]) );
  DFF \creg_reg[403]  ( .D(creg_next[403]), .CLK(clk), .RST(rst), .I(m[403]), 
        .Q(c[403]) );
  DFF \creg_reg[404]  ( .D(creg_next[404]), .CLK(clk), .RST(rst), .I(m[404]), 
        .Q(c[404]) );
  DFF \creg_reg[405]  ( .D(creg_next[405]), .CLK(clk), .RST(rst), .I(m[405]), 
        .Q(c[405]) );
  DFF \creg_reg[406]  ( .D(creg_next[406]), .CLK(clk), .RST(rst), .I(m[406]), 
        .Q(c[406]) );
  DFF \creg_reg[407]  ( .D(creg_next[407]), .CLK(clk), .RST(rst), .I(m[407]), 
        .Q(c[407]) );
  DFF \creg_reg[408]  ( .D(creg_next[408]), .CLK(clk), .RST(rst), .I(m[408]), 
        .Q(c[408]) );
  DFF \creg_reg[409]  ( .D(creg_next[409]), .CLK(clk), .RST(rst), .I(m[409]), 
        .Q(c[409]) );
  DFF \creg_reg[410]  ( .D(creg_next[410]), .CLK(clk), .RST(rst), .I(m[410]), 
        .Q(c[410]) );
  DFF \creg_reg[411]  ( .D(creg_next[411]), .CLK(clk), .RST(rst), .I(m[411]), 
        .Q(c[411]) );
  DFF \creg_reg[412]  ( .D(creg_next[412]), .CLK(clk), .RST(rst), .I(m[412]), 
        .Q(c[412]) );
  DFF \creg_reg[413]  ( .D(creg_next[413]), .CLK(clk), .RST(rst), .I(m[413]), 
        .Q(c[413]) );
  DFF \creg_reg[414]  ( .D(creg_next[414]), .CLK(clk), .RST(rst), .I(m[414]), 
        .Q(c[414]) );
  DFF \creg_reg[415]  ( .D(creg_next[415]), .CLK(clk), .RST(rst), .I(m[415]), 
        .Q(c[415]) );
  DFF \creg_reg[416]  ( .D(creg_next[416]), .CLK(clk), .RST(rst), .I(m[416]), 
        .Q(c[416]) );
  DFF \creg_reg[417]  ( .D(creg_next[417]), .CLK(clk), .RST(rst), .I(m[417]), 
        .Q(c[417]) );
  DFF \creg_reg[418]  ( .D(creg_next[418]), .CLK(clk), .RST(rst), .I(m[418]), 
        .Q(c[418]) );
  DFF \creg_reg[419]  ( .D(creg_next[419]), .CLK(clk), .RST(rst), .I(m[419]), 
        .Q(c[419]) );
  DFF \creg_reg[420]  ( .D(creg_next[420]), .CLK(clk), .RST(rst), .I(m[420]), 
        .Q(c[420]) );
  DFF \creg_reg[421]  ( .D(creg_next[421]), .CLK(clk), .RST(rst), .I(m[421]), 
        .Q(c[421]) );
  DFF \creg_reg[422]  ( .D(creg_next[422]), .CLK(clk), .RST(rst), .I(m[422]), 
        .Q(c[422]) );
  DFF \creg_reg[423]  ( .D(creg_next[423]), .CLK(clk), .RST(rst), .I(m[423]), 
        .Q(c[423]) );
  DFF \creg_reg[424]  ( .D(creg_next[424]), .CLK(clk), .RST(rst), .I(m[424]), 
        .Q(c[424]) );
  DFF \creg_reg[425]  ( .D(creg_next[425]), .CLK(clk), .RST(rst), .I(m[425]), 
        .Q(c[425]) );
  DFF \creg_reg[426]  ( .D(creg_next[426]), .CLK(clk), .RST(rst), .I(m[426]), 
        .Q(c[426]) );
  DFF \creg_reg[427]  ( .D(creg_next[427]), .CLK(clk), .RST(rst), .I(m[427]), 
        .Q(c[427]) );
  DFF \creg_reg[428]  ( .D(creg_next[428]), .CLK(clk), .RST(rst), .I(m[428]), 
        .Q(c[428]) );
  DFF \creg_reg[429]  ( .D(creg_next[429]), .CLK(clk), .RST(rst), .I(m[429]), 
        .Q(c[429]) );
  DFF \creg_reg[430]  ( .D(creg_next[430]), .CLK(clk), .RST(rst), .I(m[430]), 
        .Q(c[430]) );
  DFF \creg_reg[431]  ( .D(creg_next[431]), .CLK(clk), .RST(rst), .I(m[431]), 
        .Q(c[431]) );
  DFF \creg_reg[432]  ( .D(creg_next[432]), .CLK(clk), .RST(rst), .I(m[432]), 
        .Q(c[432]) );
  DFF \creg_reg[433]  ( .D(creg_next[433]), .CLK(clk), .RST(rst), .I(m[433]), 
        .Q(c[433]) );
  DFF \creg_reg[434]  ( .D(creg_next[434]), .CLK(clk), .RST(rst), .I(m[434]), 
        .Q(c[434]) );
  DFF \creg_reg[435]  ( .D(creg_next[435]), .CLK(clk), .RST(rst), .I(m[435]), 
        .Q(c[435]) );
  DFF \creg_reg[436]  ( .D(creg_next[436]), .CLK(clk), .RST(rst), .I(m[436]), 
        .Q(c[436]) );
  DFF \creg_reg[437]  ( .D(creg_next[437]), .CLK(clk), .RST(rst), .I(m[437]), 
        .Q(c[437]) );
  DFF \creg_reg[438]  ( .D(creg_next[438]), .CLK(clk), .RST(rst), .I(m[438]), 
        .Q(c[438]) );
  DFF \creg_reg[439]  ( .D(creg_next[439]), .CLK(clk), .RST(rst), .I(m[439]), 
        .Q(c[439]) );
  DFF \creg_reg[440]  ( .D(creg_next[440]), .CLK(clk), .RST(rst), .I(m[440]), 
        .Q(c[440]) );
  DFF \creg_reg[441]  ( .D(creg_next[441]), .CLK(clk), .RST(rst), .I(m[441]), 
        .Q(c[441]) );
  DFF \creg_reg[442]  ( .D(creg_next[442]), .CLK(clk), .RST(rst), .I(m[442]), 
        .Q(c[442]) );
  DFF \creg_reg[443]  ( .D(creg_next[443]), .CLK(clk), .RST(rst), .I(m[443]), 
        .Q(c[443]) );
  DFF \creg_reg[444]  ( .D(creg_next[444]), .CLK(clk), .RST(rst), .I(m[444]), 
        .Q(c[444]) );
  DFF \creg_reg[445]  ( .D(creg_next[445]), .CLK(clk), .RST(rst), .I(m[445]), 
        .Q(c[445]) );
  DFF \creg_reg[446]  ( .D(creg_next[446]), .CLK(clk), .RST(rst), .I(m[446]), 
        .Q(c[446]) );
  DFF \creg_reg[447]  ( .D(creg_next[447]), .CLK(clk), .RST(rst), .I(m[447]), 
        .Q(c[447]) );
  DFF \creg_reg[448]  ( .D(creg_next[448]), .CLK(clk), .RST(rst), .I(m[448]), 
        .Q(c[448]) );
  DFF \creg_reg[449]  ( .D(creg_next[449]), .CLK(clk), .RST(rst), .I(m[449]), 
        .Q(c[449]) );
  DFF \creg_reg[450]  ( .D(creg_next[450]), .CLK(clk), .RST(rst), .I(m[450]), 
        .Q(c[450]) );
  DFF \creg_reg[451]  ( .D(creg_next[451]), .CLK(clk), .RST(rst), .I(m[451]), 
        .Q(c[451]) );
  DFF \creg_reg[452]  ( .D(creg_next[452]), .CLK(clk), .RST(rst), .I(m[452]), 
        .Q(c[452]) );
  DFF \creg_reg[453]  ( .D(creg_next[453]), .CLK(clk), .RST(rst), .I(m[453]), 
        .Q(c[453]) );
  DFF \creg_reg[454]  ( .D(creg_next[454]), .CLK(clk), .RST(rst), .I(m[454]), 
        .Q(c[454]) );
  DFF \creg_reg[455]  ( .D(creg_next[455]), .CLK(clk), .RST(rst), .I(m[455]), 
        .Q(c[455]) );
  DFF \creg_reg[456]  ( .D(creg_next[456]), .CLK(clk), .RST(rst), .I(m[456]), 
        .Q(c[456]) );
  DFF \creg_reg[457]  ( .D(creg_next[457]), .CLK(clk), .RST(rst), .I(m[457]), 
        .Q(c[457]) );
  DFF \creg_reg[458]  ( .D(creg_next[458]), .CLK(clk), .RST(rst), .I(m[458]), 
        .Q(c[458]) );
  DFF \creg_reg[459]  ( .D(creg_next[459]), .CLK(clk), .RST(rst), .I(m[459]), 
        .Q(c[459]) );
  DFF \creg_reg[460]  ( .D(creg_next[460]), .CLK(clk), .RST(rst), .I(m[460]), 
        .Q(c[460]) );
  DFF \creg_reg[461]  ( .D(creg_next[461]), .CLK(clk), .RST(rst), .I(m[461]), 
        .Q(c[461]) );
  DFF \creg_reg[462]  ( .D(creg_next[462]), .CLK(clk), .RST(rst), .I(m[462]), 
        .Q(c[462]) );
  DFF \creg_reg[463]  ( .D(creg_next[463]), .CLK(clk), .RST(rst), .I(m[463]), 
        .Q(c[463]) );
  DFF \creg_reg[464]  ( .D(creg_next[464]), .CLK(clk), .RST(rst), .I(m[464]), 
        .Q(c[464]) );
  DFF \creg_reg[465]  ( .D(creg_next[465]), .CLK(clk), .RST(rst), .I(m[465]), 
        .Q(c[465]) );
  DFF \creg_reg[466]  ( .D(creg_next[466]), .CLK(clk), .RST(rst), .I(m[466]), 
        .Q(c[466]) );
  DFF \creg_reg[467]  ( .D(creg_next[467]), .CLK(clk), .RST(rst), .I(m[467]), 
        .Q(c[467]) );
  DFF \creg_reg[468]  ( .D(creg_next[468]), .CLK(clk), .RST(rst), .I(m[468]), 
        .Q(c[468]) );
  DFF \creg_reg[469]  ( .D(creg_next[469]), .CLK(clk), .RST(rst), .I(m[469]), 
        .Q(c[469]) );
  DFF \creg_reg[470]  ( .D(creg_next[470]), .CLK(clk), .RST(rst), .I(m[470]), 
        .Q(c[470]) );
  DFF \creg_reg[471]  ( .D(creg_next[471]), .CLK(clk), .RST(rst), .I(m[471]), 
        .Q(c[471]) );
  DFF \creg_reg[472]  ( .D(creg_next[472]), .CLK(clk), .RST(rst), .I(m[472]), 
        .Q(c[472]) );
  DFF \creg_reg[473]  ( .D(creg_next[473]), .CLK(clk), .RST(rst), .I(m[473]), 
        .Q(c[473]) );
  DFF \creg_reg[474]  ( .D(creg_next[474]), .CLK(clk), .RST(rst), .I(m[474]), 
        .Q(c[474]) );
  DFF \creg_reg[475]  ( .D(creg_next[475]), .CLK(clk), .RST(rst), .I(m[475]), 
        .Q(c[475]) );
  DFF \creg_reg[476]  ( .D(creg_next[476]), .CLK(clk), .RST(rst), .I(m[476]), 
        .Q(c[476]) );
  DFF \creg_reg[477]  ( .D(creg_next[477]), .CLK(clk), .RST(rst), .I(m[477]), 
        .Q(c[477]) );
  DFF \creg_reg[478]  ( .D(creg_next[478]), .CLK(clk), .RST(rst), .I(m[478]), 
        .Q(c[478]) );
  DFF \creg_reg[479]  ( .D(creg_next[479]), .CLK(clk), .RST(rst), .I(m[479]), 
        .Q(c[479]) );
  DFF \creg_reg[480]  ( .D(creg_next[480]), .CLK(clk), .RST(rst), .I(m[480]), 
        .Q(c[480]) );
  DFF \creg_reg[481]  ( .D(creg_next[481]), .CLK(clk), .RST(rst), .I(m[481]), 
        .Q(c[481]) );
  DFF \creg_reg[482]  ( .D(creg_next[482]), .CLK(clk), .RST(rst), .I(m[482]), 
        .Q(c[482]) );
  DFF \creg_reg[483]  ( .D(creg_next[483]), .CLK(clk), .RST(rst), .I(m[483]), 
        .Q(c[483]) );
  DFF \creg_reg[484]  ( .D(creg_next[484]), .CLK(clk), .RST(rst), .I(m[484]), 
        .Q(c[484]) );
  DFF \creg_reg[485]  ( .D(creg_next[485]), .CLK(clk), .RST(rst), .I(m[485]), 
        .Q(c[485]) );
  DFF \creg_reg[486]  ( .D(creg_next[486]), .CLK(clk), .RST(rst), .I(m[486]), 
        .Q(c[486]) );
  DFF \creg_reg[487]  ( .D(creg_next[487]), .CLK(clk), .RST(rst), .I(m[487]), 
        .Q(c[487]) );
  DFF \creg_reg[488]  ( .D(creg_next[488]), .CLK(clk), .RST(rst), .I(m[488]), 
        .Q(c[488]) );
  DFF \creg_reg[489]  ( .D(creg_next[489]), .CLK(clk), .RST(rst), .I(m[489]), 
        .Q(c[489]) );
  DFF \creg_reg[490]  ( .D(creg_next[490]), .CLK(clk), .RST(rst), .I(m[490]), 
        .Q(c[490]) );
  DFF \creg_reg[491]  ( .D(creg_next[491]), .CLK(clk), .RST(rst), .I(m[491]), 
        .Q(c[491]) );
  DFF \creg_reg[492]  ( .D(creg_next[492]), .CLK(clk), .RST(rst), .I(m[492]), 
        .Q(c[492]) );
  DFF \creg_reg[493]  ( .D(creg_next[493]), .CLK(clk), .RST(rst), .I(m[493]), 
        .Q(c[493]) );
  DFF \creg_reg[494]  ( .D(creg_next[494]), .CLK(clk), .RST(rst), .I(m[494]), 
        .Q(c[494]) );
  DFF \creg_reg[495]  ( .D(creg_next[495]), .CLK(clk), .RST(rst), .I(m[495]), 
        .Q(c[495]) );
  DFF \creg_reg[496]  ( .D(creg_next[496]), .CLK(clk), .RST(rst), .I(m[496]), 
        .Q(c[496]) );
  DFF \creg_reg[497]  ( .D(creg_next[497]), .CLK(clk), .RST(rst), .I(m[497]), 
        .Q(c[497]) );
  DFF \creg_reg[498]  ( .D(creg_next[498]), .CLK(clk), .RST(rst), .I(m[498]), 
        .Q(c[498]) );
  DFF \creg_reg[499]  ( .D(creg_next[499]), .CLK(clk), .RST(rst), .I(m[499]), 
        .Q(c[499]) );
  DFF \creg_reg[500]  ( .D(creg_next[500]), .CLK(clk), .RST(rst), .I(m[500]), 
        .Q(c[500]) );
  DFF \creg_reg[501]  ( .D(creg_next[501]), .CLK(clk), .RST(rst), .I(m[501]), 
        .Q(c[501]) );
  DFF \creg_reg[502]  ( .D(creg_next[502]), .CLK(clk), .RST(rst), .I(m[502]), 
        .Q(c[502]) );
  DFF \creg_reg[503]  ( .D(creg_next[503]), .CLK(clk), .RST(rst), .I(m[503]), 
        .Q(c[503]) );
  DFF \creg_reg[504]  ( .D(creg_next[504]), .CLK(clk), .RST(rst), .I(m[504]), 
        .Q(c[504]) );
  DFF \creg_reg[505]  ( .D(creg_next[505]), .CLK(clk), .RST(rst), .I(m[505]), 
        .Q(c[505]) );
  DFF \creg_reg[506]  ( .D(creg_next[506]), .CLK(clk), .RST(rst), .I(m[506]), 
        .Q(c[506]) );
  DFF \creg_reg[507]  ( .D(creg_next[507]), .CLK(clk), .RST(rst), .I(m[507]), 
        .Q(c[507]) );
  DFF \creg_reg[508]  ( .D(creg_next[508]), .CLK(clk), .RST(rst), .I(m[508]), 
        .Q(c[508]) );
  DFF \creg_reg[509]  ( .D(creg_next[509]), .CLK(clk), .RST(rst), .I(m[509]), 
        .Q(c[509]) );
  DFF \creg_reg[510]  ( .D(creg_next[510]), .CLK(clk), .RST(rst), .I(m[510]), 
        .Q(c[510]) );
  DFF \creg_reg[511]  ( .D(creg_next[511]), .CLK(clk), .RST(rst), .I(m[511]), 
        .Q(c[511]) );
  DFF \creg_reg[512]  ( .D(creg_next[512]), .CLK(clk), .RST(rst), .I(m[512]), 
        .Q(c[512]) );
  DFF \creg_reg[513]  ( .D(creg_next[513]), .CLK(clk), .RST(rst), .I(m[513]), 
        .Q(c[513]) );
  DFF \creg_reg[514]  ( .D(creg_next[514]), .CLK(clk), .RST(rst), .I(m[514]), 
        .Q(c[514]) );
  DFF \creg_reg[515]  ( .D(creg_next[515]), .CLK(clk), .RST(rst), .I(m[515]), 
        .Q(c[515]) );
  DFF \creg_reg[516]  ( .D(creg_next[516]), .CLK(clk), .RST(rst), .I(m[516]), 
        .Q(c[516]) );
  DFF \creg_reg[517]  ( .D(creg_next[517]), .CLK(clk), .RST(rst), .I(m[517]), 
        .Q(c[517]) );
  DFF \creg_reg[518]  ( .D(creg_next[518]), .CLK(clk), .RST(rst), .I(m[518]), 
        .Q(c[518]) );
  DFF \creg_reg[519]  ( .D(creg_next[519]), .CLK(clk), .RST(rst), .I(m[519]), 
        .Q(c[519]) );
  DFF \creg_reg[520]  ( .D(creg_next[520]), .CLK(clk), .RST(rst), .I(m[520]), 
        .Q(c[520]) );
  DFF \creg_reg[521]  ( .D(creg_next[521]), .CLK(clk), .RST(rst), .I(m[521]), 
        .Q(c[521]) );
  DFF \creg_reg[522]  ( .D(creg_next[522]), .CLK(clk), .RST(rst), .I(m[522]), 
        .Q(c[522]) );
  DFF \creg_reg[523]  ( .D(creg_next[523]), .CLK(clk), .RST(rst), .I(m[523]), 
        .Q(c[523]) );
  DFF \creg_reg[524]  ( .D(creg_next[524]), .CLK(clk), .RST(rst), .I(m[524]), 
        .Q(c[524]) );
  DFF \creg_reg[525]  ( .D(creg_next[525]), .CLK(clk), .RST(rst), .I(m[525]), 
        .Q(c[525]) );
  DFF \creg_reg[526]  ( .D(creg_next[526]), .CLK(clk), .RST(rst), .I(m[526]), 
        .Q(c[526]) );
  DFF \creg_reg[527]  ( .D(creg_next[527]), .CLK(clk), .RST(rst), .I(m[527]), 
        .Q(c[527]) );
  DFF \creg_reg[528]  ( .D(creg_next[528]), .CLK(clk), .RST(rst), .I(m[528]), 
        .Q(c[528]) );
  DFF \creg_reg[529]  ( .D(creg_next[529]), .CLK(clk), .RST(rst), .I(m[529]), 
        .Q(c[529]) );
  DFF \creg_reg[530]  ( .D(creg_next[530]), .CLK(clk), .RST(rst), .I(m[530]), 
        .Q(c[530]) );
  DFF \creg_reg[531]  ( .D(creg_next[531]), .CLK(clk), .RST(rst), .I(m[531]), 
        .Q(c[531]) );
  DFF \creg_reg[532]  ( .D(creg_next[532]), .CLK(clk), .RST(rst), .I(m[532]), 
        .Q(c[532]) );
  DFF \creg_reg[533]  ( .D(creg_next[533]), .CLK(clk), .RST(rst), .I(m[533]), 
        .Q(c[533]) );
  DFF \creg_reg[534]  ( .D(creg_next[534]), .CLK(clk), .RST(rst), .I(m[534]), 
        .Q(c[534]) );
  DFF \creg_reg[535]  ( .D(creg_next[535]), .CLK(clk), .RST(rst), .I(m[535]), 
        .Q(c[535]) );
  DFF \creg_reg[536]  ( .D(creg_next[536]), .CLK(clk), .RST(rst), .I(m[536]), 
        .Q(c[536]) );
  DFF \creg_reg[537]  ( .D(creg_next[537]), .CLK(clk), .RST(rst), .I(m[537]), 
        .Q(c[537]) );
  DFF \creg_reg[538]  ( .D(creg_next[538]), .CLK(clk), .RST(rst), .I(m[538]), 
        .Q(c[538]) );
  DFF \creg_reg[539]  ( .D(creg_next[539]), .CLK(clk), .RST(rst), .I(m[539]), 
        .Q(c[539]) );
  DFF \creg_reg[540]  ( .D(creg_next[540]), .CLK(clk), .RST(rst), .I(m[540]), 
        .Q(c[540]) );
  DFF \creg_reg[541]  ( .D(creg_next[541]), .CLK(clk), .RST(rst), .I(m[541]), 
        .Q(c[541]) );
  DFF \creg_reg[542]  ( .D(creg_next[542]), .CLK(clk), .RST(rst), .I(m[542]), 
        .Q(c[542]) );
  DFF \creg_reg[543]  ( .D(creg_next[543]), .CLK(clk), .RST(rst), .I(m[543]), 
        .Q(c[543]) );
  DFF \creg_reg[544]  ( .D(creg_next[544]), .CLK(clk), .RST(rst), .I(m[544]), 
        .Q(c[544]) );
  DFF \creg_reg[545]  ( .D(creg_next[545]), .CLK(clk), .RST(rst), .I(m[545]), 
        .Q(c[545]) );
  DFF \creg_reg[546]  ( .D(creg_next[546]), .CLK(clk), .RST(rst), .I(m[546]), 
        .Q(c[546]) );
  DFF \creg_reg[547]  ( .D(creg_next[547]), .CLK(clk), .RST(rst), .I(m[547]), 
        .Q(c[547]) );
  DFF \creg_reg[548]  ( .D(creg_next[548]), .CLK(clk), .RST(rst), .I(m[548]), 
        .Q(c[548]) );
  DFF \creg_reg[549]  ( .D(creg_next[549]), .CLK(clk), .RST(rst), .I(m[549]), 
        .Q(c[549]) );
  DFF \creg_reg[550]  ( .D(creg_next[550]), .CLK(clk), .RST(rst), .I(m[550]), 
        .Q(c[550]) );
  DFF \creg_reg[551]  ( .D(creg_next[551]), .CLK(clk), .RST(rst), .I(m[551]), 
        .Q(c[551]) );
  DFF \creg_reg[552]  ( .D(creg_next[552]), .CLK(clk), .RST(rst), .I(m[552]), 
        .Q(c[552]) );
  DFF \creg_reg[553]  ( .D(creg_next[553]), .CLK(clk), .RST(rst), .I(m[553]), 
        .Q(c[553]) );
  DFF \creg_reg[554]  ( .D(creg_next[554]), .CLK(clk), .RST(rst), .I(m[554]), 
        .Q(c[554]) );
  DFF \creg_reg[555]  ( .D(creg_next[555]), .CLK(clk), .RST(rst), .I(m[555]), 
        .Q(c[555]) );
  DFF \creg_reg[556]  ( .D(creg_next[556]), .CLK(clk), .RST(rst), .I(m[556]), 
        .Q(c[556]) );
  DFF \creg_reg[557]  ( .D(creg_next[557]), .CLK(clk), .RST(rst), .I(m[557]), 
        .Q(c[557]) );
  DFF \creg_reg[558]  ( .D(creg_next[558]), .CLK(clk), .RST(rst), .I(m[558]), 
        .Q(c[558]) );
  DFF \creg_reg[559]  ( .D(creg_next[559]), .CLK(clk), .RST(rst), .I(m[559]), 
        .Q(c[559]) );
  DFF \creg_reg[560]  ( .D(creg_next[560]), .CLK(clk), .RST(rst), .I(m[560]), 
        .Q(c[560]) );
  DFF \creg_reg[561]  ( .D(creg_next[561]), .CLK(clk), .RST(rst), .I(m[561]), 
        .Q(c[561]) );
  DFF \creg_reg[562]  ( .D(creg_next[562]), .CLK(clk), .RST(rst), .I(m[562]), 
        .Q(c[562]) );
  DFF \creg_reg[563]  ( .D(creg_next[563]), .CLK(clk), .RST(rst), .I(m[563]), 
        .Q(c[563]) );
  DFF \creg_reg[564]  ( .D(creg_next[564]), .CLK(clk), .RST(rst), .I(m[564]), 
        .Q(c[564]) );
  DFF \creg_reg[565]  ( .D(creg_next[565]), .CLK(clk), .RST(rst), .I(m[565]), 
        .Q(c[565]) );
  DFF \creg_reg[566]  ( .D(creg_next[566]), .CLK(clk), .RST(rst), .I(m[566]), 
        .Q(c[566]) );
  DFF \creg_reg[567]  ( .D(creg_next[567]), .CLK(clk), .RST(rst), .I(m[567]), 
        .Q(c[567]) );
  DFF \creg_reg[568]  ( .D(creg_next[568]), .CLK(clk), .RST(rst), .I(m[568]), 
        .Q(c[568]) );
  DFF \creg_reg[569]  ( .D(creg_next[569]), .CLK(clk), .RST(rst), .I(m[569]), 
        .Q(c[569]) );
  DFF \creg_reg[570]  ( .D(creg_next[570]), .CLK(clk), .RST(rst), .I(m[570]), 
        .Q(c[570]) );
  DFF \creg_reg[571]  ( .D(creg_next[571]), .CLK(clk), .RST(rst), .I(m[571]), 
        .Q(c[571]) );
  DFF \creg_reg[572]  ( .D(creg_next[572]), .CLK(clk), .RST(rst), .I(m[572]), 
        .Q(c[572]) );
  DFF \creg_reg[573]  ( .D(creg_next[573]), .CLK(clk), .RST(rst), .I(m[573]), 
        .Q(c[573]) );
  DFF \creg_reg[574]  ( .D(creg_next[574]), .CLK(clk), .RST(rst), .I(m[574]), 
        .Q(c[574]) );
  DFF \creg_reg[575]  ( .D(creg_next[575]), .CLK(clk), .RST(rst), .I(m[575]), 
        .Q(c[575]) );
  DFF \creg_reg[576]  ( .D(creg_next[576]), .CLK(clk), .RST(rst), .I(m[576]), 
        .Q(c[576]) );
  DFF \creg_reg[577]  ( .D(creg_next[577]), .CLK(clk), .RST(rst), .I(m[577]), 
        .Q(c[577]) );
  DFF \creg_reg[578]  ( .D(creg_next[578]), .CLK(clk), .RST(rst), .I(m[578]), 
        .Q(c[578]) );
  DFF \creg_reg[579]  ( .D(creg_next[579]), .CLK(clk), .RST(rst), .I(m[579]), 
        .Q(c[579]) );
  DFF \creg_reg[580]  ( .D(creg_next[580]), .CLK(clk), .RST(rst), .I(m[580]), 
        .Q(c[580]) );
  DFF \creg_reg[581]  ( .D(creg_next[581]), .CLK(clk), .RST(rst), .I(m[581]), 
        .Q(c[581]) );
  DFF \creg_reg[582]  ( .D(creg_next[582]), .CLK(clk), .RST(rst), .I(m[582]), 
        .Q(c[582]) );
  DFF \creg_reg[583]  ( .D(creg_next[583]), .CLK(clk), .RST(rst), .I(m[583]), 
        .Q(c[583]) );
  DFF \creg_reg[584]  ( .D(creg_next[584]), .CLK(clk), .RST(rst), .I(m[584]), 
        .Q(c[584]) );
  DFF \creg_reg[585]  ( .D(creg_next[585]), .CLK(clk), .RST(rst), .I(m[585]), 
        .Q(c[585]) );
  DFF \creg_reg[586]  ( .D(creg_next[586]), .CLK(clk), .RST(rst), .I(m[586]), 
        .Q(c[586]) );
  DFF \creg_reg[587]  ( .D(creg_next[587]), .CLK(clk), .RST(rst), .I(m[587]), 
        .Q(c[587]) );
  DFF \creg_reg[588]  ( .D(creg_next[588]), .CLK(clk), .RST(rst), .I(m[588]), 
        .Q(c[588]) );
  DFF \creg_reg[589]  ( .D(creg_next[589]), .CLK(clk), .RST(rst), .I(m[589]), 
        .Q(c[589]) );
  DFF \creg_reg[590]  ( .D(creg_next[590]), .CLK(clk), .RST(rst), .I(m[590]), 
        .Q(c[590]) );
  DFF \creg_reg[591]  ( .D(creg_next[591]), .CLK(clk), .RST(rst), .I(m[591]), 
        .Q(c[591]) );
  DFF \creg_reg[592]  ( .D(creg_next[592]), .CLK(clk), .RST(rst), .I(m[592]), 
        .Q(c[592]) );
  DFF \creg_reg[593]  ( .D(creg_next[593]), .CLK(clk), .RST(rst), .I(m[593]), 
        .Q(c[593]) );
  DFF \creg_reg[594]  ( .D(creg_next[594]), .CLK(clk), .RST(rst), .I(m[594]), 
        .Q(c[594]) );
  DFF \creg_reg[595]  ( .D(creg_next[595]), .CLK(clk), .RST(rst), .I(m[595]), 
        .Q(c[595]) );
  DFF \creg_reg[596]  ( .D(creg_next[596]), .CLK(clk), .RST(rst), .I(m[596]), 
        .Q(c[596]) );
  DFF \creg_reg[597]  ( .D(creg_next[597]), .CLK(clk), .RST(rst), .I(m[597]), 
        .Q(c[597]) );
  DFF \creg_reg[598]  ( .D(creg_next[598]), .CLK(clk), .RST(rst), .I(m[598]), 
        .Q(c[598]) );
  DFF \creg_reg[599]  ( .D(creg_next[599]), .CLK(clk), .RST(rst), .I(m[599]), 
        .Q(c[599]) );
  DFF \creg_reg[600]  ( .D(creg_next[600]), .CLK(clk), .RST(rst), .I(m[600]), 
        .Q(c[600]) );
  DFF \creg_reg[601]  ( .D(creg_next[601]), .CLK(clk), .RST(rst), .I(m[601]), 
        .Q(c[601]) );
  DFF \creg_reg[602]  ( .D(creg_next[602]), .CLK(clk), .RST(rst), .I(m[602]), 
        .Q(c[602]) );
  DFF \creg_reg[603]  ( .D(creg_next[603]), .CLK(clk), .RST(rst), .I(m[603]), 
        .Q(c[603]) );
  DFF \creg_reg[604]  ( .D(creg_next[604]), .CLK(clk), .RST(rst), .I(m[604]), 
        .Q(c[604]) );
  DFF \creg_reg[605]  ( .D(creg_next[605]), .CLK(clk), .RST(rst), .I(m[605]), 
        .Q(c[605]) );
  DFF \creg_reg[606]  ( .D(creg_next[606]), .CLK(clk), .RST(rst), .I(m[606]), 
        .Q(c[606]) );
  DFF \creg_reg[607]  ( .D(creg_next[607]), .CLK(clk), .RST(rst), .I(m[607]), 
        .Q(c[607]) );
  DFF \creg_reg[608]  ( .D(creg_next[608]), .CLK(clk), .RST(rst), .I(m[608]), 
        .Q(c[608]) );
  DFF \creg_reg[609]  ( .D(creg_next[609]), .CLK(clk), .RST(rst), .I(m[609]), 
        .Q(c[609]) );
  DFF \creg_reg[610]  ( .D(creg_next[610]), .CLK(clk), .RST(rst), .I(m[610]), 
        .Q(c[610]) );
  DFF \creg_reg[611]  ( .D(creg_next[611]), .CLK(clk), .RST(rst), .I(m[611]), 
        .Q(c[611]) );
  DFF \creg_reg[612]  ( .D(creg_next[612]), .CLK(clk), .RST(rst), .I(m[612]), 
        .Q(c[612]) );
  DFF \creg_reg[613]  ( .D(creg_next[613]), .CLK(clk), .RST(rst), .I(m[613]), 
        .Q(c[613]) );
  DFF \creg_reg[614]  ( .D(creg_next[614]), .CLK(clk), .RST(rst), .I(m[614]), 
        .Q(c[614]) );
  DFF \creg_reg[615]  ( .D(creg_next[615]), .CLK(clk), .RST(rst), .I(m[615]), 
        .Q(c[615]) );
  DFF \creg_reg[616]  ( .D(creg_next[616]), .CLK(clk), .RST(rst), .I(m[616]), 
        .Q(c[616]) );
  DFF \creg_reg[617]  ( .D(creg_next[617]), .CLK(clk), .RST(rst), .I(m[617]), 
        .Q(c[617]) );
  DFF \creg_reg[618]  ( .D(creg_next[618]), .CLK(clk), .RST(rst), .I(m[618]), 
        .Q(c[618]) );
  DFF \creg_reg[619]  ( .D(creg_next[619]), .CLK(clk), .RST(rst), .I(m[619]), 
        .Q(c[619]) );
  DFF \creg_reg[620]  ( .D(creg_next[620]), .CLK(clk), .RST(rst), .I(m[620]), 
        .Q(c[620]) );
  DFF \creg_reg[621]  ( .D(creg_next[621]), .CLK(clk), .RST(rst), .I(m[621]), 
        .Q(c[621]) );
  DFF \creg_reg[622]  ( .D(creg_next[622]), .CLK(clk), .RST(rst), .I(m[622]), 
        .Q(c[622]) );
  DFF \creg_reg[623]  ( .D(creg_next[623]), .CLK(clk), .RST(rst), .I(m[623]), 
        .Q(c[623]) );
  DFF \creg_reg[624]  ( .D(creg_next[624]), .CLK(clk), .RST(rst), .I(m[624]), 
        .Q(c[624]) );
  DFF \creg_reg[625]  ( .D(creg_next[625]), .CLK(clk), .RST(rst), .I(m[625]), 
        .Q(c[625]) );
  DFF \creg_reg[626]  ( .D(creg_next[626]), .CLK(clk), .RST(rst), .I(m[626]), 
        .Q(c[626]) );
  DFF \creg_reg[627]  ( .D(creg_next[627]), .CLK(clk), .RST(rst), .I(m[627]), 
        .Q(c[627]) );
  DFF \creg_reg[628]  ( .D(creg_next[628]), .CLK(clk), .RST(rst), .I(m[628]), 
        .Q(c[628]) );
  DFF \creg_reg[629]  ( .D(creg_next[629]), .CLK(clk), .RST(rst), .I(m[629]), 
        .Q(c[629]) );
  DFF \creg_reg[630]  ( .D(creg_next[630]), .CLK(clk), .RST(rst), .I(m[630]), 
        .Q(c[630]) );
  DFF \creg_reg[631]  ( .D(creg_next[631]), .CLK(clk), .RST(rst), .I(m[631]), 
        .Q(c[631]) );
  DFF \creg_reg[632]  ( .D(creg_next[632]), .CLK(clk), .RST(rst), .I(m[632]), 
        .Q(c[632]) );
  DFF \creg_reg[633]  ( .D(creg_next[633]), .CLK(clk), .RST(rst), .I(m[633]), 
        .Q(c[633]) );
  DFF \creg_reg[634]  ( .D(creg_next[634]), .CLK(clk), .RST(rst), .I(m[634]), 
        .Q(c[634]) );
  DFF \creg_reg[635]  ( .D(creg_next[635]), .CLK(clk), .RST(rst), .I(m[635]), 
        .Q(c[635]) );
  DFF \creg_reg[636]  ( .D(creg_next[636]), .CLK(clk), .RST(rst), .I(m[636]), 
        .Q(c[636]) );
  DFF \creg_reg[637]  ( .D(creg_next[637]), .CLK(clk), .RST(rst), .I(m[637]), 
        .Q(c[637]) );
  DFF \creg_reg[638]  ( .D(creg_next[638]), .CLK(clk), .RST(rst), .I(m[638]), 
        .Q(c[638]) );
  DFF \creg_reg[639]  ( .D(creg_next[639]), .CLK(clk), .RST(rst), .I(m[639]), 
        .Q(c[639]) );
  DFF \creg_reg[640]  ( .D(creg_next[640]), .CLK(clk), .RST(rst), .I(m[640]), 
        .Q(c[640]) );
  DFF \creg_reg[641]  ( .D(creg_next[641]), .CLK(clk), .RST(rst), .I(m[641]), 
        .Q(c[641]) );
  DFF \creg_reg[642]  ( .D(creg_next[642]), .CLK(clk), .RST(rst), .I(m[642]), 
        .Q(c[642]) );
  DFF \creg_reg[643]  ( .D(creg_next[643]), .CLK(clk), .RST(rst), .I(m[643]), 
        .Q(c[643]) );
  DFF \creg_reg[644]  ( .D(creg_next[644]), .CLK(clk), .RST(rst), .I(m[644]), 
        .Q(c[644]) );
  DFF \creg_reg[645]  ( .D(creg_next[645]), .CLK(clk), .RST(rst), .I(m[645]), 
        .Q(c[645]) );
  DFF \creg_reg[646]  ( .D(creg_next[646]), .CLK(clk), .RST(rst), .I(m[646]), 
        .Q(c[646]) );
  DFF \creg_reg[647]  ( .D(creg_next[647]), .CLK(clk), .RST(rst), .I(m[647]), 
        .Q(c[647]) );
  DFF \creg_reg[648]  ( .D(creg_next[648]), .CLK(clk), .RST(rst), .I(m[648]), 
        .Q(c[648]) );
  DFF \creg_reg[649]  ( .D(creg_next[649]), .CLK(clk), .RST(rst), .I(m[649]), 
        .Q(c[649]) );
  DFF \creg_reg[650]  ( .D(creg_next[650]), .CLK(clk), .RST(rst), .I(m[650]), 
        .Q(c[650]) );
  DFF \creg_reg[651]  ( .D(creg_next[651]), .CLK(clk), .RST(rst), .I(m[651]), 
        .Q(c[651]) );
  DFF \creg_reg[652]  ( .D(creg_next[652]), .CLK(clk), .RST(rst), .I(m[652]), 
        .Q(c[652]) );
  DFF \creg_reg[653]  ( .D(creg_next[653]), .CLK(clk), .RST(rst), .I(m[653]), 
        .Q(c[653]) );
  DFF \creg_reg[654]  ( .D(creg_next[654]), .CLK(clk), .RST(rst), .I(m[654]), 
        .Q(c[654]) );
  DFF \creg_reg[655]  ( .D(creg_next[655]), .CLK(clk), .RST(rst), .I(m[655]), 
        .Q(c[655]) );
  DFF \creg_reg[656]  ( .D(creg_next[656]), .CLK(clk), .RST(rst), .I(m[656]), 
        .Q(c[656]) );
  DFF \creg_reg[657]  ( .D(creg_next[657]), .CLK(clk), .RST(rst), .I(m[657]), 
        .Q(c[657]) );
  DFF \creg_reg[658]  ( .D(creg_next[658]), .CLK(clk), .RST(rst), .I(m[658]), 
        .Q(c[658]) );
  DFF \creg_reg[659]  ( .D(creg_next[659]), .CLK(clk), .RST(rst), .I(m[659]), 
        .Q(c[659]) );
  DFF \creg_reg[660]  ( .D(creg_next[660]), .CLK(clk), .RST(rst), .I(m[660]), 
        .Q(c[660]) );
  DFF \creg_reg[661]  ( .D(creg_next[661]), .CLK(clk), .RST(rst), .I(m[661]), 
        .Q(c[661]) );
  DFF \creg_reg[662]  ( .D(creg_next[662]), .CLK(clk), .RST(rst), .I(m[662]), 
        .Q(c[662]) );
  DFF \creg_reg[663]  ( .D(creg_next[663]), .CLK(clk), .RST(rst), .I(m[663]), 
        .Q(c[663]) );
  DFF \creg_reg[664]  ( .D(creg_next[664]), .CLK(clk), .RST(rst), .I(m[664]), 
        .Q(c[664]) );
  DFF \creg_reg[665]  ( .D(creg_next[665]), .CLK(clk), .RST(rst), .I(m[665]), 
        .Q(c[665]) );
  DFF \creg_reg[666]  ( .D(creg_next[666]), .CLK(clk), .RST(rst), .I(m[666]), 
        .Q(c[666]) );
  DFF \creg_reg[667]  ( .D(creg_next[667]), .CLK(clk), .RST(rst), .I(m[667]), 
        .Q(c[667]) );
  DFF \creg_reg[668]  ( .D(creg_next[668]), .CLK(clk), .RST(rst), .I(m[668]), 
        .Q(c[668]) );
  DFF \creg_reg[669]  ( .D(creg_next[669]), .CLK(clk), .RST(rst), .I(m[669]), 
        .Q(c[669]) );
  DFF \creg_reg[670]  ( .D(creg_next[670]), .CLK(clk), .RST(rst), .I(m[670]), 
        .Q(c[670]) );
  DFF \creg_reg[671]  ( .D(creg_next[671]), .CLK(clk), .RST(rst), .I(m[671]), 
        .Q(c[671]) );
  DFF \creg_reg[672]  ( .D(creg_next[672]), .CLK(clk), .RST(rst), .I(m[672]), 
        .Q(c[672]) );
  DFF \creg_reg[673]  ( .D(creg_next[673]), .CLK(clk), .RST(rst), .I(m[673]), 
        .Q(c[673]) );
  DFF \creg_reg[674]  ( .D(creg_next[674]), .CLK(clk), .RST(rst), .I(m[674]), 
        .Q(c[674]) );
  DFF \creg_reg[675]  ( .D(creg_next[675]), .CLK(clk), .RST(rst), .I(m[675]), 
        .Q(c[675]) );
  DFF \creg_reg[676]  ( .D(creg_next[676]), .CLK(clk), .RST(rst), .I(m[676]), 
        .Q(c[676]) );
  DFF \creg_reg[677]  ( .D(creg_next[677]), .CLK(clk), .RST(rst), .I(m[677]), 
        .Q(c[677]) );
  DFF \creg_reg[678]  ( .D(creg_next[678]), .CLK(clk), .RST(rst), .I(m[678]), 
        .Q(c[678]) );
  DFF \creg_reg[679]  ( .D(creg_next[679]), .CLK(clk), .RST(rst), .I(m[679]), 
        .Q(c[679]) );
  DFF \creg_reg[680]  ( .D(creg_next[680]), .CLK(clk), .RST(rst), .I(m[680]), 
        .Q(c[680]) );
  DFF \creg_reg[681]  ( .D(creg_next[681]), .CLK(clk), .RST(rst), .I(m[681]), 
        .Q(c[681]) );
  DFF \creg_reg[682]  ( .D(creg_next[682]), .CLK(clk), .RST(rst), .I(m[682]), 
        .Q(c[682]) );
  DFF \creg_reg[683]  ( .D(creg_next[683]), .CLK(clk), .RST(rst), .I(m[683]), 
        .Q(c[683]) );
  DFF \creg_reg[684]  ( .D(creg_next[684]), .CLK(clk), .RST(rst), .I(m[684]), 
        .Q(c[684]) );
  DFF \creg_reg[685]  ( .D(creg_next[685]), .CLK(clk), .RST(rst), .I(m[685]), 
        .Q(c[685]) );
  DFF \creg_reg[686]  ( .D(creg_next[686]), .CLK(clk), .RST(rst), .I(m[686]), 
        .Q(c[686]) );
  DFF \creg_reg[687]  ( .D(creg_next[687]), .CLK(clk), .RST(rst), .I(m[687]), 
        .Q(c[687]) );
  DFF \creg_reg[688]  ( .D(creg_next[688]), .CLK(clk), .RST(rst), .I(m[688]), 
        .Q(c[688]) );
  DFF \creg_reg[689]  ( .D(creg_next[689]), .CLK(clk), .RST(rst), .I(m[689]), 
        .Q(c[689]) );
  DFF \creg_reg[690]  ( .D(creg_next[690]), .CLK(clk), .RST(rst), .I(m[690]), 
        .Q(c[690]) );
  DFF \creg_reg[691]  ( .D(creg_next[691]), .CLK(clk), .RST(rst), .I(m[691]), 
        .Q(c[691]) );
  DFF \creg_reg[692]  ( .D(creg_next[692]), .CLK(clk), .RST(rst), .I(m[692]), 
        .Q(c[692]) );
  DFF \creg_reg[693]  ( .D(creg_next[693]), .CLK(clk), .RST(rst), .I(m[693]), 
        .Q(c[693]) );
  DFF \creg_reg[694]  ( .D(creg_next[694]), .CLK(clk), .RST(rst), .I(m[694]), 
        .Q(c[694]) );
  DFF \creg_reg[695]  ( .D(creg_next[695]), .CLK(clk), .RST(rst), .I(m[695]), 
        .Q(c[695]) );
  DFF \creg_reg[696]  ( .D(creg_next[696]), .CLK(clk), .RST(rst), .I(m[696]), 
        .Q(c[696]) );
  DFF \creg_reg[697]  ( .D(creg_next[697]), .CLK(clk), .RST(rst), .I(m[697]), 
        .Q(c[697]) );
  DFF \creg_reg[698]  ( .D(creg_next[698]), .CLK(clk), .RST(rst), .I(m[698]), 
        .Q(c[698]) );
  DFF \creg_reg[699]  ( .D(creg_next[699]), .CLK(clk), .RST(rst), .I(m[699]), 
        .Q(c[699]) );
  DFF \creg_reg[700]  ( .D(creg_next[700]), .CLK(clk), .RST(rst), .I(m[700]), 
        .Q(c[700]) );
  DFF \creg_reg[701]  ( .D(creg_next[701]), .CLK(clk), .RST(rst), .I(m[701]), 
        .Q(c[701]) );
  DFF \creg_reg[702]  ( .D(creg_next[702]), .CLK(clk), .RST(rst), .I(m[702]), 
        .Q(c[702]) );
  DFF \creg_reg[703]  ( .D(creg_next[703]), .CLK(clk), .RST(rst), .I(m[703]), 
        .Q(c[703]) );
  DFF \creg_reg[704]  ( .D(creg_next[704]), .CLK(clk), .RST(rst), .I(m[704]), 
        .Q(c[704]) );
  DFF \creg_reg[705]  ( .D(creg_next[705]), .CLK(clk), .RST(rst), .I(m[705]), 
        .Q(c[705]) );
  DFF \creg_reg[706]  ( .D(creg_next[706]), .CLK(clk), .RST(rst), .I(m[706]), 
        .Q(c[706]) );
  DFF \creg_reg[707]  ( .D(creg_next[707]), .CLK(clk), .RST(rst), .I(m[707]), 
        .Q(c[707]) );
  DFF \creg_reg[708]  ( .D(creg_next[708]), .CLK(clk), .RST(rst), .I(m[708]), 
        .Q(c[708]) );
  DFF \creg_reg[709]  ( .D(creg_next[709]), .CLK(clk), .RST(rst), .I(m[709]), 
        .Q(c[709]) );
  DFF \creg_reg[710]  ( .D(creg_next[710]), .CLK(clk), .RST(rst), .I(m[710]), 
        .Q(c[710]) );
  DFF \creg_reg[711]  ( .D(creg_next[711]), .CLK(clk), .RST(rst), .I(m[711]), 
        .Q(c[711]) );
  DFF \creg_reg[712]  ( .D(creg_next[712]), .CLK(clk), .RST(rst), .I(m[712]), 
        .Q(c[712]) );
  DFF \creg_reg[713]  ( .D(creg_next[713]), .CLK(clk), .RST(rst), .I(m[713]), 
        .Q(c[713]) );
  DFF \creg_reg[714]  ( .D(creg_next[714]), .CLK(clk), .RST(rst), .I(m[714]), 
        .Q(c[714]) );
  DFF \creg_reg[715]  ( .D(creg_next[715]), .CLK(clk), .RST(rst), .I(m[715]), 
        .Q(c[715]) );
  DFF \creg_reg[716]  ( .D(creg_next[716]), .CLK(clk), .RST(rst), .I(m[716]), 
        .Q(c[716]) );
  DFF \creg_reg[717]  ( .D(creg_next[717]), .CLK(clk), .RST(rst), .I(m[717]), 
        .Q(c[717]) );
  DFF \creg_reg[718]  ( .D(creg_next[718]), .CLK(clk), .RST(rst), .I(m[718]), 
        .Q(c[718]) );
  DFF \creg_reg[719]  ( .D(creg_next[719]), .CLK(clk), .RST(rst), .I(m[719]), 
        .Q(c[719]) );
  DFF \creg_reg[720]  ( .D(creg_next[720]), .CLK(clk), .RST(rst), .I(m[720]), 
        .Q(c[720]) );
  DFF \creg_reg[721]  ( .D(creg_next[721]), .CLK(clk), .RST(rst), .I(m[721]), 
        .Q(c[721]) );
  DFF \creg_reg[722]  ( .D(creg_next[722]), .CLK(clk), .RST(rst), .I(m[722]), 
        .Q(c[722]) );
  DFF \creg_reg[723]  ( .D(creg_next[723]), .CLK(clk), .RST(rst), .I(m[723]), 
        .Q(c[723]) );
  DFF \creg_reg[724]  ( .D(creg_next[724]), .CLK(clk), .RST(rst), .I(m[724]), 
        .Q(c[724]) );
  DFF \creg_reg[725]  ( .D(creg_next[725]), .CLK(clk), .RST(rst), .I(m[725]), 
        .Q(c[725]) );
  DFF \creg_reg[726]  ( .D(creg_next[726]), .CLK(clk), .RST(rst), .I(m[726]), 
        .Q(c[726]) );
  DFF \creg_reg[727]  ( .D(creg_next[727]), .CLK(clk), .RST(rst), .I(m[727]), 
        .Q(c[727]) );
  DFF \creg_reg[728]  ( .D(creg_next[728]), .CLK(clk), .RST(rst), .I(m[728]), 
        .Q(c[728]) );
  DFF \creg_reg[729]  ( .D(creg_next[729]), .CLK(clk), .RST(rst), .I(m[729]), 
        .Q(c[729]) );
  DFF \creg_reg[730]  ( .D(creg_next[730]), .CLK(clk), .RST(rst), .I(m[730]), 
        .Q(c[730]) );
  DFF \creg_reg[731]  ( .D(creg_next[731]), .CLK(clk), .RST(rst), .I(m[731]), 
        .Q(c[731]) );
  DFF \creg_reg[732]  ( .D(creg_next[732]), .CLK(clk), .RST(rst), .I(m[732]), 
        .Q(c[732]) );
  DFF \creg_reg[733]  ( .D(creg_next[733]), .CLK(clk), .RST(rst), .I(m[733]), 
        .Q(c[733]) );
  DFF \creg_reg[734]  ( .D(creg_next[734]), .CLK(clk), .RST(rst), .I(m[734]), 
        .Q(c[734]) );
  DFF \creg_reg[735]  ( .D(creg_next[735]), .CLK(clk), .RST(rst), .I(m[735]), 
        .Q(c[735]) );
  DFF \creg_reg[736]  ( .D(creg_next[736]), .CLK(clk), .RST(rst), .I(m[736]), 
        .Q(c[736]) );
  DFF \creg_reg[737]  ( .D(creg_next[737]), .CLK(clk), .RST(rst), .I(m[737]), 
        .Q(c[737]) );
  DFF \creg_reg[738]  ( .D(creg_next[738]), .CLK(clk), .RST(rst), .I(m[738]), 
        .Q(c[738]) );
  DFF \creg_reg[739]  ( .D(creg_next[739]), .CLK(clk), .RST(rst), .I(m[739]), 
        .Q(c[739]) );
  DFF \creg_reg[740]  ( .D(creg_next[740]), .CLK(clk), .RST(rst), .I(m[740]), 
        .Q(c[740]) );
  DFF \creg_reg[741]  ( .D(creg_next[741]), .CLK(clk), .RST(rst), .I(m[741]), 
        .Q(c[741]) );
  DFF \creg_reg[742]  ( .D(creg_next[742]), .CLK(clk), .RST(rst), .I(m[742]), 
        .Q(c[742]) );
  DFF \creg_reg[743]  ( .D(creg_next[743]), .CLK(clk), .RST(rst), .I(m[743]), 
        .Q(c[743]) );
  DFF \creg_reg[744]  ( .D(creg_next[744]), .CLK(clk), .RST(rst), .I(m[744]), 
        .Q(c[744]) );
  DFF \creg_reg[745]  ( .D(creg_next[745]), .CLK(clk), .RST(rst), .I(m[745]), 
        .Q(c[745]) );
  DFF \creg_reg[746]  ( .D(creg_next[746]), .CLK(clk), .RST(rst), .I(m[746]), 
        .Q(c[746]) );
  DFF \creg_reg[747]  ( .D(creg_next[747]), .CLK(clk), .RST(rst), .I(m[747]), 
        .Q(c[747]) );
  DFF \creg_reg[748]  ( .D(creg_next[748]), .CLK(clk), .RST(rst), .I(m[748]), 
        .Q(c[748]) );
  DFF \creg_reg[749]  ( .D(creg_next[749]), .CLK(clk), .RST(rst), .I(m[749]), 
        .Q(c[749]) );
  DFF \creg_reg[750]  ( .D(creg_next[750]), .CLK(clk), .RST(rst), .I(m[750]), 
        .Q(c[750]) );
  DFF \creg_reg[751]  ( .D(creg_next[751]), .CLK(clk), .RST(rst), .I(m[751]), 
        .Q(c[751]) );
  DFF \creg_reg[752]  ( .D(creg_next[752]), .CLK(clk), .RST(rst), .I(m[752]), 
        .Q(c[752]) );
  DFF \creg_reg[753]  ( .D(creg_next[753]), .CLK(clk), .RST(rst), .I(m[753]), 
        .Q(c[753]) );
  DFF \creg_reg[754]  ( .D(creg_next[754]), .CLK(clk), .RST(rst), .I(m[754]), 
        .Q(c[754]) );
  DFF \creg_reg[755]  ( .D(creg_next[755]), .CLK(clk), .RST(rst), .I(m[755]), 
        .Q(c[755]) );
  DFF \creg_reg[756]  ( .D(creg_next[756]), .CLK(clk), .RST(rst), .I(m[756]), 
        .Q(c[756]) );
  DFF \creg_reg[757]  ( .D(creg_next[757]), .CLK(clk), .RST(rst), .I(m[757]), 
        .Q(c[757]) );
  DFF \creg_reg[758]  ( .D(creg_next[758]), .CLK(clk), .RST(rst), .I(m[758]), 
        .Q(c[758]) );
  DFF \creg_reg[759]  ( .D(creg_next[759]), .CLK(clk), .RST(rst), .I(m[759]), 
        .Q(c[759]) );
  DFF \creg_reg[760]  ( .D(creg_next[760]), .CLK(clk), .RST(rst), .I(m[760]), 
        .Q(c[760]) );
  DFF \creg_reg[761]  ( .D(creg_next[761]), .CLK(clk), .RST(rst), .I(m[761]), 
        .Q(c[761]) );
  DFF \creg_reg[762]  ( .D(creg_next[762]), .CLK(clk), .RST(rst), .I(m[762]), 
        .Q(c[762]) );
  DFF \creg_reg[763]  ( .D(creg_next[763]), .CLK(clk), .RST(rst), .I(m[763]), 
        .Q(c[763]) );
  DFF \creg_reg[764]  ( .D(creg_next[764]), .CLK(clk), .RST(rst), .I(m[764]), 
        .Q(c[764]) );
  DFF \creg_reg[765]  ( .D(creg_next[765]), .CLK(clk), .RST(rst), .I(m[765]), 
        .Q(c[765]) );
  DFF \creg_reg[766]  ( .D(creg_next[766]), .CLK(clk), .RST(rst), .I(m[766]), 
        .Q(c[766]) );
  DFF \creg_reg[767]  ( .D(creg_next[767]), .CLK(clk), .RST(rst), .I(m[767]), 
        .Q(c[767]) );
  DFF \creg_reg[768]  ( .D(creg_next[768]), .CLK(clk), .RST(rst), .I(m[768]), 
        .Q(c[768]) );
  DFF \creg_reg[769]  ( .D(creg_next[769]), .CLK(clk), .RST(rst), .I(m[769]), 
        .Q(c[769]) );
  DFF \creg_reg[770]  ( .D(creg_next[770]), .CLK(clk), .RST(rst), .I(m[770]), 
        .Q(c[770]) );
  DFF \creg_reg[771]  ( .D(creg_next[771]), .CLK(clk), .RST(rst), .I(m[771]), 
        .Q(c[771]) );
  DFF \creg_reg[772]  ( .D(creg_next[772]), .CLK(clk), .RST(rst), .I(m[772]), 
        .Q(c[772]) );
  DFF \creg_reg[773]  ( .D(creg_next[773]), .CLK(clk), .RST(rst), .I(m[773]), 
        .Q(c[773]) );
  DFF \creg_reg[774]  ( .D(creg_next[774]), .CLK(clk), .RST(rst), .I(m[774]), 
        .Q(c[774]) );
  DFF \creg_reg[775]  ( .D(creg_next[775]), .CLK(clk), .RST(rst), .I(m[775]), 
        .Q(c[775]) );
  DFF \creg_reg[776]  ( .D(creg_next[776]), .CLK(clk), .RST(rst), .I(m[776]), 
        .Q(c[776]) );
  DFF \creg_reg[777]  ( .D(creg_next[777]), .CLK(clk), .RST(rst), .I(m[777]), 
        .Q(c[777]) );
  DFF \creg_reg[778]  ( .D(creg_next[778]), .CLK(clk), .RST(rst), .I(m[778]), 
        .Q(c[778]) );
  DFF \creg_reg[779]  ( .D(creg_next[779]), .CLK(clk), .RST(rst), .I(m[779]), 
        .Q(c[779]) );
  DFF \creg_reg[780]  ( .D(creg_next[780]), .CLK(clk), .RST(rst), .I(m[780]), 
        .Q(c[780]) );
  DFF \creg_reg[781]  ( .D(creg_next[781]), .CLK(clk), .RST(rst), .I(m[781]), 
        .Q(c[781]) );
  DFF \creg_reg[782]  ( .D(creg_next[782]), .CLK(clk), .RST(rst), .I(m[782]), 
        .Q(c[782]) );
  DFF \creg_reg[783]  ( .D(creg_next[783]), .CLK(clk), .RST(rst), .I(m[783]), 
        .Q(c[783]) );
  DFF \creg_reg[784]  ( .D(creg_next[784]), .CLK(clk), .RST(rst), .I(m[784]), 
        .Q(c[784]) );
  DFF \creg_reg[785]  ( .D(creg_next[785]), .CLK(clk), .RST(rst), .I(m[785]), 
        .Q(c[785]) );
  DFF \creg_reg[786]  ( .D(creg_next[786]), .CLK(clk), .RST(rst), .I(m[786]), 
        .Q(c[786]) );
  DFF \creg_reg[787]  ( .D(creg_next[787]), .CLK(clk), .RST(rst), .I(m[787]), 
        .Q(c[787]) );
  DFF \creg_reg[788]  ( .D(creg_next[788]), .CLK(clk), .RST(rst), .I(m[788]), 
        .Q(c[788]) );
  DFF \creg_reg[789]  ( .D(creg_next[789]), .CLK(clk), .RST(rst), .I(m[789]), 
        .Q(c[789]) );
  DFF \creg_reg[790]  ( .D(creg_next[790]), .CLK(clk), .RST(rst), .I(m[790]), 
        .Q(c[790]) );
  DFF \creg_reg[791]  ( .D(creg_next[791]), .CLK(clk), .RST(rst), .I(m[791]), 
        .Q(c[791]) );
  DFF \creg_reg[792]  ( .D(creg_next[792]), .CLK(clk), .RST(rst), .I(m[792]), 
        .Q(c[792]) );
  DFF \creg_reg[793]  ( .D(creg_next[793]), .CLK(clk), .RST(rst), .I(m[793]), 
        .Q(c[793]) );
  DFF \creg_reg[794]  ( .D(creg_next[794]), .CLK(clk), .RST(rst), .I(m[794]), 
        .Q(c[794]) );
  DFF \creg_reg[795]  ( .D(creg_next[795]), .CLK(clk), .RST(rst), .I(m[795]), 
        .Q(c[795]) );
  DFF \creg_reg[796]  ( .D(creg_next[796]), .CLK(clk), .RST(rst), .I(m[796]), 
        .Q(c[796]) );
  DFF \creg_reg[797]  ( .D(creg_next[797]), .CLK(clk), .RST(rst), .I(m[797]), 
        .Q(c[797]) );
  DFF \creg_reg[798]  ( .D(creg_next[798]), .CLK(clk), .RST(rst), .I(m[798]), 
        .Q(c[798]) );
  DFF \creg_reg[799]  ( .D(creg_next[799]), .CLK(clk), .RST(rst), .I(m[799]), 
        .Q(c[799]) );
  DFF \creg_reg[800]  ( .D(creg_next[800]), .CLK(clk), .RST(rst), .I(m[800]), 
        .Q(c[800]) );
  DFF \creg_reg[801]  ( .D(creg_next[801]), .CLK(clk), .RST(rst), .I(m[801]), 
        .Q(c[801]) );
  DFF \creg_reg[802]  ( .D(creg_next[802]), .CLK(clk), .RST(rst), .I(m[802]), 
        .Q(c[802]) );
  DFF \creg_reg[803]  ( .D(creg_next[803]), .CLK(clk), .RST(rst), .I(m[803]), 
        .Q(c[803]) );
  DFF \creg_reg[804]  ( .D(creg_next[804]), .CLK(clk), .RST(rst), .I(m[804]), 
        .Q(c[804]) );
  DFF \creg_reg[805]  ( .D(creg_next[805]), .CLK(clk), .RST(rst), .I(m[805]), 
        .Q(c[805]) );
  DFF \creg_reg[806]  ( .D(creg_next[806]), .CLK(clk), .RST(rst), .I(m[806]), 
        .Q(c[806]) );
  DFF \creg_reg[807]  ( .D(creg_next[807]), .CLK(clk), .RST(rst), .I(m[807]), 
        .Q(c[807]) );
  DFF \creg_reg[808]  ( .D(creg_next[808]), .CLK(clk), .RST(rst), .I(m[808]), 
        .Q(c[808]) );
  DFF \creg_reg[809]  ( .D(creg_next[809]), .CLK(clk), .RST(rst), .I(m[809]), 
        .Q(c[809]) );
  DFF \creg_reg[810]  ( .D(creg_next[810]), .CLK(clk), .RST(rst), .I(m[810]), 
        .Q(c[810]) );
  DFF \creg_reg[811]  ( .D(creg_next[811]), .CLK(clk), .RST(rst), .I(m[811]), 
        .Q(c[811]) );
  DFF \creg_reg[812]  ( .D(creg_next[812]), .CLK(clk), .RST(rst), .I(m[812]), 
        .Q(c[812]) );
  DFF \creg_reg[813]  ( .D(creg_next[813]), .CLK(clk), .RST(rst), .I(m[813]), 
        .Q(c[813]) );
  DFF \creg_reg[814]  ( .D(creg_next[814]), .CLK(clk), .RST(rst), .I(m[814]), 
        .Q(c[814]) );
  DFF \creg_reg[815]  ( .D(creg_next[815]), .CLK(clk), .RST(rst), .I(m[815]), 
        .Q(c[815]) );
  DFF \creg_reg[816]  ( .D(creg_next[816]), .CLK(clk), .RST(rst), .I(m[816]), 
        .Q(c[816]) );
  DFF \creg_reg[817]  ( .D(creg_next[817]), .CLK(clk), .RST(rst), .I(m[817]), 
        .Q(c[817]) );
  DFF \creg_reg[818]  ( .D(creg_next[818]), .CLK(clk), .RST(rst), .I(m[818]), 
        .Q(c[818]) );
  DFF \creg_reg[819]  ( .D(creg_next[819]), .CLK(clk), .RST(rst), .I(m[819]), 
        .Q(c[819]) );
  DFF \creg_reg[820]  ( .D(creg_next[820]), .CLK(clk), .RST(rst), .I(m[820]), 
        .Q(c[820]) );
  DFF \creg_reg[821]  ( .D(creg_next[821]), .CLK(clk), .RST(rst), .I(m[821]), 
        .Q(c[821]) );
  DFF \creg_reg[822]  ( .D(creg_next[822]), .CLK(clk), .RST(rst), .I(m[822]), 
        .Q(c[822]) );
  DFF \creg_reg[823]  ( .D(creg_next[823]), .CLK(clk), .RST(rst), .I(m[823]), 
        .Q(c[823]) );
  DFF \creg_reg[824]  ( .D(creg_next[824]), .CLK(clk), .RST(rst), .I(m[824]), 
        .Q(c[824]) );
  DFF \creg_reg[825]  ( .D(creg_next[825]), .CLK(clk), .RST(rst), .I(m[825]), 
        .Q(c[825]) );
  DFF \creg_reg[826]  ( .D(creg_next[826]), .CLK(clk), .RST(rst), .I(m[826]), 
        .Q(c[826]) );
  DFF \creg_reg[827]  ( .D(creg_next[827]), .CLK(clk), .RST(rst), .I(m[827]), 
        .Q(c[827]) );
  DFF \creg_reg[828]  ( .D(creg_next[828]), .CLK(clk), .RST(rst), .I(m[828]), 
        .Q(c[828]) );
  DFF \creg_reg[829]  ( .D(creg_next[829]), .CLK(clk), .RST(rst), .I(m[829]), 
        .Q(c[829]) );
  DFF \creg_reg[830]  ( .D(creg_next[830]), .CLK(clk), .RST(rst), .I(m[830]), 
        .Q(c[830]) );
  DFF \creg_reg[831]  ( .D(creg_next[831]), .CLK(clk), .RST(rst), .I(m[831]), 
        .Q(c[831]) );
  DFF \creg_reg[832]  ( .D(creg_next[832]), .CLK(clk), .RST(rst), .I(m[832]), 
        .Q(c[832]) );
  DFF \creg_reg[833]  ( .D(creg_next[833]), .CLK(clk), .RST(rst), .I(m[833]), 
        .Q(c[833]) );
  DFF \creg_reg[834]  ( .D(creg_next[834]), .CLK(clk), .RST(rst), .I(m[834]), 
        .Q(c[834]) );
  DFF \creg_reg[835]  ( .D(creg_next[835]), .CLK(clk), .RST(rst), .I(m[835]), 
        .Q(c[835]) );
  DFF \creg_reg[836]  ( .D(creg_next[836]), .CLK(clk), .RST(rst), .I(m[836]), 
        .Q(c[836]) );
  DFF \creg_reg[837]  ( .D(creg_next[837]), .CLK(clk), .RST(rst), .I(m[837]), 
        .Q(c[837]) );
  DFF \creg_reg[838]  ( .D(creg_next[838]), .CLK(clk), .RST(rst), .I(m[838]), 
        .Q(c[838]) );
  DFF \creg_reg[839]  ( .D(creg_next[839]), .CLK(clk), .RST(rst), .I(m[839]), 
        .Q(c[839]) );
  DFF \creg_reg[840]  ( .D(creg_next[840]), .CLK(clk), .RST(rst), .I(m[840]), 
        .Q(c[840]) );
  DFF \creg_reg[841]  ( .D(creg_next[841]), .CLK(clk), .RST(rst), .I(m[841]), 
        .Q(c[841]) );
  DFF \creg_reg[842]  ( .D(creg_next[842]), .CLK(clk), .RST(rst), .I(m[842]), 
        .Q(c[842]) );
  DFF \creg_reg[843]  ( .D(creg_next[843]), .CLK(clk), .RST(rst), .I(m[843]), 
        .Q(c[843]) );
  DFF \creg_reg[844]  ( .D(creg_next[844]), .CLK(clk), .RST(rst), .I(m[844]), 
        .Q(c[844]) );
  DFF \creg_reg[845]  ( .D(creg_next[845]), .CLK(clk), .RST(rst), .I(m[845]), 
        .Q(c[845]) );
  DFF \creg_reg[846]  ( .D(creg_next[846]), .CLK(clk), .RST(rst), .I(m[846]), 
        .Q(c[846]) );
  DFF \creg_reg[847]  ( .D(creg_next[847]), .CLK(clk), .RST(rst), .I(m[847]), 
        .Q(c[847]) );
  DFF \creg_reg[848]  ( .D(creg_next[848]), .CLK(clk), .RST(rst), .I(m[848]), 
        .Q(c[848]) );
  DFF \creg_reg[849]  ( .D(creg_next[849]), .CLK(clk), .RST(rst), .I(m[849]), 
        .Q(c[849]) );
  DFF \creg_reg[850]  ( .D(creg_next[850]), .CLK(clk), .RST(rst), .I(m[850]), 
        .Q(c[850]) );
  DFF \creg_reg[851]  ( .D(creg_next[851]), .CLK(clk), .RST(rst), .I(m[851]), 
        .Q(c[851]) );
  DFF \creg_reg[852]  ( .D(creg_next[852]), .CLK(clk), .RST(rst), .I(m[852]), 
        .Q(c[852]) );
  DFF \creg_reg[853]  ( .D(creg_next[853]), .CLK(clk), .RST(rst), .I(m[853]), 
        .Q(c[853]) );
  DFF \creg_reg[854]  ( .D(creg_next[854]), .CLK(clk), .RST(rst), .I(m[854]), 
        .Q(c[854]) );
  DFF \creg_reg[855]  ( .D(creg_next[855]), .CLK(clk), .RST(rst), .I(m[855]), 
        .Q(c[855]) );
  DFF \creg_reg[856]  ( .D(creg_next[856]), .CLK(clk), .RST(rst), .I(m[856]), 
        .Q(c[856]) );
  DFF \creg_reg[857]  ( .D(creg_next[857]), .CLK(clk), .RST(rst), .I(m[857]), 
        .Q(c[857]) );
  DFF \creg_reg[858]  ( .D(creg_next[858]), .CLK(clk), .RST(rst), .I(m[858]), 
        .Q(c[858]) );
  DFF \creg_reg[859]  ( .D(creg_next[859]), .CLK(clk), .RST(rst), .I(m[859]), 
        .Q(c[859]) );
  DFF \creg_reg[860]  ( .D(creg_next[860]), .CLK(clk), .RST(rst), .I(m[860]), 
        .Q(c[860]) );
  DFF \creg_reg[861]  ( .D(creg_next[861]), .CLK(clk), .RST(rst), .I(m[861]), 
        .Q(c[861]) );
  DFF \creg_reg[862]  ( .D(creg_next[862]), .CLK(clk), .RST(rst), .I(m[862]), 
        .Q(c[862]) );
  DFF \creg_reg[863]  ( .D(creg_next[863]), .CLK(clk), .RST(rst), .I(m[863]), 
        .Q(c[863]) );
  DFF \creg_reg[864]  ( .D(creg_next[864]), .CLK(clk), .RST(rst), .I(m[864]), 
        .Q(c[864]) );
  DFF \creg_reg[865]  ( .D(creg_next[865]), .CLK(clk), .RST(rst), .I(m[865]), 
        .Q(c[865]) );
  DFF \creg_reg[866]  ( .D(creg_next[866]), .CLK(clk), .RST(rst), .I(m[866]), 
        .Q(c[866]) );
  DFF \creg_reg[867]  ( .D(creg_next[867]), .CLK(clk), .RST(rst), .I(m[867]), 
        .Q(c[867]) );
  DFF \creg_reg[868]  ( .D(creg_next[868]), .CLK(clk), .RST(rst), .I(m[868]), 
        .Q(c[868]) );
  DFF \creg_reg[869]  ( .D(creg_next[869]), .CLK(clk), .RST(rst), .I(m[869]), 
        .Q(c[869]) );
  DFF \creg_reg[870]  ( .D(creg_next[870]), .CLK(clk), .RST(rst), .I(m[870]), 
        .Q(c[870]) );
  DFF \creg_reg[871]  ( .D(creg_next[871]), .CLK(clk), .RST(rst), .I(m[871]), 
        .Q(c[871]) );
  DFF \creg_reg[872]  ( .D(creg_next[872]), .CLK(clk), .RST(rst), .I(m[872]), 
        .Q(c[872]) );
  DFF \creg_reg[873]  ( .D(creg_next[873]), .CLK(clk), .RST(rst), .I(m[873]), 
        .Q(c[873]) );
  DFF \creg_reg[874]  ( .D(creg_next[874]), .CLK(clk), .RST(rst), .I(m[874]), 
        .Q(c[874]) );
  DFF \creg_reg[875]  ( .D(creg_next[875]), .CLK(clk), .RST(rst), .I(m[875]), 
        .Q(c[875]) );
  DFF \creg_reg[876]  ( .D(creg_next[876]), .CLK(clk), .RST(rst), .I(m[876]), 
        .Q(c[876]) );
  DFF \creg_reg[877]  ( .D(creg_next[877]), .CLK(clk), .RST(rst), .I(m[877]), 
        .Q(c[877]) );
  DFF \creg_reg[878]  ( .D(creg_next[878]), .CLK(clk), .RST(rst), .I(m[878]), 
        .Q(c[878]) );
  DFF \creg_reg[879]  ( .D(creg_next[879]), .CLK(clk), .RST(rst), .I(m[879]), 
        .Q(c[879]) );
  DFF \creg_reg[880]  ( .D(creg_next[880]), .CLK(clk), .RST(rst), .I(m[880]), 
        .Q(c[880]) );
  DFF \creg_reg[881]  ( .D(creg_next[881]), .CLK(clk), .RST(rst), .I(m[881]), 
        .Q(c[881]) );
  DFF \creg_reg[882]  ( .D(creg_next[882]), .CLK(clk), .RST(rst), .I(m[882]), 
        .Q(c[882]) );
  DFF \creg_reg[883]  ( .D(creg_next[883]), .CLK(clk), .RST(rst), .I(m[883]), 
        .Q(c[883]) );
  DFF \creg_reg[884]  ( .D(creg_next[884]), .CLK(clk), .RST(rst), .I(m[884]), 
        .Q(c[884]) );
  DFF \creg_reg[885]  ( .D(creg_next[885]), .CLK(clk), .RST(rst), .I(m[885]), 
        .Q(c[885]) );
  DFF \creg_reg[886]  ( .D(creg_next[886]), .CLK(clk), .RST(rst), .I(m[886]), 
        .Q(c[886]) );
  DFF \creg_reg[887]  ( .D(creg_next[887]), .CLK(clk), .RST(rst), .I(m[887]), 
        .Q(c[887]) );
  DFF \creg_reg[888]  ( .D(creg_next[888]), .CLK(clk), .RST(rst), .I(m[888]), 
        .Q(c[888]) );
  DFF \creg_reg[889]  ( .D(creg_next[889]), .CLK(clk), .RST(rst), .I(m[889]), 
        .Q(c[889]) );
  DFF \creg_reg[890]  ( .D(creg_next[890]), .CLK(clk), .RST(rst), .I(m[890]), 
        .Q(c[890]) );
  DFF \creg_reg[891]  ( .D(creg_next[891]), .CLK(clk), .RST(rst), .I(m[891]), 
        .Q(c[891]) );
  DFF \creg_reg[892]  ( .D(creg_next[892]), .CLK(clk), .RST(rst), .I(m[892]), 
        .Q(c[892]) );
  DFF \creg_reg[893]  ( .D(creg_next[893]), .CLK(clk), .RST(rst), .I(m[893]), 
        .Q(c[893]) );
  DFF \creg_reg[894]  ( .D(creg_next[894]), .CLK(clk), .RST(rst), .I(m[894]), 
        .Q(c[894]) );
  DFF \creg_reg[895]  ( .D(creg_next[895]), .CLK(clk), .RST(rst), .I(m[895]), 
        .Q(c[895]) );
  DFF \creg_reg[896]  ( .D(creg_next[896]), .CLK(clk), .RST(rst), .I(m[896]), 
        .Q(c[896]) );
  DFF \creg_reg[897]  ( .D(creg_next[897]), .CLK(clk), .RST(rst), .I(m[897]), 
        .Q(c[897]) );
  DFF \creg_reg[898]  ( .D(creg_next[898]), .CLK(clk), .RST(rst), .I(m[898]), 
        .Q(c[898]) );
  DFF \creg_reg[899]  ( .D(creg_next[899]), .CLK(clk), .RST(rst), .I(m[899]), 
        .Q(c[899]) );
  DFF \creg_reg[900]  ( .D(creg_next[900]), .CLK(clk), .RST(rst), .I(m[900]), 
        .Q(c[900]) );
  DFF \creg_reg[901]  ( .D(creg_next[901]), .CLK(clk), .RST(rst), .I(m[901]), 
        .Q(c[901]) );
  DFF \creg_reg[902]  ( .D(creg_next[902]), .CLK(clk), .RST(rst), .I(m[902]), 
        .Q(c[902]) );
  DFF \creg_reg[903]  ( .D(creg_next[903]), .CLK(clk), .RST(rst), .I(m[903]), 
        .Q(c[903]) );
  DFF \creg_reg[904]  ( .D(creg_next[904]), .CLK(clk), .RST(rst), .I(m[904]), 
        .Q(c[904]) );
  DFF \creg_reg[905]  ( .D(creg_next[905]), .CLK(clk), .RST(rst), .I(m[905]), 
        .Q(c[905]) );
  DFF \creg_reg[906]  ( .D(creg_next[906]), .CLK(clk), .RST(rst), .I(m[906]), 
        .Q(c[906]) );
  DFF \creg_reg[907]  ( .D(creg_next[907]), .CLK(clk), .RST(rst), .I(m[907]), 
        .Q(c[907]) );
  DFF \creg_reg[908]  ( .D(creg_next[908]), .CLK(clk), .RST(rst), .I(m[908]), 
        .Q(c[908]) );
  DFF \creg_reg[909]  ( .D(creg_next[909]), .CLK(clk), .RST(rst), .I(m[909]), 
        .Q(c[909]) );
  DFF \creg_reg[910]  ( .D(creg_next[910]), .CLK(clk), .RST(rst), .I(m[910]), 
        .Q(c[910]) );
  DFF \creg_reg[911]  ( .D(creg_next[911]), .CLK(clk), .RST(rst), .I(m[911]), 
        .Q(c[911]) );
  DFF \creg_reg[912]  ( .D(creg_next[912]), .CLK(clk), .RST(rst), .I(m[912]), 
        .Q(c[912]) );
  DFF \creg_reg[913]  ( .D(creg_next[913]), .CLK(clk), .RST(rst), .I(m[913]), 
        .Q(c[913]) );
  DFF \creg_reg[914]  ( .D(creg_next[914]), .CLK(clk), .RST(rst), .I(m[914]), 
        .Q(c[914]) );
  DFF \creg_reg[915]  ( .D(creg_next[915]), .CLK(clk), .RST(rst), .I(m[915]), 
        .Q(c[915]) );
  DFF \creg_reg[916]  ( .D(creg_next[916]), .CLK(clk), .RST(rst), .I(m[916]), 
        .Q(c[916]) );
  DFF \creg_reg[917]  ( .D(creg_next[917]), .CLK(clk), .RST(rst), .I(m[917]), 
        .Q(c[917]) );
  DFF \creg_reg[918]  ( .D(creg_next[918]), .CLK(clk), .RST(rst), .I(m[918]), 
        .Q(c[918]) );
  DFF \creg_reg[919]  ( .D(creg_next[919]), .CLK(clk), .RST(rst), .I(m[919]), 
        .Q(c[919]) );
  DFF \creg_reg[920]  ( .D(creg_next[920]), .CLK(clk), .RST(rst), .I(m[920]), 
        .Q(c[920]) );
  DFF \creg_reg[921]  ( .D(creg_next[921]), .CLK(clk), .RST(rst), .I(m[921]), 
        .Q(c[921]) );
  DFF \creg_reg[922]  ( .D(creg_next[922]), .CLK(clk), .RST(rst), .I(m[922]), 
        .Q(c[922]) );
  DFF \creg_reg[923]  ( .D(creg_next[923]), .CLK(clk), .RST(rst), .I(m[923]), 
        .Q(c[923]) );
  DFF \creg_reg[924]  ( .D(creg_next[924]), .CLK(clk), .RST(rst), .I(m[924]), 
        .Q(c[924]) );
  DFF \creg_reg[925]  ( .D(creg_next[925]), .CLK(clk), .RST(rst), .I(m[925]), 
        .Q(c[925]) );
  DFF \creg_reg[926]  ( .D(creg_next[926]), .CLK(clk), .RST(rst), .I(m[926]), 
        .Q(c[926]) );
  DFF \creg_reg[927]  ( .D(creg_next[927]), .CLK(clk), .RST(rst), .I(m[927]), 
        .Q(c[927]) );
  DFF \creg_reg[928]  ( .D(creg_next[928]), .CLK(clk), .RST(rst), .I(m[928]), 
        .Q(c[928]) );
  DFF \creg_reg[929]  ( .D(creg_next[929]), .CLK(clk), .RST(rst), .I(m[929]), 
        .Q(c[929]) );
  DFF \creg_reg[930]  ( .D(creg_next[930]), .CLK(clk), .RST(rst), .I(m[930]), 
        .Q(c[930]) );
  DFF \creg_reg[931]  ( .D(creg_next[931]), .CLK(clk), .RST(rst), .I(m[931]), 
        .Q(c[931]) );
  DFF \creg_reg[932]  ( .D(creg_next[932]), .CLK(clk), .RST(rst), .I(m[932]), 
        .Q(c[932]) );
  DFF \creg_reg[933]  ( .D(creg_next[933]), .CLK(clk), .RST(rst), .I(m[933]), 
        .Q(c[933]) );
  DFF \creg_reg[934]  ( .D(creg_next[934]), .CLK(clk), .RST(rst), .I(m[934]), 
        .Q(c[934]) );
  DFF \creg_reg[935]  ( .D(creg_next[935]), .CLK(clk), .RST(rst), .I(m[935]), 
        .Q(c[935]) );
  DFF \creg_reg[936]  ( .D(creg_next[936]), .CLK(clk), .RST(rst), .I(m[936]), 
        .Q(c[936]) );
  DFF \creg_reg[937]  ( .D(creg_next[937]), .CLK(clk), .RST(rst), .I(m[937]), 
        .Q(c[937]) );
  DFF \creg_reg[938]  ( .D(creg_next[938]), .CLK(clk), .RST(rst), .I(m[938]), 
        .Q(c[938]) );
  DFF \creg_reg[939]  ( .D(creg_next[939]), .CLK(clk), .RST(rst), .I(m[939]), 
        .Q(c[939]) );
  DFF \creg_reg[940]  ( .D(creg_next[940]), .CLK(clk), .RST(rst), .I(m[940]), 
        .Q(c[940]) );
  DFF \creg_reg[941]  ( .D(creg_next[941]), .CLK(clk), .RST(rst), .I(m[941]), 
        .Q(c[941]) );
  DFF \creg_reg[942]  ( .D(creg_next[942]), .CLK(clk), .RST(rst), .I(m[942]), 
        .Q(c[942]) );
  DFF \creg_reg[943]  ( .D(creg_next[943]), .CLK(clk), .RST(rst), .I(m[943]), 
        .Q(c[943]) );
  DFF \creg_reg[944]  ( .D(creg_next[944]), .CLK(clk), .RST(rst), .I(m[944]), 
        .Q(c[944]) );
  DFF \creg_reg[945]  ( .D(creg_next[945]), .CLK(clk), .RST(rst), .I(m[945]), 
        .Q(c[945]) );
  DFF \creg_reg[946]  ( .D(creg_next[946]), .CLK(clk), .RST(rst), .I(m[946]), 
        .Q(c[946]) );
  DFF \creg_reg[947]  ( .D(creg_next[947]), .CLK(clk), .RST(rst), .I(m[947]), 
        .Q(c[947]) );
  DFF \creg_reg[948]  ( .D(creg_next[948]), .CLK(clk), .RST(rst), .I(m[948]), 
        .Q(c[948]) );
  DFF \creg_reg[949]  ( .D(creg_next[949]), .CLK(clk), .RST(rst), .I(m[949]), 
        .Q(c[949]) );
  DFF \creg_reg[950]  ( .D(creg_next[950]), .CLK(clk), .RST(rst), .I(m[950]), 
        .Q(c[950]) );
  DFF \creg_reg[951]  ( .D(creg_next[951]), .CLK(clk), .RST(rst), .I(m[951]), 
        .Q(c[951]) );
  DFF \creg_reg[952]  ( .D(creg_next[952]), .CLK(clk), .RST(rst), .I(m[952]), 
        .Q(c[952]) );
  DFF \creg_reg[953]  ( .D(creg_next[953]), .CLK(clk), .RST(rst), .I(m[953]), 
        .Q(c[953]) );
  DFF \creg_reg[954]  ( .D(creg_next[954]), .CLK(clk), .RST(rst), .I(m[954]), 
        .Q(c[954]) );
  DFF \creg_reg[955]  ( .D(creg_next[955]), .CLK(clk), .RST(rst), .I(m[955]), 
        .Q(c[955]) );
  DFF \creg_reg[956]  ( .D(creg_next[956]), .CLK(clk), .RST(rst), .I(m[956]), 
        .Q(c[956]) );
  DFF \creg_reg[957]  ( .D(creg_next[957]), .CLK(clk), .RST(rst), .I(m[957]), 
        .Q(c[957]) );
  DFF \creg_reg[958]  ( .D(creg_next[958]), .CLK(clk), .RST(rst), .I(m[958]), 
        .Q(c[958]) );
  DFF \creg_reg[959]  ( .D(creg_next[959]), .CLK(clk), .RST(rst), .I(m[959]), 
        .Q(c[959]) );
  DFF \creg_reg[960]  ( .D(creg_next[960]), .CLK(clk), .RST(rst), .I(m[960]), 
        .Q(c[960]) );
  DFF \creg_reg[961]  ( .D(creg_next[961]), .CLK(clk), .RST(rst), .I(m[961]), 
        .Q(c[961]) );
  DFF \creg_reg[962]  ( .D(creg_next[962]), .CLK(clk), .RST(rst), .I(m[962]), 
        .Q(c[962]) );
  DFF \creg_reg[963]  ( .D(creg_next[963]), .CLK(clk), .RST(rst), .I(m[963]), 
        .Q(c[963]) );
  DFF \creg_reg[964]  ( .D(creg_next[964]), .CLK(clk), .RST(rst), .I(m[964]), 
        .Q(c[964]) );
  DFF \creg_reg[965]  ( .D(creg_next[965]), .CLK(clk), .RST(rst), .I(m[965]), 
        .Q(c[965]) );
  DFF \creg_reg[966]  ( .D(creg_next[966]), .CLK(clk), .RST(rst), .I(m[966]), 
        .Q(c[966]) );
  DFF \creg_reg[967]  ( .D(creg_next[967]), .CLK(clk), .RST(rst), .I(m[967]), 
        .Q(c[967]) );
  DFF \creg_reg[968]  ( .D(creg_next[968]), .CLK(clk), .RST(rst), .I(m[968]), 
        .Q(c[968]) );
  DFF \creg_reg[969]  ( .D(creg_next[969]), .CLK(clk), .RST(rst), .I(m[969]), 
        .Q(c[969]) );
  DFF \creg_reg[970]  ( .D(creg_next[970]), .CLK(clk), .RST(rst), .I(m[970]), 
        .Q(c[970]) );
  DFF \creg_reg[971]  ( .D(creg_next[971]), .CLK(clk), .RST(rst), .I(m[971]), 
        .Q(c[971]) );
  DFF \creg_reg[972]  ( .D(creg_next[972]), .CLK(clk), .RST(rst), .I(m[972]), 
        .Q(c[972]) );
  DFF \creg_reg[973]  ( .D(creg_next[973]), .CLK(clk), .RST(rst), .I(m[973]), 
        .Q(c[973]) );
  DFF \creg_reg[974]  ( .D(creg_next[974]), .CLK(clk), .RST(rst), .I(m[974]), 
        .Q(c[974]) );
  DFF \creg_reg[975]  ( .D(creg_next[975]), .CLK(clk), .RST(rst), .I(m[975]), 
        .Q(c[975]) );
  DFF \creg_reg[976]  ( .D(creg_next[976]), .CLK(clk), .RST(rst), .I(m[976]), 
        .Q(c[976]) );
  DFF \creg_reg[977]  ( .D(creg_next[977]), .CLK(clk), .RST(rst), .I(m[977]), 
        .Q(c[977]) );
  DFF \creg_reg[978]  ( .D(creg_next[978]), .CLK(clk), .RST(rst), .I(m[978]), 
        .Q(c[978]) );
  DFF \creg_reg[979]  ( .D(creg_next[979]), .CLK(clk), .RST(rst), .I(m[979]), 
        .Q(c[979]) );
  DFF \creg_reg[980]  ( .D(creg_next[980]), .CLK(clk), .RST(rst), .I(m[980]), 
        .Q(c[980]) );
  DFF \creg_reg[981]  ( .D(creg_next[981]), .CLK(clk), .RST(rst), .I(m[981]), 
        .Q(c[981]) );
  DFF \creg_reg[982]  ( .D(creg_next[982]), .CLK(clk), .RST(rst), .I(m[982]), 
        .Q(c[982]) );
  DFF \creg_reg[983]  ( .D(creg_next[983]), .CLK(clk), .RST(rst), .I(m[983]), 
        .Q(c[983]) );
  DFF \creg_reg[984]  ( .D(creg_next[984]), .CLK(clk), .RST(rst), .I(m[984]), 
        .Q(c[984]) );
  DFF \creg_reg[985]  ( .D(creg_next[985]), .CLK(clk), .RST(rst), .I(m[985]), 
        .Q(c[985]) );
  DFF \creg_reg[986]  ( .D(creg_next[986]), .CLK(clk), .RST(rst), .I(m[986]), 
        .Q(c[986]) );
  DFF \creg_reg[987]  ( .D(creg_next[987]), .CLK(clk), .RST(rst), .I(m[987]), 
        .Q(c[987]) );
  DFF \creg_reg[988]  ( .D(creg_next[988]), .CLK(clk), .RST(rst), .I(m[988]), 
        .Q(c[988]) );
  DFF \creg_reg[989]  ( .D(creg_next[989]), .CLK(clk), .RST(rst), .I(m[989]), 
        .Q(c[989]) );
  DFF \creg_reg[990]  ( .D(creg_next[990]), .CLK(clk), .RST(rst), .I(m[990]), 
        .Q(c[990]) );
  DFF \creg_reg[991]  ( .D(creg_next[991]), .CLK(clk), .RST(rst), .I(m[991]), 
        .Q(c[991]) );
  DFF \creg_reg[992]  ( .D(creg_next[992]), .CLK(clk), .RST(rst), .I(m[992]), 
        .Q(c[992]) );
  DFF \creg_reg[993]  ( .D(creg_next[993]), .CLK(clk), .RST(rst), .I(m[993]), 
        .Q(c[993]) );
  DFF \creg_reg[994]  ( .D(creg_next[994]), .CLK(clk), .RST(rst), .I(m[994]), 
        .Q(c[994]) );
  DFF \creg_reg[995]  ( .D(creg_next[995]), .CLK(clk), .RST(rst), .I(m[995]), 
        .Q(c[995]) );
  DFF \creg_reg[996]  ( .D(creg_next[996]), .CLK(clk), .RST(rst), .I(m[996]), 
        .Q(c[996]) );
  DFF \creg_reg[997]  ( .D(creg_next[997]), .CLK(clk), .RST(rst), .I(m[997]), 
        .Q(c[997]) );
  DFF \creg_reg[998]  ( .D(creg_next[998]), .CLK(clk), .RST(rst), .I(m[998]), 
        .Q(c[998]) );
  DFF \creg_reg[999]  ( .D(creg_next[999]), .CLK(clk), .RST(rst), .I(m[999]), 
        .Q(c[999]) );
  DFF \creg_reg[1000]  ( .D(creg_next[1000]), .CLK(clk), .RST(rst), .I(m[1000]), .Q(c[1000]) );
  DFF \creg_reg[1001]  ( .D(creg_next[1001]), .CLK(clk), .RST(rst), .I(m[1001]), .Q(c[1001]) );
  DFF \creg_reg[1002]  ( .D(creg_next[1002]), .CLK(clk), .RST(rst), .I(m[1002]), .Q(c[1002]) );
  DFF \creg_reg[1003]  ( .D(creg_next[1003]), .CLK(clk), .RST(rst), .I(m[1003]), .Q(c[1003]) );
  DFF \creg_reg[1004]  ( .D(creg_next[1004]), .CLK(clk), .RST(rst), .I(m[1004]), .Q(c[1004]) );
  DFF \creg_reg[1005]  ( .D(creg_next[1005]), .CLK(clk), .RST(rst), .I(m[1005]), .Q(c[1005]) );
  DFF \creg_reg[1006]  ( .D(creg_next[1006]), .CLK(clk), .RST(rst), .I(m[1006]), .Q(c[1006]) );
  DFF \creg_reg[1007]  ( .D(creg_next[1007]), .CLK(clk), .RST(rst), .I(m[1007]), .Q(c[1007]) );
  DFF \creg_reg[1008]  ( .D(creg_next[1008]), .CLK(clk), .RST(rst), .I(m[1008]), .Q(c[1008]) );
  DFF \creg_reg[1009]  ( .D(creg_next[1009]), .CLK(clk), .RST(rst), .I(m[1009]), .Q(c[1009]) );
  DFF \creg_reg[1010]  ( .D(creg_next[1010]), .CLK(clk), .RST(rst), .I(m[1010]), .Q(c[1010]) );
  DFF \creg_reg[1011]  ( .D(creg_next[1011]), .CLK(clk), .RST(rst), .I(m[1011]), .Q(c[1011]) );
  DFF \creg_reg[1012]  ( .D(creg_next[1012]), .CLK(clk), .RST(rst), .I(m[1012]), .Q(c[1012]) );
  DFF \creg_reg[1013]  ( .D(creg_next[1013]), .CLK(clk), .RST(rst), .I(m[1013]), .Q(c[1013]) );
  DFF \creg_reg[1014]  ( .D(creg_next[1014]), .CLK(clk), .RST(rst), .I(m[1014]), .Q(c[1014]) );
  DFF \creg_reg[1015]  ( .D(creg_next[1015]), .CLK(clk), .RST(rst), .I(m[1015]), .Q(c[1015]) );
  DFF \creg_reg[1016]  ( .D(creg_next[1016]), .CLK(clk), .RST(rst), .I(m[1016]), .Q(c[1016]) );
  DFF \creg_reg[1017]  ( .D(creg_next[1017]), .CLK(clk), .RST(rst), .I(m[1017]), .Q(c[1017]) );
  DFF \creg_reg[1018]  ( .D(creg_next[1018]), .CLK(clk), .RST(rst), .I(m[1018]), .Q(c[1018]) );
  DFF \creg_reg[1019]  ( .D(creg_next[1019]), .CLK(clk), .RST(rst), .I(m[1019]), .Q(c[1019]) );
  DFF \creg_reg[1020]  ( .D(creg_next[1020]), .CLK(clk), .RST(rst), .I(m[1020]), .Q(c[1020]) );
  DFF \creg_reg[1021]  ( .D(creg_next[1021]), .CLK(clk), .RST(rst), .I(m[1021]), .Q(c[1021]) );
  DFF \creg_reg[1022]  ( .D(creg_next[1022]), .CLK(clk), .RST(rst), .I(m[1022]), .Q(c[1022]) );
  DFF \creg_reg[1023]  ( .D(creg_next[1023]), .CLK(clk), .RST(rst), .I(m[1023]), .Q(c[1023]) );
  XOR U1036 ( .A(start_in[1023]), .B(mul_pow), .Z(n8) );
  NANDN U1037 ( .A(first_one), .B(n1033), .Z(n6) );
  NAND U1038 ( .A(n1034), .B(ein[1023]), .Z(n1033) );
  AND U1039 ( .A(mul_pow), .B(start_in[1023]), .Z(n1034) );
  NAND U1040 ( .A(n1035), .B(n1036), .Z(_0_net_) );
  NANDN U1041 ( .A(mul_pow), .B(first_one), .Z(n1036) );
  NAND U1042 ( .A(first_one), .B(ein[1023]), .Z(n1035) );
endmodule

