
module modmult_step_N1024_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [1025:0] A;
  input [1025:0] B;
  output [1025:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120;

  IV U1 ( .A(n5119), .Z(n1) );
  IV U2 ( .A(A[1]), .Z(n2) );
  XNOR U3 ( .A(n3), .B(n4), .Z(DIFF[9]) );
  XOR U4 ( .A(B[9]), .B(A[9]), .Z(n4) );
  XNOR U5 ( .A(n5), .B(n6), .Z(DIFF[99]) );
  XOR U6 ( .A(B[99]), .B(A[99]), .Z(n6) );
  XNOR U7 ( .A(n7), .B(n8), .Z(DIFF[999]) );
  XOR U8 ( .A(B[999]), .B(A[999]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(DIFF[998]) );
  XOR U10 ( .A(B[998]), .B(A[998]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(DIFF[997]) );
  XOR U12 ( .A(B[997]), .B(A[997]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(DIFF[996]) );
  XOR U14 ( .A(B[996]), .B(A[996]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(DIFF[995]) );
  XOR U16 ( .A(B[995]), .B(A[995]), .Z(n16) );
  XOR U17 ( .A(n17), .B(n18), .Z(DIFF[994]) );
  XOR U18 ( .A(B[994]), .B(A[994]), .Z(n18) );
  XOR U19 ( .A(n19), .B(n20), .Z(DIFF[993]) );
  XOR U20 ( .A(B[993]), .B(A[993]), .Z(n20) );
  XOR U21 ( .A(n21), .B(n22), .Z(DIFF[992]) );
  XOR U22 ( .A(B[992]), .B(A[992]), .Z(n22) );
  XOR U23 ( .A(n23), .B(n24), .Z(DIFF[991]) );
  XOR U24 ( .A(B[991]), .B(A[991]), .Z(n24) );
  XOR U25 ( .A(n25), .B(n26), .Z(DIFF[990]) );
  XOR U26 ( .A(B[990]), .B(A[990]), .Z(n26) );
  XOR U27 ( .A(n27), .B(n28), .Z(DIFF[98]) );
  XOR U28 ( .A(B[98]), .B(A[98]), .Z(n28) );
  XOR U29 ( .A(n29), .B(n30), .Z(DIFF[989]) );
  XOR U30 ( .A(B[989]), .B(A[989]), .Z(n30) );
  XOR U31 ( .A(n31), .B(n32), .Z(DIFF[988]) );
  XOR U32 ( .A(B[988]), .B(A[988]), .Z(n32) );
  XOR U33 ( .A(n33), .B(n34), .Z(DIFF[987]) );
  XOR U34 ( .A(B[987]), .B(A[987]), .Z(n34) );
  XOR U35 ( .A(n35), .B(n36), .Z(DIFF[986]) );
  XOR U36 ( .A(B[986]), .B(A[986]), .Z(n36) );
  XOR U37 ( .A(n37), .B(n38), .Z(DIFF[985]) );
  XOR U38 ( .A(B[985]), .B(A[985]), .Z(n38) );
  XOR U39 ( .A(n39), .B(n40), .Z(DIFF[984]) );
  XOR U40 ( .A(B[984]), .B(A[984]), .Z(n40) );
  XOR U41 ( .A(n41), .B(n42), .Z(DIFF[983]) );
  XOR U42 ( .A(B[983]), .B(A[983]), .Z(n42) );
  XOR U43 ( .A(n43), .B(n44), .Z(DIFF[982]) );
  XOR U44 ( .A(B[982]), .B(A[982]), .Z(n44) );
  XOR U45 ( .A(n45), .B(n46), .Z(DIFF[981]) );
  XOR U46 ( .A(B[981]), .B(A[981]), .Z(n46) );
  XOR U47 ( .A(n47), .B(n48), .Z(DIFF[980]) );
  XOR U48 ( .A(B[980]), .B(A[980]), .Z(n48) );
  XOR U49 ( .A(n49), .B(n50), .Z(DIFF[97]) );
  XOR U50 ( .A(B[97]), .B(A[97]), .Z(n50) );
  XOR U51 ( .A(n51), .B(n52), .Z(DIFF[979]) );
  XOR U52 ( .A(B[979]), .B(A[979]), .Z(n52) );
  XOR U53 ( .A(n53), .B(n54), .Z(DIFF[978]) );
  XOR U54 ( .A(B[978]), .B(A[978]), .Z(n54) );
  XOR U55 ( .A(n55), .B(n56), .Z(DIFF[977]) );
  XOR U56 ( .A(B[977]), .B(A[977]), .Z(n56) );
  XOR U57 ( .A(n57), .B(n58), .Z(DIFF[976]) );
  XOR U58 ( .A(B[976]), .B(A[976]), .Z(n58) );
  XOR U59 ( .A(n59), .B(n60), .Z(DIFF[975]) );
  XOR U60 ( .A(B[975]), .B(A[975]), .Z(n60) );
  XOR U61 ( .A(n61), .B(n62), .Z(DIFF[974]) );
  XOR U62 ( .A(B[974]), .B(A[974]), .Z(n62) );
  XOR U63 ( .A(n63), .B(n64), .Z(DIFF[973]) );
  XOR U64 ( .A(B[973]), .B(A[973]), .Z(n64) );
  XOR U65 ( .A(n65), .B(n66), .Z(DIFF[972]) );
  XOR U66 ( .A(B[972]), .B(A[972]), .Z(n66) );
  XOR U67 ( .A(n67), .B(n68), .Z(DIFF[971]) );
  XOR U68 ( .A(B[971]), .B(A[971]), .Z(n68) );
  XOR U69 ( .A(n69), .B(n70), .Z(DIFF[970]) );
  XOR U70 ( .A(B[970]), .B(A[970]), .Z(n70) );
  XOR U71 ( .A(n71), .B(n72), .Z(DIFF[96]) );
  XOR U72 ( .A(B[96]), .B(A[96]), .Z(n72) );
  XOR U73 ( .A(n73), .B(n74), .Z(DIFF[969]) );
  XOR U74 ( .A(B[969]), .B(A[969]), .Z(n74) );
  XOR U75 ( .A(n75), .B(n76), .Z(DIFF[968]) );
  XOR U76 ( .A(B[968]), .B(A[968]), .Z(n76) );
  XOR U77 ( .A(n77), .B(n78), .Z(DIFF[967]) );
  XOR U78 ( .A(B[967]), .B(A[967]), .Z(n78) );
  XOR U79 ( .A(n79), .B(n80), .Z(DIFF[966]) );
  XOR U80 ( .A(B[966]), .B(A[966]), .Z(n80) );
  XOR U81 ( .A(n81), .B(n82), .Z(DIFF[965]) );
  XOR U82 ( .A(B[965]), .B(A[965]), .Z(n82) );
  XOR U83 ( .A(n83), .B(n84), .Z(DIFF[964]) );
  XOR U84 ( .A(B[964]), .B(A[964]), .Z(n84) );
  XOR U85 ( .A(n85), .B(n86), .Z(DIFF[963]) );
  XOR U86 ( .A(B[963]), .B(A[963]), .Z(n86) );
  XOR U87 ( .A(n87), .B(n88), .Z(DIFF[962]) );
  XOR U88 ( .A(B[962]), .B(A[962]), .Z(n88) );
  XOR U89 ( .A(n89), .B(n90), .Z(DIFF[961]) );
  XOR U90 ( .A(B[961]), .B(A[961]), .Z(n90) );
  XOR U91 ( .A(n91), .B(n92), .Z(DIFF[960]) );
  XOR U92 ( .A(B[960]), .B(A[960]), .Z(n92) );
  XOR U93 ( .A(n93), .B(n94), .Z(DIFF[95]) );
  XOR U94 ( .A(B[95]), .B(A[95]), .Z(n94) );
  XOR U95 ( .A(n95), .B(n96), .Z(DIFF[959]) );
  XOR U96 ( .A(B[959]), .B(A[959]), .Z(n96) );
  XOR U97 ( .A(n97), .B(n98), .Z(DIFF[958]) );
  XOR U98 ( .A(B[958]), .B(A[958]), .Z(n98) );
  XOR U99 ( .A(n99), .B(n100), .Z(DIFF[957]) );
  XOR U100 ( .A(B[957]), .B(A[957]), .Z(n100) );
  XOR U101 ( .A(n101), .B(n102), .Z(DIFF[956]) );
  XOR U102 ( .A(B[956]), .B(A[956]), .Z(n102) );
  XOR U103 ( .A(n103), .B(n104), .Z(DIFF[955]) );
  XOR U104 ( .A(B[955]), .B(A[955]), .Z(n104) );
  XOR U105 ( .A(n105), .B(n106), .Z(DIFF[954]) );
  XOR U106 ( .A(B[954]), .B(A[954]), .Z(n106) );
  XOR U107 ( .A(n107), .B(n108), .Z(DIFF[953]) );
  XOR U108 ( .A(B[953]), .B(A[953]), .Z(n108) );
  XOR U109 ( .A(n109), .B(n110), .Z(DIFF[952]) );
  XOR U110 ( .A(B[952]), .B(A[952]), .Z(n110) );
  XOR U111 ( .A(n111), .B(n112), .Z(DIFF[951]) );
  XOR U112 ( .A(B[951]), .B(A[951]), .Z(n112) );
  XOR U113 ( .A(n113), .B(n114), .Z(DIFF[950]) );
  XOR U114 ( .A(B[950]), .B(A[950]), .Z(n114) );
  XOR U115 ( .A(n115), .B(n116), .Z(DIFF[94]) );
  XOR U116 ( .A(B[94]), .B(A[94]), .Z(n116) );
  XOR U117 ( .A(n117), .B(n118), .Z(DIFF[949]) );
  XOR U118 ( .A(B[949]), .B(A[949]), .Z(n118) );
  XOR U119 ( .A(n119), .B(n120), .Z(DIFF[948]) );
  XOR U120 ( .A(B[948]), .B(A[948]), .Z(n120) );
  XOR U121 ( .A(n121), .B(n122), .Z(DIFF[947]) );
  XOR U122 ( .A(B[947]), .B(A[947]), .Z(n122) );
  XOR U123 ( .A(n123), .B(n124), .Z(DIFF[946]) );
  XOR U124 ( .A(B[946]), .B(A[946]), .Z(n124) );
  XOR U125 ( .A(n125), .B(n126), .Z(DIFF[945]) );
  XOR U126 ( .A(B[945]), .B(A[945]), .Z(n126) );
  XOR U127 ( .A(n127), .B(n128), .Z(DIFF[944]) );
  XOR U128 ( .A(B[944]), .B(A[944]), .Z(n128) );
  XOR U129 ( .A(n129), .B(n130), .Z(DIFF[943]) );
  XOR U130 ( .A(B[943]), .B(A[943]), .Z(n130) );
  XOR U131 ( .A(n131), .B(n132), .Z(DIFF[942]) );
  XOR U132 ( .A(B[942]), .B(A[942]), .Z(n132) );
  XOR U133 ( .A(n133), .B(n134), .Z(DIFF[941]) );
  XOR U134 ( .A(B[941]), .B(A[941]), .Z(n134) );
  XOR U135 ( .A(n135), .B(n136), .Z(DIFF[940]) );
  XOR U136 ( .A(B[940]), .B(A[940]), .Z(n136) );
  XOR U137 ( .A(n137), .B(n138), .Z(DIFF[93]) );
  XOR U138 ( .A(B[93]), .B(A[93]), .Z(n138) );
  XOR U139 ( .A(n139), .B(n140), .Z(DIFF[939]) );
  XOR U140 ( .A(B[939]), .B(A[939]), .Z(n140) );
  XOR U141 ( .A(n141), .B(n142), .Z(DIFF[938]) );
  XOR U142 ( .A(B[938]), .B(A[938]), .Z(n142) );
  XOR U143 ( .A(n143), .B(n144), .Z(DIFF[937]) );
  XOR U144 ( .A(B[937]), .B(A[937]), .Z(n144) );
  XOR U145 ( .A(n145), .B(n146), .Z(DIFF[936]) );
  XOR U146 ( .A(B[936]), .B(A[936]), .Z(n146) );
  XOR U147 ( .A(n147), .B(n148), .Z(DIFF[935]) );
  XOR U148 ( .A(B[935]), .B(A[935]), .Z(n148) );
  XOR U149 ( .A(n149), .B(n150), .Z(DIFF[934]) );
  XOR U150 ( .A(B[934]), .B(A[934]), .Z(n150) );
  XOR U151 ( .A(n151), .B(n152), .Z(DIFF[933]) );
  XOR U152 ( .A(B[933]), .B(A[933]), .Z(n152) );
  XOR U153 ( .A(n153), .B(n154), .Z(DIFF[932]) );
  XOR U154 ( .A(B[932]), .B(A[932]), .Z(n154) );
  XOR U155 ( .A(n155), .B(n156), .Z(DIFF[931]) );
  XOR U156 ( .A(B[931]), .B(A[931]), .Z(n156) );
  XOR U157 ( .A(n157), .B(n158), .Z(DIFF[930]) );
  XOR U158 ( .A(B[930]), .B(A[930]), .Z(n158) );
  XOR U159 ( .A(n159), .B(n160), .Z(DIFF[92]) );
  XOR U160 ( .A(B[92]), .B(A[92]), .Z(n160) );
  XOR U161 ( .A(n161), .B(n162), .Z(DIFF[929]) );
  XOR U162 ( .A(B[929]), .B(A[929]), .Z(n162) );
  XOR U163 ( .A(n163), .B(n164), .Z(DIFF[928]) );
  XOR U164 ( .A(B[928]), .B(A[928]), .Z(n164) );
  XOR U165 ( .A(n165), .B(n166), .Z(DIFF[927]) );
  XOR U166 ( .A(B[927]), .B(A[927]), .Z(n166) );
  XOR U167 ( .A(n167), .B(n168), .Z(DIFF[926]) );
  XOR U168 ( .A(B[926]), .B(A[926]), .Z(n168) );
  XOR U169 ( .A(n169), .B(n170), .Z(DIFF[925]) );
  XOR U170 ( .A(B[925]), .B(A[925]), .Z(n170) );
  XOR U171 ( .A(n171), .B(n172), .Z(DIFF[924]) );
  XOR U172 ( .A(B[924]), .B(A[924]), .Z(n172) );
  XOR U173 ( .A(n173), .B(n174), .Z(DIFF[923]) );
  XOR U174 ( .A(B[923]), .B(A[923]), .Z(n174) );
  XOR U175 ( .A(n175), .B(n176), .Z(DIFF[922]) );
  XOR U176 ( .A(B[922]), .B(A[922]), .Z(n176) );
  XOR U177 ( .A(n177), .B(n178), .Z(DIFF[921]) );
  XOR U178 ( .A(B[921]), .B(A[921]), .Z(n178) );
  XOR U179 ( .A(n179), .B(n180), .Z(DIFF[920]) );
  XOR U180 ( .A(B[920]), .B(A[920]), .Z(n180) );
  XOR U181 ( .A(n181), .B(n182), .Z(DIFF[91]) );
  XOR U182 ( .A(B[91]), .B(A[91]), .Z(n182) );
  XOR U183 ( .A(n183), .B(n184), .Z(DIFF[919]) );
  XOR U184 ( .A(B[919]), .B(A[919]), .Z(n184) );
  XOR U185 ( .A(n185), .B(n186), .Z(DIFF[918]) );
  XOR U186 ( .A(B[918]), .B(A[918]), .Z(n186) );
  XOR U187 ( .A(n187), .B(n188), .Z(DIFF[917]) );
  XOR U188 ( .A(B[917]), .B(A[917]), .Z(n188) );
  XOR U189 ( .A(n189), .B(n190), .Z(DIFF[916]) );
  XOR U190 ( .A(B[916]), .B(A[916]), .Z(n190) );
  XOR U191 ( .A(n191), .B(n192), .Z(DIFF[915]) );
  XOR U192 ( .A(B[915]), .B(A[915]), .Z(n192) );
  XOR U193 ( .A(n193), .B(n194), .Z(DIFF[914]) );
  XOR U194 ( .A(B[914]), .B(A[914]), .Z(n194) );
  XOR U195 ( .A(n195), .B(n196), .Z(DIFF[913]) );
  XOR U196 ( .A(B[913]), .B(A[913]), .Z(n196) );
  XOR U197 ( .A(n197), .B(n198), .Z(DIFF[912]) );
  XOR U198 ( .A(B[912]), .B(A[912]), .Z(n198) );
  XOR U199 ( .A(n199), .B(n200), .Z(DIFF[911]) );
  XOR U200 ( .A(B[911]), .B(A[911]), .Z(n200) );
  XOR U201 ( .A(n201), .B(n202), .Z(DIFF[910]) );
  XOR U202 ( .A(B[910]), .B(A[910]), .Z(n202) );
  XOR U203 ( .A(n203), .B(n204), .Z(DIFF[90]) );
  XOR U204 ( .A(B[90]), .B(A[90]), .Z(n204) );
  XOR U205 ( .A(n205), .B(n206), .Z(DIFF[909]) );
  XOR U206 ( .A(B[909]), .B(A[909]), .Z(n206) );
  XOR U207 ( .A(n207), .B(n208), .Z(DIFF[908]) );
  XOR U208 ( .A(B[908]), .B(A[908]), .Z(n208) );
  XOR U209 ( .A(n209), .B(n210), .Z(DIFF[907]) );
  XOR U210 ( .A(B[907]), .B(A[907]), .Z(n210) );
  XOR U211 ( .A(n211), .B(n212), .Z(DIFF[906]) );
  XOR U212 ( .A(B[906]), .B(A[906]), .Z(n212) );
  XOR U213 ( .A(n213), .B(n214), .Z(DIFF[905]) );
  XOR U214 ( .A(B[905]), .B(A[905]), .Z(n214) );
  XOR U215 ( .A(n215), .B(n216), .Z(DIFF[904]) );
  XOR U216 ( .A(B[904]), .B(A[904]), .Z(n216) );
  XOR U217 ( .A(n217), .B(n218), .Z(DIFF[903]) );
  XOR U218 ( .A(B[903]), .B(A[903]), .Z(n218) );
  XOR U219 ( .A(n219), .B(n220), .Z(DIFF[902]) );
  XOR U220 ( .A(B[902]), .B(A[902]), .Z(n220) );
  XOR U221 ( .A(n221), .B(n222), .Z(DIFF[901]) );
  XOR U222 ( .A(B[901]), .B(A[901]), .Z(n222) );
  XOR U223 ( .A(n223), .B(n224), .Z(DIFF[900]) );
  XOR U224 ( .A(B[900]), .B(A[900]), .Z(n224) );
  XOR U225 ( .A(n225), .B(n226), .Z(DIFF[8]) );
  XOR U226 ( .A(B[8]), .B(A[8]), .Z(n226) );
  XOR U227 ( .A(n227), .B(n228), .Z(DIFF[89]) );
  XOR U228 ( .A(B[89]), .B(A[89]), .Z(n228) );
  XOR U229 ( .A(n229), .B(n230), .Z(DIFF[899]) );
  XOR U230 ( .A(B[899]), .B(A[899]), .Z(n230) );
  XOR U231 ( .A(n231), .B(n232), .Z(DIFF[898]) );
  XOR U232 ( .A(B[898]), .B(A[898]), .Z(n232) );
  XOR U233 ( .A(n233), .B(n234), .Z(DIFF[897]) );
  XOR U234 ( .A(B[897]), .B(A[897]), .Z(n234) );
  XOR U235 ( .A(n235), .B(n236), .Z(DIFF[896]) );
  XOR U236 ( .A(B[896]), .B(A[896]), .Z(n236) );
  XOR U237 ( .A(n237), .B(n238), .Z(DIFF[895]) );
  XOR U238 ( .A(B[895]), .B(A[895]), .Z(n238) );
  XOR U239 ( .A(n239), .B(n240), .Z(DIFF[894]) );
  XOR U240 ( .A(B[894]), .B(A[894]), .Z(n240) );
  XOR U241 ( .A(n241), .B(n242), .Z(DIFF[893]) );
  XOR U242 ( .A(B[893]), .B(A[893]), .Z(n242) );
  XOR U243 ( .A(n243), .B(n244), .Z(DIFF[892]) );
  XOR U244 ( .A(B[892]), .B(A[892]), .Z(n244) );
  XOR U245 ( .A(n245), .B(n246), .Z(DIFF[891]) );
  XOR U246 ( .A(B[891]), .B(A[891]), .Z(n246) );
  XOR U247 ( .A(n247), .B(n248), .Z(DIFF[890]) );
  XOR U248 ( .A(B[890]), .B(A[890]), .Z(n248) );
  XOR U249 ( .A(n249), .B(n250), .Z(DIFF[88]) );
  XOR U250 ( .A(B[88]), .B(A[88]), .Z(n250) );
  XOR U251 ( .A(n251), .B(n252), .Z(DIFF[889]) );
  XOR U252 ( .A(B[889]), .B(A[889]), .Z(n252) );
  XOR U253 ( .A(n253), .B(n254), .Z(DIFF[888]) );
  XOR U254 ( .A(B[888]), .B(A[888]), .Z(n254) );
  XOR U255 ( .A(n255), .B(n256), .Z(DIFF[887]) );
  XOR U256 ( .A(B[887]), .B(A[887]), .Z(n256) );
  XOR U257 ( .A(n257), .B(n258), .Z(DIFF[886]) );
  XOR U258 ( .A(B[886]), .B(A[886]), .Z(n258) );
  XOR U259 ( .A(n259), .B(n260), .Z(DIFF[885]) );
  XOR U260 ( .A(B[885]), .B(A[885]), .Z(n260) );
  XOR U261 ( .A(n261), .B(n262), .Z(DIFF[884]) );
  XOR U262 ( .A(B[884]), .B(A[884]), .Z(n262) );
  XOR U263 ( .A(n263), .B(n264), .Z(DIFF[883]) );
  XOR U264 ( .A(B[883]), .B(A[883]), .Z(n264) );
  XOR U265 ( .A(n265), .B(n266), .Z(DIFF[882]) );
  XOR U266 ( .A(B[882]), .B(A[882]), .Z(n266) );
  XOR U267 ( .A(n267), .B(n268), .Z(DIFF[881]) );
  XOR U268 ( .A(B[881]), .B(A[881]), .Z(n268) );
  XOR U269 ( .A(n269), .B(n270), .Z(DIFF[880]) );
  XOR U270 ( .A(B[880]), .B(A[880]), .Z(n270) );
  XOR U271 ( .A(n271), .B(n272), .Z(DIFF[87]) );
  XOR U272 ( .A(B[87]), .B(A[87]), .Z(n272) );
  XOR U273 ( .A(n273), .B(n274), .Z(DIFF[879]) );
  XOR U274 ( .A(B[879]), .B(A[879]), .Z(n274) );
  XOR U275 ( .A(n275), .B(n276), .Z(DIFF[878]) );
  XOR U276 ( .A(B[878]), .B(A[878]), .Z(n276) );
  XOR U277 ( .A(n277), .B(n278), .Z(DIFF[877]) );
  XOR U278 ( .A(B[877]), .B(A[877]), .Z(n278) );
  XOR U279 ( .A(n279), .B(n280), .Z(DIFF[876]) );
  XOR U280 ( .A(B[876]), .B(A[876]), .Z(n280) );
  XOR U281 ( .A(n281), .B(n282), .Z(DIFF[875]) );
  XOR U282 ( .A(B[875]), .B(A[875]), .Z(n282) );
  XOR U283 ( .A(n283), .B(n284), .Z(DIFF[874]) );
  XOR U284 ( .A(B[874]), .B(A[874]), .Z(n284) );
  XOR U285 ( .A(n285), .B(n286), .Z(DIFF[873]) );
  XOR U286 ( .A(B[873]), .B(A[873]), .Z(n286) );
  XOR U287 ( .A(n287), .B(n288), .Z(DIFF[872]) );
  XOR U288 ( .A(B[872]), .B(A[872]), .Z(n288) );
  XOR U289 ( .A(n289), .B(n290), .Z(DIFF[871]) );
  XOR U290 ( .A(B[871]), .B(A[871]), .Z(n290) );
  XOR U291 ( .A(n291), .B(n292), .Z(DIFF[870]) );
  XOR U292 ( .A(B[870]), .B(A[870]), .Z(n292) );
  XOR U293 ( .A(n293), .B(n294), .Z(DIFF[86]) );
  XOR U294 ( .A(B[86]), .B(A[86]), .Z(n294) );
  XOR U295 ( .A(n295), .B(n296), .Z(DIFF[869]) );
  XOR U296 ( .A(B[869]), .B(A[869]), .Z(n296) );
  XOR U297 ( .A(n297), .B(n298), .Z(DIFF[868]) );
  XOR U298 ( .A(B[868]), .B(A[868]), .Z(n298) );
  XOR U299 ( .A(n299), .B(n300), .Z(DIFF[867]) );
  XOR U300 ( .A(B[867]), .B(A[867]), .Z(n300) );
  XOR U301 ( .A(n301), .B(n302), .Z(DIFF[866]) );
  XOR U302 ( .A(B[866]), .B(A[866]), .Z(n302) );
  XOR U303 ( .A(n303), .B(n304), .Z(DIFF[865]) );
  XOR U304 ( .A(B[865]), .B(A[865]), .Z(n304) );
  XOR U305 ( .A(n305), .B(n306), .Z(DIFF[864]) );
  XOR U306 ( .A(B[864]), .B(A[864]), .Z(n306) );
  XOR U307 ( .A(n307), .B(n308), .Z(DIFF[863]) );
  XOR U308 ( .A(B[863]), .B(A[863]), .Z(n308) );
  XOR U309 ( .A(n309), .B(n310), .Z(DIFF[862]) );
  XOR U310 ( .A(B[862]), .B(A[862]), .Z(n310) );
  XOR U311 ( .A(n311), .B(n312), .Z(DIFF[861]) );
  XOR U312 ( .A(B[861]), .B(A[861]), .Z(n312) );
  XOR U313 ( .A(n313), .B(n314), .Z(DIFF[860]) );
  XOR U314 ( .A(B[860]), .B(A[860]), .Z(n314) );
  XOR U315 ( .A(n315), .B(n316), .Z(DIFF[85]) );
  XOR U316 ( .A(B[85]), .B(A[85]), .Z(n316) );
  XOR U317 ( .A(n317), .B(n318), .Z(DIFF[859]) );
  XOR U318 ( .A(B[859]), .B(A[859]), .Z(n318) );
  XOR U319 ( .A(n319), .B(n320), .Z(DIFF[858]) );
  XOR U320 ( .A(B[858]), .B(A[858]), .Z(n320) );
  XOR U321 ( .A(n321), .B(n322), .Z(DIFF[857]) );
  XOR U322 ( .A(B[857]), .B(A[857]), .Z(n322) );
  XOR U323 ( .A(n323), .B(n324), .Z(DIFF[856]) );
  XOR U324 ( .A(B[856]), .B(A[856]), .Z(n324) );
  XOR U325 ( .A(n325), .B(n326), .Z(DIFF[855]) );
  XOR U326 ( .A(B[855]), .B(A[855]), .Z(n326) );
  XOR U327 ( .A(n327), .B(n328), .Z(DIFF[854]) );
  XOR U328 ( .A(B[854]), .B(A[854]), .Z(n328) );
  XOR U329 ( .A(n329), .B(n330), .Z(DIFF[853]) );
  XOR U330 ( .A(B[853]), .B(A[853]), .Z(n330) );
  XOR U331 ( .A(n331), .B(n332), .Z(DIFF[852]) );
  XOR U332 ( .A(B[852]), .B(A[852]), .Z(n332) );
  XOR U333 ( .A(n333), .B(n334), .Z(DIFF[851]) );
  XOR U334 ( .A(B[851]), .B(A[851]), .Z(n334) );
  XOR U335 ( .A(n335), .B(n336), .Z(DIFF[850]) );
  XOR U336 ( .A(B[850]), .B(A[850]), .Z(n336) );
  XOR U337 ( .A(n337), .B(n338), .Z(DIFF[84]) );
  XOR U338 ( .A(B[84]), .B(A[84]), .Z(n338) );
  XOR U339 ( .A(n339), .B(n340), .Z(DIFF[849]) );
  XOR U340 ( .A(B[849]), .B(A[849]), .Z(n340) );
  XOR U341 ( .A(n341), .B(n342), .Z(DIFF[848]) );
  XOR U342 ( .A(B[848]), .B(A[848]), .Z(n342) );
  XOR U343 ( .A(n343), .B(n344), .Z(DIFF[847]) );
  XOR U344 ( .A(B[847]), .B(A[847]), .Z(n344) );
  XOR U345 ( .A(n345), .B(n346), .Z(DIFF[846]) );
  XOR U346 ( .A(B[846]), .B(A[846]), .Z(n346) );
  XOR U347 ( .A(n347), .B(n348), .Z(DIFF[845]) );
  XOR U348 ( .A(B[845]), .B(A[845]), .Z(n348) );
  XOR U349 ( .A(n349), .B(n350), .Z(DIFF[844]) );
  XOR U350 ( .A(B[844]), .B(A[844]), .Z(n350) );
  XOR U351 ( .A(n351), .B(n352), .Z(DIFF[843]) );
  XOR U352 ( .A(B[843]), .B(A[843]), .Z(n352) );
  XOR U353 ( .A(n353), .B(n354), .Z(DIFF[842]) );
  XOR U354 ( .A(B[842]), .B(A[842]), .Z(n354) );
  XOR U355 ( .A(n355), .B(n356), .Z(DIFF[841]) );
  XOR U356 ( .A(B[841]), .B(A[841]), .Z(n356) );
  XOR U357 ( .A(n357), .B(n358), .Z(DIFF[840]) );
  XOR U358 ( .A(B[840]), .B(A[840]), .Z(n358) );
  XOR U359 ( .A(n359), .B(n360), .Z(DIFF[83]) );
  XOR U360 ( .A(B[83]), .B(A[83]), .Z(n360) );
  XOR U361 ( .A(n361), .B(n362), .Z(DIFF[839]) );
  XOR U362 ( .A(B[839]), .B(A[839]), .Z(n362) );
  XOR U363 ( .A(n363), .B(n364), .Z(DIFF[838]) );
  XOR U364 ( .A(B[838]), .B(A[838]), .Z(n364) );
  XOR U365 ( .A(n365), .B(n366), .Z(DIFF[837]) );
  XOR U366 ( .A(B[837]), .B(A[837]), .Z(n366) );
  XOR U367 ( .A(n367), .B(n368), .Z(DIFF[836]) );
  XOR U368 ( .A(B[836]), .B(A[836]), .Z(n368) );
  XOR U369 ( .A(n369), .B(n370), .Z(DIFF[835]) );
  XOR U370 ( .A(B[835]), .B(A[835]), .Z(n370) );
  XOR U371 ( .A(n371), .B(n372), .Z(DIFF[834]) );
  XOR U372 ( .A(B[834]), .B(A[834]), .Z(n372) );
  XOR U373 ( .A(n373), .B(n374), .Z(DIFF[833]) );
  XOR U374 ( .A(B[833]), .B(A[833]), .Z(n374) );
  XOR U375 ( .A(n375), .B(n376), .Z(DIFF[832]) );
  XOR U376 ( .A(B[832]), .B(A[832]), .Z(n376) );
  XOR U377 ( .A(n377), .B(n378), .Z(DIFF[831]) );
  XOR U378 ( .A(B[831]), .B(A[831]), .Z(n378) );
  XOR U379 ( .A(n379), .B(n380), .Z(DIFF[830]) );
  XOR U380 ( .A(B[830]), .B(A[830]), .Z(n380) );
  XOR U381 ( .A(n381), .B(n382), .Z(DIFF[82]) );
  XOR U382 ( .A(B[82]), .B(A[82]), .Z(n382) );
  XOR U383 ( .A(n383), .B(n384), .Z(DIFF[829]) );
  XOR U384 ( .A(B[829]), .B(A[829]), .Z(n384) );
  XOR U385 ( .A(n385), .B(n386), .Z(DIFF[828]) );
  XOR U386 ( .A(B[828]), .B(A[828]), .Z(n386) );
  XOR U387 ( .A(n387), .B(n388), .Z(DIFF[827]) );
  XOR U388 ( .A(B[827]), .B(A[827]), .Z(n388) );
  XOR U389 ( .A(n389), .B(n390), .Z(DIFF[826]) );
  XOR U390 ( .A(B[826]), .B(A[826]), .Z(n390) );
  XOR U391 ( .A(n391), .B(n392), .Z(DIFF[825]) );
  XOR U392 ( .A(B[825]), .B(A[825]), .Z(n392) );
  XOR U393 ( .A(n393), .B(n394), .Z(DIFF[824]) );
  XOR U394 ( .A(B[824]), .B(A[824]), .Z(n394) );
  XOR U395 ( .A(n395), .B(n396), .Z(DIFF[823]) );
  XOR U396 ( .A(B[823]), .B(A[823]), .Z(n396) );
  XOR U397 ( .A(n397), .B(n398), .Z(DIFF[822]) );
  XOR U398 ( .A(B[822]), .B(A[822]), .Z(n398) );
  XOR U399 ( .A(n399), .B(n400), .Z(DIFF[821]) );
  XOR U400 ( .A(B[821]), .B(A[821]), .Z(n400) );
  XOR U401 ( .A(n401), .B(n402), .Z(DIFF[820]) );
  XOR U402 ( .A(B[820]), .B(A[820]), .Z(n402) );
  XOR U403 ( .A(n403), .B(n404), .Z(DIFF[81]) );
  XOR U404 ( .A(B[81]), .B(A[81]), .Z(n404) );
  XOR U405 ( .A(n405), .B(n406), .Z(DIFF[819]) );
  XOR U406 ( .A(B[819]), .B(A[819]), .Z(n406) );
  XOR U407 ( .A(n407), .B(n408), .Z(DIFF[818]) );
  XOR U408 ( .A(B[818]), .B(A[818]), .Z(n408) );
  XOR U409 ( .A(n409), .B(n410), .Z(DIFF[817]) );
  XOR U410 ( .A(B[817]), .B(A[817]), .Z(n410) );
  XOR U411 ( .A(n411), .B(n412), .Z(DIFF[816]) );
  XOR U412 ( .A(B[816]), .B(A[816]), .Z(n412) );
  XOR U413 ( .A(n413), .B(n414), .Z(DIFF[815]) );
  XOR U414 ( .A(B[815]), .B(A[815]), .Z(n414) );
  XOR U415 ( .A(n415), .B(n416), .Z(DIFF[814]) );
  XOR U416 ( .A(B[814]), .B(A[814]), .Z(n416) );
  XOR U417 ( .A(n417), .B(n418), .Z(DIFF[813]) );
  XOR U418 ( .A(B[813]), .B(A[813]), .Z(n418) );
  XOR U419 ( .A(n419), .B(n420), .Z(DIFF[812]) );
  XOR U420 ( .A(B[812]), .B(A[812]), .Z(n420) );
  XOR U421 ( .A(n421), .B(n422), .Z(DIFF[811]) );
  XOR U422 ( .A(B[811]), .B(A[811]), .Z(n422) );
  XOR U423 ( .A(n423), .B(n424), .Z(DIFF[810]) );
  XOR U424 ( .A(B[810]), .B(A[810]), .Z(n424) );
  XOR U425 ( .A(n425), .B(n426), .Z(DIFF[80]) );
  XOR U426 ( .A(B[80]), .B(A[80]), .Z(n426) );
  XOR U427 ( .A(n427), .B(n428), .Z(DIFF[809]) );
  XOR U428 ( .A(B[809]), .B(A[809]), .Z(n428) );
  XOR U429 ( .A(n429), .B(n430), .Z(DIFF[808]) );
  XOR U430 ( .A(B[808]), .B(A[808]), .Z(n430) );
  XOR U431 ( .A(n431), .B(n432), .Z(DIFF[807]) );
  XOR U432 ( .A(B[807]), .B(A[807]), .Z(n432) );
  XOR U433 ( .A(n433), .B(n434), .Z(DIFF[806]) );
  XOR U434 ( .A(B[806]), .B(A[806]), .Z(n434) );
  XOR U435 ( .A(n435), .B(n436), .Z(DIFF[805]) );
  XOR U436 ( .A(B[805]), .B(A[805]), .Z(n436) );
  XOR U437 ( .A(n437), .B(n438), .Z(DIFF[804]) );
  XOR U438 ( .A(B[804]), .B(A[804]), .Z(n438) );
  XOR U439 ( .A(n439), .B(n440), .Z(DIFF[803]) );
  XOR U440 ( .A(B[803]), .B(A[803]), .Z(n440) );
  XOR U441 ( .A(n441), .B(n442), .Z(DIFF[802]) );
  XOR U442 ( .A(B[802]), .B(A[802]), .Z(n442) );
  XOR U443 ( .A(n443), .B(n444), .Z(DIFF[801]) );
  XOR U444 ( .A(B[801]), .B(A[801]), .Z(n444) );
  XOR U445 ( .A(n445), .B(n446), .Z(DIFF[800]) );
  XOR U446 ( .A(B[800]), .B(A[800]), .Z(n446) );
  XOR U447 ( .A(n447), .B(n448), .Z(DIFF[7]) );
  XOR U448 ( .A(B[7]), .B(A[7]), .Z(n448) );
  XOR U449 ( .A(n449), .B(n450), .Z(DIFF[79]) );
  XOR U450 ( .A(B[79]), .B(A[79]), .Z(n450) );
  XOR U451 ( .A(n451), .B(n452), .Z(DIFF[799]) );
  XOR U452 ( .A(B[799]), .B(A[799]), .Z(n452) );
  XOR U453 ( .A(n453), .B(n454), .Z(DIFF[798]) );
  XOR U454 ( .A(B[798]), .B(A[798]), .Z(n454) );
  XOR U455 ( .A(n455), .B(n456), .Z(DIFF[797]) );
  XOR U456 ( .A(B[797]), .B(A[797]), .Z(n456) );
  XOR U457 ( .A(n457), .B(n458), .Z(DIFF[796]) );
  XOR U458 ( .A(B[796]), .B(A[796]), .Z(n458) );
  XOR U459 ( .A(n459), .B(n460), .Z(DIFF[795]) );
  XOR U460 ( .A(B[795]), .B(A[795]), .Z(n460) );
  XOR U461 ( .A(n461), .B(n462), .Z(DIFF[794]) );
  XOR U462 ( .A(B[794]), .B(A[794]), .Z(n462) );
  XOR U463 ( .A(n463), .B(n464), .Z(DIFF[793]) );
  XOR U464 ( .A(B[793]), .B(A[793]), .Z(n464) );
  XOR U465 ( .A(n465), .B(n466), .Z(DIFF[792]) );
  XOR U466 ( .A(B[792]), .B(A[792]), .Z(n466) );
  XOR U467 ( .A(n467), .B(n468), .Z(DIFF[791]) );
  XOR U468 ( .A(B[791]), .B(A[791]), .Z(n468) );
  XOR U469 ( .A(n469), .B(n470), .Z(DIFF[790]) );
  XOR U470 ( .A(B[790]), .B(A[790]), .Z(n470) );
  XOR U471 ( .A(n471), .B(n472), .Z(DIFF[78]) );
  XOR U472 ( .A(B[78]), .B(A[78]), .Z(n472) );
  XOR U473 ( .A(n473), .B(n474), .Z(DIFF[789]) );
  XOR U474 ( .A(B[789]), .B(A[789]), .Z(n474) );
  XOR U475 ( .A(n475), .B(n476), .Z(DIFF[788]) );
  XOR U476 ( .A(B[788]), .B(A[788]), .Z(n476) );
  XOR U477 ( .A(n477), .B(n478), .Z(DIFF[787]) );
  XOR U478 ( .A(B[787]), .B(A[787]), .Z(n478) );
  XOR U479 ( .A(n479), .B(n480), .Z(DIFF[786]) );
  XOR U480 ( .A(B[786]), .B(A[786]), .Z(n480) );
  XOR U481 ( .A(n481), .B(n482), .Z(DIFF[785]) );
  XOR U482 ( .A(B[785]), .B(A[785]), .Z(n482) );
  XOR U483 ( .A(n483), .B(n484), .Z(DIFF[784]) );
  XOR U484 ( .A(B[784]), .B(A[784]), .Z(n484) );
  XOR U485 ( .A(n485), .B(n486), .Z(DIFF[783]) );
  XOR U486 ( .A(B[783]), .B(A[783]), .Z(n486) );
  XOR U487 ( .A(n487), .B(n488), .Z(DIFF[782]) );
  XOR U488 ( .A(B[782]), .B(A[782]), .Z(n488) );
  XOR U489 ( .A(n489), .B(n490), .Z(DIFF[781]) );
  XOR U490 ( .A(B[781]), .B(A[781]), .Z(n490) );
  XOR U491 ( .A(n491), .B(n492), .Z(DIFF[780]) );
  XOR U492 ( .A(B[780]), .B(A[780]), .Z(n492) );
  XOR U493 ( .A(n493), .B(n494), .Z(DIFF[77]) );
  XOR U494 ( .A(B[77]), .B(A[77]), .Z(n494) );
  XOR U495 ( .A(n495), .B(n496), .Z(DIFF[779]) );
  XOR U496 ( .A(B[779]), .B(A[779]), .Z(n496) );
  XOR U497 ( .A(n497), .B(n498), .Z(DIFF[778]) );
  XOR U498 ( .A(B[778]), .B(A[778]), .Z(n498) );
  XOR U499 ( .A(n499), .B(n500), .Z(DIFF[777]) );
  XOR U500 ( .A(B[777]), .B(A[777]), .Z(n500) );
  XOR U501 ( .A(n501), .B(n502), .Z(DIFF[776]) );
  XOR U502 ( .A(B[776]), .B(A[776]), .Z(n502) );
  XOR U503 ( .A(n503), .B(n504), .Z(DIFF[775]) );
  XOR U504 ( .A(B[775]), .B(A[775]), .Z(n504) );
  XOR U505 ( .A(n505), .B(n506), .Z(DIFF[774]) );
  XOR U506 ( .A(B[774]), .B(A[774]), .Z(n506) );
  XOR U507 ( .A(n507), .B(n508), .Z(DIFF[773]) );
  XOR U508 ( .A(B[773]), .B(A[773]), .Z(n508) );
  XOR U509 ( .A(n509), .B(n510), .Z(DIFF[772]) );
  XOR U510 ( .A(B[772]), .B(A[772]), .Z(n510) );
  XOR U511 ( .A(n511), .B(n512), .Z(DIFF[771]) );
  XOR U512 ( .A(B[771]), .B(A[771]), .Z(n512) );
  XOR U513 ( .A(n513), .B(n514), .Z(DIFF[770]) );
  XOR U514 ( .A(B[770]), .B(A[770]), .Z(n514) );
  XOR U515 ( .A(n515), .B(n516), .Z(DIFF[76]) );
  XOR U516 ( .A(B[76]), .B(A[76]), .Z(n516) );
  XOR U517 ( .A(n517), .B(n518), .Z(DIFF[769]) );
  XOR U518 ( .A(B[769]), .B(A[769]), .Z(n518) );
  XOR U519 ( .A(n519), .B(n520), .Z(DIFF[768]) );
  XOR U520 ( .A(B[768]), .B(A[768]), .Z(n520) );
  XOR U521 ( .A(n521), .B(n522), .Z(DIFF[767]) );
  XOR U522 ( .A(B[767]), .B(A[767]), .Z(n522) );
  XOR U523 ( .A(n523), .B(n524), .Z(DIFF[766]) );
  XOR U524 ( .A(B[766]), .B(A[766]), .Z(n524) );
  XOR U525 ( .A(n525), .B(n526), .Z(DIFF[765]) );
  XOR U526 ( .A(B[765]), .B(A[765]), .Z(n526) );
  XOR U527 ( .A(n527), .B(n528), .Z(DIFF[764]) );
  XOR U528 ( .A(B[764]), .B(A[764]), .Z(n528) );
  XOR U529 ( .A(n529), .B(n530), .Z(DIFF[763]) );
  XOR U530 ( .A(B[763]), .B(A[763]), .Z(n530) );
  XOR U531 ( .A(n531), .B(n532), .Z(DIFF[762]) );
  XOR U532 ( .A(B[762]), .B(A[762]), .Z(n532) );
  XOR U533 ( .A(n533), .B(n534), .Z(DIFF[761]) );
  XOR U534 ( .A(B[761]), .B(A[761]), .Z(n534) );
  XOR U535 ( .A(n535), .B(n536), .Z(DIFF[760]) );
  XOR U536 ( .A(B[760]), .B(A[760]), .Z(n536) );
  XOR U537 ( .A(n537), .B(n538), .Z(DIFF[75]) );
  XOR U538 ( .A(B[75]), .B(A[75]), .Z(n538) );
  XOR U539 ( .A(n539), .B(n540), .Z(DIFF[759]) );
  XOR U540 ( .A(B[759]), .B(A[759]), .Z(n540) );
  XOR U541 ( .A(n541), .B(n542), .Z(DIFF[758]) );
  XOR U542 ( .A(B[758]), .B(A[758]), .Z(n542) );
  XOR U543 ( .A(n543), .B(n544), .Z(DIFF[757]) );
  XOR U544 ( .A(B[757]), .B(A[757]), .Z(n544) );
  XOR U545 ( .A(n545), .B(n546), .Z(DIFF[756]) );
  XOR U546 ( .A(B[756]), .B(A[756]), .Z(n546) );
  XOR U547 ( .A(n547), .B(n548), .Z(DIFF[755]) );
  XOR U548 ( .A(B[755]), .B(A[755]), .Z(n548) );
  XOR U549 ( .A(n549), .B(n550), .Z(DIFF[754]) );
  XOR U550 ( .A(B[754]), .B(A[754]), .Z(n550) );
  XOR U551 ( .A(n551), .B(n552), .Z(DIFF[753]) );
  XOR U552 ( .A(B[753]), .B(A[753]), .Z(n552) );
  XOR U553 ( .A(n553), .B(n554), .Z(DIFF[752]) );
  XOR U554 ( .A(B[752]), .B(A[752]), .Z(n554) );
  XOR U555 ( .A(n555), .B(n556), .Z(DIFF[751]) );
  XOR U556 ( .A(B[751]), .B(A[751]), .Z(n556) );
  XOR U557 ( .A(n557), .B(n558), .Z(DIFF[750]) );
  XOR U558 ( .A(B[750]), .B(A[750]), .Z(n558) );
  XOR U559 ( .A(n559), .B(n560), .Z(DIFF[74]) );
  XOR U560 ( .A(B[74]), .B(A[74]), .Z(n560) );
  XOR U561 ( .A(n561), .B(n562), .Z(DIFF[749]) );
  XOR U562 ( .A(B[749]), .B(A[749]), .Z(n562) );
  XOR U563 ( .A(n563), .B(n564), .Z(DIFF[748]) );
  XOR U564 ( .A(B[748]), .B(A[748]), .Z(n564) );
  XOR U565 ( .A(n565), .B(n566), .Z(DIFF[747]) );
  XOR U566 ( .A(B[747]), .B(A[747]), .Z(n566) );
  XOR U567 ( .A(n567), .B(n568), .Z(DIFF[746]) );
  XOR U568 ( .A(B[746]), .B(A[746]), .Z(n568) );
  XOR U569 ( .A(n569), .B(n570), .Z(DIFF[745]) );
  XOR U570 ( .A(B[745]), .B(A[745]), .Z(n570) );
  XOR U571 ( .A(n571), .B(n572), .Z(DIFF[744]) );
  XOR U572 ( .A(B[744]), .B(A[744]), .Z(n572) );
  XOR U573 ( .A(n573), .B(n574), .Z(DIFF[743]) );
  XOR U574 ( .A(B[743]), .B(A[743]), .Z(n574) );
  XOR U575 ( .A(n575), .B(n576), .Z(DIFF[742]) );
  XOR U576 ( .A(B[742]), .B(A[742]), .Z(n576) );
  XOR U577 ( .A(n577), .B(n578), .Z(DIFF[741]) );
  XOR U578 ( .A(B[741]), .B(A[741]), .Z(n578) );
  XOR U579 ( .A(n579), .B(n580), .Z(DIFF[740]) );
  XOR U580 ( .A(B[740]), .B(A[740]), .Z(n580) );
  XOR U581 ( .A(n581), .B(n582), .Z(DIFF[73]) );
  XOR U582 ( .A(B[73]), .B(A[73]), .Z(n582) );
  XOR U583 ( .A(n583), .B(n584), .Z(DIFF[739]) );
  XOR U584 ( .A(B[739]), .B(A[739]), .Z(n584) );
  XOR U585 ( .A(n585), .B(n586), .Z(DIFF[738]) );
  XOR U586 ( .A(B[738]), .B(A[738]), .Z(n586) );
  XOR U587 ( .A(n587), .B(n588), .Z(DIFF[737]) );
  XOR U588 ( .A(B[737]), .B(A[737]), .Z(n588) );
  XOR U589 ( .A(n589), .B(n590), .Z(DIFF[736]) );
  XOR U590 ( .A(B[736]), .B(A[736]), .Z(n590) );
  XOR U591 ( .A(n591), .B(n592), .Z(DIFF[735]) );
  XOR U592 ( .A(B[735]), .B(A[735]), .Z(n592) );
  XOR U593 ( .A(n593), .B(n594), .Z(DIFF[734]) );
  XOR U594 ( .A(B[734]), .B(A[734]), .Z(n594) );
  XOR U595 ( .A(n595), .B(n596), .Z(DIFF[733]) );
  XOR U596 ( .A(B[733]), .B(A[733]), .Z(n596) );
  XOR U597 ( .A(n597), .B(n598), .Z(DIFF[732]) );
  XOR U598 ( .A(B[732]), .B(A[732]), .Z(n598) );
  XOR U599 ( .A(n599), .B(n600), .Z(DIFF[731]) );
  XOR U600 ( .A(B[731]), .B(A[731]), .Z(n600) );
  XOR U601 ( .A(n601), .B(n602), .Z(DIFF[730]) );
  XOR U602 ( .A(B[730]), .B(A[730]), .Z(n602) );
  XOR U603 ( .A(n603), .B(n604), .Z(DIFF[72]) );
  XOR U604 ( .A(B[72]), .B(A[72]), .Z(n604) );
  XOR U605 ( .A(n605), .B(n606), .Z(DIFF[729]) );
  XOR U606 ( .A(B[729]), .B(A[729]), .Z(n606) );
  XOR U607 ( .A(n607), .B(n608), .Z(DIFF[728]) );
  XOR U608 ( .A(B[728]), .B(A[728]), .Z(n608) );
  XOR U609 ( .A(n609), .B(n610), .Z(DIFF[727]) );
  XOR U610 ( .A(B[727]), .B(A[727]), .Z(n610) );
  XOR U611 ( .A(n611), .B(n612), .Z(DIFF[726]) );
  XOR U612 ( .A(B[726]), .B(A[726]), .Z(n612) );
  XOR U613 ( .A(n613), .B(n614), .Z(DIFF[725]) );
  XOR U614 ( .A(B[725]), .B(A[725]), .Z(n614) );
  XOR U615 ( .A(n615), .B(n616), .Z(DIFF[724]) );
  XOR U616 ( .A(B[724]), .B(A[724]), .Z(n616) );
  XOR U617 ( .A(n617), .B(n618), .Z(DIFF[723]) );
  XOR U618 ( .A(B[723]), .B(A[723]), .Z(n618) );
  XOR U619 ( .A(n619), .B(n620), .Z(DIFF[722]) );
  XOR U620 ( .A(B[722]), .B(A[722]), .Z(n620) );
  XOR U621 ( .A(n621), .B(n622), .Z(DIFF[721]) );
  XOR U622 ( .A(B[721]), .B(A[721]), .Z(n622) );
  XOR U623 ( .A(n623), .B(n624), .Z(DIFF[720]) );
  XOR U624 ( .A(B[720]), .B(A[720]), .Z(n624) );
  XOR U625 ( .A(n625), .B(n626), .Z(DIFF[71]) );
  XOR U626 ( .A(B[71]), .B(A[71]), .Z(n626) );
  XOR U627 ( .A(n627), .B(n628), .Z(DIFF[719]) );
  XOR U628 ( .A(B[719]), .B(A[719]), .Z(n628) );
  XOR U629 ( .A(n629), .B(n630), .Z(DIFF[718]) );
  XOR U630 ( .A(B[718]), .B(A[718]), .Z(n630) );
  XOR U631 ( .A(n631), .B(n632), .Z(DIFF[717]) );
  XOR U632 ( .A(B[717]), .B(A[717]), .Z(n632) );
  XOR U633 ( .A(n633), .B(n634), .Z(DIFF[716]) );
  XOR U634 ( .A(B[716]), .B(A[716]), .Z(n634) );
  XOR U635 ( .A(n635), .B(n636), .Z(DIFF[715]) );
  XOR U636 ( .A(B[715]), .B(A[715]), .Z(n636) );
  XOR U637 ( .A(n637), .B(n638), .Z(DIFF[714]) );
  XOR U638 ( .A(B[714]), .B(A[714]), .Z(n638) );
  XOR U639 ( .A(n639), .B(n640), .Z(DIFF[713]) );
  XOR U640 ( .A(B[713]), .B(A[713]), .Z(n640) );
  XOR U641 ( .A(n641), .B(n642), .Z(DIFF[712]) );
  XOR U642 ( .A(B[712]), .B(A[712]), .Z(n642) );
  XOR U643 ( .A(n643), .B(n644), .Z(DIFF[711]) );
  XOR U644 ( .A(B[711]), .B(A[711]), .Z(n644) );
  XOR U645 ( .A(n645), .B(n646), .Z(DIFF[710]) );
  XOR U646 ( .A(B[710]), .B(A[710]), .Z(n646) );
  XOR U647 ( .A(n647), .B(n648), .Z(DIFF[70]) );
  XOR U648 ( .A(B[70]), .B(A[70]), .Z(n648) );
  XOR U649 ( .A(n649), .B(n650), .Z(DIFF[709]) );
  XOR U650 ( .A(B[709]), .B(A[709]), .Z(n650) );
  XOR U651 ( .A(n651), .B(n652), .Z(DIFF[708]) );
  XOR U652 ( .A(B[708]), .B(A[708]), .Z(n652) );
  XOR U653 ( .A(n653), .B(n654), .Z(DIFF[707]) );
  XOR U654 ( .A(B[707]), .B(A[707]), .Z(n654) );
  XOR U655 ( .A(n655), .B(n656), .Z(DIFF[706]) );
  XOR U656 ( .A(B[706]), .B(A[706]), .Z(n656) );
  XOR U657 ( .A(n657), .B(n658), .Z(DIFF[705]) );
  XOR U658 ( .A(B[705]), .B(A[705]), .Z(n658) );
  XOR U659 ( .A(n659), .B(n660), .Z(DIFF[704]) );
  XOR U660 ( .A(B[704]), .B(A[704]), .Z(n660) );
  XOR U661 ( .A(n661), .B(n662), .Z(DIFF[703]) );
  XOR U662 ( .A(B[703]), .B(A[703]), .Z(n662) );
  XOR U663 ( .A(n663), .B(n664), .Z(DIFF[702]) );
  XOR U664 ( .A(B[702]), .B(A[702]), .Z(n664) );
  XOR U665 ( .A(n665), .B(n666), .Z(DIFF[701]) );
  XOR U666 ( .A(B[701]), .B(A[701]), .Z(n666) );
  XOR U667 ( .A(n667), .B(n668), .Z(DIFF[700]) );
  XOR U668 ( .A(B[700]), .B(A[700]), .Z(n668) );
  XOR U669 ( .A(n669), .B(n670), .Z(DIFF[6]) );
  XOR U670 ( .A(B[6]), .B(A[6]), .Z(n670) );
  XOR U671 ( .A(n671), .B(n672), .Z(DIFF[69]) );
  XOR U672 ( .A(B[69]), .B(A[69]), .Z(n672) );
  XOR U673 ( .A(n673), .B(n674), .Z(DIFF[699]) );
  XOR U674 ( .A(B[699]), .B(A[699]), .Z(n674) );
  XOR U675 ( .A(n675), .B(n676), .Z(DIFF[698]) );
  XOR U676 ( .A(B[698]), .B(A[698]), .Z(n676) );
  XOR U677 ( .A(n677), .B(n678), .Z(DIFF[697]) );
  XOR U678 ( .A(B[697]), .B(A[697]), .Z(n678) );
  XOR U679 ( .A(n679), .B(n680), .Z(DIFF[696]) );
  XOR U680 ( .A(B[696]), .B(A[696]), .Z(n680) );
  XOR U681 ( .A(n681), .B(n682), .Z(DIFF[695]) );
  XOR U682 ( .A(B[695]), .B(A[695]), .Z(n682) );
  XOR U683 ( .A(n683), .B(n684), .Z(DIFF[694]) );
  XOR U684 ( .A(B[694]), .B(A[694]), .Z(n684) );
  XOR U685 ( .A(n685), .B(n686), .Z(DIFF[693]) );
  XOR U686 ( .A(B[693]), .B(A[693]), .Z(n686) );
  XOR U687 ( .A(n687), .B(n688), .Z(DIFF[692]) );
  XOR U688 ( .A(B[692]), .B(A[692]), .Z(n688) );
  XOR U689 ( .A(n689), .B(n690), .Z(DIFF[691]) );
  XOR U690 ( .A(B[691]), .B(A[691]), .Z(n690) );
  XOR U691 ( .A(n691), .B(n692), .Z(DIFF[690]) );
  XOR U692 ( .A(B[690]), .B(A[690]), .Z(n692) );
  XOR U693 ( .A(n693), .B(n694), .Z(DIFF[68]) );
  XOR U694 ( .A(B[68]), .B(A[68]), .Z(n694) );
  XOR U695 ( .A(n695), .B(n696), .Z(DIFF[689]) );
  XOR U696 ( .A(B[689]), .B(A[689]), .Z(n696) );
  XOR U697 ( .A(n697), .B(n698), .Z(DIFF[688]) );
  XOR U698 ( .A(B[688]), .B(A[688]), .Z(n698) );
  XOR U699 ( .A(n699), .B(n700), .Z(DIFF[687]) );
  XOR U700 ( .A(B[687]), .B(A[687]), .Z(n700) );
  XOR U701 ( .A(n701), .B(n702), .Z(DIFF[686]) );
  XOR U702 ( .A(B[686]), .B(A[686]), .Z(n702) );
  XOR U703 ( .A(n703), .B(n704), .Z(DIFF[685]) );
  XOR U704 ( .A(B[685]), .B(A[685]), .Z(n704) );
  XOR U705 ( .A(n705), .B(n706), .Z(DIFF[684]) );
  XOR U706 ( .A(B[684]), .B(A[684]), .Z(n706) );
  XOR U707 ( .A(n707), .B(n708), .Z(DIFF[683]) );
  XOR U708 ( .A(B[683]), .B(A[683]), .Z(n708) );
  XOR U709 ( .A(n709), .B(n710), .Z(DIFF[682]) );
  XOR U710 ( .A(B[682]), .B(A[682]), .Z(n710) );
  XOR U711 ( .A(n711), .B(n712), .Z(DIFF[681]) );
  XOR U712 ( .A(B[681]), .B(A[681]), .Z(n712) );
  XOR U713 ( .A(n713), .B(n714), .Z(DIFF[680]) );
  XOR U714 ( .A(B[680]), .B(A[680]), .Z(n714) );
  XOR U715 ( .A(n715), .B(n716), .Z(DIFF[67]) );
  XOR U716 ( .A(B[67]), .B(A[67]), .Z(n716) );
  XOR U717 ( .A(n717), .B(n718), .Z(DIFF[679]) );
  XOR U718 ( .A(B[679]), .B(A[679]), .Z(n718) );
  XOR U719 ( .A(n719), .B(n720), .Z(DIFF[678]) );
  XOR U720 ( .A(B[678]), .B(A[678]), .Z(n720) );
  XOR U721 ( .A(n721), .B(n722), .Z(DIFF[677]) );
  XOR U722 ( .A(B[677]), .B(A[677]), .Z(n722) );
  XOR U723 ( .A(n723), .B(n724), .Z(DIFF[676]) );
  XOR U724 ( .A(B[676]), .B(A[676]), .Z(n724) );
  XOR U725 ( .A(n725), .B(n726), .Z(DIFF[675]) );
  XOR U726 ( .A(B[675]), .B(A[675]), .Z(n726) );
  XOR U727 ( .A(n727), .B(n728), .Z(DIFF[674]) );
  XOR U728 ( .A(B[674]), .B(A[674]), .Z(n728) );
  XOR U729 ( .A(n729), .B(n730), .Z(DIFF[673]) );
  XOR U730 ( .A(B[673]), .B(A[673]), .Z(n730) );
  XOR U731 ( .A(n731), .B(n732), .Z(DIFF[672]) );
  XOR U732 ( .A(B[672]), .B(A[672]), .Z(n732) );
  XOR U733 ( .A(n733), .B(n734), .Z(DIFF[671]) );
  XOR U734 ( .A(B[671]), .B(A[671]), .Z(n734) );
  XOR U735 ( .A(n735), .B(n736), .Z(DIFF[670]) );
  XOR U736 ( .A(B[670]), .B(A[670]), .Z(n736) );
  XOR U737 ( .A(n737), .B(n738), .Z(DIFF[66]) );
  XOR U738 ( .A(B[66]), .B(A[66]), .Z(n738) );
  XOR U739 ( .A(n739), .B(n740), .Z(DIFF[669]) );
  XOR U740 ( .A(B[669]), .B(A[669]), .Z(n740) );
  XOR U741 ( .A(n741), .B(n742), .Z(DIFF[668]) );
  XOR U742 ( .A(B[668]), .B(A[668]), .Z(n742) );
  XOR U743 ( .A(n743), .B(n744), .Z(DIFF[667]) );
  XOR U744 ( .A(B[667]), .B(A[667]), .Z(n744) );
  XOR U745 ( .A(n745), .B(n746), .Z(DIFF[666]) );
  XOR U746 ( .A(B[666]), .B(A[666]), .Z(n746) );
  XOR U747 ( .A(n747), .B(n748), .Z(DIFF[665]) );
  XOR U748 ( .A(B[665]), .B(A[665]), .Z(n748) );
  XOR U749 ( .A(n749), .B(n750), .Z(DIFF[664]) );
  XOR U750 ( .A(B[664]), .B(A[664]), .Z(n750) );
  XOR U751 ( .A(n751), .B(n752), .Z(DIFF[663]) );
  XOR U752 ( .A(B[663]), .B(A[663]), .Z(n752) );
  XOR U753 ( .A(n753), .B(n754), .Z(DIFF[662]) );
  XOR U754 ( .A(B[662]), .B(A[662]), .Z(n754) );
  XOR U755 ( .A(n755), .B(n756), .Z(DIFF[661]) );
  XOR U756 ( .A(B[661]), .B(A[661]), .Z(n756) );
  XOR U757 ( .A(n757), .B(n758), .Z(DIFF[660]) );
  XOR U758 ( .A(B[660]), .B(A[660]), .Z(n758) );
  XOR U759 ( .A(n759), .B(n760), .Z(DIFF[65]) );
  XOR U760 ( .A(B[65]), .B(A[65]), .Z(n760) );
  XOR U761 ( .A(n761), .B(n762), .Z(DIFF[659]) );
  XOR U762 ( .A(B[659]), .B(A[659]), .Z(n762) );
  XOR U763 ( .A(n763), .B(n764), .Z(DIFF[658]) );
  XOR U764 ( .A(B[658]), .B(A[658]), .Z(n764) );
  XOR U765 ( .A(n765), .B(n766), .Z(DIFF[657]) );
  XOR U766 ( .A(B[657]), .B(A[657]), .Z(n766) );
  XOR U767 ( .A(n767), .B(n768), .Z(DIFF[656]) );
  XOR U768 ( .A(B[656]), .B(A[656]), .Z(n768) );
  XOR U769 ( .A(n769), .B(n770), .Z(DIFF[655]) );
  XOR U770 ( .A(B[655]), .B(A[655]), .Z(n770) );
  XOR U771 ( .A(n771), .B(n772), .Z(DIFF[654]) );
  XOR U772 ( .A(B[654]), .B(A[654]), .Z(n772) );
  XOR U773 ( .A(n773), .B(n774), .Z(DIFF[653]) );
  XOR U774 ( .A(B[653]), .B(A[653]), .Z(n774) );
  XOR U775 ( .A(n775), .B(n776), .Z(DIFF[652]) );
  XOR U776 ( .A(B[652]), .B(A[652]), .Z(n776) );
  XOR U777 ( .A(n777), .B(n778), .Z(DIFF[651]) );
  XOR U778 ( .A(B[651]), .B(A[651]), .Z(n778) );
  XOR U779 ( .A(n779), .B(n780), .Z(DIFF[650]) );
  XOR U780 ( .A(B[650]), .B(A[650]), .Z(n780) );
  XOR U781 ( .A(n781), .B(n782), .Z(DIFF[64]) );
  XOR U782 ( .A(B[64]), .B(A[64]), .Z(n782) );
  XOR U783 ( .A(n783), .B(n784), .Z(DIFF[649]) );
  XOR U784 ( .A(B[649]), .B(A[649]), .Z(n784) );
  XOR U785 ( .A(n785), .B(n786), .Z(DIFF[648]) );
  XOR U786 ( .A(B[648]), .B(A[648]), .Z(n786) );
  XOR U787 ( .A(n787), .B(n788), .Z(DIFF[647]) );
  XOR U788 ( .A(B[647]), .B(A[647]), .Z(n788) );
  XOR U789 ( .A(n789), .B(n790), .Z(DIFF[646]) );
  XOR U790 ( .A(B[646]), .B(A[646]), .Z(n790) );
  XOR U791 ( .A(n791), .B(n792), .Z(DIFF[645]) );
  XOR U792 ( .A(B[645]), .B(A[645]), .Z(n792) );
  XOR U793 ( .A(n793), .B(n794), .Z(DIFF[644]) );
  XOR U794 ( .A(B[644]), .B(A[644]), .Z(n794) );
  XOR U795 ( .A(n795), .B(n796), .Z(DIFF[643]) );
  XOR U796 ( .A(B[643]), .B(A[643]), .Z(n796) );
  XOR U797 ( .A(n797), .B(n798), .Z(DIFF[642]) );
  XOR U798 ( .A(B[642]), .B(A[642]), .Z(n798) );
  XOR U799 ( .A(n799), .B(n800), .Z(DIFF[641]) );
  XOR U800 ( .A(B[641]), .B(A[641]), .Z(n800) );
  XOR U801 ( .A(n801), .B(n802), .Z(DIFF[640]) );
  XOR U802 ( .A(B[640]), .B(A[640]), .Z(n802) );
  XOR U803 ( .A(n803), .B(n804), .Z(DIFF[63]) );
  XOR U804 ( .A(B[63]), .B(A[63]), .Z(n804) );
  XOR U805 ( .A(n805), .B(n806), .Z(DIFF[639]) );
  XOR U806 ( .A(B[639]), .B(A[639]), .Z(n806) );
  XOR U807 ( .A(n807), .B(n808), .Z(DIFF[638]) );
  XOR U808 ( .A(B[638]), .B(A[638]), .Z(n808) );
  XOR U809 ( .A(n809), .B(n810), .Z(DIFF[637]) );
  XOR U810 ( .A(B[637]), .B(A[637]), .Z(n810) );
  XOR U811 ( .A(n811), .B(n812), .Z(DIFF[636]) );
  XOR U812 ( .A(B[636]), .B(A[636]), .Z(n812) );
  XOR U813 ( .A(n813), .B(n814), .Z(DIFF[635]) );
  XOR U814 ( .A(B[635]), .B(A[635]), .Z(n814) );
  XOR U815 ( .A(n815), .B(n816), .Z(DIFF[634]) );
  XOR U816 ( .A(B[634]), .B(A[634]), .Z(n816) );
  XOR U817 ( .A(n817), .B(n818), .Z(DIFF[633]) );
  XOR U818 ( .A(B[633]), .B(A[633]), .Z(n818) );
  XOR U819 ( .A(n819), .B(n820), .Z(DIFF[632]) );
  XOR U820 ( .A(B[632]), .B(A[632]), .Z(n820) );
  XOR U821 ( .A(n821), .B(n822), .Z(DIFF[631]) );
  XOR U822 ( .A(B[631]), .B(A[631]), .Z(n822) );
  XOR U823 ( .A(n823), .B(n824), .Z(DIFF[630]) );
  XOR U824 ( .A(B[630]), .B(A[630]), .Z(n824) );
  XOR U825 ( .A(n825), .B(n826), .Z(DIFF[62]) );
  XOR U826 ( .A(B[62]), .B(A[62]), .Z(n826) );
  XOR U827 ( .A(n827), .B(n828), .Z(DIFF[629]) );
  XOR U828 ( .A(B[629]), .B(A[629]), .Z(n828) );
  XOR U829 ( .A(n829), .B(n830), .Z(DIFF[628]) );
  XOR U830 ( .A(B[628]), .B(A[628]), .Z(n830) );
  XOR U831 ( .A(n831), .B(n832), .Z(DIFF[627]) );
  XOR U832 ( .A(B[627]), .B(A[627]), .Z(n832) );
  XOR U833 ( .A(n833), .B(n834), .Z(DIFF[626]) );
  XOR U834 ( .A(B[626]), .B(A[626]), .Z(n834) );
  XOR U835 ( .A(n835), .B(n836), .Z(DIFF[625]) );
  XOR U836 ( .A(B[625]), .B(A[625]), .Z(n836) );
  XOR U837 ( .A(n837), .B(n838), .Z(DIFF[624]) );
  XOR U838 ( .A(B[624]), .B(A[624]), .Z(n838) );
  XOR U839 ( .A(n839), .B(n840), .Z(DIFF[623]) );
  XOR U840 ( .A(B[623]), .B(A[623]), .Z(n840) );
  XOR U841 ( .A(n841), .B(n842), .Z(DIFF[622]) );
  XOR U842 ( .A(B[622]), .B(A[622]), .Z(n842) );
  XOR U843 ( .A(n843), .B(n844), .Z(DIFF[621]) );
  XOR U844 ( .A(B[621]), .B(A[621]), .Z(n844) );
  XOR U845 ( .A(n845), .B(n846), .Z(DIFF[620]) );
  XOR U846 ( .A(B[620]), .B(A[620]), .Z(n846) );
  XOR U847 ( .A(n847), .B(n848), .Z(DIFF[61]) );
  XOR U848 ( .A(B[61]), .B(A[61]), .Z(n848) );
  XOR U849 ( .A(n849), .B(n850), .Z(DIFF[619]) );
  XOR U850 ( .A(B[619]), .B(A[619]), .Z(n850) );
  XOR U851 ( .A(n851), .B(n852), .Z(DIFF[618]) );
  XOR U852 ( .A(B[618]), .B(A[618]), .Z(n852) );
  XOR U853 ( .A(n853), .B(n854), .Z(DIFF[617]) );
  XOR U854 ( .A(B[617]), .B(A[617]), .Z(n854) );
  XOR U855 ( .A(n855), .B(n856), .Z(DIFF[616]) );
  XOR U856 ( .A(B[616]), .B(A[616]), .Z(n856) );
  XOR U857 ( .A(n857), .B(n858), .Z(DIFF[615]) );
  XOR U858 ( .A(B[615]), .B(A[615]), .Z(n858) );
  XOR U859 ( .A(n859), .B(n860), .Z(DIFF[614]) );
  XOR U860 ( .A(B[614]), .B(A[614]), .Z(n860) );
  XOR U861 ( .A(n861), .B(n862), .Z(DIFF[613]) );
  XOR U862 ( .A(B[613]), .B(A[613]), .Z(n862) );
  XOR U863 ( .A(n863), .B(n864), .Z(DIFF[612]) );
  XOR U864 ( .A(B[612]), .B(A[612]), .Z(n864) );
  XOR U865 ( .A(n865), .B(n866), .Z(DIFF[611]) );
  XOR U866 ( .A(B[611]), .B(A[611]), .Z(n866) );
  XOR U867 ( .A(n867), .B(n868), .Z(DIFF[610]) );
  XOR U868 ( .A(B[610]), .B(A[610]), .Z(n868) );
  XOR U869 ( .A(n869), .B(n870), .Z(DIFF[60]) );
  XOR U870 ( .A(B[60]), .B(A[60]), .Z(n870) );
  XOR U871 ( .A(n871), .B(n872), .Z(DIFF[609]) );
  XOR U872 ( .A(B[609]), .B(A[609]), .Z(n872) );
  XOR U873 ( .A(n873), .B(n874), .Z(DIFF[608]) );
  XOR U874 ( .A(B[608]), .B(A[608]), .Z(n874) );
  XOR U875 ( .A(n875), .B(n876), .Z(DIFF[607]) );
  XOR U876 ( .A(B[607]), .B(A[607]), .Z(n876) );
  XOR U877 ( .A(n877), .B(n878), .Z(DIFF[606]) );
  XOR U878 ( .A(B[606]), .B(A[606]), .Z(n878) );
  XOR U879 ( .A(n879), .B(n880), .Z(DIFF[605]) );
  XOR U880 ( .A(B[605]), .B(A[605]), .Z(n880) );
  XOR U881 ( .A(n881), .B(n882), .Z(DIFF[604]) );
  XOR U882 ( .A(B[604]), .B(A[604]), .Z(n882) );
  XOR U883 ( .A(n883), .B(n884), .Z(DIFF[603]) );
  XOR U884 ( .A(B[603]), .B(A[603]), .Z(n884) );
  XOR U885 ( .A(n885), .B(n886), .Z(DIFF[602]) );
  XOR U886 ( .A(B[602]), .B(A[602]), .Z(n886) );
  XOR U887 ( .A(n887), .B(n888), .Z(DIFF[601]) );
  XOR U888 ( .A(B[601]), .B(A[601]), .Z(n888) );
  XOR U889 ( .A(n889), .B(n890), .Z(DIFF[600]) );
  XOR U890 ( .A(B[600]), .B(A[600]), .Z(n890) );
  XOR U891 ( .A(n891), .B(n892), .Z(DIFF[5]) );
  XOR U892 ( .A(B[5]), .B(A[5]), .Z(n892) );
  XOR U893 ( .A(n893), .B(n894), .Z(DIFF[59]) );
  XOR U894 ( .A(B[59]), .B(A[59]), .Z(n894) );
  XOR U895 ( .A(n895), .B(n896), .Z(DIFF[599]) );
  XOR U896 ( .A(B[599]), .B(A[599]), .Z(n896) );
  XOR U897 ( .A(n897), .B(n898), .Z(DIFF[598]) );
  XOR U898 ( .A(B[598]), .B(A[598]), .Z(n898) );
  XOR U899 ( .A(n899), .B(n900), .Z(DIFF[597]) );
  XOR U900 ( .A(B[597]), .B(A[597]), .Z(n900) );
  XOR U901 ( .A(n901), .B(n902), .Z(DIFF[596]) );
  XOR U902 ( .A(B[596]), .B(A[596]), .Z(n902) );
  XOR U903 ( .A(n903), .B(n904), .Z(DIFF[595]) );
  XOR U904 ( .A(B[595]), .B(A[595]), .Z(n904) );
  XOR U905 ( .A(n905), .B(n906), .Z(DIFF[594]) );
  XOR U906 ( .A(B[594]), .B(A[594]), .Z(n906) );
  XOR U907 ( .A(n907), .B(n908), .Z(DIFF[593]) );
  XOR U908 ( .A(B[593]), .B(A[593]), .Z(n908) );
  XOR U909 ( .A(n909), .B(n910), .Z(DIFF[592]) );
  XOR U910 ( .A(B[592]), .B(A[592]), .Z(n910) );
  XOR U911 ( .A(n911), .B(n912), .Z(DIFF[591]) );
  XOR U912 ( .A(B[591]), .B(A[591]), .Z(n912) );
  XOR U913 ( .A(n913), .B(n914), .Z(DIFF[590]) );
  XOR U914 ( .A(B[590]), .B(A[590]), .Z(n914) );
  XOR U915 ( .A(n915), .B(n916), .Z(DIFF[58]) );
  XOR U916 ( .A(B[58]), .B(A[58]), .Z(n916) );
  XOR U917 ( .A(n917), .B(n918), .Z(DIFF[589]) );
  XOR U918 ( .A(B[589]), .B(A[589]), .Z(n918) );
  XOR U919 ( .A(n919), .B(n920), .Z(DIFF[588]) );
  XOR U920 ( .A(B[588]), .B(A[588]), .Z(n920) );
  XOR U921 ( .A(n921), .B(n922), .Z(DIFF[587]) );
  XOR U922 ( .A(B[587]), .B(A[587]), .Z(n922) );
  XOR U923 ( .A(n923), .B(n924), .Z(DIFF[586]) );
  XOR U924 ( .A(B[586]), .B(A[586]), .Z(n924) );
  XOR U925 ( .A(n925), .B(n926), .Z(DIFF[585]) );
  XOR U926 ( .A(B[585]), .B(A[585]), .Z(n926) );
  XOR U927 ( .A(n927), .B(n928), .Z(DIFF[584]) );
  XOR U928 ( .A(B[584]), .B(A[584]), .Z(n928) );
  XOR U929 ( .A(n929), .B(n930), .Z(DIFF[583]) );
  XOR U930 ( .A(B[583]), .B(A[583]), .Z(n930) );
  XOR U931 ( .A(n931), .B(n932), .Z(DIFF[582]) );
  XOR U932 ( .A(B[582]), .B(A[582]), .Z(n932) );
  XOR U933 ( .A(n933), .B(n934), .Z(DIFF[581]) );
  XOR U934 ( .A(B[581]), .B(A[581]), .Z(n934) );
  XOR U935 ( .A(n935), .B(n936), .Z(DIFF[580]) );
  XOR U936 ( .A(B[580]), .B(A[580]), .Z(n936) );
  XOR U937 ( .A(n937), .B(n938), .Z(DIFF[57]) );
  XOR U938 ( .A(B[57]), .B(A[57]), .Z(n938) );
  XOR U939 ( .A(n939), .B(n940), .Z(DIFF[579]) );
  XOR U940 ( .A(B[579]), .B(A[579]), .Z(n940) );
  XOR U941 ( .A(n941), .B(n942), .Z(DIFF[578]) );
  XOR U942 ( .A(B[578]), .B(A[578]), .Z(n942) );
  XOR U943 ( .A(n943), .B(n944), .Z(DIFF[577]) );
  XOR U944 ( .A(B[577]), .B(A[577]), .Z(n944) );
  XOR U945 ( .A(n945), .B(n946), .Z(DIFF[576]) );
  XOR U946 ( .A(B[576]), .B(A[576]), .Z(n946) );
  XOR U947 ( .A(n947), .B(n948), .Z(DIFF[575]) );
  XOR U948 ( .A(B[575]), .B(A[575]), .Z(n948) );
  XOR U949 ( .A(n949), .B(n950), .Z(DIFF[574]) );
  XOR U950 ( .A(B[574]), .B(A[574]), .Z(n950) );
  XOR U951 ( .A(n951), .B(n952), .Z(DIFF[573]) );
  XOR U952 ( .A(B[573]), .B(A[573]), .Z(n952) );
  XOR U953 ( .A(n953), .B(n954), .Z(DIFF[572]) );
  XOR U954 ( .A(B[572]), .B(A[572]), .Z(n954) );
  XOR U955 ( .A(n955), .B(n956), .Z(DIFF[571]) );
  XOR U956 ( .A(B[571]), .B(A[571]), .Z(n956) );
  XOR U957 ( .A(n957), .B(n958), .Z(DIFF[570]) );
  XOR U958 ( .A(B[570]), .B(A[570]), .Z(n958) );
  XOR U959 ( .A(n959), .B(n960), .Z(DIFF[56]) );
  XOR U960 ( .A(B[56]), .B(A[56]), .Z(n960) );
  XOR U961 ( .A(n961), .B(n962), .Z(DIFF[569]) );
  XOR U962 ( .A(B[569]), .B(A[569]), .Z(n962) );
  XOR U963 ( .A(n963), .B(n964), .Z(DIFF[568]) );
  XOR U964 ( .A(B[568]), .B(A[568]), .Z(n964) );
  XOR U965 ( .A(n965), .B(n966), .Z(DIFF[567]) );
  XOR U966 ( .A(B[567]), .B(A[567]), .Z(n966) );
  XOR U967 ( .A(n967), .B(n968), .Z(DIFF[566]) );
  XOR U968 ( .A(B[566]), .B(A[566]), .Z(n968) );
  XOR U969 ( .A(n969), .B(n970), .Z(DIFF[565]) );
  XOR U970 ( .A(B[565]), .B(A[565]), .Z(n970) );
  XOR U971 ( .A(n971), .B(n972), .Z(DIFF[564]) );
  XOR U972 ( .A(B[564]), .B(A[564]), .Z(n972) );
  XOR U973 ( .A(n973), .B(n974), .Z(DIFF[563]) );
  XOR U974 ( .A(B[563]), .B(A[563]), .Z(n974) );
  XOR U975 ( .A(n975), .B(n976), .Z(DIFF[562]) );
  XOR U976 ( .A(B[562]), .B(A[562]), .Z(n976) );
  XOR U977 ( .A(n977), .B(n978), .Z(DIFF[561]) );
  XOR U978 ( .A(B[561]), .B(A[561]), .Z(n978) );
  XOR U979 ( .A(n979), .B(n980), .Z(DIFF[560]) );
  XOR U980 ( .A(B[560]), .B(A[560]), .Z(n980) );
  XOR U981 ( .A(n981), .B(n982), .Z(DIFF[55]) );
  XOR U982 ( .A(B[55]), .B(A[55]), .Z(n982) );
  XOR U983 ( .A(n983), .B(n984), .Z(DIFF[559]) );
  XOR U984 ( .A(B[559]), .B(A[559]), .Z(n984) );
  XOR U985 ( .A(n985), .B(n986), .Z(DIFF[558]) );
  XOR U986 ( .A(B[558]), .B(A[558]), .Z(n986) );
  XOR U987 ( .A(n987), .B(n988), .Z(DIFF[557]) );
  XOR U988 ( .A(B[557]), .B(A[557]), .Z(n988) );
  XOR U989 ( .A(n989), .B(n990), .Z(DIFF[556]) );
  XOR U990 ( .A(B[556]), .B(A[556]), .Z(n990) );
  XOR U991 ( .A(n991), .B(n992), .Z(DIFF[555]) );
  XOR U992 ( .A(B[555]), .B(A[555]), .Z(n992) );
  XOR U993 ( .A(n993), .B(n994), .Z(DIFF[554]) );
  XOR U994 ( .A(B[554]), .B(A[554]), .Z(n994) );
  XOR U995 ( .A(n995), .B(n996), .Z(DIFF[553]) );
  XOR U996 ( .A(B[553]), .B(A[553]), .Z(n996) );
  XOR U997 ( .A(n997), .B(n998), .Z(DIFF[552]) );
  XOR U998 ( .A(B[552]), .B(A[552]), .Z(n998) );
  XOR U999 ( .A(n999), .B(n1000), .Z(DIFF[551]) );
  XOR U1000 ( .A(B[551]), .B(A[551]), .Z(n1000) );
  XOR U1001 ( .A(n1001), .B(n1002), .Z(DIFF[550]) );
  XOR U1002 ( .A(B[550]), .B(A[550]), .Z(n1002) );
  XOR U1003 ( .A(n1003), .B(n1004), .Z(DIFF[54]) );
  XOR U1004 ( .A(B[54]), .B(A[54]), .Z(n1004) );
  XOR U1005 ( .A(n1005), .B(n1006), .Z(DIFF[549]) );
  XOR U1006 ( .A(B[549]), .B(A[549]), .Z(n1006) );
  XOR U1007 ( .A(n1007), .B(n1008), .Z(DIFF[548]) );
  XOR U1008 ( .A(B[548]), .B(A[548]), .Z(n1008) );
  XOR U1009 ( .A(n1009), .B(n1010), .Z(DIFF[547]) );
  XOR U1010 ( .A(B[547]), .B(A[547]), .Z(n1010) );
  XOR U1011 ( .A(n1011), .B(n1012), .Z(DIFF[546]) );
  XOR U1012 ( .A(B[546]), .B(A[546]), .Z(n1012) );
  XOR U1013 ( .A(n1013), .B(n1014), .Z(DIFF[545]) );
  XOR U1014 ( .A(B[545]), .B(A[545]), .Z(n1014) );
  XOR U1015 ( .A(n1015), .B(n1016), .Z(DIFF[544]) );
  XOR U1016 ( .A(B[544]), .B(A[544]), .Z(n1016) );
  XOR U1017 ( .A(n1017), .B(n1018), .Z(DIFF[543]) );
  XOR U1018 ( .A(B[543]), .B(A[543]), .Z(n1018) );
  XOR U1019 ( .A(n1019), .B(n1020), .Z(DIFF[542]) );
  XOR U1020 ( .A(B[542]), .B(A[542]), .Z(n1020) );
  XOR U1021 ( .A(n1021), .B(n1022), .Z(DIFF[541]) );
  XOR U1022 ( .A(B[541]), .B(A[541]), .Z(n1022) );
  XOR U1023 ( .A(n1023), .B(n1024), .Z(DIFF[540]) );
  XOR U1024 ( .A(B[540]), .B(A[540]), .Z(n1024) );
  XOR U1025 ( .A(n1025), .B(n1026), .Z(DIFF[53]) );
  XOR U1026 ( .A(B[53]), .B(A[53]), .Z(n1026) );
  XOR U1027 ( .A(n1027), .B(n1028), .Z(DIFF[539]) );
  XOR U1028 ( .A(B[539]), .B(A[539]), .Z(n1028) );
  XOR U1029 ( .A(n1029), .B(n1030), .Z(DIFF[538]) );
  XOR U1030 ( .A(B[538]), .B(A[538]), .Z(n1030) );
  XOR U1031 ( .A(n1031), .B(n1032), .Z(DIFF[537]) );
  XOR U1032 ( .A(B[537]), .B(A[537]), .Z(n1032) );
  XOR U1033 ( .A(n1033), .B(n1034), .Z(DIFF[536]) );
  XOR U1034 ( .A(B[536]), .B(A[536]), .Z(n1034) );
  XOR U1035 ( .A(n1035), .B(n1036), .Z(DIFF[535]) );
  XOR U1036 ( .A(B[535]), .B(A[535]), .Z(n1036) );
  XOR U1037 ( .A(n1037), .B(n1038), .Z(DIFF[534]) );
  XOR U1038 ( .A(B[534]), .B(A[534]), .Z(n1038) );
  XOR U1039 ( .A(n1039), .B(n1040), .Z(DIFF[533]) );
  XOR U1040 ( .A(B[533]), .B(A[533]), .Z(n1040) );
  XOR U1041 ( .A(n1041), .B(n1042), .Z(DIFF[532]) );
  XOR U1042 ( .A(B[532]), .B(A[532]), .Z(n1042) );
  XOR U1043 ( .A(n1043), .B(n1044), .Z(DIFF[531]) );
  XOR U1044 ( .A(B[531]), .B(A[531]), .Z(n1044) );
  XOR U1045 ( .A(n1045), .B(n1046), .Z(DIFF[530]) );
  XOR U1046 ( .A(B[530]), .B(A[530]), .Z(n1046) );
  XOR U1047 ( .A(n1047), .B(n1048), .Z(DIFF[52]) );
  XOR U1048 ( .A(B[52]), .B(A[52]), .Z(n1048) );
  XOR U1049 ( .A(n1049), .B(n1050), .Z(DIFF[529]) );
  XOR U1050 ( .A(B[529]), .B(A[529]), .Z(n1050) );
  XOR U1051 ( .A(n1051), .B(n1052), .Z(DIFF[528]) );
  XOR U1052 ( .A(B[528]), .B(A[528]), .Z(n1052) );
  XOR U1053 ( .A(n1053), .B(n1054), .Z(DIFF[527]) );
  XOR U1054 ( .A(B[527]), .B(A[527]), .Z(n1054) );
  XOR U1055 ( .A(n1055), .B(n1056), .Z(DIFF[526]) );
  XOR U1056 ( .A(B[526]), .B(A[526]), .Z(n1056) );
  XOR U1057 ( .A(n1057), .B(n1058), .Z(DIFF[525]) );
  XOR U1058 ( .A(B[525]), .B(A[525]), .Z(n1058) );
  XOR U1059 ( .A(n1059), .B(n1060), .Z(DIFF[524]) );
  XOR U1060 ( .A(B[524]), .B(A[524]), .Z(n1060) );
  XOR U1061 ( .A(n1061), .B(n1062), .Z(DIFF[523]) );
  XOR U1062 ( .A(B[523]), .B(A[523]), .Z(n1062) );
  XOR U1063 ( .A(n1063), .B(n1064), .Z(DIFF[522]) );
  XOR U1064 ( .A(B[522]), .B(A[522]), .Z(n1064) );
  XOR U1065 ( .A(n1065), .B(n1066), .Z(DIFF[521]) );
  XOR U1066 ( .A(B[521]), .B(A[521]), .Z(n1066) );
  XOR U1067 ( .A(n1067), .B(n1068), .Z(DIFF[520]) );
  XOR U1068 ( .A(B[520]), .B(A[520]), .Z(n1068) );
  XOR U1069 ( .A(n1069), .B(n1070), .Z(DIFF[51]) );
  XOR U1070 ( .A(B[51]), .B(A[51]), .Z(n1070) );
  XOR U1071 ( .A(n1071), .B(n1072), .Z(DIFF[519]) );
  XOR U1072 ( .A(B[519]), .B(A[519]), .Z(n1072) );
  XOR U1073 ( .A(n1073), .B(n1074), .Z(DIFF[518]) );
  XOR U1074 ( .A(B[518]), .B(A[518]), .Z(n1074) );
  XOR U1075 ( .A(n1075), .B(n1076), .Z(DIFF[517]) );
  XOR U1076 ( .A(B[517]), .B(A[517]), .Z(n1076) );
  XOR U1077 ( .A(n1077), .B(n1078), .Z(DIFF[516]) );
  XOR U1078 ( .A(B[516]), .B(A[516]), .Z(n1078) );
  XOR U1079 ( .A(n1079), .B(n1080), .Z(DIFF[515]) );
  XOR U1080 ( .A(B[515]), .B(A[515]), .Z(n1080) );
  XOR U1081 ( .A(n1081), .B(n1082), .Z(DIFF[514]) );
  XOR U1082 ( .A(B[514]), .B(A[514]), .Z(n1082) );
  XOR U1083 ( .A(n1083), .B(n1084), .Z(DIFF[513]) );
  XOR U1084 ( .A(B[513]), .B(A[513]), .Z(n1084) );
  XOR U1085 ( .A(n1085), .B(n1086), .Z(DIFF[512]) );
  XOR U1086 ( .A(B[512]), .B(A[512]), .Z(n1086) );
  XOR U1087 ( .A(n1087), .B(n1088), .Z(DIFF[511]) );
  XOR U1088 ( .A(B[511]), .B(A[511]), .Z(n1088) );
  XOR U1089 ( .A(n1089), .B(n1090), .Z(DIFF[510]) );
  XOR U1090 ( .A(B[510]), .B(A[510]), .Z(n1090) );
  XOR U1091 ( .A(n1091), .B(n1092), .Z(DIFF[50]) );
  XOR U1092 ( .A(B[50]), .B(A[50]), .Z(n1092) );
  XOR U1093 ( .A(n1093), .B(n1094), .Z(DIFF[509]) );
  XOR U1094 ( .A(B[509]), .B(A[509]), .Z(n1094) );
  XOR U1095 ( .A(n1095), .B(n1096), .Z(DIFF[508]) );
  XOR U1096 ( .A(B[508]), .B(A[508]), .Z(n1096) );
  XOR U1097 ( .A(n1097), .B(n1098), .Z(DIFF[507]) );
  XOR U1098 ( .A(B[507]), .B(A[507]), .Z(n1098) );
  XOR U1099 ( .A(n1099), .B(n1100), .Z(DIFF[506]) );
  XOR U1100 ( .A(B[506]), .B(A[506]), .Z(n1100) );
  XOR U1101 ( .A(n1101), .B(n1102), .Z(DIFF[505]) );
  XOR U1102 ( .A(B[505]), .B(A[505]), .Z(n1102) );
  XOR U1103 ( .A(n1103), .B(n1104), .Z(DIFF[504]) );
  XOR U1104 ( .A(B[504]), .B(A[504]), .Z(n1104) );
  XOR U1105 ( .A(n1105), .B(n1106), .Z(DIFF[503]) );
  XOR U1106 ( .A(B[503]), .B(A[503]), .Z(n1106) );
  XOR U1107 ( .A(n1107), .B(n1108), .Z(DIFF[502]) );
  XOR U1108 ( .A(B[502]), .B(A[502]), .Z(n1108) );
  XOR U1109 ( .A(n1109), .B(n1110), .Z(DIFF[501]) );
  XOR U1110 ( .A(B[501]), .B(A[501]), .Z(n1110) );
  XOR U1111 ( .A(n1111), .B(n1112), .Z(DIFF[500]) );
  XOR U1112 ( .A(B[500]), .B(A[500]), .Z(n1112) );
  XOR U1113 ( .A(n1113), .B(n1114), .Z(DIFF[4]) );
  XOR U1114 ( .A(B[4]), .B(A[4]), .Z(n1114) );
  XOR U1115 ( .A(n1115), .B(n1116), .Z(DIFF[49]) );
  XOR U1116 ( .A(B[49]), .B(A[49]), .Z(n1116) );
  XOR U1117 ( .A(n1117), .B(n1118), .Z(DIFF[499]) );
  XOR U1118 ( .A(B[499]), .B(A[499]), .Z(n1118) );
  XOR U1119 ( .A(n1119), .B(n1120), .Z(DIFF[498]) );
  XOR U1120 ( .A(B[498]), .B(A[498]), .Z(n1120) );
  XOR U1121 ( .A(n1121), .B(n1122), .Z(DIFF[497]) );
  XOR U1122 ( .A(B[497]), .B(A[497]), .Z(n1122) );
  XOR U1123 ( .A(n1123), .B(n1124), .Z(DIFF[496]) );
  XOR U1124 ( .A(B[496]), .B(A[496]), .Z(n1124) );
  XOR U1125 ( .A(n1125), .B(n1126), .Z(DIFF[495]) );
  XOR U1126 ( .A(B[495]), .B(A[495]), .Z(n1126) );
  XOR U1127 ( .A(n1127), .B(n1128), .Z(DIFF[494]) );
  XOR U1128 ( .A(B[494]), .B(A[494]), .Z(n1128) );
  XOR U1129 ( .A(n1129), .B(n1130), .Z(DIFF[493]) );
  XOR U1130 ( .A(B[493]), .B(A[493]), .Z(n1130) );
  XOR U1131 ( .A(n1131), .B(n1132), .Z(DIFF[492]) );
  XOR U1132 ( .A(B[492]), .B(A[492]), .Z(n1132) );
  XOR U1133 ( .A(n1133), .B(n1134), .Z(DIFF[491]) );
  XOR U1134 ( .A(B[491]), .B(A[491]), .Z(n1134) );
  XOR U1135 ( .A(n1135), .B(n1136), .Z(DIFF[490]) );
  XOR U1136 ( .A(B[490]), .B(A[490]), .Z(n1136) );
  XOR U1137 ( .A(n1137), .B(n1138), .Z(DIFF[48]) );
  XOR U1138 ( .A(B[48]), .B(A[48]), .Z(n1138) );
  XOR U1139 ( .A(n1139), .B(n1140), .Z(DIFF[489]) );
  XOR U1140 ( .A(B[489]), .B(A[489]), .Z(n1140) );
  XOR U1141 ( .A(n1141), .B(n1142), .Z(DIFF[488]) );
  XOR U1142 ( .A(B[488]), .B(A[488]), .Z(n1142) );
  XOR U1143 ( .A(n1143), .B(n1144), .Z(DIFF[487]) );
  XOR U1144 ( .A(B[487]), .B(A[487]), .Z(n1144) );
  XOR U1145 ( .A(n1145), .B(n1146), .Z(DIFF[486]) );
  XOR U1146 ( .A(B[486]), .B(A[486]), .Z(n1146) );
  XOR U1147 ( .A(n1147), .B(n1148), .Z(DIFF[485]) );
  XOR U1148 ( .A(B[485]), .B(A[485]), .Z(n1148) );
  XOR U1149 ( .A(n1149), .B(n1150), .Z(DIFF[484]) );
  XOR U1150 ( .A(B[484]), .B(A[484]), .Z(n1150) );
  XOR U1151 ( .A(n1151), .B(n1152), .Z(DIFF[483]) );
  XOR U1152 ( .A(B[483]), .B(A[483]), .Z(n1152) );
  XOR U1153 ( .A(n1153), .B(n1154), .Z(DIFF[482]) );
  XOR U1154 ( .A(B[482]), .B(A[482]), .Z(n1154) );
  XOR U1155 ( .A(n1155), .B(n1156), .Z(DIFF[481]) );
  XOR U1156 ( .A(B[481]), .B(A[481]), .Z(n1156) );
  XOR U1157 ( .A(n1157), .B(n1158), .Z(DIFF[480]) );
  XOR U1158 ( .A(B[480]), .B(A[480]), .Z(n1158) );
  XOR U1159 ( .A(n1159), .B(n1160), .Z(DIFF[47]) );
  XOR U1160 ( .A(B[47]), .B(A[47]), .Z(n1160) );
  XOR U1161 ( .A(n1161), .B(n1162), .Z(DIFF[479]) );
  XOR U1162 ( .A(B[479]), .B(A[479]), .Z(n1162) );
  XOR U1163 ( .A(n1163), .B(n1164), .Z(DIFF[478]) );
  XOR U1164 ( .A(B[478]), .B(A[478]), .Z(n1164) );
  XOR U1165 ( .A(n1165), .B(n1166), .Z(DIFF[477]) );
  XOR U1166 ( .A(B[477]), .B(A[477]), .Z(n1166) );
  XOR U1167 ( .A(n1167), .B(n1168), .Z(DIFF[476]) );
  XOR U1168 ( .A(B[476]), .B(A[476]), .Z(n1168) );
  XOR U1169 ( .A(n1169), .B(n1170), .Z(DIFF[475]) );
  XOR U1170 ( .A(B[475]), .B(A[475]), .Z(n1170) );
  XOR U1171 ( .A(n1171), .B(n1172), .Z(DIFF[474]) );
  XOR U1172 ( .A(B[474]), .B(A[474]), .Z(n1172) );
  XOR U1173 ( .A(n1173), .B(n1174), .Z(DIFF[473]) );
  XOR U1174 ( .A(B[473]), .B(A[473]), .Z(n1174) );
  XOR U1175 ( .A(n1175), .B(n1176), .Z(DIFF[472]) );
  XOR U1176 ( .A(B[472]), .B(A[472]), .Z(n1176) );
  XOR U1177 ( .A(n1177), .B(n1178), .Z(DIFF[471]) );
  XOR U1178 ( .A(B[471]), .B(A[471]), .Z(n1178) );
  XOR U1179 ( .A(n1179), .B(n1180), .Z(DIFF[470]) );
  XOR U1180 ( .A(B[470]), .B(A[470]), .Z(n1180) );
  XOR U1181 ( .A(n1181), .B(n1182), .Z(DIFF[46]) );
  XOR U1182 ( .A(B[46]), .B(A[46]), .Z(n1182) );
  XOR U1183 ( .A(n1183), .B(n1184), .Z(DIFF[469]) );
  XOR U1184 ( .A(B[469]), .B(A[469]), .Z(n1184) );
  XOR U1185 ( .A(n1185), .B(n1186), .Z(DIFF[468]) );
  XOR U1186 ( .A(B[468]), .B(A[468]), .Z(n1186) );
  XOR U1187 ( .A(n1187), .B(n1188), .Z(DIFF[467]) );
  XOR U1188 ( .A(B[467]), .B(A[467]), .Z(n1188) );
  XOR U1189 ( .A(n1189), .B(n1190), .Z(DIFF[466]) );
  XOR U1190 ( .A(B[466]), .B(A[466]), .Z(n1190) );
  XOR U1191 ( .A(n1191), .B(n1192), .Z(DIFF[465]) );
  XOR U1192 ( .A(B[465]), .B(A[465]), .Z(n1192) );
  XOR U1193 ( .A(n1193), .B(n1194), .Z(DIFF[464]) );
  XOR U1194 ( .A(B[464]), .B(A[464]), .Z(n1194) );
  XOR U1195 ( .A(n1195), .B(n1196), .Z(DIFF[463]) );
  XOR U1196 ( .A(B[463]), .B(A[463]), .Z(n1196) );
  XOR U1197 ( .A(n1197), .B(n1198), .Z(DIFF[462]) );
  XOR U1198 ( .A(B[462]), .B(A[462]), .Z(n1198) );
  XOR U1199 ( .A(n1199), .B(n1200), .Z(DIFF[461]) );
  XOR U1200 ( .A(B[461]), .B(A[461]), .Z(n1200) );
  XOR U1201 ( .A(n1201), .B(n1202), .Z(DIFF[460]) );
  XOR U1202 ( .A(B[460]), .B(A[460]), .Z(n1202) );
  XOR U1203 ( .A(n1203), .B(n1204), .Z(DIFF[45]) );
  XOR U1204 ( .A(B[45]), .B(A[45]), .Z(n1204) );
  XOR U1205 ( .A(n1205), .B(n1206), .Z(DIFF[459]) );
  XOR U1206 ( .A(B[459]), .B(A[459]), .Z(n1206) );
  XOR U1207 ( .A(n1207), .B(n1208), .Z(DIFF[458]) );
  XOR U1208 ( .A(B[458]), .B(A[458]), .Z(n1208) );
  XOR U1209 ( .A(n1209), .B(n1210), .Z(DIFF[457]) );
  XOR U1210 ( .A(B[457]), .B(A[457]), .Z(n1210) );
  XOR U1211 ( .A(n1211), .B(n1212), .Z(DIFF[456]) );
  XOR U1212 ( .A(B[456]), .B(A[456]), .Z(n1212) );
  XOR U1213 ( .A(n1213), .B(n1214), .Z(DIFF[455]) );
  XOR U1214 ( .A(B[455]), .B(A[455]), .Z(n1214) );
  XOR U1215 ( .A(n1215), .B(n1216), .Z(DIFF[454]) );
  XOR U1216 ( .A(B[454]), .B(A[454]), .Z(n1216) );
  XOR U1217 ( .A(n1217), .B(n1218), .Z(DIFF[453]) );
  XOR U1218 ( .A(B[453]), .B(A[453]), .Z(n1218) );
  XOR U1219 ( .A(n1219), .B(n1220), .Z(DIFF[452]) );
  XOR U1220 ( .A(B[452]), .B(A[452]), .Z(n1220) );
  XOR U1221 ( .A(n1221), .B(n1222), .Z(DIFF[451]) );
  XOR U1222 ( .A(B[451]), .B(A[451]), .Z(n1222) );
  XOR U1223 ( .A(n1223), .B(n1224), .Z(DIFF[450]) );
  XOR U1224 ( .A(B[450]), .B(A[450]), .Z(n1224) );
  XOR U1225 ( .A(n1225), .B(n1226), .Z(DIFF[44]) );
  XOR U1226 ( .A(B[44]), .B(A[44]), .Z(n1226) );
  XOR U1227 ( .A(n1227), .B(n1228), .Z(DIFF[449]) );
  XOR U1228 ( .A(B[449]), .B(A[449]), .Z(n1228) );
  XOR U1229 ( .A(n1229), .B(n1230), .Z(DIFF[448]) );
  XOR U1230 ( .A(B[448]), .B(A[448]), .Z(n1230) );
  XOR U1231 ( .A(n1231), .B(n1232), .Z(DIFF[447]) );
  XOR U1232 ( .A(B[447]), .B(A[447]), .Z(n1232) );
  XOR U1233 ( .A(n1233), .B(n1234), .Z(DIFF[446]) );
  XOR U1234 ( .A(B[446]), .B(A[446]), .Z(n1234) );
  XOR U1235 ( .A(n1235), .B(n1236), .Z(DIFF[445]) );
  XOR U1236 ( .A(B[445]), .B(A[445]), .Z(n1236) );
  XOR U1237 ( .A(n1237), .B(n1238), .Z(DIFF[444]) );
  XOR U1238 ( .A(B[444]), .B(A[444]), .Z(n1238) );
  XOR U1239 ( .A(n1239), .B(n1240), .Z(DIFF[443]) );
  XOR U1240 ( .A(B[443]), .B(A[443]), .Z(n1240) );
  XOR U1241 ( .A(n1241), .B(n1242), .Z(DIFF[442]) );
  XOR U1242 ( .A(B[442]), .B(A[442]), .Z(n1242) );
  XOR U1243 ( .A(n1243), .B(n1244), .Z(DIFF[441]) );
  XOR U1244 ( .A(B[441]), .B(A[441]), .Z(n1244) );
  XOR U1245 ( .A(n1245), .B(n1246), .Z(DIFF[440]) );
  XOR U1246 ( .A(B[440]), .B(A[440]), .Z(n1246) );
  XOR U1247 ( .A(n1247), .B(n1248), .Z(DIFF[43]) );
  XOR U1248 ( .A(B[43]), .B(A[43]), .Z(n1248) );
  XOR U1249 ( .A(n1249), .B(n1250), .Z(DIFF[439]) );
  XOR U1250 ( .A(B[439]), .B(A[439]), .Z(n1250) );
  XOR U1251 ( .A(n1251), .B(n1252), .Z(DIFF[438]) );
  XOR U1252 ( .A(B[438]), .B(A[438]), .Z(n1252) );
  XOR U1253 ( .A(n1253), .B(n1254), .Z(DIFF[437]) );
  XOR U1254 ( .A(B[437]), .B(A[437]), .Z(n1254) );
  XOR U1255 ( .A(n1255), .B(n1256), .Z(DIFF[436]) );
  XOR U1256 ( .A(B[436]), .B(A[436]), .Z(n1256) );
  XOR U1257 ( .A(n1257), .B(n1258), .Z(DIFF[435]) );
  XOR U1258 ( .A(B[435]), .B(A[435]), .Z(n1258) );
  XOR U1259 ( .A(n1259), .B(n1260), .Z(DIFF[434]) );
  XOR U1260 ( .A(B[434]), .B(A[434]), .Z(n1260) );
  XOR U1261 ( .A(n1261), .B(n1262), .Z(DIFF[433]) );
  XOR U1262 ( .A(B[433]), .B(A[433]), .Z(n1262) );
  XOR U1263 ( .A(n1263), .B(n1264), .Z(DIFF[432]) );
  XOR U1264 ( .A(B[432]), .B(A[432]), .Z(n1264) );
  XOR U1265 ( .A(n1265), .B(n1266), .Z(DIFF[431]) );
  XOR U1266 ( .A(B[431]), .B(A[431]), .Z(n1266) );
  XOR U1267 ( .A(n1267), .B(n1268), .Z(DIFF[430]) );
  XOR U1268 ( .A(B[430]), .B(A[430]), .Z(n1268) );
  XOR U1269 ( .A(n1269), .B(n1270), .Z(DIFF[42]) );
  XOR U1270 ( .A(B[42]), .B(A[42]), .Z(n1270) );
  XOR U1271 ( .A(n1271), .B(n1272), .Z(DIFF[429]) );
  XOR U1272 ( .A(B[429]), .B(A[429]), .Z(n1272) );
  XOR U1273 ( .A(n1273), .B(n1274), .Z(DIFF[428]) );
  XOR U1274 ( .A(B[428]), .B(A[428]), .Z(n1274) );
  XOR U1275 ( .A(n1275), .B(n1276), .Z(DIFF[427]) );
  XOR U1276 ( .A(B[427]), .B(A[427]), .Z(n1276) );
  XOR U1277 ( .A(n1277), .B(n1278), .Z(DIFF[426]) );
  XOR U1278 ( .A(B[426]), .B(A[426]), .Z(n1278) );
  XOR U1279 ( .A(n1279), .B(n1280), .Z(DIFF[425]) );
  XOR U1280 ( .A(B[425]), .B(A[425]), .Z(n1280) );
  XOR U1281 ( .A(n1281), .B(n1282), .Z(DIFF[424]) );
  XOR U1282 ( .A(B[424]), .B(A[424]), .Z(n1282) );
  XOR U1283 ( .A(n1283), .B(n1284), .Z(DIFF[423]) );
  XOR U1284 ( .A(B[423]), .B(A[423]), .Z(n1284) );
  XOR U1285 ( .A(n1285), .B(n1286), .Z(DIFF[422]) );
  XOR U1286 ( .A(B[422]), .B(A[422]), .Z(n1286) );
  XOR U1287 ( .A(n1287), .B(n1288), .Z(DIFF[421]) );
  XOR U1288 ( .A(B[421]), .B(A[421]), .Z(n1288) );
  XOR U1289 ( .A(n1289), .B(n1290), .Z(DIFF[420]) );
  XOR U1290 ( .A(B[420]), .B(A[420]), .Z(n1290) );
  XOR U1291 ( .A(n1291), .B(n1292), .Z(DIFF[41]) );
  XOR U1292 ( .A(B[41]), .B(A[41]), .Z(n1292) );
  XOR U1293 ( .A(n1293), .B(n1294), .Z(DIFF[419]) );
  XOR U1294 ( .A(B[419]), .B(A[419]), .Z(n1294) );
  XOR U1295 ( .A(n1295), .B(n1296), .Z(DIFF[418]) );
  XOR U1296 ( .A(B[418]), .B(A[418]), .Z(n1296) );
  XOR U1297 ( .A(n1297), .B(n1298), .Z(DIFF[417]) );
  XOR U1298 ( .A(B[417]), .B(A[417]), .Z(n1298) );
  XOR U1299 ( .A(n1299), .B(n1300), .Z(DIFF[416]) );
  XOR U1300 ( .A(B[416]), .B(A[416]), .Z(n1300) );
  XOR U1301 ( .A(n1301), .B(n1302), .Z(DIFF[415]) );
  XOR U1302 ( .A(B[415]), .B(A[415]), .Z(n1302) );
  XOR U1303 ( .A(n1303), .B(n1304), .Z(DIFF[414]) );
  XOR U1304 ( .A(B[414]), .B(A[414]), .Z(n1304) );
  XOR U1305 ( .A(n1305), .B(n1306), .Z(DIFF[413]) );
  XOR U1306 ( .A(B[413]), .B(A[413]), .Z(n1306) );
  XOR U1307 ( .A(n1307), .B(n1308), .Z(DIFF[412]) );
  XOR U1308 ( .A(B[412]), .B(A[412]), .Z(n1308) );
  XOR U1309 ( .A(n1309), .B(n1310), .Z(DIFF[411]) );
  XOR U1310 ( .A(B[411]), .B(A[411]), .Z(n1310) );
  XOR U1311 ( .A(n1311), .B(n1312), .Z(DIFF[410]) );
  XOR U1312 ( .A(B[410]), .B(A[410]), .Z(n1312) );
  XOR U1313 ( .A(n1313), .B(n1314), .Z(DIFF[40]) );
  XOR U1314 ( .A(B[40]), .B(A[40]), .Z(n1314) );
  XOR U1315 ( .A(n1315), .B(n1316), .Z(DIFF[409]) );
  XOR U1316 ( .A(B[409]), .B(A[409]), .Z(n1316) );
  XOR U1317 ( .A(n1317), .B(n1318), .Z(DIFF[408]) );
  XOR U1318 ( .A(B[408]), .B(A[408]), .Z(n1318) );
  XOR U1319 ( .A(n1319), .B(n1320), .Z(DIFF[407]) );
  XOR U1320 ( .A(B[407]), .B(A[407]), .Z(n1320) );
  XOR U1321 ( .A(n1321), .B(n1322), .Z(DIFF[406]) );
  XOR U1322 ( .A(B[406]), .B(A[406]), .Z(n1322) );
  XOR U1323 ( .A(n1323), .B(n1324), .Z(DIFF[405]) );
  XOR U1324 ( .A(B[405]), .B(A[405]), .Z(n1324) );
  XOR U1325 ( .A(n1325), .B(n1326), .Z(DIFF[404]) );
  XOR U1326 ( .A(B[404]), .B(A[404]), .Z(n1326) );
  XOR U1327 ( .A(n1327), .B(n1328), .Z(DIFF[403]) );
  XOR U1328 ( .A(B[403]), .B(A[403]), .Z(n1328) );
  XOR U1329 ( .A(n1329), .B(n1330), .Z(DIFF[402]) );
  XOR U1330 ( .A(B[402]), .B(A[402]), .Z(n1330) );
  XOR U1331 ( .A(n1331), .B(n1332), .Z(DIFF[401]) );
  XOR U1332 ( .A(B[401]), .B(A[401]), .Z(n1332) );
  XOR U1333 ( .A(n1333), .B(n1334), .Z(DIFF[400]) );
  XOR U1334 ( .A(B[400]), .B(A[400]), .Z(n1334) );
  XOR U1335 ( .A(n1335), .B(n1336), .Z(DIFF[3]) );
  XOR U1336 ( .A(B[3]), .B(A[3]), .Z(n1336) );
  XOR U1337 ( .A(n1337), .B(n1338), .Z(DIFF[39]) );
  XOR U1338 ( .A(B[39]), .B(A[39]), .Z(n1338) );
  XOR U1339 ( .A(n1339), .B(n1340), .Z(DIFF[399]) );
  XOR U1340 ( .A(B[399]), .B(A[399]), .Z(n1340) );
  XOR U1341 ( .A(n1341), .B(n1342), .Z(DIFF[398]) );
  XOR U1342 ( .A(B[398]), .B(A[398]), .Z(n1342) );
  XOR U1343 ( .A(n1343), .B(n1344), .Z(DIFF[397]) );
  XOR U1344 ( .A(B[397]), .B(A[397]), .Z(n1344) );
  XOR U1345 ( .A(n1345), .B(n1346), .Z(DIFF[396]) );
  XOR U1346 ( .A(B[396]), .B(A[396]), .Z(n1346) );
  XOR U1347 ( .A(n1347), .B(n1348), .Z(DIFF[395]) );
  XOR U1348 ( .A(B[395]), .B(A[395]), .Z(n1348) );
  XOR U1349 ( .A(n1349), .B(n1350), .Z(DIFF[394]) );
  XOR U1350 ( .A(B[394]), .B(A[394]), .Z(n1350) );
  XOR U1351 ( .A(n1351), .B(n1352), .Z(DIFF[393]) );
  XOR U1352 ( .A(B[393]), .B(A[393]), .Z(n1352) );
  XOR U1353 ( .A(n1353), .B(n1354), .Z(DIFF[392]) );
  XOR U1354 ( .A(B[392]), .B(A[392]), .Z(n1354) );
  XOR U1355 ( .A(n1355), .B(n1356), .Z(DIFF[391]) );
  XOR U1356 ( .A(B[391]), .B(A[391]), .Z(n1356) );
  XOR U1357 ( .A(n1357), .B(n1358), .Z(DIFF[390]) );
  XOR U1358 ( .A(B[390]), .B(A[390]), .Z(n1358) );
  XOR U1359 ( .A(n1359), .B(n1360), .Z(DIFF[38]) );
  XOR U1360 ( .A(B[38]), .B(A[38]), .Z(n1360) );
  XOR U1361 ( .A(n1361), .B(n1362), .Z(DIFF[389]) );
  XOR U1362 ( .A(B[389]), .B(A[389]), .Z(n1362) );
  XOR U1363 ( .A(n1363), .B(n1364), .Z(DIFF[388]) );
  XOR U1364 ( .A(B[388]), .B(A[388]), .Z(n1364) );
  XOR U1365 ( .A(n1365), .B(n1366), .Z(DIFF[387]) );
  XOR U1366 ( .A(B[387]), .B(A[387]), .Z(n1366) );
  XOR U1367 ( .A(n1367), .B(n1368), .Z(DIFF[386]) );
  XOR U1368 ( .A(B[386]), .B(A[386]), .Z(n1368) );
  XOR U1369 ( .A(n1369), .B(n1370), .Z(DIFF[385]) );
  XOR U1370 ( .A(B[385]), .B(A[385]), .Z(n1370) );
  XOR U1371 ( .A(n1371), .B(n1372), .Z(DIFF[384]) );
  XOR U1372 ( .A(B[384]), .B(A[384]), .Z(n1372) );
  XOR U1373 ( .A(n1373), .B(n1374), .Z(DIFF[383]) );
  XOR U1374 ( .A(B[383]), .B(A[383]), .Z(n1374) );
  XOR U1375 ( .A(n1375), .B(n1376), .Z(DIFF[382]) );
  XOR U1376 ( .A(B[382]), .B(A[382]), .Z(n1376) );
  XOR U1377 ( .A(n1377), .B(n1378), .Z(DIFF[381]) );
  XOR U1378 ( .A(B[381]), .B(A[381]), .Z(n1378) );
  XOR U1379 ( .A(n1379), .B(n1380), .Z(DIFF[380]) );
  XOR U1380 ( .A(B[380]), .B(A[380]), .Z(n1380) );
  XOR U1381 ( .A(n1381), .B(n1382), .Z(DIFF[37]) );
  XOR U1382 ( .A(B[37]), .B(A[37]), .Z(n1382) );
  XOR U1383 ( .A(n1383), .B(n1384), .Z(DIFF[379]) );
  XOR U1384 ( .A(B[379]), .B(A[379]), .Z(n1384) );
  XOR U1385 ( .A(n1385), .B(n1386), .Z(DIFF[378]) );
  XOR U1386 ( .A(B[378]), .B(A[378]), .Z(n1386) );
  XOR U1387 ( .A(n1387), .B(n1388), .Z(DIFF[377]) );
  XOR U1388 ( .A(B[377]), .B(A[377]), .Z(n1388) );
  XOR U1389 ( .A(n1389), .B(n1390), .Z(DIFF[376]) );
  XOR U1390 ( .A(B[376]), .B(A[376]), .Z(n1390) );
  XOR U1391 ( .A(n1391), .B(n1392), .Z(DIFF[375]) );
  XOR U1392 ( .A(B[375]), .B(A[375]), .Z(n1392) );
  XOR U1393 ( .A(n1393), .B(n1394), .Z(DIFF[374]) );
  XOR U1394 ( .A(B[374]), .B(A[374]), .Z(n1394) );
  XOR U1395 ( .A(n1395), .B(n1396), .Z(DIFF[373]) );
  XOR U1396 ( .A(B[373]), .B(A[373]), .Z(n1396) );
  XOR U1397 ( .A(n1397), .B(n1398), .Z(DIFF[372]) );
  XOR U1398 ( .A(B[372]), .B(A[372]), .Z(n1398) );
  XOR U1399 ( .A(n1399), .B(n1400), .Z(DIFF[371]) );
  XOR U1400 ( .A(B[371]), .B(A[371]), .Z(n1400) );
  XOR U1401 ( .A(n1401), .B(n1402), .Z(DIFF[370]) );
  XOR U1402 ( .A(B[370]), .B(A[370]), .Z(n1402) );
  XOR U1403 ( .A(n1403), .B(n1404), .Z(DIFF[36]) );
  XOR U1404 ( .A(B[36]), .B(A[36]), .Z(n1404) );
  XOR U1405 ( .A(n1405), .B(n1406), .Z(DIFF[369]) );
  XOR U1406 ( .A(B[369]), .B(A[369]), .Z(n1406) );
  XOR U1407 ( .A(n1407), .B(n1408), .Z(DIFF[368]) );
  XOR U1408 ( .A(B[368]), .B(A[368]), .Z(n1408) );
  XOR U1409 ( .A(n1409), .B(n1410), .Z(DIFF[367]) );
  XOR U1410 ( .A(B[367]), .B(A[367]), .Z(n1410) );
  XOR U1411 ( .A(n1411), .B(n1412), .Z(DIFF[366]) );
  XOR U1412 ( .A(B[366]), .B(A[366]), .Z(n1412) );
  XOR U1413 ( .A(n1413), .B(n1414), .Z(DIFF[365]) );
  XOR U1414 ( .A(B[365]), .B(A[365]), .Z(n1414) );
  XOR U1415 ( .A(n1415), .B(n1416), .Z(DIFF[364]) );
  XOR U1416 ( .A(B[364]), .B(A[364]), .Z(n1416) );
  XOR U1417 ( .A(n1417), .B(n1418), .Z(DIFF[363]) );
  XOR U1418 ( .A(B[363]), .B(A[363]), .Z(n1418) );
  XOR U1419 ( .A(n1419), .B(n1420), .Z(DIFF[362]) );
  XOR U1420 ( .A(B[362]), .B(A[362]), .Z(n1420) );
  XOR U1421 ( .A(n1421), .B(n1422), .Z(DIFF[361]) );
  XOR U1422 ( .A(B[361]), .B(A[361]), .Z(n1422) );
  XOR U1423 ( .A(n1423), .B(n1424), .Z(DIFF[360]) );
  XOR U1424 ( .A(B[360]), .B(A[360]), .Z(n1424) );
  XOR U1425 ( .A(n1425), .B(n1426), .Z(DIFF[35]) );
  XOR U1426 ( .A(B[35]), .B(A[35]), .Z(n1426) );
  XOR U1427 ( .A(n1427), .B(n1428), .Z(DIFF[359]) );
  XOR U1428 ( .A(B[359]), .B(A[359]), .Z(n1428) );
  XOR U1429 ( .A(n1429), .B(n1430), .Z(DIFF[358]) );
  XOR U1430 ( .A(B[358]), .B(A[358]), .Z(n1430) );
  XOR U1431 ( .A(n1431), .B(n1432), .Z(DIFF[357]) );
  XOR U1432 ( .A(B[357]), .B(A[357]), .Z(n1432) );
  XOR U1433 ( .A(n1433), .B(n1434), .Z(DIFF[356]) );
  XOR U1434 ( .A(B[356]), .B(A[356]), .Z(n1434) );
  XOR U1435 ( .A(n1435), .B(n1436), .Z(DIFF[355]) );
  XOR U1436 ( .A(B[355]), .B(A[355]), .Z(n1436) );
  XOR U1437 ( .A(n1437), .B(n1438), .Z(DIFF[354]) );
  XOR U1438 ( .A(B[354]), .B(A[354]), .Z(n1438) );
  XOR U1439 ( .A(n1439), .B(n1440), .Z(DIFF[353]) );
  XOR U1440 ( .A(B[353]), .B(A[353]), .Z(n1440) );
  XOR U1441 ( .A(n1441), .B(n1442), .Z(DIFF[352]) );
  XOR U1442 ( .A(B[352]), .B(A[352]), .Z(n1442) );
  XOR U1443 ( .A(n1443), .B(n1444), .Z(DIFF[351]) );
  XOR U1444 ( .A(B[351]), .B(A[351]), .Z(n1444) );
  XOR U1445 ( .A(n1445), .B(n1446), .Z(DIFF[350]) );
  XOR U1446 ( .A(B[350]), .B(A[350]), .Z(n1446) );
  XOR U1447 ( .A(n1447), .B(n1448), .Z(DIFF[34]) );
  XOR U1448 ( .A(B[34]), .B(A[34]), .Z(n1448) );
  XOR U1449 ( .A(n1449), .B(n1450), .Z(DIFF[349]) );
  XOR U1450 ( .A(B[349]), .B(A[349]), .Z(n1450) );
  XOR U1451 ( .A(n1451), .B(n1452), .Z(DIFF[348]) );
  XOR U1452 ( .A(B[348]), .B(A[348]), .Z(n1452) );
  XOR U1453 ( .A(n1453), .B(n1454), .Z(DIFF[347]) );
  XOR U1454 ( .A(B[347]), .B(A[347]), .Z(n1454) );
  XOR U1455 ( .A(n1455), .B(n1456), .Z(DIFF[346]) );
  XOR U1456 ( .A(B[346]), .B(A[346]), .Z(n1456) );
  XOR U1457 ( .A(n1457), .B(n1458), .Z(DIFF[345]) );
  XOR U1458 ( .A(B[345]), .B(A[345]), .Z(n1458) );
  XOR U1459 ( .A(n1459), .B(n1460), .Z(DIFF[344]) );
  XOR U1460 ( .A(B[344]), .B(A[344]), .Z(n1460) );
  XOR U1461 ( .A(n1461), .B(n1462), .Z(DIFF[343]) );
  XOR U1462 ( .A(B[343]), .B(A[343]), .Z(n1462) );
  XOR U1463 ( .A(n1463), .B(n1464), .Z(DIFF[342]) );
  XOR U1464 ( .A(B[342]), .B(A[342]), .Z(n1464) );
  XOR U1465 ( .A(n1465), .B(n1466), .Z(DIFF[341]) );
  XOR U1466 ( .A(B[341]), .B(A[341]), .Z(n1466) );
  XOR U1467 ( .A(n1467), .B(n1468), .Z(DIFF[340]) );
  XOR U1468 ( .A(B[340]), .B(A[340]), .Z(n1468) );
  XOR U1469 ( .A(n1469), .B(n1470), .Z(DIFF[33]) );
  XOR U1470 ( .A(B[33]), .B(A[33]), .Z(n1470) );
  XOR U1471 ( .A(n1471), .B(n1472), .Z(DIFF[339]) );
  XOR U1472 ( .A(B[339]), .B(A[339]), .Z(n1472) );
  XOR U1473 ( .A(n1473), .B(n1474), .Z(DIFF[338]) );
  XOR U1474 ( .A(B[338]), .B(A[338]), .Z(n1474) );
  XOR U1475 ( .A(n1475), .B(n1476), .Z(DIFF[337]) );
  XOR U1476 ( .A(B[337]), .B(A[337]), .Z(n1476) );
  XOR U1477 ( .A(n1477), .B(n1478), .Z(DIFF[336]) );
  XOR U1478 ( .A(B[336]), .B(A[336]), .Z(n1478) );
  XOR U1479 ( .A(n1479), .B(n1480), .Z(DIFF[335]) );
  XOR U1480 ( .A(B[335]), .B(A[335]), .Z(n1480) );
  XOR U1481 ( .A(n1481), .B(n1482), .Z(DIFF[334]) );
  XOR U1482 ( .A(B[334]), .B(A[334]), .Z(n1482) );
  XOR U1483 ( .A(n1483), .B(n1484), .Z(DIFF[333]) );
  XOR U1484 ( .A(B[333]), .B(A[333]), .Z(n1484) );
  XOR U1485 ( .A(n1485), .B(n1486), .Z(DIFF[332]) );
  XOR U1486 ( .A(B[332]), .B(A[332]), .Z(n1486) );
  XOR U1487 ( .A(n1487), .B(n1488), .Z(DIFF[331]) );
  XOR U1488 ( .A(B[331]), .B(A[331]), .Z(n1488) );
  XOR U1489 ( .A(n1489), .B(n1490), .Z(DIFF[330]) );
  XOR U1490 ( .A(B[330]), .B(A[330]), .Z(n1490) );
  XOR U1491 ( .A(n1491), .B(n1492), .Z(DIFF[32]) );
  XOR U1492 ( .A(B[32]), .B(A[32]), .Z(n1492) );
  XOR U1493 ( .A(n1493), .B(n1494), .Z(DIFF[329]) );
  XOR U1494 ( .A(B[329]), .B(A[329]), .Z(n1494) );
  XOR U1495 ( .A(n1495), .B(n1496), .Z(DIFF[328]) );
  XOR U1496 ( .A(B[328]), .B(A[328]), .Z(n1496) );
  XOR U1497 ( .A(n1497), .B(n1498), .Z(DIFF[327]) );
  XOR U1498 ( .A(B[327]), .B(A[327]), .Z(n1498) );
  XOR U1499 ( .A(n1499), .B(n1500), .Z(DIFF[326]) );
  XOR U1500 ( .A(B[326]), .B(A[326]), .Z(n1500) );
  XOR U1501 ( .A(n1501), .B(n1502), .Z(DIFF[325]) );
  XOR U1502 ( .A(B[325]), .B(A[325]), .Z(n1502) );
  XOR U1503 ( .A(n1503), .B(n1504), .Z(DIFF[324]) );
  XOR U1504 ( .A(B[324]), .B(A[324]), .Z(n1504) );
  XOR U1505 ( .A(n1505), .B(n1506), .Z(DIFF[323]) );
  XOR U1506 ( .A(B[323]), .B(A[323]), .Z(n1506) );
  XOR U1507 ( .A(n1507), .B(n1508), .Z(DIFF[322]) );
  XOR U1508 ( .A(B[322]), .B(A[322]), .Z(n1508) );
  XOR U1509 ( .A(n1509), .B(n1510), .Z(DIFF[321]) );
  XOR U1510 ( .A(B[321]), .B(A[321]), .Z(n1510) );
  XOR U1511 ( .A(n1511), .B(n1512), .Z(DIFF[320]) );
  XOR U1512 ( .A(B[320]), .B(A[320]), .Z(n1512) );
  XOR U1513 ( .A(n1513), .B(n1514), .Z(DIFF[31]) );
  XOR U1514 ( .A(B[31]), .B(A[31]), .Z(n1514) );
  XOR U1515 ( .A(n1515), .B(n1516), .Z(DIFF[319]) );
  XOR U1516 ( .A(B[319]), .B(A[319]), .Z(n1516) );
  XOR U1517 ( .A(n1517), .B(n1518), .Z(DIFF[318]) );
  XOR U1518 ( .A(B[318]), .B(A[318]), .Z(n1518) );
  XOR U1519 ( .A(n1519), .B(n1520), .Z(DIFF[317]) );
  XOR U1520 ( .A(B[317]), .B(A[317]), .Z(n1520) );
  XOR U1521 ( .A(n1521), .B(n1522), .Z(DIFF[316]) );
  XOR U1522 ( .A(B[316]), .B(A[316]), .Z(n1522) );
  XOR U1523 ( .A(n1523), .B(n1524), .Z(DIFF[315]) );
  XOR U1524 ( .A(B[315]), .B(A[315]), .Z(n1524) );
  XOR U1525 ( .A(n1525), .B(n1526), .Z(DIFF[314]) );
  XOR U1526 ( .A(B[314]), .B(A[314]), .Z(n1526) );
  XOR U1527 ( .A(n1527), .B(n1528), .Z(DIFF[313]) );
  XOR U1528 ( .A(B[313]), .B(A[313]), .Z(n1528) );
  XOR U1529 ( .A(n1529), .B(n1530), .Z(DIFF[312]) );
  XOR U1530 ( .A(B[312]), .B(A[312]), .Z(n1530) );
  XOR U1531 ( .A(n1531), .B(n1532), .Z(DIFF[311]) );
  XOR U1532 ( .A(B[311]), .B(A[311]), .Z(n1532) );
  XOR U1533 ( .A(n1533), .B(n1534), .Z(DIFF[310]) );
  XOR U1534 ( .A(B[310]), .B(A[310]), .Z(n1534) );
  XOR U1535 ( .A(n1535), .B(n1536), .Z(DIFF[30]) );
  XOR U1536 ( .A(B[30]), .B(A[30]), .Z(n1536) );
  XOR U1537 ( .A(n1537), .B(n1538), .Z(DIFF[309]) );
  XOR U1538 ( .A(B[309]), .B(A[309]), .Z(n1538) );
  XOR U1539 ( .A(n1539), .B(n1540), .Z(DIFF[308]) );
  XOR U1540 ( .A(B[308]), .B(A[308]), .Z(n1540) );
  XOR U1541 ( .A(n1541), .B(n1542), .Z(DIFF[307]) );
  XOR U1542 ( .A(B[307]), .B(A[307]), .Z(n1542) );
  XOR U1543 ( .A(n1543), .B(n1544), .Z(DIFF[306]) );
  XOR U1544 ( .A(B[306]), .B(A[306]), .Z(n1544) );
  XOR U1545 ( .A(n1545), .B(n1546), .Z(DIFF[305]) );
  XOR U1546 ( .A(B[305]), .B(A[305]), .Z(n1546) );
  XOR U1547 ( .A(n1547), .B(n1548), .Z(DIFF[304]) );
  XOR U1548 ( .A(B[304]), .B(A[304]), .Z(n1548) );
  XOR U1549 ( .A(n1549), .B(n1550), .Z(DIFF[303]) );
  XOR U1550 ( .A(B[303]), .B(A[303]), .Z(n1550) );
  XOR U1551 ( .A(n1551), .B(n1552), .Z(DIFF[302]) );
  XOR U1552 ( .A(B[302]), .B(A[302]), .Z(n1552) );
  XOR U1553 ( .A(n1553), .B(n1554), .Z(DIFF[301]) );
  XOR U1554 ( .A(B[301]), .B(A[301]), .Z(n1554) );
  XOR U1555 ( .A(n1555), .B(n1556), .Z(DIFF[300]) );
  XOR U1556 ( .A(B[300]), .B(A[300]), .Z(n1556) );
  XOR U1557 ( .A(n1557), .B(n1558), .Z(DIFF[2]) );
  XOR U1558 ( .A(B[2]), .B(A[2]), .Z(n1558) );
  XOR U1559 ( .A(n1559), .B(n1560), .Z(DIFF[29]) );
  XOR U1560 ( .A(B[29]), .B(A[29]), .Z(n1560) );
  XOR U1561 ( .A(n1561), .B(n1562), .Z(DIFF[299]) );
  XOR U1562 ( .A(B[299]), .B(A[299]), .Z(n1562) );
  XOR U1563 ( .A(n1563), .B(n1564), .Z(DIFF[298]) );
  XOR U1564 ( .A(B[298]), .B(A[298]), .Z(n1564) );
  XOR U1565 ( .A(n1565), .B(n1566), .Z(DIFF[297]) );
  XOR U1566 ( .A(B[297]), .B(A[297]), .Z(n1566) );
  XOR U1567 ( .A(n1567), .B(n1568), .Z(DIFF[296]) );
  XOR U1568 ( .A(B[296]), .B(A[296]), .Z(n1568) );
  XOR U1569 ( .A(n1569), .B(n1570), .Z(DIFF[295]) );
  XOR U1570 ( .A(B[295]), .B(A[295]), .Z(n1570) );
  XOR U1571 ( .A(n1571), .B(n1572), .Z(DIFF[294]) );
  XOR U1572 ( .A(B[294]), .B(A[294]), .Z(n1572) );
  XOR U1573 ( .A(n1573), .B(n1574), .Z(DIFF[293]) );
  XOR U1574 ( .A(B[293]), .B(A[293]), .Z(n1574) );
  XOR U1575 ( .A(n1575), .B(n1576), .Z(DIFF[292]) );
  XOR U1576 ( .A(B[292]), .B(A[292]), .Z(n1576) );
  XOR U1577 ( .A(n1577), .B(n1578), .Z(DIFF[291]) );
  XOR U1578 ( .A(B[291]), .B(A[291]), .Z(n1578) );
  XOR U1579 ( .A(n1579), .B(n1580), .Z(DIFF[290]) );
  XOR U1580 ( .A(B[290]), .B(A[290]), .Z(n1580) );
  XOR U1581 ( .A(n1581), .B(n1582), .Z(DIFF[28]) );
  XOR U1582 ( .A(B[28]), .B(A[28]), .Z(n1582) );
  XOR U1583 ( .A(n1583), .B(n1584), .Z(DIFF[289]) );
  XOR U1584 ( .A(B[289]), .B(A[289]), .Z(n1584) );
  XOR U1585 ( .A(n1585), .B(n1586), .Z(DIFF[288]) );
  XOR U1586 ( .A(B[288]), .B(A[288]), .Z(n1586) );
  XOR U1587 ( .A(n1587), .B(n1588), .Z(DIFF[287]) );
  XOR U1588 ( .A(B[287]), .B(A[287]), .Z(n1588) );
  XOR U1589 ( .A(n1589), .B(n1590), .Z(DIFF[286]) );
  XOR U1590 ( .A(B[286]), .B(A[286]), .Z(n1590) );
  XOR U1591 ( .A(n1591), .B(n1592), .Z(DIFF[285]) );
  XOR U1592 ( .A(B[285]), .B(A[285]), .Z(n1592) );
  XOR U1593 ( .A(n1593), .B(n1594), .Z(DIFF[284]) );
  XOR U1594 ( .A(B[284]), .B(A[284]), .Z(n1594) );
  XOR U1595 ( .A(n1595), .B(n1596), .Z(DIFF[283]) );
  XOR U1596 ( .A(B[283]), .B(A[283]), .Z(n1596) );
  XOR U1597 ( .A(n1597), .B(n1598), .Z(DIFF[282]) );
  XOR U1598 ( .A(B[282]), .B(A[282]), .Z(n1598) );
  XOR U1599 ( .A(n1599), .B(n1600), .Z(DIFF[281]) );
  XOR U1600 ( .A(B[281]), .B(A[281]), .Z(n1600) );
  XOR U1601 ( .A(n1601), .B(n1602), .Z(DIFF[280]) );
  XOR U1602 ( .A(B[280]), .B(A[280]), .Z(n1602) );
  XOR U1603 ( .A(n1603), .B(n1604), .Z(DIFF[27]) );
  XOR U1604 ( .A(B[27]), .B(A[27]), .Z(n1604) );
  XOR U1605 ( .A(n1605), .B(n1606), .Z(DIFF[279]) );
  XOR U1606 ( .A(B[279]), .B(A[279]), .Z(n1606) );
  XOR U1607 ( .A(n1607), .B(n1608), .Z(DIFF[278]) );
  XOR U1608 ( .A(B[278]), .B(A[278]), .Z(n1608) );
  XOR U1609 ( .A(n1609), .B(n1610), .Z(DIFF[277]) );
  XOR U1610 ( .A(B[277]), .B(A[277]), .Z(n1610) );
  XOR U1611 ( .A(n1611), .B(n1612), .Z(DIFF[276]) );
  XOR U1612 ( .A(B[276]), .B(A[276]), .Z(n1612) );
  XOR U1613 ( .A(n1613), .B(n1614), .Z(DIFF[275]) );
  XOR U1614 ( .A(B[275]), .B(A[275]), .Z(n1614) );
  XOR U1615 ( .A(n1615), .B(n1616), .Z(DIFF[274]) );
  XOR U1616 ( .A(B[274]), .B(A[274]), .Z(n1616) );
  XOR U1617 ( .A(n1617), .B(n1618), .Z(DIFF[273]) );
  XOR U1618 ( .A(B[273]), .B(A[273]), .Z(n1618) );
  XOR U1619 ( .A(n1619), .B(n1620), .Z(DIFF[272]) );
  XOR U1620 ( .A(B[272]), .B(A[272]), .Z(n1620) );
  XOR U1621 ( .A(n1621), .B(n1622), .Z(DIFF[271]) );
  XOR U1622 ( .A(B[271]), .B(A[271]), .Z(n1622) );
  XOR U1623 ( .A(n1623), .B(n1624), .Z(DIFF[270]) );
  XOR U1624 ( .A(B[270]), .B(A[270]), .Z(n1624) );
  XOR U1625 ( .A(n1625), .B(n1626), .Z(DIFF[26]) );
  XOR U1626 ( .A(B[26]), .B(A[26]), .Z(n1626) );
  XOR U1627 ( .A(n1627), .B(n1628), .Z(DIFF[269]) );
  XOR U1628 ( .A(B[269]), .B(A[269]), .Z(n1628) );
  XOR U1629 ( .A(n1629), .B(n1630), .Z(DIFF[268]) );
  XOR U1630 ( .A(B[268]), .B(A[268]), .Z(n1630) );
  XOR U1631 ( .A(n1631), .B(n1632), .Z(DIFF[267]) );
  XOR U1632 ( .A(B[267]), .B(A[267]), .Z(n1632) );
  XOR U1633 ( .A(n1633), .B(n1634), .Z(DIFF[266]) );
  XOR U1634 ( .A(B[266]), .B(A[266]), .Z(n1634) );
  XOR U1635 ( .A(n1635), .B(n1636), .Z(DIFF[265]) );
  XOR U1636 ( .A(B[265]), .B(A[265]), .Z(n1636) );
  XOR U1637 ( .A(n1637), .B(n1638), .Z(DIFF[264]) );
  XOR U1638 ( .A(B[264]), .B(A[264]), .Z(n1638) );
  XOR U1639 ( .A(n1639), .B(n1640), .Z(DIFF[263]) );
  XOR U1640 ( .A(B[263]), .B(A[263]), .Z(n1640) );
  XOR U1641 ( .A(n1641), .B(n1642), .Z(DIFF[262]) );
  XOR U1642 ( .A(B[262]), .B(A[262]), .Z(n1642) );
  XOR U1643 ( .A(n1643), .B(n1644), .Z(DIFF[261]) );
  XOR U1644 ( .A(B[261]), .B(A[261]), .Z(n1644) );
  XOR U1645 ( .A(n1645), .B(n1646), .Z(DIFF[260]) );
  XOR U1646 ( .A(B[260]), .B(A[260]), .Z(n1646) );
  XOR U1647 ( .A(n1647), .B(n1648), .Z(DIFF[25]) );
  XOR U1648 ( .A(B[25]), .B(A[25]), .Z(n1648) );
  XOR U1649 ( .A(n1649), .B(n1650), .Z(DIFF[259]) );
  XOR U1650 ( .A(B[259]), .B(A[259]), .Z(n1650) );
  XOR U1651 ( .A(n1651), .B(n1652), .Z(DIFF[258]) );
  XOR U1652 ( .A(B[258]), .B(A[258]), .Z(n1652) );
  XOR U1653 ( .A(n1653), .B(n1654), .Z(DIFF[257]) );
  XOR U1654 ( .A(B[257]), .B(A[257]), .Z(n1654) );
  XOR U1655 ( .A(n1655), .B(n1656), .Z(DIFF[256]) );
  XOR U1656 ( .A(B[256]), .B(A[256]), .Z(n1656) );
  XOR U1657 ( .A(n1657), .B(n1658), .Z(DIFF[255]) );
  XOR U1658 ( .A(B[255]), .B(A[255]), .Z(n1658) );
  XOR U1659 ( .A(n1659), .B(n1660), .Z(DIFF[254]) );
  XOR U1660 ( .A(B[254]), .B(A[254]), .Z(n1660) );
  XOR U1661 ( .A(n1661), .B(n1662), .Z(DIFF[253]) );
  XOR U1662 ( .A(B[253]), .B(A[253]), .Z(n1662) );
  XOR U1663 ( .A(n1663), .B(n1664), .Z(DIFF[252]) );
  XOR U1664 ( .A(B[252]), .B(A[252]), .Z(n1664) );
  XOR U1665 ( .A(n1665), .B(n1666), .Z(DIFF[251]) );
  XOR U1666 ( .A(B[251]), .B(A[251]), .Z(n1666) );
  XOR U1667 ( .A(n1667), .B(n1668), .Z(DIFF[250]) );
  XOR U1668 ( .A(B[250]), .B(A[250]), .Z(n1668) );
  XOR U1669 ( .A(n1669), .B(n1670), .Z(DIFF[24]) );
  XOR U1670 ( .A(B[24]), .B(A[24]), .Z(n1670) );
  XOR U1671 ( .A(n1671), .B(n1672), .Z(DIFF[249]) );
  XOR U1672 ( .A(B[249]), .B(A[249]), .Z(n1672) );
  XOR U1673 ( .A(n1673), .B(n1674), .Z(DIFF[248]) );
  XOR U1674 ( .A(B[248]), .B(A[248]), .Z(n1674) );
  XOR U1675 ( .A(n1675), .B(n1676), .Z(DIFF[247]) );
  XOR U1676 ( .A(B[247]), .B(A[247]), .Z(n1676) );
  XOR U1677 ( .A(n1677), .B(n1678), .Z(DIFF[246]) );
  XOR U1678 ( .A(B[246]), .B(A[246]), .Z(n1678) );
  XOR U1679 ( .A(n1679), .B(n1680), .Z(DIFF[245]) );
  XOR U1680 ( .A(B[245]), .B(A[245]), .Z(n1680) );
  XOR U1681 ( .A(n1681), .B(n1682), .Z(DIFF[244]) );
  XOR U1682 ( .A(B[244]), .B(A[244]), .Z(n1682) );
  XOR U1683 ( .A(n1683), .B(n1684), .Z(DIFF[243]) );
  XOR U1684 ( .A(B[243]), .B(A[243]), .Z(n1684) );
  XOR U1685 ( .A(n1685), .B(n1686), .Z(DIFF[242]) );
  XOR U1686 ( .A(B[242]), .B(A[242]), .Z(n1686) );
  XOR U1687 ( .A(n1687), .B(n1688), .Z(DIFF[241]) );
  XOR U1688 ( .A(B[241]), .B(A[241]), .Z(n1688) );
  XOR U1689 ( .A(n1689), .B(n1690), .Z(DIFF[240]) );
  XOR U1690 ( .A(B[240]), .B(A[240]), .Z(n1690) );
  XOR U1691 ( .A(n1691), .B(n1692), .Z(DIFF[23]) );
  XOR U1692 ( .A(B[23]), .B(A[23]), .Z(n1692) );
  XOR U1693 ( .A(n1693), .B(n1694), .Z(DIFF[239]) );
  XOR U1694 ( .A(B[239]), .B(A[239]), .Z(n1694) );
  XOR U1695 ( .A(n1695), .B(n1696), .Z(DIFF[238]) );
  XOR U1696 ( .A(B[238]), .B(A[238]), .Z(n1696) );
  XOR U1697 ( .A(n1697), .B(n1698), .Z(DIFF[237]) );
  XOR U1698 ( .A(B[237]), .B(A[237]), .Z(n1698) );
  XOR U1699 ( .A(n1699), .B(n1700), .Z(DIFF[236]) );
  XOR U1700 ( .A(B[236]), .B(A[236]), .Z(n1700) );
  XOR U1701 ( .A(n1701), .B(n1702), .Z(DIFF[235]) );
  XOR U1702 ( .A(B[235]), .B(A[235]), .Z(n1702) );
  XOR U1703 ( .A(n1703), .B(n1704), .Z(DIFF[234]) );
  XOR U1704 ( .A(B[234]), .B(A[234]), .Z(n1704) );
  XOR U1705 ( .A(n1705), .B(n1706), .Z(DIFF[233]) );
  XOR U1706 ( .A(B[233]), .B(A[233]), .Z(n1706) );
  XOR U1707 ( .A(n1707), .B(n1708), .Z(DIFF[232]) );
  XOR U1708 ( .A(B[232]), .B(A[232]), .Z(n1708) );
  XOR U1709 ( .A(n1709), .B(n1710), .Z(DIFF[231]) );
  XOR U1710 ( .A(B[231]), .B(A[231]), .Z(n1710) );
  XOR U1711 ( .A(n1711), .B(n1712), .Z(DIFF[230]) );
  XOR U1712 ( .A(B[230]), .B(A[230]), .Z(n1712) );
  XOR U1713 ( .A(n1713), .B(n1714), .Z(DIFF[22]) );
  XOR U1714 ( .A(B[22]), .B(A[22]), .Z(n1714) );
  XOR U1715 ( .A(n1715), .B(n1716), .Z(DIFF[229]) );
  XOR U1716 ( .A(B[229]), .B(A[229]), .Z(n1716) );
  XOR U1717 ( .A(n1717), .B(n1718), .Z(DIFF[228]) );
  XOR U1718 ( .A(B[228]), .B(A[228]), .Z(n1718) );
  XOR U1719 ( .A(n1719), .B(n1720), .Z(DIFF[227]) );
  XOR U1720 ( .A(B[227]), .B(A[227]), .Z(n1720) );
  XOR U1721 ( .A(n1721), .B(n1722), .Z(DIFF[226]) );
  XOR U1722 ( .A(B[226]), .B(A[226]), .Z(n1722) );
  XOR U1723 ( .A(n1723), .B(n1724), .Z(DIFF[225]) );
  XOR U1724 ( .A(B[225]), .B(A[225]), .Z(n1724) );
  XOR U1725 ( .A(n1725), .B(n1726), .Z(DIFF[224]) );
  XOR U1726 ( .A(B[224]), .B(A[224]), .Z(n1726) );
  XOR U1727 ( .A(n1727), .B(n1728), .Z(DIFF[223]) );
  XOR U1728 ( .A(B[223]), .B(A[223]), .Z(n1728) );
  XOR U1729 ( .A(n1729), .B(n1730), .Z(DIFF[222]) );
  XOR U1730 ( .A(B[222]), .B(A[222]), .Z(n1730) );
  XOR U1731 ( .A(n1731), .B(n1732), .Z(DIFF[221]) );
  XOR U1732 ( .A(B[221]), .B(A[221]), .Z(n1732) );
  XOR U1733 ( .A(n1733), .B(n1734), .Z(DIFF[220]) );
  XOR U1734 ( .A(B[220]), .B(A[220]), .Z(n1734) );
  XOR U1735 ( .A(n1735), .B(n1736), .Z(DIFF[21]) );
  XOR U1736 ( .A(B[21]), .B(A[21]), .Z(n1736) );
  XOR U1737 ( .A(n1737), .B(n1738), .Z(DIFF[219]) );
  XOR U1738 ( .A(B[219]), .B(A[219]), .Z(n1738) );
  XOR U1739 ( .A(n1739), .B(n1740), .Z(DIFF[218]) );
  XOR U1740 ( .A(B[218]), .B(A[218]), .Z(n1740) );
  XOR U1741 ( .A(n1741), .B(n1742), .Z(DIFF[217]) );
  XOR U1742 ( .A(B[217]), .B(A[217]), .Z(n1742) );
  XOR U1743 ( .A(n1743), .B(n1744), .Z(DIFF[216]) );
  XOR U1744 ( .A(B[216]), .B(A[216]), .Z(n1744) );
  XOR U1745 ( .A(n1745), .B(n1746), .Z(DIFF[215]) );
  XOR U1746 ( .A(B[215]), .B(A[215]), .Z(n1746) );
  XOR U1747 ( .A(n1747), .B(n1748), .Z(DIFF[214]) );
  XOR U1748 ( .A(B[214]), .B(A[214]), .Z(n1748) );
  XOR U1749 ( .A(n1749), .B(n1750), .Z(DIFF[213]) );
  XOR U1750 ( .A(B[213]), .B(A[213]), .Z(n1750) );
  XOR U1751 ( .A(n1751), .B(n1752), .Z(DIFF[212]) );
  XOR U1752 ( .A(B[212]), .B(A[212]), .Z(n1752) );
  XOR U1753 ( .A(n1753), .B(n1754), .Z(DIFF[211]) );
  XOR U1754 ( .A(B[211]), .B(A[211]), .Z(n1754) );
  XOR U1755 ( .A(n1755), .B(n1756), .Z(DIFF[210]) );
  XOR U1756 ( .A(B[210]), .B(A[210]), .Z(n1756) );
  XOR U1757 ( .A(n1757), .B(n1758), .Z(DIFF[20]) );
  XOR U1758 ( .A(B[20]), .B(A[20]), .Z(n1758) );
  XOR U1759 ( .A(n1759), .B(n1760), .Z(DIFF[209]) );
  XOR U1760 ( .A(B[209]), .B(A[209]), .Z(n1760) );
  XOR U1761 ( .A(n1761), .B(n1762), .Z(DIFF[208]) );
  XOR U1762 ( .A(B[208]), .B(A[208]), .Z(n1762) );
  XOR U1763 ( .A(n1763), .B(n1764), .Z(DIFF[207]) );
  XOR U1764 ( .A(B[207]), .B(A[207]), .Z(n1764) );
  XOR U1765 ( .A(n1765), .B(n1766), .Z(DIFF[206]) );
  XOR U1766 ( .A(B[206]), .B(A[206]), .Z(n1766) );
  XOR U1767 ( .A(n1767), .B(n1768), .Z(DIFF[205]) );
  XOR U1768 ( .A(B[205]), .B(A[205]), .Z(n1768) );
  XOR U1769 ( .A(n1769), .B(n1770), .Z(DIFF[204]) );
  XOR U1770 ( .A(B[204]), .B(A[204]), .Z(n1770) );
  XOR U1771 ( .A(n1771), .B(n1772), .Z(DIFF[203]) );
  XOR U1772 ( .A(B[203]), .B(A[203]), .Z(n1772) );
  XOR U1773 ( .A(n1773), .B(n1774), .Z(DIFF[202]) );
  XOR U1774 ( .A(B[202]), .B(A[202]), .Z(n1774) );
  XOR U1775 ( .A(n1775), .B(n1776), .Z(DIFF[201]) );
  XOR U1776 ( .A(B[201]), .B(A[201]), .Z(n1776) );
  XOR U1777 ( .A(n1777), .B(n1778), .Z(DIFF[200]) );
  XOR U1778 ( .A(B[200]), .B(A[200]), .Z(n1778) );
  XOR U1779 ( .A(n1), .B(n1779), .Z(DIFF[1]) );
  XOR U1780 ( .A(B[1]), .B(A[1]), .Z(n1779) );
  XOR U1781 ( .A(n1780), .B(n1781), .Z(DIFF[19]) );
  XOR U1782 ( .A(B[19]), .B(A[19]), .Z(n1781) );
  XOR U1783 ( .A(n1782), .B(n1783), .Z(DIFF[199]) );
  XOR U1784 ( .A(B[199]), .B(A[199]), .Z(n1783) );
  XOR U1785 ( .A(n1784), .B(n1785), .Z(DIFF[198]) );
  XOR U1786 ( .A(B[198]), .B(A[198]), .Z(n1785) );
  XOR U1787 ( .A(n1786), .B(n1787), .Z(DIFF[197]) );
  XOR U1788 ( .A(B[197]), .B(A[197]), .Z(n1787) );
  XOR U1789 ( .A(n1788), .B(n1789), .Z(DIFF[196]) );
  XOR U1790 ( .A(B[196]), .B(A[196]), .Z(n1789) );
  XOR U1791 ( .A(n1790), .B(n1791), .Z(DIFF[195]) );
  XOR U1792 ( .A(B[195]), .B(A[195]), .Z(n1791) );
  XOR U1793 ( .A(n1792), .B(n1793), .Z(DIFF[194]) );
  XOR U1794 ( .A(B[194]), .B(A[194]), .Z(n1793) );
  XOR U1795 ( .A(n1794), .B(n1795), .Z(DIFF[193]) );
  XOR U1796 ( .A(B[193]), .B(A[193]), .Z(n1795) );
  XOR U1797 ( .A(n1796), .B(n1797), .Z(DIFF[192]) );
  XOR U1798 ( .A(B[192]), .B(A[192]), .Z(n1797) );
  XOR U1799 ( .A(n1798), .B(n1799), .Z(DIFF[191]) );
  XOR U1800 ( .A(B[191]), .B(A[191]), .Z(n1799) );
  XOR U1801 ( .A(n1800), .B(n1801), .Z(DIFF[190]) );
  XOR U1802 ( .A(B[190]), .B(A[190]), .Z(n1801) );
  XOR U1803 ( .A(n1802), .B(n1803), .Z(DIFF[18]) );
  XOR U1804 ( .A(B[18]), .B(A[18]), .Z(n1803) );
  XOR U1805 ( .A(n1804), .B(n1805), .Z(DIFF[189]) );
  XOR U1806 ( .A(B[189]), .B(A[189]), .Z(n1805) );
  XOR U1807 ( .A(n1806), .B(n1807), .Z(DIFF[188]) );
  XOR U1808 ( .A(B[188]), .B(A[188]), .Z(n1807) );
  XOR U1809 ( .A(n1808), .B(n1809), .Z(DIFF[187]) );
  XOR U1810 ( .A(B[187]), .B(A[187]), .Z(n1809) );
  XOR U1811 ( .A(n1810), .B(n1811), .Z(DIFF[186]) );
  XOR U1812 ( .A(B[186]), .B(A[186]), .Z(n1811) );
  XOR U1813 ( .A(n1812), .B(n1813), .Z(DIFF[185]) );
  XOR U1814 ( .A(B[185]), .B(A[185]), .Z(n1813) );
  XOR U1815 ( .A(n1814), .B(n1815), .Z(DIFF[184]) );
  XOR U1816 ( .A(B[184]), .B(A[184]), .Z(n1815) );
  XOR U1817 ( .A(n1816), .B(n1817), .Z(DIFF[183]) );
  XOR U1818 ( .A(B[183]), .B(A[183]), .Z(n1817) );
  XOR U1819 ( .A(n1818), .B(n1819), .Z(DIFF[182]) );
  XOR U1820 ( .A(B[182]), .B(A[182]), .Z(n1819) );
  XOR U1821 ( .A(n1820), .B(n1821), .Z(DIFF[181]) );
  XOR U1822 ( .A(B[181]), .B(A[181]), .Z(n1821) );
  XOR U1823 ( .A(n1822), .B(n1823), .Z(DIFF[180]) );
  XOR U1824 ( .A(B[180]), .B(A[180]), .Z(n1823) );
  XOR U1825 ( .A(n1824), .B(n1825), .Z(DIFF[17]) );
  XOR U1826 ( .A(B[17]), .B(A[17]), .Z(n1825) );
  XOR U1827 ( .A(n1826), .B(n1827), .Z(DIFF[179]) );
  XOR U1828 ( .A(B[179]), .B(A[179]), .Z(n1827) );
  XOR U1829 ( .A(n1828), .B(n1829), .Z(DIFF[178]) );
  XOR U1830 ( .A(B[178]), .B(A[178]), .Z(n1829) );
  XOR U1831 ( .A(n1830), .B(n1831), .Z(DIFF[177]) );
  XOR U1832 ( .A(B[177]), .B(A[177]), .Z(n1831) );
  XOR U1833 ( .A(n1832), .B(n1833), .Z(DIFF[176]) );
  XOR U1834 ( .A(B[176]), .B(A[176]), .Z(n1833) );
  XOR U1835 ( .A(n1834), .B(n1835), .Z(DIFF[175]) );
  XOR U1836 ( .A(B[175]), .B(A[175]), .Z(n1835) );
  XOR U1837 ( .A(n1836), .B(n1837), .Z(DIFF[174]) );
  XOR U1838 ( .A(B[174]), .B(A[174]), .Z(n1837) );
  XOR U1839 ( .A(n1838), .B(n1839), .Z(DIFF[173]) );
  XOR U1840 ( .A(B[173]), .B(A[173]), .Z(n1839) );
  XOR U1841 ( .A(n1840), .B(n1841), .Z(DIFF[172]) );
  XOR U1842 ( .A(B[172]), .B(A[172]), .Z(n1841) );
  XOR U1843 ( .A(n1842), .B(n1843), .Z(DIFF[171]) );
  XOR U1844 ( .A(B[171]), .B(A[171]), .Z(n1843) );
  XOR U1845 ( .A(n1844), .B(n1845), .Z(DIFF[170]) );
  XOR U1846 ( .A(B[170]), .B(A[170]), .Z(n1845) );
  XOR U1847 ( .A(n1846), .B(n1847), .Z(DIFF[16]) );
  XOR U1848 ( .A(B[16]), .B(A[16]), .Z(n1847) );
  XOR U1849 ( .A(n1848), .B(n1849), .Z(DIFF[169]) );
  XOR U1850 ( .A(B[169]), .B(A[169]), .Z(n1849) );
  XOR U1851 ( .A(n1850), .B(n1851), .Z(DIFF[168]) );
  XOR U1852 ( .A(B[168]), .B(A[168]), .Z(n1851) );
  XOR U1853 ( .A(n1852), .B(n1853), .Z(DIFF[167]) );
  XOR U1854 ( .A(B[167]), .B(A[167]), .Z(n1853) );
  XOR U1855 ( .A(n1854), .B(n1855), .Z(DIFF[166]) );
  XOR U1856 ( .A(B[166]), .B(A[166]), .Z(n1855) );
  XOR U1857 ( .A(n1856), .B(n1857), .Z(DIFF[165]) );
  XOR U1858 ( .A(B[165]), .B(A[165]), .Z(n1857) );
  XOR U1859 ( .A(n1858), .B(n1859), .Z(DIFF[164]) );
  XOR U1860 ( .A(B[164]), .B(A[164]), .Z(n1859) );
  XOR U1861 ( .A(n1860), .B(n1861), .Z(DIFF[163]) );
  XOR U1862 ( .A(B[163]), .B(A[163]), .Z(n1861) );
  XOR U1863 ( .A(n1862), .B(n1863), .Z(DIFF[162]) );
  XOR U1864 ( .A(B[162]), .B(A[162]), .Z(n1863) );
  XOR U1865 ( .A(n1864), .B(n1865), .Z(DIFF[161]) );
  XOR U1866 ( .A(B[161]), .B(A[161]), .Z(n1865) );
  XOR U1867 ( .A(n1866), .B(n1867), .Z(DIFF[160]) );
  XOR U1868 ( .A(B[160]), .B(A[160]), .Z(n1867) );
  XOR U1869 ( .A(n1868), .B(n1869), .Z(DIFF[15]) );
  XOR U1870 ( .A(B[15]), .B(A[15]), .Z(n1869) );
  XOR U1871 ( .A(n1870), .B(n1871), .Z(DIFF[159]) );
  XOR U1872 ( .A(B[159]), .B(A[159]), .Z(n1871) );
  XOR U1873 ( .A(n1872), .B(n1873), .Z(DIFF[158]) );
  XOR U1874 ( .A(B[158]), .B(A[158]), .Z(n1873) );
  XOR U1875 ( .A(n1874), .B(n1875), .Z(DIFF[157]) );
  XOR U1876 ( .A(B[157]), .B(A[157]), .Z(n1875) );
  XOR U1877 ( .A(n1876), .B(n1877), .Z(DIFF[156]) );
  XOR U1878 ( .A(B[156]), .B(A[156]), .Z(n1877) );
  XOR U1879 ( .A(n1878), .B(n1879), .Z(DIFF[155]) );
  XOR U1880 ( .A(B[155]), .B(A[155]), .Z(n1879) );
  XOR U1881 ( .A(n1880), .B(n1881), .Z(DIFF[154]) );
  XOR U1882 ( .A(B[154]), .B(A[154]), .Z(n1881) );
  XOR U1883 ( .A(n1882), .B(n1883), .Z(DIFF[153]) );
  XOR U1884 ( .A(B[153]), .B(A[153]), .Z(n1883) );
  XOR U1885 ( .A(n1884), .B(n1885), .Z(DIFF[152]) );
  XOR U1886 ( .A(B[152]), .B(A[152]), .Z(n1885) );
  XOR U1887 ( .A(n1886), .B(n1887), .Z(DIFF[151]) );
  XOR U1888 ( .A(B[151]), .B(A[151]), .Z(n1887) );
  XOR U1889 ( .A(n1888), .B(n1889), .Z(DIFF[150]) );
  XOR U1890 ( .A(B[150]), .B(A[150]), .Z(n1889) );
  XOR U1891 ( .A(n1890), .B(n1891), .Z(DIFF[14]) );
  XOR U1892 ( .A(B[14]), .B(A[14]), .Z(n1891) );
  XOR U1893 ( .A(n1892), .B(n1893), .Z(DIFF[149]) );
  XOR U1894 ( .A(B[149]), .B(A[149]), .Z(n1893) );
  XOR U1895 ( .A(n1894), .B(n1895), .Z(DIFF[148]) );
  XOR U1896 ( .A(B[148]), .B(A[148]), .Z(n1895) );
  XOR U1897 ( .A(n1896), .B(n1897), .Z(DIFF[147]) );
  XOR U1898 ( .A(B[147]), .B(A[147]), .Z(n1897) );
  XOR U1899 ( .A(n1898), .B(n1899), .Z(DIFF[146]) );
  XOR U1900 ( .A(B[146]), .B(A[146]), .Z(n1899) );
  XOR U1901 ( .A(n1900), .B(n1901), .Z(DIFF[145]) );
  XOR U1902 ( .A(B[145]), .B(A[145]), .Z(n1901) );
  XOR U1903 ( .A(n1902), .B(n1903), .Z(DIFF[144]) );
  XOR U1904 ( .A(B[144]), .B(A[144]), .Z(n1903) );
  XOR U1905 ( .A(n1904), .B(n1905), .Z(DIFF[143]) );
  XOR U1906 ( .A(B[143]), .B(A[143]), .Z(n1905) );
  XOR U1907 ( .A(n1906), .B(n1907), .Z(DIFF[142]) );
  XOR U1908 ( .A(B[142]), .B(A[142]), .Z(n1907) );
  XOR U1909 ( .A(n1908), .B(n1909), .Z(DIFF[141]) );
  XOR U1910 ( .A(B[141]), .B(A[141]), .Z(n1909) );
  XOR U1911 ( .A(n1910), .B(n1911), .Z(DIFF[140]) );
  XOR U1912 ( .A(B[140]), .B(A[140]), .Z(n1911) );
  XOR U1913 ( .A(n1912), .B(n1913), .Z(DIFF[13]) );
  XOR U1914 ( .A(B[13]), .B(A[13]), .Z(n1913) );
  XOR U1915 ( .A(n1914), .B(n1915), .Z(DIFF[139]) );
  XOR U1916 ( .A(B[139]), .B(A[139]), .Z(n1915) );
  XOR U1917 ( .A(n1916), .B(n1917), .Z(DIFF[138]) );
  XOR U1918 ( .A(B[138]), .B(A[138]), .Z(n1917) );
  XOR U1919 ( .A(n1918), .B(n1919), .Z(DIFF[137]) );
  XOR U1920 ( .A(B[137]), .B(A[137]), .Z(n1919) );
  XOR U1921 ( .A(n1920), .B(n1921), .Z(DIFF[136]) );
  XOR U1922 ( .A(B[136]), .B(A[136]), .Z(n1921) );
  XOR U1923 ( .A(n1922), .B(n1923), .Z(DIFF[135]) );
  XOR U1924 ( .A(B[135]), .B(A[135]), .Z(n1923) );
  XOR U1925 ( .A(n1924), .B(n1925), .Z(DIFF[134]) );
  XOR U1926 ( .A(B[134]), .B(A[134]), .Z(n1925) );
  XOR U1927 ( .A(n1926), .B(n1927), .Z(DIFF[133]) );
  XOR U1928 ( .A(B[133]), .B(A[133]), .Z(n1927) );
  XOR U1929 ( .A(n1928), .B(n1929), .Z(DIFF[132]) );
  XOR U1930 ( .A(B[132]), .B(A[132]), .Z(n1929) );
  XOR U1931 ( .A(n1930), .B(n1931), .Z(DIFF[131]) );
  XOR U1932 ( .A(B[131]), .B(A[131]), .Z(n1931) );
  XOR U1933 ( .A(n1932), .B(n1933), .Z(DIFF[130]) );
  XOR U1934 ( .A(B[130]), .B(A[130]), .Z(n1933) );
  XOR U1935 ( .A(n1934), .B(n1935), .Z(DIFF[12]) );
  XOR U1936 ( .A(B[12]), .B(A[12]), .Z(n1935) );
  XOR U1937 ( .A(n1936), .B(n1937), .Z(DIFF[129]) );
  XOR U1938 ( .A(B[129]), .B(A[129]), .Z(n1937) );
  XOR U1939 ( .A(n1938), .B(n1939), .Z(DIFF[128]) );
  XOR U1940 ( .A(B[128]), .B(A[128]), .Z(n1939) );
  XOR U1941 ( .A(n1940), .B(n1941), .Z(DIFF[127]) );
  XOR U1942 ( .A(B[127]), .B(A[127]), .Z(n1941) );
  XOR U1943 ( .A(n1942), .B(n1943), .Z(DIFF[126]) );
  XOR U1944 ( .A(B[126]), .B(A[126]), .Z(n1943) );
  XOR U1945 ( .A(n1944), .B(n1945), .Z(DIFF[125]) );
  XOR U1946 ( .A(B[125]), .B(A[125]), .Z(n1945) );
  XOR U1947 ( .A(n1946), .B(n1947), .Z(DIFF[124]) );
  XOR U1948 ( .A(B[124]), .B(A[124]), .Z(n1947) );
  XOR U1949 ( .A(n1948), .B(n1949), .Z(DIFF[123]) );
  XOR U1950 ( .A(B[123]), .B(A[123]), .Z(n1949) );
  XOR U1951 ( .A(n1950), .B(n1951), .Z(DIFF[122]) );
  XOR U1952 ( .A(B[122]), .B(A[122]), .Z(n1951) );
  XOR U1953 ( .A(n1952), .B(n1953), .Z(DIFF[121]) );
  XOR U1954 ( .A(B[121]), .B(A[121]), .Z(n1953) );
  XOR U1955 ( .A(n1954), .B(n1955), .Z(DIFF[120]) );
  XOR U1956 ( .A(B[120]), .B(A[120]), .Z(n1955) );
  XOR U1957 ( .A(n1956), .B(n1957), .Z(DIFF[11]) );
  XOR U1958 ( .A(B[11]), .B(A[11]), .Z(n1957) );
  XOR U1959 ( .A(n1958), .B(n1959), .Z(DIFF[119]) );
  XOR U1960 ( .A(B[119]), .B(A[119]), .Z(n1959) );
  XOR U1961 ( .A(n1960), .B(n1961), .Z(DIFF[118]) );
  XOR U1962 ( .A(B[118]), .B(A[118]), .Z(n1961) );
  XOR U1963 ( .A(n1962), .B(n1963), .Z(DIFF[117]) );
  XOR U1964 ( .A(B[117]), .B(A[117]), .Z(n1963) );
  XOR U1965 ( .A(n1964), .B(n1965), .Z(DIFF[116]) );
  XOR U1966 ( .A(B[116]), .B(A[116]), .Z(n1965) );
  XOR U1967 ( .A(n1966), .B(n1967), .Z(DIFF[115]) );
  XOR U1968 ( .A(B[115]), .B(A[115]), .Z(n1967) );
  XOR U1969 ( .A(n1968), .B(n1969), .Z(DIFF[114]) );
  XOR U1970 ( .A(B[114]), .B(A[114]), .Z(n1969) );
  XOR U1971 ( .A(n1970), .B(n1971), .Z(DIFF[113]) );
  XOR U1972 ( .A(B[113]), .B(A[113]), .Z(n1971) );
  XOR U1973 ( .A(n1972), .B(n1973), .Z(DIFF[112]) );
  XOR U1974 ( .A(B[112]), .B(A[112]), .Z(n1973) );
  XOR U1975 ( .A(n1974), .B(n1975), .Z(DIFF[111]) );
  XOR U1976 ( .A(B[111]), .B(A[111]), .Z(n1975) );
  XOR U1977 ( .A(n1976), .B(n1977), .Z(DIFF[110]) );
  XOR U1978 ( .A(B[110]), .B(A[110]), .Z(n1977) );
  XOR U1979 ( .A(n1978), .B(n1979), .Z(DIFF[10]) );
  XOR U1980 ( .A(B[10]), .B(A[10]), .Z(n1979) );
  XOR U1981 ( .A(n1980), .B(n1981), .Z(DIFF[109]) );
  XOR U1982 ( .A(B[109]), .B(A[109]), .Z(n1981) );
  XOR U1983 ( .A(n1982), .B(n1983), .Z(DIFF[108]) );
  XOR U1984 ( .A(B[108]), .B(A[108]), .Z(n1983) );
  XOR U1985 ( .A(n1984), .B(n1985), .Z(DIFF[107]) );
  XOR U1986 ( .A(B[107]), .B(A[107]), .Z(n1985) );
  XOR U1987 ( .A(n1986), .B(n1987), .Z(DIFF[106]) );
  XOR U1988 ( .A(B[106]), .B(A[106]), .Z(n1987) );
  XOR U1989 ( .A(n1988), .B(n1989), .Z(DIFF[105]) );
  XOR U1990 ( .A(B[105]), .B(A[105]), .Z(n1989) );
  XOR U1991 ( .A(n1990), .B(n1991), .Z(DIFF[104]) );
  XOR U1992 ( .A(B[104]), .B(A[104]), .Z(n1991) );
  XOR U1993 ( .A(n1992), .B(n1993), .Z(DIFF[103]) );
  XOR U1994 ( .A(B[103]), .B(A[103]), .Z(n1993) );
  XOR U1995 ( .A(n1994), .B(n1995), .Z(DIFF[102]) );
  XOR U1996 ( .A(B[102]), .B(A[102]), .Z(n1995) );
  XOR U1997 ( .A(A[1025]), .B(n1996), .Z(DIFF[1025]) );
  ANDN U1998 ( .B(n1997), .A(A[1024]), .Z(n1996) );
  XOR U1999 ( .A(A[1024]), .B(n1997), .Z(DIFF[1024]) );
  AND U2000 ( .A(n1998), .B(n1999), .Z(n1997) );
  NANDN U2001 ( .A(B[1023]), .B(n2000), .Z(n1999) );
  NANDN U2002 ( .A(A[1023]), .B(n2001), .Z(n2000) );
  NANDN U2003 ( .A(n2001), .B(A[1023]), .Z(n1998) );
  XOR U2004 ( .A(n2001), .B(n2002), .Z(DIFF[1023]) );
  XOR U2005 ( .A(B[1023]), .B(A[1023]), .Z(n2002) );
  AND U2006 ( .A(n2003), .B(n2004), .Z(n2001) );
  NANDN U2007 ( .A(B[1022]), .B(n2005), .Z(n2004) );
  NANDN U2008 ( .A(A[1022]), .B(n2006), .Z(n2005) );
  NANDN U2009 ( .A(n2006), .B(A[1022]), .Z(n2003) );
  XOR U2010 ( .A(n2006), .B(n2007), .Z(DIFF[1022]) );
  XOR U2011 ( .A(B[1022]), .B(A[1022]), .Z(n2007) );
  AND U2012 ( .A(n2008), .B(n2009), .Z(n2006) );
  NANDN U2013 ( .A(B[1021]), .B(n2010), .Z(n2009) );
  NANDN U2014 ( .A(A[1021]), .B(n2011), .Z(n2010) );
  NANDN U2015 ( .A(n2011), .B(A[1021]), .Z(n2008) );
  XOR U2016 ( .A(n2011), .B(n2012), .Z(DIFF[1021]) );
  XOR U2017 ( .A(B[1021]), .B(A[1021]), .Z(n2012) );
  AND U2018 ( .A(n2013), .B(n2014), .Z(n2011) );
  NANDN U2019 ( .A(B[1020]), .B(n2015), .Z(n2014) );
  NANDN U2020 ( .A(A[1020]), .B(n2016), .Z(n2015) );
  NANDN U2021 ( .A(n2016), .B(A[1020]), .Z(n2013) );
  XOR U2022 ( .A(n2016), .B(n2017), .Z(DIFF[1020]) );
  XOR U2023 ( .A(B[1020]), .B(A[1020]), .Z(n2017) );
  AND U2024 ( .A(n2018), .B(n2019), .Z(n2016) );
  NANDN U2025 ( .A(B[1019]), .B(n2020), .Z(n2019) );
  NANDN U2026 ( .A(A[1019]), .B(n2021), .Z(n2020) );
  NANDN U2027 ( .A(n2021), .B(A[1019]), .Z(n2018) );
  XOR U2028 ( .A(n2022), .B(n2023), .Z(DIFF[101]) );
  XOR U2029 ( .A(B[101]), .B(A[101]), .Z(n2023) );
  XOR U2030 ( .A(n2021), .B(n2024), .Z(DIFF[1019]) );
  XOR U2031 ( .A(B[1019]), .B(A[1019]), .Z(n2024) );
  AND U2032 ( .A(n2025), .B(n2026), .Z(n2021) );
  NANDN U2033 ( .A(B[1018]), .B(n2027), .Z(n2026) );
  NANDN U2034 ( .A(A[1018]), .B(n2028), .Z(n2027) );
  NANDN U2035 ( .A(n2028), .B(A[1018]), .Z(n2025) );
  XOR U2036 ( .A(n2028), .B(n2029), .Z(DIFF[1018]) );
  XOR U2037 ( .A(B[1018]), .B(A[1018]), .Z(n2029) );
  AND U2038 ( .A(n2030), .B(n2031), .Z(n2028) );
  NANDN U2039 ( .A(B[1017]), .B(n2032), .Z(n2031) );
  NANDN U2040 ( .A(A[1017]), .B(n2033), .Z(n2032) );
  NANDN U2041 ( .A(n2033), .B(A[1017]), .Z(n2030) );
  XOR U2042 ( .A(n2033), .B(n2034), .Z(DIFF[1017]) );
  XOR U2043 ( .A(B[1017]), .B(A[1017]), .Z(n2034) );
  AND U2044 ( .A(n2035), .B(n2036), .Z(n2033) );
  NANDN U2045 ( .A(B[1016]), .B(n2037), .Z(n2036) );
  NANDN U2046 ( .A(A[1016]), .B(n2038), .Z(n2037) );
  NANDN U2047 ( .A(n2038), .B(A[1016]), .Z(n2035) );
  XOR U2048 ( .A(n2038), .B(n2039), .Z(DIFF[1016]) );
  XOR U2049 ( .A(B[1016]), .B(A[1016]), .Z(n2039) );
  AND U2050 ( .A(n2040), .B(n2041), .Z(n2038) );
  NANDN U2051 ( .A(B[1015]), .B(n2042), .Z(n2041) );
  NANDN U2052 ( .A(A[1015]), .B(n2043), .Z(n2042) );
  NANDN U2053 ( .A(n2043), .B(A[1015]), .Z(n2040) );
  XOR U2054 ( .A(n2043), .B(n2044), .Z(DIFF[1015]) );
  XOR U2055 ( .A(B[1015]), .B(A[1015]), .Z(n2044) );
  AND U2056 ( .A(n2045), .B(n2046), .Z(n2043) );
  NANDN U2057 ( .A(B[1014]), .B(n2047), .Z(n2046) );
  NANDN U2058 ( .A(A[1014]), .B(n2048), .Z(n2047) );
  NANDN U2059 ( .A(n2048), .B(A[1014]), .Z(n2045) );
  XOR U2060 ( .A(n2048), .B(n2049), .Z(DIFF[1014]) );
  XOR U2061 ( .A(B[1014]), .B(A[1014]), .Z(n2049) );
  AND U2062 ( .A(n2050), .B(n2051), .Z(n2048) );
  NANDN U2063 ( .A(B[1013]), .B(n2052), .Z(n2051) );
  NANDN U2064 ( .A(A[1013]), .B(n2053), .Z(n2052) );
  NANDN U2065 ( .A(n2053), .B(A[1013]), .Z(n2050) );
  XOR U2066 ( .A(n2053), .B(n2054), .Z(DIFF[1013]) );
  XOR U2067 ( .A(B[1013]), .B(A[1013]), .Z(n2054) );
  AND U2068 ( .A(n2055), .B(n2056), .Z(n2053) );
  NANDN U2069 ( .A(B[1012]), .B(n2057), .Z(n2056) );
  NANDN U2070 ( .A(A[1012]), .B(n2058), .Z(n2057) );
  NANDN U2071 ( .A(n2058), .B(A[1012]), .Z(n2055) );
  XOR U2072 ( .A(n2058), .B(n2059), .Z(DIFF[1012]) );
  XOR U2073 ( .A(B[1012]), .B(A[1012]), .Z(n2059) );
  AND U2074 ( .A(n2060), .B(n2061), .Z(n2058) );
  NANDN U2075 ( .A(B[1011]), .B(n2062), .Z(n2061) );
  NANDN U2076 ( .A(A[1011]), .B(n2063), .Z(n2062) );
  NANDN U2077 ( .A(n2063), .B(A[1011]), .Z(n2060) );
  XOR U2078 ( .A(n2063), .B(n2064), .Z(DIFF[1011]) );
  XOR U2079 ( .A(B[1011]), .B(A[1011]), .Z(n2064) );
  AND U2080 ( .A(n2065), .B(n2066), .Z(n2063) );
  NANDN U2081 ( .A(B[1010]), .B(n2067), .Z(n2066) );
  NANDN U2082 ( .A(A[1010]), .B(n2068), .Z(n2067) );
  NANDN U2083 ( .A(n2068), .B(A[1010]), .Z(n2065) );
  XOR U2084 ( .A(n2068), .B(n2069), .Z(DIFF[1010]) );
  XOR U2085 ( .A(B[1010]), .B(A[1010]), .Z(n2069) );
  AND U2086 ( .A(n2070), .B(n2071), .Z(n2068) );
  NANDN U2087 ( .A(B[1009]), .B(n2072), .Z(n2071) );
  NANDN U2088 ( .A(A[1009]), .B(n2073), .Z(n2072) );
  NANDN U2089 ( .A(n2073), .B(A[1009]), .Z(n2070) );
  XOR U2090 ( .A(n2074), .B(n2075), .Z(DIFF[100]) );
  XOR U2091 ( .A(B[100]), .B(A[100]), .Z(n2075) );
  XOR U2092 ( .A(n2073), .B(n2076), .Z(DIFF[1009]) );
  XOR U2093 ( .A(B[1009]), .B(A[1009]), .Z(n2076) );
  AND U2094 ( .A(n2077), .B(n2078), .Z(n2073) );
  NANDN U2095 ( .A(B[1008]), .B(n2079), .Z(n2078) );
  NANDN U2096 ( .A(A[1008]), .B(n2080), .Z(n2079) );
  NANDN U2097 ( .A(n2080), .B(A[1008]), .Z(n2077) );
  XOR U2098 ( .A(n2080), .B(n2081), .Z(DIFF[1008]) );
  XOR U2099 ( .A(B[1008]), .B(A[1008]), .Z(n2081) );
  AND U2100 ( .A(n2082), .B(n2083), .Z(n2080) );
  NANDN U2101 ( .A(B[1007]), .B(n2084), .Z(n2083) );
  NANDN U2102 ( .A(A[1007]), .B(n2085), .Z(n2084) );
  NANDN U2103 ( .A(n2085), .B(A[1007]), .Z(n2082) );
  XOR U2104 ( .A(n2085), .B(n2086), .Z(DIFF[1007]) );
  XOR U2105 ( .A(B[1007]), .B(A[1007]), .Z(n2086) );
  AND U2106 ( .A(n2087), .B(n2088), .Z(n2085) );
  NANDN U2107 ( .A(B[1006]), .B(n2089), .Z(n2088) );
  NANDN U2108 ( .A(A[1006]), .B(n2090), .Z(n2089) );
  NANDN U2109 ( .A(n2090), .B(A[1006]), .Z(n2087) );
  XOR U2110 ( .A(n2090), .B(n2091), .Z(DIFF[1006]) );
  XOR U2111 ( .A(B[1006]), .B(A[1006]), .Z(n2091) );
  AND U2112 ( .A(n2092), .B(n2093), .Z(n2090) );
  NANDN U2113 ( .A(B[1005]), .B(n2094), .Z(n2093) );
  NANDN U2114 ( .A(A[1005]), .B(n2095), .Z(n2094) );
  NANDN U2115 ( .A(n2095), .B(A[1005]), .Z(n2092) );
  XOR U2116 ( .A(n2095), .B(n2096), .Z(DIFF[1005]) );
  XOR U2117 ( .A(B[1005]), .B(A[1005]), .Z(n2096) );
  AND U2118 ( .A(n2097), .B(n2098), .Z(n2095) );
  NANDN U2119 ( .A(B[1004]), .B(n2099), .Z(n2098) );
  NANDN U2120 ( .A(A[1004]), .B(n2100), .Z(n2099) );
  NANDN U2121 ( .A(n2100), .B(A[1004]), .Z(n2097) );
  XOR U2122 ( .A(n2100), .B(n2101), .Z(DIFF[1004]) );
  XOR U2123 ( .A(B[1004]), .B(A[1004]), .Z(n2101) );
  AND U2124 ( .A(n2102), .B(n2103), .Z(n2100) );
  NANDN U2125 ( .A(B[1003]), .B(n2104), .Z(n2103) );
  NANDN U2126 ( .A(A[1003]), .B(n2105), .Z(n2104) );
  NANDN U2127 ( .A(n2105), .B(A[1003]), .Z(n2102) );
  XOR U2128 ( .A(n2105), .B(n2106), .Z(DIFF[1003]) );
  XOR U2129 ( .A(B[1003]), .B(A[1003]), .Z(n2106) );
  AND U2130 ( .A(n2107), .B(n2108), .Z(n2105) );
  NANDN U2131 ( .A(B[1002]), .B(n2109), .Z(n2108) );
  NANDN U2132 ( .A(A[1002]), .B(n2110), .Z(n2109) );
  NANDN U2133 ( .A(n2110), .B(A[1002]), .Z(n2107) );
  XOR U2134 ( .A(n2110), .B(n2111), .Z(DIFF[1002]) );
  XOR U2135 ( .A(B[1002]), .B(A[1002]), .Z(n2111) );
  AND U2136 ( .A(n2112), .B(n2113), .Z(n2110) );
  NANDN U2137 ( .A(B[1001]), .B(n2114), .Z(n2113) );
  NANDN U2138 ( .A(A[1001]), .B(n2115), .Z(n2114) );
  NANDN U2139 ( .A(n2115), .B(A[1001]), .Z(n2112) );
  XOR U2140 ( .A(n2115), .B(n2116), .Z(DIFF[1001]) );
  XOR U2141 ( .A(B[1001]), .B(A[1001]), .Z(n2116) );
  AND U2142 ( .A(n2117), .B(n2118), .Z(n2115) );
  NANDN U2143 ( .A(B[1000]), .B(n2119), .Z(n2118) );
  NANDN U2144 ( .A(A[1000]), .B(n2120), .Z(n2119) );
  NANDN U2145 ( .A(n2120), .B(A[1000]), .Z(n2117) );
  XOR U2146 ( .A(n2120), .B(n2121), .Z(DIFF[1000]) );
  XOR U2147 ( .A(B[1000]), .B(A[1000]), .Z(n2121) );
  AND U2148 ( .A(n2122), .B(n2123), .Z(n2120) );
  NANDN U2149 ( .A(B[999]), .B(n2124), .Z(n2123) );
  OR U2150 ( .A(n7), .B(A[999]), .Z(n2124) );
  NAND U2151 ( .A(A[999]), .B(n7), .Z(n2122) );
  NAND U2152 ( .A(n2125), .B(n2126), .Z(n7) );
  NANDN U2153 ( .A(B[998]), .B(n2127), .Z(n2126) );
  NANDN U2154 ( .A(A[998]), .B(n9), .Z(n2127) );
  NANDN U2155 ( .A(n9), .B(A[998]), .Z(n2125) );
  AND U2156 ( .A(n2128), .B(n2129), .Z(n9) );
  NANDN U2157 ( .A(B[997]), .B(n2130), .Z(n2129) );
  NANDN U2158 ( .A(A[997]), .B(n11), .Z(n2130) );
  NANDN U2159 ( .A(n11), .B(A[997]), .Z(n2128) );
  AND U2160 ( .A(n2131), .B(n2132), .Z(n11) );
  NANDN U2161 ( .A(B[996]), .B(n2133), .Z(n2132) );
  NANDN U2162 ( .A(A[996]), .B(n13), .Z(n2133) );
  NANDN U2163 ( .A(n13), .B(A[996]), .Z(n2131) );
  AND U2164 ( .A(n2134), .B(n2135), .Z(n13) );
  NANDN U2165 ( .A(B[995]), .B(n2136), .Z(n2135) );
  NANDN U2166 ( .A(A[995]), .B(n15), .Z(n2136) );
  NANDN U2167 ( .A(n15), .B(A[995]), .Z(n2134) );
  AND U2168 ( .A(n2137), .B(n2138), .Z(n15) );
  NANDN U2169 ( .A(B[994]), .B(n2139), .Z(n2138) );
  NANDN U2170 ( .A(A[994]), .B(n17), .Z(n2139) );
  NANDN U2171 ( .A(n17), .B(A[994]), .Z(n2137) );
  AND U2172 ( .A(n2140), .B(n2141), .Z(n17) );
  NANDN U2173 ( .A(B[993]), .B(n2142), .Z(n2141) );
  NANDN U2174 ( .A(A[993]), .B(n19), .Z(n2142) );
  NANDN U2175 ( .A(n19), .B(A[993]), .Z(n2140) );
  AND U2176 ( .A(n2143), .B(n2144), .Z(n19) );
  NANDN U2177 ( .A(B[992]), .B(n2145), .Z(n2144) );
  NANDN U2178 ( .A(A[992]), .B(n21), .Z(n2145) );
  NANDN U2179 ( .A(n21), .B(A[992]), .Z(n2143) );
  AND U2180 ( .A(n2146), .B(n2147), .Z(n21) );
  NANDN U2181 ( .A(B[991]), .B(n2148), .Z(n2147) );
  NANDN U2182 ( .A(A[991]), .B(n23), .Z(n2148) );
  NANDN U2183 ( .A(n23), .B(A[991]), .Z(n2146) );
  AND U2184 ( .A(n2149), .B(n2150), .Z(n23) );
  NANDN U2185 ( .A(B[990]), .B(n2151), .Z(n2150) );
  NANDN U2186 ( .A(A[990]), .B(n25), .Z(n2151) );
  NANDN U2187 ( .A(n25), .B(A[990]), .Z(n2149) );
  AND U2188 ( .A(n2152), .B(n2153), .Z(n25) );
  NANDN U2189 ( .A(B[989]), .B(n2154), .Z(n2153) );
  NANDN U2190 ( .A(A[989]), .B(n29), .Z(n2154) );
  NANDN U2191 ( .A(n29), .B(A[989]), .Z(n2152) );
  AND U2192 ( .A(n2155), .B(n2156), .Z(n29) );
  NANDN U2193 ( .A(B[988]), .B(n2157), .Z(n2156) );
  NANDN U2194 ( .A(A[988]), .B(n31), .Z(n2157) );
  NANDN U2195 ( .A(n31), .B(A[988]), .Z(n2155) );
  AND U2196 ( .A(n2158), .B(n2159), .Z(n31) );
  NANDN U2197 ( .A(B[987]), .B(n2160), .Z(n2159) );
  NANDN U2198 ( .A(A[987]), .B(n33), .Z(n2160) );
  NANDN U2199 ( .A(n33), .B(A[987]), .Z(n2158) );
  AND U2200 ( .A(n2161), .B(n2162), .Z(n33) );
  NANDN U2201 ( .A(B[986]), .B(n2163), .Z(n2162) );
  NANDN U2202 ( .A(A[986]), .B(n35), .Z(n2163) );
  NANDN U2203 ( .A(n35), .B(A[986]), .Z(n2161) );
  AND U2204 ( .A(n2164), .B(n2165), .Z(n35) );
  NANDN U2205 ( .A(B[985]), .B(n2166), .Z(n2165) );
  NANDN U2206 ( .A(A[985]), .B(n37), .Z(n2166) );
  NANDN U2207 ( .A(n37), .B(A[985]), .Z(n2164) );
  AND U2208 ( .A(n2167), .B(n2168), .Z(n37) );
  NANDN U2209 ( .A(B[984]), .B(n2169), .Z(n2168) );
  NANDN U2210 ( .A(A[984]), .B(n39), .Z(n2169) );
  NANDN U2211 ( .A(n39), .B(A[984]), .Z(n2167) );
  AND U2212 ( .A(n2170), .B(n2171), .Z(n39) );
  NANDN U2213 ( .A(B[983]), .B(n2172), .Z(n2171) );
  NANDN U2214 ( .A(A[983]), .B(n41), .Z(n2172) );
  NANDN U2215 ( .A(n41), .B(A[983]), .Z(n2170) );
  AND U2216 ( .A(n2173), .B(n2174), .Z(n41) );
  NANDN U2217 ( .A(B[982]), .B(n2175), .Z(n2174) );
  NANDN U2218 ( .A(A[982]), .B(n43), .Z(n2175) );
  NANDN U2219 ( .A(n43), .B(A[982]), .Z(n2173) );
  AND U2220 ( .A(n2176), .B(n2177), .Z(n43) );
  NANDN U2221 ( .A(B[981]), .B(n2178), .Z(n2177) );
  NANDN U2222 ( .A(A[981]), .B(n45), .Z(n2178) );
  NANDN U2223 ( .A(n45), .B(A[981]), .Z(n2176) );
  AND U2224 ( .A(n2179), .B(n2180), .Z(n45) );
  NANDN U2225 ( .A(B[980]), .B(n2181), .Z(n2180) );
  NANDN U2226 ( .A(A[980]), .B(n47), .Z(n2181) );
  NANDN U2227 ( .A(n47), .B(A[980]), .Z(n2179) );
  AND U2228 ( .A(n2182), .B(n2183), .Z(n47) );
  NANDN U2229 ( .A(B[979]), .B(n2184), .Z(n2183) );
  NANDN U2230 ( .A(A[979]), .B(n51), .Z(n2184) );
  NANDN U2231 ( .A(n51), .B(A[979]), .Z(n2182) );
  AND U2232 ( .A(n2185), .B(n2186), .Z(n51) );
  NANDN U2233 ( .A(B[978]), .B(n2187), .Z(n2186) );
  NANDN U2234 ( .A(A[978]), .B(n53), .Z(n2187) );
  NANDN U2235 ( .A(n53), .B(A[978]), .Z(n2185) );
  AND U2236 ( .A(n2188), .B(n2189), .Z(n53) );
  NANDN U2237 ( .A(B[977]), .B(n2190), .Z(n2189) );
  NANDN U2238 ( .A(A[977]), .B(n55), .Z(n2190) );
  NANDN U2239 ( .A(n55), .B(A[977]), .Z(n2188) );
  AND U2240 ( .A(n2191), .B(n2192), .Z(n55) );
  NANDN U2241 ( .A(B[976]), .B(n2193), .Z(n2192) );
  NANDN U2242 ( .A(A[976]), .B(n57), .Z(n2193) );
  NANDN U2243 ( .A(n57), .B(A[976]), .Z(n2191) );
  AND U2244 ( .A(n2194), .B(n2195), .Z(n57) );
  NANDN U2245 ( .A(B[975]), .B(n2196), .Z(n2195) );
  NANDN U2246 ( .A(A[975]), .B(n59), .Z(n2196) );
  NANDN U2247 ( .A(n59), .B(A[975]), .Z(n2194) );
  AND U2248 ( .A(n2197), .B(n2198), .Z(n59) );
  NANDN U2249 ( .A(B[974]), .B(n2199), .Z(n2198) );
  NANDN U2250 ( .A(A[974]), .B(n61), .Z(n2199) );
  NANDN U2251 ( .A(n61), .B(A[974]), .Z(n2197) );
  AND U2252 ( .A(n2200), .B(n2201), .Z(n61) );
  NANDN U2253 ( .A(B[973]), .B(n2202), .Z(n2201) );
  NANDN U2254 ( .A(A[973]), .B(n63), .Z(n2202) );
  NANDN U2255 ( .A(n63), .B(A[973]), .Z(n2200) );
  AND U2256 ( .A(n2203), .B(n2204), .Z(n63) );
  NANDN U2257 ( .A(B[972]), .B(n2205), .Z(n2204) );
  NANDN U2258 ( .A(A[972]), .B(n65), .Z(n2205) );
  NANDN U2259 ( .A(n65), .B(A[972]), .Z(n2203) );
  AND U2260 ( .A(n2206), .B(n2207), .Z(n65) );
  NANDN U2261 ( .A(B[971]), .B(n2208), .Z(n2207) );
  NANDN U2262 ( .A(A[971]), .B(n67), .Z(n2208) );
  NANDN U2263 ( .A(n67), .B(A[971]), .Z(n2206) );
  AND U2264 ( .A(n2209), .B(n2210), .Z(n67) );
  NANDN U2265 ( .A(B[970]), .B(n2211), .Z(n2210) );
  NANDN U2266 ( .A(A[970]), .B(n69), .Z(n2211) );
  NANDN U2267 ( .A(n69), .B(A[970]), .Z(n2209) );
  AND U2268 ( .A(n2212), .B(n2213), .Z(n69) );
  NANDN U2269 ( .A(B[969]), .B(n2214), .Z(n2213) );
  NANDN U2270 ( .A(A[969]), .B(n73), .Z(n2214) );
  NANDN U2271 ( .A(n73), .B(A[969]), .Z(n2212) );
  AND U2272 ( .A(n2215), .B(n2216), .Z(n73) );
  NANDN U2273 ( .A(B[968]), .B(n2217), .Z(n2216) );
  NANDN U2274 ( .A(A[968]), .B(n75), .Z(n2217) );
  NANDN U2275 ( .A(n75), .B(A[968]), .Z(n2215) );
  AND U2276 ( .A(n2218), .B(n2219), .Z(n75) );
  NANDN U2277 ( .A(B[967]), .B(n2220), .Z(n2219) );
  NANDN U2278 ( .A(A[967]), .B(n77), .Z(n2220) );
  NANDN U2279 ( .A(n77), .B(A[967]), .Z(n2218) );
  AND U2280 ( .A(n2221), .B(n2222), .Z(n77) );
  NANDN U2281 ( .A(B[966]), .B(n2223), .Z(n2222) );
  NANDN U2282 ( .A(A[966]), .B(n79), .Z(n2223) );
  NANDN U2283 ( .A(n79), .B(A[966]), .Z(n2221) );
  AND U2284 ( .A(n2224), .B(n2225), .Z(n79) );
  NANDN U2285 ( .A(B[965]), .B(n2226), .Z(n2225) );
  NANDN U2286 ( .A(A[965]), .B(n81), .Z(n2226) );
  NANDN U2287 ( .A(n81), .B(A[965]), .Z(n2224) );
  AND U2288 ( .A(n2227), .B(n2228), .Z(n81) );
  NANDN U2289 ( .A(B[964]), .B(n2229), .Z(n2228) );
  NANDN U2290 ( .A(A[964]), .B(n83), .Z(n2229) );
  NANDN U2291 ( .A(n83), .B(A[964]), .Z(n2227) );
  AND U2292 ( .A(n2230), .B(n2231), .Z(n83) );
  NANDN U2293 ( .A(B[963]), .B(n2232), .Z(n2231) );
  NANDN U2294 ( .A(A[963]), .B(n85), .Z(n2232) );
  NANDN U2295 ( .A(n85), .B(A[963]), .Z(n2230) );
  AND U2296 ( .A(n2233), .B(n2234), .Z(n85) );
  NANDN U2297 ( .A(B[962]), .B(n2235), .Z(n2234) );
  NANDN U2298 ( .A(A[962]), .B(n87), .Z(n2235) );
  NANDN U2299 ( .A(n87), .B(A[962]), .Z(n2233) );
  AND U2300 ( .A(n2236), .B(n2237), .Z(n87) );
  NANDN U2301 ( .A(B[961]), .B(n2238), .Z(n2237) );
  NANDN U2302 ( .A(A[961]), .B(n89), .Z(n2238) );
  NANDN U2303 ( .A(n89), .B(A[961]), .Z(n2236) );
  AND U2304 ( .A(n2239), .B(n2240), .Z(n89) );
  NANDN U2305 ( .A(B[960]), .B(n2241), .Z(n2240) );
  NANDN U2306 ( .A(A[960]), .B(n91), .Z(n2241) );
  NANDN U2307 ( .A(n91), .B(A[960]), .Z(n2239) );
  AND U2308 ( .A(n2242), .B(n2243), .Z(n91) );
  NANDN U2309 ( .A(B[959]), .B(n2244), .Z(n2243) );
  NANDN U2310 ( .A(A[959]), .B(n95), .Z(n2244) );
  NANDN U2311 ( .A(n95), .B(A[959]), .Z(n2242) );
  AND U2312 ( .A(n2245), .B(n2246), .Z(n95) );
  NANDN U2313 ( .A(B[958]), .B(n2247), .Z(n2246) );
  NANDN U2314 ( .A(A[958]), .B(n97), .Z(n2247) );
  NANDN U2315 ( .A(n97), .B(A[958]), .Z(n2245) );
  AND U2316 ( .A(n2248), .B(n2249), .Z(n97) );
  NANDN U2317 ( .A(B[957]), .B(n2250), .Z(n2249) );
  NANDN U2318 ( .A(A[957]), .B(n99), .Z(n2250) );
  NANDN U2319 ( .A(n99), .B(A[957]), .Z(n2248) );
  AND U2320 ( .A(n2251), .B(n2252), .Z(n99) );
  NANDN U2321 ( .A(B[956]), .B(n2253), .Z(n2252) );
  NANDN U2322 ( .A(A[956]), .B(n101), .Z(n2253) );
  NANDN U2323 ( .A(n101), .B(A[956]), .Z(n2251) );
  AND U2324 ( .A(n2254), .B(n2255), .Z(n101) );
  NANDN U2325 ( .A(B[955]), .B(n2256), .Z(n2255) );
  NANDN U2326 ( .A(A[955]), .B(n103), .Z(n2256) );
  NANDN U2327 ( .A(n103), .B(A[955]), .Z(n2254) );
  AND U2328 ( .A(n2257), .B(n2258), .Z(n103) );
  NANDN U2329 ( .A(B[954]), .B(n2259), .Z(n2258) );
  NANDN U2330 ( .A(A[954]), .B(n105), .Z(n2259) );
  NANDN U2331 ( .A(n105), .B(A[954]), .Z(n2257) );
  AND U2332 ( .A(n2260), .B(n2261), .Z(n105) );
  NANDN U2333 ( .A(B[953]), .B(n2262), .Z(n2261) );
  NANDN U2334 ( .A(A[953]), .B(n107), .Z(n2262) );
  NANDN U2335 ( .A(n107), .B(A[953]), .Z(n2260) );
  AND U2336 ( .A(n2263), .B(n2264), .Z(n107) );
  NANDN U2337 ( .A(B[952]), .B(n2265), .Z(n2264) );
  NANDN U2338 ( .A(A[952]), .B(n109), .Z(n2265) );
  NANDN U2339 ( .A(n109), .B(A[952]), .Z(n2263) );
  AND U2340 ( .A(n2266), .B(n2267), .Z(n109) );
  NANDN U2341 ( .A(B[951]), .B(n2268), .Z(n2267) );
  NANDN U2342 ( .A(A[951]), .B(n111), .Z(n2268) );
  NANDN U2343 ( .A(n111), .B(A[951]), .Z(n2266) );
  AND U2344 ( .A(n2269), .B(n2270), .Z(n111) );
  NANDN U2345 ( .A(B[950]), .B(n2271), .Z(n2270) );
  NANDN U2346 ( .A(A[950]), .B(n113), .Z(n2271) );
  NANDN U2347 ( .A(n113), .B(A[950]), .Z(n2269) );
  AND U2348 ( .A(n2272), .B(n2273), .Z(n113) );
  NANDN U2349 ( .A(B[949]), .B(n2274), .Z(n2273) );
  NANDN U2350 ( .A(A[949]), .B(n117), .Z(n2274) );
  NANDN U2351 ( .A(n117), .B(A[949]), .Z(n2272) );
  AND U2352 ( .A(n2275), .B(n2276), .Z(n117) );
  NANDN U2353 ( .A(B[948]), .B(n2277), .Z(n2276) );
  NANDN U2354 ( .A(A[948]), .B(n119), .Z(n2277) );
  NANDN U2355 ( .A(n119), .B(A[948]), .Z(n2275) );
  AND U2356 ( .A(n2278), .B(n2279), .Z(n119) );
  NANDN U2357 ( .A(B[947]), .B(n2280), .Z(n2279) );
  NANDN U2358 ( .A(A[947]), .B(n121), .Z(n2280) );
  NANDN U2359 ( .A(n121), .B(A[947]), .Z(n2278) );
  AND U2360 ( .A(n2281), .B(n2282), .Z(n121) );
  NANDN U2361 ( .A(B[946]), .B(n2283), .Z(n2282) );
  NANDN U2362 ( .A(A[946]), .B(n123), .Z(n2283) );
  NANDN U2363 ( .A(n123), .B(A[946]), .Z(n2281) );
  AND U2364 ( .A(n2284), .B(n2285), .Z(n123) );
  NANDN U2365 ( .A(B[945]), .B(n2286), .Z(n2285) );
  NANDN U2366 ( .A(A[945]), .B(n125), .Z(n2286) );
  NANDN U2367 ( .A(n125), .B(A[945]), .Z(n2284) );
  AND U2368 ( .A(n2287), .B(n2288), .Z(n125) );
  NANDN U2369 ( .A(B[944]), .B(n2289), .Z(n2288) );
  NANDN U2370 ( .A(A[944]), .B(n127), .Z(n2289) );
  NANDN U2371 ( .A(n127), .B(A[944]), .Z(n2287) );
  AND U2372 ( .A(n2290), .B(n2291), .Z(n127) );
  NANDN U2373 ( .A(B[943]), .B(n2292), .Z(n2291) );
  NANDN U2374 ( .A(A[943]), .B(n129), .Z(n2292) );
  NANDN U2375 ( .A(n129), .B(A[943]), .Z(n2290) );
  AND U2376 ( .A(n2293), .B(n2294), .Z(n129) );
  NANDN U2377 ( .A(B[942]), .B(n2295), .Z(n2294) );
  NANDN U2378 ( .A(A[942]), .B(n131), .Z(n2295) );
  NANDN U2379 ( .A(n131), .B(A[942]), .Z(n2293) );
  AND U2380 ( .A(n2296), .B(n2297), .Z(n131) );
  NANDN U2381 ( .A(B[941]), .B(n2298), .Z(n2297) );
  NANDN U2382 ( .A(A[941]), .B(n133), .Z(n2298) );
  NANDN U2383 ( .A(n133), .B(A[941]), .Z(n2296) );
  AND U2384 ( .A(n2299), .B(n2300), .Z(n133) );
  NANDN U2385 ( .A(B[940]), .B(n2301), .Z(n2300) );
  NANDN U2386 ( .A(A[940]), .B(n135), .Z(n2301) );
  NANDN U2387 ( .A(n135), .B(A[940]), .Z(n2299) );
  AND U2388 ( .A(n2302), .B(n2303), .Z(n135) );
  NANDN U2389 ( .A(B[939]), .B(n2304), .Z(n2303) );
  NANDN U2390 ( .A(A[939]), .B(n139), .Z(n2304) );
  NANDN U2391 ( .A(n139), .B(A[939]), .Z(n2302) );
  AND U2392 ( .A(n2305), .B(n2306), .Z(n139) );
  NANDN U2393 ( .A(B[938]), .B(n2307), .Z(n2306) );
  NANDN U2394 ( .A(A[938]), .B(n141), .Z(n2307) );
  NANDN U2395 ( .A(n141), .B(A[938]), .Z(n2305) );
  AND U2396 ( .A(n2308), .B(n2309), .Z(n141) );
  NANDN U2397 ( .A(B[937]), .B(n2310), .Z(n2309) );
  NANDN U2398 ( .A(A[937]), .B(n143), .Z(n2310) );
  NANDN U2399 ( .A(n143), .B(A[937]), .Z(n2308) );
  AND U2400 ( .A(n2311), .B(n2312), .Z(n143) );
  NANDN U2401 ( .A(B[936]), .B(n2313), .Z(n2312) );
  NANDN U2402 ( .A(A[936]), .B(n145), .Z(n2313) );
  NANDN U2403 ( .A(n145), .B(A[936]), .Z(n2311) );
  AND U2404 ( .A(n2314), .B(n2315), .Z(n145) );
  NANDN U2405 ( .A(B[935]), .B(n2316), .Z(n2315) );
  NANDN U2406 ( .A(A[935]), .B(n147), .Z(n2316) );
  NANDN U2407 ( .A(n147), .B(A[935]), .Z(n2314) );
  AND U2408 ( .A(n2317), .B(n2318), .Z(n147) );
  NANDN U2409 ( .A(B[934]), .B(n2319), .Z(n2318) );
  NANDN U2410 ( .A(A[934]), .B(n149), .Z(n2319) );
  NANDN U2411 ( .A(n149), .B(A[934]), .Z(n2317) );
  AND U2412 ( .A(n2320), .B(n2321), .Z(n149) );
  NANDN U2413 ( .A(B[933]), .B(n2322), .Z(n2321) );
  NANDN U2414 ( .A(A[933]), .B(n151), .Z(n2322) );
  NANDN U2415 ( .A(n151), .B(A[933]), .Z(n2320) );
  AND U2416 ( .A(n2323), .B(n2324), .Z(n151) );
  NANDN U2417 ( .A(B[932]), .B(n2325), .Z(n2324) );
  NANDN U2418 ( .A(A[932]), .B(n153), .Z(n2325) );
  NANDN U2419 ( .A(n153), .B(A[932]), .Z(n2323) );
  AND U2420 ( .A(n2326), .B(n2327), .Z(n153) );
  NANDN U2421 ( .A(B[931]), .B(n2328), .Z(n2327) );
  NANDN U2422 ( .A(A[931]), .B(n155), .Z(n2328) );
  NANDN U2423 ( .A(n155), .B(A[931]), .Z(n2326) );
  AND U2424 ( .A(n2329), .B(n2330), .Z(n155) );
  NANDN U2425 ( .A(B[930]), .B(n2331), .Z(n2330) );
  NANDN U2426 ( .A(A[930]), .B(n157), .Z(n2331) );
  NANDN U2427 ( .A(n157), .B(A[930]), .Z(n2329) );
  AND U2428 ( .A(n2332), .B(n2333), .Z(n157) );
  NANDN U2429 ( .A(B[929]), .B(n2334), .Z(n2333) );
  NANDN U2430 ( .A(A[929]), .B(n161), .Z(n2334) );
  NANDN U2431 ( .A(n161), .B(A[929]), .Z(n2332) );
  AND U2432 ( .A(n2335), .B(n2336), .Z(n161) );
  NANDN U2433 ( .A(B[928]), .B(n2337), .Z(n2336) );
  NANDN U2434 ( .A(A[928]), .B(n163), .Z(n2337) );
  NANDN U2435 ( .A(n163), .B(A[928]), .Z(n2335) );
  AND U2436 ( .A(n2338), .B(n2339), .Z(n163) );
  NANDN U2437 ( .A(B[927]), .B(n2340), .Z(n2339) );
  NANDN U2438 ( .A(A[927]), .B(n165), .Z(n2340) );
  NANDN U2439 ( .A(n165), .B(A[927]), .Z(n2338) );
  AND U2440 ( .A(n2341), .B(n2342), .Z(n165) );
  NANDN U2441 ( .A(B[926]), .B(n2343), .Z(n2342) );
  NANDN U2442 ( .A(A[926]), .B(n167), .Z(n2343) );
  NANDN U2443 ( .A(n167), .B(A[926]), .Z(n2341) );
  AND U2444 ( .A(n2344), .B(n2345), .Z(n167) );
  NANDN U2445 ( .A(B[925]), .B(n2346), .Z(n2345) );
  NANDN U2446 ( .A(A[925]), .B(n169), .Z(n2346) );
  NANDN U2447 ( .A(n169), .B(A[925]), .Z(n2344) );
  AND U2448 ( .A(n2347), .B(n2348), .Z(n169) );
  NANDN U2449 ( .A(B[924]), .B(n2349), .Z(n2348) );
  NANDN U2450 ( .A(A[924]), .B(n171), .Z(n2349) );
  NANDN U2451 ( .A(n171), .B(A[924]), .Z(n2347) );
  AND U2452 ( .A(n2350), .B(n2351), .Z(n171) );
  NANDN U2453 ( .A(B[923]), .B(n2352), .Z(n2351) );
  NANDN U2454 ( .A(A[923]), .B(n173), .Z(n2352) );
  NANDN U2455 ( .A(n173), .B(A[923]), .Z(n2350) );
  AND U2456 ( .A(n2353), .B(n2354), .Z(n173) );
  NANDN U2457 ( .A(B[922]), .B(n2355), .Z(n2354) );
  NANDN U2458 ( .A(A[922]), .B(n175), .Z(n2355) );
  NANDN U2459 ( .A(n175), .B(A[922]), .Z(n2353) );
  AND U2460 ( .A(n2356), .B(n2357), .Z(n175) );
  NANDN U2461 ( .A(B[921]), .B(n2358), .Z(n2357) );
  NANDN U2462 ( .A(A[921]), .B(n177), .Z(n2358) );
  NANDN U2463 ( .A(n177), .B(A[921]), .Z(n2356) );
  AND U2464 ( .A(n2359), .B(n2360), .Z(n177) );
  NANDN U2465 ( .A(B[920]), .B(n2361), .Z(n2360) );
  NANDN U2466 ( .A(A[920]), .B(n179), .Z(n2361) );
  NANDN U2467 ( .A(n179), .B(A[920]), .Z(n2359) );
  AND U2468 ( .A(n2362), .B(n2363), .Z(n179) );
  NANDN U2469 ( .A(B[919]), .B(n2364), .Z(n2363) );
  NANDN U2470 ( .A(A[919]), .B(n183), .Z(n2364) );
  NANDN U2471 ( .A(n183), .B(A[919]), .Z(n2362) );
  AND U2472 ( .A(n2365), .B(n2366), .Z(n183) );
  NANDN U2473 ( .A(B[918]), .B(n2367), .Z(n2366) );
  NANDN U2474 ( .A(A[918]), .B(n185), .Z(n2367) );
  NANDN U2475 ( .A(n185), .B(A[918]), .Z(n2365) );
  AND U2476 ( .A(n2368), .B(n2369), .Z(n185) );
  NANDN U2477 ( .A(B[917]), .B(n2370), .Z(n2369) );
  NANDN U2478 ( .A(A[917]), .B(n187), .Z(n2370) );
  NANDN U2479 ( .A(n187), .B(A[917]), .Z(n2368) );
  AND U2480 ( .A(n2371), .B(n2372), .Z(n187) );
  NANDN U2481 ( .A(B[916]), .B(n2373), .Z(n2372) );
  NANDN U2482 ( .A(A[916]), .B(n189), .Z(n2373) );
  NANDN U2483 ( .A(n189), .B(A[916]), .Z(n2371) );
  AND U2484 ( .A(n2374), .B(n2375), .Z(n189) );
  NANDN U2485 ( .A(B[915]), .B(n2376), .Z(n2375) );
  NANDN U2486 ( .A(A[915]), .B(n191), .Z(n2376) );
  NANDN U2487 ( .A(n191), .B(A[915]), .Z(n2374) );
  AND U2488 ( .A(n2377), .B(n2378), .Z(n191) );
  NANDN U2489 ( .A(B[914]), .B(n2379), .Z(n2378) );
  NANDN U2490 ( .A(A[914]), .B(n193), .Z(n2379) );
  NANDN U2491 ( .A(n193), .B(A[914]), .Z(n2377) );
  AND U2492 ( .A(n2380), .B(n2381), .Z(n193) );
  NANDN U2493 ( .A(B[913]), .B(n2382), .Z(n2381) );
  NANDN U2494 ( .A(A[913]), .B(n195), .Z(n2382) );
  NANDN U2495 ( .A(n195), .B(A[913]), .Z(n2380) );
  AND U2496 ( .A(n2383), .B(n2384), .Z(n195) );
  NANDN U2497 ( .A(B[912]), .B(n2385), .Z(n2384) );
  NANDN U2498 ( .A(A[912]), .B(n197), .Z(n2385) );
  NANDN U2499 ( .A(n197), .B(A[912]), .Z(n2383) );
  AND U2500 ( .A(n2386), .B(n2387), .Z(n197) );
  NANDN U2501 ( .A(B[911]), .B(n2388), .Z(n2387) );
  NANDN U2502 ( .A(A[911]), .B(n199), .Z(n2388) );
  NANDN U2503 ( .A(n199), .B(A[911]), .Z(n2386) );
  AND U2504 ( .A(n2389), .B(n2390), .Z(n199) );
  NANDN U2505 ( .A(B[910]), .B(n2391), .Z(n2390) );
  NANDN U2506 ( .A(A[910]), .B(n201), .Z(n2391) );
  NANDN U2507 ( .A(n201), .B(A[910]), .Z(n2389) );
  AND U2508 ( .A(n2392), .B(n2393), .Z(n201) );
  NANDN U2509 ( .A(B[909]), .B(n2394), .Z(n2393) );
  NANDN U2510 ( .A(A[909]), .B(n205), .Z(n2394) );
  NANDN U2511 ( .A(n205), .B(A[909]), .Z(n2392) );
  AND U2512 ( .A(n2395), .B(n2396), .Z(n205) );
  NANDN U2513 ( .A(B[908]), .B(n2397), .Z(n2396) );
  NANDN U2514 ( .A(A[908]), .B(n207), .Z(n2397) );
  NANDN U2515 ( .A(n207), .B(A[908]), .Z(n2395) );
  AND U2516 ( .A(n2398), .B(n2399), .Z(n207) );
  NANDN U2517 ( .A(B[907]), .B(n2400), .Z(n2399) );
  NANDN U2518 ( .A(A[907]), .B(n209), .Z(n2400) );
  NANDN U2519 ( .A(n209), .B(A[907]), .Z(n2398) );
  AND U2520 ( .A(n2401), .B(n2402), .Z(n209) );
  NANDN U2521 ( .A(B[906]), .B(n2403), .Z(n2402) );
  NANDN U2522 ( .A(A[906]), .B(n211), .Z(n2403) );
  NANDN U2523 ( .A(n211), .B(A[906]), .Z(n2401) );
  AND U2524 ( .A(n2404), .B(n2405), .Z(n211) );
  NANDN U2525 ( .A(B[905]), .B(n2406), .Z(n2405) );
  NANDN U2526 ( .A(A[905]), .B(n213), .Z(n2406) );
  NANDN U2527 ( .A(n213), .B(A[905]), .Z(n2404) );
  AND U2528 ( .A(n2407), .B(n2408), .Z(n213) );
  NANDN U2529 ( .A(B[904]), .B(n2409), .Z(n2408) );
  NANDN U2530 ( .A(A[904]), .B(n215), .Z(n2409) );
  NANDN U2531 ( .A(n215), .B(A[904]), .Z(n2407) );
  AND U2532 ( .A(n2410), .B(n2411), .Z(n215) );
  NANDN U2533 ( .A(B[903]), .B(n2412), .Z(n2411) );
  NANDN U2534 ( .A(A[903]), .B(n217), .Z(n2412) );
  NANDN U2535 ( .A(n217), .B(A[903]), .Z(n2410) );
  AND U2536 ( .A(n2413), .B(n2414), .Z(n217) );
  NANDN U2537 ( .A(B[902]), .B(n2415), .Z(n2414) );
  NANDN U2538 ( .A(A[902]), .B(n219), .Z(n2415) );
  NANDN U2539 ( .A(n219), .B(A[902]), .Z(n2413) );
  AND U2540 ( .A(n2416), .B(n2417), .Z(n219) );
  NANDN U2541 ( .A(B[901]), .B(n2418), .Z(n2417) );
  NANDN U2542 ( .A(A[901]), .B(n221), .Z(n2418) );
  NANDN U2543 ( .A(n221), .B(A[901]), .Z(n2416) );
  AND U2544 ( .A(n2419), .B(n2420), .Z(n221) );
  NANDN U2545 ( .A(B[900]), .B(n2421), .Z(n2420) );
  NANDN U2546 ( .A(A[900]), .B(n223), .Z(n2421) );
  NANDN U2547 ( .A(n223), .B(A[900]), .Z(n2419) );
  AND U2548 ( .A(n2422), .B(n2423), .Z(n223) );
  NANDN U2549 ( .A(B[899]), .B(n2424), .Z(n2423) );
  NANDN U2550 ( .A(A[899]), .B(n229), .Z(n2424) );
  NANDN U2551 ( .A(n229), .B(A[899]), .Z(n2422) );
  AND U2552 ( .A(n2425), .B(n2426), .Z(n229) );
  NANDN U2553 ( .A(B[898]), .B(n2427), .Z(n2426) );
  NANDN U2554 ( .A(A[898]), .B(n231), .Z(n2427) );
  NANDN U2555 ( .A(n231), .B(A[898]), .Z(n2425) );
  AND U2556 ( .A(n2428), .B(n2429), .Z(n231) );
  NANDN U2557 ( .A(B[897]), .B(n2430), .Z(n2429) );
  NANDN U2558 ( .A(A[897]), .B(n233), .Z(n2430) );
  NANDN U2559 ( .A(n233), .B(A[897]), .Z(n2428) );
  AND U2560 ( .A(n2431), .B(n2432), .Z(n233) );
  NANDN U2561 ( .A(B[896]), .B(n2433), .Z(n2432) );
  NANDN U2562 ( .A(A[896]), .B(n235), .Z(n2433) );
  NANDN U2563 ( .A(n235), .B(A[896]), .Z(n2431) );
  AND U2564 ( .A(n2434), .B(n2435), .Z(n235) );
  NANDN U2565 ( .A(B[895]), .B(n2436), .Z(n2435) );
  NANDN U2566 ( .A(A[895]), .B(n237), .Z(n2436) );
  NANDN U2567 ( .A(n237), .B(A[895]), .Z(n2434) );
  AND U2568 ( .A(n2437), .B(n2438), .Z(n237) );
  NANDN U2569 ( .A(B[894]), .B(n2439), .Z(n2438) );
  NANDN U2570 ( .A(A[894]), .B(n239), .Z(n2439) );
  NANDN U2571 ( .A(n239), .B(A[894]), .Z(n2437) );
  AND U2572 ( .A(n2440), .B(n2441), .Z(n239) );
  NANDN U2573 ( .A(B[893]), .B(n2442), .Z(n2441) );
  NANDN U2574 ( .A(A[893]), .B(n241), .Z(n2442) );
  NANDN U2575 ( .A(n241), .B(A[893]), .Z(n2440) );
  AND U2576 ( .A(n2443), .B(n2444), .Z(n241) );
  NANDN U2577 ( .A(B[892]), .B(n2445), .Z(n2444) );
  NANDN U2578 ( .A(A[892]), .B(n243), .Z(n2445) );
  NANDN U2579 ( .A(n243), .B(A[892]), .Z(n2443) );
  AND U2580 ( .A(n2446), .B(n2447), .Z(n243) );
  NANDN U2581 ( .A(B[891]), .B(n2448), .Z(n2447) );
  NANDN U2582 ( .A(A[891]), .B(n245), .Z(n2448) );
  NANDN U2583 ( .A(n245), .B(A[891]), .Z(n2446) );
  AND U2584 ( .A(n2449), .B(n2450), .Z(n245) );
  NANDN U2585 ( .A(B[890]), .B(n2451), .Z(n2450) );
  NANDN U2586 ( .A(A[890]), .B(n247), .Z(n2451) );
  NANDN U2587 ( .A(n247), .B(A[890]), .Z(n2449) );
  AND U2588 ( .A(n2452), .B(n2453), .Z(n247) );
  NANDN U2589 ( .A(B[889]), .B(n2454), .Z(n2453) );
  NANDN U2590 ( .A(A[889]), .B(n251), .Z(n2454) );
  NANDN U2591 ( .A(n251), .B(A[889]), .Z(n2452) );
  AND U2592 ( .A(n2455), .B(n2456), .Z(n251) );
  NANDN U2593 ( .A(B[888]), .B(n2457), .Z(n2456) );
  NANDN U2594 ( .A(A[888]), .B(n253), .Z(n2457) );
  NANDN U2595 ( .A(n253), .B(A[888]), .Z(n2455) );
  AND U2596 ( .A(n2458), .B(n2459), .Z(n253) );
  NANDN U2597 ( .A(B[887]), .B(n2460), .Z(n2459) );
  NANDN U2598 ( .A(A[887]), .B(n255), .Z(n2460) );
  NANDN U2599 ( .A(n255), .B(A[887]), .Z(n2458) );
  AND U2600 ( .A(n2461), .B(n2462), .Z(n255) );
  NANDN U2601 ( .A(B[886]), .B(n2463), .Z(n2462) );
  NANDN U2602 ( .A(A[886]), .B(n257), .Z(n2463) );
  NANDN U2603 ( .A(n257), .B(A[886]), .Z(n2461) );
  AND U2604 ( .A(n2464), .B(n2465), .Z(n257) );
  NANDN U2605 ( .A(B[885]), .B(n2466), .Z(n2465) );
  NANDN U2606 ( .A(A[885]), .B(n259), .Z(n2466) );
  NANDN U2607 ( .A(n259), .B(A[885]), .Z(n2464) );
  AND U2608 ( .A(n2467), .B(n2468), .Z(n259) );
  NANDN U2609 ( .A(B[884]), .B(n2469), .Z(n2468) );
  NANDN U2610 ( .A(A[884]), .B(n261), .Z(n2469) );
  NANDN U2611 ( .A(n261), .B(A[884]), .Z(n2467) );
  AND U2612 ( .A(n2470), .B(n2471), .Z(n261) );
  NANDN U2613 ( .A(B[883]), .B(n2472), .Z(n2471) );
  NANDN U2614 ( .A(A[883]), .B(n263), .Z(n2472) );
  NANDN U2615 ( .A(n263), .B(A[883]), .Z(n2470) );
  AND U2616 ( .A(n2473), .B(n2474), .Z(n263) );
  NANDN U2617 ( .A(B[882]), .B(n2475), .Z(n2474) );
  NANDN U2618 ( .A(A[882]), .B(n265), .Z(n2475) );
  NANDN U2619 ( .A(n265), .B(A[882]), .Z(n2473) );
  AND U2620 ( .A(n2476), .B(n2477), .Z(n265) );
  NANDN U2621 ( .A(B[881]), .B(n2478), .Z(n2477) );
  NANDN U2622 ( .A(A[881]), .B(n267), .Z(n2478) );
  NANDN U2623 ( .A(n267), .B(A[881]), .Z(n2476) );
  AND U2624 ( .A(n2479), .B(n2480), .Z(n267) );
  NANDN U2625 ( .A(B[880]), .B(n2481), .Z(n2480) );
  NANDN U2626 ( .A(A[880]), .B(n269), .Z(n2481) );
  NANDN U2627 ( .A(n269), .B(A[880]), .Z(n2479) );
  AND U2628 ( .A(n2482), .B(n2483), .Z(n269) );
  NANDN U2629 ( .A(B[879]), .B(n2484), .Z(n2483) );
  NANDN U2630 ( .A(A[879]), .B(n273), .Z(n2484) );
  NANDN U2631 ( .A(n273), .B(A[879]), .Z(n2482) );
  AND U2632 ( .A(n2485), .B(n2486), .Z(n273) );
  NANDN U2633 ( .A(B[878]), .B(n2487), .Z(n2486) );
  NANDN U2634 ( .A(A[878]), .B(n275), .Z(n2487) );
  NANDN U2635 ( .A(n275), .B(A[878]), .Z(n2485) );
  AND U2636 ( .A(n2488), .B(n2489), .Z(n275) );
  NANDN U2637 ( .A(B[877]), .B(n2490), .Z(n2489) );
  NANDN U2638 ( .A(A[877]), .B(n277), .Z(n2490) );
  NANDN U2639 ( .A(n277), .B(A[877]), .Z(n2488) );
  AND U2640 ( .A(n2491), .B(n2492), .Z(n277) );
  NANDN U2641 ( .A(B[876]), .B(n2493), .Z(n2492) );
  NANDN U2642 ( .A(A[876]), .B(n279), .Z(n2493) );
  NANDN U2643 ( .A(n279), .B(A[876]), .Z(n2491) );
  AND U2644 ( .A(n2494), .B(n2495), .Z(n279) );
  NANDN U2645 ( .A(B[875]), .B(n2496), .Z(n2495) );
  NANDN U2646 ( .A(A[875]), .B(n281), .Z(n2496) );
  NANDN U2647 ( .A(n281), .B(A[875]), .Z(n2494) );
  AND U2648 ( .A(n2497), .B(n2498), .Z(n281) );
  NANDN U2649 ( .A(B[874]), .B(n2499), .Z(n2498) );
  NANDN U2650 ( .A(A[874]), .B(n283), .Z(n2499) );
  NANDN U2651 ( .A(n283), .B(A[874]), .Z(n2497) );
  AND U2652 ( .A(n2500), .B(n2501), .Z(n283) );
  NANDN U2653 ( .A(B[873]), .B(n2502), .Z(n2501) );
  NANDN U2654 ( .A(A[873]), .B(n285), .Z(n2502) );
  NANDN U2655 ( .A(n285), .B(A[873]), .Z(n2500) );
  AND U2656 ( .A(n2503), .B(n2504), .Z(n285) );
  NANDN U2657 ( .A(B[872]), .B(n2505), .Z(n2504) );
  NANDN U2658 ( .A(A[872]), .B(n287), .Z(n2505) );
  NANDN U2659 ( .A(n287), .B(A[872]), .Z(n2503) );
  AND U2660 ( .A(n2506), .B(n2507), .Z(n287) );
  NANDN U2661 ( .A(B[871]), .B(n2508), .Z(n2507) );
  NANDN U2662 ( .A(A[871]), .B(n289), .Z(n2508) );
  NANDN U2663 ( .A(n289), .B(A[871]), .Z(n2506) );
  AND U2664 ( .A(n2509), .B(n2510), .Z(n289) );
  NANDN U2665 ( .A(B[870]), .B(n2511), .Z(n2510) );
  NANDN U2666 ( .A(A[870]), .B(n291), .Z(n2511) );
  NANDN U2667 ( .A(n291), .B(A[870]), .Z(n2509) );
  AND U2668 ( .A(n2512), .B(n2513), .Z(n291) );
  NANDN U2669 ( .A(B[869]), .B(n2514), .Z(n2513) );
  NANDN U2670 ( .A(A[869]), .B(n295), .Z(n2514) );
  NANDN U2671 ( .A(n295), .B(A[869]), .Z(n2512) );
  AND U2672 ( .A(n2515), .B(n2516), .Z(n295) );
  NANDN U2673 ( .A(B[868]), .B(n2517), .Z(n2516) );
  NANDN U2674 ( .A(A[868]), .B(n297), .Z(n2517) );
  NANDN U2675 ( .A(n297), .B(A[868]), .Z(n2515) );
  AND U2676 ( .A(n2518), .B(n2519), .Z(n297) );
  NANDN U2677 ( .A(B[867]), .B(n2520), .Z(n2519) );
  NANDN U2678 ( .A(A[867]), .B(n299), .Z(n2520) );
  NANDN U2679 ( .A(n299), .B(A[867]), .Z(n2518) );
  AND U2680 ( .A(n2521), .B(n2522), .Z(n299) );
  NANDN U2681 ( .A(B[866]), .B(n2523), .Z(n2522) );
  NANDN U2682 ( .A(A[866]), .B(n301), .Z(n2523) );
  NANDN U2683 ( .A(n301), .B(A[866]), .Z(n2521) );
  AND U2684 ( .A(n2524), .B(n2525), .Z(n301) );
  NANDN U2685 ( .A(B[865]), .B(n2526), .Z(n2525) );
  NANDN U2686 ( .A(A[865]), .B(n303), .Z(n2526) );
  NANDN U2687 ( .A(n303), .B(A[865]), .Z(n2524) );
  AND U2688 ( .A(n2527), .B(n2528), .Z(n303) );
  NANDN U2689 ( .A(B[864]), .B(n2529), .Z(n2528) );
  NANDN U2690 ( .A(A[864]), .B(n305), .Z(n2529) );
  NANDN U2691 ( .A(n305), .B(A[864]), .Z(n2527) );
  AND U2692 ( .A(n2530), .B(n2531), .Z(n305) );
  NANDN U2693 ( .A(B[863]), .B(n2532), .Z(n2531) );
  NANDN U2694 ( .A(A[863]), .B(n307), .Z(n2532) );
  NANDN U2695 ( .A(n307), .B(A[863]), .Z(n2530) );
  AND U2696 ( .A(n2533), .B(n2534), .Z(n307) );
  NANDN U2697 ( .A(B[862]), .B(n2535), .Z(n2534) );
  NANDN U2698 ( .A(A[862]), .B(n309), .Z(n2535) );
  NANDN U2699 ( .A(n309), .B(A[862]), .Z(n2533) );
  AND U2700 ( .A(n2536), .B(n2537), .Z(n309) );
  NANDN U2701 ( .A(B[861]), .B(n2538), .Z(n2537) );
  NANDN U2702 ( .A(A[861]), .B(n311), .Z(n2538) );
  NANDN U2703 ( .A(n311), .B(A[861]), .Z(n2536) );
  AND U2704 ( .A(n2539), .B(n2540), .Z(n311) );
  NANDN U2705 ( .A(B[860]), .B(n2541), .Z(n2540) );
  NANDN U2706 ( .A(A[860]), .B(n313), .Z(n2541) );
  NANDN U2707 ( .A(n313), .B(A[860]), .Z(n2539) );
  AND U2708 ( .A(n2542), .B(n2543), .Z(n313) );
  NANDN U2709 ( .A(B[859]), .B(n2544), .Z(n2543) );
  NANDN U2710 ( .A(A[859]), .B(n317), .Z(n2544) );
  NANDN U2711 ( .A(n317), .B(A[859]), .Z(n2542) );
  AND U2712 ( .A(n2545), .B(n2546), .Z(n317) );
  NANDN U2713 ( .A(B[858]), .B(n2547), .Z(n2546) );
  NANDN U2714 ( .A(A[858]), .B(n319), .Z(n2547) );
  NANDN U2715 ( .A(n319), .B(A[858]), .Z(n2545) );
  AND U2716 ( .A(n2548), .B(n2549), .Z(n319) );
  NANDN U2717 ( .A(B[857]), .B(n2550), .Z(n2549) );
  NANDN U2718 ( .A(A[857]), .B(n321), .Z(n2550) );
  NANDN U2719 ( .A(n321), .B(A[857]), .Z(n2548) );
  AND U2720 ( .A(n2551), .B(n2552), .Z(n321) );
  NANDN U2721 ( .A(B[856]), .B(n2553), .Z(n2552) );
  NANDN U2722 ( .A(A[856]), .B(n323), .Z(n2553) );
  NANDN U2723 ( .A(n323), .B(A[856]), .Z(n2551) );
  AND U2724 ( .A(n2554), .B(n2555), .Z(n323) );
  NANDN U2725 ( .A(B[855]), .B(n2556), .Z(n2555) );
  NANDN U2726 ( .A(A[855]), .B(n325), .Z(n2556) );
  NANDN U2727 ( .A(n325), .B(A[855]), .Z(n2554) );
  AND U2728 ( .A(n2557), .B(n2558), .Z(n325) );
  NANDN U2729 ( .A(B[854]), .B(n2559), .Z(n2558) );
  NANDN U2730 ( .A(A[854]), .B(n327), .Z(n2559) );
  NANDN U2731 ( .A(n327), .B(A[854]), .Z(n2557) );
  AND U2732 ( .A(n2560), .B(n2561), .Z(n327) );
  NANDN U2733 ( .A(B[853]), .B(n2562), .Z(n2561) );
  NANDN U2734 ( .A(A[853]), .B(n329), .Z(n2562) );
  NANDN U2735 ( .A(n329), .B(A[853]), .Z(n2560) );
  AND U2736 ( .A(n2563), .B(n2564), .Z(n329) );
  NANDN U2737 ( .A(B[852]), .B(n2565), .Z(n2564) );
  NANDN U2738 ( .A(A[852]), .B(n331), .Z(n2565) );
  NANDN U2739 ( .A(n331), .B(A[852]), .Z(n2563) );
  AND U2740 ( .A(n2566), .B(n2567), .Z(n331) );
  NANDN U2741 ( .A(B[851]), .B(n2568), .Z(n2567) );
  NANDN U2742 ( .A(A[851]), .B(n333), .Z(n2568) );
  NANDN U2743 ( .A(n333), .B(A[851]), .Z(n2566) );
  AND U2744 ( .A(n2569), .B(n2570), .Z(n333) );
  NANDN U2745 ( .A(B[850]), .B(n2571), .Z(n2570) );
  NANDN U2746 ( .A(A[850]), .B(n335), .Z(n2571) );
  NANDN U2747 ( .A(n335), .B(A[850]), .Z(n2569) );
  AND U2748 ( .A(n2572), .B(n2573), .Z(n335) );
  NANDN U2749 ( .A(B[849]), .B(n2574), .Z(n2573) );
  NANDN U2750 ( .A(A[849]), .B(n339), .Z(n2574) );
  NANDN U2751 ( .A(n339), .B(A[849]), .Z(n2572) );
  AND U2752 ( .A(n2575), .B(n2576), .Z(n339) );
  NANDN U2753 ( .A(B[848]), .B(n2577), .Z(n2576) );
  NANDN U2754 ( .A(A[848]), .B(n341), .Z(n2577) );
  NANDN U2755 ( .A(n341), .B(A[848]), .Z(n2575) );
  AND U2756 ( .A(n2578), .B(n2579), .Z(n341) );
  NANDN U2757 ( .A(B[847]), .B(n2580), .Z(n2579) );
  NANDN U2758 ( .A(A[847]), .B(n343), .Z(n2580) );
  NANDN U2759 ( .A(n343), .B(A[847]), .Z(n2578) );
  AND U2760 ( .A(n2581), .B(n2582), .Z(n343) );
  NANDN U2761 ( .A(B[846]), .B(n2583), .Z(n2582) );
  NANDN U2762 ( .A(A[846]), .B(n345), .Z(n2583) );
  NANDN U2763 ( .A(n345), .B(A[846]), .Z(n2581) );
  AND U2764 ( .A(n2584), .B(n2585), .Z(n345) );
  NANDN U2765 ( .A(B[845]), .B(n2586), .Z(n2585) );
  NANDN U2766 ( .A(A[845]), .B(n347), .Z(n2586) );
  NANDN U2767 ( .A(n347), .B(A[845]), .Z(n2584) );
  AND U2768 ( .A(n2587), .B(n2588), .Z(n347) );
  NANDN U2769 ( .A(B[844]), .B(n2589), .Z(n2588) );
  NANDN U2770 ( .A(A[844]), .B(n349), .Z(n2589) );
  NANDN U2771 ( .A(n349), .B(A[844]), .Z(n2587) );
  AND U2772 ( .A(n2590), .B(n2591), .Z(n349) );
  NANDN U2773 ( .A(B[843]), .B(n2592), .Z(n2591) );
  NANDN U2774 ( .A(A[843]), .B(n351), .Z(n2592) );
  NANDN U2775 ( .A(n351), .B(A[843]), .Z(n2590) );
  AND U2776 ( .A(n2593), .B(n2594), .Z(n351) );
  NANDN U2777 ( .A(B[842]), .B(n2595), .Z(n2594) );
  NANDN U2778 ( .A(A[842]), .B(n353), .Z(n2595) );
  NANDN U2779 ( .A(n353), .B(A[842]), .Z(n2593) );
  AND U2780 ( .A(n2596), .B(n2597), .Z(n353) );
  NANDN U2781 ( .A(B[841]), .B(n2598), .Z(n2597) );
  NANDN U2782 ( .A(A[841]), .B(n355), .Z(n2598) );
  NANDN U2783 ( .A(n355), .B(A[841]), .Z(n2596) );
  AND U2784 ( .A(n2599), .B(n2600), .Z(n355) );
  NANDN U2785 ( .A(B[840]), .B(n2601), .Z(n2600) );
  NANDN U2786 ( .A(A[840]), .B(n357), .Z(n2601) );
  NANDN U2787 ( .A(n357), .B(A[840]), .Z(n2599) );
  AND U2788 ( .A(n2602), .B(n2603), .Z(n357) );
  NANDN U2789 ( .A(B[839]), .B(n2604), .Z(n2603) );
  NANDN U2790 ( .A(A[839]), .B(n361), .Z(n2604) );
  NANDN U2791 ( .A(n361), .B(A[839]), .Z(n2602) );
  AND U2792 ( .A(n2605), .B(n2606), .Z(n361) );
  NANDN U2793 ( .A(B[838]), .B(n2607), .Z(n2606) );
  NANDN U2794 ( .A(A[838]), .B(n363), .Z(n2607) );
  NANDN U2795 ( .A(n363), .B(A[838]), .Z(n2605) );
  AND U2796 ( .A(n2608), .B(n2609), .Z(n363) );
  NANDN U2797 ( .A(B[837]), .B(n2610), .Z(n2609) );
  NANDN U2798 ( .A(A[837]), .B(n365), .Z(n2610) );
  NANDN U2799 ( .A(n365), .B(A[837]), .Z(n2608) );
  AND U2800 ( .A(n2611), .B(n2612), .Z(n365) );
  NANDN U2801 ( .A(B[836]), .B(n2613), .Z(n2612) );
  NANDN U2802 ( .A(A[836]), .B(n367), .Z(n2613) );
  NANDN U2803 ( .A(n367), .B(A[836]), .Z(n2611) );
  AND U2804 ( .A(n2614), .B(n2615), .Z(n367) );
  NANDN U2805 ( .A(B[835]), .B(n2616), .Z(n2615) );
  NANDN U2806 ( .A(A[835]), .B(n369), .Z(n2616) );
  NANDN U2807 ( .A(n369), .B(A[835]), .Z(n2614) );
  AND U2808 ( .A(n2617), .B(n2618), .Z(n369) );
  NANDN U2809 ( .A(B[834]), .B(n2619), .Z(n2618) );
  NANDN U2810 ( .A(A[834]), .B(n371), .Z(n2619) );
  NANDN U2811 ( .A(n371), .B(A[834]), .Z(n2617) );
  AND U2812 ( .A(n2620), .B(n2621), .Z(n371) );
  NANDN U2813 ( .A(B[833]), .B(n2622), .Z(n2621) );
  NANDN U2814 ( .A(A[833]), .B(n373), .Z(n2622) );
  NANDN U2815 ( .A(n373), .B(A[833]), .Z(n2620) );
  AND U2816 ( .A(n2623), .B(n2624), .Z(n373) );
  NANDN U2817 ( .A(B[832]), .B(n2625), .Z(n2624) );
  NANDN U2818 ( .A(A[832]), .B(n375), .Z(n2625) );
  NANDN U2819 ( .A(n375), .B(A[832]), .Z(n2623) );
  AND U2820 ( .A(n2626), .B(n2627), .Z(n375) );
  NANDN U2821 ( .A(B[831]), .B(n2628), .Z(n2627) );
  NANDN U2822 ( .A(A[831]), .B(n377), .Z(n2628) );
  NANDN U2823 ( .A(n377), .B(A[831]), .Z(n2626) );
  AND U2824 ( .A(n2629), .B(n2630), .Z(n377) );
  NANDN U2825 ( .A(B[830]), .B(n2631), .Z(n2630) );
  NANDN U2826 ( .A(A[830]), .B(n379), .Z(n2631) );
  NANDN U2827 ( .A(n379), .B(A[830]), .Z(n2629) );
  AND U2828 ( .A(n2632), .B(n2633), .Z(n379) );
  NANDN U2829 ( .A(B[829]), .B(n2634), .Z(n2633) );
  NANDN U2830 ( .A(A[829]), .B(n383), .Z(n2634) );
  NANDN U2831 ( .A(n383), .B(A[829]), .Z(n2632) );
  AND U2832 ( .A(n2635), .B(n2636), .Z(n383) );
  NANDN U2833 ( .A(B[828]), .B(n2637), .Z(n2636) );
  NANDN U2834 ( .A(A[828]), .B(n385), .Z(n2637) );
  NANDN U2835 ( .A(n385), .B(A[828]), .Z(n2635) );
  AND U2836 ( .A(n2638), .B(n2639), .Z(n385) );
  NANDN U2837 ( .A(B[827]), .B(n2640), .Z(n2639) );
  NANDN U2838 ( .A(A[827]), .B(n387), .Z(n2640) );
  NANDN U2839 ( .A(n387), .B(A[827]), .Z(n2638) );
  AND U2840 ( .A(n2641), .B(n2642), .Z(n387) );
  NANDN U2841 ( .A(B[826]), .B(n2643), .Z(n2642) );
  NANDN U2842 ( .A(A[826]), .B(n389), .Z(n2643) );
  NANDN U2843 ( .A(n389), .B(A[826]), .Z(n2641) );
  AND U2844 ( .A(n2644), .B(n2645), .Z(n389) );
  NANDN U2845 ( .A(B[825]), .B(n2646), .Z(n2645) );
  NANDN U2846 ( .A(A[825]), .B(n391), .Z(n2646) );
  NANDN U2847 ( .A(n391), .B(A[825]), .Z(n2644) );
  AND U2848 ( .A(n2647), .B(n2648), .Z(n391) );
  NANDN U2849 ( .A(B[824]), .B(n2649), .Z(n2648) );
  NANDN U2850 ( .A(A[824]), .B(n393), .Z(n2649) );
  NANDN U2851 ( .A(n393), .B(A[824]), .Z(n2647) );
  AND U2852 ( .A(n2650), .B(n2651), .Z(n393) );
  NANDN U2853 ( .A(B[823]), .B(n2652), .Z(n2651) );
  NANDN U2854 ( .A(A[823]), .B(n395), .Z(n2652) );
  NANDN U2855 ( .A(n395), .B(A[823]), .Z(n2650) );
  AND U2856 ( .A(n2653), .B(n2654), .Z(n395) );
  NANDN U2857 ( .A(B[822]), .B(n2655), .Z(n2654) );
  NANDN U2858 ( .A(A[822]), .B(n397), .Z(n2655) );
  NANDN U2859 ( .A(n397), .B(A[822]), .Z(n2653) );
  AND U2860 ( .A(n2656), .B(n2657), .Z(n397) );
  NANDN U2861 ( .A(B[821]), .B(n2658), .Z(n2657) );
  NANDN U2862 ( .A(A[821]), .B(n399), .Z(n2658) );
  NANDN U2863 ( .A(n399), .B(A[821]), .Z(n2656) );
  AND U2864 ( .A(n2659), .B(n2660), .Z(n399) );
  NANDN U2865 ( .A(B[820]), .B(n2661), .Z(n2660) );
  NANDN U2866 ( .A(A[820]), .B(n401), .Z(n2661) );
  NANDN U2867 ( .A(n401), .B(A[820]), .Z(n2659) );
  AND U2868 ( .A(n2662), .B(n2663), .Z(n401) );
  NANDN U2869 ( .A(B[819]), .B(n2664), .Z(n2663) );
  NANDN U2870 ( .A(A[819]), .B(n405), .Z(n2664) );
  NANDN U2871 ( .A(n405), .B(A[819]), .Z(n2662) );
  AND U2872 ( .A(n2665), .B(n2666), .Z(n405) );
  NANDN U2873 ( .A(B[818]), .B(n2667), .Z(n2666) );
  NANDN U2874 ( .A(A[818]), .B(n407), .Z(n2667) );
  NANDN U2875 ( .A(n407), .B(A[818]), .Z(n2665) );
  AND U2876 ( .A(n2668), .B(n2669), .Z(n407) );
  NANDN U2877 ( .A(B[817]), .B(n2670), .Z(n2669) );
  NANDN U2878 ( .A(A[817]), .B(n409), .Z(n2670) );
  NANDN U2879 ( .A(n409), .B(A[817]), .Z(n2668) );
  AND U2880 ( .A(n2671), .B(n2672), .Z(n409) );
  NANDN U2881 ( .A(B[816]), .B(n2673), .Z(n2672) );
  NANDN U2882 ( .A(A[816]), .B(n411), .Z(n2673) );
  NANDN U2883 ( .A(n411), .B(A[816]), .Z(n2671) );
  AND U2884 ( .A(n2674), .B(n2675), .Z(n411) );
  NANDN U2885 ( .A(B[815]), .B(n2676), .Z(n2675) );
  NANDN U2886 ( .A(A[815]), .B(n413), .Z(n2676) );
  NANDN U2887 ( .A(n413), .B(A[815]), .Z(n2674) );
  AND U2888 ( .A(n2677), .B(n2678), .Z(n413) );
  NANDN U2889 ( .A(B[814]), .B(n2679), .Z(n2678) );
  NANDN U2890 ( .A(A[814]), .B(n415), .Z(n2679) );
  NANDN U2891 ( .A(n415), .B(A[814]), .Z(n2677) );
  AND U2892 ( .A(n2680), .B(n2681), .Z(n415) );
  NANDN U2893 ( .A(B[813]), .B(n2682), .Z(n2681) );
  NANDN U2894 ( .A(A[813]), .B(n417), .Z(n2682) );
  NANDN U2895 ( .A(n417), .B(A[813]), .Z(n2680) );
  AND U2896 ( .A(n2683), .B(n2684), .Z(n417) );
  NANDN U2897 ( .A(B[812]), .B(n2685), .Z(n2684) );
  NANDN U2898 ( .A(A[812]), .B(n419), .Z(n2685) );
  NANDN U2899 ( .A(n419), .B(A[812]), .Z(n2683) );
  AND U2900 ( .A(n2686), .B(n2687), .Z(n419) );
  NANDN U2901 ( .A(B[811]), .B(n2688), .Z(n2687) );
  NANDN U2902 ( .A(A[811]), .B(n421), .Z(n2688) );
  NANDN U2903 ( .A(n421), .B(A[811]), .Z(n2686) );
  AND U2904 ( .A(n2689), .B(n2690), .Z(n421) );
  NANDN U2905 ( .A(B[810]), .B(n2691), .Z(n2690) );
  NANDN U2906 ( .A(A[810]), .B(n423), .Z(n2691) );
  NANDN U2907 ( .A(n423), .B(A[810]), .Z(n2689) );
  AND U2908 ( .A(n2692), .B(n2693), .Z(n423) );
  NANDN U2909 ( .A(B[809]), .B(n2694), .Z(n2693) );
  NANDN U2910 ( .A(A[809]), .B(n427), .Z(n2694) );
  NANDN U2911 ( .A(n427), .B(A[809]), .Z(n2692) );
  AND U2912 ( .A(n2695), .B(n2696), .Z(n427) );
  NANDN U2913 ( .A(B[808]), .B(n2697), .Z(n2696) );
  NANDN U2914 ( .A(A[808]), .B(n429), .Z(n2697) );
  NANDN U2915 ( .A(n429), .B(A[808]), .Z(n2695) );
  AND U2916 ( .A(n2698), .B(n2699), .Z(n429) );
  NANDN U2917 ( .A(B[807]), .B(n2700), .Z(n2699) );
  NANDN U2918 ( .A(A[807]), .B(n431), .Z(n2700) );
  NANDN U2919 ( .A(n431), .B(A[807]), .Z(n2698) );
  AND U2920 ( .A(n2701), .B(n2702), .Z(n431) );
  NANDN U2921 ( .A(B[806]), .B(n2703), .Z(n2702) );
  NANDN U2922 ( .A(A[806]), .B(n433), .Z(n2703) );
  NANDN U2923 ( .A(n433), .B(A[806]), .Z(n2701) );
  AND U2924 ( .A(n2704), .B(n2705), .Z(n433) );
  NANDN U2925 ( .A(B[805]), .B(n2706), .Z(n2705) );
  NANDN U2926 ( .A(A[805]), .B(n435), .Z(n2706) );
  NANDN U2927 ( .A(n435), .B(A[805]), .Z(n2704) );
  AND U2928 ( .A(n2707), .B(n2708), .Z(n435) );
  NANDN U2929 ( .A(B[804]), .B(n2709), .Z(n2708) );
  NANDN U2930 ( .A(A[804]), .B(n437), .Z(n2709) );
  NANDN U2931 ( .A(n437), .B(A[804]), .Z(n2707) );
  AND U2932 ( .A(n2710), .B(n2711), .Z(n437) );
  NANDN U2933 ( .A(B[803]), .B(n2712), .Z(n2711) );
  NANDN U2934 ( .A(A[803]), .B(n439), .Z(n2712) );
  NANDN U2935 ( .A(n439), .B(A[803]), .Z(n2710) );
  AND U2936 ( .A(n2713), .B(n2714), .Z(n439) );
  NANDN U2937 ( .A(B[802]), .B(n2715), .Z(n2714) );
  NANDN U2938 ( .A(A[802]), .B(n441), .Z(n2715) );
  NANDN U2939 ( .A(n441), .B(A[802]), .Z(n2713) );
  AND U2940 ( .A(n2716), .B(n2717), .Z(n441) );
  NANDN U2941 ( .A(B[801]), .B(n2718), .Z(n2717) );
  NANDN U2942 ( .A(A[801]), .B(n443), .Z(n2718) );
  NANDN U2943 ( .A(n443), .B(A[801]), .Z(n2716) );
  AND U2944 ( .A(n2719), .B(n2720), .Z(n443) );
  NANDN U2945 ( .A(B[800]), .B(n2721), .Z(n2720) );
  NANDN U2946 ( .A(A[800]), .B(n445), .Z(n2721) );
  NANDN U2947 ( .A(n445), .B(A[800]), .Z(n2719) );
  AND U2948 ( .A(n2722), .B(n2723), .Z(n445) );
  NANDN U2949 ( .A(B[799]), .B(n2724), .Z(n2723) );
  NANDN U2950 ( .A(A[799]), .B(n451), .Z(n2724) );
  NANDN U2951 ( .A(n451), .B(A[799]), .Z(n2722) );
  AND U2952 ( .A(n2725), .B(n2726), .Z(n451) );
  NANDN U2953 ( .A(B[798]), .B(n2727), .Z(n2726) );
  NANDN U2954 ( .A(A[798]), .B(n453), .Z(n2727) );
  NANDN U2955 ( .A(n453), .B(A[798]), .Z(n2725) );
  AND U2956 ( .A(n2728), .B(n2729), .Z(n453) );
  NANDN U2957 ( .A(B[797]), .B(n2730), .Z(n2729) );
  NANDN U2958 ( .A(A[797]), .B(n455), .Z(n2730) );
  NANDN U2959 ( .A(n455), .B(A[797]), .Z(n2728) );
  AND U2960 ( .A(n2731), .B(n2732), .Z(n455) );
  NANDN U2961 ( .A(B[796]), .B(n2733), .Z(n2732) );
  NANDN U2962 ( .A(A[796]), .B(n457), .Z(n2733) );
  NANDN U2963 ( .A(n457), .B(A[796]), .Z(n2731) );
  AND U2964 ( .A(n2734), .B(n2735), .Z(n457) );
  NANDN U2965 ( .A(B[795]), .B(n2736), .Z(n2735) );
  NANDN U2966 ( .A(A[795]), .B(n459), .Z(n2736) );
  NANDN U2967 ( .A(n459), .B(A[795]), .Z(n2734) );
  AND U2968 ( .A(n2737), .B(n2738), .Z(n459) );
  NANDN U2969 ( .A(B[794]), .B(n2739), .Z(n2738) );
  NANDN U2970 ( .A(A[794]), .B(n461), .Z(n2739) );
  NANDN U2971 ( .A(n461), .B(A[794]), .Z(n2737) );
  AND U2972 ( .A(n2740), .B(n2741), .Z(n461) );
  NANDN U2973 ( .A(B[793]), .B(n2742), .Z(n2741) );
  NANDN U2974 ( .A(A[793]), .B(n463), .Z(n2742) );
  NANDN U2975 ( .A(n463), .B(A[793]), .Z(n2740) );
  AND U2976 ( .A(n2743), .B(n2744), .Z(n463) );
  NANDN U2977 ( .A(B[792]), .B(n2745), .Z(n2744) );
  NANDN U2978 ( .A(A[792]), .B(n465), .Z(n2745) );
  NANDN U2979 ( .A(n465), .B(A[792]), .Z(n2743) );
  AND U2980 ( .A(n2746), .B(n2747), .Z(n465) );
  NANDN U2981 ( .A(B[791]), .B(n2748), .Z(n2747) );
  NANDN U2982 ( .A(A[791]), .B(n467), .Z(n2748) );
  NANDN U2983 ( .A(n467), .B(A[791]), .Z(n2746) );
  AND U2984 ( .A(n2749), .B(n2750), .Z(n467) );
  NANDN U2985 ( .A(B[790]), .B(n2751), .Z(n2750) );
  NANDN U2986 ( .A(A[790]), .B(n469), .Z(n2751) );
  NANDN U2987 ( .A(n469), .B(A[790]), .Z(n2749) );
  AND U2988 ( .A(n2752), .B(n2753), .Z(n469) );
  NANDN U2989 ( .A(B[789]), .B(n2754), .Z(n2753) );
  NANDN U2990 ( .A(A[789]), .B(n473), .Z(n2754) );
  NANDN U2991 ( .A(n473), .B(A[789]), .Z(n2752) );
  AND U2992 ( .A(n2755), .B(n2756), .Z(n473) );
  NANDN U2993 ( .A(B[788]), .B(n2757), .Z(n2756) );
  NANDN U2994 ( .A(A[788]), .B(n475), .Z(n2757) );
  NANDN U2995 ( .A(n475), .B(A[788]), .Z(n2755) );
  AND U2996 ( .A(n2758), .B(n2759), .Z(n475) );
  NANDN U2997 ( .A(B[787]), .B(n2760), .Z(n2759) );
  NANDN U2998 ( .A(A[787]), .B(n477), .Z(n2760) );
  NANDN U2999 ( .A(n477), .B(A[787]), .Z(n2758) );
  AND U3000 ( .A(n2761), .B(n2762), .Z(n477) );
  NANDN U3001 ( .A(B[786]), .B(n2763), .Z(n2762) );
  NANDN U3002 ( .A(A[786]), .B(n479), .Z(n2763) );
  NANDN U3003 ( .A(n479), .B(A[786]), .Z(n2761) );
  AND U3004 ( .A(n2764), .B(n2765), .Z(n479) );
  NANDN U3005 ( .A(B[785]), .B(n2766), .Z(n2765) );
  NANDN U3006 ( .A(A[785]), .B(n481), .Z(n2766) );
  NANDN U3007 ( .A(n481), .B(A[785]), .Z(n2764) );
  AND U3008 ( .A(n2767), .B(n2768), .Z(n481) );
  NANDN U3009 ( .A(B[784]), .B(n2769), .Z(n2768) );
  NANDN U3010 ( .A(A[784]), .B(n483), .Z(n2769) );
  NANDN U3011 ( .A(n483), .B(A[784]), .Z(n2767) );
  AND U3012 ( .A(n2770), .B(n2771), .Z(n483) );
  NANDN U3013 ( .A(B[783]), .B(n2772), .Z(n2771) );
  NANDN U3014 ( .A(A[783]), .B(n485), .Z(n2772) );
  NANDN U3015 ( .A(n485), .B(A[783]), .Z(n2770) );
  AND U3016 ( .A(n2773), .B(n2774), .Z(n485) );
  NANDN U3017 ( .A(B[782]), .B(n2775), .Z(n2774) );
  NANDN U3018 ( .A(A[782]), .B(n487), .Z(n2775) );
  NANDN U3019 ( .A(n487), .B(A[782]), .Z(n2773) );
  AND U3020 ( .A(n2776), .B(n2777), .Z(n487) );
  NANDN U3021 ( .A(B[781]), .B(n2778), .Z(n2777) );
  NANDN U3022 ( .A(A[781]), .B(n489), .Z(n2778) );
  NANDN U3023 ( .A(n489), .B(A[781]), .Z(n2776) );
  AND U3024 ( .A(n2779), .B(n2780), .Z(n489) );
  NANDN U3025 ( .A(B[780]), .B(n2781), .Z(n2780) );
  NANDN U3026 ( .A(A[780]), .B(n491), .Z(n2781) );
  NANDN U3027 ( .A(n491), .B(A[780]), .Z(n2779) );
  AND U3028 ( .A(n2782), .B(n2783), .Z(n491) );
  NANDN U3029 ( .A(B[779]), .B(n2784), .Z(n2783) );
  NANDN U3030 ( .A(A[779]), .B(n495), .Z(n2784) );
  NANDN U3031 ( .A(n495), .B(A[779]), .Z(n2782) );
  AND U3032 ( .A(n2785), .B(n2786), .Z(n495) );
  NANDN U3033 ( .A(B[778]), .B(n2787), .Z(n2786) );
  NANDN U3034 ( .A(A[778]), .B(n497), .Z(n2787) );
  NANDN U3035 ( .A(n497), .B(A[778]), .Z(n2785) );
  AND U3036 ( .A(n2788), .B(n2789), .Z(n497) );
  NANDN U3037 ( .A(B[777]), .B(n2790), .Z(n2789) );
  NANDN U3038 ( .A(A[777]), .B(n499), .Z(n2790) );
  NANDN U3039 ( .A(n499), .B(A[777]), .Z(n2788) );
  AND U3040 ( .A(n2791), .B(n2792), .Z(n499) );
  NANDN U3041 ( .A(B[776]), .B(n2793), .Z(n2792) );
  NANDN U3042 ( .A(A[776]), .B(n501), .Z(n2793) );
  NANDN U3043 ( .A(n501), .B(A[776]), .Z(n2791) );
  AND U3044 ( .A(n2794), .B(n2795), .Z(n501) );
  NANDN U3045 ( .A(B[775]), .B(n2796), .Z(n2795) );
  NANDN U3046 ( .A(A[775]), .B(n503), .Z(n2796) );
  NANDN U3047 ( .A(n503), .B(A[775]), .Z(n2794) );
  AND U3048 ( .A(n2797), .B(n2798), .Z(n503) );
  NANDN U3049 ( .A(B[774]), .B(n2799), .Z(n2798) );
  NANDN U3050 ( .A(A[774]), .B(n505), .Z(n2799) );
  NANDN U3051 ( .A(n505), .B(A[774]), .Z(n2797) );
  AND U3052 ( .A(n2800), .B(n2801), .Z(n505) );
  NANDN U3053 ( .A(B[773]), .B(n2802), .Z(n2801) );
  NANDN U3054 ( .A(A[773]), .B(n507), .Z(n2802) );
  NANDN U3055 ( .A(n507), .B(A[773]), .Z(n2800) );
  AND U3056 ( .A(n2803), .B(n2804), .Z(n507) );
  NANDN U3057 ( .A(B[772]), .B(n2805), .Z(n2804) );
  NANDN U3058 ( .A(A[772]), .B(n509), .Z(n2805) );
  NANDN U3059 ( .A(n509), .B(A[772]), .Z(n2803) );
  AND U3060 ( .A(n2806), .B(n2807), .Z(n509) );
  NANDN U3061 ( .A(B[771]), .B(n2808), .Z(n2807) );
  NANDN U3062 ( .A(A[771]), .B(n511), .Z(n2808) );
  NANDN U3063 ( .A(n511), .B(A[771]), .Z(n2806) );
  AND U3064 ( .A(n2809), .B(n2810), .Z(n511) );
  NANDN U3065 ( .A(B[770]), .B(n2811), .Z(n2810) );
  NANDN U3066 ( .A(A[770]), .B(n513), .Z(n2811) );
  NANDN U3067 ( .A(n513), .B(A[770]), .Z(n2809) );
  AND U3068 ( .A(n2812), .B(n2813), .Z(n513) );
  NANDN U3069 ( .A(B[769]), .B(n2814), .Z(n2813) );
  NANDN U3070 ( .A(A[769]), .B(n517), .Z(n2814) );
  NANDN U3071 ( .A(n517), .B(A[769]), .Z(n2812) );
  AND U3072 ( .A(n2815), .B(n2816), .Z(n517) );
  NANDN U3073 ( .A(B[768]), .B(n2817), .Z(n2816) );
  NANDN U3074 ( .A(A[768]), .B(n519), .Z(n2817) );
  NANDN U3075 ( .A(n519), .B(A[768]), .Z(n2815) );
  AND U3076 ( .A(n2818), .B(n2819), .Z(n519) );
  NANDN U3077 ( .A(B[767]), .B(n2820), .Z(n2819) );
  NANDN U3078 ( .A(A[767]), .B(n521), .Z(n2820) );
  NANDN U3079 ( .A(n521), .B(A[767]), .Z(n2818) );
  AND U3080 ( .A(n2821), .B(n2822), .Z(n521) );
  NANDN U3081 ( .A(B[766]), .B(n2823), .Z(n2822) );
  NANDN U3082 ( .A(A[766]), .B(n523), .Z(n2823) );
  NANDN U3083 ( .A(n523), .B(A[766]), .Z(n2821) );
  AND U3084 ( .A(n2824), .B(n2825), .Z(n523) );
  NANDN U3085 ( .A(B[765]), .B(n2826), .Z(n2825) );
  NANDN U3086 ( .A(A[765]), .B(n525), .Z(n2826) );
  NANDN U3087 ( .A(n525), .B(A[765]), .Z(n2824) );
  AND U3088 ( .A(n2827), .B(n2828), .Z(n525) );
  NANDN U3089 ( .A(B[764]), .B(n2829), .Z(n2828) );
  NANDN U3090 ( .A(A[764]), .B(n527), .Z(n2829) );
  NANDN U3091 ( .A(n527), .B(A[764]), .Z(n2827) );
  AND U3092 ( .A(n2830), .B(n2831), .Z(n527) );
  NANDN U3093 ( .A(B[763]), .B(n2832), .Z(n2831) );
  NANDN U3094 ( .A(A[763]), .B(n529), .Z(n2832) );
  NANDN U3095 ( .A(n529), .B(A[763]), .Z(n2830) );
  AND U3096 ( .A(n2833), .B(n2834), .Z(n529) );
  NANDN U3097 ( .A(B[762]), .B(n2835), .Z(n2834) );
  NANDN U3098 ( .A(A[762]), .B(n531), .Z(n2835) );
  NANDN U3099 ( .A(n531), .B(A[762]), .Z(n2833) );
  AND U3100 ( .A(n2836), .B(n2837), .Z(n531) );
  NANDN U3101 ( .A(B[761]), .B(n2838), .Z(n2837) );
  NANDN U3102 ( .A(A[761]), .B(n533), .Z(n2838) );
  NANDN U3103 ( .A(n533), .B(A[761]), .Z(n2836) );
  AND U3104 ( .A(n2839), .B(n2840), .Z(n533) );
  NANDN U3105 ( .A(B[760]), .B(n2841), .Z(n2840) );
  NANDN U3106 ( .A(A[760]), .B(n535), .Z(n2841) );
  NANDN U3107 ( .A(n535), .B(A[760]), .Z(n2839) );
  AND U3108 ( .A(n2842), .B(n2843), .Z(n535) );
  NANDN U3109 ( .A(B[759]), .B(n2844), .Z(n2843) );
  NANDN U3110 ( .A(A[759]), .B(n539), .Z(n2844) );
  NANDN U3111 ( .A(n539), .B(A[759]), .Z(n2842) );
  AND U3112 ( .A(n2845), .B(n2846), .Z(n539) );
  NANDN U3113 ( .A(B[758]), .B(n2847), .Z(n2846) );
  NANDN U3114 ( .A(A[758]), .B(n541), .Z(n2847) );
  NANDN U3115 ( .A(n541), .B(A[758]), .Z(n2845) );
  AND U3116 ( .A(n2848), .B(n2849), .Z(n541) );
  NANDN U3117 ( .A(B[757]), .B(n2850), .Z(n2849) );
  NANDN U3118 ( .A(A[757]), .B(n543), .Z(n2850) );
  NANDN U3119 ( .A(n543), .B(A[757]), .Z(n2848) );
  AND U3120 ( .A(n2851), .B(n2852), .Z(n543) );
  NANDN U3121 ( .A(B[756]), .B(n2853), .Z(n2852) );
  NANDN U3122 ( .A(A[756]), .B(n545), .Z(n2853) );
  NANDN U3123 ( .A(n545), .B(A[756]), .Z(n2851) );
  AND U3124 ( .A(n2854), .B(n2855), .Z(n545) );
  NANDN U3125 ( .A(B[755]), .B(n2856), .Z(n2855) );
  NANDN U3126 ( .A(A[755]), .B(n547), .Z(n2856) );
  NANDN U3127 ( .A(n547), .B(A[755]), .Z(n2854) );
  AND U3128 ( .A(n2857), .B(n2858), .Z(n547) );
  NANDN U3129 ( .A(B[754]), .B(n2859), .Z(n2858) );
  NANDN U3130 ( .A(A[754]), .B(n549), .Z(n2859) );
  NANDN U3131 ( .A(n549), .B(A[754]), .Z(n2857) );
  AND U3132 ( .A(n2860), .B(n2861), .Z(n549) );
  NANDN U3133 ( .A(B[753]), .B(n2862), .Z(n2861) );
  NANDN U3134 ( .A(A[753]), .B(n551), .Z(n2862) );
  NANDN U3135 ( .A(n551), .B(A[753]), .Z(n2860) );
  AND U3136 ( .A(n2863), .B(n2864), .Z(n551) );
  NANDN U3137 ( .A(B[752]), .B(n2865), .Z(n2864) );
  NANDN U3138 ( .A(A[752]), .B(n553), .Z(n2865) );
  NANDN U3139 ( .A(n553), .B(A[752]), .Z(n2863) );
  AND U3140 ( .A(n2866), .B(n2867), .Z(n553) );
  NANDN U3141 ( .A(B[751]), .B(n2868), .Z(n2867) );
  NANDN U3142 ( .A(A[751]), .B(n555), .Z(n2868) );
  NANDN U3143 ( .A(n555), .B(A[751]), .Z(n2866) );
  AND U3144 ( .A(n2869), .B(n2870), .Z(n555) );
  NANDN U3145 ( .A(B[750]), .B(n2871), .Z(n2870) );
  NANDN U3146 ( .A(A[750]), .B(n557), .Z(n2871) );
  NANDN U3147 ( .A(n557), .B(A[750]), .Z(n2869) );
  AND U3148 ( .A(n2872), .B(n2873), .Z(n557) );
  NANDN U3149 ( .A(B[749]), .B(n2874), .Z(n2873) );
  NANDN U3150 ( .A(A[749]), .B(n561), .Z(n2874) );
  NANDN U3151 ( .A(n561), .B(A[749]), .Z(n2872) );
  AND U3152 ( .A(n2875), .B(n2876), .Z(n561) );
  NANDN U3153 ( .A(B[748]), .B(n2877), .Z(n2876) );
  NANDN U3154 ( .A(A[748]), .B(n563), .Z(n2877) );
  NANDN U3155 ( .A(n563), .B(A[748]), .Z(n2875) );
  AND U3156 ( .A(n2878), .B(n2879), .Z(n563) );
  NANDN U3157 ( .A(B[747]), .B(n2880), .Z(n2879) );
  NANDN U3158 ( .A(A[747]), .B(n565), .Z(n2880) );
  NANDN U3159 ( .A(n565), .B(A[747]), .Z(n2878) );
  AND U3160 ( .A(n2881), .B(n2882), .Z(n565) );
  NANDN U3161 ( .A(B[746]), .B(n2883), .Z(n2882) );
  NANDN U3162 ( .A(A[746]), .B(n567), .Z(n2883) );
  NANDN U3163 ( .A(n567), .B(A[746]), .Z(n2881) );
  AND U3164 ( .A(n2884), .B(n2885), .Z(n567) );
  NANDN U3165 ( .A(B[745]), .B(n2886), .Z(n2885) );
  NANDN U3166 ( .A(A[745]), .B(n569), .Z(n2886) );
  NANDN U3167 ( .A(n569), .B(A[745]), .Z(n2884) );
  AND U3168 ( .A(n2887), .B(n2888), .Z(n569) );
  NANDN U3169 ( .A(B[744]), .B(n2889), .Z(n2888) );
  NANDN U3170 ( .A(A[744]), .B(n571), .Z(n2889) );
  NANDN U3171 ( .A(n571), .B(A[744]), .Z(n2887) );
  AND U3172 ( .A(n2890), .B(n2891), .Z(n571) );
  NANDN U3173 ( .A(B[743]), .B(n2892), .Z(n2891) );
  NANDN U3174 ( .A(A[743]), .B(n573), .Z(n2892) );
  NANDN U3175 ( .A(n573), .B(A[743]), .Z(n2890) );
  AND U3176 ( .A(n2893), .B(n2894), .Z(n573) );
  NANDN U3177 ( .A(B[742]), .B(n2895), .Z(n2894) );
  NANDN U3178 ( .A(A[742]), .B(n575), .Z(n2895) );
  NANDN U3179 ( .A(n575), .B(A[742]), .Z(n2893) );
  AND U3180 ( .A(n2896), .B(n2897), .Z(n575) );
  NANDN U3181 ( .A(B[741]), .B(n2898), .Z(n2897) );
  NANDN U3182 ( .A(A[741]), .B(n577), .Z(n2898) );
  NANDN U3183 ( .A(n577), .B(A[741]), .Z(n2896) );
  AND U3184 ( .A(n2899), .B(n2900), .Z(n577) );
  NANDN U3185 ( .A(B[740]), .B(n2901), .Z(n2900) );
  NANDN U3186 ( .A(A[740]), .B(n579), .Z(n2901) );
  NANDN U3187 ( .A(n579), .B(A[740]), .Z(n2899) );
  AND U3188 ( .A(n2902), .B(n2903), .Z(n579) );
  NANDN U3189 ( .A(B[739]), .B(n2904), .Z(n2903) );
  NANDN U3190 ( .A(A[739]), .B(n583), .Z(n2904) );
  NANDN U3191 ( .A(n583), .B(A[739]), .Z(n2902) );
  AND U3192 ( .A(n2905), .B(n2906), .Z(n583) );
  NANDN U3193 ( .A(B[738]), .B(n2907), .Z(n2906) );
  NANDN U3194 ( .A(A[738]), .B(n585), .Z(n2907) );
  NANDN U3195 ( .A(n585), .B(A[738]), .Z(n2905) );
  AND U3196 ( .A(n2908), .B(n2909), .Z(n585) );
  NANDN U3197 ( .A(B[737]), .B(n2910), .Z(n2909) );
  NANDN U3198 ( .A(A[737]), .B(n587), .Z(n2910) );
  NANDN U3199 ( .A(n587), .B(A[737]), .Z(n2908) );
  AND U3200 ( .A(n2911), .B(n2912), .Z(n587) );
  NANDN U3201 ( .A(B[736]), .B(n2913), .Z(n2912) );
  NANDN U3202 ( .A(A[736]), .B(n589), .Z(n2913) );
  NANDN U3203 ( .A(n589), .B(A[736]), .Z(n2911) );
  AND U3204 ( .A(n2914), .B(n2915), .Z(n589) );
  NANDN U3205 ( .A(B[735]), .B(n2916), .Z(n2915) );
  NANDN U3206 ( .A(A[735]), .B(n591), .Z(n2916) );
  NANDN U3207 ( .A(n591), .B(A[735]), .Z(n2914) );
  AND U3208 ( .A(n2917), .B(n2918), .Z(n591) );
  NANDN U3209 ( .A(B[734]), .B(n2919), .Z(n2918) );
  NANDN U3210 ( .A(A[734]), .B(n593), .Z(n2919) );
  NANDN U3211 ( .A(n593), .B(A[734]), .Z(n2917) );
  AND U3212 ( .A(n2920), .B(n2921), .Z(n593) );
  NANDN U3213 ( .A(B[733]), .B(n2922), .Z(n2921) );
  NANDN U3214 ( .A(A[733]), .B(n595), .Z(n2922) );
  NANDN U3215 ( .A(n595), .B(A[733]), .Z(n2920) );
  AND U3216 ( .A(n2923), .B(n2924), .Z(n595) );
  NANDN U3217 ( .A(B[732]), .B(n2925), .Z(n2924) );
  NANDN U3218 ( .A(A[732]), .B(n597), .Z(n2925) );
  NANDN U3219 ( .A(n597), .B(A[732]), .Z(n2923) );
  AND U3220 ( .A(n2926), .B(n2927), .Z(n597) );
  NANDN U3221 ( .A(B[731]), .B(n2928), .Z(n2927) );
  NANDN U3222 ( .A(A[731]), .B(n599), .Z(n2928) );
  NANDN U3223 ( .A(n599), .B(A[731]), .Z(n2926) );
  AND U3224 ( .A(n2929), .B(n2930), .Z(n599) );
  NANDN U3225 ( .A(B[730]), .B(n2931), .Z(n2930) );
  NANDN U3226 ( .A(A[730]), .B(n601), .Z(n2931) );
  NANDN U3227 ( .A(n601), .B(A[730]), .Z(n2929) );
  AND U3228 ( .A(n2932), .B(n2933), .Z(n601) );
  NANDN U3229 ( .A(B[729]), .B(n2934), .Z(n2933) );
  NANDN U3230 ( .A(A[729]), .B(n605), .Z(n2934) );
  NANDN U3231 ( .A(n605), .B(A[729]), .Z(n2932) );
  AND U3232 ( .A(n2935), .B(n2936), .Z(n605) );
  NANDN U3233 ( .A(B[728]), .B(n2937), .Z(n2936) );
  NANDN U3234 ( .A(A[728]), .B(n607), .Z(n2937) );
  NANDN U3235 ( .A(n607), .B(A[728]), .Z(n2935) );
  AND U3236 ( .A(n2938), .B(n2939), .Z(n607) );
  NANDN U3237 ( .A(B[727]), .B(n2940), .Z(n2939) );
  NANDN U3238 ( .A(A[727]), .B(n609), .Z(n2940) );
  NANDN U3239 ( .A(n609), .B(A[727]), .Z(n2938) );
  AND U3240 ( .A(n2941), .B(n2942), .Z(n609) );
  NANDN U3241 ( .A(B[726]), .B(n2943), .Z(n2942) );
  NANDN U3242 ( .A(A[726]), .B(n611), .Z(n2943) );
  NANDN U3243 ( .A(n611), .B(A[726]), .Z(n2941) );
  AND U3244 ( .A(n2944), .B(n2945), .Z(n611) );
  NANDN U3245 ( .A(B[725]), .B(n2946), .Z(n2945) );
  NANDN U3246 ( .A(A[725]), .B(n613), .Z(n2946) );
  NANDN U3247 ( .A(n613), .B(A[725]), .Z(n2944) );
  AND U3248 ( .A(n2947), .B(n2948), .Z(n613) );
  NANDN U3249 ( .A(B[724]), .B(n2949), .Z(n2948) );
  NANDN U3250 ( .A(A[724]), .B(n615), .Z(n2949) );
  NANDN U3251 ( .A(n615), .B(A[724]), .Z(n2947) );
  AND U3252 ( .A(n2950), .B(n2951), .Z(n615) );
  NANDN U3253 ( .A(B[723]), .B(n2952), .Z(n2951) );
  NANDN U3254 ( .A(A[723]), .B(n617), .Z(n2952) );
  NANDN U3255 ( .A(n617), .B(A[723]), .Z(n2950) );
  AND U3256 ( .A(n2953), .B(n2954), .Z(n617) );
  NANDN U3257 ( .A(B[722]), .B(n2955), .Z(n2954) );
  NANDN U3258 ( .A(A[722]), .B(n619), .Z(n2955) );
  NANDN U3259 ( .A(n619), .B(A[722]), .Z(n2953) );
  AND U3260 ( .A(n2956), .B(n2957), .Z(n619) );
  NANDN U3261 ( .A(B[721]), .B(n2958), .Z(n2957) );
  NANDN U3262 ( .A(A[721]), .B(n621), .Z(n2958) );
  NANDN U3263 ( .A(n621), .B(A[721]), .Z(n2956) );
  AND U3264 ( .A(n2959), .B(n2960), .Z(n621) );
  NANDN U3265 ( .A(B[720]), .B(n2961), .Z(n2960) );
  NANDN U3266 ( .A(A[720]), .B(n623), .Z(n2961) );
  NANDN U3267 ( .A(n623), .B(A[720]), .Z(n2959) );
  AND U3268 ( .A(n2962), .B(n2963), .Z(n623) );
  NANDN U3269 ( .A(B[719]), .B(n2964), .Z(n2963) );
  NANDN U3270 ( .A(A[719]), .B(n627), .Z(n2964) );
  NANDN U3271 ( .A(n627), .B(A[719]), .Z(n2962) );
  AND U3272 ( .A(n2965), .B(n2966), .Z(n627) );
  NANDN U3273 ( .A(B[718]), .B(n2967), .Z(n2966) );
  NANDN U3274 ( .A(A[718]), .B(n629), .Z(n2967) );
  NANDN U3275 ( .A(n629), .B(A[718]), .Z(n2965) );
  AND U3276 ( .A(n2968), .B(n2969), .Z(n629) );
  NANDN U3277 ( .A(B[717]), .B(n2970), .Z(n2969) );
  NANDN U3278 ( .A(A[717]), .B(n631), .Z(n2970) );
  NANDN U3279 ( .A(n631), .B(A[717]), .Z(n2968) );
  AND U3280 ( .A(n2971), .B(n2972), .Z(n631) );
  NANDN U3281 ( .A(B[716]), .B(n2973), .Z(n2972) );
  NANDN U3282 ( .A(A[716]), .B(n633), .Z(n2973) );
  NANDN U3283 ( .A(n633), .B(A[716]), .Z(n2971) );
  AND U3284 ( .A(n2974), .B(n2975), .Z(n633) );
  NANDN U3285 ( .A(B[715]), .B(n2976), .Z(n2975) );
  NANDN U3286 ( .A(A[715]), .B(n635), .Z(n2976) );
  NANDN U3287 ( .A(n635), .B(A[715]), .Z(n2974) );
  AND U3288 ( .A(n2977), .B(n2978), .Z(n635) );
  NANDN U3289 ( .A(B[714]), .B(n2979), .Z(n2978) );
  NANDN U3290 ( .A(A[714]), .B(n637), .Z(n2979) );
  NANDN U3291 ( .A(n637), .B(A[714]), .Z(n2977) );
  AND U3292 ( .A(n2980), .B(n2981), .Z(n637) );
  NANDN U3293 ( .A(B[713]), .B(n2982), .Z(n2981) );
  NANDN U3294 ( .A(A[713]), .B(n639), .Z(n2982) );
  NANDN U3295 ( .A(n639), .B(A[713]), .Z(n2980) );
  AND U3296 ( .A(n2983), .B(n2984), .Z(n639) );
  NANDN U3297 ( .A(B[712]), .B(n2985), .Z(n2984) );
  NANDN U3298 ( .A(A[712]), .B(n641), .Z(n2985) );
  NANDN U3299 ( .A(n641), .B(A[712]), .Z(n2983) );
  AND U3300 ( .A(n2986), .B(n2987), .Z(n641) );
  NANDN U3301 ( .A(B[711]), .B(n2988), .Z(n2987) );
  NANDN U3302 ( .A(A[711]), .B(n643), .Z(n2988) );
  NANDN U3303 ( .A(n643), .B(A[711]), .Z(n2986) );
  AND U3304 ( .A(n2989), .B(n2990), .Z(n643) );
  NANDN U3305 ( .A(B[710]), .B(n2991), .Z(n2990) );
  NANDN U3306 ( .A(A[710]), .B(n645), .Z(n2991) );
  NANDN U3307 ( .A(n645), .B(A[710]), .Z(n2989) );
  AND U3308 ( .A(n2992), .B(n2993), .Z(n645) );
  NANDN U3309 ( .A(B[709]), .B(n2994), .Z(n2993) );
  NANDN U3310 ( .A(A[709]), .B(n649), .Z(n2994) );
  NANDN U3311 ( .A(n649), .B(A[709]), .Z(n2992) );
  AND U3312 ( .A(n2995), .B(n2996), .Z(n649) );
  NANDN U3313 ( .A(B[708]), .B(n2997), .Z(n2996) );
  NANDN U3314 ( .A(A[708]), .B(n651), .Z(n2997) );
  NANDN U3315 ( .A(n651), .B(A[708]), .Z(n2995) );
  AND U3316 ( .A(n2998), .B(n2999), .Z(n651) );
  NANDN U3317 ( .A(B[707]), .B(n3000), .Z(n2999) );
  NANDN U3318 ( .A(A[707]), .B(n653), .Z(n3000) );
  NANDN U3319 ( .A(n653), .B(A[707]), .Z(n2998) );
  AND U3320 ( .A(n3001), .B(n3002), .Z(n653) );
  NANDN U3321 ( .A(B[706]), .B(n3003), .Z(n3002) );
  NANDN U3322 ( .A(A[706]), .B(n655), .Z(n3003) );
  NANDN U3323 ( .A(n655), .B(A[706]), .Z(n3001) );
  AND U3324 ( .A(n3004), .B(n3005), .Z(n655) );
  NANDN U3325 ( .A(B[705]), .B(n3006), .Z(n3005) );
  NANDN U3326 ( .A(A[705]), .B(n657), .Z(n3006) );
  NANDN U3327 ( .A(n657), .B(A[705]), .Z(n3004) );
  AND U3328 ( .A(n3007), .B(n3008), .Z(n657) );
  NANDN U3329 ( .A(B[704]), .B(n3009), .Z(n3008) );
  NANDN U3330 ( .A(A[704]), .B(n659), .Z(n3009) );
  NANDN U3331 ( .A(n659), .B(A[704]), .Z(n3007) );
  AND U3332 ( .A(n3010), .B(n3011), .Z(n659) );
  NANDN U3333 ( .A(B[703]), .B(n3012), .Z(n3011) );
  NANDN U3334 ( .A(A[703]), .B(n661), .Z(n3012) );
  NANDN U3335 ( .A(n661), .B(A[703]), .Z(n3010) );
  AND U3336 ( .A(n3013), .B(n3014), .Z(n661) );
  NANDN U3337 ( .A(B[702]), .B(n3015), .Z(n3014) );
  NANDN U3338 ( .A(A[702]), .B(n663), .Z(n3015) );
  NANDN U3339 ( .A(n663), .B(A[702]), .Z(n3013) );
  AND U3340 ( .A(n3016), .B(n3017), .Z(n663) );
  NANDN U3341 ( .A(B[701]), .B(n3018), .Z(n3017) );
  NANDN U3342 ( .A(A[701]), .B(n665), .Z(n3018) );
  NANDN U3343 ( .A(n665), .B(A[701]), .Z(n3016) );
  AND U3344 ( .A(n3019), .B(n3020), .Z(n665) );
  NANDN U3345 ( .A(B[700]), .B(n3021), .Z(n3020) );
  NANDN U3346 ( .A(A[700]), .B(n667), .Z(n3021) );
  NANDN U3347 ( .A(n667), .B(A[700]), .Z(n3019) );
  AND U3348 ( .A(n3022), .B(n3023), .Z(n667) );
  NANDN U3349 ( .A(B[699]), .B(n3024), .Z(n3023) );
  NANDN U3350 ( .A(A[699]), .B(n673), .Z(n3024) );
  NANDN U3351 ( .A(n673), .B(A[699]), .Z(n3022) );
  AND U3352 ( .A(n3025), .B(n3026), .Z(n673) );
  NANDN U3353 ( .A(B[698]), .B(n3027), .Z(n3026) );
  NANDN U3354 ( .A(A[698]), .B(n675), .Z(n3027) );
  NANDN U3355 ( .A(n675), .B(A[698]), .Z(n3025) );
  AND U3356 ( .A(n3028), .B(n3029), .Z(n675) );
  NANDN U3357 ( .A(B[697]), .B(n3030), .Z(n3029) );
  NANDN U3358 ( .A(A[697]), .B(n677), .Z(n3030) );
  NANDN U3359 ( .A(n677), .B(A[697]), .Z(n3028) );
  AND U3360 ( .A(n3031), .B(n3032), .Z(n677) );
  NANDN U3361 ( .A(B[696]), .B(n3033), .Z(n3032) );
  NANDN U3362 ( .A(A[696]), .B(n679), .Z(n3033) );
  NANDN U3363 ( .A(n679), .B(A[696]), .Z(n3031) );
  AND U3364 ( .A(n3034), .B(n3035), .Z(n679) );
  NANDN U3365 ( .A(B[695]), .B(n3036), .Z(n3035) );
  NANDN U3366 ( .A(A[695]), .B(n681), .Z(n3036) );
  NANDN U3367 ( .A(n681), .B(A[695]), .Z(n3034) );
  AND U3368 ( .A(n3037), .B(n3038), .Z(n681) );
  NANDN U3369 ( .A(B[694]), .B(n3039), .Z(n3038) );
  NANDN U3370 ( .A(A[694]), .B(n683), .Z(n3039) );
  NANDN U3371 ( .A(n683), .B(A[694]), .Z(n3037) );
  AND U3372 ( .A(n3040), .B(n3041), .Z(n683) );
  NANDN U3373 ( .A(B[693]), .B(n3042), .Z(n3041) );
  NANDN U3374 ( .A(A[693]), .B(n685), .Z(n3042) );
  NANDN U3375 ( .A(n685), .B(A[693]), .Z(n3040) );
  AND U3376 ( .A(n3043), .B(n3044), .Z(n685) );
  NANDN U3377 ( .A(B[692]), .B(n3045), .Z(n3044) );
  NANDN U3378 ( .A(A[692]), .B(n687), .Z(n3045) );
  NANDN U3379 ( .A(n687), .B(A[692]), .Z(n3043) );
  AND U3380 ( .A(n3046), .B(n3047), .Z(n687) );
  NANDN U3381 ( .A(B[691]), .B(n3048), .Z(n3047) );
  NANDN U3382 ( .A(A[691]), .B(n689), .Z(n3048) );
  NANDN U3383 ( .A(n689), .B(A[691]), .Z(n3046) );
  AND U3384 ( .A(n3049), .B(n3050), .Z(n689) );
  NANDN U3385 ( .A(B[690]), .B(n3051), .Z(n3050) );
  NANDN U3386 ( .A(A[690]), .B(n691), .Z(n3051) );
  NANDN U3387 ( .A(n691), .B(A[690]), .Z(n3049) );
  AND U3388 ( .A(n3052), .B(n3053), .Z(n691) );
  NANDN U3389 ( .A(B[689]), .B(n3054), .Z(n3053) );
  NANDN U3390 ( .A(A[689]), .B(n695), .Z(n3054) );
  NANDN U3391 ( .A(n695), .B(A[689]), .Z(n3052) );
  AND U3392 ( .A(n3055), .B(n3056), .Z(n695) );
  NANDN U3393 ( .A(B[688]), .B(n3057), .Z(n3056) );
  NANDN U3394 ( .A(A[688]), .B(n697), .Z(n3057) );
  NANDN U3395 ( .A(n697), .B(A[688]), .Z(n3055) );
  AND U3396 ( .A(n3058), .B(n3059), .Z(n697) );
  NANDN U3397 ( .A(B[687]), .B(n3060), .Z(n3059) );
  NANDN U3398 ( .A(A[687]), .B(n699), .Z(n3060) );
  NANDN U3399 ( .A(n699), .B(A[687]), .Z(n3058) );
  AND U3400 ( .A(n3061), .B(n3062), .Z(n699) );
  NANDN U3401 ( .A(B[686]), .B(n3063), .Z(n3062) );
  NANDN U3402 ( .A(A[686]), .B(n701), .Z(n3063) );
  NANDN U3403 ( .A(n701), .B(A[686]), .Z(n3061) );
  AND U3404 ( .A(n3064), .B(n3065), .Z(n701) );
  NANDN U3405 ( .A(B[685]), .B(n3066), .Z(n3065) );
  NANDN U3406 ( .A(A[685]), .B(n703), .Z(n3066) );
  NANDN U3407 ( .A(n703), .B(A[685]), .Z(n3064) );
  AND U3408 ( .A(n3067), .B(n3068), .Z(n703) );
  NANDN U3409 ( .A(B[684]), .B(n3069), .Z(n3068) );
  NANDN U3410 ( .A(A[684]), .B(n705), .Z(n3069) );
  NANDN U3411 ( .A(n705), .B(A[684]), .Z(n3067) );
  AND U3412 ( .A(n3070), .B(n3071), .Z(n705) );
  NANDN U3413 ( .A(B[683]), .B(n3072), .Z(n3071) );
  NANDN U3414 ( .A(A[683]), .B(n707), .Z(n3072) );
  NANDN U3415 ( .A(n707), .B(A[683]), .Z(n3070) );
  AND U3416 ( .A(n3073), .B(n3074), .Z(n707) );
  NANDN U3417 ( .A(B[682]), .B(n3075), .Z(n3074) );
  NANDN U3418 ( .A(A[682]), .B(n709), .Z(n3075) );
  NANDN U3419 ( .A(n709), .B(A[682]), .Z(n3073) );
  AND U3420 ( .A(n3076), .B(n3077), .Z(n709) );
  NANDN U3421 ( .A(B[681]), .B(n3078), .Z(n3077) );
  NANDN U3422 ( .A(A[681]), .B(n711), .Z(n3078) );
  NANDN U3423 ( .A(n711), .B(A[681]), .Z(n3076) );
  AND U3424 ( .A(n3079), .B(n3080), .Z(n711) );
  NANDN U3425 ( .A(B[680]), .B(n3081), .Z(n3080) );
  NANDN U3426 ( .A(A[680]), .B(n713), .Z(n3081) );
  NANDN U3427 ( .A(n713), .B(A[680]), .Z(n3079) );
  AND U3428 ( .A(n3082), .B(n3083), .Z(n713) );
  NANDN U3429 ( .A(B[679]), .B(n3084), .Z(n3083) );
  NANDN U3430 ( .A(A[679]), .B(n717), .Z(n3084) );
  NANDN U3431 ( .A(n717), .B(A[679]), .Z(n3082) );
  AND U3432 ( .A(n3085), .B(n3086), .Z(n717) );
  NANDN U3433 ( .A(B[678]), .B(n3087), .Z(n3086) );
  NANDN U3434 ( .A(A[678]), .B(n719), .Z(n3087) );
  NANDN U3435 ( .A(n719), .B(A[678]), .Z(n3085) );
  AND U3436 ( .A(n3088), .B(n3089), .Z(n719) );
  NANDN U3437 ( .A(B[677]), .B(n3090), .Z(n3089) );
  NANDN U3438 ( .A(A[677]), .B(n721), .Z(n3090) );
  NANDN U3439 ( .A(n721), .B(A[677]), .Z(n3088) );
  AND U3440 ( .A(n3091), .B(n3092), .Z(n721) );
  NANDN U3441 ( .A(B[676]), .B(n3093), .Z(n3092) );
  NANDN U3442 ( .A(A[676]), .B(n723), .Z(n3093) );
  NANDN U3443 ( .A(n723), .B(A[676]), .Z(n3091) );
  AND U3444 ( .A(n3094), .B(n3095), .Z(n723) );
  NANDN U3445 ( .A(B[675]), .B(n3096), .Z(n3095) );
  NANDN U3446 ( .A(A[675]), .B(n725), .Z(n3096) );
  NANDN U3447 ( .A(n725), .B(A[675]), .Z(n3094) );
  AND U3448 ( .A(n3097), .B(n3098), .Z(n725) );
  NANDN U3449 ( .A(B[674]), .B(n3099), .Z(n3098) );
  NANDN U3450 ( .A(A[674]), .B(n727), .Z(n3099) );
  NANDN U3451 ( .A(n727), .B(A[674]), .Z(n3097) );
  AND U3452 ( .A(n3100), .B(n3101), .Z(n727) );
  NANDN U3453 ( .A(B[673]), .B(n3102), .Z(n3101) );
  NANDN U3454 ( .A(A[673]), .B(n729), .Z(n3102) );
  NANDN U3455 ( .A(n729), .B(A[673]), .Z(n3100) );
  AND U3456 ( .A(n3103), .B(n3104), .Z(n729) );
  NANDN U3457 ( .A(B[672]), .B(n3105), .Z(n3104) );
  NANDN U3458 ( .A(A[672]), .B(n731), .Z(n3105) );
  NANDN U3459 ( .A(n731), .B(A[672]), .Z(n3103) );
  AND U3460 ( .A(n3106), .B(n3107), .Z(n731) );
  NANDN U3461 ( .A(B[671]), .B(n3108), .Z(n3107) );
  NANDN U3462 ( .A(A[671]), .B(n733), .Z(n3108) );
  NANDN U3463 ( .A(n733), .B(A[671]), .Z(n3106) );
  AND U3464 ( .A(n3109), .B(n3110), .Z(n733) );
  NANDN U3465 ( .A(B[670]), .B(n3111), .Z(n3110) );
  NANDN U3466 ( .A(A[670]), .B(n735), .Z(n3111) );
  NANDN U3467 ( .A(n735), .B(A[670]), .Z(n3109) );
  AND U3468 ( .A(n3112), .B(n3113), .Z(n735) );
  NANDN U3469 ( .A(B[669]), .B(n3114), .Z(n3113) );
  NANDN U3470 ( .A(A[669]), .B(n739), .Z(n3114) );
  NANDN U3471 ( .A(n739), .B(A[669]), .Z(n3112) );
  AND U3472 ( .A(n3115), .B(n3116), .Z(n739) );
  NANDN U3473 ( .A(B[668]), .B(n3117), .Z(n3116) );
  NANDN U3474 ( .A(A[668]), .B(n741), .Z(n3117) );
  NANDN U3475 ( .A(n741), .B(A[668]), .Z(n3115) );
  AND U3476 ( .A(n3118), .B(n3119), .Z(n741) );
  NANDN U3477 ( .A(B[667]), .B(n3120), .Z(n3119) );
  NANDN U3478 ( .A(A[667]), .B(n743), .Z(n3120) );
  NANDN U3479 ( .A(n743), .B(A[667]), .Z(n3118) );
  AND U3480 ( .A(n3121), .B(n3122), .Z(n743) );
  NANDN U3481 ( .A(B[666]), .B(n3123), .Z(n3122) );
  NANDN U3482 ( .A(A[666]), .B(n745), .Z(n3123) );
  NANDN U3483 ( .A(n745), .B(A[666]), .Z(n3121) );
  AND U3484 ( .A(n3124), .B(n3125), .Z(n745) );
  NANDN U3485 ( .A(B[665]), .B(n3126), .Z(n3125) );
  NANDN U3486 ( .A(A[665]), .B(n747), .Z(n3126) );
  NANDN U3487 ( .A(n747), .B(A[665]), .Z(n3124) );
  AND U3488 ( .A(n3127), .B(n3128), .Z(n747) );
  NANDN U3489 ( .A(B[664]), .B(n3129), .Z(n3128) );
  NANDN U3490 ( .A(A[664]), .B(n749), .Z(n3129) );
  NANDN U3491 ( .A(n749), .B(A[664]), .Z(n3127) );
  AND U3492 ( .A(n3130), .B(n3131), .Z(n749) );
  NANDN U3493 ( .A(B[663]), .B(n3132), .Z(n3131) );
  NANDN U3494 ( .A(A[663]), .B(n751), .Z(n3132) );
  NANDN U3495 ( .A(n751), .B(A[663]), .Z(n3130) );
  AND U3496 ( .A(n3133), .B(n3134), .Z(n751) );
  NANDN U3497 ( .A(B[662]), .B(n3135), .Z(n3134) );
  NANDN U3498 ( .A(A[662]), .B(n753), .Z(n3135) );
  NANDN U3499 ( .A(n753), .B(A[662]), .Z(n3133) );
  AND U3500 ( .A(n3136), .B(n3137), .Z(n753) );
  NANDN U3501 ( .A(B[661]), .B(n3138), .Z(n3137) );
  NANDN U3502 ( .A(A[661]), .B(n755), .Z(n3138) );
  NANDN U3503 ( .A(n755), .B(A[661]), .Z(n3136) );
  AND U3504 ( .A(n3139), .B(n3140), .Z(n755) );
  NANDN U3505 ( .A(B[660]), .B(n3141), .Z(n3140) );
  NANDN U3506 ( .A(A[660]), .B(n757), .Z(n3141) );
  NANDN U3507 ( .A(n757), .B(A[660]), .Z(n3139) );
  AND U3508 ( .A(n3142), .B(n3143), .Z(n757) );
  NANDN U3509 ( .A(B[659]), .B(n3144), .Z(n3143) );
  NANDN U3510 ( .A(A[659]), .B(n761), .Z(n3144) );
  NANDN U3511 ( .A(n761), .B(A[659]), .Z(n3142) );
  AND U3512 ( .A(n3145), .B(n3146), .Z(n761) );
  NANDN U3513 ( .A(B[658]), .B(n3147), .Z(n3146) );
  NANDN U3514 ( .A(A[658]), .B(n763), .Z(n3147) );
  NANDN U3515 ( .A(n763), .B(A[658]), .Z(n3145) );
  AND U3516 ( .A(n3148), .B(n3149), .Z(n763) );
  NANDN U3517 ( .A(B[657]), .B(n3150), .Z(n3149) );
  NANDN U3518 ( .A(A[657]), .B(n765), .Z(n3150) );
  NANDN U3519 ( .A(n765), .B(A[657]), .Z(n3148) );
  AND U3520 ( .A(n3151), .B(n3152), .Z(n765) );
  NANDN U3521 ( .A(B[656]), .B(n3153), .Z(n3152) );
  NANDN U3522 ( .A(A[656]), .B(n767), .Z(n3153) );
  NANDN U3523 ( .A(n767), .B(A[656]), .Z(n3151) );
  AND U3524 ( .A(n3154), .B(n3155), .Z(n767) );
  NANDN U3525 ( .A(B[655]), .B(n3156), .Z(n3155) );
  NANDN U3526 ( .A(A[655]), .B(n769), .Z(n3156) );
  NANDN U3527 ( .A(n769), .B(A[655]), .Z(n3154) );
  AND U3528 ( .A(n3157), .B(n3158), .Z(n769) );
  NANDN U3529 ( .A(B[654]), .B(n3159), .Z(n3158) );
  NANDN U3530 ( .A(A[654]), .B(n771), .Z(n3159) );
  NANDN U3531 ( .A(n771), .B(A[654]), .Z(n3157) );
  AND U3532 ( .A(n3160), .B(n3161), .Z(n771) );
  NANDN U3533 ( .A(B[653]), .B(n3162), .Z(n3161) );
  NANDN U3534 ( .A(A[653]), .B(n773), .Z(n3162) );
  NANDN U3535 ( .A(n773), .B(A[653]), .Z(n3160) );
  AND U3536 ( .A(n3163), .B(n3164), .Z(n773) );
  NANDN U3537 ( .A(B[652]), .B(n3165), .Z(n3164) );
  NANDN U3538 ( .A(A[652]), .B(n775), .Z(n3165) );
  NANDN U3539 ( .A(n775), .B(A[652]), .Z(n3163) );
  AND U3540 ( .A(n3166), .B(n3167), .Z(n775) );
  NANDN U3541 ( .A(B[651]), .B(n3168), .Z(n3167) );
  NANDN U3542 ( .A(A[651]), .B(n777), .Z(n3168) );
  NANDN U3543 ( .A(n777), .B(A[651]), .Z(n3166) );
  AND U3544 ( .A(n3169), .B(n3170), .Z(n777) );
  NANDN U3545 ( .A(B[650]), .B(n3171), .Z(n3170) );
  NANDN U3546 ( .A(A[650]), .B(n779), .Z(n3171) );
  NANDN U3547 ( .A(n779), .B(A[650]), .Z(n3169) );
  AND U3548 ( .A(n3172), .B(n3173), .Z(n779) );
  NANDN U3549 ( .A(B[649]), .B(n3174), .Z(n3173) );
  NANDN U3550 ( .A(A[649]), .B(n783), .Z(n3174) );
  NANDN U3551 ( .A(n783), .B(A[649]), .Z(n3172) );
  AND U3552 ( .A(n3175), .B(n3176), .Z(n783) );
  NANDN U3553 ( .A(B[648]), .B(n3177), .Z(n3176) );
  NANDN U3554 ( .A(A[648]), .B(n785), .Z(n3177) );
  NANDN U3555 ( .A(n785), .B(A[648]), .Z(n3175) );
  AND U3556 ( .A(n3178), .B(n3179), .Z(n785) );
  NANDN U3557 ( .A(B[647]), .B(n3180), .Z(n3179) );
  NANDN U3558 ( .A(A[647]), .B(n787), .Z(n3180) );
  NANDN U3559 ( .A(n787), .B(A[647]), .Z(n3178) );
  AND U3560 ( .A(n3181), .B(n3182), .Z(n787) );
  NANDN U3561 ( .A(B[646]), .B(n3183), .Z(n3182) );
  NANDN U3562 ( .A(A[646]), .B(n789), .Z(n3183) );
  NANDN U3563 ( .A(n789), .B(A[646]), .Z(n3181) );
  AND U3564 ( .A(n3184), .B(n3185), .Z(n789) );
  NANDN U3565 ( .A(B[645]), .B(n3186), .Z(n3185) );
  NANDN U3566 ( .A(A[645]), .B(n791), .Z(n3186) );
  NANDN U3567 ( .A(n791), .B(A[645]), .Z(n3184) );
  AND U3568 ( .A(n3187), .B(n3188), .Z(n791) );
  NANDN U3569 ( .A(B[644]), .B(n3189), .Z(n3188) );
  NANDN U3570 ( .A(A[644]), .B(n793), .Z(n3189) );
  NANDN U3571 ( .A(n793), .B(A[644]), .Z(n3187) );
  AND U3572 ( .A(n3190), .B(n3191), .Z(n793) );
  NANDN U3573 ( .A(B[643]), .B(n3192), .Z(n3191) );
  NANDN U3574 ( .A(A[643]), .B(n795), .Z(n3192) );
  NANDN U3575 ( .A(n795), .B(A[643]), .Z(n3190) );
  AND U3576 ( .A(n3193), .B(n3194), .Z(n795) );
  NANDN U3577 ( .A(B[642]), .B(n3195), .Z(n3194) );
  NANDN U3578 ( .A(A[642]), .B(n797), .Z(n3195) );
  NANDN U3579 ( .A(n797), .B(A[642]), .Z(n3193) );
  AND U3580 ( .A(n3196), .B(n3197), .Z(n797) );
  NANDN U3581 ( .A(B[641]), .B(n3198), .Z(n3197) );
  NANDN U3582 ( .A(A[641]), .B(n799), .Z(n3198) );
  NANDN U3583 ( .A(n799), .B(A[641]), .Z(n3196) );
  AND U3584 ( .A(n3199), .B(n3200), .Z(n799) );
  NANDN U3585 ( .A(B[640]), .B(n3201), .Z(n3200) );
  NANDN U3586 ( .A(A[640]), .B(n801), .Z(n3201) );
  NANDN U3587 ( .A(n801), .B(A[640]), .Z(n3199) );
  AND U3588 ( .A(n3202), .B(n3203), .Z(n801) );
  NANDN U3589 ( .A(B[639]), .B(n3204), .Z(n3203) );
  NANDN U3590 ( .A(A[639]), .B(n805), .Z(n3204) );
  NANDN U3591 ( .A(n805), .B(A[639]), .Z(n3202) );
  AND U3592 ( .A(n3205), .B(n3206), .Z(n805) );
  NANDN U3593 ( .A(B[638]), .B(n3207), .Z(n3206) );
  NANDN U3594 ( .A(A[638]), .B(n807), .Z(n3207) );
  NANDN U3595 ( .A(n807), .B(A[638]), .Z(n3205) );
  AND U3596 ( .A(n3208), .B(n3209), .Z(n807) );
  NANDN U3597 ( .A(B[637]), .B(n3210), .Z(n3209) );
  NANDN U3598 ( .A(A[637]), .B(n809), .Z(n3210) );
  NANDN U3599 ( .A(n809), .B(A[637]), .Z(n3208) );
  AND U3600 ( .A(n3211), .B(n3212), .Z(n809) );
  NANDN U3601 ( .A(B[636]), .B(n3213), .Z(n3212) );
  NANDN U3602 ( .A(A[636]), .B(n811), .Z(n3213) );
  NANDN U3603 ( .A(n811), .B(A[636]), .Z(n3211) );
  AND U3604 ( .A(n3214), .B(n3215), .Z(n811) );
  NANDN U3605 ( .A(B[635]), .B(n3216), .Z(n3215) );
  NANDN U3606 ( .A(A[635]), .B(n813), .Z(n3216) );
  NANDN U3607 ( .A(n813), .B(A[635]), .Z(n3214) );
  AND U3608 ( .A(n3217), .B(n3218), .Z(n813) );
  NANDN U3609 ( .A(B[634]), .B(n3219), .Z(n3218) );
  NANDN U3610 ( .A(A[634]), .B(n815), .Z(n3219) );
  NANDN U3611 ( .A(n815), .B(A[634]), .Z(n3217) );
  AND U3612 ( .A(n3220), .B(n3221), .Z(n815) );
  NANDN U3613 ( .A(B[633]), .B(n3222), .Z(n3221) );
  NANDN U3614 ( .A(A[633]), .B(n817), .Z(n3222) );
  NANDN U3615 ( .A(n817), .B(A[633]), .Z(n3220) );
  AND U3616 ( .A(n3223), .B(n3224), .Z(n817) );
  NANDN U3617 ( .A(B[632]), .B(n3225), .Z(n3224) );
  NANDN U3618 ( .A(A[632]), .B(n819), .Z(n3225) );
  NANDN U3619 ( .A(n819), .B(A[632]), .Z(n3223) );
  AND U3620 ( .A(n3226), .B(n3227), .Z(n819) );
  NANDN U3621 ( .A(B[631]), .B(n3228), .Z(n3227) );
  NANDN U3622 ( .A(A[631]), .B(n821), .Z(n3228) );
  NANDN U3623 ( .A(n821), .B(A[631]), .Z(n3226) );
  AND U3624 ( .A(n3229), .B(n3230), .Z(n821) );
  NANDN U3625 ( .A(B[630]), .B(n3231), .Z(n3230) );
  NANDN U3626 ( .A(A[630]), .B(n823), .Z(n3231) );
  NANDN U3627 ( .A(n823), .B(A[630]), .Z(n3229) );
  AND U3628 ( .A(n3232), .B(n3233), .Z(n823) );
  NANDN U3629 ( .A(B[629]), .B(n3234), .Z(n3233) );
  NANDN U3630 ( .A(A[629]), .B(n827), .Z(n3234) );
  NANDN U3631 ( .A(n827), .B(A[629]), .Z(n3232) );
  AND U3632 ( .A(n3235), .B(n3236), .Z(n827) );
  NANDN U3633 ( .A(B[628]), .B(n3237), .Z(n3236) );
  NANDN U3634 ( .A(A[628]), .B(n829), .Z(n3237) );
  NANDN U3635 ( .A(n829), .B(A[628]), .Z(n3235) );
  AND U3636 ( .A(n3238), .B(n3239), .Z(n829) );
  NANDN U3637 ( .A(B[627]), .B(n3240), .Z(n3239) );
  NANDN U3638 ( .A(A[627]), .B(n831), .Z(n3240) );
  NANDN U3639 ( .A(n831), .B(A[627]), .Z(n3238) );
  AND U3640 ( .A(n3241), .B(n3242), .Z(n831) );
  NANDN U3641 ( .A(B[626]), .B(n3243), .Z(n3242) );
  NANDN U3642 ( .A(A[626]), .B(n833), .Z(n3243) );
  NANDN U3643 ( .A(n833), .B(A[626]), .Z(n3241) );
  AND U3644 ( .A(n3244), .B(n3245), .Z(n833) );
  NANDN U3645 ( .A(B[625]), .B(n3246), .Z(n3245) );
  NANDN U3646 ( .A(A[625]), .B(n835), .Z(n3246) );
  NANDN U3647 ( .A(n835), .B(A[625]), .Z(n3244) );
  AND U3648 ( .A(n3247), .B(n3248), .Z(n835) );
  NANDN U3649 ( .A(B[624]), .B(n3249), .Z(n3248) );
  NANDN U3650 ( .A(A[624]), .B(n837), .Z(n3249) );
  NANDN U3651 ( .A(n837), .B(A[624]), .Z(n3247) );
  AND U3652 ( .A(n3250), .B(n3251), .Z(n837) );
  NANDN U3653 ( .A(B[623]), .B(n3252), .Z(n3251) );
  NANDN U3654 ( .A(A[623]), .B(n839), .Z(n3252) );
  NANDN U3655 ( .A(n839), .B(A[623]), .Z(n3250) );
  AND U3656 ( .A(n3253), .B(n3254), .Z(n839) );
  NANDN U3657 ( .A(B[622]), .B(n3255), .Z(n3254) );
  NANDN U3658 ( .A(A[622]), .B(n841), .Z(n3255) );
  NANDN U3659 ( .A(n841), .B(A[622]), .Z(n3253) );
  AND U3660 ( .A(n3256), .B(n3257), .Z(n841) );
  NANDN U3661 ( .A(B[621]), .B(n3258), .Z(n3257) );
  NANDN U3662 ( .A(A[621]), .B(n843), .Z(n3258) );
  NANDN U3663 ( .A(n843), .B(A[621]), .Z(n3256) );
  AND U3664 ( .A(n3259), .B(n3260), .Z(n843) );
  NANDN U3665 ( .A(B[620]), .B(n3261), .Z(n3260) );
  NANDN U3666 ( .A(A[620]), .B(n845), .Z(n3261) );
  NANDN U3667 ( .A(n845), .B(A[620]), .Z(n3259) );
  AND U3668 ( .A(n3262), .B(n3263), .Z(n845) );
  NANDN U3669 ( .A(B[619]), .B(n3264), .Z(n3263) );
  NANDN U3670 ( .A(A[619]), .B(n849), .Z(n3264) );
  NANDN U3671 ( .A(n849), .B(A[619]), .Z(n3262) );
  AND U3672 ( .A(n3265), .B(n3266), .Z(n849) );
  NANDN U3673 ( .A(B[618]), .B(n3267), .Z(n3266) );
  NANDN U3674 ( .A(A[618]), .B(n851), .Z(n3267) );
  NANDN U3675 ( .A(n851), .B(A[618]), .Z(n3265) );
  AND U3676 ( .A(n3268), .B(n3269), .Z(n851) );
  NANDN U3677 ( .A(B[617]), .B(n3270), .Z(n3269) );
  NANDN U3678 ( .A(A[617]), .B(n853), .Z(n3270) );
  NANDN U3679 ( .A(n853), .B(A[617]), .Z(n3268) );
  AND U3680 ( .A(n3271), .B(n3272), .Z(n853) );
  NANDN U3681 ( .A(B[616]), .B(n3273), .Z(n3272) );
  NANDN U3682 ( .A(A[616]), .B(n855), .Z(n3273) );
  NANDN U3683 ( .A(n855), .B(A[616]), .Z(n3271) );
  AND U3684 ( .A(n3274), .B(n3275), .Z(n855) );
  NANDN U3685 ( .A(B[615]), .B(n3276), .Z(n3275) );
  NANDN U3686 ( .A(A[615]), .B(n857), .Z(n3276) );
  NANDN U3687 ( .A(n857), .B(A[615]), .Z(n3274) );
  AND U3688 ( .A(n3277), .B(n3278), .Z(n857) );
  NANDN U3689 ( .A(B[614]), .B(n3279), .Z(n3278) );
  NANDN U3690 ( .A(A[614]), .B(n859), .Z(n3279) );
  NANDN U3691 ( .A(n859), .B(A[614]), .Z(n3277) );
  AND U3692 ( .A(n3280), .B(n3281), .Z(n859) );
  NANDN U3693 ( .A(B[613]), .B(n3282), .Z(n3281) );
  NANDN U3694 ( .A(A[613]), .B(n861), .Z(n3282) );
  NANDN U3695 ( .A(n861), .B(A[613]), .Z(n3280) );
  AND U3696 ( .A(n3283), .B(n3284), .Z(n861) );
  NANDN U3697 ( .A(B[612]), .B(n3285), .Z(n3284) );
  NANDN U3698 ( .A(A[612]), .B(n863), .Z(n3285) );
  NANDN U3699 ( .A(n863), .B(A[612]), .Z(n3283) );
  AND U3700 ( .A(n3286), .B(n3287), .Z(n863) );
  NANDN U3701 ( .A(B[611]), .B(n3288), .Z(n3287) );
  NANDN U3702 ( .A(A[611]), .B(n865), .Z(n3288) );
  NANDN U3703 ( .A(n865), .B(A[611]), .Z(n3286) );
  AND U3704 ( .A(n3289), .B(n3290), .Z(n865) );
  NANDN U3705 ( .A(B[610]), .B(n3291), .Z(n3290) );
  NANDN U3706 ( .A(A[610]), .B(n867), .Z(n3291) );
  NANDN U3707 ( .A(n867), .B(A[610]), .Z(n3289) );
  AND U3708 ( .A(n3292), .B(n3293), .Z(n867) );
  NANDN U3709 ( .A(B[609]), .B(n3294), .Z(n3293) );
  NANDN U3710 ( .A(A[609]), .B(n871), .Z(n3294) );
  NANDN U3711 ( .A(n871), .B(A[609]), .Z(n3292) );
  AND U3712 ( .A(n3295), .B(n3296), .Z(n871) );
  NANDN U3713 ( .A(B[608]), .B(n3297), .Z(n3296) );
  NANDN U3714 ( .A(A[608]), .B(n873), .Z(n3297) );
  NANDN U3715 ( .A(n873), .B(A[608]), .Z(n3295) );
  AND U3716 ( .A(n3298), .B(n3299), .Z(n873) );
  NANDN U3717 ( .A(B[607]), .B(n3300), .Z(n3299) );
  NANDN U3718 ( .A(A[607]), .B(n875), .Z(n3300) );
  NANDN U3719 ( .A(n875), .B(A[607]), .Z(n3298) );
  AND U3720 ( .A(n3301), .B(n3302), .Z(n875) );
  NANDN U3721 ( .A(B[606]), .B(n3303), .Z(n3302) );
  NANDN U3722 ( .A(A[606]), .B(n877), .Z(n3303) );
  NANDN U3723 ( .A(n877), .B(A[606]), .Z(n3301) );
  AND U3724 ( .A(n3304), .B(n3305), .Z(n877) );
  NANDN U3725 ( .A(B[605]), .B(n3306), .Z(n3305) );
  NANDN U3726 ( .A(A[605]), .B(n879), .Z(n3306) );
  NANDN U3727 ( .A(n879), .B(A[605]), .Z(n3304) );
  AND U3728 ( .A(n3307), .B(n3308), .Z(n879) );
  NANDN U3729 ( .A(B[604]), .B(n3309), .Z(n3308) );
  NANDN U3730 ( .A(A[604]), .B(n881), .Z(n3309) );
  NANDN U3731 ( .A(n881), .B(A[604]), .Z(n3307) );
  AND U3732 ( .A(n3310), .B(n3311), .Z(n881) );
  NANDN U3733 ( .A(B[603]), .B(n3312), .Z(n3311) );
  NANDN U3734 ( .A(A[603]), .B(n883), .Z(n3312) );
  NANDN U3735 ( .A(n883), .B(A[603]), .Z(n3310) );
  AND U3736 ( .A(n3313), .B(n3314), .Z(n883) );
  NANDN U3737 ( .A(B[602]), .B(n3315), .Z(n3314) );
  NANDN U3738 ( .A(A[602]), .B(n885), .Z(n3315) );
  NANDN U3739 ( .A(n885), .B(A[602]), .Z(n3313) );
  AND U3740 ( .A(n3316), .B(n3317), .Z(n885) );
  NANDN U3741 ( .A(B[601]), .B(n3318), .Z(n3317) );
  NANDN U3742 ( .A(A[601]), .B(n887), .Z(n3318) );
  NANDN U3743 ( .A(n887), .B(A[601]), .Z(n3316) );
  AND U3744 ( .A(n3319), .B(n3320), .Z(n887) );
  NANDN U3745 ( .A(B[600]), .B(n3321), .Z(n3320) );
  NANDN U3746 ( .A(A[600]), .B(n889), .Z(n3321) );
  NANDN U3747 ( .A(n889), .B(A[600]), .Z(n3319) );
  AND U3748 ( .A(n3322), .B(n3323), .Z(n889) );
  NANDN U3749 ( .A(B[599]), .B(n3324), .Z(n3323) );
  NANDN U3750 ( .A(A[599]), .B(n895), .Z(n3324) );
  NANDN U3751 ( .A(n895), .B(A[599]), .Z(n3322) );
  AND U3752 ( .A(n3325), .B(n3326), .Z(n895) );
  NANDN U3753 ( .A(B[598]), .B(n3327), .Z(n3326) );
  NANDN U3754 ( .A(A[598]), .B(n897), .Z(n3327) );
  NANDN U3755 ( .A(n897), .B(A[598]), .Z(n3325) );
  AND U3756 ( .A(n3328), .B(n3329), .Z(n897) );
  NANDN U3757 ( .A(B[597]), .B(n3330), .Z(n3329) );
  NANDN U3758 ( .A(A[597]), .B(n899), .Z(n3330) );
  NANDN U3759 ( .A(n899), .B(A[597]), .Z(n3328) );
  AND U3760 ( .A(n3331), .B(n3332), .Z(n899) );
  NANDN U3761 ( .A(B[596]), .B(n3333), .Z(n3332) );
  NANDN U3762 ( .A(A[596]), .B(n901), .Z(n3333) );
  NANDN U3763 ( .A(n901), .B(A[596]), .Z(n3331) );
  AND U3764 ( .A(n3334), .B(n3335), .Z(n901) );
  NANDN U3765 ( .A(B[595]), .B(n3336), .Z(n3335) );
  NANDN U3766 ( .A(A[595]), .B(n903), .Z(n3336) );
  NANDN U3767 ( .A(n903), .B(A[595]), .Z(n3334) );
  AND U3768 ( .A(n3337), .B(n3338), .Z(n903) );
  NANDN U3769 ( .A(B[594]), .B(n3339), .Z(n3338) );
  NANDN U3770 ( .A(A[594]), .B(n905), .Z(n3339) );
  NANDN U3771 ( .A(n905), .B(A[594]), .Z(n3337) );
  AND U3772 ( .A(n3340), .B(n3341), .Z(n905) );
  NANDN U3773 ( .A(B[593]), .B(n3342), .Z(n3341) );
  NANDN U3774 ( .A(A[593]), .B(n907), .Z(n3342) );
  NANDN U3775 ( .A(n907), .B(A[593]), .Z(n3340) );
  AND U3776 ( .A(n3343), .B(n3344), .Z(n907) );
  NANDN U3777 ( .A(B[592]), .B(n3345), .Z(n3344) );
  NANDN U3778 ( .A(A[592]), .B(n909), .Z(n3345) );
  NANDN U3779 ( .A(n909), .B(A[592]), .Z(n3343) );
  AND U3780 ( .A(n3346), .B(n3347), .Z(n909) );
  NANDN U3781 ( .A(B[591]), .B(n3348), .Z(n3347) );
  NANDN U3782 ( .A(A[591]), .B(n911), .Z(n3348) );
  NANDN U3783 ( .A(n911), .B(A[591]), .Z(n3346) );
  AND U3784 ( .A(n3349), .B(n3350), .Z(n911) );
  NANDN U3785 ( .A(B[590]), .B(n3351), .Z(n3350) );
  NANDN U3786 ( .A(A[590]), .B(n913), .Z(n3351) );
  NANDN U3787 ( .A(n913), .B(A[590]), .Z(n3349) );
  AND U3788 ( .A(n3352), .B(n3353), .Z(n913) );
  NANDN U3789 ( .A(B[589]), .B(n3354), .Z(n3353) );
  NANDN U3790 ( .A(A[589]), .B(n917), .Z(n3354) );
  NANDN U3791 ( .A(n917), .B(A[589]), .Z(n3352) );
  AND U3792 ( .A(n3355), .B(n3356), .Z(n917) );
  NANDN U3793 ( .A(B[588]), .B(n3357), .Z(n3356) );
  NANDN U3794 ( .A(A[588]), .B(n919), .Z(n3357) );
  NANDN U3795 ( .A(n919), .B(A[588]), .Z(n3355) );
  AND U3796 ( .A(n3358), .B(n3359), .Z(n919) );
  NANDN U3797 ( .A(B[587]), .B(n3360), .Z(n3359) );
  NANDN U3798 ( .A(A[587]), .B(n921), .Z(n3360) );
  NANDN U3799 ( .A(n921), .B(A[587]), .Z(n3358) );
  AND U3800 ( .A(n3361), .B(n3362), .Z(n921) );
  NANDN U3801 ( .A(B[586]), .B(n3363), .Z(n3362) );
  NANDN U3802 ( .A(A[586]), .B(n923), .Z(n3363) );
  NANDN U3803 ( .A(n923), .B(A[586]), .Z(n3361) );
  AND U3804 ( .A(n3364), .B(n3365), .Z(n923) );
  NANDN U3805 ( .A(B[585]), .B(n3366), .Z(n3365) );
  NANDN U3806 ( .A(A[585]), .B(n925), .Z(n3366) );
  NANDN U3807 ( .A(n925), .B(A[585]), .Z(n3364) );
  AND U3808 ( .A(n3367), .B(n3368), .Z(n925) );
  NANDN U3809 ( .A(B[584]), .B(n3369), .Z(n3368) );
  NANDN U3810 ( .A(A[584]), .B(n927), .Z(n3369) );
  NANDN U3811 ( .A(n927), .B(A[584]), .Z(n3367) );
  AND U3812 ( .A(n3370), .B(n3371), .Z(n927) );
  NANDN U3813 ( .A(B[583]), .B(n3372), .Z(n3371) );
  NANDN U3814 ( .A(A[583]), .B(n929), .Z(n3372) );
  NANDN U3815 ( .A(n929), .B(A[583]), .Z(n3370) );
  AND U3816 ( .A(n3373), .B(n3374), .Z(n929) );
  NANDN U3817 ( .A(B[582]), .B(n3375), .Z(n3374) );
  NANDN U3818 ( .A(A[582]), .B(n931), .Z(n3375) );
  NANDN U3819 ( .A(n931), .B(A[582]), .Z(n3373) );
  AND U3820 ( .A(n3376), .B(n3377), .Z(n931) );
  NANDN U3821 ( .A(B[581]), .B(n3378), .Z(n3377) );
  NANDN U3822 ( .A(A[581]), .B(n933), .Z(n3378) );
  NANDN U3823 ( .A(n933), .B(A[581]), .Z(n3376) );
  AND U3824 ( .A(n3379), .B(n3380), .Z(n933) );
  NANDN U3825 ( .A(B[580]), .B(n3381), .Z(n3380) );
  NANDN U3826 ( .A(A[580]), .B(n935), .Z(n3381) );
  NANDN U3827 ( .A(n935), .B(A[580]), .Z(n3379) );
  AND U3828 ( .A(n3382), .B(n3383), .Z(n935) );
  NANDN U3829 ( .A(B[579]), .B(n3384), .Z(n3383) );
  NANDN U3830 ( .A(A[579]), .B(n939), .Z(n3384) );
  NANDN U3831 ( .A(n939), .B(A[579]), .Z(n3382) );
  AND U3832 ( .A(n3385), .B(n3386), .Z(n939) );
  NANDN U3833 ( .A(B[578]), .B(n3387), .Z(n3386) );
  NANDN U3834 ( .A(A[578]), .B(n941), .Z(n3387) );
  NANDN U3835 ( .A(n941), .B(A[578]), .Z(n3385) );
  AND U3836 ( .A(n3388), .B(n3389), .Z(n941) );
  NANDN U3837 ( .A(B[577]), .B(n3390), .Z(n3389) );
  NANDN U3838 ( .A(A[577]), .B(n943), .Z(n3390) );
  NANDN U3839 ( .A(n943), .B(A[577]), .Z(n3388) );
  AND U3840 ( .A(n3391), .B(n3392), .Z(n943) );
  NANDN U3841 ( .A(B[576]), .B(n3393), .Z(n3392) );
  NANDN U3842 ( .A(A[576]), .B(n945), .Z(n3393) );
  NANDN U3843 ( .A(n945), .B(A[576]), .Z(n3391) );
  AND U3844 ( .A(n3394), .B(n3395), .Z(n945) );
  NANDN U3845 ( .A(B[575]), .B(n3396), .Z(n3395) );
  NANDN U3846 ( .A(A[575]), .B(n947), .Z(n3396) );
  NANDN U3847 ( .A(n947), .B(A[575]), .Z(n3394) );
  AND U3848 ( .A(n3397), .B(n3398), .Z(n947) );
  NANDN U3849 ( .A(B[574]), .B(n3399), .Z(n3398) );
  NANDN U3850 ( .A(A[574]), .B(n949), .Z(n3399) );
  NANDN U3851 ( .A(n949), .B(A[574]), .Z(n3397) );
  AND U3852 ( .A(n3400), .B(n3401), .Z(n949) );
  NANDN U3853 ( .A(B[573]), .B(n3402), .Z(n3401) );
  NANDN U3854 ( .A(A[573]), .B(n951), .Z(n3402) );
  NANDN U3855 ( .A(n951), .B(A[573]), .Z(n3400) );
  AND U3856 ( .A(n3403), .B(n3404), .Z(n951) );
  NANDN U3857 ( .A(B[572]), .B(n3405), .Z(n3404) );
  NANDN U3858 ( .A(A[572]), .B(n953), .Z(n3405) );
  NANDN U3859 ( .A(n953), .B(A[572]), .Z(n3403) );
  AND U3860 ( .A(n3406), .B(n3407), .Z(n953) );
  NANDN U3861 ( .A(B[571]), .B(n3408), .Z(n3407) );
  NANDN U3862 ( .A(A[571]), .B(n955), .Z(n3408) );
  NANDN U3863 ( .A(n955), .B(A[571]), .Z(n3406) );
  AND U3864 ( .A(n3409), .B(n3410), .Z(n955) );
  NANDN U3865 ( .A(B[570]), .B(n3411), .Z(n3410) );
  NANDN U3866 ( .A(A[570]), .B(n957), .Z(n3411) );
  NANDN U3867 ( .A(n957), .B(A[570]), .Z(n3409) );
  AND U3868 ( .A(n3412), .B(n3413), .Z(n957) );
  NANDN U3869 ( .A(B[569]), .B(n3414), .Z(n3413) );
  NANDN U3870 ( .A(A[569]), .B(n961), .Z(n3414) );
  NANDN U3871 ( .A(n961), .B(A[569]), .Z(n3412) );
  AND U3872 ( .A(n3415), .B(n3416), .Z(n961) );
  NANDN U3873 ( .A(B[568]), .B(n3417), .Z(n3416) );
  NANDN U3874 ( .A(A[568]), .B(n963), .Z(n3417) );
  NANDN U3875 ( .A(n963), .B(A[568]), .Z(n3415) );
  AND U3876 ( .A(n3418), .B(n3419), .Z(n963) );
  NANDN U3877 ( .A(B[567]), .B(n3420), .Z(n3419) );
  NANDN U3878 ( .A(A[567]), .B(n965), .Z(n3420) );
  NANDN U3879 ( .A(n965), .B(A[567]), .Z(n3418) );
  AND U3880 ( .A(n3421), .B(n3422), .Z(n965) );
  NANDN U3881 ( .A(B[566]), .B(n3423), .Z(n3422) );
  NANDN U3882 ( .A(A[566]), .B(n967), .Z(n3423) );
  NANDN U3883 ( .A(n967), .B(A[566]), .Z(n3421) );
  AND U3884 ( .A(n3424), .B(n3425), .Z(n967) );
  NANDN U3885 ( .A(B[565]), .B(n3426), .Z(n3425) );
  NANDN U3886 ( .A(A[565]), .B(n969), .Z(n3426) );
  NANDN U3887 ( .A(n969), .B(A[565]), .Z(n3424) );
  AND U3888 ( .A(n3427), .B(n3428), .Z(n969) );
  NANDN U3889 ( .A(B[564]), .B(n3429), .Z(n3428) );
  NANDN U3890 ( .A(A[564]), .B(n971), .Z(n3429) );
  NANDN U3891 ( .A(n971), .B(A[564]), .Z(n3427) );
  AND U3892 ( .A(n3430), .B(n3431), .Z(n971) );
  NANDN U3893 ( .A(B[563]), .B(n3432), .Z(n3431) );
  NANDN U3894 ( .A(A[563]), .B(n973), .Z(n3432) );
  NANDN U3895 ( .A(n973), .B(A[563]), .Z(n3430) );
  AND U3896 ( .A(n3433), .B(n3434), .Z(n973) );
  NANDN U3897 ( .A(B[562]), .B(n3435), .Z(n3434) );
  NANDN U3898 ( .A(A[562]), .B(n975), .Z(n3435) );
  NANDN U3899 ( .A(n975), .B(A[562]), .Z(n3433) );
  AND U3900 ( .A(n3436), .B(n3437), .Z(n975) );
  NANDN U3901 ( .A(B[561]), .B(n3438), .Z(n3437) );
  NANDN U3902 ( .A(A[561]), .B(n977), .Z(n3438) );
  NANDN U3903 ( .A(n977), .B(A[561]), .Z(n3436) );
  AND U3904 ( .A(n3439), .B(n3440), .Z(n977) );
  NANDN U3905 ( .A(B[560]), .B(n3441), .Z(n3440) );
  NANDN U3906 ( .A(A[560]), .B(n979), .Z(n3441) );
  NANDN U3907 ( .A(n979), .B(A[560]), .Z(n3439) );
  AND U3908 ( .A(n3442), .B(n3443), .Z(n979) );
  NANDN U3909 ( .A(B[559]), .B(n3444), .Z(n3443) );
  NANDN U3910 ( .A(A[559]), .B(n983), .Z(n3444) );
  NANDN U3911 ( .A(n983), .B(A[559]), .Z(n3442) );
  AND U3912 ( .A(n3445), .B(n3446), .Z(n983) );
  NANDN U3913 ( .A(B[558]), .B(n3447), .Z(n3446) );
  NANDN U3914 ( .A(A[558]), .B(n985), .Z(n3447) );
  NANDN U3915 ( .A(n985), .B(A[558]), .Z(n3445) );
  AND U3916 ( .A(n3448), .B(n3449), .Z(n985) );
  NANDN U3917 ( .A(B[557]), .B(n3450), .Z(n3449) );
  NANDN U3918 ( .A(A[557]), .B(n987), .Z(n3450) );
  NANDN U3919 ( .A(n987), .B(A[557]), .Z(n3448) );
  AND U3920 ( .A(n3451), .B(n3452), .Z(n987) );
  NANDN U3921 ( .A(B[556]), .B(n3453), .Z(n3452) );
  NANDN U3922 ( .A(A[556]), .B(n989), .Z(n3453) );
  NANDN U3923 ( .A(n989), .B(A[556]), .Z(n3451) );
  AND U3924 ( .A(n3454), .B(n3455), .Z(n989) );
  NANDN U3925 ( .A(B[555]), .B(n3456), .Z(n3455) );
  NANDN U3926 ( .A(A[555]), .B(n991), .Z(n3456) );
  NANDN U3927 ( .A(n991), .B(A[555]), .Z(n3454) );
  AND U3928 ( .A(n3457), .B(n3458), .Z(n991) );
  NANDN U3929 ( .A(B[554]), .B(n3459), .Z(n3458) );
  NANDN U3930 ( .A(A[554]), .B(n993), .Z(n3459) );
  NANDN U3931 ( .A(n993), .B(A[554]), .Z(n3457) );
  AND U3932 ( .A(n3460), .B(n3461), .Z(n993) );
  NANDN U3933 ( .A(B[553]), .B(n3462), .Z(n3461) );
  NANDN U3934 ( .A(A[553]), .B(n995), .Z(n3462) );
  NANDN U3935 ( .A(n995), .B(A[553]), .Z(n3460) );
  AND U3936 ( .A(n3463), .B(n3464), .Z(n995) );
  NANDN U3937 ( .A(B[552]), .B(n3465), .Z(n3464) );
  NANDN U3938 ( .A(A[552]), .B(n997), .Z(n3465) );
  NANDN U3939 ( .A(n997), .B(A[552]), .Z(n3463) );
  AND U3940 ( .A(n3466), .B(n3467), .Z(n997) );
  NANDN U3941 ( .A(B[551]), .B(n3468), .Z(n3467) );
  NANDN U3942 ( .A(A[551]), .B(n999), .Z(n3468) );
  NANDN U3943 ( .A(n999), .B(A[551]), .Z(n3466) );
  AND U3944 ( .A(n3469), .B(n3470), .Z(n999) );
  NANDN U3945 ( .A(B[550]), .B(n3471), .Z(n3470) );
  NANDN U3946 ( .A(A[550]), .B(n1001), .Z(n3471) );
  NANDN U3947 ( .A(n1001), .B(A[550]), .Z(n3469) );
  AND U3948 ( .A(n3472), .B(n3473), .Z(n1001) );
  NANDN U3949 ( .A(B[549]), .B(n3474), .Z(n3473) );
  NANDN U3950 ( .A(A[549]), .B(n1005), .Z(n3474) );
  NANDN U3951 ( .A(n1005), .B(A[549]), .Z(n3472) );
  AND U3952 ( .A(n3475), .B(n3476), .Z(n1005) );
  NANDN U3953 ( .A(B[548]), .B(n3477), .Z(n3476) );
  NANDN U3954 ( .A(A[548]), .B(n1007), .Z(n3477) );
  NANDN U3955 ( .A(n1007), .B(A[548]), .Z(n3475) );
  AND U3956 ( .A(n3478), .B(n3479), .Z(n1007) );
  NANDN U3957 ( .A(B[547]), .B(n3480), .Z(n3479) );
  NANDN U3958 ( .A(A[547]), .B(n1009), .Z(n3480) );
  NANDN U3959 ( .A(n1009), .B(A[547]), .Z(n3478) );
  AND U3960 ( .A(n3481), .B(n3482), .Z(n1009) );
  NANDN U3961 ( .A(B[546]), .B(n3483), .Z(n3482) );
  NANDN U3962 ( .A(A[546]), .B(n1011), .Z(n3483) );
  NANDN U3963 ( .A(n1011), .B(A[546]), .Z(n3481) );
  AND U3964 ( .A(n3484), .B(n3485), .Z(n1011) );
  NANDN U3965 ( .A(B[545]), .B(n3486), .Z(n3485) );
  NANDN U3966 ( .A(A[545]), .B(n1013), .Z(n3486) );
  NANDN U3967 ( .A(n1013), .B(A[545]), .Z(n3484) );
  AND U3968 ( .A(n3487), .B(n3488), .Z(n1013) );
  NANDN U3969 ( .A(B[544]), .B(n3489), .Z(n3488) );
  NANDN U3970 ( .A(A[544]), .B(n1015), .Z(n3489) );
  NANDN U3971 ( .A(n1015), .B(A[544]), .Z(n3487) );
  AND U3972 ( .A(n3490), .B(n3491), .Z(n1015) );
  NANDN U3973 ( .A(B[543]), .B(n3492), .Z(n3491) );
  NANDN U3974 ( .A(A[543]), .B(n1017), .Z(n3492) );
  NANDN U3975 ( .A(n1017), .B(A[543]), .Z(n3490) );
  AND U3976 ( .A(n3493), .B(n3494), .Z(n1017) );
  NANDN U3977 ( .A(B[542]), .B(n3495), .Z(n3494) );
  NANDN U3978 ( .A(A[542]), .B(n1019), .Z(n3495) );
  NANDN U3979 ( .A(n1019), .B(A[542]), .Z(n3493) );
  AND U3980 ( .A(n3496), .B(n3497), .Z(n1019) );
  NANDN U3981 ( .A(B[541]), .B(n3498), .Z(n3497) );
  NANDN U3982 ( .A(A[541]), .B(n1021), .Z(n3498) );
  NANDN U3983 ( .A(n1021), .B(A[541]), .Z(n3496) );
  AND U3984 ( .A(n3499), .B(n3500), .Z(n1021) );
  NANDN U3985 ( .A(B[540]), .B(n3501), .Z(n3500) );
  NANDN U3986 ( .A(A[540]), .B(n1023), .Z(n3501) );
  NANDN U3987 ( .A(n1023), .B(A[540]), .Z(n3499) );
  AND U3988 ( .A(n3502), .B(n3503), .Z(n1023) );
  NANDN U3989 ( .A(B[539]), .B(n3504), .Z(n3503) );
  NANDN U3990 ( .A(A[539]), .B(n1027), .Z(n3504) );
  NANDN U3991 ( .A(n1027), .B(A[539]), .Z(n3502) );
  AND U3992 ( .A(n3505), .B(n3506), .Z(n1027) );
  NANDN U3993 ( .A(B[538]), .B(n3507), .Z(n3506) );
  NANDN U3994 ( .A(A[538]), .B(n1029), .Z(n3507) );
  NANDN U3995 ( .A(n1029), .B(A[538]), .Z(n3505) );
  AND U3996 ( .A(n3508), .B(n3509), .Z(n1029) );
  NANDN U3997 ( .A(B[537]), .B(n3510), .Z(n3509) );
  NANDN U3998 ( .A(A[537]), .B(n1031), .Z(n3510) );
  NANDN U3999 ( .A(n1031), .B(A[537]), .Z(n3508) );
  AND U4000 ( .A(n3511), .B(n3512), .Z(n1031) );
  NANDN U4001 ( .A(B[536]), .B(n3513), .Z(n3512) );
  NANDN U4002 ( .A(A[536]), .B(n1033), .Z(n3513) );
  NANDN U4003 ( .A(n1033), .B(A[536]), .Z(n3511) );
  AND U4004 ( .A(n3514), .B(n3515), .Z(n1033) );
  NANDN U4005 ( .A(B[535]), .B(n3516), .Z(n3515) );
  NANDN U4006 ( .A(A[535]), .B(n1035), .Z(n3516) );
  NANDN U4007 ( .A(n1035), .B(A[535]), .Z(n3514) );
  AND U4008 ( .A(n3517), .B(n3518), .Z(n1035) );
  NANDN U4009 ( .A(B[534]), .B(n3519), .Z(n3518) );
  NANDN U4010 ( .A(A[534]), .B(n1037), .Z(n3519) );
  NANDN U4011 ( .A(n1037), .B(A[534]), .Z(n3517) );
  AND U4012 ( .A(n3520), .B(n3521), .Z(n1037) );
  NANDN U4013 ( .A(B[533]), .B(n3522), .Z(n3521) );
  NANDN U4014 ( .A(A[533]), .B(n1039), .Z(n3522) );
  NANDN U4015 ( .A(n1039), .B(A[533]), .Z(n3520) );
  AND U4016 ( .A(n3523), .B(n3524), .Z(n1039) );
  NANDN U4017 ( .A(B[532]), .B(n3525), .Z(n3524) );
  NANDN U4018 ( .A(A[532]), .B(n1041), .Z(n3525) );
  NANDN U4019 ( .A(n1041), .B(A[532]), .Z(n3523) );
  AND U4020 ( .A(n3526), .B(n3527), .Z(n1041) );
  NANDN U4021 ( .A(B[531]), .B(n3528), .Z(n3527) );
  NANDN U4022 ( .A(A[531]), .B(n1043), .Z(n3528) );
  NANDN U4023 ( .A(n1043), .B(A[531]), .Z(n3526) );
  AND U4024 ( .A(n3529), .B(n3530), .Z(n1043) );
  NANDN U4025 ( .A(B[530]), .B(n3531), .Z(n3530) );
  NANDN U4026 ( .A(A[530]), .B(n1045), .Z(n3531) );
  NANDN U4027 ( .A(n1045), .B(A[530]), .Z(n3529) );
  AND U4028 ( .A(n3532), .B(n3533), .Z(n1045) );
  NANDN U4029 ( .A(B[529]), .B(n3534), .Z(n3533) );
  NANDN U4030 ( .A(A[529]), .B(n1049), .Z(n3534) );
  NANDN U4031 ( .A(n1049), .B(A[529]), .Z(n3532) );
  AND U4032 ( .A(n3535), .B(n3536), .Z(n1049) );
  NANDN U4033 ( .A(B[528]), .B(n3537), .Z(n3536) );
  NANDN U4034 ( .A(A[528]), .B(n1051), .Z(n3537) );
  NANDN U4035 ( .A(n1051), .B(A[528]), .Z(n3535) );
  AND U4036 ( .A(n3538), .B(n3539), .Z(n1051) );
  NANDN U4037 ( .A(B[527]), .B(n3540), .Z(n3539) );
  NANDN U4038 ( .A(A[527]), .B(n1053), .Z(n3540) );
  NANDN U4039 ( .A(n1053), .B(A[527]), .Z(n3538) );
  AND U4040 ( .A(n3541), .B(n3542), .Z(n1053) );
  NANDN U4041 ( .A(B[526]), .B(n3543), .Z(n3542) );
  NANDN U4042 ( .A(A[526]), .B(n1055), .Z(n3543) );
  NANDN U4043 ( .A(n1055), .B(A[526]), .Z(n3541) );
  AND U4044 ( .A(n3544), .B(n3545), .Z(n1055) );
  NANDN U4045 ( .A(B[525]), .B(n3546), .Z(n3545) );
  NANDN U4046 ( .A(A[525]), .B(n1057), .Z(n3546) );
  NANDN U4047 ( .A(n1057), .B(A[525]), .Z(n3544) );
  AND U4048 ( .A(n3547), .B(n3548), .Z(n1057) );
  NANDN U4049 ( .A(B[524]), .B(n3549), .Z(n3548) );
  NANDN U4050 ( .A(A[524]), .B(n1059), .Z(n3549) );
  NANDN U4051 ( .A(n1059), .B(A[524]), .Z(n3547) );
  AND U4052 ( .A(n3550), .B(n3551), .Z(n1059) );
  NANDN U4053 ( .A(B[523]), .B(n3552), .Z(n3551) );
  NANDN U4054 ( .A(A[523]), .B(n1061), .Z(n3552) );
  NANDN U4055 ( .A(n1061), .B(A[523]), .Z(n3550) );
  AND U4056 ( .A(n3553), .B(n3554), .Z(n1061) );
  NANDN U4057 ( .A(B[522]), .B(n3555), .Z(n3554) );
  NANDN U4058 ( .A(A[522]), .B(n1063), .Z(n3555) );
  NANDN U4059 ( .A(n1063), .B(A[522]), .Z(n3553) );
  AND U4060 ( .A(n3556), .B(n3557), .Z(n1063) );
  NANDN U4061 ( .A(B[521]), .B(n3558), .Z(n3557) );
  NANDN U4062 ( .A(A[521]), .B(n1065), .Z(n3558) );
  NANDN U4063 ( .A(n1065), .B(A[521]), .Z(n3556) );
  AND U4064 ( .A(n3559), .B(n3560), .Z(n1065) );
  NANDN U4065 ( .A(B[520]), .B(n3561), .Z(n3560) );
  NANDN U4066 ( .A(A[520]), .B(n1067), .Z(n3561) );
  NANDN U4067 ( .A(n1067), .B(A[520]), .Z(n3559) );
  AND U4068 ( .A(n3562), .B(n3563), .Z(n1067) );
  NANDN U4069 ( .A(B[519]), .B(n3564), .Z(n3563) );
  NANDN U4070 ( .A(A[519]), .B(n1071), .Z(n3564) );
  NANDN U4071 ( .A(n1071), .B(A[519]), .Z(n3562) );
  AND U4072 ( .A(n3565), .B(n3566), .Z(n1071) );
  NANDN U4073 ( .A(B[518]), .B(n3567), .Z(n3566) );
  NANDN U4074 ( .A(A[518]), .B(n1073), .Z(n3567) );
  NANDN U4075 ( .A(n1073), .B(A[518]), .Z(n3565) );
  AND U4076 ( .A(n3568), .B(n3569), .Z(n1073) );
  NANDN U4077 ( .A(B[517]), .B(n3570), .Z(n3569) );
  NANDN U4078 ( .A(A[517]), .B(n1075), .Z(n3570) );
  NANDN U4079 ( .A(n1075), .B(A[517]), .Z(n3568) );
  AND U4080 ( .A(n3571), .B(n3572), .Z(n1075) );
  NANDN U4081 ( .A(B[516]), .B(n3573), .Z(n3572) );
  NANDN U4082 ( .A(A[516]), .B(n1077), .Z(n3573) );
  NANDN U4083 ( .A(n1077), .B(A[516]), .Z(n3571) );
  AND U4084 ( .A(n3574), .B(n3575), .Z(n1077) );
  NANDN U4085 ( .A(B[515]), .B(n3576), .Z(n3575) );
  NANDN U4086 ( .A(A[515]), .B(n1079), .Z(n3576) );
  NANDN U4087 ( .A(n1079), .B(A[515]), .Z(n3574) );
  AND U4088 ( .A(n3577), .B(n3578), .Z(n1079) );
  NANDN U4089 ( .A(B[514]), .B(n3579), .Z(n3578) );
  NANDN U4090 ( .A(A[514]), .B(n1081), .Z(n3579) );
  NANDN U4091 ( .A(n1081), .B(A[514]), .Z(n3577) );
  AND U4092 ( .A(n3580), .B(n3581), .Z(n1081) );
  NANDN U4093 ( .A(B[513]), .B(n3582), .Z(n3581) );
  NANDN U4094 ( .A(A[513]), .B(n1083), .Z(n3582) );
  NANDN U4095 ( .A(n1083), .B(A[513]), .Z(n3580) );
  AND U4096 ( .A(n3583), .B(n3584), .Z(n1083) );
  NANDN U4097 ( .A(B[512]), .B(n3585), .Z(n3584) );
  NANDN U4098 ( .A(A[512]), .B(n1085), .Z(n3585) );
  NANDN U4099 ( .A(n1085), .B(A[512]), .Z(n3583) );
  AND U4100 ( .A(n3586), .B(n3587), .Z(n1085) );
  NANDN U4101 ( .A(B[511]), .B(n3588), .Z(n3587) );
  NANDN U4102 ( .A(A[511]), .B(n1087), .Z(n3588) );
  NANDN U4103 ( .A(n1087), .B(A[511]), .Z(n3586) );
  AND U4104 ( .A(n3589), .B(n3590), .Z(n1087) );
  NANDN U4105 ( .A(B[510]), .B(n3591), .Z(n3590) );
  NANDN U4106 ( .A(A[510]), .B(n1089), .Z(n3591) );
  NANDN U4107 ( .A(n1089), .B(A[510]), .Z(n3589) );
  AND U4108 ( .A(n3592), .B(n3593), .Z(n1089) );
  NANDN U4109 ( .A(B[509]), .B(n3594), .Z(n3593) );
  NANDN U4110 ( .A(A[509]), .B(n1093), .Z(n3594) );
  NANDN U4111 ( .A(n1093), .B(A[509]), .Z(n3592) );
  AND U4112 ( .A(n3595), .B(n3596), .Z(n1093) );
  NANDN U4113 ( .A(B[508]), .B(n3597), .Z(n3596) );
  NANDN U4114 ( .A(A[508]), .B(n1095), .Z(n3597) );
  NANDN U4115 ( .A(n1095), .B(A[508]), .Z(n3595) );
  AND U4116 ( .A(n3598), .B(n3599), .Z(n1095) );
  NANDN U4117 ( .A(B[507]), .B(n3600), .Z(n3599) );
  NANDN U4118 ( .A(A[507]), .B(n1097), .Z(n3600) );
  NANDN U4119 ( .A(n1097), .B(A[507]), .Z(n3598) );
  AND U4120 ( .A(n3601), .B(n3602), .Z(n1097) );
  NANDN U4121 ( .A(B[506]), .B(n3603), .Z(n3602) );
  NANDN U4122 ( .A(A[506]), .B(n1099), .Z(n3603) );
  NANDN U4123 ( .A(n1099), .B(A[506]), .Z(n3601) );
  AND U4124 ( .A(n3604), .B(n3605), .Z(n1099) );
  NANDN U4125 ( .A(B[505]), .B(n3606), .Z(n3605) );
  NANDN U4126 ( .A(A[505]), .B(n1101), .Z(n3606) );
  NANDN U4127 ( .A(n1101), .B(A[505]), .Z(n3604) );
  AND U4128 ( .A(n3607), .B(n3608), .Z(n1101) );
  NANDN U4129 ( .A(B[504]), .B(n3609), .Z(n3608) );
  NANDN U4130 ( .A(A[504]), .B(n1103), .Z(n3609) );
  NANDN U4131 ( .A(n1103), .B(A[504]), .Z(n3607) );
  AND U4132 ( .A(n3610), .B(n3611), .Z(n1103) );
  NANDN U4133 ( .A(B[503]), .B(n3612), .Z(n3611) );
  NANDN U4134 ( .A(A[503]), .B(n1105), .Z(n3612) );
  NANDN U4135 ( .A(n1105), .B(A[503]), .Z(n3610) );
  AND U4136 ( .A(n3613), .B(n3614), .Z(n1105) );
  NANDN U4137 ( .A(B[502]), .B(n3615), .Z(n3614) );
  NANDN U4138 ( .A(A[502]), .B(n1107), .Z(n3615) );
  NANDN U4139 ( .A(n1107), .B(A[502]), .Z(n3613) );
  AND U4140 ( .A(n3616), .B(n3617), .Z(n1107) );
  NANDN U4141 ( .A(B[501]), .B(n3618), .Z(n3617) );
  NANDN U4142 ( .A(A[501]), .B(n1109), .Z(n3618) );
  NANDN U4143 ( .A(n1109), .B(A[501]), .Z(n3616) );
  AND U4144 ( .A(n3619), .B(n3620), .Z(n1109) );
  NANDN U4145 ( .A(B[500]), .B(n3621), .Z(n3620) );
  NANDN U4146 ( .A(A[500]), .B(n1111), .Z(n3621) );
  NANDN U4147 ( .A(n1111), .B(A[500]), .Z(n3619) );
  AND U4148 ( .A(n3622), .B(n3623), .Z(n1111) );
  NANDN U4149 ( .A(B[499]), .B(n3624), .Z(n3623) );
  NANDN U4150 ( .A(A[499]), .B(n1117), .Z(n3624) );
  NANDN U4151 ( .A(n1117), .B(A[499]), .Z(n3622) );
  AND U4152 ( .A(n3625), .B(n3626), .Z(n1117) );
  NANDN U4153 ( .A(B[498]), .B(n3627), .Z(n3626) );
  NANDN U4154 ( .A(A[498]), .B(n1119), .Z(n3627) );
  NANDN U4155 ( .A(n1119), .B(A[498]), .Z(n3625) );
  AND U4156 ( .A(n3628), .B(n3629), .Z(n1119) );
  NANDN U4157 ( .A(B[497]), .B(n3630), .Z(n3629) );
  NANDN U4158 ( .A(A[497]), .B(n1121), .Z(n3630) );
  NANDN U4159 ( .A(n1121), .B(A[497]), .Z(n3628) );
  AND U4160 ( .A(n3631), .B(n3632), .Z(n1121) );
  NANDN U4161 ( .A(B[496]), .B(n3633), .Z(n3632) );
  NANDN U4162 ( .A(A[496]), .B(n1123), .Z(n3633) );
  NANDN U4163 ( .A(n1123), .B(A[496]), .Z(n3631) );
  AND U4164 ( .A(n3634), .B(n3635), .Z(n1123) );
  NANDN U4165 ( .A(B[495]), .B(n3636), .Z(n3635) );
  NANDN U4166 ( .A(A[495]), .B(n1125), .Z(n3636) );
  NANDN U4167 ( .A(n1125), .B(A[495]), .Z(n3634) );
  AND U4168 ( .A(n3637), .B(n3638), .Z(n1125) );
  NANDN U4169 ( .A(B[494]), .B(n3639), .Z(n3638) );
  NANDN U4170 ( .A(A[494]), .B(n1127), .Z(n3639) );
  NANDN U4171 ( .A(n1127), .B(A[494]), .Z(n3637) );
  AND U4172 ( .A(n3640), .B(n3641), .Z(n1127) );
  NANDN U4173 ( .A(B[493]), .B(n3642), .Z(n3641) );
  NANDN U4174 ( .A(A[493]), .B(n1129), .Z(n3642) );
  NANDN U4175 ( .A(n1129), .B(A[493]), .Z(n3640) );
  AND U4176 ( .A(n3643), .B(n3644), .Z(n1129) );
  NANDN U4177 ( .A(B[492]), .B(n3645), .Z(n3644) );
  NANDN U4178 ( .A(A[492]), .B(n1131), .Z(n3645) );
  NANDN U4179 ( .A(n1131), .B(A[492]), .Z(n3643) );
  AND U4180 ( .A(n3646), .B(n3647), .Z(n1131) );
  NANDN U4181 ( .A(B[491]), .B(n3648), .Z(n3647) );
  NANDN U4182 ( .A(A[491]), .B(n1133), .Z(n3648) );
  NANDN U4183 ( .A(n1133), .B(A[491]), .Z(n3646) );
  AND U4184 ( .A(n3649), .B(n3650), .Z(n1133) );
  NANDN U4185 ( .A(B[490]), .B(n3651), .Z(n3650) );
  NANDN U4186 ( .A(A[490]), .B(n1135), .Z(n3651) );
  NANDN U4187 ( .A(n1135), .B(A[490]), .Z(n3649) );
  AND U4188 ( .A(n3652), .B(n3653), .Z(n1135) );
  NANDN U4189 ( .A(B[489]), .B(n3654), .Z(n3653) );
  NANDN U4190 ( .A(A[489]), .B(n1139), .Z(n3654) );
  NANDN U4191 ( .A(n1139), .B(A[489]), .Z(n3652) );
  AND U4192 ( .A(n3655), .B(n3656), .Z(n1139) );
  NANDN U4193 ( .A(B[488]), .B(n3657), .Z(n3656) );
  NANDN U4194 ( .A(A[488]), .B(n1141), .Z(n3657) );
  NANDN U4195 ( .A(n1141), .B(A[488]), .Z(n3655) );
  AND U4196 ( .A(n3658), .B(n3659), .Z(n1141) );
  NANDN U4197 ( .A(B[487]), .B(n3660), .Z(n3659) );
  NANDN U4198 ( .A(A[487]), .B(n1143), .Z(n3660) );
  NANDN U4199 ( .A(n1143), .B(A[487]), .Z(n3658) );
  AND U4200 ( .A(n3661), .B(n3662), .Z(n1143) );
  NANDN U4201 ( .A(B[486]), .B(n3663), .Z(n3662) );
  NANDN U4202 ( .A(A[486]), .B(n1145), .Z(n3663) );
  NANDN U4203 ( .A(n1145), .B(A[486]), .Z(n3661) );
  AND U4204 ( .A(n3664), .B(n3665), .Z(n1145) );
  NANDN U4205 ( .A(B[485]), .B(n3666), .Z(n3665) );
  NANDN U4206 ( .A(A[485]), .B(n1147), .Z(n3666) );
  NANDN U4207 ( .A(n1147), .B(A[485]), .Z(n3664) );
  AND U4208 ( .A(n3667), .B(n3668), .Z(n1147) );
  NANDN U4209 ( .A(B[484]), .B(n3669), .Z(n3668) );
  NANDN U4210 ( .A(A[484]), .B(n1149), .Z(n3669) );
  NANDN U4211 ( .A(n1149), .B(A[484]), .Z(n3667) );
  AND U4212 ( .A(n3670), .B(n3671), .Z(n1149) );
  NANDN U4213 ( .A(B[483]), .B(n3672), .Z(n3671) );
  NANDN U4214 ( .A(A[483]), .B(n1151), .Z(n3672) );
  NANDN U4215 ( .A(n1151), .B(A[483]), .Z(n3670) );
  AND U4216 ( .A(n3673), .B(n3674), .Z(n1151) );
  NANDN U4217 ( .A(B[482]), .B(n3675), .Z(n3674) );
  NANDN U4218 ( .A(A[482]), .B(n1153), .Z(n3675) );
  NANDN U4219 ( .A(n1153), .B(A[482]), .Z(n3673) );
  AND U4220 ( .A(n3676), .B(n3677), .Z(n1153) );
  NANDN U4221 ( .A(B[481]), .B(n3678), .Z(n3677) );
  NANDN U4222 ( .A(A[481]), .B(n1155), .Z(n3678) );
  NANDN U4223 ( .A(n1155), .B(A[481]), .Z(n3676) );
  AND U4224 ( .A(n3679), .B(n3680), .Z(n1155) );
  NANDN U4225 ( .A(B[480]), .B(n3681), .Z(n3680) );
  NANDN U4226 ( .A(A[480]), .B(n1157), .Z(n3681) );
  NANDN U4227 ( .A(n1157), .B(A[480]), .Z(n3679) );
  AND U4228 ( .A(n3682), .B(n3683), .Z(n1157) );
  NANDN U4229 ( .A(B[479]), .B(n3684), .Z(n3683) );
  NANDN U4230 ( .A(A[479]), .B(n1161), .Z(n3684) );
  NANDN U4231 ( .A(n1161), .B(A[479]), .Z(n3682) );
  AND U4232 ( .A(n3685), .B(n3686), .Z(n1161) );
  NANDN U4233 ( .A(B[478]), .B(n3687), .Z(n3686) );
  NANDN U4234 ( .A(A[478]), .B(n1163), .Z(n3687) );
  NANDN U4235 ( .A(n1163), .B(A[478]), .Z(n3685) );
  AND U4236 ( .A(n3688), .B(n3689), .Z(n1163) );
  NANDN U4237 ( .A(B[477]), .B(n3690), .Z(n3689) );
  NANDN U4238 ( .A(A[477]), .B(n1165), .Z(n3690) );
  NANDN U4239 ( .A(n1165), .B(A[477]), .Z(n3688) );
  AND U4240 ( .A(n3691), .B(n3692), .Z(n1165) );
  NANDN U4241 ( .A(B[476]), .B(n3693), .Z(n3692) );
  NANDN U4242 ( .A(A[476]), .B(n1167), .Z(n3693) );
  NANDN U4243 ( .A(n1167), .B(A[476]), .Z(n3691) );
  AND U4244 ( .A(n3694), .B(n3695), .Z(n1167) );
  NANDN U4245 ( .A(B[475]), .B(n3696), .Z(n3695) );
  NANDN U4246 ( .A(A[475]), .B(n1169), .Z(n3696) );
  NANDN U4247 ( .A(n1169), .B(A[475]), .Z(n3694) );
  AND U4248 ( .A(n3697), .B(n3698), .Z(n1169) );
  NANDN U4249 ( .A(B[474]), .B(n3699), .Z(n3698) );
  NANDN U4250 ( .A(A[474]), .B(n1171), .Z(n3699) );
  NANDN U4251 ( .A(n1171), .B(A[474]), .Z(n3697) );
  AND U4252 ( .A(n3700), .B(n3701), .Z(n1171) );
  NANDN U4253 ( .A(B[473]), .B(n3702), .Z(n3701) );
  NANDN U4254 ( .A(A[473]), .B(n1173), .Z(n3702) );
  NANDN U4255 ( .A(n1173), .B(A[473]), .Z(n3700) );
  AND U4256 ( .A(n3703), .B(n3704), .Z(n1173) );
  NANDN U4257 ( .A(B[472]), .B(n3705), .Z(n3704) );
  NANDN U4258 ( .A(A[472]), .B(n1175), .Z(n3705) );
  NANDN U4259 ( .A(n1175), .B(A[472]), .Z(n3703) );
  AND U4260 ( .A(n3706), .B(n3707), .Z(n1175) );
  NANDN U4261 ( .A(B[471]), .B(n3708), .Z(n3707) );
  NANDN U4262 ( .A(A[471]), .B(n1177), .Z(n3708) );
  NANDN U4263 ( .A(n1177), .B(A[471]), .Z(n3706) );
  AND U4264 ( .A(n3709), .B(n3710), .Z(n1177) );
  NANDN U4265 ( .A(B[470]), .B(n3711), .Z(n3710) );
  NANDN U4266 ( .A(A[470]), .B(n1179), .Z(n3711) );
  NANDN U4267 ( .A(n1179), .B(A[470]), .Z(n3709) );
  AND U4268 ( .A(n3712), .B(n3713), .Z(n1179) );
  NANDN U4269 ( .A(B[469]), .B(n3714), .Z(n3713) );
  NANDN U4270 ( .A(A[469]), .B(n1183), .Z(n3714) );
  NANDN U4271 ( .A(n1183), .B(A[469]), .Z(n3712) );
  AND U4272 ( .A(n3715), .B(n3716), .Z(n1183) );
  NANDN U4273 ( .A(B[468]), .B(n3717), .Z(n3716) );
  NANDN U4274 ( .A(A[468]), .B(n1185), .Z(n3717) );
  NANDN U4275 ( .A(n1185), .B(A[468]), .Z(n3715) );
  AND U4276 ( .A(n3718), .B(n3719), .Z(n1185) );
  NANDN U4277 ( .A(B[467]), .B(n3720), .Z(n3719) );
  NANDN U4278 ( .A(A[467]), .B(n1187), .Z(n3720) );
  NANDN U4279 ( .A(n1187), .B(A[467]), .Z(n3718) );
  AND U4280 ( .A(n3721), .B(n3722), .Z(n1187) );
  NANDN U4281 ( .A(B[466]), .B(n3723), .Z(n3722) );
  NANDN U4282 ( .A(A[466]), .B(n1189), .Z(n3723) );
  NANDN U4283 ( .A(n1189), .B(A[466]), .Z(n3721) );
  AND U4284 ( .A(n3724), .B(n3725), .Z(n1189) );
  NANDN U4285 ( .A(B[465]), .B(n3726), .Z(n3725) );
  NANDN U4286 ( .A(A[465]), .B(n1191), .Z(n3726) );
  NANDN U4287 ( .A(n1191), .B(A[465]), .Z(n3724) );
  AND U4288 ( .A(n3727), .B(n3728), .Z(n1191) );
  NANDN U4289 ( .A(B[464]), .B(n3729), .Z(n3728) );
  NANDN U4290 ( .A(A[464]), .B(n1193), .Z(n3729) );
  NANDN U4291 ( .A(n1193), .B(A[464]), .Z(n3727) );
  AND U4292 ( .A(n3730), .B(n3731), .Z(n1193) );
  NANDN U4293 ( .A(B[463]), .B(n3732), .Z(n3731) );
  NANDN U4294 ( .A(A[463]), .B(n1195), .Z(n3732) );
  NANDN U4295 ( .A(n1195), .B(A[463]), .Z(n3730) );
  AND U4296 ( .A(n3733), .B(n3734), .Z(n1195) );
  NANDN U4297 ( .A(B[462]), .B(n3735), .Z(n3734) );
  NANDN U4298 ( .A(A[462]), .B(n1197), .Z(n3735) );
  NANDN U4299 ( .A(n1197), .B(A[462]), .Z(n3733) );
  AND U4300 ( .A(n3736), .B(n3737), .Z(n1197) );
  NANDN U4301 ( .A(B[461]), .B(n3738), .Z(n3737) );
  NANDN U4302 ( .A(A[461]), .B(n1199), .Z(n3738) );
  NANDN U4303 ( .A(n1199), .B(A[461]), .Z(n3736) );
  AND U4304 ( .A(n3739), .B(n3740), .Z(n1199) );
  NANDN U4305 ( .A(B[460]), .B(n3741), .Z(n3740) );
  NANDN U4306 ( .A(A[460]), .B(n1201), .Z(n3741) );
  NANDN U4307 ( .A(n1201), .B(A[460]), .Z(n3739) );
  AND U4308 ( .A(n3742), .B(n3743), .Z(n1201) );
  NANDN U4309 ( .A(B[459]), .B(n3744), .Z(n3743) );
  NANDN U4310 ( .A(A[459]), .B(n1205), .Z(n3744) );
  NANDN U4311 ( .A(n1205), .B(A[459]), .Z(n3742) );
  AND U4312 ( .A(n3745), .B(n3746), .Z(n1205) );
  NANDN U4313 ( .A(B[458]), .B(n3747), .Z(n3746) );
  NANDN U4314 ( .A(A[458]), .B(n1207), .Z(n3747) );
  NANDN U4315 ( .A(n1207), .B(A[458]), .Z(n3745) );
  AND U4316 ( .A(n3748), .B(n3749), .Z(n1207) );
  NANDN U4317 ( .A(B[457]), .B(n3750), .Z(n3749) );
  NANDN U4318 ( .A(A[457]), .B(n1209), .Z(n3750) );
  NANDN U4319 ( .A(n1209), .B(A[457]), .Z(n3748) );
  AND U4320 ( .A(n3751), .B(n3752), .Z(n1209) );
  NANDN U4321 ( .A(B[456]), .B(n3753), .Z(n3752) );
  NANDN U4322 ( .A(A[456]), .B(n1211), .Z(n3753) );
  NANDN U4323 ( .A(n1211), .B(A[456]), .Z(n3751) );
  AND U4324 ( .A(n3754), .B(n3755), .Z(n1211) );
  NANDN U4325 ( .A(B[455]), .B(n3756), .Z(n3755) );
  NANDN U4326 ( .A(A[455]), .B(n1213), .Z(n3756) );
  NANDN U4327 ( .A(n1213), .B(A[455]), .Z(n3754) );
  AND U4328 ( .A(n3757), .B(n3758), .Z(n1213) );
  NANDN U4329 ( .A(B[454]), .B(n3759), .Z(n3758) );
  NANDN U4330 ( .A(A[454]), .B(n1215), .Z(n3759) );
  NANDN U4331 ( .A(n1215), .B(A[454]), .Z(n3757) );
  AND U4332 ( .A(n3760), .B(n3761), .Z(n1215) );
  NANDN U4333 ( .A(B[453]), .B(n3762), .Z(n3761) );
  NANDN U4334 ( .A(A[453]), .B(n1217), .Z(n3762) );
  NANDN U4335 ( .A(n1217), .B(A[453]), .Z(n3760) );
  AND U4336 ( .A(n3763), .B(n3764), .Z(n1217) );
  NANDN U4337 ( .A(B[452]), .B(n3765), .Z(n3764) );
  NANDN U4338 ( .A(A[452]), .B(n1219), .Z(n3765) );
  NANDN U4339 ( .A(n1219), .B(A[452]), .Z(n3763) );
  AND U4340 ( .A(n3766), .B(n3767), .Z(n1219) );
  NANDN U4341 ( .A(B[451]), .B(n3768), .Z(n3767) );
  NANDN U4342 ( .A(A[451]), .B(n1221), .Z(n3768) );
  NANDN U4343 ( .A(n1221), .B(A[451]), .Z(n3766) );
  AND U4344 ( .A(n3769), .B(n3770), .Z(n1221) );
  NANDN U4345 ( .A(B[450]), .B(n3771), .Z(n3770) );
  NANDN U4346 ( .A(A[450]), .B(n1223), .Z(n3771) );
  NANDN U4347 ( .A(n1223), .B(A[450]), .Z(n3769) );
  AND U4348 ( .A(n3772), .B(n3773), .Z(n1223) );
  NANDN U4349 ( .A(B[449]), .B(n3774), .Z(n3773) );
  NANDN U4350 ( .A(A[449]), .B(n1227), .Z(n3774) );
  NANDN U4351 ( .A(n1227), .B(A[449]), .Z(n3772) );
  AND U4352 ( .A(n3775), .B(n3776), .Z(n1227) );
  NANDN U4353 ( .A(B[448]), .B(n3777), .Z(n3776) );
  NANDN U4354 ( .A(A[448]), .B(n1229), .Z(n3777) );
  NANDN U4355 ( .A(n1229), .B(A[448]), .Z(n3775) );
  AND U4356 ( .A(n3778), .B(n3779), .Z(n1229) );
  NANDN U4357 ( .A(B[447]), .B(n3780), .Z(n3779) );
  NANDN U4358 ( .A(A[447]), .B(n1231), .Z(n3780) );
  NANDN U4359 ( .A(n1231), .B(A[447]), .Z(n3778) );
  AND U4360 ( .A(n3781), .B(n3782), .Z(n1231) );
  NANDN U4361 ( .A(B[446]), .B(n3783), .Z(n3782) );
  NANDN U4362 ( .A(A[446]), .B(n1233), .Z(n3783) );
  NANDN U4363 ( .A(n1233), .B(A[446]), .Z(n3781) );
  AND U4364 ( .A(n3784), .B(n3785), .Z(n1233) );
  NANDN U4365 ( .A(B[445]), .B(n3786), .Z(n3785) );
  NANDN U4366 ( .A(A[445]), .B(n1235), .Z(n3786) );
  NANDN U4367 ( .A(n1235), .B(A[445]), .Z(n3784) );
  AND U4368 ( .A(n3787), .B(n3788), .Z(n1235) );
  NANDN U4369 ( .A(B[444]), .B(n3789), .Z(n3788) );
  NANDN U4370 ( .A(A[444]), .B(n1237), .Z(n3789) );
  NANDN U4371 ( .A(n1237), .B(A[444]), .Z(n3787) );
  AND U4372 ( .A(n3790), .B(n3791), .Z(n1237) );
  NANDN U4373 ( .A(B[443]), .B(n3792), .Z(n3791) );
  NANDN U4374 ( .A(A[443]), .B(n1239), .Z(n3792) );
  NANDN U4375 ( .A(n1239), .B(A[443]), .Z(n3790) );
  AND U4376 ( .A(n3793), .B(n3794), .Z(n1239) );
  NANDN U4377 ( .A(B[442]), .B(n3795), .Z(n3794) );
  NANDN U4378 ( .A(A[442]), .B(n1241), .Z(n3795) );
  NANDN U4379 ( .A(n1241), .B(A[442]), .Z(n3793) );
  AND U4380 ( .A(n3796), .B(n3797), .Z(n1241) );
  NANDN U4381 ( .A(B[441]), .B(n3798), .Z(n3797) );
  NANDN U4382 ( .A(A[441]), .B(n1243), .Z(n3798) );
  NANDN U4383 ( .A(n1243), .B(A[441]), .Z(n3796) );
  AND U4384 ( .A(n3799), .B(n3800), .Z(n1243) );
  NANDN U4385 ( .A(B[440]), .B(n3801), .Z(n3800) );
  NANDN U4386 ( .A(A[440]), .B(n1245), .Z(n3801) );
  NANDN U4387 ( .A(n1245), .B(A[440]), .Z(n3799) );
  AND U4388 ( .A(n3802), .B(n3803), .Z(n1245) );
  NANDN U4389 ( .A(B[439]), .B(n3804), .Z(n3803) );
  NANDN U4390 ( .A(A[439]), .B(n1249), .Z(n3804) );
  NANDN U4391 ( .A(n1249), .B(A[439]), .Z(n3802) );
  AND U4392 ( .A(n3805), .B(n3806), .Z(n1249) );
  NANDN U4393 ( .A(B[438]), .B(n3807), .Z(n3806) );
  NANDN U4394 ( .A(A[438]), .B(n1251), .Z(n3807) );
  NANDN U4395 ( .A(n1251), .B(A[438]), .Z(n3805) );
  AND U4396 ( .A(n3808), .B(n3809), .Z(n1251) );
  NANDN U4397 ( .A(B[437]), .B(n3810), .Z(n3809) );
  NANDN U4398 ( .A(A[437]), .B(n1253), .Z(n3810) );
  NANDN U4399 ( .A(n1253), .B(A[437]), .Z(n3808) );
  AND U4400 ( .A(n3811), .B(n3812), .Z(n1253) );
  NANDN U4401 ( .A(B[436]), .B(n3813), .Z(n3812) );
  NANDN U4402 ( .A(A[436]), .B(n1255), .Z(n3813) );
  NANDN U4403 ( .A(n1255), .B(A[436]), .Z(n3811) );
  AND U4404 ( .A(n3814), .B(n3815), .Z(n1255) );
  NANDN U4405 ( .A(B[435]), .B(n3816), .Z(n3815) );
  NANDN U4406 ( .A(A[435]), .B(n1257), .Z(n3816) );
  NANDN U4407 ( .A(n1257), .B(A[435]), .Z(n3814) );
  AND U4408 ( .A(n3817), .B(n3818), .Z(n1257) );
  NANDN U4409 ( .A(B[434]), .B(n3819), .Z(n3818) );
  NANDN U4410 ( .A(A[434]), .B(n1259), .Z(n3819) );
  NANDN U4411 ( .A(n1259), .B(A[434]), .Z(n3817) );
  AND U4412 ( .A(n3820), .B(n3821), .Z(n1259) );
  NANDN U4413 ( .A(B[433]), .B(n3822), .Z(n3821) );
  NANDN U4414 ( .A(A[433]), .B(n1261), .Z(n3822) );
  NANDN U4415 ( .A(n1261), .B(A[433]), .Z(n3820) );
  AND U4416 ( .A(n3823), .B(n3824), .Z(n1261) );
  NANDN U4417 ( .A(B[432]), .B(n3825), .Z(n3824) );
  NANDN U4418 ( .A(A[432]), .B(n1263), .Z(n3825) );
  NANDN U4419 ( .A(n1263), .B(A[432]), .Z(n3823) );
  AND U4420 ( .A(n3826), .B(n3827), .Z(n1263) );
  NANDN U4421 ( .A(B[431]), .B(n3828), .Z(n3827) );
  NANDN U4422 ( .A(A[431]), .B(n1265), .Z(n3828) );
  NANDN U4423 ( .A(n1265), .B(A[431]), .Z(n3826) );
  AND U4424 ( .A(n3829), .B(n3830), .Z(n1265) );
  NANDN U4425 ( .A(B[430]), .B(n3831), .Z(n3830) );
  NANDN U4426 ( .A(A[430]), .B(n1267), .Z(n3831) );
  NANDN U4427 ( .A(n1267), .B(A[430]), .Z(n3829) );
  AND U4428 ( .A(n3832), .B(n3833), .Z(n1267) );
  NANDN U4429 ( .A(B[429]), .B(n3834), .Z(n3833) );
  NANDN U4430 ( .A(A[429]), .B(n1271), .Z(n3834) );
  NANDN U4431 ( .A(n1271), .B(A[429]), .Z(n3832) );
  AND U4432 ( .A(n3835), .B(n3836), .Z(n1271) );
  NANDN U4433 ( .A(B[428]), .B(n3837), .Z(n3836) );
  NANDN U4434 ( .A(A[428]), .B(n1273), .Z(n3837) );
  NANDN U4435 ( .A(n1273), .B(A[428]), .Z(n3835) );
  AND U4436 ( .A(n3838), .B(n3839), .Z(n1273) );
  NANDN U4437 ( .A(B[427]), .B(n3840), .Z(n3839) );
  NANDN U4438 ( .A(A[427]), .B(n1275), .Z(n3840) );
  NANDN U4439 ( .A(n1275), .B(A[427]), .Z(n3838) );
  AND U4440 ( .A(n3841), .B(n3842), .Z(n1275) );
  NANDN U4441 ( .A(B[426]), .B(n3843), .Z(n3842) );
  NANDN U4442 ( .A(A[426]), .B(n1277), .Z(n3843) );
  NANDN U4443 ( .A(n1277), .B(A[426]), .Z(n3841) );
  AND U4444 ( .A(n3844), .B(n3845), .Z(n1277) );
  NANDN U4445 ( .A(B[425]), .B(n3846), .Z(n3845) );
  NANDN U4446 ( .A(A[425]), .B(n1279), .Z(n3846) );
  NANDN U4447 ( .A(n1279), .B(A[425]), .Z(n3844) );
  AND U4448 ( .A(n3847), .B(n3848), .Z(n1279) );
  NANDN U4449 ( .A(B[424]), .B(n3849), .Z(n3848) );
  NANDN U4450 ( .A(A[424]), .B(n1281), .Z(n3849) );
  NANDN U4451 ( .A(n1281), .B(A[424]), .Z(n3847) );
  AND U4452 ( .A(n3850), .B(n3851), .Z(n1281) );
  NANDN U4453 ( .A(B[423]), .B(n3852), .Z(n3851) );
  NANDN U4454 ( .A(A[423]), .B(n1283), .Z(n3852) );
  NANDN U4455 ( .A(n1283), .B(A[423]), .Z(n3850) );
  AND U4456 ( .A(n3853), .B(n3854), .Z(n1283) );
  NANDN U4457 ( .A(B[422]), .B(n3855), .Z(n3854) );
  NANDN U4458 ( .A(A[422]), .B(n1285), .Z(n3855) );
  NANDN U4459 ( .A(n1285), .B(A[422]), .Z(n3853) );
  AND U4460 ( .A(n3856), .B(n3857), .Z(n1285) );
  NANDN U4461 ( .A(B[421]), .B(n3858), .Z(n3857) );
  NANDN U4462 ( .A(A[421]), .B(n1287), .Z(n3858) );
  NANDN U4463 ( .A(n1287), .B(A[421]), .Z(n3856) );
  AND U4464 ( .A(n3859), .B(n3860), .Z(n1287) );
  NANDN U4465 ( .A(B[420]), .B(n3861), .Z(n3860) );
  NANDN U4466 ( .A(A[420]), .B(n1289), .Z(n3861) );
  NANDN U4467 ( .A(n1289), .B(A[420]), .Z(n3859) );
  AND U4468 ( .A(n3862), .B(n3863), .Z(n1289) );
  NANDN U4469 ( .A(B[419]), .B(n3864), .Z(n3863) );
  NANDN U4470 ( .A(A[419]), .B(n1293), .Z(n3864) );
  NANDN U4471 ( .A(n1293), .B(A[419]), .Z(n3862) );
  AND U4472 ( .A(n3865), .B(n3866), .Z(n1293) );
  NANDN U4473 ( .A(B[418]), .B(n3867), .Z(n3866) );
  NANDN U4474 ( .A(A[418]), .B(n1295), .Z(n3867) );
  NANDN U4475 ( .A(n1295), .B(A[418]), .Z(n3865) );
  AND U4476 ( .A(n3868), .B(n3869), .Z(n1295) );
  NANDN U4477 ( .A(B[417]), .B(n3870), .Z(n3869) );
  NANDN U4478 ( .A(A[417]), .B(n1297), .Z(n3870) );
  NANDN U4479 ( .A(n1297), .B(A[417]), .Z(n3868) );
  AND U4480 ( .A(n3871), .B(n3872), .Z(n1297) );
  NANDN U4481 ( .A(B[416]), .B(n3873), .Z(n3872) );
  NANDN U4482 ( .A(A[416]), .B(n1299), .Z(n3873) );
  NANDN U4483 ( .A(n1299), .B(A[416]), .Z(n3871) );
  AND U4484 ( .A(n3874), .B(n3875), .Z(n1299) );
  NANDN U4485 ( .A(B[415]), .B(n3876), .Z(n3875) );
  NANDN U4486 ( .A(A[415]), .B(n1301), .Z(n3876) );
  NANDN U4487 ( .A(n1301), .B(A[415]), .Z(n3874) );
  AND U4488 ( .A(n3877), .B(n3878), .Z(n1301) );
  NANDN U4489 ( .A(B[414]), .B(n3879), .Z(n3878) );
  NANDN U4490 ( .A(A[414]), .B(n1303), .Z(n3879) );
  NANDN U4491 ( .A(n1303), .B(A[414]), .Z(n3877) );
  AND U4492 ( .A(n3880), .B(n3881), .Z(n1303) );
  NANDN U4493 ( .A(B[413]), .B(n3882), .Z(n3881) );
  NANDN U4494 ( .A(A[413]), .B(n1305), .Z(n3882) );
  NANDN U4495 ( .A(n1305), .B(A[413]), .Z(n3880) );
  AND U4496 ( .A(n3883), .B(n3884), .Z(n1305) );
  NANDN U4497 ( .A(B[412]), .B(n3885), .Z(n3884) );
  NANDN U4498 ( .A(A[412]), .B(n1307), .Z(n3885) );
  NANDN U4499 ( .A(n1307), .B(A[412]), .Z(n3883) );
  AND U4500 ( .A(n3886), .B(n3887), .Z(n1307) );
  NANDN U4501 ( .A(B[411]), .B(n3888), .Z(n3887) );
  NANDN U4502 ( .A(A[411]), .B(n1309), .Z(n3888) );
  NANDN U4503 ( .A(n1309), .B(A[411]), .Z(n3886) );
  AND U4504 ( .A(n3889), .B(n3890), .Z(n1309) );
  NANDN U4505 ( .A(B[410]), .B(n3891), .Z(n3890) );
  NANDN U4506 ( .A(A[410]), .B(n1311), .Z(n3891) );
  NANDN U4507 ( .A(n1311), .B(A[410]), .Z(n3889) );
  AND U4508 ( .A(n3892), .B(n3893), .Z(n1311) );
  NANDN U4509 ( .A(B[409]), .B(n3894), .Z(n3893) );
  NANDN U4510 ( .A(A[409]), .B(n1315), .Z(n3894) );
  NANDN U4511 ( .A(n1315), .B(A[409]), .Z(n3892) );
  AND U4512 ( .A(n3895), .B(n3896), .Z(n1315) );
  NANDN U4513 ( .A(B[408]), .B(n3897), .Z(n3896) );
  NANDN U4514 ( .A(A[408]), .B(n1317), .Z(n3897) );
  NANDN U4515 ( .A(n1317), .B(A[408]), .Z(n3895) );
  AND U4516 ( .A(n3898), .B(n3899), .Z(n1317) );
  NANDN U4517 ( .A(B[407]), .B(n3900), .Z(n3899) );
  NANDN U4518 ( .A(A[407]), .B(n1319), .Z(n3900) );
  NANDN U4519 ( .A(n1319), .B(A[407]), .Z(n3898) );
  AND U4520 ( .A(n3901), .B(n3902), .Z(n1319) );
  NANDN U4521 ( .A(B[406]), .B(n3903), .Z(n3902) );
  NANDN U4522 ( .A(A[406]), .B(n1321), .Z(n3903) );
  NANDN U4523 ( .A(n1321), .B(A[406]), .Z(n3901) );
  AND U4524 ( .A(n3904), .B(n3905), .Z(n1321) );
  NANDN U4525 ( .A(B[405]), .B(n3906), .Z(n3905) );
  NANDN U4526 ( .A(A[405]), .B(n1323), .Z(n3906) );
  NANDN U4527 ( .A(n1323), .B(A[405]), .Z(n3904) );
  AND U4528 ( .A(n3907), .B(n3908), .Z(n1323) );
  NANDN U4529 ( .A(B[404]), .B(n3909), .Z(n3908) );
  NANDN U4530 ( .A(A[404]), .B(n1325), .Z(n3909) );
  NANDN U4531 ( .A(n1325), .B(A[404]), .Z(n3907) );
  AND U4532 ( .A(n3910), .B(n3911), .Z(n1325) );
  NANDN U4533 ( .A(B[403]), .B(n3912), .Z(n3911) );
  NANDN U4534 ( .A(A[403]), .B(n1327), .Z(n3912) );
  NANDN U4535 ( .A(n1327), .B(A[403]), .Z(n3910) );
  AND U4536 ( .A(n3913), .B(n3914), .Z(n1327) );
  NANDN U4537 ( .A(B[402]), .B(n3915), .Z(n3914) );
  NANDN U4538 ( .A(A[402]), .B(n1329), .Z(n3915) );
  NANDN U4539 ( .A(n1329), .B(A[402]), .Z(n3913) );
  AND U4540 ( .A(n3916), .B(n3917), .Z(n1329) );
  NANDN U4541 ( .A(B[401]), .B(n3918), .Z(n3917) );
  NANDN U4542 ( .A(A[401]), .B(n1331), .Z(n3918) );
  NANDN U4543 ( .A(n1331), .B(A[401]), .Z(n3916) );
  AND U4544 ( .A(n3919), .B(n3920), .Z(n1331) );
  NANDN U4545 ( .A(B[400]), .B(n3921), .Z(n3920) );
  NANDN U4546 ( .A(A[400]), .B(n1333), .Z(n3921) );
  NANDN U4547 ( .A(n1333), .B(A[400]), .Z(n3919) );
  AND U4548 ( .A(n3922), .B(n3923), .Z(n1333) );
  NANDN U4549 ( .A(B[399]), .B(n3924), .Z(n3923) );
  NANDN U4550 ( .A(A[399]), .B(n1339), .Z(n3924) );
  NANDN U4551 ( .A(n1339), .B(A[399]), .Z(n3922) );
  AND U4552 ( .A(n3925), .B(n3926), .Z(n1339) );
  NANDN U4553 ( .A(B[398]), .B(n3927), .Z(n3926) );
  NANDN U4554 ( .A(A[398]), .B(n1341), .Z(n3927) );
  NANDN U4555 ( .A(n1341), .B(A[398]), .Z(n3925) );
  AND U4556 ( .A(n3928), .B(n3929), .Z(n1341) );
  NANDN U4557 ( .A(B[397]), .B(n3930), .Z(n3929) );
  NANDN U4558 ( .A(A[397]), .B(n1343), .Z(n3930) );
  NANDN U4559 ( .A(n1343), .B(A[397]), .Z(n3928) );
  AND U4560 ( .A(n3931), .B(n3932), .Z(n1343) );
  NANDN U4561 ( .A(B[396]), .B(n3933), .Z(n3932) );
  NANDN U4562 ( .A(A[396]), .B(n1345), .Z(n3933) );
  NANDN U4563 ( .A(n1345), .B(A[396]), .Z(n3931) );
  AND U4564 ( .A(n3934), .B(n3935), .Z(n1345) );
  NANDN U4565 ( .A(B[395]), .B(n3936), .Z(n3935) );
  NANDN U4566 ( .A(A[395]), .B(n1347), .Z(n3936) );
  NANDN U4567 ( .A(n1347), .B(A[395]), .Z(n3934) );
  AND U4568 ( .A(n3937), .B(n3938), .Z(n1347) );
  NANDN U4569 ( .A(B[394]), .B(n3939), .Z(n3938) );
  NANDN U4570 ( .A(A[394]), .B(n1349), .Z(n3939) );
  NANDN U4571 ( .A(n1349), .B(A[394]), .Z(n3937) );
  AND U4572 ( .A(n3940), .B(n3941), .Z(n1349) );
  NANDN U4573 ( .A(B[393]), .B(n3942), .Z(n3941) );
  NANDN U4574 ( .A(A[393]), .B(n1351), .Z(n3942) );
  NANDN U4575 ( .A(n1351), .B(A[393]), .Z(n3940) );
  AND U4576 ( .A(n3943), .B(n3944), .Z(n1351) );
  NANDN U4577 ( .A(B[392]), .B(n3945), .Z(n3944) );
  NANDN U4578 ( .A(A[392]), .B(n1353), .Z(n3945) );
  NANDN U4579 ( .A(n1353), .B(A[392]), .Z(n3943) );
  AND U4580 ( .A(n3946), .B(n3947), .Z(n1353) );
  NANDN U4581 ( .A(B[391]), .B(n3948), .Z(n3947) );
  NANDN U4582 ( .A(A[391]), .B(n1355), .Z(n3948) );
  NANDN U4583 ( .A(n1355), .B(A[391]), .Z(n3946) );
  AND U4584 ( .A(n3949), .B(n3950), .Z(n1355) );
  NANDN U4585 ( .A(B[390]), .B(n3951), .Z(n3950) );
  NANDN U4586 ( .A(A[390]), .B(n1357), .Z(n3951) );
  NANDN U4587 ( .A(n1357), .B(A[390]), .Z(n3949) );
  AND U4588 ( .A(n3952), .B(n3953), .Z(n1357) );
  NANDN U4589 ( .A(B[389]), .B(n3954), .Z(n3953) );
  NANDN U4590 ( .A(A[389]), .B(n1361), .Z(n3954) );
  NANDN U4591 ( .A(n1361), .B(A[389]), .Z(n3952) );
  AND U4592 ( .A(n3955), .B(n3956), .Z(n1361) );
  NANDN U4593 ( .A(B[388]), .B(n3957), .Z(n3956) );
  NANDN U4594 ( .A(A[388]), .B(n1363), .Z(n3957) );
  NANDN U4595 ( .A(n1363), .B(A[388]), .Z(n3955) );
  AND U4596 ( .A(n3958), .B(n3959), .Z(n1363) );
  NANDN U4597 ( .A(B[387]), .B(n3960), .Z(n3959) );
  NANDN U4598 ( .A(A[387]), .B(n1365), .Z(n3960) );
  NANDN U4599 ( .A(n1365), .B(A[387]), .Z(n3958) );
  AND U4600 ( .A(n3961), .B(n3962), .Z(n1365) );
  NANDN U4601 ( .A(B[386]), .B(n3963), .Z(n3962) );
  NANDN U4602 ( .A(A[386]), .B(n1367), .Z(n3963) );
  NANDN U4603 ( .A(n1367), .B(A[386]), .Z(n3961) );
  AND U4604 ( .A(n3964), .B(n3965), .Z(n1367) );
  NANDN U4605 ( .A(B[385]), .B(n3966), .Z(n3965) );
  NANDN U4606 ( .A(A[385]), .B(n1369), .Z(n3966) );
  NANDN U4607 ( .A(n1369), .B(A[385]), .Z(n3964) );
  AND U4608 ( .A(n3967), .B(n3968), .Z(n1369) );
  NANDN U4609 ( .A(B[384]), .B(n3969), .Z(n3968) );
  NANDN U4610 ( .A(A[384]), .B(n1371), .Z(n3969) );
  NANDN U4611 ( .A(n1371), .B(A[384]), .Z(n3967) );
  AND U4612 ( .A(n3970), .B(n3971), .Z(n1371) );
  NANDN U4613 ( .A(B[383]), .B(n3972), .Z(n3971) );
  NANDN U4614 ( .A(A[383]), .B(n1373), .Z(n3972) );
  NANDN U4615 ( .A(n1373), .B(A[383]), .Z(n3970) );
  AND U4616 ( .A(n3973), .B(n3974), .Z(n1373) );
  NANDN U4617 ( .A(B[382]), .B(n3975), .Z(n3974) );
  NANDN U4618 ( .A(A[382]), .B(n1375), .Z(n3975) );
  NANDN U4619 ( .A(n1375), .B(A[382]), .Z(n3973) );
  AND U4620 ( .A(n3976), .B(n3977), .Z(n1375) );
  NANDN U4621 ( .A(B[381]), .B(n3978), .Z(n3977) );
  NANDN U4622 ( .A(A[381]), .B(n1377), .Z(n3978) );
  NANDN U4623 ( .A(n1377), .B(A[381]), .Z(n3976) );
  AND U4624 ( .A(n3979), .B(n3980), .Z(n1377) );
  NANDN U4625 ( .A(B[380]), .B(n3981), .Z(n3980) );
  NANDN U4626 ( .A(A[380]), .B(n1379), .Z(n3981) );
  NANDN U4627 ( .A(n1379), .B(A[380]), .Z(n3979) );
  AND U4628 ( .A(n3982), .B(n3983), .Z(n1379) );
  NANDN U4629 ( .A(B[379]), .B(n3984), .Z(n3983) );
  NANDN U4630 ( .A(A[379]), .B(n1383), .Z(n3984) );
  NANDN U4631 ( .A(n1383), .B(A[379]), .Z(n3982) );
  AND U4632 ( .A(n3985), .B(n3986), .Z(n1383) );
  NANDN U4633 ( .A(B[378]), .B(n3987), .Z(n3986) );
  NANDN U4634 ( .A(A[378]), .B(n1385), .Z(n3987) );
  NANDN U4635 ( .A(n1385), .B(A[378]), .Z(n3985) );
  AND U4636 ( .A(n3988), .B(n3989), .Z(n1385) );
  NANDN U4637 ( .A(B[377]), .B(n3990), .Z(n3989) );
  NANDN U4638 ( .A(A[377]), .B(n1387), .Z(n3990) );
  NANDN U4639 ( .A(n1387), .B(A[377]), .Z(n3988) );
  AND U4640 ( .A(n3991), .B(n3992), .Z(n1387) );
  NANDN U4641 ( .A(B[376]), .B(n3993), .Z(n3992) );
  NANDN U4642 ( .A(A[376]), .B(n1389), .Z(n3993) );
  NANDN U4643 ( .A(n1389), .B(A[376]), .Z(n3991) );
  AND U4644 ( .A(n3994), .B(n3995), .Z(n1389) );
  NANDN U4645 ( .A(B[375]), .B(n3996), .Z(n3995) );
  NANDN U4646 ( .A(A[375]), .B(n1391), .Z(n3996) );
  NANDN U4647 ( .A(n1391), .B(A[375]), .Z(n3994) );
  AND U4648 ( .A(n3997), .B(n3998), .Z(n1391) );
  NANDN U4649 ( .A(B[374]), .B(n3999), .Z(n3998) );
  NANDN U4650 ( .A(A[374]), .B(n1393), .Z(n3999) );
  NANDN U4651 ( .A(n1393), .B(A[374]), .Z(n3997) );
  AND U4652 ( .A(n4000), .B(n4001), .Z(n1393) );
  NANDN U4653 ( .A(B[373]), .B(n4002), .Z(n4001) );
  NANDN U4654 ( .A(A[373]), .B(n1395), .Z(n4002) );
  NANDN U4655 ( .A(n1395), .B(A[373]), .Z(n4000) );
  AND U4656 ( .A(n4003), .B(n4004), .Z(n1395) );
  NANDN U4657 ( .A(B[372]), .B(n4005), .Z(n4004) );
  NANDN U4658 ( .A(A[372]), .B(n1397), .Z(n4005) );
  NANDN U4659 ( .A(n1397), .B(A[372]), .Z(n4003) );
  AND U4660 ( .A(n4006), .B(n4007), .Z(n1397) );
  NANDN U4661 ( .A(B[371]), .B(n4008), .Z(n4007) );
  NANDN U4662 ( .A(A[371]), .B(n1399), .Z(n4008) );
  NANDN U4663 ( .A(n1399), .B(A[371]), .Z(n4006) );
  AND U4664 ( .A(n4009), .B(n4010), .Z(n1399) );
  NANDN U4665 ( .A(B[370]), .B(n4011), .Z(n4010) );
  NANDN U4666 ( .A(A[370]), .B(n1401), .Z(n4011) );
  NANDN U4667 ( .A(n1401), .B(A[370]), .Z(n4009) );
  AND U4668 ( .A(n4012), .B(n4013), .Z(n1401) );
  NANDN U4669 ( .A(B[369]), .B(n4014), .Z(n4013) );
  NANDN U4670 ( .A(A[369]), .B(n1405), .Z(n4014) );
  NANDN U4671 ( .A(n1405), .B(A[369]), .Z(n4012) );
  AND U4672 ( .A(n4015), .B(n4016), .Z(n1405) );
  NANDN U4673 ( .A(B[368]), .B(n4017), .Z(n4016) );
  NANDN U4674 ( .A(A[368]), .B(n1407), .Z(n4017) );
  NANDN U4675 ( .A(n1407), .B(A[368]), .Z(n4015) );
  AND U4676 ( .A(n4018), .B(n4019), .Z(n1407) );
  NANDN U4677 ( .A(B[367]), .B(n4020), .Z(n4019) );
  NANDN U4678 ( .A(A[367]), .B(n1409), .Z(n4020) );
  NANDN U4679 ( .A(n1409), .B(A[367]), .Z(n4018) );
  AND U4680 ( .A(n4021), .B(n4022), .Z(n1409) );
  NANDN U4681 ( .A(B[366]), .B(n4023), .Z(n4022) );
  NANDN U4682 ( .A(A[366]), .B(n1411), .Z(n4023) );
  NANDN U4683 ( .A(n1411), .B(A[366]), .Z(n4021) );
  AND U4684 ( .A(n4024), .B(n4025), .Z(n1411) );
  NANDN U4685 ( .A(B[365]), .B(n4026), .Z(n4025) );
  NANDN U4686 ( .A(A[365]), .B(n1413), .Z(n4026) );
  NANDN U4687 ( .A(n1413), .B(A[365]), .Z(n4024) );
  AND U4688 ( .A(n4027), .B(n4028), .Z(n1413) );
  NANDN U4689 ( .A(B[364]), .B(n4029), .Z(n4028) );
  NANDN U4690 ( .A(A[364]), .B(n1415), .Z(n4029) );
  NANDN U4691 ( .A(n1415), .B(A[364]), .Z(n4027) );
  AND U4692 ( .A(n4030), .B(n4031), .Z(n1415) );
  NANDN U4693 ( .A(B[363]), .B(n4032), .Z(n4031) );
  NANDN U4694 ( .A(A[363]), .B(n1417), .Z(n4032) );
  NANDN U4695 ( .A(n1417), .B(A[363]), .Z(n4030) );
  AND U4696 ( .A(n4033), .B(n4034), .Z(n1417) );
  NANDN U4697 ( .A(B[362]), .B(n4035), .Z(n4034) );
  NANDN U4698 ( .A(A[362]), .B(n1419), .Z(n4035) );
  NANDN U4699 ( .A(n1419), .B(A[362]), .Z(n4033) );
  AND U4700 ( .A(n4036), .B(n4037), .Z(n1419) );
  NANDN U4701 ( .A(B[361]), .B(n4038), .Z(n4037) );
  NANDN U4702 ( .A(A[361]), .B(n1421), .Z(n4038) );
  NANDN U4703 ( .A(n1421), .B(A[361]), .Z(n4036) );
  AND U4704 ( .A(n4039), .B(n4040), .Z(n1421) );
  NANDN U4705 ( .A(B[360]), .B(n4041), .Z(n4040) );
  NANDN U4706 ( .A(A[360]), .B(n1423), .Z(n4041) );
  NANDN U4707 ( .A(n1423), .B(A[360]), .Z(n4039) );
  AND U4708 ( .A(n4042), .B(n4043), .Z(n1423) );
  NANDN U4709 ( .A(B[359]), .B(n4044), .Z(n4043) );
  NANDN U4710 ( .A(A[359]), .B(n1427), .Z(n4044) );
  NANDN U4711 ( .A(n1427), .B(A[359]), .Z(n4042) );
  AND U4712 ( .A(n4045), .B(n4046), .Z(n1427) );
  NANDN U4713 ( .A(B[358]), .B(n4047), .Z(n4046) );
  NANDN U4714 ( .A(A[358]), .B(n1429), .Z(n4047) );
  NANDN U4715 ( .A(n1429), .B(A[358]), .Z(n4045) );
  AND U4716 ( .A(n4048), .B(n4049), .Z(n1429) );
  NANDN U4717 ( .A(B[357]), .B(n4050), .Z(n4049) );
  NANDN U4718 ( .A(A[357]), .B(n1431), .Z(n4050) );
  NANDN U4719 ( .A(n1431), .B(A[357]), .Z(n4048) );
  AND U4720 ( .A(n4051), .B(n4052), .Z(n1431) );
  NANDN U4721 ( .A(B[356]), .B(n4053), .Z(n4052) );
  NANDN U4722 ( .A(A[356]), .B(n1433), .Z(n4053) );
  NANDN U4723 ( .A(n1433), .B(A[356]), .Z(n4051) );
  AND U4724 ( .A(n4054), .B(n4055), .Z(n1433) );
  NANDN U4725 ( .A(B[355]), .B(n4056), .Z(n4055) );
  NANDN U4726 ( .A(A[355]), .B(n1435), .Z(n4056) );
  NANDN U4727 ( .A(n1435), .B(A[355]), .Z(n4054) );
  AND U4728 ( .A(n4057), .B(n4058), .Z(n1435) );
  NANDN U4729 ( .A(B[354]), .B(n4059), .Z(n4058) );
  NANDN U4730 ( .A(A[354]), .B(n1437), .Z(n4059) );
  NANDN U4731 ( .A(n1437), .B(A[354]), .Z(n4057) );
  AND U4732 ( .A(n4060), .B(n4061), .Z(n1437) );
  NANDN U4733 ( .A(B[353]), .B(n4062), .Z(n4061) );
  NANDN U4734 ( .A(A[353]), .B(n1439), .Z(n4062) );
  NANDN U4735 ( .A(n1439), .B(A[353]), .Z(n4060) );
  AND U4736 ( .A(n4063), .B(n4064), .Z(n1439) );
  NANDN U4737 ( .A(B[352]), .B(n4065), .Z(n4064) );
  NANDN U4738 ( .A(A[352]), .B(n1441), .Z(n4065) );
  NANDN U4739 ( .A(n1441), .B(A[352]), .Z(n4063) );
  AND U4740 ( .A(n4066), .B(n4067), .Z(n1441) );
  NANDN U4741 ( .A(B[351]), .B(n4068), .Z(n4067) );
  NANDN U4742 ( .A(A[351]), .B(n1443), .Z(n4068) );
  NANDN U4743 ( .A(n1443), .B(A[351]), .Z(n4066) );
  AND U4744 ( .A(n4069), .B(n4070), .Z(n1443) );
  NANDN U4745 ( .A(B[350]), .B(n4071), .Z(n4070) );
  NANDN U4746 ( .A(A[350]), .B(n1445), .Z(n4071) );
  NANDN U4747 ( .A(n1445), .B(A[350]), .Z(n4069) );
  AND U4748 ( .A(n4072), .B(n4073), .Z(n1445) );
  NANDN U4749 ( .A(B[349]), .B(n4074), .Z(n4073) );
  NANDN U4750 ( .A(A[349]), .B(n1449), .Z(n4074) );
  NANDN U4751 ( .A(n1449), .B(A[349]), .Z(n4072) );
  AND U4752 ( .A(n4075), .B(n4076), .Z(n1449) );
  NANDN U4753 ( .A(B[348]), .B(n4077), .Z(n4076) );
  NANDN U4754 ( .A(A[348]), .B(n1451), .Z(n4077) );
  NANDN U4755 ( .A(n1451), .B(A[348]), .Z(n4075) );
  AND U4756 ( .A(n4078), .B(n4079), .Z(n1451) );
  NANDN U4757 ( .A(B[347]), .B(n4080), .Z(n4079) );
  NANDN U4758 ( .A(A[347]), .B(n1453), .Z(n4080) );
  NANDN U4759 ( .A(n1453), .B(A[347]), .Z(n4078) );
  AND U4760 ( .A(n4081), .B(n4082), .Z(n1453) );
  NANDN U4761 ( .A(B[346]), .B(n4083), .Z(n4082) );
  NANDN U4762 ( .A(A[346]), .B(n1455), .Z(n4083) );
  NANDN U4763 ( .A(n1455), .B(A[346]), .Z(n4081) );
  AND U4764 ( .A(n4084), .B(n4085), .Z(n1455) );
  NANDN U4765 ( .A(B[345]), .B(n4086), .Z(n4085) );
  NANDN U4766 ( .A(A[345]), .B(n1457), .Z(n4086) );
  NANDN U4767 ( .A(n1457), .B(A[345]), .Z(n4084) );
  AND U4768 ( .A(n4087), .B(n4088), .Z(n1457) );
  NANDN U4769 ( .A(B[344]), .B(n4089), .Z(n4088) );
  NANDN U4770 ( .A(A[344]), .B(n1459), .Z(n4089) );
  NANDN U4771 ( .A(n1459), .B(A[344]), .Z(n4087) );
  AND U4772 ( .A(n4090), .B(n4091), .Z(n1459) );
  NANDN U4773 ( .A(B[343]), .B(n4092), .Z(n4091) );
  NANDN U4774 ( .A(A[343]), .B(n1461), .Z(n4092) );
  NANDN U4775 ( .A(n1461), .B(A[343]), .Z(n4090) );
  AND U4776 ( .A(n4093), .B(n4094), .Z(n1461) );
  NANDN U4777 ( .A(B[342]), .B(n4095), .Z(n4094) );
  NANDN U4778 ( .A(A[342]), .B(n1463), .Z(n4095) );
  NANDN U4779 ( .A(n1463), .B(A[342]), .Z(n4093) );
  AND U4780 ( .A(n4096), .B(n4097), .Z(n1463) );
  NANDN U4781 ( .A(B[341]), .B(n4098), .Z(n4097) );
  NANDN U4782 ( .A(A[341]), .B(n1465), .Z(n4098) );
  NANDN U4783 ( .A(n1465), .B(A[341]), .Z(n4096) );
  AND U4784 ( .A(n4099), .B(n4100), .Z(n1465) );
  NANDN U4785 ( .A(B[340]), .B(n4101), .Z(n4100) );
  NANDN U4786 ( .A(A[340]), .B(n1467), .Z(n4101) );
  NANDN U4787 ( .A(n1467), .B(A[340]), .Z(n4099) );
  AND U4788 ( .A(n4102), .B(n4103), .Z(n1467) );
  NANDN U4789 ( .A(B[339]), .B(n4104), .Z(n4103) );
  NANDN U4790 ( .A(A[339]), .B(n1471), .Z(n4104) );
  NANDN U4791 ( .A(n1471), .B(A[339]), .Z(n4102) );
  AND U4792 ( .A(n4105), .B(n4106), .Z(n1471) );
  NANDN U4793 ( .A(B[338]), .B(n4107), .Z(n4106) );
  NANDN U4794 ( .A(A[338]), .B(n1473), .Z(n4107) );
  NANDN U4795 ( .A(n1473), .B(A[338]), .Z(n4105) );
  AND U4796 ( .A(n4108), .B(n4109), .Z(n1473) );
  NANDN U4797 ( .A(B[337]), .B(n4110), .Z(n4109) );
  NANDN U4798 ( .A(A[337]), .B(n1475), .Z(n4110) );
  NANDN U4799 ( .A(n1475), .B(A[337]), .Z(n4108) );
  AND U4800 ( .A(n4111), .B(n4112), .Z(n1475) );
  NANDN U4801 ( .A(B[336]), .B(n4113), .Z(n4112) );
  NANDN U4802 ( .A(A[336]), .B(n1477), .Z(n4113) );
  NANDN U4803 ( .A(n1477), .B(A[336]), .Z(n4111) );
  AND U4804 ( .A(n4114), .B(n4115), .Z(n1477) );
  NANDN U4805 ( .A(B[335]), .B(n4116), .Z(n4115) );
  NANDN U4806 ( .A(A[335]), .B(n1479), .Z(n4116) );
  NANDN U4807 ( .A(n1479), .B(A[335]), .Z(n4114) );
  AND U4808 ( .A(n4117), .B(n4118), .Z(n1479) );
  NANDN U4809 ( .A(B[334]), .B(n4119), .Z(n4118) );
  NANDN U4810 ( .A(A[334]), .B(n1481), .Z(n4119) );
  NANDN U4811 ( .A(n1481), .B(A[334]), .Z(n4117) );
  AND U4812 ( .A(n4120), .B(n4121), .Z(n1481) );
  NANDN U4813 ( .A(B[333]), .B(n4122), .Z(n4121) );
  NANDN U4814 ( .A(A[333]), .B(n1483), .Z(n4122) );
  NANDN U4815 ( .A(n1483), .B(A[333]), .Z(n4120) );
  AND U4816 ( .A(n4123), .B(n4124), .Z(n1483) );
  NANDN U4817 ( .A(B[332]), .B(n4125), .Z(n4124) );
  NANDN U4818 ( .A(A[332]), .B(n1485), .Z(n4125) );
  NANDN U4819 ( .A(n1485), .B(A[332]), .Z(n4123) );
  AND U4820 ( .A(n4126), .B(n4127), .Z(n1485) );
  NANDN U4821 ( .A(B[331]), .B(n4128), .Z(n4127) );
  NANDN U4822 ( .A(A[331]), .B(n1487), .Z(n4128) );
  NANDN U4823 ( .A(n1487), .B(A[331]), .Z(n4126) );
  AND U4824 ( .A(n4129), .B(n4130), .Z(n1487) );
  NANDN U4825 ( .A(B[330]), .B(n4131), .Z(n4130) );
  NANDN U4826 ( .A(A[330]), .B(n1489), .Z(n4131) );
  NANDN U4827 ( .A(n1489), .B(A[330]), .Z(n4129) );
  AND U4828 ( .A(n4132), .B(n4133), .Z(n1489) );
  NANDN U4829 ( .A(B[329]), .B(n4134), .Z(n4133) );
  NANDN U4830 ( .A(A[329]), .B(n1493), .Z(n4134) );
  NANDN U4831 ( .A(n1493), .B(A[329]), .Z(n4132) );
  AND U4832 ( .A(n4135), .B(n4136), .Z(n1493) );
  NANDN U4833 ( .A(B[328]), .B(n4137), .Z(n4136) );
  NANDN U4834 ( .A(A[328]), .B(n1495), .Z(n4137) );
  NANDN U4835 ( .A(n1495), .B(A[328]), .Z(n4135) );
  AND U4836 ( .A(n4138), .B(n4139), .Z(n1495) );
  NANDN U4837 ( .A(B[327]), .B(n4140), .Z(n4139) );
  NANDN U4838 ( .A(A[327]), .B(n1497), .Z(n4140) );
  NANDN U4839 ( .A(n1497), .B(A[327]), .Z(n4138) );
  AND U4840 ( .A(n4141), .B(n4142), .Z(n1497) );
  NANDN U4841 ( .A(B[326]), .B(n4143), .Z(n4142) );
  NANDN U4842 ( .A(A[326]), .B(n1499), .Z(n4143) );
  NANDN U4843 ( .A(n1499), .B(A[326]), .Z(n4141) );
  AND U4844 ( .A(n4144), .B(n4145), .Z(n1499) );
  NANDN U4845 ( .A(B[325]), .B(n4146), .Z(n4145) );
  NANDN U4846 ( .A(A[325]), .B(n1501), .Z(n4146) );
  NANDN U4847 ( .A(n1501), .B(A[325]), .Z(n4144) );
  AND U4848 ( .A(n4147), .B(n4148), .Z(n1501) );
  NANDN U4849 ( .A(B[324]), .B(n4149), .Z(n4148) );
  NANDN U4850 ( .A(A[324]), .B(n1503), .Z(n4149) );
  NANDN U4851 ( .A(n1503), .B(A[324]), .Z(n4147) );
  AND U4852 ( .A(n4150), .B(n4151), .Z(n1503) );
  NANDN U4853 ( .A(B[323]), .B(n4152), .Z(n4151) );
  NANDN U4854 ( .A(A[323]), .B(n1505), .Z(n4152) );
  NANDN U4855 ( .A(n1505), .B(A[323]), .Z(n4150) );
  AND U4856 ( .A(n4153), .B(n4154), .Z(n1505) );
  NANDN U4857 ( .A(B[322]), .B(n4155), .Z(n4154) );
  NANDN U4858 ( .A(A[322]), .B(n1507), .Z(n4155) );
  NANDN U4859 ( .A(n1507), .B(A[322]), .Z(n4153) );
  AND U4860 ( .A(n4156), .B(n4157), .Z(n1507) );
  NANDN U4861 ( .A(B[321]), .B(n4158), .Z(n4157) );
  NANDN U4862 ( .A(A[321]), .B(n1509), .Z(n4158) );
  NANDN U4863 ( .A(n1509), .B(A[321]), .Z(n4156) );
  AND U4864 ( .A(n4159), .B(n4160), .Z(n1509) );
  NANDN U4865 ( .A(B[320]), .B(n4161), .Z(n4160) );
  NANDN U4866 ( .A(A[320]), .B(n1511), .Z(n4161) );
  NANDN U4867 ( .A(n1511), .B(A[320]), .Z(n4159) );
  AND U4868 ( .A(n4162), .B(n4163), .Z(n1511) );
  NANDN U4869 ( .A(B[319]), .B(n4164), .Z(n4163) );
  NANDN U4870 ( .A(A[319]), .B(n1515), .Z(n4164) );
  NANDN U4871 ( .A(n1515), .B(A[319]), .Z(n4162) );
  AND U4872 ( .A(n4165), .B(n4166), .Z(n1515) );
  NANDN U4873 ( .A(B[318]), .B(n4167), .Z(n4166) );
  NANDN U4874 ( .A(A[318]), .B(n1517), .Z(n4167) );
  NANDN U4875 ( .A(n1517), .B(A[318]), .Z(n4165) );
  AND U4876 ( .A(n4168), .B(n4169), .Z(n1517) );
  NANDN U4877 ( .A(B[317]), .B(n4170), .Z(n4169) );
  NANDN U4878 ( .A(A[317]), .B(n1519), .Z(n4170) );
  NANDN U4879 ( .A(n1519), .B(A[317]), .Z(n4168) );
  AND U4880 ( .A(n4171), .B(n4172), .Z(n1519) );
  NANDN U4881 ( .A(B[316]), .B(n4173), .Z(n4172) );
  NANDN U4882 ( .A(A[316]), .B(n1521), .Z(n4173) );
  NANDN U4883 ( .A(n1521), .B(A[316]), .Z(n4171) );
  AND U4884 ( .A(n4174), .B(n4175), .Z(n1521) );
  NANDN U4885 ( .A(B[315]), .B(n4176), .Z(n4175) );
  NANDN U4886 ( .A(A[315]), .B(n1523), .Z(n4176) );
  NANDN U4887 ( .A(n1523), .B(A[315]), .Z(n4174) );
  AND U4888 ( .A(n4177), .B(n4178), .Z(n1523) );
  NANDN U4889 ( .A(B[314]), .B(n4179), .Z(n4178) );
  NANDN U4890 ( .A(A[314]), .B(n1525), .Z(n4179) );
  NANDN U4891 ( .A(n1525), .B(A[314]), .Z(n4177) );
  AND U4892 ( .A(n4180), .B(n4181), .Z(n1525) );
  NANDN U4893 ( .A(B[313]), .B(n4182), .Z(n4181) );
  NANDN U4894 ( .A(A[313]), .B(n1527), .Z(n4182) );
  NANDN U4895 ( .A(n1527), .B(A[313]), .Z(n4180) );
  AND U4896 ( .A(n4183), .B(n4184), .Z(n1527) );
  NANDN U4897 ( .A(B[312]), .B(n4185), .Z(n4184) );
  NANDN U4898 ( .A(A[312]), .B(n1529), .Z(n4185) );
  NANDN U4899 ( .A(n1529), .B(A[312]), .Z(n4183) );
  AND U4900 ( .A(n4186), .B(n4187), .Z(n1529) );
  NANDN U4901 ( .A(B[311]), .B(n4188), .Z(n4187) );
  NANDN U4902 ( .A(A[311]), .B(n1531), .Z(n4188) );
  NANDN U4903 ( .A(n1531), .B(A[311]), .Z(n4186) );
  AND U4904 ( .A(n4189), .B(n4190), .Z(n1531) );
  NANDN U4905 ( .A(B[310]), .B(n4191), .Z(n4190) );
  NANDN U4906 ( .A(A[310]), .B(n1533), .Z(n4191) );
  NANDN U4907 ( .A(n1533), .B(A[310]), .Z(n4189) );
  AND U4908 ( .A(n4192), .B(n4193), .Z(n1533) );
  NANDN U4909 ( .A(B[309]), .B(n4194), .Z(n4193) );
  NANDN U4910 ( .A(A[309]), .B(n1537), .Z(n4194) );
  NANDN U4911 ( .A(n1537), .B(A[309]), .Z(n4192) );
  AND U4912 ( .A(n4195), .B(n4196), .Z(n1537) );
  NANDN U4913 ( .A(B[308]), .B(n4197), .Z(n4196) );
  NANDN U4914 ( .A(A[308]), .B(n1539), .Z(n4197) );
  NANDN U4915 ( .A(n1539), .B(A[308]), .Z(n4195) );
  AND U4916 ( .A(n4198), .B(n4199), .Z(n1539) );
  NANDN U4917 ( .A(B[307]), .B(n4200), .Z(n4199) );
  NANDN U4918 ( .A(A[307]), .B(n1541), .Z(n4200) );
  NANDN U4919 ( .A(n1541), .B(A[307]), .Z(n4198) );
  AND U4920 ( .A(n4201), .B(n4202), .Z(n1541) );
  NANDN U4921 ( .A(B[306]), .B(n4203), .Z(n4202) );
  NANDN U4922 ( .A(A[306]), .B(n1543), .Z(n4203) );
  NANDN U4923 ( .A(n1543), .B(A[306]), .Z(n4201) );
  AND U4924 ( .A(n4204), .B(n4205), .Z(n1543) );
  NANDN U4925 ( .A(B[305]), .B(n4206), .Z(n4205) );
  NANDN U4926 ( .A(A[305]), .B(n1545), .Z(n4206) );
  NANDN U4927 ( .A(n1545), .B(A[305]), .Z(n4204) );
  AND U4928 ( .A(n4207), .B(n4208), .Z(n1545) );
  NANDN U4929 ( .A(B[304]), .B(n4209), .Z(n4208) );
  NANDN U4930 ( .A(A[304]), .B(n1547), .Z(n4209) );
  NANDN U4931 ( .A(n1547), .B(A[304]), .Z(n4207) );
  AND U4932 ( .A(n4210), .B(n4211), .Z(n1547) );
  NANDN U4933 ( .A(B[303]), .B(n4212), .Z(n4211) );
  NANDN U4934 ( .A(A[303]), .B(n1549), .Z(n4212) );
  NANDN U4935 ( .A(n1549), .B(A[303]), .Z(n4210) );
  AND U4936 ( .A(n4213), .B(n4214), .Z(n1549) );
  NANDN U4937 ( .A(B[302]), .B(n4215), .Z(n4214) );
  NANDN U4938 ( .A(A[302]), .B(n1551), .Z(n4215) );
  NANDN U4939 ( .A(n1551), .B(A[302]), .Z(n4213) );
  AND U4940 ( .A(n4216), .B(n4217), .Z(n1551) );
  NANDN U4941 ( .A(B[301]), .B(n4218), .Z(n4217) );
  NANDN U4942 ( .A(A[301]), .B(n1553), .Z(n4218) );
  NANDN U4943 ( .A(n1553), .B(A[301]), .Z(n4216) );
  AND U4944 ( .A(n4219), .B(n4220), .Z(n1553) );
  NANDN U4945 ( .A(B[300]), .B(n4221), .Z(n4220) );
  NANDN U4946 ( .A(A[300]), .B(n1555), .Z(n4221) );
  NANDN U4947 ( .A(n1555), .B(A[300]), .Z(n4219) );
  AND U4948 ( .A(n4222), .B(n4223), .Z(n1555) );
  NANDN U4949 ( .A(B[299]), .B(n4224), .Z(n4223) );
  NANDN U4950 ( .A(A[299]), .B(n1561), .Z(n4224) );
  NANDN U4951 ( .A(n1561), .B(A[299]), .Z(n4222) );
  AND U4952 ( .A(n4225), .B(n4226), .Z(n1561) );
  NANDN U4953 ( .A(B[298]), .B(n4227), .Z(n4226) );
  NANDN U4954 ( .A(A[298]), .B(n1563), .Z(n4227) );
  NANDN U4955 ( .A(n1563), .B(A[298]), .Z(n4225) );
  AND U4956 ( .A(n4228), .B(n4229), .Z(n1563) );
  NANDN U4957 ( .A(B[297]), .B(n4230), .Z(n4229) );
  NANDN U4958 ( .A(A[297]), .B(n1565), .Z(n4230) );
  NANDN U4959 ( .A(n1565), .B(A[297]), .Z(n4228) );
  AND U4960 ( .A(n4231), .B(n4232), .Z(n1565) );
  NANDN U4961 ( .A(B[296]), .B(n4233), .Z(n4232) );
  NANDN U4962 ( .A(A[296]), .B(n1567), .Z(n4233) );
  NANDN U4963 ( .A(n1567), .B(A[296]), .Z(n4231) );
  AND U4964 ( .A(n4234), .B(n4235), .Z(n1567) );
  NANDN U4965 ( .A(B[295]), .B(n4236), .Z(n4235) );
  NANDN U4966 ( .A(A[295]), .B(n1569), .Z(n4236) );
  NANDN U4967 ( .A(n1569), .B(A[295]), .Z(n4234) );
  AND U4968 ( .A(n4237), .B(n4238), .Z(n1569) );
  NANDN U4969 ( .A(B[294]), .B(n4239), .Z(n4238) );
  NANDN U4970 ( .A(A[294]), .B(n1571), .Z(n4239) );
  NANDN U4971 ( .A(n1571), .B(A[294]), .Z(n4237) );
  AND U4972 ( .A(n4240), .B(n4241), .Z(n1571) );
  NANDN U4973 ( .A(B[293]), .B(n4242), .Z(n4241) );
  NANDN U4974 ( .A(A[293]), .B(n1573), .Z(n4242) );
  NANDN U4975 ( .A(n1573), .B(A[293]), .Z(n4240) );
  AND U4976 ( .A(n4243), .B(n4244), .Z(n1573) );
  NANDN U4977 ( .A(B[292]), .B(n4245), .Z(n4244) );
  NANDN U4978 ( .A(A[292]), .B(n1575), .Z(n4245) );
  NANDN U4979 ( .A(n1575), .B(A[292]), .Z(n4243) );
  AND U4980 ( .A(n4246), .B(n4247), .Z(n1575) );
  NANDN U4981 ( .A(B[291]), .B(n4248), .Z(n4247) );
  NANDN U4982 ( .A(A[291]), .B(n1577), .Z(n4248) );
  NANDN U4983 ( .A(n1577), .B(A[291]), .Z(n4246) );
  AND U4984 ( .A(n4249), .B(n4250), .Z(n1577) );
  NANDN U4985 ( .A(B[290]), .B(n4251), .Z(n4250) );
  NANDN U4986 ( .A(A[290]), .B(n1579), .Z(n4251) );
  NANDN U4987 ( .A(n1579), .B(A[290]), .Z(n4249) );
  AND U4988 ( .A(n4252), .B(n4253), .Z(n1579) );
  NANDN U4989 ( .A(B[289]), .B(n4254), .Z(n4253) );
  NANDN U4990 ( .A(A[289]), .B(n1583), .Z(n4254) );
  NANDN U4991 ( .A(n1583), .B(A[289]), .Z(n4252) );
  AND U4992 ( .A(n4255), .B(n4256), .Z(n1583) );
  NANDN U4993 ( .A(B[288]), .B(n4257), .Z(n4256) );
  NANDN U4994 ( .A(A[288]), .B(n1585), .Z(n4257) );
  NANDN U4995 ( .A(n1585), .B(A[288]), .Z(n4255) );
  AND U4996 ( .A(n4258), .B(n4259), .Z(n1585) );
  NANDN U4997 ( .A(B[287]), .B(n4260), .Z(n4259) );
  NANDN U4998 ( .A(A[287]), .B(n1587), .Z(n4260) );
  NANDN U4999 ( .A(n1587), .B(A[287]), .Z(n4258) );
  AND U5000 ( .A(n4261), .B(n4262), .Z(n1587) );
  NANDN U5001 ( .A(B[286]), .B(n4263), .Z(n4262) );
  NANDN U5002 ( .A(A[286]), .B(n1589), .Z(n4263) );
  NANDN U5003 ( .A(n1589), .B(A[286]), .Z(n4261) );
  AND U5004 ( .A(n4264), .B(n4265), .Z(n1589) );
  NANDN U5005 ( .A(B[285]), .B(n4266), .Z(n4265) );
  NANDN U5006 ( .A(A[285]), .B(n1591), .Z(n4266) );
  NANDN U5007 ( .A(n1591), .B(A[285]), .Z(n4264) );
  AND U5008 ( .A(n4267), .B(n4268), .Z(n1591) );
  NANDN U5009 ( .A(B[284]), .B(n4269), .Z(n4268) );
  NANDN U5010 ( .A(A[284]), .B(n1593), .Z(n4269) );
  NANDN U5011 ( .A(n1593), .B(A[284]), .Z(n4267) );
  AND U5012 ( .A(n4270), .B(n4271), .Z(n1593) );
  NANDN U5013 ( .A(B[283]), .B(n4272), .Z(n4271) );
  NANDN U5014 ( .A(A[283]), .B(n1595), .Z(n4272) );
  NANDN U5015 ( .A(n1595), .B(A[283]), .Z(n4270) );
  AND U5016 ( .A(n4273), .B(n4274), .Z(n1595) );
  NANDN U5017 ( .A(B[282]), .B(n4275), .Z(n4274) );
  NANDN U5018 ( .A(A[282]), .B(n1597), .Z(n4275) );
  NANDN U5019 ( .A(n1597), .B(A[282]), .Z(n4273) );
  AND U5020 ( .A(n4276), .B(n4277), .Z(n1597) );
  NANDN U5021 ( .A(B[281]), .B(n4278), .Z(n4277) );
  NANDN U5022 ( .A(A[281]), .B(n1599), .Z(n4278) );
  NANDN U5023 ( .A(n1599), .B(A[281]), .Z(n4276) );
  AND U5024 ( .A(n4279), .B(n4280), .Z(n1599) );
  NANDN U5025 ( .A(B[280]), .B(n4281), .Z(n4280) );
  NANDN U5026 ( .A(A[280]), .B(n1601), .Z(n4281) );
  NANDN U5027 ( .A(n1601), .B(A[280]), .Z(n4279) );
  AND U5028 ( .A(n4282), .B(n4283), .Z(n1601) );
  NANDN U5029 ( .A(B[279]), .B(n4284), .Z(n4283) );
  NANDN U5030 ( .A(A[279]), .B(n1605), .Z(n4284) );
  NANDN U5031 ( .A(n1605), .B(A[279]), .Z(n4282) );
  AND U5032 ( .A(n4285), .B(n4286), .Z(n1605) );
  NANDN U5033 ( .A(B[278]), .B(n4287), .Z(n4286) );
  NANDN U5034 ( .A(A[278]), .B(n1607), .Z(n4287) );
  NANDN U5035 ( .A(n1607), .B(A[278]), .Z(n4285) );
  AND U5036 ( .A(n4288), .B(n4289), .Z(n1607) );
  NANDN U5037 ( .A(B[277]), .B(n4290), .Z(n4289) );
  NANDN U5038 ( .A(A[277]), .B(n1609), .Z(n4290) );
  NANDN U5039 ( .A(n1609), .B(A[277]), .Z(n4288) );
  AND U5040 ( .A(n4291), .B(n4292), .Z(n1609) );
  NANDN U5041 ( .A(B[276]), .B(n4293), .Z(n4292) );
  NANDN U5042 ( .A(A[276]), .B(n1611), .Z(n4293) );
  NANDN U5043 ( .A(n1611), .B(A[276]), .Z(n4291) );
  AND U5044 ( .A(n4294), .B(n4295), .Z(n1611) );
  NANDN U5045 ( .A(B[275]), .B(n4296), .Z(n4295) );
  NANDN U5046 ( .A(A[275]), .B(n1613), .Z(n4296) );
  NANDN U5047 ( .A(n1613), .B(A[275]), .Z(n4294) );
  AND U5048 ( .A(n4297), .B(n4298), .Z(n1613) );
  NANDN U5049 ( .A(B[274]), .B(n4299), .Z(n4298) );
  NANDN U5050 ( .A(A[274]), .B(n1615), .Z(n4299) );
  NANDN U5051 ( .A(n1615), .B(A[274]), .Z(n4297) );
  AND U5052 ( .A(n4300), .B(n4301), .Z(n1615) );
  NANDN U5053 ( .A(B[273]), .B(n4302), .Z(n4301) );
  NANDN U5054 ( .A(A[273]), .B(n1617), .Z(n4302) );
  NANDN U5055 ( .A(n1617), .B(A[273]), .Z(n4300) );
  AND U5056 ( .A(n4303), .B(n4304), .Z(n1617) );
  NANDN U5057 ( .A(B[272]), .B(n4305), .Z(n4304) );
  NANDN U5058 ( .A(A[272]), .B(n1619), .Z(n4305) );
  NANDN U5059 ( .A(n1619), .B(A[272]), .Z(n4303) );
  AND U5060 ( .A(n4306), .B(n4307), .Z(n1619) );
  NANDN U5061 ( .A(B[271]), .B(n4308), .Z(n4307) );
  NANDN U5062 ( .A(A[271]), .B(n1621), .Z(n4308) );
  NANDN U5063 ( .A(n1621), .B(A[271]), .Z(n4306) );
  AND U5064 ( .A(n4309), .B(n4310), .Z(n1621) );
  NANDN U5065 ( .A(B[270]), .B(n4311), .Z(n4310) );
  NANDN U5066 ( .A(A[270]), .B(n1623), .Z(n4311) );
  NANDN U5067 ( .A(n1623), .B(A[270]), .Z(n4309) );
  AND U5068 ( .A(n4312), .B(n4313), .Z(n1623) );
  NANDN U5069 ( .A(B[269]), .B(n4314), .Z(n4313) );
  NANDN U5070 ( .A(A[269]), .B(n1627), .Z(n4314) );
  NANDN U5071 ( .A(n1627), .B(A[269]), .Z(n4312) );
  AND U5072 ( .A(n4315), .B(n4316), .Z(n1627) );
  NANDN U5073 ( .A(B[268]), .B(n4317), .Z(n4316) );
  NANDN U5074 ( .A(A[268]), .B(n1629), .Z(n4317) );
  NANDN U5075 ( .A(n1629), .B(A[268]), .Z(n4315) );
  AND U5076 ( .A(n4318), .B(n4319), .Z(n1629) );
  NANDN U5077 ( .A(B[267]), .B(n4320), .Z(n4319) );
  NANDN U5078 ( .A(A[267]), .B(n1631), .Z(n4320) );
  NANDN U5079 ( .A(n1631), .B(A[267]), .Z(n4318) );
  AND U5080 ( .A(n4321), .B(n4322), .Z(n1631) );
  NANDN U5081 ( .A(B[266]), .B(n4323), .Z(n4322) );
  NANDN U5082 ( .A(A[266]), .B(n1633), .Z(n4323) );
  NANDN U5083 ( .A(n1633), .B(A[266]), .Z(n4321) );
  AND U5084 ( .A(n4324), .B(n4325), .Z(n1633) );
  NANDN U5085 ( .A(B[265]), .B(n4326), .Z(n4325) );
  NANDN U5086 ( .A(A[265]), .B(n1635), .Z(n4326) );
  NANDN U5087 ( .A(n1635), .B(A[265]), .Z(n4324) );
  AND U5088 ( .A(n4327), .B(n4328), .Z(n1635) );
  NANDN U5089 ( .A(B[264]), .B(n4329), .Z(n4328) );
  NANDN U5090 ( .A(A[264]), .B(n1637), .Z(n4329) );
  NANDN U5091 ( .A(n1637), .B(A[264]), .Z(n4327) );
  AND U5092 ( .A(n4330), .B(n4331), .Z(n1637) );
  NANDN U5093 ( .A(B[263]), .B(n4332), .Z(n4331) );
  NANDN U5094 ( .A(A[263]), .B(n1639), .Z(n4332) );
  NANDN U5095 ( .A(n1639), .B(A[263]), .Z(n4330) );
  AND U5096 ( .A(n4333), .B(n4334), .Z(n1639) );
  NANDN U5097 ( .A(B[262]), .B(n4335), .Z(n4334) );
  NANDN U5098 ( .A(A[262]), .B(n1641), .Z(n4335) );
  NANDN U5099 ( .A(n1641), .B(A[262]), .Z(n4333) );
  AND U5100 ( .A(n4336), .B(n4337), .Z(n1641) );
  NANDN U5101 ( .A(B[261]), .B(n4338), .Z(n4337) );
  NANDN U5102 ( .A(A[261]), .B(n1643), .Z(n4338) );
  NANDN U5103 ( .A(n1643), .B(A[261]), .Z(n4336) );
  AND U5104 ( .A(n4339), .B(n4340), .Z(n1643) );
  NANDN U5105 ( .A(B[260]), .B(n4341), .Z(n4340) );
  NANDN U5106 ( .A(A[260]), .B(n1645), .Z(n4341) );
  NANDN U5107 ( .A(n1645), .B(A[260]), .Z(n4339) );
  AND U5108 ( .A(n4342), .B(n4343), .Z(n1645) );
  NANDN U5109 ( .A(B[259]), .B(n4344), .Z(n4343) );
  NANDN U5110 ( .A(A[259]), .B(n1649), .Z(n4344) );
  NANDN U5111 ( .A(n1649), .B(A[259]), .Z(n4342) );
  AND U5112 ( .A(n4345), .B(n4346), .Z(n1649) );
  NANDN U5113 ( .A(B[258]), .B(n4347), .Z(n4346) );
  NANDN U5114 ( .A(A[258]), .B(n1651), .Z(n4347) );
  NANDN U5115 ( .A(n1651), .B(A[258]), .Z(n4345) );
  AND U5116 ( .A(n4348), .B(n4349), .Z(n1651) );
  NANDN U5117 ( .A(B[257]), .B(n4350), .Z(n4349) );
  NANDN U5118 ( .A(A[257]), .B(n1653), .Z(n4350) );
  NANDN U5119 ( .A(n1653), .B(A[257]), .Z(n4348) );
  AND U5120 ( .A(n4351), .B(n4352), .Z(n1653) );
  NANDN U5121 ( .A(B[256]), .B(n4353), .Z(n4352) );
  NANDN U5122 ( .A(A[256]), .B(n1655), .Z(n4353) );
  NANDN U5123 ( .A(n1655), .B(A[256]), .Z(n4351) );
  AND U5124 ( .A(n4354), .B(n4355), .Z(n1655) );
  NANDN U5125 ( .A(B[255]), .B(n4356), .Z(n4355) );
  NANDN U5126 ( .A(A[255]), .B(n1657), .Z(n4356) );
  NANDN U5127 ( .A(n1657), .B(A[255]), .Z(n4354) );
  AND U5128 ( .A(n4357), .B(n4358), .Z(n1657) );
  NANDN U5129 ( .A(B[254]), .B(n4359), .Z(n4358) );
  NANDN U5130 ( .A(A[254]), .B(n1659), .Z(n4359) );
  NANDN U5131 ( .A(n1659), .B(A[254]), .Z(n4357) );
  AND U5132 ( .A(n4360), .B(n4361), .Z(n1659) );
  NANDN U5133 ( .A(B[253]), .B(n4362), .Z(n4361) );
  NANDN U5134 ( .A(A[253]), .B(n1661), .Z(n4362) );
  NANDN U5135 ( .A(n1661), .B(A[253]), .Z(n4360) );
  AND U5136 ( .A(n4363), .B(n4364), .Z(n1661) );
  NANDN U5137 ( .A(B[252]), .B(n4365), .Z(n4364) );
  NANDN U5138 ( .A(A[252]), .B(n1663), .Z(n4365) );
  NANDN U5139 ( .A(n1663), .B(A[252]), .Z(n4363) );
  AND U5140 ( .A(n4366), .B(n4367), .Z(n1663) );
  NANDN U5141 ( .A(B[251]), .B(n4368), .Z(n4367) );
  NANDN U5142 ( .A(A[251]), .B(n1665), .Z(n4368) );
  NANDN U5143 ( .A(n1665), .B(A[251]), .Z(n4366) );
  AND U5144 ( .A(n4369), .B(n4370), .Z(n1665) );
  NANDN U5145 ( .A(B[250]), .B(n4371), .Z(n4370) );
  NANDN U5146 ( .A(A[250]), .B(n1667), .Z(n4371) );
  NANDN U5147 ( .A(n1667), .B(A[250]), .Z(n4369) );
  AND U5148 ( .A(n4372), .B(n4373), .Z(n1667) );
  NANDN U5149 ( .A(B[249]), .B(n4374), .Z(n4373) );
  NANDN U5150 ( .A(A[249]), .B(n1671), .Z(n4374) );
  NANDN U5151 ( .A(n1671), .B(A[249]), .Z(n4372) );
  AND U5152 ( .A(n4375), .B(n4376), .Z(n1671) );
  NANDN U5153 ( .A(B[248]), .B(n4377), .Z(n4376) );
  NANDN U5154 ( .A(A[248]), .B(n1673), .Z(n4377) );
  NANDN U5155 ( .A(n1673), .B(A[248]), .Z(n4375) );
  AND U5156 ( .A(n4378), .B(n4379), .Z(n1673) );
  NANDN U5157 ( .A(B[247]), .B(n4380), .Z(n4379) );
  NANDN U5158 ( .A(A[247]), .B(n1675), .Z(n4380) );
  NANDN U5159 ( .A(n1675), .B(A[247]), .Z(n4378) );
  AND U5160 ( .A(n4381), .B(n4382), .Z(n1675) );
  NANDN U5161 ( .A(B[246]), .B(n4383), .Z(n4382) );
  NANDN U5162 ( .A(A[246]), .B(n1677), .Z(n4383) );
  NANDN U5163 ( .A(n1677), .B(A[246]), .Z(n4381) );
  AND U5164 ( .A(n4384), .B(n4385), .Z(n1677) );
  NANDN U5165 ( .A(B[245]), .B(n4386), .Z(n4385) );
  NANDN U5166 ( .A(A[245]), .B(n1679), .Z(n4386) );
  NANDN U5167 ( .A(n1679), .B(A[245]), .Z(n4384) );
  AND U5168 ( .A(n4387), .B(n4388), .Z(n1679) );
  NANDN U5169 ( .A(B[244]), .B(n4389), .Z(n4388) );
  NANDN U5170 ( .A(A[244]), .B(n1681), .Z(n4389) );
  NANDN U5171 ( .A(n1681), .B(A[244]), .Z(n4387) );
  AND U5172 ( .A(n4390), .B(n4391), .Z(n1681) );
  NANDN U5173 ( .A(B[243]), .B(n4392), .Z(n4391) );
  NANDN U5174 ( .A(A[243]), .B(n1683), .Z(n4392) );
  NANDN U5175 ( .A(n1683), .B(A[243]), .Z(n4390) );
  AND U5176 ( .A(n4393), .B(n4394), .Z(n1683) );
  NANDN U5177 ( .A(B[242]), .B(n4395), .Z(n4394) );
  NANDN U5178 ( .A(A[242]), .B(n1685), .Z(n4395) );
  NANDN U5179 ( .A(n1685), .B(A[242]), .Z(n4393) );
  AND U5180 ( .A(n4396), .B(n4397), .Z(n1685) );
  NANDN U5181 ( .A(B[241]), .B(n4398), .Z(n4397) );
  NANDN U5182 ( .A(A[241]), .B(n1687), .Z(n4398) );
  NANDN U5183 ( .A(n1687), .B(A[241]), .Z(n4396) );
  AND U5184 ( .A(n4399), .B(n4400), .Z(n1687) );
  NANDN U5185 ( .A(B[240]), .B(n4401), .Z(n4400) );
  NANDN U5186 ( .A(A[240]), .B(n1689), .Z(n4401) );
  NANDN U5187 ( .A(n1689), .B(A[240]), .Z(n4399) );
  AND U5188 ( .A(n4402), .B(n4403), .Z(n1689) );
  NANDN U5189 ( .A(B[239]), .B(n4404), .Z(n4403) );
  NANDN U5190 ( .A(A[239]), .B(n1693), .Z(n4404) );
  NANDN U5191 ( .A(n1693), .B(A[239]), .Z(n4402) );
  AND U5192 ( .A(n4405), .B(n4406), .Z(n1693) );
  NANDN U5193 ( .A(B[238]), .B(n4407), .Z(n4406) );
  NANDN U5194 ( .A(A[238]), .B(n1695), .Z(n4407) );
  NANDN U5195 ( .A(n1695), .B(A[238]), .Z(n4405) );
  AND U5196 ( .A(n4408), .B(n4409), .Z(n1695) );
  NANDN U5197 ( .A(B[237]), .B(n4410), .Z(n4409) );
  NANDN U5198 ( .A(A[237]), .B(n1697), .Z(n4410) );
  NANDN U5199 ( .A(n1697), .B(A[237]), .Z(n4408) );
  AND U5200 ( .A(n4411), .B(n4412), .Z(n1697) );
  NANDN U5201 ( .A(B[236]), .B(n4413), .Z(n4412) );
  NANDN U5202 ( .A(A[236]), .B(n1699), .Z(n4413) );
  NANDN U5203 ( .A(n1699), .B(A[236]), .Z(n4411) );
  AND U5204 ( .A(n4414), .B(n4415), .Z(n1699) );
  NANDN U5205 ( .A(B[235]), .B(n4416), .Z(n4415) );
  NANDN U5206 ( .A(A[235]), .B(n1701), .Z(n4416) );
  NANDN U5207 ( .A(n1701), .B(A[235]), .Z(n4414) );
  AND U5208 ( .A(n4417), .B(n4418), .Z(n1701) );
  NANDN U5209 ( .A(B[234]), .B(n4419), .Z(n4418) );
  NANDN U5210 ( .A(A[234]), .B(n1703), .Z(n4419) );
  NANDN U5211 ( .A(n1703), .B(A[234]), .Z(n4417) );
  AND U5212 ( .A(n4420), .B(n4421), .Z(n1703) );
  NANDN U5213 ( .A(B[233]), .B(n4422), .Z(n4421) );
  NANDN U5214 ( .A(A[233]), .B(n1705), .Z(n4422) );
  NANDN U5215 ( .A(n1705), .B(A[233]), .Z(n4420) );
  AND U5216 ( .A(n4423), .B(n4424), .Z(n1705) );
  NANDN U5217 ( .A(B[232]), .B(n4425), .Z(n4424) );
  NANDN U5218 ( .A(A[232]), .B(n1707), .Z(n4425) );
  NANDN U5219 ( .A(n1707), .B(A[232]), .Z(n4423) );
  AND U5220 ( .A(n4426), .B(n4427), .Z(n1707) );
  NANDN U5221 ( .A(B[231]), .B(n4428), .Z(n4427) );
  NANDN U5222 ( .A(A[231]), .B(n1709), .Z(n4428) );
  NANDN U5223 ( .A(n1709), .B(A[231]), .Z(n4426) );
  AND U5224 ( .A(n4429), .B(n4430), .Z(n1709) );
  NANDN U5225 ( .A(B[230]), .B(n4431), .Z(n4430) );
  NANDN U5226 ( .A(A[230]), .B(n1711), .Z(n4431) );
  NANDN U5227 ( .A(n1711), .B(A[230]), .Z(n4429) );
  AND U5228 ( .A(n4432), .B(n4433), .Z(n1711) );
  NANDN U5229 ( .A(B[229]), .B(n4434), .Z(n4433) );
  NANDN U5230 ( .A(A[229]), .B(n1715), .Z(n4434) );
  NANDN U5231 ( .A(n1715), .B(A[229]), .Z(n4432) );
  AND U5232 ( .A(n4435), .B(n4436), .Z(n1715) );
  NANDN U5233 ( .A(B[228]), .B(n4437), .Z(n4436) );
  NANDN U5234 ( .A(A[228]), .B(n1717), .Z(n4437) );
  NANDN U5235 ( .A(n1717), .B(A[228]), .Z(n4435) );
  AND U5236 ( .A(n4438), .B(n4439), .Z(n1717) );
  NANDN U5237 ( .A(B[227]), .B(n4440), .Z(n4439) );
  NANDN U5238 ( .A(A[227]), .B(n1719), .Z(n4440) );
  NANDN U5239 ( .A(n1719), .B(A[227]), .Z(n4438) );
  AND U5240 ( .A(n4441), .B(n4442), .Z(n1719) );
  NANDN U5241 ( .A(B[226]), .B(n4443), .Z(n4442) );
  NANDN U5242 ( .A(A[226]), .B(n1721), .Z(n4443) );
  NANDN U5243 ( .A(n1721), .B(A[226]), .Z(n4441) );
  AND U5244 ( .A(n4444), .B(n4445), .Z(n1721) );
  NANDN U5245 ( .A(B[225]), .B(n4446), .Z(n4445) );
  NANDN U5246 ( .A(A[225]), .B(n1723), .Z(n4446) );
  NANDN U5247 ( .A(n1723), .B(A[225]), .Z(n4444) );
  AND U5248 ( .A(n4447), .B(n4448), .Z(n1723) );
  NANDN U5249 ( .A(B[224]), .B(n4449), .Z(n4448) );
  NANDN U5250 ( .A(A[224]), .B(n1725), .Z(n4449) );
  NANDN U5251 ( .A(n1725), .B(A[224]), .Z(n4447) );
  AND U5252 ( .A(n4450), .B(n4451), .Z(n1725) );
  NANDN U5253 ( .A(B[223]), .B(n4452), .Z(n4451) );
  NANDN U5254 ( .A(A[223]), .B(n1727), .Z(n4452) );
  NANDN U5255 ( .A(n1727), .B(A[223]), .Z(n4450) );
  AND U5256 ( .A(n4453), .B(n4454), .Z(n1727) );
  NANDN U5257 ( .A(B[222]), .B(n4455), .Z(n4454) );
  NANDN U5258 ( .A(A[222]), .B(n1729), .Z(n4455) );
  NANDN U5259 ( .A(n1729), .B(A[222]), .Z(n4453) );
  AND U5260 ( .A(n4456), .B(n4457), .Z(n1729) );
  NANDN U5261 ( .A(B[221]), .B(n4458), .Z(n4457) );
  NANDN U5262 ( .A(A[221]), .B(n1731), .Z(n4458) );
  NANDN U5263 ( .A(n1731), .B(A[221]), .Z(n4456) );
  AND U5264 ( .A(n4459), .B(n4460), .Z(n1731) );
  NANDN U5265 ( .A(B[220]), .B(n4461), .Z(n4460) );
  NANDN U5266 ( .A(A[220]), .B(n1733), .Z(n4461) );
  NANDN U5267 ( .A(n1733), .B(A[220]), .Z(n4459) );
  AND U5268 ( .A(n4462), .B(n4463), .Z(n1733) );
  NANDN U5269 ( .A(B[219]), .B(n4464), .Z(n4463) );
  NANDN U5270 ( .A(A[219]), .B(n1737), .Z(n4464) );
  NANDN U5271 ( .A(n1737), .B(A[219]), .Z(n4462) );
  AND U5272 ( .A(n4465), .B(n4466), .Z(n1737) );
  NANDN U5273 ( .A(B[218]), .B(n4467), .Z(n4466) );
  NANDN U5274 ( .A(A[218]), .B(n1739), .Z(n4467) );
  NANDN U5275 ( .A(n1739), .B(A[218]), .Z(n4465) );
  AND U5276 ( .A(n4468), .B(n4469), .Z(n1739) );
  NANDN U5277 ( .A(B[217]), .B(n4470), .Z(n4469) );
  NANDN U5278 ( .A(A[217]), .B(n1741), .Z(n4470) );
  NANDN U5279 ( .A(n1741), .B(A[217]), .Z(n4468) );
  AND U5280 ( .A(n4471), .B(n4472), .Z(n1741) );
  NANDN U5281 ( .A(B[216]), .B(n4473), .Z(n4472) );
  NANDN U5282 ( .A(A[216]), .B(n1743), .Z(n4473) );
  NANDN U5283 ( .A(n1743), .B(A[216]), .Z(n4471) );
  AND U5284 ( .A(n4474), .B(n4475), .Z(n1743) );
  NANDN U5285 ( .A(B[215]), .B(n4476), .Z(n4475) );
  NANDN U5286 ( .A(A[215]), .B(n1745), .Z(n4476) );
  NANDN U5287 ( .A(n1745), .B(A[215]), .Z(n4474) );
  AND U5288 ( .A(n4477), .B(n4478), .Z(n1745) );
  NANDN U5289 ( .A(B[214]), .B(n4479), .Z(n4478) );
  NANDN U5290 ( .A(A[214]), .B(n1747), .Z(n4479) );
  NANDN U5291 ( .A(n1747), .B(A[214]), .Z(n4477) );
  AND U5292 ( .A(n4480), .B(n4481), .Z(n1747) );
  NANDN U5293 ( .A(B[213]), .B(n4482), .Z(n4481) );
  NANDN U5294 ( .A(A[213]), .B(n1749), .Z(n4482) );
  NANDN U5295 ( .A(n1749), .B(A[213]), .Z(n4480) );
  AND U5296 ( .A(n4483), .B(n4484), .Z(n1749) );
  NANDN U5297 ( .A(B[212]), .B(n4485), .Z(n4484) );
  NANDN U5298 ( .A(A[212]), .B(n1751), .Z(n4485) );
  NANDN U5299 ( .A(n1751), .B(A[212]), .Z(n4483) );
  AND U5300 ( .A(n4486), .B(n4487), .Z(n1751) );
  NANDN U5301 ( .A(B[211]), .B(n4488), .Z(n4487) );
  NANDN U5302 ( .A(A[211]), .B(n1753), .Z(n4488) );
  NANDN U5303 ( .A(n1753), .B(A[211]), .Z(n4486) );
  AND U5304 ( .A(n4489), .B(n4490), .Z(n1753) );
  NANDN U5305 ( .A(B[210]), .B(n4491), .Z(n4490) );
  NANDN U5306 ( .A(A[210]), .B(n1755), .Z(n4491) );
  NANDN U5307 ( .A(n1755), .B(A[210]), .Z(n4489) );
  AND U5308 ( .A(n4492), .B(n4493), .Z(n1755) );
  NANDN U5309 ( .A(B[209]), .B(n4494), .Z(n4493) );
  NANDN U5310 ( .A(A[209]), .B(n1759), .Z(n4494) );
  NANDN U5311 ( .A(n1759), .B(A[209]), .Z(n4492) );
  AND U5312 ( .A(n4495), .B(n4496), .Z(n1759) );
  NANDN U5313 ( .A(B[208]), .B(n4497), .Z(n4496) );
  NANDN U5314 ( .A(A[208]), .B(n1761), .Z(n4497) );
  NANDN U5315 ( .A(n1761), .B(A[208]), .Z(n4495) );
  AND U5316 ( .A(n4498), .B(n4499), .Z(n1761) );
  NANDN U5317 ( .A(B[207]), .B(n4500), .Z(n4499) );
  NANDN U5318 ( .A(A[207]), .B(n1763), .Z(n4500) );
  NANDN U5319 ( .A(n1763), .B(A[207]), .Z(n4498) );
  AND U5320 ( .A(n4501), .B(n4502), .Z(n1763) );
  NANDN U5321 ( .A(B[206]), .B(n4503), .Z(n4502) );
  NANDN U5322 ( .A(A[206]), .B(n1765), .Z(n4503) );
  NANDN U5323 ( .A(n1765), .B(A[206]), .Z(n4501) );
  AND U5324 ( .A(n4504), .B(n4505), .Z(n1765) );
  NANDN U5325 ( .A(B[205]), .B(n4506), .Z(n4505) );
  NANDN U5326 ( .A(A[205]), .B(n1767), .Z(n4506) );
  NANDN U5327 ( .A(n1767), .B(A[205]), .Z(n4504) );
  AND U5328 ( .A(n4507), .B(n4508), .Z(n1767) );
  NANDN U5329 ( .A(B[204]), .B(n4509), .Z(n4508) );
  NANDN U5330 ( .A(A[204]), .B(n1769), .Z(n4509) );
  NANDN U5331 ( .A(n1769), .B(A[204]), .Z(n4507) );
  AND U5332 ( .A(n4510), .B(n4511), .Z(n1769) );
  NANDN U5333 ( .A(B[203]), .B(n4512), .Z(n4511) );
  NANDN U5334 ( .A(A[203]), .B(n1771), .Z(n4512) );
  NANDN U5335 ( .A(n1771), .B(A[203]), .Z(n4510) );
  AND U5336 ( .A(n4513), .B(n4514), .Z(n1771) );
  NANDN U5337 ( .A(B[202]), .B(n4515), .Z(n4514) );
  NANDN U5338 ( .A(A[202]), .B(n1773), .Z(n4515) );
  NANDN U5339 ( .A(n1773), .B(A[202]), .Z(n4513) );
  AND U5340 ( .A(n4516), .B(n4517), .Z(n1773) );
  NANDN U5341 ( .A(B[201]), .B(n4518), .Z(n4517) );
  NANDN U5342 ( .A(A[201]), .B(n1775), .Z(n4518) );
  NANDN U5343 ( .A(n1775), .B(A[201]), .Z(n4516) );
  AND U5344 ( .A(n4519), .B(n4520), .Z(n1775) );
  NANDN U5345 ( .A(B[200]), .B(n4521), .Z(n4520) );
  NANDN U5346 ( .A(A[200]), .B(n1777), .Z(n4521) );
  NANDN U5347 ( .A(n1777), .B(A[200]), .Z(n4519) );
  AND U5348 ( .A(n4522), .B(n4523), .Z(n1777) );
  NANDN U5349 ( .A(B[199]), .B(n4524), .Z(n4523) );
  NANDN U5350 ( .A(A[199]), .B(n1782), .Z(n4524) );
  NANDN U5351 ( .A(n1782), .B(A[199]), .Z(n4522) );
  AND U5352 ( .A(n4525), .B(n4526), .Z(n1782) );
  NANDN U5353 ( .A(B[198]), .B(n4527), .Z(n4526) );
  NANDN U5354 ( .A(A[198]), .B(n1784), .Z(n4527) );
  NANDN U5355 ( .A(n1784), .B(A[198]), .Z(n4525) );
  AND U5356 ( .A(n4528), .B(n4529), .Z(n1784) );
  NANDN U5357 ( .A(B[197]), .B(n4530), .Z(n4529) );
  NANDN U5358 ( .A(A[197]), .B(n1786), .Z(n4530) );
  NANDN U5359 ( .A(n1786), .B(A[197]), .Z(n4528) );
  AND U5360 ( .A(n4531), .B(n4532), .Z(n1786) );
  NANDN U5361 ( .A(B[196]), .B(n4533), .Z(n4532) );
  NANDN U5362 ( .A(A[196]), .B(n1788), .Z(n4533) );
  NANDN U5363 ( .A(n1788), .B(A[196]), .Z(n4531) );
  AND U5364 ( .A(n4534), .B(n4535), .Z(n1788) );
  NANDN U5365 ( .A(B[195]), .B(n4536), .Z(n4535) );
  NANDN U5366 ( .A(A[195]), .B(n1790), .Z(n4536) );
  NANDN U5367 ( .A(n1790), .B(A[195]), .Z(n4534) );
  AND U5368 ( .A(n4537), .B(n4538), .Z(n1790) );
  NANDN U5369 ( .A(B[194]), .B(n4539), .Z(n4538) );
  NANDN U5370 ( .A(A[194]), .B(n1792), .Z(n4539) );
  NANDN U5371 ( .A(n1792), .B(A[194]), .Z(n4537) );
  AND U5372 ( .A(n4540), .B(n4541), .Z(n1792) );
  NANDN U5373 ( .A(B[193]), .B(n4542), .Z(n4541) );
  NANDN U5374 ( .A(A[193]), .B(n1794), .Z(n4542) );
  NANDN U5375 ( .A(n1794), .B(A[193]), .Z(n4540) );
  AND U5376 ( .A(n4543), .B(n4544), .Z(n1794) );
  NANDN U5377 ( .A(B[192]), .B(n4545), .Z(n4544) );
  NANDN U5378 ( .A(A[192]), .B(n1796), .Z(n4545) );
  NANDN U5379 ( .A(n1796), .B(A[192]), .Z(n4543) );
  AND U5380 ( .A(n4546), .B(n4547), .Z(n1796) );
  NANDN U5381 ( .A(B[191]), .B(n4548), .Z(n4547) );
  NANDN U5382 ( .A(A[191]), .B(n1798), .Z(n4548) );
  NANDN U5383 ( .A(n1798), .B(A[191]), .Z(n4546) );
  AND U5384 ( .A(n4549), .B(n4550), .Z(n1798) );
  NANDN U5385 ( .A(B[190]), .B(n4551), .Z(n4550) );
  NANDN U5386 ( .A(A[190]), .B(n1800), .Z(n4551) );
  NANDN U5387 ( .A(n1800), .B(A[190]), .Z(n4549) );
  AND U5388 ( .A(n4552), .B(n4553), .Z(n1800) );
  NANDN U5389 ( .A(B[189]), .B(n4554), .Z(n4553) );
  NANDN U5390 ( .A(A[189]), .B(n1804), .Z(n4554) );
  NANDN U5391 ( .A(n1804), .B(A[189]), .Z(n4552) );
  AND U5392 ( .A(n4555), .B(n4556), .Z(n1804) );
  NANDN U5393 ( .A(B[188]), .B(n4557), .Z(n4556) );
  NANDN U5394 ( .A(A[188]), .B(n1806), .Z(n4557) );
  NANDN U5395 ( .A(n1806), .B(A[188]), .Z(n4555) );
  AND U5396 ( .A(n4558), .B(n4559), .Z(n1806) );
  NANDN U5397 ( .A(B[187]), .B(n4560), .Z(n4559) );
  NANDN U5398 ( .A(A[187]), .B(n1808), .Z(n4560) );
  NANDN U5399 ( .A(n1808), .B(A[187]), .Z(n4558) );
  AND U5400 ( .A(n4561), .B(n4562), .Z(n1808) );
  NANDN U5401 ( .A(B[186]), .B(n4563), .Z(n4562) );
  NANDN U5402 ( .A(A[186]), .B(n1810), .Z(n4563) );
  NANDN U5403 ( .A(n1810), .B(A[186]), .Z(n4561) );
  AND U5404 ( .A(n4564), .B(n4565), .Z(n1810) );
  NANDN U5405 ( .A(B[185]), .B(n4566), .Z(n4565) );
  NANDN U5406 ( .A(A[185]), .B(n1812), .Z(n4566) );
  NANDN U5407 ( .A(n1812), .B(A[185]), .Z(n4564) );
  AND U5408 ( .A(n4567), .B(n4568), .Z(n1812) );
  NANDN U5409 ( .A(B[184]), .B(n4569), .Z(n4568) );
  NANDN U5410 ( .A(A[184]), .B(n1814), .Z(n4569) );
  NANDN U5411 ( .A(n1814), .B(A[184]), .Z(n4567) );
  AND U5412 ( .A(n4570), .B(n4571), .Z(n1814) );
  NANDN U5413 ( .A(B[183]), .B(n4572), .Z(n4571) );
  NANDN U5414 ( .A(A[183]), .B(n1816), .Z(n4572) );
  NANDN U5415 ( .A(n1816), .B(A[183]), .Z(n4570) );
  AND U5416 ( .A(n4573), .B(n4574), .Z(n1816) );
  NANDN U5417 ( .A(B[182]), .B(n4575), .Z(n4574) );
  NANDN U5418 ( .A(A[182]), .B(n1818), .Z(n4575) );
  NANDN U5419 ( .A(n1818), .B(A[182]), .Z(n4573) );
  AND U5420 ( .A(n4576), .B(n4577), .Z(n1818) );
  NANDN U5421 ( .A(B[181]), .B(n4578), .Z(n4577) );
  NANDN U5422 ( .A(A[181]), .B(n1820), .Z(n4578) );
  NANDN U5423 ( .A(n1820), .B(A[181]), .Z(n4576) );
  AND U5424 ( .A(n4579), .B(n4580), .Z(n1820) );
  NANDN U5425 ( .A(B[180]), .B(n4581), .Z(n4580) );
  NANDN U5426 ( .A(A[180]), .B(n1822), .Z(n4581) );
  NANDN U5427 ( .A(n1822), .B(A[180]), .Z(n4579) );
  AND U5428 ( .A(n4582), .B(n4583), .Z(n1822) );
  NANDN U5429 ( .A(B[179]), .B(n4584), .Z(n4583) );
  NANDN U5430 ( .A(A[179]), .B(n1826), .Z(n4584) );
  NANDN U5431 ( .A(n1826), .B(A[179]), .Z(n4582) );
  AND U5432 ( .A(n4585), .B(n4586), .Z(n1826) );
  NANDN U5433 ( .A(B[178]), .B(n4587), .Z(n4586) );
  NANDN U5434 ( .A(A[178]), .B(n1828), .Z(n4587) );
  NANDN U5435 ( .A(n1828), .B(A[178]), .Z(n4585) );
  AND U5436 ( .A(n4588), .B(n4589), .Z(n1828) );
  NANDN U5437 ( .A(B[177]), .B(n4590), .Z(n4589) );
  NANDN U5438 ( .A(A[177]), .B(n1830), .Z(n4590) );
  NANDN U5439 ( .A(n1830), .B(A[177]), .Z(n4588) );
  AND U5440 ( .A(n4591), .B(n4592), .Z(n1830) );
  NANDN U5441 ( .A(B[176]), .B(n4593), .Z(n4592) );
  NANDN U5442 ( .A(A[176]), .B(n1832), .Z(n4593) );
  NANDN U5443 ( .A(n1832), .B(A[176]), .Z(n4591) );
  AND U5444 ( .A(n4594), .B(n4595), .Z(n1832) );
  NANDN U5445 ( .A(B[175]), .B(n4596), .Z(n4595) );
  NANDN U5446 ( .A(A[175]), .B(n1834), .Z(n4596) );
  NANDN U5447 ( .A(n1834), .B(A[175]), .Z(n4594) );
  AND U5448 ( .A(n4597), .B(n4598), .Z(n1834) );
  NANDN U5449 ( .A(B[174]), .B(n4599), .Z(n4598) );
  NANDN U5450 ( .A(A[174]), .B(n1836), .Z(n4599) );
  NANDN U5451 ( .A(n1836), .B(A[174]), .Z(n4597) );
  AND U5452 ( .A(n4600), .B(n4601), .Z(n1836) );
  NANDN U5453 ( .A(B[173]), .B(n4602), .Z(n4601) );
  NANDN U5454 ( .A(A[173]), .B(n1838), .Z(n4602) );
  NANDN U5455 ( .A(n1838), .B(A[173]), .Z(n4600) );
  AND U5456 ( .A(n4603), .B(n4604), .Z(n1838) );
  NANDN U5457 ( .A(B[172]), .B(n4605), .Z(n4604) );
  NANDN U5458 ( .A(A[172]), .B(n1840), .Z(n4605) );
  NANDN U5459 ( .A(n1840), .B(A[172]), .Z(n4603) );
  AND U5460 ( .A(n4606), .B(n4607), .Z(n1840) );
  NANDN U5461 ( .A(B[171]), .B(n4608), .Z(n4607) );
  NANDN U5462 ( .A(A[171]), .B(n1842), .Z(n4608) );
  NANDN U5463 ( .A(n1842), .B(A[171]), .Z(n4606) );
  AND U5464 ( .A(n4609), .B(n4610), .Z(n1842) );
  NANDN U5465 ( .A(B[170]), .B(n4611), .Z(n4610) );
  NANDN U5466 ( .A(A[170]), .B(n1844), .Z(n4611) );
  NANDN U5467 ( .A(n1844), .B(A[170]), .Z(n4609) );
  AND U5468 ( .A(n4612), .B(n4613), .Z(n1844) );
  NANDN U5469 ( .A(B[169]), .B(n4614), .Z(n4613) );
  NANDN U5470 ( .A(A[169]), .B(n1848), .Z(n4614) );
  NANDN U5471 ( .A(n1848), .B(A[169]), .Z(n4612) );
  AND U5472 ( .A(n4615), .B(n4616), .Z(n1848) );
  NANDN U5473 ( .A(B[168]), .B(n4617), .Z(n4616) );
  NANDN U5474 ( .A(A[168]), .B(n1850), .Z(n4617) );
  NANDN U5475 ( .A(n1850), .B(A[168]), .Z(n4615) );
  AND U5476 ( .A(n4618), .B(n4619), .Z(n1850) );
  NANDN U5477 ( .A(B[167]), .B(n4620), .Z(n4619) );
  NANDN U5478 ( .A(A[167]), .B(n1852), .Z(n4620) );
  NANDN U5479 ( .A(n1852), .B(A[167]), .Z(n4618) );
  AND U5480 ( .A(n4621), .B(n4622), .Z(n1852) );
  NANDN U5481 ( .A(B[166]), .B(n4623), .Z(n4622) );
  NANDN U5482 ( .A(A[166]), .B(n1854), .Z(n4623) );
  NANDN U5483 ( .A(n1854), .B(A[166]), .Z(n4621) );
  AND U5484 ( .A(n4624), .B(n4625), .Z(n1854) );
  NANDN U5485 ( .A(B[165]), .B(n4626), .Z(n4625) );
  NANDN U5486 ( .A(A[165]), .B(n1856), .Z(n4626) );
  NANDN U5487 ( .A(n1856), .B(A[165]), .Z(n4624) );
  AND U5488 ( .A(n4627), .B(n4628), .Z(n1856) );
  NANDN U5489 ( .A(B[164]), .B(n4629), .Z(n4628) );
  NANDN U5490 ( .A(A[164]), .B(n1858), .Z(n4629) );
  NANDN U5491 ( .A(n1858), .B(A[164]), .Z(n4627) );
  AND U5492 ( .A(n4630), .B(n4631), .Z(n1858) );
  NANDN U5493 ( .A(B[163]), .B(n4632), .Z(n4631) );
  NANDN U5494 ( .A(A[163]), .B(n1860), .Z(n4632) );
  NANDN U5495 ( .A(n1860), .B(A[163]), .Z(n4630) );
  AND U5496 ( .A(n4633), .B(n4634), .Z(n1860) );
  NANDN U5497 ( .A(B[162]), .B(n4635), .Z(n4634) );
  NANDN U5498 ( .A(A[162]), .B(n1862), .Z(n4635) );
  NANDN U5499 ( .A(n1862), .B(A[162]), .Z(n4633) );
  AND U5500 ( .A(n4636), .B(n4637), .Z(n1862) );
  NANDN U5501 ( .A(B[161]), .B(n4638), .Z(n4637) );
  NANDN U5502 ( .A(A[161]), .B(n1864), .Z(n4638) );
  NANDN U5503 ( .A(n1864), .B(A[161]), .Z(n4636) );
  AND U5504 ( .A(n4639), .B(n4640), .Z(n1864) );
  NANDN U5505 ( .A(B[160]), .B(n4641), .Z(n4640) );
  NANDN U5506 ( .A(A[160]), .B(n1866), .Z(n4641) );
  NANDN U5507 ( .A(n1866), .B(A[160]), .Z(n4639) );
  AND U5508 ( .A(n4642), .B(n4643), .Z(n1866) );
  NANDN U5509 ( .A(B[159]), .B(n4644), .Z(n4643) );
  NANDN U5510 ( .A(A[159]), .B(n1870), .Z(n4644) );
  NANDN U5511 ( .A(n1870), .B(A[159]), .Z(n4642) );
  AND U5512 ( .A(n4645), .B(n4646), .Z(n1870) );
  NANDN U5513 ( .A(B[158]), .B(n4647), .Z(n4646) );
  NANDN U5514 ( .A(A[158]), .B(n1872), .Z(n4647) );
  NANDN U5515 ( .A(n1872), .B(A[158]), .Z(n4645) );
  AND U5516 ( .A(n4648), .B(n4649), .Z(n1872) );
  NANDN U5517 ( .A(B[157]), .B(n4650), .Z(n4649) );
  NANDN U5518 ( .A(A[157]), .B(n1874), .Z(n4650) );
  NANDN U5519 ( .A(n1874), .B(A[157]), .Z(n4648) );
  AND U5520 ( .A(n4651), .B(n4652), .Z(n1874) );
  NANDN U5521 ( .A(B[156]), .B(n4653), .Z(n4652) );
  NANDN U5522 ( .A(A[156]), .B(n1876), .Z(n4653) );
  NANDN U5523 ( .A(n1876), .B(A[156]), .Z(n4651) );
  AND U5524 ( .A(n4654), .B(n4655), .Z(n1876) );
  NANDN U5525 ( .A(B[155]), .B(n4656), .Z(n4655) );
  NANDN U5526 ( .A(A[155]), .B(n1878), .Z(n4656) );
  NANDN U5527 ( .A(n1878), .B(A[155]), .Z(n4654) );
  AND U5528 ( .A(n4657), .B(n4658), .Z(n1878) );
  NANDN U5529 ( .A(B[154]), .B(n4659), .Z(n4658) );
  NANDN U5530 ( .A(A[154]), .B(n1880), .Z(n4659) );
  NANDN U5531 ( .A(n1880), .B(A[154]), .Z(n4657) );
  AND U5532 ( .A(n4660), .B(n4661), .Z(n1880) );
  NANDN U5533 ( .A(B[153]), .B(n4662), .Z(n4661) );
  NANDN U5534 ( .A(A[153]), .B(n1882), .Z(n4662) );
  NANDN U5535 ( .A(n1882), .B(A[153]), .Z(n4660) );
  AND U5536 ( .A(n4663), .B(n4664), .Z(n1882) );
  NANDN U5537 ( .A(B[152]), .B(n4665), .Z(n4664) );
  NANDN U5538 ( .A(A[152]), .B(n1884), .Z(n4665) );
  NANDN U5539 ( .A(n1884), .B(A[152]), .Z(n4663) );
  AND U5540 ( .A(n4666), .B(n4667), .Z(n1884) );
  NANDN U5541 ( .A(B[151]), .B(n4668), .Z(n4667) );
  NANDN U5542 ( .A(A[151]), .B(n1886), .Z(n4668) );
  NANDN U5543 ( .A(n1886), .B(A[151]), .Z(n4666) );
  AND U5544 ( .A(n4669), .B(n4670), .Z(n1886) );
  NANDN U5545 ( .A(B[150]), .B(n4671), .Z(n4670) );
  NANDN U5546 ( .A(A[150]), .B(n1888), .Z(n4671) );
  NANDN U5547 ( .A(n1888), .B(A[150]), .Z(n4669) );
  AND U5548 ( .A(n4672), .B(n4673), .Z(n1888) );
  NANDN U5549 ( .A(B[149]), .B(n4674), .Z(n4673) );
  NANDN U5550 ( .A(A[149]), .B(n1892), .Z(n4674) );
  NANDN U5551 ( .A(n1892), .B(A[149]), .Z(n4672) );
  AND U5552 ( .A(n4675), .B(n4676), .Z(n1892) );
  NANDN U5553 ( .A(B[148]), .B(n4677), .Z(n4676) );
  NANDN U5554 ( .A(A[148]), .B(n1894), .Z(n4677) );
  NANDN U5555 ( .A(n1894), .B(A[148]), .Z(n4675) );
  AND U5556 ( .A(n4678), .B(n4679), .Z(n1894) );
  NANDN U5557 ( .A(B[147]), .B(n4680), .Z(n4679) );
  NANDN U5558 ( .A(A[147]), .B(n1896), .Z(n4680) );
  NANDN U5559 ( .A(n1896), .B(A[147]), .Z(n4678) );
  AND U5560 ( .A(n4681), .B(n4682), .Z(n1896) );
  NANDN U5561 ( .A(B[146]), .B(n4683), .Z(n4682) );
  NANDN U5562 ( .A(A[146]), .B(n1898), .Z(n4683) );
  NANDN U5563 ( .A(n1898), .B(A[146]), .Z(n4681) );
  AND U5564 ( .A(n4684), .B(n4685), .Z(n1898) );
  NANDN U5565 ( .A(B[145]), .B(n4686), .Z(n4685) );
  NANDN U5566 ( .A(A[145]), .B(n1900), .Z(n4686) );
  NANDN U5567 ( .A(n1900), .B(A[145]), .Z(n4684) );
  AND U5568 ( .A(n4687), .B(n4688), .Z(n1900) );
  NANDN U5569 ( .A(B[144]), .B(n4689), .Z(n4688) );
  NANDN U5570 ( .A(A[144]), .B(n1902), .Z(n4689) );
  NANDN U5571 ( .A(n1902), .B(A[144]), .Z(n4687) );
  AND U5572 ( .A(n4690), .B(n4691), .Z(n1902) );
  NANDN U5573 ( .A(B[143]), .B(n4692), .Z(n4691) );
  NANDN U5574 ( .A(A[143]), .B(n1904), .Z(n4692) );
  NANDN U5575 ( .A(n1904), .B(A[143]), .Z(n4690) );
  AND U5576 ( .A(n4693), .B(n4694), .Z(n1904) );
  NANDN U5577 ( .A(B[142]), .B(n4695), .Z(n4694) );
  NANDN U5578 ( .A(A[142]), .B(n1906), .Z(n4695) );
  NANDN U5579 ( .A(n1906), .B(A[142]), .Z(n4693) );
  AND U5580 ( .A(n4696), .B(n4697), .Z(n1906) );
  NANDN U5581 ( .A(B[141]), .B(n4698), .Z(n4697) );
  NANDN U5582 ( .A(A[141]), .B(n1908), .Z(n4698) );
  NANDN U5583 ( .A(n1908), .B(A[141]), .Z(n4696) );
  AND U5584 ( .A(n4699), .B(n4700), .Z(n1908) );
  NANDN U5585 ( .A(B[140]), .B(n4701), .Z(n4700) );
  NANDN U5586 ( .A(A[140]), .B(n1910), .Z(n4701) );
  NANDN U5587 ( .A(n1910), .B(A[140]), .Z(n4699) );
  AND U5588 ( .A(n4702), .B(n4703), .Z(n1910) );
  NANDN U5589 ( .A(B[139]), .B(n4704), .Z(n4703) );
  NANDN U5590 ( .A(A[139]), .B(n1914), .Z(n4704) );
  NANDN U5591 ( .A(n1914), .B(A[139]), .Z(n4702) );
  AND U5592 ( .A(n4705), .B(n4706), .Z(n1914) );
  NANDN U5593 ( .A(B[138]), .B(n4707), .Z(n4706) );
  NANDN U5594 ( .A(A[138]), .B(n1916), .Z(n4707) );
  NANDN U5595 ( .A(n1916), .B(A[138]), .Z(n4705) );
  AND U5596 ( .A(n4708), .B(n4709), .Z(n1916) );
  NANDN U5597 ( .A(B[137]), .B(n4710), .Z(n4709) );
  NANDN U5598 ( .A(A[137]), .B(n1918), .Z(n4710) );
  NANDN U5599 ( .A(n1918), .B(A[137]), .Z(n4708) );
  AND U5600 ( .A(n4711), .B(n4712), .Z(n1918) );
  NANDN U5601 ( .A(B[136]), .B(n4713), .Z(n4712) );
  NANDN U5602 ( .A(A[136]), .B(n1920), .Z(n4713) );
  NANDN U5603 ( .A(n1920), .B(A[136]), .Z(n4711) );
  AND U5604 ( .A(n4714), .B(n4715), .Z(n1920) );
  NANDN U5605 ( .A(B[135]), .B(n4716), .Z(n4715) );
  NANDN U5606 ( .A(A[135]), .B(n1922), .Z(n4716) );
  NANDN U5607 ( .A(n1922), .B(A[135]), .Z(n4714) );
  AND U5608 ( .A(n4717), .B(n4718), .Z(n1922) );
  NANDN U5609 ( .A(B[134]), .B(n4719), .Z(n4718) );
  NANDN U5610 ( .A(A[134]), .B(n1924), .Z(n4719) );
  NANDN U5611 ( .A(n1924), .B(A[134]), .Z(n4717) );
  AND U5612 ( .A(n4720), .B(n4721), .Z(n1924) );
  NANDN U5613 ( .A(B[133]), .B(n4722), .Z(n4721) );
  NANDN U5614 ( .A(A[133]), .B(n1926), .Z(n4722) );
  NANDN U5615 ( .A(n1926), .B(A[133]), .Z(n4720) );
  AND U5616 ( .A(n4723), .B(n4724), .Z(n1926) );
  NANDN U5617 ( .A(B[132]), .B(n4725), .Z(n4724) );
  NANDN U5618 ( .A(A[132]), .B(n1928), .Z(n4725) );
  NANDN U5619 ( .A(n1928), .B(A[132]), .Z(n4723) );
  AND U5620 ( .A(n4726), .B(n4727), .Z(n1928) );
  NANDN U5621 ( .A(B[131]), .B(n4728), .Z(n4727) );
  NANDN U5622 ( .A(A[131]), .B(n1930), .Z(n4728) );
  NANDN U5623 ( .A(n1930), .B(A[131]), .Z(n4726) );
  AND U5624 ( .A(n4729), .B(n4730), .Z(n1930) );
  NANDN U5625 ( .A(B[130]), .B(n4731), .Z(n4730) );
  NANDN U5626 ( .A(A[130]), .B(n1932), .Z(n4731) );
  NANDN U5627 ( .A(n1932), .B(A[130]), .Z(n4729) );
  AND U5628 ( .A(n4732), .B(n4733), .Z(n1932) );
  NANDN U5629 ( .A(B[129]), .B(n4734), .Z(n4733) );
  NANDN U5630 ( .A(A[129]), .B(n1936), .Z(n4734) );
  NANDN U5631 ( .A(n1936), .B(A[129]), .Z(n4732) );
  AND U5632 ( .A(n4735), .B(n4736), .Z(n1936) );
  NANDN U5633 ( .A(B[128]), .B(n4737), .Z(n4736) );
  NANDN U5634 ( .A(A[128]), .B(n1938), .Z(n4737) );
  NANDN U5635 ( .A(n1938), .B(A[128]), .Z(n4735) );
  AND U5636 ( .A(n4738), .B(n4739), .Z(n1938) );
  NANDN U5637 ( .A(B[127]), .B(n4740), .Z(n4739) );
  NANDN U5638 ( .A(A[127]), .B(n1940), .Z(n4740) );
  NANDN U5639 ( .A(n1940), .B(A[127]), .Z(n4738) );
  AND U5640 ( .A(n4741), .B(n4742), .Z(n1940) );
  NANDN U5641 ( .A(B[126]), .B(n4743), .Z(n4742) );
  NANDN U5642 ( .A(A[126]), .B(n1942), .Z(n4743) );
  NANDN U5643 ( .A(n1942), .B(A[126]), .Z(n4741) );
  AND U5644 ( .A(n4744), .B(n4745), .Z(n1942) );
  NANDN U5645 ( .A(B[125]), .B(n4746), .Z(n4745) );
  NANDN U5646 ( .A(A[125]), .B(n1944), .Z(n4746) );
  NANDN U5647 ( .A(n1944), .B(A[125]), .Z(n4744) );
  AND U5648 ( .A(n4747), .B(n4748), .Z(n1944) );
  NANDN U5649 ( .A(B[124]), .B(n4749), .Z(n4748) );
  NANDN U5650 ( .A(A[124]), .B(n1946), .Z(n4749) );
  NANDN U5651 ( .A(n1946), .B(A[124]), .Z(n4747) );
  AND U5652 ( .A(n4750), .B(n4751), .Z(n1946) );
  NANDN U5653 ( .A(B[123]), .B(n4752), .Z(n4751) );
  NANDN U5654 ( .A(A[123]), .B(n1948), .Z(n4752) );
  NANDN U5655 ( .A(n1948), .B(A[123]), .Z(n4750) );
  AND U5656 ( .A(n4753), .B(n4754), .Z(n1948) );
  NANDN U5657 ( .A(B[122]), .B(n4755), .Z(n4754) );
  NANDN U5658 ( .A(A[122]), .B(n1950), .Z(n4755) );
  NANDN U5659 ( .A(n1950), .B(A[122]), .Z(n4753) );
  AND U5660 ( .A(n4756), .B(n4757), .Z(n1950) );
  NANDN U5661 ( .A(B[121]), .B(n4758), .Z(n4757) );
  NANDN U5662 ( .A(A[121]), .B(n1952), .Z(n4758) );
  NANDN U5663 ( .A(n1952), .B(A[121]), .Z(n4756) );
  AND U5664 ( .A(n4759), .B(n4760), .Z(n1952) );
  NANDN U5665 ( .A(B[120]), .B(n4761), .Z(n4760) );
  NANDN U5666 ( .A(A[120]), .B(n1954), .Z(n4761) );
  NANDN U5667 ( .A(n1954), .B(A[120]), .Z(n4759) );
  AND U5668 ( .A(n4762), .B(n4763), .Z(n1954) );
  NANDN U5669 ( .A(B[119]), .B(n4764), .Z(n4763) );
  NANDN U5670 ( .A(A[119]), .B(n1958), .Z(n4764) );
  NANDN U5671 ( .A(n1958), .B(A[119]), .Z(n4762) );
  AND U5672 ( .A(n4765), .B(n4766), .Z(n1958) );
  NANDN U5673 ( .A(B[118]), .B(n4767), .Z(n4766) );
  NANDN U5674 ( .A(A[118]), .B(n1960), .Z(n4767) );
  NANDN U5675 ( .A(n1960), .B(A[118]), .Z(n4765) );
  AND U5676 ( .A(n4768), .B(n4769), .Z(n1960) );
  NANDN U5677 ( .A(B[117]), .B(n4770), .Z(n4769) );
  NANDN U5678 ( .A(A[117]), .B(n1962), .Z(n4770) );
  NANDN U5679 ( .A(n1962), .B(A[117]), .Z(n4768) );
  AND U5680 ( .A(n4771), .B(n4772), .Z(n1962) );
  NANDN U5681 ( .A(B[116]), .B(n4773), .Z(n4772) );
  NANDN U5682 ( .A(A[116]), .B(n1964), .Z(n4773) );
  NANDN U5683 ( .A(n1964), .B(A[116]), .Z(n4771) );
  AND U5684 ( .A(n4774), .B(n4775), .Z(n1964) );
  NANDN U5685 ( .A(B[115]), .B(n4776), .Z(n4775) );
  NANDN U5686 ( .A(A[115]), .B(n1966), .Z(n4776) );
  NANDN U5687 ( .A(n1966), .B(A[115]), .Z(n4774) );
  AND U5688 ( .A(n4777), .B(n4778), .Z(n1966) );
  NANDN U5689 ( .A(B[114]), .B(n4779), .Z(n4778) );
  NANDN U5690 ( .A(A[114]), .B(n1968), .Z(n4779) );
  NANDN U5691 ( .A(n1968), .B(A[114]), .Z(n4777) );
  AND U5692 ( .A(n4780), .B(n4781), .Z(n1968) );
  NANDN U5693 ( .A(B[113]), .B(n4782), .Z(n4781) );
  NANDN U5694 ( .A(A[113]), .B(n1970), .Z(n4782) );
  NANDN U5695 ( .A(n1970), .B(A[113]), .Z(n4780) );
  AND U5696 ( .A(n4783), .B(n4784), .Z(n1970) );
  NANDN U5697 ( .A(B[112]), .B(n4785), .Z(n4784) );
  NANDN U5698 ( .A(A[112]), .B(n1972), .Z(n4785) );
  NANDN U5699 ( .A(n1972), .B(A[112]), .Z(n4783) );
  AND U5700 ( .A(n4786), .B(n4787), .Z(n1972) );
  NANDN U5701 ( .A(B[111]), .B(n4788), .Z(n4787) );
  NANDN U5702 ( .A(A[111]), .B(n1974), .Z(n4788) );
  NANDN U5703 ( .A(n1974), .B(A[111]), .Z(n4786) );
  AND U5704 ( .A(n4789), .B(n4790), .Z(n1974) );
  NANDN U5705 ( .A(B[110]), .B(n4791), .Z(n4790) );
  NANDN U5706 ( .A(A[110]), .B(n1976), .Z(n4791) );
  NANDN U5707 ( .A(n1976), .B(A[110]), .Z(n4789) );
  AND U5708 ( .A(n4792), .B(n4793), .Z(n1976) );
  NANDN U5709 ( .A(B[109]), .B(n4794), .Z(n4793) );
  NANDN U5710 ( .A(A[109]), .B(n1980), .Z(n4794) );
  NANDN U5711 ( .A(n1980), .B(A[109]), .Z(n4792) );
  AND U5712 ( .A(n4795), .B(n4796), .Z(n1980) );
  NANDN U5713 ( .A(B[108]), .B(n4797), .Z(n4796) );
  NANDN U5714 ( .A(A[108]), .B(n1982), .Z(n4797) );
  NANDN U5715 ( .A(n1982), .B(A[108]), .Z(n4795) );
  AND U5716 ( .A(n4798), .B(n4799), .Z(n1982) );
  NANDN U5717 ( .A(B[107]), .B(n4800), .Z(n4799) );
  NANDN U5718 ( .A(A[107]), .B(n1984), .Z(n4800) );
  NANDN U5719 ( .A(n1984), .B(A[107]), .Z(n4798) );
  AND U5720 ( .A(n4801), .B(n4802), .Z(n1984) );
  NANDN U5721 ( .A(B[106]), .B(n4803), .Z(n4802) );
  NANDN U5722 ( .A(A[106]), .B(n1986), .Z(n4803) );
  NANDN U5723 ( .A(n1986), .B(A[106]), .Z(n4801) );
  AND U5724 ( .A(n4804), .B(n4805), .Z(n1986) );
  NANDN U5725 ( .A(B[105]), .B(n4806), .Z(n4805) );
  NANDN U5726 ( .A(A[105]), .B(n1988), .Z(n4806) );
  NANDN U5727 ( .A(n1988), .B(A[105]), .Z(n4804) );
  AND U5728 ( .A(n4807), .B(n4808), .Z(n1988) );
  NANDN U5729 ( .A(B[104]), .B(n4809), .Z(n4808) );
  NANDN U5730 ( .A(A[104]), .B(n1990), .Z(n4809) );
  NANDN U5731 ( .A(n1990), .B(A[104]), .Z(n4807) );
  AND U5732 ( .A(n4810), .B(n4811), .Z(n1990) );
  NANDN U5733 ( .A(B[103]), .B(n4812), .Z(n4811) );
  NANDN U5734 ( .A(A[103]), .B(n1992), .Z(n4812) );
  NANDN U5735 ( .A(n1992), .B(A[103]), .Z(n4810) );
  AND U5736 ( .A(n4813), .B(n4814), .Z(n1992) );
  NANDN U5737 ( .A(B[102]), .B(n4815), .Z(n4814) );
  NANDN U5738 ( .A(A[102]), .B(n1994), .Z(n4815) );
  NANDN U5739 ( .A(n1994), .B(A[102]), .Z(n4813) );
  AND U5740 ( .A(n4816), .B(n4817), .Z(n1994) );
  NANDN U5741 ( .A(B[101]), .B(n4818), .Z(n4817) );
  NANDN U5742 ( .A(A[101]), .B(n2022), .Z(n4818) );
  NANDN U5743 ( .A(n2022), .B(A[101]), .Z(n4816) );
  AND U5744 ( .A(n4819), .B(n4820), .Z(n2022) );
  NANDN U5745 ( .A(B[100]), .B(n4821), .Z(n4820) );
  NANDN U5746 ( .A(A[100]), .B(n2074), .Z(n4821) );
  NANDN U5747 ( .A(n2074), .B(A[100]), .Z(n4819) );
  AND U5748 ( .A(n4822), .B(n4823), .Z(n2074) );
  NANDN U5749 ( .A(B[99]), .B(n4824), .Z(n4823) );
  OR U5750 ( .A(n5), .B(A[99]), .Z(n4824) );
  NAND U5751 ( .A(A[99]), .B(n5), .Z(n4822) );
  NAND U5752 ( .A(n4825), .B(n4826), .Z(n5) );
  NANDN U5753 ( .A(B[98]), .B(n4827), .Z(n4826) );
  NANDN U5754 ( .A(A[98]), .B(n27), .Z(n4827) );
  NANDN U5755 ( .A(n27), .B(A[98]), .Z(n4825) );
  AND U5756 ( .A(n4828), .B(n4829), .Z(n27) );
  NANDN U5757 ( .A(B[97]), .B(n4830), .Z(n4829) );
  NANDN U5758 ( .A(A[97]), .B(n49), .Z(n4830) );
  NANDN U5759 ( .A(n49), .B(A[97]), .Z(n4828) );
  AND U5760 ( .A(n4831), .B(n4832), .Z(n49) );
  NANDN U5761 ( .A(B[96]), .B(n4833), .Z(n4832) );
  NANDN U5762 ( .A(A[96]), .B(n71), .Z(n4833) );
  NANDN U5763 ( .A(n71), .B(A[96]), .Z(n4831) );
  AND U5764 ( .A(n4834), .B(n4835), .Z(n71) );
  NANDN U5765 ( .A(B[95]), .B(n4836), .Z(n4835) );
  NANDN U5766 ( .A(A[95]), .B(n93), .Z(n4836) );
  NANDN U5767 ( .A(n93), .B(A[95]), .Z(n4834) );
  AND U5768 ( .A(n4837), .B(n4838), .Z(n93) );
  NANDN U5769 ( .A(B[94]), .B(n4839), .Z(n4838) );
  NANDN U5770 ( .A(A[94]), .B(n115), .Z(n4839) );
  NANDN U5771 ( .A(n115), .B(A[94]), .Z(n4837) );
  AND U5772 ( .A(n4840), .B(n4841), .Z(n115) );
  NANDN U5773 ( .A(B[93]), .B(n4842), .Z(n4841) );
  NANDN U5774 ( .A(A[93]), .B(n137), .Z(n4842) );
  NANDN U5775 ( .A(n137), .B(A[93]), .Z(n4840) );
  AND U5776 ( .A(n4843), .B(n4844), .Z(n137) );
  NANDN U5777 ( .A(B[92]), .B(n4845), .Z(n4844) );
  NANDN U5778 ( .A(A[92]), .B(n159), .Z(n4845) );
  NANDN U5779 ( .A(n159), .B(A[92]), .Z(n4843) );
  AND U5780 ( .A(n4846), .B(n4847), .Z(n159) );
  NANDN U5781 ( .A(B[91]), .B(n4848), .Z(n4847) );
  NANDN U5782 ( .A(A[91]), .B(n181), .Z(n4848) );
  NANDN U5783 ( .A(n181), .B(A[91]), .Z(n4846) );
  AND U5784 ( .A(n4849), .B(n4850), .Z(n181) );
  NANDN U5785 ( .A(B[90]), .B(n4851), .Z(n4850) );
  NANDN U5786 ( .A(A[90]), .B(n203), .Z(n4851) );
  NANDN U5787 ( .A(n203), .B(A[90]), .Z(n4849) );
  AND U5788 ( .A(n4852), .B(n4853), .Z(n203) );
  NANDN U5789 ( .A(B[89]), .B(n4854), .Z(n4853) );
  NANDN U5790 ( .A(A[89]), .B(n227), .Z(n4854) );
  NANDN U5791 ( .A(n227), .B(A[89]), .Z(n4852) );
  AND U5792 ( .A(n4855), .B(n4856), .Z(n227) );
  NANDN U5793 ( .A(B[88]), .B(n4857), .Z(n4856) );
  NANDN U5794 ( .A(A[88]), .B(n249), .Z(n4857) );
  NANDN U5795 ( .A(n249), .B(A[88]), .Z(n4855) );
  AND U5796 ( .A(n4858), .B(n4859), .Z(n249) );
  NANDN U5797 ( .A(B[87]), .B(n4860), .Z(n4859) );
  NANDN U5798 ( .A(A[87]), .B(n271), .Z(n4860) );
  NANDN U5799 ( .A(n271), .B(A[87]), .Z(n4858) );
  AND U5800 ( .A(n4861), .B(n4862), .Z(n271) );
  NANDN U5801 ( .A(B[86]), .B(n4863), .Z(n4862) );
  NANDN U5802 ( .A(A[86]), .B(n293), .Z(n4863) );
  NANDN U5803 ( .A(n293), .B(A[86]), .Z(n4861) );
  AND U5804 ( .A(n4864), .B(n4865), .Z(n293) );
  NANDN U5805 ( .A(B[85]), .B(n4866), .Z(n4865) );
  NANDN U5806 ( .A(A[85]), .B(n315), .Z(n4866) );
  NANDN U5807 ( .A(n315), .B(A[85]), .Z(n4864) );
  AND U5808 ( .A(n4867), .B(n4868), .Z(n315) );
  NANDN U5809 ( .A(B[84]), .B(n4869), .Z(n4868) );
  NANDN U5810 ( .A(A[84]), .B(n337), .Z(n4869) );
  NANDN U5811 ( .A(n337), .B(A[84]), .Z(n4867) );
  AND U5812 ( .A(n4870), .B(n4871), .Z(n337) );
  NANDN U5813 ( .A(B[83]), .B(n4872), .Z(n4871) );
  NANDN U5814 ( .A(A[83]), .B(n359), .Z(n4872) );
  NANDN U5815 ( .A(n359), .B(A[83]), .Z(n4870) );
  AND U5816 ( .A(n4873), .B(n4874), .Z(n359) );
  NANDN U5817 ( .A(B[82]), .B(n4875), .Z(n4874) );
  NANDN U5818 ( .A(A[82]), .B(n381), .Z(n4875) );
  NANDN U5819 ( .A(n381), .B(A[82]), .Z(n4873) );
  AND U5820 ( .A(n4876), .B(n4877), .Z(n381) );
  NANDN U5821 ( .A(B[81]), .B(n4878), .Z(n4877) );
  NANDN U5822 ( .A(A[81]), .B(n403), .Z(n4878) );
  NANDN U5823 ( .A(n403), .B(A[81]), .Z(n4876) );
  AND U5824 ( .A(n4879), .B(n4880), .Z(n403) );
  NANDN U5825 ( .A(B[80]), .B(n4881), .Z(n4880) );
  NANDN U5826 ( .A(A[80]), .B(n425), .Z(n4881) );
  NANDN U5827 ( .A(n425), .B(A[80]), .Z(n4879) );
  AND U5828 ( .A(n4882), .B(n4883), .Z(n425) );
  NANDN U5829 ( .A(B[79]), .B(n4884), .Z(n4883) );
  NANDN U5830 ( .A(A[79]), .B(n449), .Z(n4884) );
  NANDN U5831 ( .A(n449), .B(A[79]), .Z(n4882) );
  AND U5832 ( .A(n4885), .B(n4886), .Z(n449) );
  NANDN U5833 ( .A(B[78]), .B(n4887), .Z(n4886) );
  NANDN U5834 ( .A(A[78]), .B(n471), .Z(n4887) );
  NANDN U5835 ( .A(n471), .B(A[78]), .Z(n4885) );
  AND U5836 ( .A(n4888), .B(n4889), .Z(n471) );
  NANDN U5837 ( .A(B[77]), .B(n4890), .Z(n4889) );
  NANDN U5838 ( .A(A[77]), .B(n493), .Z(n4890) );
  NANDN U5839 ( .A(n493), .B(A[77]), .Z(n4888) );
  AND U5840 ( .A(n4891), .B(n4892), .Z(n493) );
  NANDN U5841 ( .A(B[76]), .B(n4893), .Z(n4892) );
  NANDN U5842 ( .A(A[76]), .B(n515), .Z(n4893) );
  NANDN U5843 ( .A(n515), .B(A[76]), .Z(n4891) );
  AND U5844 ( .A(n4894), .B(n4895), .Z(n515) );
  NANDN U5845 ( .A(B[75]), .B(n4896), .Z(n4895) );
  NANDN U5846 ( .A(A[75]), .B(n537), .Z(n4896) );
  NANDN U5847 ( .A(n537), .B(A[75]), .Z(n4894) );
  AND U5848 ( .A(n4897), .B(n4898), .Z(n537) );
  NANDN U5849 ( .A(B[74]), .B(n4899), .Z(n4898) );
  NANDN U5850 ( .A(A[74]), .B(n559), .Z(n4899) );
  NANDN U5851 ( .A(n559), .B(A[74]), .Z(n4897) );
  AND U5852 ( .A(n4900), .B(n4901), .Z(n559) );
  NANDN U5853 ( .A(B[73]), .B(n4902), .Z(n4901) );
  NANDN U5854 ( .A(A[73]), .B(n581), .Z(n4902) );
  NANDN U5855 ( .A(n581), .B(A[73]), .Z(n4900) );
  AND U5856 ( .A(n4903), .B(n4904), .Z(n581) );
  NANDN U5857 ( .A(B[72]), .B(n4905), .Z(n4904) );
  NANDN U5858 ( .A(A[72]), .B(n603), .Z(n4905) );
  NANDN U5859 ( .A(n603), .B(A[72]), .Z(n4903) );
  AND U5860 ( .A(n4906), .B(n4907), .Z(n603) );
  NANDN U5861 ( .A(B[71]), .B(n4908), .Z(n4907) );
  NANDN U5862 ( .A(A[71]), .B(n625), .Z(n4908) );
  NANDN U5863 ( .A(n625), .B(A[71]), .Z(n4906) );
  AND U5864 ( .A(n4909), .B(n4910), .Z(n625) );
  NANDN U5865 ( .A(B[70]), .B(n4911), .Z(n4910) );
  NANDN U5866 ( .A(A[70]), .B(n647), .Z(n4911) );
  NANDN U5867 ( .A(n647), .B(A[70]), .Z(n4909) );
  AND U5868 ( .A(n4912), .B(n4913), .Z(n647) );
  NANDN U5869 ( .A(B[69]), .B(n4914), .Z(n4913) );
  NANDN U5870 ( .A(A[69]), .B(n671), .Z(n4914) );
  NANDN U5871 ( .A(n671), .B(A[69]), .Z(n4912) );
  AND U5872 ( .A(n4915), .B(n4916), .Z(n671) );
  NANDN U5873 ( .A(B[68]), .B(n4917), .Z(n4916) );
  NANDN U5874 ( .A(A[68]), .B(n693), .Z(n4917) );
  NANDN U5875 ( .A(n693), .B(A[68]), .Z(n4915) );
  AND U5876 ( .A(n4918), .B(n4919), .Z(n693) );
  NANDN U5877 ( .A(B[67]), .B(n4920), .Z(n4919) );
  NANDN U5878 ( .A(A[67]), .B(n715), .Z(n4920) );
  NANDN U5879 ( .A(n715), .B(A[67]), .Z(n4918) );
  AND U5880 ( .A(n4921), .B(n4922), .Z(n715) );
  NANDN U5881 ( .A(B[66]), .B(n4923), .Z(n4922) );
  NANDN U5882 ( .A(A[66]), .B(n737), .Z(n4923) );
  NANDN U5883 ( .A(n737), .B(A[66]), .Z(n4921) );
  AND U5884 ( .A(n4924), .B(n4925), .Z(n737) );
  NANDN U5885 ( .A(B[65]), .B(n4926), .Z(n4925) );
  NANDN U5886 ( .A(A[65]), .B(n759), .Z(n4926) );
  NANDN U5887 ( .A(n759), .B(A[65]), .Z(n4924) );
  AND U5888 ( .A(n4927), .B(n4928), .Z(n759) );
  NANDN U5889 ( .A(B[64]), .B(n4929), .Z(n4928) );
  NANDN U5890 ( .A(A[64]), .B(n781), .Z(n4929) );
  NANDN U5891 ( .A(n781), .B(A[64]), .Z(n4927) );
  AND U5892 ( .A(n4930), .B(n4931), .Z(n781) );
  NANDN U5893 ( .A(B[63]), .B(n4932), .Z(n4931) );
  NANDN U5894 ( .A(A[63]), .B(n803), .Z(n4932) );
  NANDN U5895 ( .A(n803), .B(A[63]), .Z(n4930) );
  AND U5896 ( .A(n4933), .B(n4934), .Z(n803) );
  NANDN U5897 ( .A(B[62]), .B(n4935), .Z(n4934) );
  NANDN U5898 ( .A(A[62]), .B(n825), .Z(n4935) );
  NANDN U5899 ( .A(n825), .B(A[62]), .Z(n4933) );
  AND U5900 ( .A(n4936), .B(n4937), .Z(n825) );
  NANDN U5901 ( .A(B[61]), .B(n4938), .Z(n4937) );
  NANDN U5902 ( .A(A[61]), .B(n847), .Z(n4938) );
  NANDN U5903 ( .A(n847), .B(A[61]), .Z(n4936) );
  AND U5904 ( .A(n4939), .B(n4940), .Z(n847) );
  NANDN U5905 ( .A(B[60]), .B(n4941), .Z(n4940) );
  NANDN U5906 ( .A(A[60]), .B(n869), .Z(n4941) );
  NANDN U5907 ( .A(n869), .B(A[60]), .Z(n4939) );
  AND U5908 ( .A(n4942), .B(n4943), .Z(n869) );
  NANDN U5909 ( .A(B[59]), .B(n4944), .Z(n4943) );
  NANDN U5910 ( .A(A[59]), .B(n893), .Z(n4944) );
  NANDN U5911 ( .A(n893), .B(A[59]), .Z(n4942) );
  AND U5912 ( .A(n4945), .B(n4946), .Z(n893) );
  NANDN U5913 ( .A(B[58]), .B(n4947), .Z(n4946) );
  NANDN U5914 ( .A(A[58]), .B(n915), .Z(n4947) );
  NANDN U5915 ( .A(n915), .B(A[58]), .Z(n4945) );
  AND U5916 ( .A(n4948), .B(n4949), .Z(n915) );
  NANDN U5917 ( .A(B[57]), .B(n4950), .Z(n4949) );
  NANDN U5918 ( .A(A[57]), .B(n937), .Z(n4950) );
  NANDN U5919 ( .A(n937), .B(A[57]), .Z(n4948) );
  AND U5920 ( .A(n4951), .B(n4952), .Z(n937) );
  NANDN U5921 ( .A(B[56]), .B(n4953), .Z(n4952) );
  NANDN U5922 ( .A(A[56]), .B(n959), .Z(n4953) );
  NANDN U5923 ( .A(n959), .B(A[56]), .Z(n4951) );
  AND U5924 ( .A(n4954), .B(n4955), .Z(n959) );
  NANDN U5925 ( .A(B[55]), .B(n4956), .Z(n4955) );
  NANDN U5926 ( .A(A[55]), .B(n981), .Z(n4956) );
  NANDN U5927 ( .A(n981), .B(A[55]), .Z(n4954) );
  AND U5928 ( .A(n4957), .B(n4958), .Z(n981) );
  NANDN U5929 ( .A(B[54]), .B(n4959), .Z(n4958) );
  NANDN U5930 ( .A(A[54]), .B(n1003), .Z(n4959) );
  NANDN U5931 ( .A(n1003), .B(A[54]), .Z(n4957) );
  AND U5932 ( .A(n4960), .B(n4961), .Z(n1003) );
  NANDN U5933 ( .A(B[53]), .B(n4962), .Z(n4961) );
  NANDN U5934 ( .A(A[53]), .B(n1025), .Z(n4962) );
  NANDN U5935 ( .A(n1025), .B(A[53]), .Z(n4960) );
  AND U5936 ( .A(n4963), .B(n4964), .Z(n1025) );
  NANDN U5937 ( .A(B[52]), .B(n4965), .Z(n4964) );
  NANDN U5938 ( .A(A[52]), .B(n1047), .Z(n4965) );
  NANDN U5939 ( .A(n1047), .B(A[52]), .Z(n4963) );
  AND U5940 ( .A(n4966), .B(n4967), .Z(n1047) );
  NANDN U5941 ( .A(B[51]), .B(n4968), .Z(n4967) );
  NANDN U5942 ( .A(A[51]), .B(n1069), .Z(n4968) );
  NANDN U5943 ( .A(n1069), .B(A[51]), .Z(n4966) );
  AND U5944 ( .A(n4969), .B(n4970), .Z(n1069) );
  NANDN U5945 ( .A(B[50]), .B(n4971), .Z(n4970) );
  NANDN U5946 ( .A(A[50]), .B(n1091), .Z(n4971) );
  NANDN U5947 ( .A(n1091), .B(A[50]), .Z(n4969) );
  AND U5948 ( .A(n4972), .B(n4973), .Z(n1091) );
  NANDN U5949 ( .A(B[49]), .B(n4974), .Z(n4973) );
  NANDN U5950 ( .A(A[49]), .B(n1115), .Z(n4974) );
  NANDN U5951 ( .A(n1115), .B(A[49]), .Z(n4972) );
  AND U5952 ( .A(n4975), .B(n4976), .Z(n1115) );
  NANDN U5953 ( .A(B[48]), .B(n4977), .Z(n4976) );
  NANDN U5954 ( .A(A[48]), .B(n1137), .Z(n4977) );
  NANDN U5955 ( .A(n1137), .B(A[48]), .Z(n4975) );
  AND U5956 ( .A(n4978), .B(n4979), .Z(n1137) );
  NANDN U5957 ( .A(B[47]), .B(n4980), .Z(n4979) );
  NANDN U5958 ( .A(A[47]), .B(n1159), .Z(n4980) );
  NANDN U5959 ( .A(n1159), .B(A[47]), .Z(n4978) );
  AND U5960 ( .A(n4981), .B(n4982), .Z(n1159) );
  NANDN U5961 ( .A(B[46]), .B(n4983), .Z(n4982) );
  NANDN U5962 ( .A(A[46]), .B(n1181), .Z(n4983) );
  NANDN U5963 ( .A(n1181), .B(A[46]), .Z(n4981) );
  AND U5964 ( .A(n4984), .B(n4985), .Z(n1181) );
  NANDN U5965 ( .A(B[45]), .B(n4986), .Z(n4985) );
  NANDN U5966 ( .A(A[45]), .B(n1203), .Z(n4986) );
  NANDN U5967 ( .A(n1203), .B(A[45]), .Z(n4984) );
  AND U5968 ( .A(n4987), .B(n4988), .Z(n1203) );
  NANDN U5969 ( .A(B[44]), .B(n4989), .Z(n4988) );
  NANDN U5970 ( .A(A[44]), .B(n1225), .Z(n4989) );
  NANDN U5971 ( .A(n1225), .B(A[44]), .Z(n4987) );
  AND U5972 ( .A(n4990), .B(n4991), .Z(n1225) );
  NANDN U5973 ( .A(B[43]), .B(n4992), .Z(n4991) );
  NANDN U5974 ( .A(A[43]), .B(n1247), .Z(n4992) );
  NANDN U5975 ( .A(n1247), .B(A[43]), .Z(n4990) );
  AND U5976 ( .A(n4993), .B(n4994), .Z(n1247) );
  NANDN U5977 ( .A(B[42]), .B(n4995), .Z(n4994) );
  NANDN U5978 ( .A(A[42]), .B(n1269), .Z(n4995) );
  NANDN U5979 ( .A(n1269), .B(A[42]), .Z(n4993) );
  AND U5980 ( .A(n4996), .B(n4997), .Z(n1269) );
  NANDN U5981 ( .A(B[41]), .B(n4998), .Z(n4997) );
  NANDN U5982 ( .A(A[41]), .B(n1291), .Z(n4998) );
  NANDN U5983 ( .A(n1291), .B(A[41]), .Z(n4996) );
  AND U5984 ( .A(n4999), .B(n5000), .Z(n1291) );
  NANDN U5985 ( .A(B[40]), .B(n5001), .Z(n5000) );
  NANDN U5986 ( .A(A[40]), .B(n1313), .Z(n5001) );
  NANDN U5987 ( .A(n1313), .B(A[40]), .Z(n4999) );
  AND U5988 ( .A(n5002), .B(n5003), .Z(n1313) );
  NANDN U5989 ( .A(B[39]), .B(n5004), .Z(n5003) );
  NANDN U5990 ( .A(A[39]), .B(n1337), .Z(n5004) );
  NANDN U5991 ( .A(n1337), .B(A[39]), .Z(n5002) );
  AND U5992 ( .A(n5005), .B(n5006), .Z(n1337) );
  NANDN U5993 ( .A(B[38]), .B(n5007), .Z(n5006) );
  NANDN U5994 ( .A(A[38]), .B(n1359), .Z(n5007) );
  NANDN U5995 ( .A(n1359), .B(A[38]), .Z(n5005) );
  AND U5996 ( .A(n5008), .B(n5009), .Z(n1359) );
  NANDN U5997 ( .A(B[37]), .B(n5010), .Z(n5009) );
  NANDN U5998 ( .A(A[37]), .B(n1381), .Z(n5010) );
  NANDN U5999 ( .A(n1381), .B(A[37]), .Z(n5008) );
  AND U6000 ( .A(n5011), .B(n5012), .Z(n1381) );
  NANDN U6001 ( .A(B[36]), .B(n5013), .Z(n5012) );
  NANDN U6002 ( .A(A[36]), .B(n1403), .Z(n5013) );
  NANDN U6003 ( .A(n1403), .B(A[36]), .Z(n5011) );
  AND U6004 ( .A(n5014), .B(n5015), .Z(n1403) );
  NANDN U6005 ( .A(B[35]), .B(n5016), .Z(n5015) );
  NANDN U6006 ( .A(A[35]), .B(n1425), .Z(n5016) );
  NANDN U6007 ( .A(n1425), .B(A[35]), .Z(n5014) );
  AND U6008 ( .A(n5017), .B(n5018), .Z(n1425) );
  NANDN U6009 ( .A(B[34]), .B(n5019), .Z(n5018) );
  NANDN U6010 ( .A(A[34]), .B(n1447), .Z(n5019) );
  NANDN U6011 ( .A(n1447), .B(A[34]), .Z(n5017) );
  AND U6012 ( .A(n5020), .B(n5021), .Z(n1447) );
  NANDN U6013 ( .A(B[33]), .B(n5022), .Z(n5021) );
  NANDN U6014 ( .A(A[33]), .B(n1469), .Z(n5022) );
  NANDN U6015 ( .A(n1469), .B(A[33]), .Z(n5020) );
  AND U6016 ( .A(n5023), .B(n5024), .Z(n1469) );
  NANDN U6017 ( .A(B[32]), .B(n5025), .Z(n5024) );
  NANDN U6018 ( .A(A[32]), .B(n1491), .Z(n5025) );
  NANDN U6019 ( .A(n1491), .B(A[32]), .Z(n5023) );
  AND U6020 ( .A(n5026), .B(n5027), .Z(n1491) );
  NANDN U6021 ( .A(B[31]), .B(n5028), .Z(n5027) );
  NANDN U6022 ( .A(A[31]), .B(n1513), .Z(n5028) );
  NANDN U6023 ( .A(n1513), .B(A[31]), .Z(n5026) );
  AND U6024 ( .A(n5029), .B(n5030), .Z(n1513) );
  NANDN U6025 ( .A(B[30]), .B(n5031), .Z(n5030) );
  NANDN U6026 ( .A(A[30]), .B(n1535), .Z(n5031) );
  NANDN U6027 ( .A(n1535), .B(A[30]), .Z(n5029) );
  AND U6028 ( .A(n5032), .B(n5033), .Z(n1535) );
  NANDN U6029 ( .A(B[29]), .B(n5034), .Z(n5033) );
  NANDN U6030 ( .A(A[29]), .B(n1559), .Z(n5034) );
  NANDN U6031 ( .A(n1559), .B(A[29]), .Z(n5032) );
  AND U6032 ( .A(n5035), .B(n5036), .Z(n1559) );
  NANDN U6033 ( .A(B[28]), .B(n5037), .Z(n5036) );
  NANDN U6034 ( .A(A[28]), .B(n1581), .Z(n5037) );
  NANDN U6035 ( .A(n1581), .B(A[28]), .Z(n5035) );
  AND U6036 ( .A(n5038), .B(n5039), .Z(n1581) );
  NANDN U6037 ( .A(B[27]), .B(n5040), .Z(n5039) );
  NANDN U6038 ( .A(A[27]), .B(n1603), .Z(n5040) );
  NANDN U6039 ( .A(n1603), .B(A[27]), .Z(n5038) );
  AND U6040 ( .A(n5041), .B(n5042), .Z(n1603) );
  NANDN U6041 ( .A(B[26]), .B(n5043), .Z(n5042) );
  NANDN U6042 ( .A(A[26]), .B(n1625), .Z(n5043) );
  NANDN U6043 ( .A(n1625), .B(A[26]), .Z(n5041) );
  AND U6044 ( .A(n5044), .B(n5045), .Z(n1625) );
  NANDN U6045 ( .A(B[25]), .B(n5046), .Z(n5045) );
  NANDN U6046 ( .A(A[25]), .B(n1647), .Z(n5046) );
  NANDN U6047 ( .A(n1647), .B(A[25]), .Z(n5044) );
  AND U6048 ( .A(n5047), .B(n5048), .Z(n1647) );
  NANDN U6049 ( .A(B[24]), .B(n5049), .Z(n5048) );
  NANDN U6050 ( .A(A[24]), .B(n1669), .Z(n5049) );
  NANDN U6051 ( .A(n1669), .B(A[24]), .Z(n5047) );
  AND U6052 ( .A(n5050), .B(n5051), .Z(n1669) );
  NANDN U6053 ( .A(B[23]), .B(n5052), .Z(n5051) );
  NANDN U6054 ( .A(A[23]), .B(n1691), .Z(n5052) );
  NANDN U6055 ( .A(n1691), .B(A[23]), .Z(n5050) );
  AND U6056 ( .A(n5053), .B(n5054), .Z(n1691) );
  NANDN U6057 ( .A(B[22]), .B(n5055), .Z(n5054) );
  NANDN U6058 ( .A(A[22]), .B(n1713), .Z(n5055) );
  NANDN U6059 ( .A(n1713), .B(A[22]), .Z(n5053) );
  AND U6060 ( .A(n5056), .B(n5057), .Z(n1713) );
  NANDN U6061 ( .A(B[21]), .B(n5058), .Z(n5057) );
  NANDN U6062 ( .A(A[21]), .B(n1735), .Z(n5058) );
  NANDN U6063 ( .A(n1735), .B(A[21]), .Z(n5056) );
  AND U6064 ( .A(n5059), .B(n5060), .Z(n1735) );
  NANDN U6065 ( .A(B[20]), .B(n5061), .Z(n5060) );
  NANDN U6066 ( .A(A[20]), .B(n1757), .Z(n5061) );
  NANDN U6067 ( .A(n1757), .B(A[20]), .Z(n5059) );
  AND U6068 ( .A(n5062), .B(n5063), .Z(n1757) );
  NANDN U6069 ( .A(B[19]), .B(n5064), .Z(n5063) );
  NANDN U6070 ( .A(A[19]), .B(n1780), .Z(n5064) );
  NANDN U6071 ( .A(n1780), .B(A[19]), .Z(n5062) );
  AND U6072 ( .A(n5065), .B(n5066), .Z(n1780) );
  NANDN U6073 ( .A(B[18]), .B(n5067), .Z(n5066) );
  NANDN U6074 ( .A(A[18]), .B(n1802), .Z(n5067) );
  NANDN U6075 ( .A(n1802), .B(A[18]), .Z(n5065) );
  AND U6076 ( .A(n5068), .B(n5069), .Z(n1802) );
  NANDN U6077 ( .A(B[17]), .B(n5070), .Z(n5069) );
  NANDN U6078 ( .A(A[17]), .B(n1824), .Z(n5070) );
  NANDN U6079 ( .A(n1824), .B(A[17]), .Z(n5068) );
  AND U6080 ( .A(n5071), .B(n5072), .Z(n1824) );
  NANDN U6081 ( .A(B[16]), .B(n5073), .Z(n5072) );
  NANDN U6082 ( .A(A[16]), .B(n1846), .Z(n5073) );
  NANDN U6083 ( .A(n1846), .B(A[16]), .Z(n5071) );
  AND U6084 ( .A(n5074), .B(n5075), .Z(n1846) );
  NANDN U6085 ( .A(B[15]), .B(n5076), .Z(n5075) );
  NANDN U6086 ( .A(A[15]), .B(n1868), .Z(n5076) );
  NANDN U6087 ( .A(n1868), .B(A[15]), .Z(n5074) );
  AND U6088 ( .A(n5077), .B(n5078), .Z(n1868) );
  NANDN U6089 ( .A(B[14]), .B(n5079), .Z(n5078) );
  NANDN U6090 ( .A(A[14]), .B(n1890), .Z(n5079) );
  NANDN U6091 ( .A(n1890), .B(A[14]), .Z(n5077) );
  AND U6092 ( .A(n5080), .B(n5081), .Z(n1890) );
  NANDN U6093 ( .A(B[13]), .B(n5082), .Z(n5081) );
  NANDN U6094 ( .A(A[13]), .B(n1912), .Z(n5082) );
  NANDN U6095 ( .A(n1912), .B(A[13]), .Z(n5080) );
  AND U6096 ( .A(n5083), .B(n5084), .Z(n1912) );
  NANDN U6097 ( .A(B[12]), .B(n5085), .Z(n5084) );
  NANDN U6098 ( .A(A[12]), .B(n1934), .Z(n5085) );
  NANDN U6099 ( .A(n1934), .B(A[12]), .Z(n5083) );
  AND U6100 ( .A(n5086), .B(n5087), .Z(n1934) );
  NANDN U6101 ( .A(B[11]), .B(n5088), .Z(n5087) );
  NANDN U6102 ( .A(A[11]), .B(n1956), .Z(n5088) );
  NANDN U6103 ( .A(n1956), .B(A[11]), .Z(n5086) );
  AND U6104 ( .A(n5089), .B(n5090), .Z(n1956) );
  NANDN U6105 ( .A(B[10]), .B(n5091), .Z(n5090) );
  NANDN U6106 ( .A(A[10]), .B(n1978), .Z(n5091) );
  NANDN U6107 ( .A(n1978), .B(A[10]), .Z(n5089) );
  AND U6108 ( .A(n5092), .B(n5093), .Z(n1978) );
  NANDN U6109 ( .A(B[9]), .B(n5094), .Z(n5093) );
  OR U6110 ( .A(n3), .B(A[9]), .Z(n5094) );
  NAND U6111 ( .A(A[9]), .B(n3), .Z(n5092) );
  NAND U6112 ( .A(n5095), .B(n5096), .Z(n3) );
  NANDN U6113 ( .A(B[8]), .B(n5097), .Z(n5096) );
  NANDN U6114 ( .A(A[8]), .B(n225), .Z(n5097) );
  NANDN U6115 ( .A(n225), .B(A[8]), .Z(n5095) );
  AND U6116 ( .A(n5098), .B(n5099), .Z(n225) );
  NANDN U6117 ( .A(B[7]), .B(n5100), .Z(n5099) );
  NANDN U6118 ( .A(A[7]), .B(n447), .Z(n5100) );
  NANDN U6119 ( .A(n447), .B(A[7]), .Z(n5098) );
  AND U6120 ( .A(n5101), .B(n5102), .Z(n447) );
  NANDN U6121 ( .A(B[6]), .B(n5103), .Z(n5102) );
  NANDN U6122 ( .A(A[6]), .B(n669), .Z(n5103) );
  NANDN U6123 ( .A(n669), .B(A[6]), .Z(n5101) );
  AND U6124 ( .A(n5104), .B(n5105), .Z(n669) );
  NANDN U6125 ( .A(B[5]), .B(n5106), .Z(n5105) );
  NANDN U6126 ( .A(A[5]), .B(n891), .Z(n5106) );
  NANDN U6127 ( .A(n891), .B(A[5]), .Z(n5104) );
  AND U6128 ( .A(n5107), .B(n5108), .Z(n891) );
  NANDN U6129 ( .A(B[4]), .B(n5109), .Z(n5108) );
  NANDN U6130 ( .A(A[4]), .B(n1113), .Z(n5109) );
  NANDN U6131 ( .A(n1113), .B(A[4]), .Z(n5107) );
  AND U6132 ( .A(n5110), .B(n5111), .Z(n1113) );
  NANDN U6133 ( .A(B[3]), .B(n5112), .Z(n5111) );
  NANDN U6134 ( .A(A[3]), .B(n1335), .Z(n5112) );
  NANDN U6135 ( .A(n1335), .B(A[3]), .Z(n5110) );
  AND U6136 ( .A(n5113), .B(n5114), .Z(n1335) );
  NANDN U6137 ( .A(B[2]), .B(n5115), .Z(n5114) );
  NANDN U6138 ( .A(A[2]), .B(n1557), .Z(n5115) );
  NANDN U6139 ( .A(n1557), .B(A[2]), .Z(n5113) );
  AND U6140 ( .A(n5116), .B(n5117), .Z(n1557) );
  NANDN U6141 ( .A(B[1]), .B(n5118), .Z(n5117) );
  NAND U6142 ( .A(n1), .B(n2), .Z(n5118) );
  NAND U6143 ( .A(A[1]), .B(n5119), .Z(n5116) );
  NAND U6144 ( .A(n5119), .B(n5120), .Z(DIFF[0]) );
  NANDN U6145 ( .A(B[0]), .B(A[0]), .Z(n5120) );
  NANDN U6146 ( .A(A[0]), .B(B[0]), .Z(n5119) );
endmodule


module modmult_step_N1024_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [1023:0] A;
  input [0:0] B;
  output [1024:0] PRODUCT;
  input TC;


  AND U2 ( .A(A[1023]), .B(B[0]), .Z(PRODUCT[1023]) );
  AND U3 ( .A(A[1022]), .B(B[0]), .Z(PRODUCT[1022]) );
  AND U4 ( .A(A[1021]), .B(B[0]), .Z(PRODUCT[1021]) );
  AND U5 ( .A(A[1020]), .B(B[0]), .Z(PRODUCT[1020]) );
  AND U6 ( .A(A[1019]), .B(B[0]), .Z(PRODUCT[1019]) );
  AND U7 ( .A(A[1018]), .B(B[0]), .Z(PRODUCT[1018]) );
  AND U8 ( .A(A[1017]), .B(B[0]), .Z(PRODUCT[1017]) );
  AND U9 ( .A(A[1016]), .B(B[0]), .Z(PRODUCT[1016]) );
  AND U10 ( .A(A[1015]), .B(B[0]), .Z(PRODUCT[1015]) );
  AND U11 ( .A(A[1014]), .B(B[0]), .Z(PRODUCT[1014]) );
  AND U12 ( .A(A[1013]), .B(B[0]), .Z(PRODUCT[1013]) );
  AND U13 ( .A(A[1012]), .B(B[0]), .Z(PRODUCT[1012]) );
  AND U14 ( .A(A[1011]), .B(B[0]), .Z(PRODUCT[1011]) );
  AND U15 ( .A(A[1010]), .B(B[0]), .Z(PRODUCT[1010]) );
  AND U16 ( .A(A[1009]), .B(B[0]), .Z(PRODUCT[1009]) );
  AND U17 ( .A(A[1008]), .B(B[0]), .Z(PRODUCT[1008]) );
  AND U18 ( .A(A[1007]), .B(B[0]), .Z(PRODUCT[1007]) );
  AND U19 ( .A(A[1006]), .B(B[0]), .Z(PRODUCT[1006]) );
  AND U20 ( .A(A[1005]), .B(B[0]), .Z(PRODUCT[1005]) );
  AND U21 ( .A(A[1004]), .B(B[0]), .Z(PRODUCT[1004]) );
  AND U22 ( .A(A[1003]), .B(B[0]), .Z(PRODUCT[1003]) );
  AND U23 ( .A(A[1002]), .B(B[0]), .Z(PRODUCT[1002]) );
  AND U24 ( .A(A[1001]), .B(B[0]), .Z(PRODUCT[1001]) );
  AND U25 ( .A(A[1000]), .B(B[0]), .Z(PRODUCT[1000]) );
  AND U26 ( .A(A[999]), .B(B[0]), .Z(PRODUCT[999]) );
  AND U27 ( .A(A[998]), .B(B[0]), .Z(PRODUCT[998]) );
  AND U28 ( .A(A[997]), .B(B[0]), .Z(PRODUCT[997]) );
  AND U29 ( .A(A[996]), .B(B[0]), .Z(PRODUCT[996]) );
  AND U30 ( .A(A[995]), .B(B[0]), .Z(PRODUCT[995]) );
  AND U31 ( .A(A[994]), .B(B[0]), .Z(PRODUCT[994]) );
  AND U32 ( .A(A[993]), .B(B[0]), .Z(PRODUCT[993]) );
  AND U33 ( .A(A[992]), .B(B[0]), .Z(PRODUCT[992]) );
  AND U34 ( .A(A[991]), .B(B[0]), .Z(PRODUCT[991]) );
  AND U35 ( .A(A[990]), .B(B[0]), .Z(PRODUCT[990]) );
  AND U36 ( .A(A[989]), .B(B[0]), .Z(PRODUCT[989]) );
  AND U37 ( .A(A[988]), .B(B[0]), .Z(PRODUCT[988]) );
  AND U38 ( .A(A[987]), .B(B[0]), .Z(PRODUCT[987]) );
  AND U39 ( .A(A[986]), .B(B[0]), .Z(PRODUCT[986]) );
  AND U40 ( .A(A[985]), .B(B[0]), .Z(PRODUCT[985]) );
  AND U41 ( .A(A[984]), .B(B[0]), .Z(PRODUCT[984]) );
  AND U42 ( .A(A[983]), .B(B[0]), .Z(PRODUCT[983]) );
  AND U43 ( .A(A[982]), .B(B[0]), .Z(PRODUCT[982]) );
  AND U44 ( .A(A[981]), .B(B[0]), .Z(PRODUCT[981]) );
  AND U45 ( .A(A[980]), .B(B[0]), .Z(PRODUCT[980]) );
  AND U46 ( .A(A[979]), .B(B[0]), .Z(PRODUCT[979]) );
  AND U47 ( .A(A[978]), .B(B[0]), .Z(PRODUCT[978]) );
  AND U48 ( .A(A[977]), .B(B[0]), .Z(PRODUCT[977]) );
  AND U49 ( .A(A[976]), .B(B[0]), .Z(PRODUCT[976]) );
  AND U50 ( .A(A[975]), .B(B[0]), .Z(PRODUCT[975]) );
  AND U51 ( .A(A[974]), .B(B[0]), .Z(PRODUCT[974]) );
  AND U52 ( .A(A[973]), .B(B[0]), .Z(PRODUCT[973]) );
  AND U53 ( .A(A[972]), .B(B[0]), .Z(PRODUCT[972]) );
  AND U54 ( .A(A[971]), .B(B[0]), .Z(PRODUCT[971]) );
  AND U55 ( .A(A[970]), .B(B[0]), .Z(PRODUCT[970]) );
  AND U56 ( .A(A[969]), .B(B[0]), .Z(PRODUCT[969]) );
  AND U57 ( .A(A[968]), .B(B[0]), .Z(PRODUCT[968]) );
  AND U58 ( .A(A[967]), .B(B[0]), .Z(PRODUCT[967]) );
  AND U59 ( .A(A[966]), .B(B[0]), .Z(PRODUCT[966]) );
  AND U60 ( .A(A[965]), .B(B[0]), .Z(PRODUCT[965]) );
  AND U61 ( .A(A[964]), .B(B[0]), .Z(PRODUCT[964]) );
  AND U62 ( .A(A[963]), .B(B[0]), .Z(PRODUCT[963]) );
  AND U63 ( .A(A[962]), .B(B[0]), .Z(PRODUCT[962]) );
  AND U64 ( .A(A[961]), .B(B[0]), .Z(PRODUCT[961]) );
  AND U65 ( .A(A[960]), .B(B[0]), .Z(PRODUCT[960]) );
  AND U66 ( .A(A[959]), .B(B[0]), .Z(PRODUCT[959]) );
  AND U67 ( .A(A[958]), .B(B[0]), .Z(PRODUCT[958]) );
  AND U68 ( .A(A[957]), .B(B[0]), .Z(PRODUCT[957]) );
  AND U69 ( .A(A[956]), .B(B[0]), .Z(PRODUCT[956]) );
  AND U70 ( .A(A[955]), .B(B[0]), .Z(PRODUCT[955]) );
  AND U71 ( .A(A[954]), .B(B[0]), .Z(PRODUCT[954]) );
  AND U72 ( .A(A[953]), .B(B[0]), .Z(PRODUCT[953]) );
  AND U73 ( .A(A[952]), .B(B[0]), .Z(PRODUCT[952]) );
  AND U74 ( .A(A[951]), .B(B[0]), .Z(PRODUCT[951]) );
  AND U75 ( .A(A[950]), .B(B[0]), .Z(PRODUCT[950]) );
  AND U76 ( .A(A[949]), .B(B[0]), .Z(PRODUCT[949]) );
  AND U77 ( .A(A[948]), .B(B[0]), .Z(PRODUCT[948]) );
  AND U78 ( .A(A[947]), .B(B[0]), .Z(PRODUCT[947]) );
  AND U79 ( .A(A[946]), .B(B[0]), .Z(PRODUCT[946]) );
  AND U80 ( .A(A[945]), .B(B[0]), .Z(PRODUCT[945]) );
  AND U81 ( .A(A[944]), .B(B[0]), .Z(PRODUCT[944]) );
  AND U82 ( .A(A[943]), .B(B[0]), .Z(PRODUCT[943]) );
  AND U83 ( .A(A[942]), .B(B[0]), .Z(PRODUCT[942]) );
  AND U84 ( .A(A[941]), .B(B[0]), .Z(PRODUCT[941]) );
  AND U85 ( .A(A[940]), .B(B[0]), .Z(PRODUCT[940]) );
  AND U86 ( .A(A[939]), .B(B[0]), .Z(PRODUCT[939]) );
  AND U87 ( .A(A[938]), .B(B[0]), .Z(PRODUCT[938]) );
  AND U88 ( .A(A[937]), .B(B[0]), .Z(PRODUCT[937]) );
  AND U89 ( .A(A[936]), .B(B[0]), .Z(PRODUCT[936]) );
  AND U90 ( .A(A[935]), .B(B[0]), .Z(PRODUCT[935]) );
  AND U91 ( .A(A[934]), .B(B[0]), .Z(PRODUCT[934]) );
  AND U92 ( .A(A[933]), .B(B[0]), .Z(PRODUCT[933]) );
  AND U93 ( .A(A[932]), .B(B[0]), .Z(PRODUCT[932]) );
  AND U94 ( .A(A[931]), .B(B[0]), .Z(PRODUCT[931]) );
  AND U95 ( .A(A[930]), .B(B[0]), .Z(PRODUCT[930]) );
  AND U96 ( .A(A[929]), .B(B[0]), .Z(PRODUCT[929]) );
  AND U97 ( .A(A[928]), .B(B[0]), .Z(PRODUCT[928]) );
  AND U98 ( .A(A[927]), .B(B[0]), .Z(PRODUCT[927]) );
  AND U99 ( .A(A[926]), .B(B[0]), .Z(PRODUCT[926]) );
  AND U100 ( .A(A[925]), .B(B[0]), .Z(PRODUCT[925]) );
  AND U101 ( .A(A[924]), .B(B[0]), .Z(PRODUCT[924]) );
  AND U102 ( .A(A[923]), .B(B[0]), .Z(PRODUCT[923]) );
  AND U103 ( .A(A[922]), .B(B[0]), .Z(PRODUCT[922]) );
  AND U104 ( .A(A[921]), .B(B[0]), .Z(PRODUCT[921]) );
  AND U105 ( .A(A[920]), .B(B[0]), .Z(PRODUCT[920]) );
  AND U106 ( .A(A[919]), .B(B[0]), .Z(PRODUCT[919]) );
  AND U107 ( .A(A[918]), .B(B[0]), .Z(PRODUCT[918]) );
  AND U108 ( .A(A[917]), .B(B[0]), .Z(PRODUCT[917]) );
  AND U109 ( .A(A[916]), .B(B[0]), .Z(PRODUCT[916]) );
  AND U110 ( .A(A[915]), .B(B[0]), .Z(PRODUCT[915]) );
  AND U111 ( .A(A[914]), .B(B[0]), .Z(PRODUCT[914]) );
  AND U112 ( .A(A[913]), .B(B[0]), .Z(PRODUCT[913]) );
  AND U113 ( .A(A[912]), .B(B[0]), .Z(PRODUCT[912]) );
  AND U114 ( .A(A[911]), .B(B[0]), .Z(PRODUCT[911]) );
  AND U115 ( .A(A[910]), .B(B[0]), .Z(PRODUCT[910]) );
  AND U116 ( .A(A[909]), .B(B[0]), .Z(PRODUCT[909]) );
  AND U117 ( .A(A[908]), .B(B[0]), .Z(PRODUCT[908]) );
  AND U118 ( .A(A[907]), .B(B[0]), .Z(PRODUCT[907]) );
  AND U119 ( .A(A[906]), .B(B[0]), .Z(PRODUCT[906]) );
  AND U120 ( .A(A[905]), .B(B[0]), .Z(PRODUCT[905]) );
  AND U121 ( .A(A[904]), .B(B[0]), .Z(PRODUCT[904]) );
  AND U122 ( .A(A[903]), .B(B[0]), .Z(PRODUCT[903]) );
  AND U123 ( .A(A[902]), .B(B[0]), .Z(PRODUCT[902]) );
  AND U124 ( .A(A[901]), .B(B[0]), .Z(PRODUCT[901]) );
  AND U125 ( .A(A[900]), .B(B[0]), .Z(PRODUCT[900]) );
  AND U126 ( .A(A[899]), .B(B[0]), .Z(PRODUCT[899]) );
  AND U127 ( .A(A[898]), .B(B[0]), .Z(PRODUCT[898]) );
  AND U128 ( .A(A[897]), .B(B[0]), .Z(PRODUCT[897]) );
  AND U129 ( .A(A[896]), .B(B[0]), .Z(PRODUCT[896]) );
  AND U130 ( .A(A[895]), .B(B[0]), .Z(PRODUCT[895]) );
  AND U131 ( .A(A[894]), .B(B[0]), .Z(PRODUCT[894]) );
  AND U132 ( .A(A[893]), .B(B[0]), .Z(PRODUCT[893]) );
  AND U133 ( .A(A[892]), .B(B[0]), .Z(PRODUCT[892]) );
  AND U134 ( .A(A[891]), .B(B[0]), .Z(PRODUCT[891]) );
  AND U135 ( .A(A[890]), .B(B[0]), .Z(PRODUCT[890]) );
  AND U136 ( .A(A[889]), .B(B[0]), .Z(PRODUCT[889]) );
  AND U137 ( .A(A[888]), .B(B[0]), .Z(PRODUCT[888]) );
  AND U138 ( .A(A[887]), .B(B[0]), .Z(PRODUCT[887]) );
  AND U139 ( .A(A[886]), .B(B[0]), .Z(PRODUCT[886]) );
  AND U140 ( .A(A[885]), .B(B[0]), .Z(PRODUCT[885]) );
  AND U141 ( .A(A[884]), .B(B[0]), .Z(PRODUCT[884]) );
  AND U142 ( .A(A[883]), .B(B[0]), .Z(PRODUCT[883]) );
  AND U143 ( .A(A[882]), .B(B[0]), .Z(PRODUCT[882]) );
  AND U144 ( .A(A[881]), .B(B[0]), .Z(PRODUCT[881]) );
  AND U145 ( .A(A[880]), .B(B[0]), .Z(PRODUCT[880]) );
  AND U146 ( .A(A[879]), .B(B[0]), .Z(PRODUCT[879]) );
  AND U147 ( .A(A[878]), .B(B[0]), .Z(PRODUCT[878]) );
  AND U148 ( .A(A[877]), .B(B[0]), .Z(PRODUCT[877]) );
  AND U149 ( .A(A[876]), .B(B[0]), .Z(PRODUCT[876]) );
  AND U150 ( .A(A[875]), .B(B[0]), .Z(PRODUCT[875]) );
  AND U151 ( .A(A[874]), .B(B[0]), .Z(PRODUCT[874]) );
  AND U152 ( .A(A[873]), .B(B[0]), .Z(PRODUCT[873]) );
  AND U153 ( .A(A[872]), .B(B[0]), .Z(PRODUCT[872]) );
  AND U154 ( .A(A[871]), .B(B[0]), .Z(PRODUCT[871]) );
  AND U155 ( .A(A[870]), .B(B[0]), .Z(PRODUCT[870]) );
  AND U156 ( .A(A[869]), .B(B[0]), .Z(PRODUCT[869]) );
  AND U157 ( .A(A[868]), .B(B[0]), .Z(PRODUCT[868]) );
  AND U158 ( .A(A[867]), .B(B[0]), .Z(PRODUCT[867]) );
  AND U159 ( .A(A[866]), .B(B[0]), .Z(PRODUCT[866]) );
  AND U160 ( .A(A[865]), .B(B[0]), .Z(PRODUCT[865]) );
  AND U161 ( .A(A[864]), .B(B[0]), .Z(PRODUCT[864]) );
  AND U162 ( .A(A[863]), .B(B[0]), .Z(PRODUCT[863]) );
  AND U163 ( .A(A[862]), .B(B[0]), .Z(PRODUCT[862]) );
  AND U164 ( .A(A[861]), .B(B[0]), .Z(PRODUCT[861]) );
  AND U165 ( .A(A[860]), .B(B[0]), .Z(PRODUCT[860]) );
  AND U166 ( .A(A[859]), .B(B[0]), .Z(PRODUCT[859]) );
  AND U167 ( .A(A[858]), .B(B[0]), .Z(PRODUCT[858]) );
  AND U168 ( .A(A[857]), .B(B[0]), .Z(PRODUCT[857]) );
  AND U169 ( .A(A[856]), .B(B[0]), .Z(PRODUCT[856]) );
  AND U170 ( .A(A[855]), .B(B[0]), .Z(PRODUCT[855]) );
  AND U171 ( .A(A[854]), .B(B[0]), .Z(PRODUCT[854]) );
  AND U172 ( .A(A[853]), .B(B[0]), .Z(PRODUCT[853]) );
  AND U173 ( .A(A[852]), .B(B[0]), .Z(PRODUCT[852]) );
  AND U174 ( .A(A[851]), .B(B[0]), .Z(PRODUCT[851]) );
  AND U175 ( .A(A[850]), .B(B[0]), .Z(PRODUCT[850]) );
  AND U176 ( .A(A[849]), .B(B[0]), .Z(PRODUCT[849]) );
  AND U177 ( .A(A[848]), .B(B[0]), .Z(PRODUCT[848]) );
  AND U178 ( .A(A[847]), .B(B[0]), .Z(PRODUCT[847]) );
  AND U179 ( .A(A[846]), .B(B[0]), .Z(PRODUCT[846]) );
  AND U180 ( .A(A[845]), .B(B[0]), .Z(PRODUCT[845]) );
  AND U181 ( .A(A[844]), .B(B[0]), .Z(PRODUCT[844]) );
  AND U182 ( .A(A[843]), .B(B[0]), .Z(PRODUCT[843]) );
  AND U183 ( .A(A[842]), .B(B[0]), .Z(PRODUCT[842]) );
  AND U184 ( .A(A[841]), .B(B[0]), .Z(PRODUCT[841]) );
  AND U185 ( .A(A[840]), .B(B[0]), .Z(PRODUCT[840]) );
  AND U186 ( .A(A[839]), .B(B[0]), .Z(PRODUCT[839]) );
  AND U187 ( .A(A[838]), .B(B[0]), .Z(PRODUCT[838]) );
  AND U188 ( .A(A[837]), .B(B[0]), .Z(PRODUCT[837]) );
  AND U189 ( .A(A[836]), .B(B[0]), .Z(PRODUCT[836]) );
  AND U190 ( .A(A[835]), .B(B[0]), .Z(PRODUCT[835]) );
  AND U191 ( .A(A[834]), .B(B[0]), .Z(PRODUCT[834]) );
  AND U192 ( .A(A[833]), .B(B[0]), .Z(PRODUCT[833]) );
  AND U193 ( .A(A[832]), .B(B[0]), .Z(PRODUCT[832]) );
  AND U194 ( .A(A[831]), .B(B[0]), .Z(PRODUCT[831]) );
  AND U195 ( .A(A[830]), .B(B[0]), .Z(PRODUCT[830]) );
  AND U196 ( .A(A[829]), .B(B[0]), .Z(PRODUCT[829]) );
  AND U197 ( .A(A[828]), .B(B[0]), .Z(PRODUCT[828]) );
  AND U198 ( .A(A[827]), .B(B[0]), .Z(PRODUCT[827]) );
  AND U199 ( .A(A[826]), .B(B[0]), .Z(PRODUCT[826]) );
  AND U200 ( .A(A[825]), .B(B[0]), .Z(PRODUCT[825]) );
  AND U201 ( .A(A[824]), .B(B[0]), .Z(PRODUCT[824]) );
  AND U202 ( .A(A[823]), .B(B[0]), .Z(PRODUCT[823]) );
  AND U203 ( .A(A[822]), .B(B[0]), .Z(PRODUCT[822]) );
  AND U204 ( .A(A[821]), .B(B[0]), .Z(PRODUCT[821]) );
  AND U205 ( .A(A[820]), .B(B[0]), .Z(PRODUCT[820]) );
  AND U206 ( .A(A[819]), .B(B[0]), .Z(PRODUCT[819]) );
  AND U207 ( .A(A[818]), .B(B[0]), .Z(PRODUCT[818]) );
  AND U208 ( .A(A[817]), .B(B[0]), .Z(PRODUCT[817]) );
  AND U209 ( .A(A[816]), .B(B[0]), .Z(PRODUCT[816]) );
  AND U210 ( .A(A[815]), .B(B[0]), .Z(PRODUCT[815]) );
  AND U211 ( .A(A[814]), .B(B[0]), .Z(PRODUCT[814]) );
  AND U212 ( .A(A[813]), .B(B[0]), .Z(PRODUCT[813]) );
  AND U213 ( .A(A[812]), .B(B[0]), .Z(PRODUCT[812]) );
  AND U214 ( .A(A[811]), .B(B[0]), .Z(PRODUCT[811]) );
  AND U215 ( .A(A[810]), .B(B[0]), .Z(PRODUCT[810]) );
  AND U216 ( .A(A[809]), .B(B[0]), .Z(PRODUCT[809]) );
  AND U217 ( .A(A[808]), .B(B[0]), .Z(PRODUCT[808]) );
  AND U218 ( .A(A[807]), .B(B[0]), .Z(PRODUCT[807]) );
  AND U219 ( .A(A[806]), .B(B[0]), .Z(PRODUCT[806]) );
  AND U220 ( .A(A[805]), .B(B[0]), .Z(PRODUCT[805]) );
  AND U221 ( .A(A[804]), .B(B[0]), .Z(PRODUCT[804]) );
  AND U222 ( .A(A[803]), .B(B[0]), .Z(PRODUCT[803]) );
  AND U223 ( .A(A[802]), .B(B[0]), .Z(PRODUCT[802]) );
  AND U224 ( .A(A[801]), .B(B[0]), .Z(PRODUCT[801]) );
  AND U225 ( .A(A[800]), .B(B[0]), .Z(PRODUCT[800]) );
  AND U226 ( .A(A[799]), .B(B[0]), .Z(PRODUCT[799]) );
  AND U227 ( .A(A[798]), .B(B[0]), .Z(PRODUCT[798]) );
  AND U228 ( .A(A[797]), .B(B[0]), .Z(PRODUCT[797]) );
  AND U229 ( .A(A[796]), .B(B[0]), .Z(PRODUCT[796]) );
  AND U230 ( .A(A[795]), .B(B[0]), .Z(PRODUCT[795]) );
  AND U231 ( .A(A[794]), .B(B[0]), .Z(PRODUCT[794]) );
  AND U232 ( .A(A[793]), .B(B[0]), .Z(PRODUCT[793]) );
  AND U233 ( .A(A[792]), .B(B[0]), .Z(PRODUCT[792]) );
  AND U234 ( .A(A[791]), .B(B[0]), .Z(PRODUCT[791]) );
  AND U235 ( .A(A[790]), .B(B[0]), .Z(PRODUCT[790]) );
  AND U236 ( .A(A[789]), .B(B[0]), .Z(PRODUCT[789]) );
  AND U237 ( .A(A[788]), .B(B[0]), .Z(PRODUCT[788]) );
  AND U238 ( .A(A[787]), .B(B[0]), .Z(PRODUCT[787]) );
  AND U239 ( .A(A[786]), .B(B[0]), .Z(PRODUCT[786]) );
  AND U240 ( .A(A[785]), .B(B[0]), .Z(PRODUCT[785]) );
  AND U241 ( .A(A[784]), .B(B[0]), .Z(PRODUCT[784]) );
  AND U242 ( .A(A[783]), .B(B[0]), .Z(PRODUCT[783]) );
  AND U243 ( .A(A[782]), .B(B[0]), .Z(PRODUCT[782]) );
  AND U244 ( .A(A[781]), .B(B[0]), .Z(PRODUCT[781]) );
  AND U245 ( .A(A[780]), .B(B[0]), .Z(PRODUCT[780]) );
  AND U246 ( .A(A[779]), .B(B[0]), .Z(PRODUCT[779]) );
  AND U247 ( .A(A[778]), .B(B[0]), .Z(PRODUCT[778]) );
  AND U248 ( .A(A[777]), .B(B[0]), .Z(PRODUCT[777]) );
  AND U249 ( .A(A[776]), .B(B[0]), .Z(PRODUCT[776]) );
  AND U250 ( .A(A[775]), .B(B[0]), .Z(PRODUCT[775]) );
  AND U251 ( .A(A[774]), .B(B[0]), .Z(PRODUCT[774]) );
  AND U252 ( .A(A[773]), .B(B[0]), .Z(PRODUCT[773]) );
  AND U253 ( .A(A[772]), .B(B[0]), .Z(PRODUCT[772]) );
  AND U254 ( .A(A[771]), .B(B[0]), .Z(PRODUCT[771]) );
  AND U255 ( .A(A[770]), .B(B[0]), .Z(PRODUCT[770]) );
  AND U256 ( .A(A[769]), .B(B[0]), .Z(PRODUCT[769]) );
  AND U257 ( .A(A[768]), .B(B[0]), .Z(PRODUCT[768]) );
  AND U258 ( .A(A[767]), .B(B[0]), .Z(PRODUCT[767]) );
  AND U259 ( .A(A[766]), .B(B[0]), .Z(PRODUCT[766]) );
  AND U260 ( .A(A[765]), .B(B[0]), .Z(PRODUCT[765]) );
  AND U261 ( .A(A[764]), .B(B[0]), .Z(PRODUCT[764]) );
  AND U262 ( .A(A[763]), .B(B[0]), .Z(PRODUCT[763]) );
  AND U263 ( .A(A[762]), .B(B[0]), .Z(PRODUCT[762]) );
  AND U264 ( .A(A[761]), .B(B[0]), .Z(PRODUCT[761]) );
  AND U265 ( .A(A[760]), .B(B[0]), .Z(PRODUCT[760]) );
  AND U266 ( .A(A[759]), .B(B[0]), .Z(PRODUCT[759]) );
  AND U267 ( .A(A[758]), .B(B[0]), .Z(PRODUCT[758]) );
  AND U268 ( .A(A[757]), .B(B[0]), .Z(PRODUCT[757]) );
  AND U269 ( .A(A[756]), .B(B[0]), .Z(PRODUCT[756]) );
  AND U270 ( .A(A[755]), .B(B[0]), .Z(PRODUCT[755]) );
  AND U271 ( .A(A[754]), .B(B[0]), .Z(PRODUCT[754]) );
  AND U272 ( .A(A[753]), .B(B[0]), .Z(PRODUCT[753]) );
  AND U273 ( .A(A[752]), .B(B[0]), .Z(PRODUCT[752]) );
  AND U274 ( .A(A[751]), .B(B[0]), .Z(PRODUCT[751]) );
  AND U275 ( .A(A[750]), .B(B[0]), .Z(PRODUCT[750]) );
  AND U276 ( .A(A[749]), .B(B[0]), .Z(PRODUCT[749]) );
  AND U277 ( .A(A[748]), .B(B[0]), .Z(PRODUCT[748]) );
  AND U278 ( .A(A[747]), .B(B[0]), .Z(PRODUCT[747]) );
  AND U279 ( .A(A[746]), .B(B[0]), .Z(PRODUCT[746]) );
  AND U280 ( .A(A[745]), .B(B[0]), .Z(PRODUCT[745]) );
  AND U281 ( .A(A[744]), .B(B[0]), .Z(PRODUCT[744]) );
  AND U282 ( .A(A[743]), .B(B[0]), .Z(PRODUCT[743]) );
  AND U283 ( .A(A[742]), .B(B[0]), .Z(PRODUCT[742]) );
  AND U284 ( .A(A[741]), .B(B[0]), .Z(PRODUCT[741]) );
  AND U285 ( .A(A[740]), .B(B[0]), .Z(PRODUCT[740]) );
  AND U286 ( .A(A[739]), .B(B[0]), .Z(PRODUCT[739]) );
  AND U287 ( .A(A[738]), .B(B[0]), .Z(PRODUCT[738]) );
  AND U288 ( .A(A[737]), .B(B[0]), .Z(PRODUCT[737]) );
  AND U289 ( .A(A[736]), .B(B[0]), .Z(PRODUCT[736]) );
  AND U290 ( .A(A[735]), .B(B[0]), .Z(PRODUCT[735]) );
  AND U291 ( .A(A[734]), .B(B[0]), .Z(PRODUCT[734]) );
  AND U292 ( .A(A[733]), .B(B[0]), .Z(PRODUCT[733]) );
  AND U293 ( .A(A[732]), .B(B[0]), .Z(PRODUCT[732]) );
  AND U294 ( .A(A[731]), .B(B[0]), .Z(PRODUCT[731]) );
  AND U295 ( .A(A[730]), .B(B[0]), .Z(PRODUCT[730]) );
  AND U296 ( .A(A[729]), .B(B[0]), .Z(PRODUCT[729]) );
  AND U297 ( .A(A[728]), .B(B[0]), .Z(PRODUCT[728]) );
  AND U298 ( .A(A[727]), .B(B[0]), .Z(PRODUCT[727]) );
  AND U299 ( .A(A[726]), .B(B[0]), .Z(PRODUCT[726]) );
  AND U300 ( .A(A[725]), .B(B[0]), .Z(PRODUCT[725]) );
  AND U301 ( .A(A[724]), .B(B[0]), .Z(PRODUCT[724]) );
  AND U302 ( .A(A[723]), .B(B[0]), .Z(PRODUCT[723]) );
  AND U303 ( .A(A[722]), .B(B[0]), .Z(PRODUCT[722]) );
  AND U304 ( .A(A[721]), .B(B[0]), .Z(PRODUCT[721]) );
  AND U305 ( .A(A[720]), .B(B[0]), .Z(PRODUCT[720]) );
  AND U306 ( .A(A[719]), .B(B[0]), .Z(PRODUCT[719]) );
  AND U307 ( .A(A[718]), .B(B[0]), .Z(PRODUCT[718]) );
  AND U308 ( .A(A[717]), .B(B[0]), .Z(PRODUCT[717]) );
  AND U309 ( .A(A[716]), .B(B[0]), .Z(PRODUCT[716]) );
  AND U310 ( .A(A[715]), .B(B[0]), .Z(PRODUCT[715]) );
  AND U311 ( .A(A[714]), .B(B[0]), .Z(PRODUCT[714]) );
  AND U312 ( .A(A[713]), .B(B[0]), .Z(PRODUCT[713]) );
  AND U313 ( .A(A[712]), .B(B[0]), .Z(PRODUCT[712]) );
  AND U314 ( .A(A[711]), .B(B[0]), .Z(PRODUCT[711]) );
  AND U315 ( .A(A[710]), .B(B[0]), .Z(PRODUCT[710]) );
  AND U316 ( .A(A[709]), .B(B[0]), .Z(PRODUCT[709]) );
  AND U317 ( .A(A[708]), .B(B[0]), .Z(PRODUCT[708]) );
  AND U318 ( .A(A[707]), .B(B[0]), .Z(PRODUCT[707]) );
  AND U319 ( .A(A[706]), .B(B[0]), .Z(PRODUCT[706]) );
  AND U320 ( .A(A[705]), .B(B[0]), .Z(PRODUCT[705]) );
  AND U321 ( .A(A[704]), .B(B[0]), .Z(PRODUCT[704]) );
  AND U322 ( .A(A[703]), .B(B[0]), .Z(PRODUCT[703]) );
  AND U323 ( .A(A[702]), .B(B[0]), .Z(PRODUCT[702]) );
  AND U324 ( .A(A[701]), .B(B[0]), .Z(PRODUCT[701]) );
  AND U325 ( .A(A[700]), .B(B[0]), .Z(PRODUCT[700]) );
  AND U326 ( .A(A[699]), .B(B[0]), .Z(PRODUCT[699]) );
  AND U327 ( .A(A[698]), .B(B[0]), .Z(PRODUCT[698]) );
  AND U328 ( .A(A[697]), .B(B[0]), .Z(PRODUCT[697]) );
  AND U329 ( .A(A[696]), .B(B[0]), .Z(PRODUCT[696]) );
  AND U330 ( .A(A[695]), .B(B[0]), .Z(PRODUCT[695]) );
  AND U331 ( .A(A[694]), .B(B[0]), .Z(PRODUCT[694]) );
  AND U332 ( .A(A[693]), .B(B[0]), .Z(PRODUCT[693]) );
  AND U333 ( .A(A[692]), .B(B[0]), .Z(PRODUCT[692]) );
  AND U334 ( .A(A[691]), .B(B[0]), .Z(PRODUCT[691]) );
  AND U335 ( .A(A[690]), .B(B[0]), .Z(PRODUCT[690]) );
  AND U336 ( .A(A[689]), .B(B[0]), .Z(PRODUCT[689]) );
  AND U337 ( .A(A[688]), .B(B[0]), .Z(PRODUCT[688]) );
  AND U338 ( .A(A[687]), .B(B[0]), .Z(PRODUCT[687]) );
  AND U339 ( .A(A[686]), .B(B[0]), .Z(PRODUCT[686]) );
  AND U340 ( .A(A[685]), .B(B[0]), .Z(PRODUCT[685]) );
  AND U341 ( .A(A[684]), .B(B[0]), .Z(PRODUCT[684]) );
  AND U342 ( .A(A[683]), .B(B[0]), .Z(PRODUCT[683]) );
  AND U343 ( .A(A[682]), .B(B[0]), .Z(PRODUCT[682]) );
  AND U344 ( .A(A[681]), .B(B[0]), .Z(PRODUCT[681]) );
  AND U345 ( .A(A[680]), .B(B[0]), .Z(PRODUCT[680]) );
  AND U346 ( .A(A[679]), .B(B[0]), .Z(PRODUCT[679]) );
  AND U347 ( .A(A[678]), .B(B[0]), .Z(PRODUCT[678]) );
  AND U348 ( .A(A[677]), .B(B[0]), .Z(PRODUCT[677]) );
  AND U349 ( .A(A[676]), .B(B[0]), .Z(PRODUCT[676]) );
  AND U350 ( .A(A[675]), .B(B[0]), .Z(PRODUCT[675]) );
  AND U351 ( .A(A[674]), .B(B[0]), .Z(PRODUCT[674]) );
  AND U352 ( .A(A[673]), .B(B[0]), .Z(PRODUCT[673]) );
  AND U353 ( .A(A[672]), .B(B[0]), .Z(PRODUCT[672]) );
  AND U354 ( .A(A[671]), .B(B[0]), .Z(PRODUCT[671]) );
  AND U355 ( .A(A[670]), .B(B[0]), .Z(PRODUCT[670]) );
  AND U356 ( .A(A[669]), .B(B[0]), .Z(PRODUCT[669]) );
  AND U357 ( .A(A[668]), .B(B[0]), .Z(PRODUCT[668]) );
  AND U358 ( .A(A[667]), .B(B[0]), .Z(PRODUCT[667]) );
  AND U359 ( .A(A[666]), .B(B[0]), .Z(PRODUCT[666]) );
  AND U360 ( .A(A[665]), .B(B[0]), .Z(PRODUCT[665]) );
  AND U361 ( .A(A[664]), .B(B[0]), .Z(PRODUCT[664]) );
  AND U362 ( .A(A[663]), .B(B[0]), .Z(PRODUCT[663]) );
  AND U363 ( .A(A[662]), .B(B[0]), .Z(PRODUCT[662]) );
  AND U364 ( .A(A[661]), .B(B[0]), .Z(PRODUCT[661]) );
  AND U365 ( .A(A[660]), .B(B[0]), .Z(PRODUCT[660]) );
  AND U366 ( .A(A[659]), .B(B[0]), .Z(PRODUCT[659]) );
  AND U367 ( .A(A[658]), .B(B[0]), .Z(PRODUCT[658]) );
  AND U368 ( .A(A[657]), .B(B[0]), .Z(PRODUCT[657]) );
  AND U369 ( .A(A[656]), .B(B[0]), .Z(PRODUCT[656]) );
  AND U370 ( .A(A[655]), .B(B[0]), .Z(PRODUCT[655]) );
  AND U371 ( .A(A[654]), .B(B[0]), .Z(PRODUCT[654]) );
  AND U372 ( .A(A[653]), .B(B[0]), .Z(PRODUCT[653]) );
  AND U373 ( .A(A[652]), .B(B[0]), .Z(PRODUCT[652]) );
  AND U374 ( .A(A[651]), .B(B[0]), .Z(PRODUCT[651]) );
  AND U375 ( .A(A[650]), .B(B[0]), .Z(PRODUCT[650]) );
  AND U376 ( .A(A[649]), .B(B[0]), .Z(PRODUCT[649]) );
  AND U377 ( .A(A[648]), .B(B[0]), .Z(PRODUCT[648]) );
  AND U378 ( .A(A[647]), .B(B[0]), .Z(PRODUCT[647]) );
  AND U379 ( .A(A[646]), .B(B[0]), .Z(PRODUCT[646]) );
  AND U380 ( .A(A[645]), .B(B[0]), .Z(PRODUCT[645]) );
  AND U381 ( .A(A[644]), .B(B[0]), .Z(PRODUCT[644]) );
  AND U382 ( .A(A[643]), .B(B[0]), .Z(PRODUCT[643]) );
  AND U383 ( .A(A[642]), .B(B[0]), .Z(PRODUCT[642]) );
  AND U384 ( .A(A[641]), .B(B[0]), .Z(PRODUCT[641]) );
  AND U385 ( .A(A[640]), .B(B[0]), .Z(PRODUCT[640]) );
  AND U386 ( .A(A[639]), .B(B[0]), .Z(PRODUCT[639]) );
  AND U387 ( .A(A[638]), .B(B[0]), .Z(PRODUCT[638]) );
  AND U388 ( .A(A[637]), .B(B[0]), .Z(PRODUCT[637]) );
  AND U389 ( .A(A[636]), .B(B[0]), .Z(PRODUCT[636]) );
  AND U390 ( .A(A[635]), .B(B[0]), .Z(PRODUCT[635]) );
  AND U391 ( .A(A[634]), .B(B[0]), .Z(PRODUCT[634]) );
  AND U392 ( .A(A[633]), .B(B[0]), .Z(PRODUCT[633]) );
  AND U393 ( .A(A[632]), .B(B[0]), .Z(PRODUCT[632]) );
  AND U394 ( .A(A[631]), .B(B[0]), .Z(PRODUCT[631]) );
  AND U395 ( .A(A[630]), .B(B[0]), .Z(PRODUCT[630]) );
  AND U396 ( .A(A[629]), .B(B[0]), .Z(PRODUCT[629]) );
  AND U397 ( .A(A[628]), .B(B[0]), .Z(PRODUCT[628]) );
  AND U398 ( .A(A[627]), .B(B[0]), .Z(PRODUCT[627]) );
  AND U399 ( .A(A[626]), .B(B[0]), .Z(PRODUCT[626]) );
  AND U400 ( .A(A[625]), .B(B[0]), .Z(PRODUCT[625]) );
  AND U401 ( .A(A[624]), .B(B[0]), .Z(PRODUCT[624]) );
  AND U402 ( .A(A[623]), .B(B[0]), .Z(PRODUCT[623]) );
  AND U403 ( .A(A[622]), .B(B[0]), .Z(PRODUCT[622]) );
  AND U404 ( .A(A[621]), .B(B[0]), .Z(PRODUCT[621]) );
  AND U405 ( .A(A[620]), .B(B[0]), .Z(PRODUCT[620]) );
  AND U406 ( .A(A[619]), .B(B[0]), .Z(PRODUCT[619]) );
  AND U407 ( .A(A[618]), .B(B[0]), .Z(PRODUCT[618]) );
  AND U408 ( .A(A[617]), .B(B[0]), .Z(PRODUCT[617]) );
  AND U409 ( .A(A[616]), .B(B[0]), .Z(PRODUCT[616]) );
  AND U410 ( .A(A[615]), .B(B[0]), .Z(PRODUCT[615]) );
  AND U411 ( .A(A[614]), .B(B[0]), .Z(PRODUCT[614]) );
  AND U412 ( .A(A[613]), .B(B[0]), .Z(PRODUCT[613]) );
  AND U413 ( .A(A[612]), .B(B[0]), .Z(PRODUCT[612]) );
  AND U414 ( .A(A[611]), .B(B[0]), .Z(PRODUCT[611]) );
  AND U415 ( .A(A[610]), .B(B[0]), .Z(PRODUCT[610]) );
  AND U416 ( .A(A[609]), .B(B[0]), .Z(PRODUCT[609]) );
  AND U417 ( .A(A[608]), .B(B[0]), .Z(PRODUCT[608]) );
  AND U418 ( .A(A[607]), .B(B[0]), .Z(PRODUCT[607]) );
  AND U419 ( .A(A[606]), .B(B[0]), .Z(PRODUCT[606]) );
  AND U420 ( .A(A[605]), .B(B[0]), .Z(PRODUCT[605]) );
  AND U421 ( .A(A[604]), .B(B[0]), .Z(PRODUCT[604]) );
  AND U422 ( .A(A[603]), .B(B[0]), .Z(PRODUCT[603]) );
  AND U423 ( .A(A[602]), .B(B[0]), .Z(PRODUCT[602]) );
  AND U424 ( .A(A[601]), .B(B[0]), .Z(PRODUCT[601]) );
  AND U425 ( .A(A[600]), .B(B[0]), .Z(PRODUCT[600]) );
  AND U426 ( .A(A[599]), .B(B[0]), .Z(PRODUCT[599]) );
  AND U427 ( .A(A[598]), .B(B[0]), .Z(PRODUCT[598]) );
  AND U428 ( .A(A[597]), .B(B[0]), .Z(PRODUCT[597]) );
  AND U429 ( .A(A[596]), .B(B[0]), .Z(PRODUCT[596]) );
  AND U430 ( .A(A[595]), .B(B[0]), .Z(PRODUCT[595]) );
  AND U431 ( .A(A[594]), .B(B[0]), .Z(PRODUCT[594]) );
  AND U432 ( .A(A[593]), .B(B[0]), .Z(PRODUCT[593]) );
  AND U433 ( .A(A[592]), .B(B[0]), .Z(PRODUCT[592]) );
  AND U434 ( .A(A[591]), .B(B[0]), .Z(PRODUCT[591]) );
  AND U435 ( .A(A[590]), .B(B[0]), .Z(PRODUCT[590]) );
  AND U436 ( .A(A[589]), .B(B[0]), .Z(PRODUCT[589]) );
  AND U437 ( .A(A[588]), .B(B[0]), .Z(PRODUCT[588]) );
  AND U438 ( .A(A[587]), .B(B[0]), .Z(PRODUCT[587]) );
  AND U439 ( .A(A[586]), .B(B[0]), .Z(PRODUCT[586]) );
  AND U440 ( .A(A[585]), .B(B[0]), .Z(PRODUCT[585]) );
  AND U441 ( .A(A[584]), .B(B[0]), .Z(PRODUCT[584]) );
  AND U442 ( .A(A[583]), .B(B[0]), .Z(PRODUCT[583]) );
  AND U443 ( .A(A[582]), .B(B[0]), .Z(PRODUCT[582]) );
  AND U444 ( .A(A[581]), .B(B[0]), .Z(PRODUCT[581]) );
  AND U445 ( .A(A[580]), .B(B[0]), .Z(PRODUCT[580]) );
  AND U446 ( .A(A[579]), .B(B[0]), .Z(PRODUCT[579]) );
  AND U447 ( .A(A[578]), .B(B[0]), .Z(PRODUCT[578]) );
  AND U448 ( .A(A[577]), .B(B[0]), .Z(PRODUCT[577]) );
  AND U449 ( .A(A[576]), .B(B[0]), .Z(PRODUCT[576]) );
  AND U450 ( .A(A[575]), .B(B[0]), .Z(PRODUCT[575]) );
  AND U451 ( .A(A[574]), .B(B[0]), .Z(PRODUCT[574]) );
  AND U452 ( .A(A[573]), .B(B[0]), .Z(PRODUCT[573]) );
  AND U453 ( .A(A[572]), .B(B[0]), .Z(PRODUCT[572]) );
  AND U454 ( .A(A[571]), .B(B[0]), .Z(PRODUCT[571]) );
  AND U455 ( .A(A[570]), .B(B[0]), .Z(PRODUCT[570]) );
  AND U456 ( .A(A[569]), .B(B[0]), .Z(PRODUCT[569]) );
  AND U457 ( .A(A[568]), .B(B[0]), .Z(PRODUCT[568]) );
  AND U458 ( .A(A[567]), .B(B[0]), .Z(PRODUCT[567]) );
  AND U459 ( .A(A[566]), .B(B[0]), .Z(PRODUCT[566]) );
  AND U460 ( .A(A[565]), .B(B[0]), .Z(PRODUCT[565]) );
  AND U461 ( .A(A[564]), .B(B[0]), .Z(PRODUCT[564]) );
  AND U462 ( .A(A[563]), .B(B[0]), .Z(PRODUCT[563]) );
  AND U463 ( .A(A[562]), .B(B[0]), .Z(PRODUCT[562]) );
  AND U464 ( .A(A[561]), .B(B[0]), .Z(PRODUCT[561]) );
  AND U465 ( .A(A[560]), .B(B[0]), .Z(PRODUCT[560]) );
  AND U466 ( .A(A[559]), .B(B[0]), .Z(PRODUCT[559]) );
  AND U467 ( .A(A[558]), .B(B[0]), .Z(PRODUCT[558]) );
  AND U468 ( .A(A[557]), .B(B[0]), .Z(PRODUCT[557]) );
  AND U469 ( .A(A[556]), .B(B[0]), .Z(PRODUCT[556]) );
  AND U470 ( .A(A[555]), .B(B[0]), .Z(PRODUCT[555]) );
  AND U471 ( .A(A[554]), .B(B[0]), .Z(PRODUCT[554]) );
  AND U472 ( .A(A[553]), .B(B[0]), .Z(PRODUCT[553]) );
  AND U473 ( .A(A[552]), .B(B[0]), .Z(PRODUCT[552]) );
  AND U474 ( .A(A[551]), .B(B[0]), .Z(PRODUCT[551]) );
  AND U475 ( .A(A[550]), .B(B[0]), .Z(PRODUCT[550]) );
  AND U476 ( .A(A[549]), .B(B[0]), .Z(PRODUCT[549]) );
  AND U477 ( .A(A[548]), .B(B[0]), .Z(PRODUCT[548]) );
  AND U478 ( .A(A[547]), .B(B[0]), .Z(PRODUCT[547]) );
  AND U479 ( .A(A[546]), .B(B[0]), .Z(PRODUCT[546]) );
  AND U480 ( .A(A[545]), .B(B[0]), .Z(PRODUCT[545]) );
  AND U481 ( .A(A[544]), .B(B[0]), .Z(PRODUCT[544]) );
  AND U482 ( .A(A[543]), .B(B[0]), .Z(PRODUCT[543]) );
  AND U483 ( .A(A[542]), .B(B[0]), .Z(PRODUCT[542]) );
  AND U484 ( .A(A[541]), .B(B[0]), .Z(PRODUCT[541]) );
  AND U485 ( .A(A[540]), .B(B[0]), .Z(PRODUCT[540]) );
  AND U486 ( .A(A[539]), .B(B[0]), .Z(PRODUCT[539]) );
  AND U487 ( .A(A[538]), .B(B[0]), .Z(PRODUCT[538]) );
  AND U488 ( .A(A[537]), .B(B[0]), .Z(PRODUCT[537]) );
  AND U489 ( .A(A[536]), .B(B[0]), .Z(PRODUCT[536]) );
  AND U490 ( .A(A[535]), .B(B[0]), .Z(PRODUCT[535]) );
  AND U491 ( .A(A[534]), .B(B[0]), .Z(PRODUCT[534]) );
  AND U492 ( .A(A[533]), .B(B[0]), .Z(PRODUCT[533]) );
  AND U493 ( .A(A[532]), .B(B[0]), .Z(PRODUCT[532]) );
  AND U494 ( .A(A[531]), .B(B[0]), .Z(PRODUCT[531]) );
  AND U495 ( .A(A[530]), .B(B[0]), .Z(PRODUCT[530]) );
  AND U496 ( .A(A[529]), .B(B[0]), .Z(PRODUCT[529]) );
  AND U497 ( .A(A[528]), .B(B[0]), .Z(PRODUCT[528]) );
  AND U498 ( .A(A[527]), .B(B[0]), .Z(PRODUCT[527]) );
  AND U499 ( .A(A[526]), .B(B[0]), .Z(PRODUCT[526]) );
  AND U500 ( .A(A[525]), .B(B[0]), .Z(PRODUCT[525]) );
  AND U501 ( .A(A[524]), .B(B[0]), .Z(PRODUCT[524]) );
  AND U502 ( .A(A[523]), .B(B[0]), .Z(PRODUCT[523]) );
  AND U503 ( .A(A[522]), .B(B[0]), .Z(PRODUCT[522]) );
  AND U504 ( .A(A[521]), .B(B[0]), .Z(PRODUCT[521]) );
  AND U505 ( .A(A[520]), .B(B[0]), .Z(PRODUCT[520]) );
  AND U506 ( .A(A[519]), .B(B[0]), .Z(PRODUCT[519]) );
  AND U507 ( .A(A[518]), .B(B[0]), .Z(PRODUCT[518]) );
  AND U508 ( .A(A[517]), .B(B[0]), .Z(PRODUCT[517]) );
  AND U509 ( .A(A[516]), .B(B[0]), .Z(PRODUCT[516]) );
  AND U510 ( .A(A[515]), .B(B[0]), .Z(PRODUCT[515]) );
  AND U511 ( .A(A[514]), .B(B[0]), .Z(PRODUCT[514]) );
  AND U512 ( .A(A[513]), .B(B[0]), .Z(PRODUCT[513]) );
  AND U513 ( .A(A[512]), .B(B[0]), .Z(PRODUCT[512]) );
  AND U514 ( .A(A[511]), .B(B[0]), .Z(PRODUCT[511]) );
  AND U515 ( .A(A[510]), .B(B[0]), .Z(PRODUCT[510]) );
  AND U516 ( .A(A[509]), .B(B[0]), .Z(PRODUCT[509]) );
  AND U517 ( .A(A[508]), .B(B[0]), .Z(PRODUCT[508]) );
  AND U518 ( .A(A[507]), .B(B[0]), .Z(PRODUCT[507]) );
  AND U519 ( .A(A[506]), .B(B[0]), .Z(PRODUCT[506]) );
  AND U520 ( .A(A[505]), .B(B[0]), .Z(PRODUCT[505]) );
  AND U521 ( .A(A[504]), .B(B[0]), .Z(PRODUCT[504]) );
  AND U522 ( .A(A[503]), .B(B[0]), .Z(PRODUCT[503]) );
  AND U523 ( .A(A[502]), .B(B[0]), .Z(PRODUCT[502]) );
  AND U524 ( .A(A[501]), .B(B[0]), .Z(PRODUCT[501]) );
  AND U525 ( .A(A[500]), .B(B[0]), .Z(PRODUCT[500]) );
  AND U526 ( .A(A[499]), .B(B[0]), .Z(PRODUCT[499]) );
  AND U527 ( .A(A[498]), .B(B[0]), .Z(PRODUCT[498]) );
  AND U528 ( .A(A[497]), .B(B[0]), .Z(PRODUCT[497]) );
  AND U529 ( .A(A[496]), .B(B[0]), .Z(PRODUCT[496]) );
  AND U530 ( .A(A[495]), .B(B[0]), .Z(PRODUCT[495]) );
  AND U531 ( .A(A[494]), .B(B[0]), .Z(PRODUCT[494]) );
  AND U532 ( .A(A[493]), .B(B[0]), .Z(PRODUCT[493]) );
  AND U533 ( .A(A[492]), .B(B[0]), .Z(PRODUCT[492]) );
  AND U534 ( .A(A[491]), .B(B[0]), .Z(PRODUCT[491]) );
  AND U535 ( .A(A[490]), .B(B[0]), .Z(PRODUCT[490]) );
  AND U536 ( .A(A[489]), .B(B[0]), .Z(PRODUCT[489]) );
  AND U537 ( .A(A[488]), .B(B[0]), .Z(PRODUCT[488]) );
  AND U538 ( .A(A[487]), .B(B[0]), .Z(PRODUCT[487]) );
  AND U539 ( .A(A[486]), .B(B[0]), .Z(PRODUCT[486]) );
  AND U540 ( .A(A[485]), .B(B[0]), .Z(PRODUCT[485]) );
  AND U541 ( .A(A[484]), .B(B[0]), .Z(PRODUCT[484]) );
  AND U542 ( .A(A[483]), .B(B[0]), .Z(PRODUCT[483]) );
  AND U543 ( .A(A[482]), .B(B[0]), .Z(PRODUCT[482]) );
  AND U544 ( .A(A[481]), .B(B[0]), .Z(PRODUCT[481]) );
  AND U545 ( .A(A[480]), .B(B[0]), .Z(PRODUCT[480]) );
  AND U546 ( .A(A[479]), .B(B[0]), .Z(PRODUCT[479]) );
  AND U547 ( .A(A[478]), .B(B[0]), .Z(PRODUCT[478]) );
  AND U548 ( .A(A[477]), .B(B[0]), .Z(PRODUCT[477]) );
  AND U549 ( .A(A[476]), .B(B[0]), .Z(PRODUCT[476]) );
  AND U550 ( .A(A[475]), .B(B[0]), .Z(PRODUCT[475]) );
  AND U551 ( .A(A[474]), .B(B[0]), .Z(PRODUCT[474]) );
  AND U552 ( .A(A[473]), .B(B[0]), .Z(PRODUCT[473]) );
  AND U553 ( .A(A[472]), .B(B[0]), .Z(PRODUCT[472]) );
  AND U554 ( .A(A[471]), .B(B[0]), .Z(PRODUCT[471]) );
  AND U555 ( .A(A[470]), .B(B[0]), .Z(PRODUCT[470]) );
  AND U556 ( .A(A[469]), .B(B[0]), .Z(PRODUCT[469]) );
  AND U557 ( .A(A[468]), .B(B[0]), .Z(PRODUCT[468]) );
  AND U558 ( .A(A[467]), .B(B[0]), .Z(PRODUCT[467]) );
  AND U559 ( .A(A[466]), .B(B[0]), .Z(PRODUCT[466]) );
  AND U560 ( .A(A[465]), .B(B[0]), .Z(PRODUCT[465]) );
  AND U561 ( .A(A[464]), .B(B[0]), .Z(PRODUCT[464]) );
  AND U562 ( .A(A[463]), .B(B[0]), .Z(PRODUCT[463]) );
  AND U563 ( .A(A[462]), .B(B[0]), .Z(PRODUCT[462]) );
  AND U564 ( .A(A[461]), .B(B[0]), .Z(PRODUCT[461]) );
  AND U565 ( .A(A[460]), .B(B[0]), .Z(PRODUCT[460]) );
  AND U566 ( .A(A[459]), .B(B[0]), .Z(PRODUCT[459]) );
  AND U567 ( .A(A[458]), .B(B[0]), .Z(PRODUCT[458]) );
  AND U568 ( .A(A[457]), .B(B[0]), .Z(PRODUCT[457]) );
  AND U569 ( .A(A[456]), .B(B[0]), .Z(PRODUCT[456]) );
  AND U570 ( .A(A[455]), .B(B[0]), .Z(PRODUCT[455]) );
  AND U571 ( .A(A[454]), .B(B[0]), .Z(PRODUCT[454]) );
  AND U572 ( .A(A[453]), .B(B[0]), .Z(PRODUCT[453]) );
  AND U573 ( .A(A[452]), .B(B[0]), .Z(PRODUCT[452]) );
  AND U574 ( .A(A[451]), .B(B[0]), .Z(PRODUCT[451]) );
  AND U575 ( .A(A[450]), .B(B[0]), .Z(PRODUCT[450]) );
  AND U576 ( .A(A[449]), .B(B[0]), .Z(PRODUCT[449]) );
  AND U577 ( .A(A[448]), .B(B[0]), .Z(PRODUCT[448]) );
  AND U578 ( .A(A[447]), .B(B[0]), .Z(PRODUCT[447]) );
  AND U579 ( .A(A[446]), .B(B[0]), .Z(PRODUCT[446]) );
  AND U580 ( .A(A[445]), .B(B[0]), .Z(PRODUCT[445]) );
  AND U581 ( .A(A[444]), .B(B[0]), .Z(PRODUCT[444]) );
  AND U582 ( .A(A[443]), .B(B[0]), .Z(PRODUCT[443]) );
  AND U583 ( .A(A[442]), .B(B[0]), .Z(PRODUCT[442]) );
  AND U584 ( .A(A[441]), .B(B[0]), .Z(PRODUCT[441]) );
  AND U585 ( .A(A[440]), .B(B[0]), .Z(PRODUCT[440]) );
  AND U586 ( .A(A[439]), .B(B[0]), .Z(PRODUCT[439]) );
  AND U587 ( .A(A[438]), .B(B[0]), .Z(PRODUCT[438]) );
  AND U588 ( .A(A[437]), .B(B[0]), .Z(PRODUCT[437]) );
  AND U589 ( .A(A[436]), .B(B[0]), .Z(PRODUCT[436]) );
  AND U590 ( .A(A[435]), .B(B[0]), .Z(PRODUCT[435]) );
  AND U591 ( .A(A[434]), .B(B[0]), .Z(PRODUCT[434]) );
  AND U592 ( .A(A[433]), .B(B[0]), .Z(PRODUCT[433]) );
  AND U593 ( .A(A[432]), .B(B[0]), .Z(PRODUCT[432]) );
  AND U594 ( .A(A[431]), .B(B[0]), .Z(PRODUCT[431]) );
  AND U595 ( .A(A[430]), .B(B[0]), .Z(PRODUCT[430]) );
  AND U596 ( .A(A[429]), .B(B[0]), .Z(PRODUCT[429]) );
  AND U597 ( .A(A[428]), .B(B[0]), .Z(PRODUCT[428]) );
  AND U598 ( .A(A[427]), .B(B[0]), .Z(PRODUCT[427]) );
  AND U599 ( .A(A[426]), .B(B[0]), .Z(PRODUCT[426]) );
  AND U600 ( .A(A[425]), .B(B[0]), .Z(PRODUCT[425]) );
  AND U601 ( .A(A[424]), .B(B[0]), .Z(PRODUCT[424]) );
  AND U602 ( .A(A[423]), .B(B[0]), .Z(PRODUCT[423]) );
  AND U603 ( .A(A[422]), .B(B[0]), .Z(PRODUCT[422]) );
  AND U604 ( .A(A[421]), .B(B[0]), .Z(PRODUCT[421]) );
  AND U605 ( .A(A[420]), .B(B[0]), .Z(PRODUCT[420]) );
  AND U606 ( .A(A[419]), .B(B[0]), .Z(PRODUCT[419]) );
  AND U607 ( .A(A[418]), .B(B[0]), .Z(PRODUCT[418]) );
  AND U608 ( .A(A[417]), .B(B[0]), .Z(PRODUCT[417]) );
  AND U609 ( .A(A[416]), .B(B[0]), .Z(PRODUCT[416]) );
  AND U610 ( .A(A[415]), .B(B[0]), .Z(PRODUCT[415]) );
  AND U611 ( .A(A[414]), .B(B[0]), .Z(PRODUCT[414]) );
  AND U612 ( .A(A[413]), .B(B[0]), .Z(PRODUCT[413]) );
  AND U613 ( .A(A[412]), .B(B[0]), .Z(PRODUCT[412]) );
  AND U614 ( .A(A[411]), .B(B[0]), .Z(PRODUCT[411]) );
  AND U615 ( .A(A[410]), .B(B[0]), .Z(PRODUCT[410]) );
  AND U616 ( .A(A[409]), .B(B[0]), .Z(PRODUCT[409]) );
  AND U617 ( .A(A[408]), .B(B[0]), .Z(PRODUCT[408]) );
  AND U618 ( .A(A[407]), .B(B[0]), .Z(PRODUCT[407]) );
  AND U619 ( .A(A[406]), .B(B[0]), .Z(PRODUCT[406]) );
  AND U620 ( .A(A[405]), .B(B[0]), .Z(PRODUCT[405]) );
  AND U621 ( .A(A[404]), .B(B[0]), .Z(PRODUCT[404]) );
  AND U622 ( .A(A[403]), .B(B[0]), .Z(PRODUCT[403]) );
  AND U623 ( .A(A[402]), .B(B[0]), .Z(PRODUCT[402]) );
  AND U624 ( .A(A[401]), .B(B[0]), .Z(PRODUCT[401]) );
  AND U625 ( .A(A[400]), .B(B[0]), .Z(PRODUCT[400]) );
  AND U626 ( .A(A[399]), .B(B[0]), .Z(PRODUCT[399]) );
  AND U627 ( .A(A[398]), .B(B[0]), .Z(PRODUCT[398]) );
  AND U628 ( .A(A[397]), .B(B[0]), .Z(PRODUCT[397]) );
  AND U629 ( .A(A[396]), .B(B[0]), .Z(PRODUCT[396]) );
  AND U630 ( .A(A[395]), .B(B[0]), .Z(PRODUCT[395]) );
  AND U631 ( .A(A[394]), .B(B[0]), .Z(PRODUCT[394]) );
  AND U632 ( .A(A[393]), .B(B[0]), .Z(PRODUCT[393]) );
  AND U633 ( .A(A[392]), .B(B[0]), .Z(PRODUCT[392]) );
  AND U634 ( .A(A[391]), .B(B[0]), .Z(PRODUCT[391]) );
  AND U635 ( .A(A[390]), .B(B[0]), .Z(PRODUCT[390]) );
  AND U636 ( .A(A[389]), .B(B[0]), .Z(PRODUCT[389]) );
  AND U637 ( .A(A[388]), .B(B[0]), .Z(PRODUCT[388]) );
  AND U638 ( .A(A[387]), .B(B[0]), .Z(PRODUCT[387]) );
  AND U639 ( .A(A[386]), .B(B[0]), .Z(PRODUCT[386]) );
  AND U640 ( .A(A[385]), .B(B[0]), .Z(PRODUCT[385]) );
  AND U641 ( .A(A[384]), .B(B[0]), .Z(PRODUCT[384]) );
  AND U642 ( .A(A[383]), .B(B[0]), .Z(PRODUCT[383]) );
  AND U643 ( .A(A[382]), .B(B[0]), .Z(PRODUCT[382]) );
  AND U644 ( .A(A[381]), .B(B[0]), .Z(PRODUCT[381]) );
  AND U645 ( .A(A[380]), .B(B[0]), .Z(PRODUCT[380]) );
  AND U646 ( .A(A[379]), .B(B[0]), .Z(PRODUCT[379]) );
  AND U647 ( .A(A[378]), .B(B[0]), .Z(PRODUCT[378]) );
  AND U648 ( .A(A[377]), .B(B[0]), .Z(PRODUCT[377]) );
  AND U649 ( .A(A[376]), .B(B[0]), .Z(PRODUCT[376]) );
  AND U650 ( .A(A[375]), .B(B[0]), .Z(PRODUCT[375]) );
  AND U651 ( .A(A[374]), .B(B[0]), .Z(PRODUCT[374]) );
  AND U652 ( .A(A[373]), .B(B[0]), .Z(PRODUCT[373]) );
  AND U653 ( .A(A[372]), .B(B[0]), .Z(PRODUCT[372]) );
  AND U654 ( .A(A[371]), .B(B[0]), .Z(PRODUCT[371]) );
  AND U655 ( .A(A[370]), .B(B[0]), .Z(PRODUCT[370]) );
  AND U656 ( .A(A[369]), .B(B[0]), .Z(PRODUCT[369]) );
  AND U657 ( .A(A[368]), .B(B[0]), .Z(PRODUCT[368]) );
  AND U658 ( .A(A[367]), .B(B[0]), .Z(PRODUCT[367]) );
  AND U659 ( .A(A[366]), .B(B[0]), .Z(PRODUCT[366]) );
  AND U660 ( .A(A[365]), .B(B[0]), .Z(PRODUCT[365]) );
  AND U661 ( .A(A[364]), .B(B[0]), .Z(PRODUCT[364]) );
  AND U662 ( .A(A[363]), .B(B[0]), .Z(PRODUCT[363]) );
  AND U663 ( .A(A[362]), .B(B[0]), .Z(PRODUCT[362]) );
  AND U664 ( .A(A[361]), .B(B[0]), .Z(PRODUCT[361]) );
  AND U665 ( .A(A[360]), .B(B[0]), .Z(PRODUCT[360]) );
  AND U666 ( .A(A[359]), .B(B[0]), .Z(PRODUCT[359]) );
  AND U667 ( .A(A[358]), .B(B[0]), .Z(PRODUCT[358]) );
  AND U668 ( .A(A[357]), .B(B[0]), .Z(PRODUCT[357]) );
  AND U669 ( .A(A[356]), .B(B[0]), .Z(PRODUCT[356]) );
  AND U670 ( .A(A[355]), .B(B[0]), .Z(PRODUCT[355]) );
  AND U671 ( .A(A[354]), .B(B[0]), .Z(PRODUCT[354]) );
  AND U672 ( .A(A[353]), .B(B[0]), .Z(PRODUCT[353]) );
  AND U673 ( .A(A[352]), .B(B[0]), .Z(PRODUCT[352]) );
  AND U674 ( .A(A[351]), .B(B[0]), .Z(PRODUCT[351]) );
  AND U675 ( .A(A[350]), .B(B[0]), .Z(PRODUCT[350]) );
  AND U676 ( .A(A[349]), .B(B[0]), .Z(PRODUCT[349]) );
  AND U677 ( .A(A[348]), .B(B[0]), .Z(PRODUCT[348]) );
  AND U678 ( .A(A[347]), .B(B[0]), .Z(PRODUCT[347]) );
  AND U679 ( .A(A[346]), .B(B[0]), .Z(PRODUCT[346]) );
  AND U680 ( .A(A[345]), .B(B[0]), .Z(PRODUCT[345]) );
  AND U681 ( .A(A[344]), .B(B[0]), .Z(PRODUCT[344]) );
  AND U682 ( .A(A[343]), .B(B[0]), .Z(PRODUCT[343]) );
  AND U683 ( .A(A[342]), .B(B[0]), .Z(PRODUCT[342]) );
  AND U684 ( .A(A[341]), .B(B[0]), .Z(PRODUCT[341]) );
  AND U685 ( .A(A[340]), .B(B[0]), .Z(PRODUCT[340]) );
  AND U686 ( .A(A[339]), .B(B[0]), .Z(PRODUCT[339]) );
  AND U687 ( .A(A[338]), .B(B[0]), .Z(PRODUCT[338]) );
  AND U688 ( .A(A[337]), .B(B[0]), .Z(PRODUCT[337]) );
  AND U689 ( .A(A[336]), .B(B[0]), .Z(PRODUCT[336]) );
  AND U690 ( .A(A[335]), .B(B[0]), .Z(PRODUCT[335]) );
  AND U691 ( .A(A[334]), .B(B[0]), .Z(PRODUCT[334]) );
  AND U692 ( .A(A[333]), .B(B[0]), .Z(PRODUCT[333]) );
  AND U693 ( .A(A[332]), .B(B[0]), .Z(PRODUCT[332]) );
  AND U694 ( .A(A[331]), .B(B[0]), .Z(PRODUCT[331]) );
  AND U695 ( .A(A[330]), .B(B[0]), .Z(PRODUCT[330]) );
  AND U696 ( .A(A[329]), .B(B[0]), .Z(PRODUCT[329]) );
  AND U697 ( .A(A[328]), .B(B[0]), .Z(PRODUCT[328]) );
  AND U698 ( .A(A[327]), .B(B[0]), .Z(PRODUCT[327]) );
  AND U699 ( .A(A[326]), .B(B[0]), .Z(PRODUCT[326]) );
  AND U700 ( .A(A[325]), .B(B[0]), .Z(PRODUCT[325]) );
  AND U701 ( .A(A[324]), .B(B[0]), .Z(PRODUCT[324]) );
  AND U702 ( .A(A[323]), .B(B[0]), .Z(PRODUCT[323]) );
  AND U703 ( .A(A[322]), .B(B[0]), .Z(PRODUCT[322]) );
  AND U704 ( .A(A[321]), .B(B[0]), .Z(PRODUCT[321]) );
  AND U705 ( .A(A[320]), .B(B[0]), .Z(PRODUCT[320]) );
  AND U706 ( .A(A[319]), .B(B[0]), .Z(PRODUCT[319]) );
  AND U707 ( .A(A[318]), .B(B[0]), .Z(PRODUCT[318]) );
  AND U708 ( .A(A[317]), .B(B[0]), .Z(PRODUCT[317]) );
  AND U709 ( .A(A[316]), .B(B[0]), .Z(PRODUCT[316]) );
  AND U710 ( .A(A[315]), .B(B[0]), .Z(PRODUCT[315]) );
  AND U711 ( .A(A[314]), .B(B[0]), .Z(PRODUCT[314]) );
  AND U712 ( .A(A[313]), .B(B[0]), .Z(PRODUCT[313]) );
  AND U713 ( .A(A[312]), .B(B[0]), .Z(PRODUCT[312]) );
  AND U714 ( .A(A[311]), .B(B[0]), .Z(PRODUCT[311]) );
  AND U715 ( .A(A[310]), .B(B[0]), .Z(PRODUCT[310]) );
  AND U716 ( .A(A[309]), .B(B[0]), .Z(PRODUCT[309]) );
  AND U717 ( .A(A[308]), .B(B[0]), .Z(PRODUCT[308]) );
  AND U718 ( .A(A[307]), .B(B[0]), .Z(PRODUCT[307]) );
  AND U719 ( .A(A[306]), .B(B[0]), .Z(PRODUCT[306]) );
  AND U720 ( .A(A[305]), .B(B[0]), .Z(PRODUCT[305]) );
  AND U721 ( .A(A[304]), .B(B[0]), .Z(PRODUCT[304]) );
  AND U722 ( .A(A[303]), .B(B[0]), .Z(PRODUCT[303]) );
  AND U723 ( .A(A[302]), .B(B[0]), .Z(PRODUCT[302]) );
  AND U724 ( .A(A[301]), .B(B[0]), .Z(PRODUCT[301]) );
  AND U725 ( .A(A[300]), .B(B[0]), .Z(PRODUCT[300]) );
  AND U726 ( .A(A[299]), .B(B[0]), .Z(PRODUCT[299]) );
  AND U727 ( .A(A[298]), .B(B[0]), .Z(PRODUCT[298]) );
  AND U728 ( .A(A[297]), .B(B[0]), .Z(PRODUCT[297]) );
  AND U729 ( .A(A[296]), .B(B[0]), .Z(PRODUCT[296]) );
  AND U730 ( .A(A[295]), .B(B[0]), .Z(PRODUCT[295]) );
  AND U731 ( .A(A[294]), .B(B[0]), .Z(PRODUCT[294]) );
  AND U732 ( .A(A[293]), .B(B[0]), .Z(PRODUCT[293]) );
  AND U733 ( .A(A[292]), .B(B[0]), .Z(PRODUCT[292]) );
  AND U734 ( .A(A[291]), .B(B[0]), .Z(PRODUCT[291]) );
  AND U735 ( .A(A[290]), .B(B[0]), .Z(PRODUCT[290]) );
  AND U736 ( .A(A[289]), .B(B[0]), .Z(PRODUCT[289]) );
  AND U737 ( .A(A[288]), .B(B[0]), .Z(PRODUCT[288]) );
  AND U738 ( .A(A[287]), .B(B[0]), .Z(PRODUCT[287]) );
  AND U739 ( .A(A[286]), .B(B[0]), .Z(PRODUCT[286]) );
  AND U740 ( .A(A[285]), .B(B[0]), .Z(PRODUCT[285]) );
  AND U741 ( .A(A[284]), .B(B[0]), .Z(PRODUCT[284]) );
  AND U742 ( .A(A[283]), .B(B[0]), .Z(PRODUCT[283]) );
  AND U743 ( .A(A[282]), .B(B[0]), .Z(PRODUCT[282]) );
  AND U744 ( .A(A[281]), .B(B[0]), .Z(PRODUCT[281]) );
  AND U745 ( .A(A[280]), .B(B[0]), .Z(PRODUCT[280]) );
  AND U746 ( .A(A[279]), .B(B[0]), .Z(PRODUCT[279]) );
  AND U747 ( .A(A[278]), .B(B[0]), .Z(PRODUCT[278]) );
  AND U748 ( .A(A[277]), .B(B[0]), .Z(PRODUCT[277]) );
  AND U749 ( .A(A[276]), .B(B[0]), .Z(PRODUCT[276]) );
  AND U750 ( .A(A[275]), .B(B[0]), .Z(PRODUCT[275]) );
  AND U751 ( .A(A[274]), .B(B[0]), .Z(PRODUCT[274]) );
  AND U752 ( .A(A[273]), .B(B[0]), .Z(PRODUCT[273]) );
  AND U753 ( .A(A[272]), .B(B[0]), .Z(PRODUCT[272]) );
  AND U754 ( .A(A[271]), .B(B[0]), .Z(PRODUCT[271]) );
  AND U755 ( .A(A[270]), .B(B[0]), .Z(PRODUCT[270]) );
  AND U756 ( .A(A[269]), .B(B[0]), .Z(PRODUCT[269]) );
  AND U757 ( .A(A[268]), .B(B[0]), .Z(PRODUCT[268]) );
  AND U758 ( .A(A[267]), .B(B[0]), .Z(PRODUCT[267]) );
  AND U759 ( .A(A[266]), .B(B[0]), .Z(PRODUCT[266]) );
  AND U760 ( .A(A[265]), .B(B[0]), .Z(PRODUCT[265]) );
  AND U761 ( .A(A[264]), .B(B[0]), .Z(PRODUCT[264]) );
  AND U762 ( .A(A[263]), .B(B[0]), .Z(PRODUCT[263]) );
  AND U763 ( .A(A[262]), .B(B[0]), .Z(PRODUCT[262]) );
  AND U764 ( .A(A[261]), .B(B[0]), .Z(PRODUCT[261]) );
  AND U765 ( .A(A[260]), .B(B[0]), .Z(PRODUCT[260]) );
  AND U766 ( .A(A[259]), .B(B[0]), .Z(PRODUCT[259]) );
  AND U767 ( .A(A[258]), .B(B[0]), .Z(PRODUCT[258]) );
  AND U768 ( .A(A[257]), .B(B[0]), .Z(PRODUCT[257]) );
  AND U769 ( .A(A[256]), .B(B[0]), .Z(PRODUCT[256]) );
  AND U770 ( .A(A[255]), .B(B[0]), .Z(PRODUCT[255]) );
  AND U771 ( .A(A[254]), .B(B[0]), .Z(PRODUCT[254]) );
  AND U772 ( .A(A[253]), .B(B[0]), .Z(PRODUCT[253]) );
  AND U773 ( .A(A[252]), .B(B[0]), .Z(PRODUCT[252]) );
  AND U774 ( .A(A[251]), .B(B[0]), .Z(PRODUCT[251]) );
  AND U775 ( .A(A[250]), .B(B[0]), .Z(PRODUCT[250]) );
  AND U776 ( .A(A[249]), .B(B[0]), .Z(PRODUCT[249]) );
  AND U777 ( .A(A[248]), .B(B[0]), .Z(PRODUCT[248]) );
  AND U778 ( .A(A[247]), .B(B[0]), .Z(PRODUCT[247]) );
  AND U779 ( .A(A[246]), .B(B[0]), .Z(PRODUCT[246]) );
  AND U780 ( .A(A[245]), .B(B[0]), .Z(PRODUCT[245]) );
  AND U781 ( .A(A[244]), .B(B[0]), .Z(PRODUCT[244]) );
  AND U782 ( .A(A[243]), .B(B[0]), .Z(PRODUCT[243]) );
  AND U783 ( .A(A[242]), .B(B[0]), .Z(PRODUCT[242]) );
  AND U784 ( .A(A[241]), .B(B[0]), .Z(PRODUCT[241]) );
  AND U785 ( .A(A[240]), .B(B[0]), .Z(PRODUCT[240]) );
  AND U786 ( .A(A[239]), .B(B[0]), .Z(PRODUCT[239]) );
  AND U787 ( .A(A[238]), .B(B[0]), .Z(PRODUCT[238]) );
  AND U788 ( .A(A[237]), .B(B[0]), .Z(PRODUCT[237]) );
  AND U789 ( .A(A[236]), .B(B[0]), .Z(PRODUCT[236]) );
  AND U790 ( .A(A[235]), .B(B[0]), .Z(PRODUCT[235]) );
  AND U791 ( .A(A[234]), .B(B[0]), .Z(PRODUCT[234]) );
  AND U792 ( .A(A[233]), .B(B[0]), .Z(PRODUCT[233]) );
  AND U793 ( .A(A[232]), .B(B[0]), .Z(PRODUCT[232]) );
  AND U794 ( .A(A[231]), .B(B[0]), .Z(PRODUCT[231]) );
  AND U795 ( .A(A[230]), .B(B[0]), .Z(PRODUCT[230]) );
  AND U796 ( .A(A[229]), .B(B[0]), .Z(PRODUCT[229]) );
  AND U797 ( .A(A[228]), .B(B[0]), .Z(PRODUCT[228]) );
  AND U798 ( .A(A[227]), .B(B[0]), .Z(PRODUCT[227]) );
  AND U799 ( .A(A[226]), .B(B[0]), .Z(PRODUCT[226]) );
  AND U800 ( .A(A[225]), .B(B[0]), .Z(PRODUCT[225]) );
  AND U801 ( .A(A[224]), .B(B[0]), .Z(PRODUCT[224]) );
  AND U802 ( .A(A[223]), .B(B[0]), .Z(PRODUCT[223]) );
  AND U803 ( .A(A[222]), .B(B[0]), .Z(PRODUCT[222]) );
  AND U804 ( .A(A[221]), .B(B[0]), .Z(PRODUCT[221]) );
  AND U805 ( .A(A[220]), .B(B[0]), .Z(PRODUCT[220]) );
  AND U806 ( .A(A[219]), .B(B[0]), .Z(PRODUCT[219]) );
  AND U807 ( .A(A[218]), .B(B[0]), .Z(PRODUCT[218]) );
  AND U808 ( .A(A[217]), .B(B[0]), .Z(PRODUCT[217]) );
  AND U809 ( .A(A[216]), .B(B[0]), .Z(PRODUCT[216]) );
  AND U810 ( .A(A[215]), .B(B[0]), .Z(PRODUCT[215]) );
  AND U811 ( .A(A[214]), .B(B[0]), .Z(PRODUCT[214]) );
  AND U812 ( .A(A[213]), .B(B[0]), .Z(PRODUCT[213]) );
  AND U813 ( .A(A[212]), .B(B[0]), .Z(PRODUCT[212]) );
  AND U814 ( .A(A[211]), .B(B[0]), .Z(PRODUCT[211]) );
  AND U815 ( .A(A[210]), .B(B[0]), .Z(PRODUCT[210]) );
  AND U816 ( .A(A[209]), .B(B[0]), .Z(PRODUCT[209]) );
  AND U817 ( .A(A[208]), .B(B[0]), .Z(PRODUCT[208]) );
  AND U818 ( .A(A[207]), .B(B[0]), .Z(PRODUCT[207]) );
  AND U819 ( .A(A[206]), .B(B[0]), .Z(PRODUCT[206]) );
  AND U820 ( .A(A[205]), .B(B[0]), .Z(PRODUCT[205]) );
  AND U821 ( .A(A[204]), .B(B[0]), .Z(PRODUCT[204]) );
  AND U822 ( .A(A[203]), .B(B[0]), .Z(PRODUCT[203]) );
  AND U823 ( .A(A[202]), .B(B[0]), .Z(PRODUCT[202]) );
  AND U824 ( .A(A[201]), .B(B[0]), .Z(PRODUCT[201]) );
  AND U825 ( .A(A[200]), .B(B[0]), .Z(PRODUCT[200]) );
  AND U826 ( .A(A[199]), .B(B[0]), .Z(PRODUCT[199]) );
  AND U827 ( .A(A[198]), .B(B[0]), .Z(PRODUCT[198]) );
  AND U828 ( .A(A[197]), .B(B[0]), .Z(PRODUCT[197]) );
  AND U829 ( .A(A[196]), .B(B[0]), .Z(PRODUCT[196]) );
  AND U830 ( .A(A[195]), .B(B[0]), .Z(PRODUCT[195]) );
  AND U831 ( .A(A[194]), .B(B[0]), .Z(PRODUCT[194]) );
  AND U832 ( .A(A[193]), .B(B[0]), .Z(PRODUCT[193]) );
  AND U833 ( .A(A[192]), .B(B[0]), .Z(PRODUCT[192]) );
  AND U834 ( .A(A[191]), .B(B[0]), .Z(PRODUCT[191]) );
  AND U835 ( .A(A[190]), .B(B[0]), .Z(PRODUCT[190]) );
  AND U836 ( .A(A[189]), .B(B[0]), .Z(PRODUCT[189]) );
  AND U837 ( .A(A[188]), .B(B[0]), .Z(PRODUCT[188]) );
  AND U838 ( .A(A[187]), .B(B[0]), .Z(PRODUCT[187]) );
  AND U839 ( .A(A[186]), .B(B[0]), .Z(PRODUCT[186]) );
  AND U840 ( .A(A[185]), .B(B[0]), .Z(PRODUCT[185]) );
  AND U841 ( .A(A[184]), .B(B[0]), .Z(PRODUCT[184]) );
  AND U842 ( .A(A[183]), .B(B[0]), .Z(PRODUCT[183]) );
  AND U843 ( .A(A[182]), .B(B[0]), .Z(PRODUCT[182]) );
  AND U844 ( .A(A[181]), .B(B[0]), .Z(PRODUCT[181]) );
  AND U845 ( .A(A[180]), .B(B[0]), .Z(PRODUCT[180]) );
  AND U846 ( .A(A[179]), .B(B[0]), .Z(PRODUCT[179]) );
  AND U847 ( .A(A[178]), .B(B[0]), .Z(PRODUCT[178]) );
  AND U848 ( .A(A[177]), .B(B[0]), .Z(PRODUCT[177]) );
  AND U849 ( .A(A[176]), .B(B[0]), .Z(PRODUCT[176]) );
  AND U850 ( .A(A[175]), .B(B[0]), .Z(PRODUCT[175]) );
  AND U851 ( .A(A[174]), .B(B[0]), .Z(PRODUCT[174]) );
  AND U852 ( .A(A[173]), .B(B[0]), .Z(PRODUCT[173]) );
  AND U853 ( .A(A[172]), .B(B[0]), .Z(PRODUCT[172]) );
  AND U854 ( .A(A[171]), .B(B[0]), .Z(PRODUCT[171]) );
  AND U855 ( .A(A[170]), .B(B[0]), .Z(PRODUCT[170]) );
  AND U856 ( .A(A[169]), .B(B[0]), .Z(PRODUCT[169]) );
  AND U857 ( .A(A[168]), .B(B[0]), .Z(PRODUCT[168]) );
  AND U858 ( .A(A[167]), .B(B[0]), .Z(PRODUCT[167]) );
  AND U859 ( .A(A[166]), .B(B[0]), .Z(PRODUCT[166]) );
  AND U860 ( .A(A[165]), .B(B[0]), .Z(PRODUCT[165]) );
  AND U861 ( .A(A[164]), .B(B[0]), .Z(PRODUCT[164]) );
  AND U862 ( .A(A[163]), .B(B[0]), .Z(PRODUCT[163]) );
  AND U863 ( .A(A[162]), .B(B[0]), .Z(PRODUCT[162]) );
  AND U864 ( .A(A[161]), .B(B[0]), .Z(PRODUCT[161]) );
  AND U865 ( .A(A[160]), .B(B[0]), .Z(PRODUCT[160]) );
  AND U866 ( .A(A[159]), .B(B[0]), .Z(PRODUCT[159]) );
  AND U867 ( .A(A[158]), .B(B[0]), .Z(PRODUCT[158]) );
  AND U868 ( .A(A[157]), .B(B[0]), .Z(PRODUCT[157]) );
  AND U869 ( .A(A[156]), .B(B[0]), .Z(PRODUCT[156]) );
  AND U870 ( .A(A[155]), .B(B[0]), .Z(PRODUCT[155]) );
  AND U871 ( .A(A[154]), .B(B[0]), .Z(PRODUCT[154]) );
  AND U872 ( .A(A[153]), .B(B[0]), .Z(PRODUCT[153]) );
  AND U873 ( .A(A[152]), .B(B[0]), .Z(PRODUCT[152]) );
  AND U874 ( .A(A[151]), .B(B[0]), .Z(PRODUCT[151]) );
  AND U875 ( .A(A[150]), .B(B[0]), .Z(PRODUCT[150]) );
  AND U876 ( .A(A[149]), .B(B[0]), .Z(PRODUCT[149]) );
  AND U877 ( .A(A[148]), .B(B[0]), .Z(PRODUCT[148]) );
  AND U878 ( .A(A[147]), .B(B[0]), .Z(PRODUCT[147]) );
  AND U879 ( .A(A[146]), .B(B[0]), .Z(PRODUCT[146]) );
  AND U880 ( .A(A[145]), .B(B[0]), .Z(PRODUCT[145]) );
  AND U881 ( .A(A[144]), .B(B[0]), .Z(PRODUCT[144]) );
  AND U882 ( .A(A[143]), .B(B[0]), .Z(PRODUCT[143]) );
  AND U883 ( .A(A[142]), .B(B[0]), .Z(PRODUCT[142]) );
  AND U884 ( .A(A[141]), .B(B[0]), .Z(PRODUCT[141]) );
  AND U885 ( .A(A[140]), .B(B[0]), .Z(PRODUCT[140]) );
  AND U886 ( .A(A[139]), .B(B[0]), .Z(PRODUCT[139]) );
  AND U887 ( .A(A[138]), .B(B[0]), .Z(PRODUCT[138]) );
  AND U888 ( .A(A[137]), .B(B[0]), .Z(PRODUCT[137]) );
  AND U889 ( .A(A[136]), .B(B[0]), .Z(PRODUCT[136]) );
  AND U890 ( .A(A[135]), .B(B[0]), .Z(PRODUCT[135]) );
  AND U891 ( .A(A[134]), .B(B[0]), .Z(PRODUCT[134]) );
  AND U892 ( .A(A[133]), .B(B[0]), .Z(PRODUCT[133]) );
  AND U893 ( .A(A[132]), .B(B[0]), .Z(PRODUCT[132]) );
  AND U894 ( .A(A[131]), .B(B[0]), .Z(PRODUCT[131]) );
  AND U895 ( .A(A[130]), .B(B[0]), .Z(PRODUCT[130]) );
  AND U896 ( .A(A[129]), .B(B[0]), .Z(PRODUCT[129]) );
  AND U897 ( .A(A[128]), .B(B[0]), .Z(PRODUCT[128]) );
  AND U898 ( .A(A[127]), .B(B[0]), .Z(PRODUCT[127]) );
  AND U899 ( .A(A[126]), .B(B[0]), .Z(PRODUCT[126]) );
  AND U900 ( .A(A[125]), .B(B[0]), .Z(PRODUCT[125]) );
  AND U901 ( .A(A[124]), .B(B[0]), .Z(PRODUCT[124]) );
  AND U902 ( .A(A[123]), .B(B[0]), .Z(PRODUCT[123]) );
  AND U903 ( .A(A[122]), .B(B[0]), .Z(PRODUCT[122]) );
  AND U904 ( .A(A[121]), .B(B[0]), .Z(PRODUCT[121]) );
  AND U905 ( .A(A[120]), .B(B[0]), .Z(PRODUCT[120]) );
  AND U906 ( .A(A[119]), .B(B[0]), .Z(PRODUCT[119]) );
  AND U907 ( .A(A[118]), .B(B[0]), .Z(PRODUCT[118]) );
  AND U908 ( .A(A[117]), .B(B[0]), .Z(PRODUCT[117]) );
  AND U909 ( .A(A[116]), .B(B[0]), .Z(PRODUCT[116]) );
  AND U910 ( .A(A[115]), .B(B[0]), .Z(PRODUCT[115]) );
  AND U911 ( .A(A[114]), .B(B[0]), .Z(PRODUCT[114]) );
  AND U912 ( .A(A[113]), .B(B[0]), .Z(PRODUCT[113]) );
  AND U913 ( .A(A[112]), .B(B[0]), .Z(PRODUCT[112]) );
  AND U914 ( .A(A[111]), .B(B[0]), .Z(PRODUCT[111]) );
  AND U915 ( .A(A[110]), .B(B[0]), .Z(PRODUCT[110]) );
  AND U916 ( .A(A[109]), .B(B[0]), .Z(PRODUCT[109]) );
  AND U917 ( .A(A[108]), .B(B[0]), .Z(PRODUCT[108]) );
  AND U918 ( .A(A[107]), .B(B[0]), .Z(PRODUCT[107]) );
  AND U919 ( .A(A[106]), .B(B[0]), .Z(PRODUCT[106]) );
  AND U920 ( .A(A[105]), .B(B[0]), .Z(PRODUCT[105]) );
  AND U921 ( .A(A[104]), .B(B[0]), .Z(PRODUCT[104]) );
  AND U922 ( .A(A[103]), .B(B[0]), .Z(PRODUCT[103]) );
  AND U923 ( .A(A[102]), .B(B[0]), .Z(PRODUCT[102]) );
  AND U924 ( .A(A[101]), .B(B[0]), .Z(PRODUCT[101]) );
  AND U925 ( .A(A[100]), .B(B[0]), .Z(PRODUCT[100]) );
  AND U926 ( .A(A[99]), .B(B[0]), .Z(PRODUCT[99]) );
  AND U927 ( .A(A[98]), .B(B[0]), .Z(PRODUCT[98]) );
  AND U928 ( .A(A[97]), .B(B[0]), .Z(PRODUCT[97]) );
  AND U929 ( .A(A[96]), .B(B[0]), .Z(PRODUCT[96]) );
  AND U930 ( .A(A[95]), .B(B[0]), .Z(PRODUCT[95]) );
  AND U931 ( .A(A[94]), .B(B[0]), .Z(PRODUCT[94]) );
  AND U932 ( .A(A[93]), .B(B[0]), .Z(PRODUCT[93]) );
  AND U933 ( .A(A[92]), .B(B[0]), .Z(PRODUCT[92]) );
  AND U934 ( .A(A[91]), .B(B[0]), .Z(PRODUCT[91]) );
  AND U935 ( .A(A[90]), .B(B[0]), .Z(PRODUCT[90]) );
  AND U936 ( .A(A[89]), .B(B[0]), .Z(PRODUCT[89]) );
  AND U937 ( .A(A[88]), .B(B[0]), .Z(PRODUCT[88]) );
  AND U938 ( .A(A[87]), .B(B[0]), .Z(PRODUCT[87]) );
  AND U939 ( .A(A[86]), .B(B[0]), .Z(PRODUCT[86]) );
  AND U940 ( .A(A[85]), .B(B[0]), .Z(PRODUCT[85]) );
  AND U941 ( .A(A[84]), .B(B[0]), .Z(PRODUCT[84]) );
  AND U942 ( .A(A[83]), .B(B[0]), .Z(PRODUCT[83]) );
  AND U943 ( .A(A[82]), .B(B[0]), .Z(PRODUCT[82]) );
  AND U944 ( .A(A[81]), .B(B[0]), .Z(PRODUCT[81]) );
  AND U945 ( .A(A[80]), .B(B[0]), .Z(PRODUCT[80]) );
  AND U946 ( .A(A[79]), .B(B[0]), .Z(PRODUCT[79]) );
  AND U947 ( .A(A[78]), .B(B[0]), .Z(PRODUCT[78]) );
  AND U948 ( .A(A[77]), .B(B[0]), .Z(PRODUCT[77]) );
  AND U949 ( .A(A[76]), .B(B[0]), .Z(PRODUCT[76]) );
  AND U950 ( .A(A[75]), .B(B[0]), .Z(PRODUCT[75]) );
  AND U951 ( .A(A[74]), .B(B[0]), .Z(PRODUCT[74]) );
  AND U952 ( .A(A[73]), .B(B[0]), .Z(PRODUCT[73]) );
  AND U953 ( .A(A[72]), .B(B[0]), .Z(PRODUCT[72]) );
  AND U954 ( .A(A[71]), .B(B[0]), .Z(PRODUCT[71]) );
  AND U955 ( .A(A[70]), .B(B[0]), .Z(PRODUCT[70]) );
  AND U956 ( .A(A[69]), .B(B[0]), .Z(PRODUCT[69]) );
  AND U957 ( .A(A[68]), .B(B[0]), .Z(PRODUCT[68]) );
  AND U958 ( .A(A[67]), .B(B[0]), .Z(PRODUCT[67]) );
  AND U959 ( .A(A[66]), .B(B[0]), .Z(PRODUCT[66]) );
  AND U960 ( .A(A[65]), .B(B[0]), .Z(PRODUCT[65]) );
  AND U961 ( .A(A[64]), .B(B[0]), .Z(PRODUCT[64]) );
  AND U962 ( .A(A[63]), .B(B[0]), .Z(PRODUCT[63]) );
  AND U963 ( .A(A[62]), .B(B[0]), .Z(PRODUCT[62]) );
  AND U964 ( .A(A[61]), .B(B[0]), .Z(PRODUCT[61]) );
  AND U965 ( .A(A[60]), .B(B[0]), .Z(PRODUCT[60]) );
  AND U966 ( .A(A[59]), .B(B[0]), .Z(PRODUCT[59]) );
  AND U967 ( .A(A[58]), .B(B[0]), .Z(PRODUCT[58]) );
  AND U968 ( .A(A[57]), .B(B[0]), .Z(PRODUCT[57]) );
  AND U969 ( .A(A[56]), .B(B[0]), .Z(PRODUCT[56]) );
  AND U970 ( .A(A[55]), .B(B[0]), .Z(PRODUCT[55]) );
  AND U971 ( .A(A[54]), .B(B[0]), .Z(PRODUCT[54]) );
  AND U972 ( .A(A[53]), .B(B[0]), .Z(PRODUCT[53]) );
  AND U973 ( .A(A[52]), .B(B[0]), .Z(PRODUCT[52]) );
  AND U974 ( .A(A[51]), .B(B[0]), .Z(PRODUCT[51]) );
  AND U975 ( .A(A[50]), .B(B[0]), .Z(PRODUCT[50]) );
  AND U976 ( .A(A[49]), .B(B[0]), .Z(PRODUCT[49]) );
  AND U977 ( .A(A[48]), .B(B[0]), .Z(PRODUCT[48]) );
  AND U978 ( .A(A[47]), .B(B[0]), .Z(PRODUCT[47]) );
  AND U979 ( .A(A[46]), .B(B[0]), .Z(PRODUCT[46]) );
  AND U980 ( .A(A[45]), .B(B[0]), .Z(PRODUCT[45]) );
  AND U981 ( .A(A[44]), .B(B[0]), .Z(PRODUCT[44]) );
  AND U982 ( .A(A[43]), .B(B[0]), .Z(PRODUCT[43]) );
  AND U983 ( .A(A[42]), .B(B[0]), .Z(PRODUCT[42]) );
  AND U984 ( .A(A[41]), .B(B[0]), .Z(PRODUCT[41]) );
  AND U985 ( .A(A[40]), .B(B[0]), .Z(PRODUCT[40]) );
  AND U986 ( .A(A[39]), .B(B[0]), .Z(PRODUCT[39]) );
  AND U987 ( .A(A[38]), .B(B[0]), .Z(PRODUCT[38]) );
  AND U988 ( .A(A[37]), .B(B[0]), .Z(PRODUCT[37]) );
  AND U989 ( .A(A[36]), .B(B[0]), .Z(PRODUCT[36]) );
  AND U990 ( .A(A[35]), .B(B[0]), .Z(PRODUCT[35]) );
  AND U991 ( .A(A[34]), .B(B[0]), .Z(PRODUCT[34]) );
  AND U992 ( .A(A[33]), .B(B[0]), .Z(PRODUCT[33]) );
  AND U993 ( .A(A[32]), .B(B[0]), .Z(PRODUCT[32]) );
  AND U994 ( .A(A[31]), .B(B[0]), .Z(PRODUCT[31]) );
  AND U995 ( .A(A[30]), .B(B[0]), .Z(PRODUCT[30]) );
  AND U996 ( .A(A[29]), .B(B[0]), .Z(PRODUCT[29]) );
  AND U997 ( .A(A[28]), .B(B[0]), .Z(PRODUCT[28]) );
  AND U998 ( .A(A[27]), .B(B[0]), .Z(PRODUCT[27]) );
  AND U999 ( .A(A[26]), .B(B[0]), .Z(PRODUCT[26]) );
  AND U1000 ( .A(A[25]), .B(B[0]), .Z(PRODUCT[25]) );
  AND U1001 ( .A(A[24]), .B(B[0]), .Z(PRODUCT[24]) );
  AND U1002 ( .A(A[23]), .B(B[0]), .Z(PRODUCT[23]) );
  AND U1003 ( .A(A[22]), .B(B[0]), .Z(PRODUCT[22]) );
  AND U1004 ( .A(A[21]), .B(B[0]), .Z(PRODUCT[21]) );
  AND U1005 ( .A(A[20]), .B(B[0]), .Z(PRODUCT[20]) );
  AND U1006 ( .A(A[19]), .B(B[0]), .Z(PRODUCT[19]) );
  AND U1007 ( .A(A[18]), .B(B[0]), .Z(PRODUCT[18]) );
  AND U1008 ( .A(A[17]), .B(B[0]), .Z(PRODUCT[17]) );
  AND U1009 ( .A(A[16]), .B(B[0]), .Z(PRODUCT[16]) );
  AND U1010 ( .A(A[15]), .B(B[0]), .Z(PRODUCT[15]) );
  AND U1011 ( .A(A[14]), .B(B[0]), .Z(PRODUCT[14]) );
  AND U1012 ( .A(A[13]), .B(B[0]), .Z(PRODUCT[13]) );
  AND U1013 ( .A(A[12]), .B(B[0]), .Z(PRODUCT[12]) );
  AND U1014 ( .A(A[11]), .B(B[0]), .Z(PRODUCT[11]) );
  AND U1015 ( .A(A[10]), .B(B[0]), .Z(PRODUCT[10]) );
  AND U1016 ( .A(B[0]), .B(A[9]), .Z(PRODUCT[9]) );
  AND U1017 ( .A(A[8]), .B(B[0]), .Z(PRODUCT[8]) );
  AND U1018 ( .A(A[7]), .B(B[0]), .Z(PRODUCT[7]) );
  AND U1019 ( .A(A[6]), .B(B[0]), .Z(PRODUCT[6]) );
  AND U1020 ( .A(A[5]), .B(B[0]), .Z(PRODUCT[5]) );
  AND U1021 ( .A(A[4]), .B(B[0]), .Z(PRODUCT[4]) );
  AND U1022 ( .A(A[3]), .B(B[0]), .Z(PRODUCT[3]) );
  AND U1023 ( .A(A[2]), .B(B[0]), .Z(PRODUCT[2]) );
  AND U1024 ( .A(A[1]), .B(B[0]), .Z(PRODUCT[1]) );
  AND U1025 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
endmodule


module modmult_step_N1024_DW01_cmp2_0 ( A, B, LEQ, TC, LT_LE, GE_GT );
  input [1025:0] A;
  input [1025:0] B;
  input LEQ, TC;
  output LT_LE, GE_GT;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094;

  NAND U1 ( .A(n1), .B(n2), .Z(LT_LE) );
  NOR U2 ( .A(B[1025]), .B(B[1024]), .Z(n2) );
  AND U3 ( .A(n3), .B(n4), .Z(n1) );
  NAND U4 ( .A(n5), .B(n6), .Z(n4) );
  NANDN U5 ( .A(B[1023]), .B(A[1023]), .Z(n6) );
  NAND U6 ( .A(n7), .B(n8), .Z(n5) );
  NANDN U7 ( .A(A[1022]), .B(B[1022]), .Z(n8) );
  NAND U8 ( .A(n9), .B(n10), .Z(n7) );
  NANDN U9 ( .A(B[1022]), .B(A[1022]), .Z(n10) );
  AND U10 ( .A(n11), .B(n12), .Z(n9) );
  NAND U11 ( .A(n13), .B(n14), .Z(n12) );
  NANDN U12 ( .A(A[1021]), .B(B[1021]), .Z(n14) );
  AND U13 ( .A(n15), .B(n16), .Z(n13) );
  NANDN U14 ( .A(A[1020]), .B(B[1020]), .Z(n16) );
  NAND U15 ( .A(n17), .B(n18), .Z(n15) );
  NANDN U16 ( .A(B[1020]), .B(A[1020]), .Z(n18) );
  AND U17 ( .A(n19), .B(n20), .Z(n17) );
  NAND U18 ( .A(n21), .B(n22), .Z(n20) );
  NANDN U19 ( .A(A[1019]), .B(B[1019]), .Z(n22) );
  AND U20 ( .A(n23), .B(n24), .Z(n21) );
  NANDN U21 ( .A(A[1018]), .B(B[1018]), .Z(n24) );
  NAND U22 ( .A(n25), .B(n26), .Z(n23) );
  NANDN U23 ( .A(B[1018]), .B(A[1018]), .Z(n26) );
  AND U24 ( .A(n27), .B(n28), .Z(n25) );
  NAND U25 ( .A(n29), .B(n30), .Z(n28) );
  NANDN U26 ( .A(A[1017]), .B(B[1017]), .Z(n30) );
  AND U27 ( .A(n31), .B(n32), .Z(n29) );
  NANDN U28 ( .A(A[1016]), .B(B[1016]), .Z(n32) );
  NAND U29 ( .A(n33), .B(n34), .Z(n31) );
  NANDN U30 ( .A(B[1016]), .B(A[1016]), .Z(n34) );
  AND U31 ( .A(n35), .B(n36), .Z(n33) );
  NAND U32 ( .A(n37), .B(n38), .Z(n36) );
  NANDN U33 ( .A(A[1015]), .B(B[1015]), .Z(n38) );
  AND U34 ( .A(n39), .B(n40), .Z(n37) );
  NANDN U35 ( .A(A[1014]), .B(B[1014]), .Z(n40) );
  NAND U36 ( .A(n41), .B(n42), .Z(n39) );
  NANDN U37 ( .A(B[1014]), .B(A[1014]), .Z(n42) );
  AND U38 ( .A(n43), .B(n44), .Z(n41) );
  NAND U39 ( .A(n45), .B(n46), .Z(n44) );
  NANDN U40 ( .A(A[1013]), .B(B[1013]), .Z(n46) );
  AND U41 ( .A(n47), .B(n48), .Z(n45) );
  NANDN U42 ( .A(A[1012]), .B(B[1012]), .Z(n48) );
  NAND U43 ( .A(n49), .B(n50), .Z(n47) );
  NANDN U44 ( .A(B[1012]), .B(A[1012]), .Z(n50) );
  AND U45 ( .A(n51), .B(n52), .Z(n49) );
  NAND U46 ( .A(n53), .B(n54), .Z(n52) );
  NANDN U47 ( .A(A[1011]), .B(B[1011]), .Z(n54) );
  AND U48 ( .A(n55), .B(n56), .Z(n53) );
  NANDN U49 ( .A(A[1010]), .B(B[1010]), .Z(n56) );
  NAND U50 ( .A(n57), .B(n58), .Z(n55) );
  NANDN U51 ( .A(B[1010]), .B(A[1010]), .Z(n58) );
  AND U52 ( .A(n59), .B(n60), .Z(n57) );
  NAND U53 ( .A(n61), .B(n62), .Z(n60) );
  NANDN U54 ( .A(A[1009]), .B(B[1009]), .Z(n62) );
  AND U55 ( .A(n63), .B(n64), .Z(n61) );
  NANDN U56 ( .A(A[1008]), .B(B[1008]), .Z(n64) );
  NAND U57 ( .A(n65), .B(n66), .Z(n63) );
  NANDN U58 ( .A(B[1008]), .B(A[1008]), .Z(n66) );
  AND U59 ( .A(n67), .B(n68), .Z(n65) );
  NAND U60 ( .A(n69), .B(n70), .Z(n68) );
  NANDN U61 ( .A(A[1007]), .B(B[1007]), .Z(n70) );
  AND U62 ( .A(n71), .B(n72), .Z(n69) );
  NANDN U63 ( .A(A[1006]), .B(B[1006]), .Z(n72) );
  NAND U64 ( .A(n73), .B(n74), .Z(n71) );
  NANDN U65 ( .A(B[1006]), .B(A[1006]), .Z(n74) );
  AND U66 ( .A(n75), .B(n76), .Z(n73) );
  NAND U67 ( .A(n77), .B(n78), .Z(n76) );
  NANDN U68 ( .A(A[1005]), .B(B[1005]), .Z(n78) );
  AND U69 ( .A(n79), .B(n80), .Z(n77) );
  NANDN U70 ( .A(A[1004]), .B(B[1004]), .Z(n80) );
  NAND U71 ( .A(n81), .B(n82), .Z(n79) );
  NANDN U72 ( .A(B[1004]), .B(A[1004]), .Z(n82) );
  AND U73 ( .A(n83), .B(n84), .Z(n81) );
  NAND U74 ( .A(n85), .B(n86), .Z(n84) );
  NANDN U75 ( .A(A[1003]), .B(B[1003]), .Z(n86) );
  AND U76 ( .A(n87), .B(n88), .Z(n85) );
  NANDN U77 ( .A(A[1002]), .B(B[1002]), .Z(n88) );
  NAND U78 ( .A(n89), .B(n90), .Z(n87) );
  NANDN U79 ( .A(B[1002]), .B(A[1002]), .Z(n90) );
  AND U80 ( .A(n91), .B(n92), .Z(n89) );
  NAND U81 ( .A(n93), .B(n94), .Z(n92) );
  NANDN U82 ( .A(A[1001]), .B(B[1001]), .Z(n94) );
  AND U83 ( .A(n95), .B(n96), .Z(n93) );
  NANDN U84 ( .A(A[1000]), .B(B[1000]), .Z(n96) );
  NAND U85 ( .A(n97), .B(n98), .Z(n95) );
  NANDN U86 ( .A(B[999]), .B(A[999]), .Z(n98) );
  AND U87 ( .A(n99), .B(n100), .Z(n97) );
  NAND U88 ( .A(n101), .B(n102), .Z(n100) );
  NANDN U89 ( .A(A[999]), .B(B[999]), .Z(n102) );
  AND U90 ( .A(n103), .B(n104), .Z(n101) );
  NANDN U91 ( .A(A[998]), .B(B[998]), .Z(n104) );
  NAND U92 ( .A(n105), .B(n106), .Z(n103) );
  NANDN U93 ( .A(B[998]), .B(A[998]), .Z(n106) );
  AND U94 ( .A(n107), .B(n108), .Z(n105) );
  NAND U95 ( .A(n109), .B(n110), .Z(n108) );
  NANDN U96 ( .A(A[997]), .B(B[997]), .Z(n110) );
  AND U97 ( .A(n111), .B(n112), .Z(n109) );
  NANDN U98 ( .A(A[996]), .B(B[996]), .Z(n112) );
  NAND U99 ( .A(n113), .B(n114), .Z(n111) );
  NANDN U100 ( .A(B[996]), .B(A[996]), .Z(n114) );
  AND U101 ( .A(n115), .B(n116), .Z(n113) );
  NAND U102 ( .A(n117), .B(n118), .Z(n116) );
  NANDN U103 ( .A(A[995]), .B(B[995]), .Z(n118) );
  AND U104 ( .A(n119), .B(n120), .Z(n117) );
  NANDN U105 ( .A(A[994]), .B(B[994]), .Z(n120) );
  NAND U106 ( .A(n121), .B(n122), .Z(n119) );
  NANDN U107 ( .A(B[994]), .B(A[994]), .Z(n122) );
  AND U108 ( .A(n123), .B(n124), .Z(n121) );
  NAND U109 ( .A(n125), .B(n126), .Z(n124) );
  NANDN U110 ( .A(A[993]), .B(B[993]), .Z(n126) );
  AND U111 ( .A(n127), .B(n128), .Z(n125) );
  NANDN U112 ( .A(A[992]), .B(B[992]), .Z(n128) );
  NAND U113 ( .A(n129), .B(n130), .Z(n127) );
  NANDN U114 ( .A(B[992]), .B(A[992]), .Z(n130) );
  AND U115 ( .A(n131), .B(n132), .Z(n129) );
  NAND U116 ( .A(n133), .B(n134), .Z(n132) );
  NANDN U117 ( .A(A[991]), .B(B[991]), .Z(n134) );
  AND U118 ( .A(n135), .B(n136), .Z(n133) );
  NANDN U119 ( .A(A[990]), .B(B[990]), .Z(n136) );
  NAND U120 ( .A(n137), .B(n138), .Z(n135) );
  NANDN U121 ( .A(B[990]), .B(A[990]), .Z(n138) );
  AND U122 ( .A(n139), .B(n140), .Z(n137) );
  NAND U123 ( .A(n141), .B(n142), .Z(n140) );
  NANDN U124 ( .A(A[989]), .B(B[989]), .Z(n142) );
  AND U125 ( .A(n143), .B(n144), .Z(n141) );
  NANDN U126 ( .A(A[988]), .B(B[988]), .Z(n144) );
  NAND U127 ( .A(n145), .B(n146), .Z(n143) );
  NANDN U128 ( .A(B[988]), .B(A[988]), .Z(n146) );
  AND U129 ( .A(n147), .B(n148), .Z(n145) );
  NAND U130 ( .A(n149), .B(n150), .Z(n148) );
  NANDN U131 ( .A(A[987]), .B(B[987]), .Z(n150) );
  AND U132 ( .A(n151), .B(n152), .Z(n149) );
  NANDN U133 ( .A(A[986]), .B(B[986]), .Z(n152) );
  NAND U134 ( .A(n153), .B(n154), .Z(n151) );
  NANDN U135 ( .A(B[986]), .B(A[986]), .Z(n154) );
  AND U136 ( .A(n155), .B(n156), .Z(n153) );
  NAND U137 ( .A(n157), .B(n158), .Z(n156) );
  NANDN U138 ( .A(A[985]), .B(B[985]), .Z(n158) );
  AND U139 ( .A(n159), .B(n160), .Z(n157) );
  NANDN U140 ( .A(A[984]), .B(B[984]), .Z(n160) );
  NAND U141 ( .A(n161), .B(n162), .Z(n159) );
  NANDN U142 ( .A(B[984]), .B(A[984]), .Z(n162) );
  AND U143 ( .A(n163), .B(n164), .Z(n161) );
  NAND U144 ( .A(n165), .B(n166), .Z(n164) );
  NANDN U145 ( .A(A[983]), .B(B[983]), .Z(n166) );
  AND U146 ( .A(n167), .B(n168), .Z(n165) );
  NANDN U147 ( .A(A[982]), .B(B[982]), .Z(n168) );
  NAND U148 ( .A(n169), .B(n170), .Z(n167) );
  NANDN U149 ( .A(B[982]), .B(A[982]), .Z(n170) );
  AND U150 ( .A(n171), .B(n172), .Z(n169) );
  NAND U151 ( .A(n173), .B(n174), .Z(n172) );
  NANDN U152 ( .A(A[981]), .B(B[981]), .Z(n174) );
  AND U153 ( .A(n175), .B(n176), .Z(n173) );
  NANDN U154 ( .A(A[980]), .B(B[980]), .Z(n176) );
  NAND U155 ( .A(n177), .B(n178), .Z(n175) );
  NANDN U156 ( .A(B[980]), .B(A[980]), .Z(n178) );
  AND U157 ( .A(n179), .B(n180), .Z(n177) );
  NAND U158 ( .A(n181), .B(n182), .Z(n180) );
  NANDN U159 ( .A(A[979]), .B(B[979]), .Z(n182) );
  AND U160 ( .A(n183), .B(n184), .Z(n181) );
  NANDN U161 ( .A(A[978]), .B(B[978]), .Z(n184) );
  NAND U162 ( .A(n185), .B(n186), .Z(n183) );
  NANDN U163 ( .A(B[978]), .B(A[978]), .Z(n186) );
  AND U164 ( .A(n187), .B(n188), .Z(n185) );
  NAND U165 ( .A(n189), .B(n190), .Z(n188) );
  NANDN U166 ( .A(A[977]), .B(B[977]), .Z(n190) );
  AND U167 ( .A(n191), .B(n192), .Z(n189) );
  NANDN U168 ( .A(A[976]), .B(B[976]), .Z(n192) );
  NAND U169 ( .A(n193), .B(n194), .Z(n191) );
  NANDN U170 ( .A(B[976]), .B(A[976]), .Z(n194) );
  AND U171 ( .A(n195), .B(n196), .Z(n193) );
  NAND U172 ( .A(n197), .B(n198), .Z(n196) );
  NANDN U173 ( .A(A[975]), .B(B[975]), .Z(n198) );
  AND U174 ( .A(n199), .B(n200), .Z(n197) );
  NANDN U175 ( .A(A[974]), .B(B[974]), .Z(n200) );
  NAND U176 ( .A(n201), .B(n202), .Z(n199) );
  NANDN U177 ( .A(B[974]), .B(A[974]), .Z(n202) );
  AND U178 ( .A(n203), .B(n204), .Z(n201) );
  NAND U179 ( .A(n205), .B(n206), .Z(n204) );
  NANDN U180 ( .A(A[973]), .B(B[973]), .Z(n206) );
  AND U181 ( .A(n207), .B(n208), .Z(n205) );
  NANDN U182 ( .A(A[972]), .B(B[972]), .Z(n208) );
  NAND U183 ( .A(n209), .B(n210), .Z(n207) );
  NANDN U184 ( .A(B[972]), .B(A[972]), .Z(n210) );
  AND U185 ( .A(n211), .B(n212), .Z(n209) );
  NAND U186 ( .A(n213), .B(n214), .Z(n212) );
  NANDN U187 ( .A(A[971]), .B(B[971]), .Z(n214) );
  AND U188 ( .A(n215), .B(n216), .Z(n213) );
  NANDN U189 ( .A(A[970]), .B(B[970]), .Z(n216) );
  NAND U190 ( .A(n217), .B(n218), .Z(n215) );
  NANDN U191 ( .A(B[970]), .B(A[970]), .Z(n218) );
  AND U192 ( .A(n219), .B(n220), .Z(n217) );
  NAND U193 ( .A(n221), .B(n222), .Z(n220) );
  NANDN U194 ( .A(A[969]), .B(B[969]), .Z(n222) );
  AND U195 ( .A(n223), .B(n224), .Z(n221) );
  NANDN U196 ( .A(A[968]), .B(B[968]), .Z(n224) );
  NAND U197 ( .A(n225), .B(n226), .Z(n223) );
  NANDN U198 ( .A(B[968]), .B(A[968]), .Z(n226) );
  AND U199 ( .A(n227), .B(n228), .Z(n225) );
  NAND U200 ( .A(n229), .B(n230), .Z(n228) );
  NANDN U201 ( .A(A[967]), .B(B[967]), .Z(n230) );
  AND U202 ( .A(n231), .B(n232), .Z(n229) );
  NANDN U203 ( .A(A[966]), .B(B[966]), .Z(n232) );
  NAND U204 ( .A(n233), .B(n234), .Z(n231) );
  NANDN U205 ( .A(B[966]), .B(A[966]), .Z(n234) );
  AND U206 ( .A(n235), .B(n236), .Z(n233) );
  NAND U207 ( .A(n237), .B(n238), .Z(n236) );
  NANDN U208 ( .A(A[965]), .B(B[965]), .Z(n238) );
  AND U209 ( .A(n239), .B(n240), .Z(n237) );
  NANDN U210 ( .A(A[964]), .B(B[964]), .Z(n240) );
  NAND U211 ( .A(n241), .B(n242), .Z(n239) );
  NANDN U212 ( .A(B[964]), .B(A[964]), .Z(n242) );
  AND U213 ( .A(n243), .B(n244), .Z(n241) );
  NAND U214 ( .A(n245), .B(n246), .Z(n244) );
  NANDN U215 ( .A(A[963]), .B(B[963]), .Z(n246) );
  AND U216 ( .A(n247), .B(n248), .Z(n245) );
  NANDN U217 ( .A(A[962]), .B(B[962]), .Z(n248) );
  NAND U218 ( .A(n249), .B(n250), .Z(n247) );
  NANDN U219 ( .A(B[962]), .B(A[962]), .Z(n250) );
  AND U220 ( .A(n251), .B(n252), .Z(n249) );
  NAND U221 ( .A(n253), .B(n254), .Z(n252) );
  NANDN U222 ( .A(A[961]), .B(B[961]), .Z(n254) );
  AND U223 ( .A(n255), .B(n256), .Z(n253) );
  NANDN U224 ( .A(A[960]), .B(B[960]), .Z(n256) );
  NAND U225 ( .A(n257), .B(n258), .Z(n255) );
  NANDN U226 ( .A(B[960]), .B(A[960]), .Z(n258) );
  AND U227 ( .A(n259), .B(n260), .Z(n257) );
  NAND U228 ( .A(n261), .B(n262), .Z(n260) );
  NANDN U229 ( .A(A[959]), .B(B[959]), .Z(n262) );
  AND U230 ( .A(n263), .B(n264), .Z(n261) );
  NANDN U231 ( .A(A[958]), .B(B[958]), .Z(n264) );
  NAND U232 ( .A(n265), .B(n266), .Z(n263) );
  NANDN U233 ( .A(B[958]), .B(A[958]), .Z(n266) );
  AND U234 ( .A(n267), .B(n268), .Z(n265) );
  NAND U235 ( .A(n269), .B(n270), .Z(n268) );
  NANDN U236 ( .A(A[957]), .B(B[957]), .Z(n270) );
  AND U237 ( .A(n271), .B(n272), .Z(n269) );
  NANDN U238 ( .A(A[956]), .B(B[956]), .Z(n272) );
  NAND U239 ( .A(n273), .B(n274), .Z(n271) );
  NANDN U240 ( .A(B[956]), .B(A[956]), .Z(n274) );
  AND U241 ( .A(n275), .B(n276), .Z(n273) );
  NAND U242 ( .A(n277), .B(n278), .Z(n276) );
  NANDN U243 ( .A(A[955]), .B(B[955]), .Z(n278) );
  AND U244 ( .A(n279), .B(n280), .Z(n277) );
  NANDN U245 ( .A(A[954]), .B(B[954]), .Z(n280) );
  NAND U246 ( .A(n281), .B(n282), .Z(n279) );
  NANDN U247 ( .A(B[954]), .B(A[954]), .Z(n282) );
  AND U248 ( .A(n283), .B(n284), .Z(n281) );
  NAND U249 ( .A(n285), .B(n286), .Z(n284) );
  NANDN U250 ( .A(A[953]), .B(B[953]), .Z(n286) );
  AND U251 ( .A(n287), .B(n288), .Z(n285) );
  NANDN U252 ( .A(A[952]), .B(B[952]), .Z(n288) );
  NAND U253 ( .A(n289), .B(n290), .Z(n287) );
  NANDN U254 ( .A(B[952]), .B(A[952]), .Z(n290) );
  AND U255 ( .A(n291), .B(n292), .Z(n289) );
  NAND U256 ( .A(n293), .B(n294), .Z(n292) );
  NANDN U257 ( .A(A[951]), .B(B[951]), .Z(n294) );
  AND U258 ( .A(n295), .B(n296), .Z(n293) );
  NANDN U259 ( .A(A[950]), .B(B[950]), .Z(n296) );
  NAND U260 ( .A(n297), .B(n298), .Z(n295) );
  NANDN U261 ( .A(B[950]), .B(A[950]), .Z(n298) );
  AND U262 ( .A(n299), .B(n300), .Z(n297) );
  NAND U263 ( .A(n301), .B(n302), .Z(n300) );
  NANDN U264 ( .A(A[949]), .B(B[949]), .Z(n302) );
  AND U265 ( .A(n303), .B(n304), .Z(n301) );
  NANDN U266 ( .A(A[948]), .B(B[948]), .Z(n304) );
  NAND U267 ( .A(n305), .B(n306), .Z(n303) );
  NANDN U268 ( .A(B[948]), .B(A[948]), .Z(n306) );
  AND U269 ( .A(n307), .B(n308), .Z(n305) );
  NAND U270 ( .A(n309), .B(n310), .Z(n308) );
  NANDN U271 ( .A(A[947]), .B(B[947]), .Z(n310) );
  AND U272 ( .A(n311), .B(n312), .Z(n309) );
  NANDN U273 ( .A(A[946]), .B(B[946]), .Z(n312) );
  NAND U274 ( .A(n313), .B(n314), .Z(n311) );
  NANDN U275 ( .A(B[946]), .B(A[946]), .Z(n314) );
  AND U276 ( .A(n315), .B(n316), .Z(n313) );
  NAND U277 ( .A(n317), .B(n318), .Z(n316) );
  NANDN U278 ( .A(A[945]), .B(B[945]), .Z(n318) );
  AND U279 ( .A(n319), .B(n320), .Z(n317) );
  NANDN U280 ( .A(A[944]), .B(B[944]), .Z(n320) );
  NAND U281 ( .A(n321), .B(n322), .Z(n319) );
  NANDN U282 ( .A(B[944]), .B(A[944]), .Z(n322) );
  AND U283 ( .A(n323), .B(n324), .Z(n321) );
  NAND U284 ( .A(n325), .B(n326), .Z(n324) );
  NANDN U285 ( .A(A[943]), .B(B[943]), .Z(n326) );
  AND U286 ( .A(n327), .B(n328), .Z(n325) );
  NANDN U287 ( .A(A[942]), .B(B[942]), .Z(n328) );
  NAND U288 ( .A(n329), .B(n330), .Z(n327) );
  NANDN U289 ( .A(B[942]), .B(A[942]), .Z(n330) );
  AND U290 ( .A(n331), .B(n332), .Z(n329) );
  NAND U291 ( .A(n333), .B(n334), .Z(n332) );
  NANDN U292 ( .A(A[941]), .B(B[941]), .Z(n334) );
  AND U293 ( .A(n335), .B(n336), .Z(n333) );
  NANDN U294 ( .A(A[940]), .B(B[940]), .Z(n336) );
  NAND U295 ( .A(n337), .B(n338), .Z(n335) );
  NANDN U296 ( .A(B[940]), .B(A[940]), .Z(n338) );
  AND U297 ( .A(n339), .B(n340), .Z(n337) );
  NAND U298 ( .A(n341), .B(n342), .Z(n340) );
  NANDN U299 ( .A(A[939]), .B(B[939]), .Z(n342) );
  AND U300 ( .A(n343), .B(n344), .Z(n341) );
  NANDN U301 ( .A(A[938]), .B(B[938]), .Z(n344) );
  NAND U302 ( .A(n345), .B(n346), .Z(n343) );
  NANDN U303 ( .A(B[938]), .B(A[938]), .Z(n346) );
  AND U304 ( .A(n347), .B(n348), .Z(n345) );
  NAND U305 ( .A(n349), .B(n350), .Z(n348) );
  NANDN U306 ( .A(A[937]), .B(B[937]), .Z(n350) );
  AND U307 ( .A(n351), .B(n352), .Z(n349) );
  NANDN U308 ( .A(A[936]), .B(B[936]), .Z(n352) );
  NAND U309 ( .A(n353), .B(n354), .Z(n351) );
  NANDN U310 ( .A(B[936]), .B(A[936]), .Z(n354) );
  AND U311 ( .A(n355), .B(n356), .Z(n353) );
  NAND U312 ( .A(n357), .B(n358), .Z(n356) );
  NANDN U313 ( .A(A[935]), .B(B[935]), .Z(n358) );
  AND U314 ( .A(n359), .B(n360), .Z(n357) );
  NANDN U315 ( .A(A[934]), .B(B[934]), .Z(n360) );
  NAND U316 ( .A(n361), .B(n362), .Z(n359) );
  NANDN U317 ( .A(B[934]), .B(A[934]), .Z(n362) );
  AND U318 ( .A(n363), .B(n364), .Z(n361) );
  NAND U319 ( .A(n365), .B(n366), .Z(n364) );
  NANDN U320 ( .A(A[933]), .B(B[933]), .Z(n366) );
  AND U321 ( .A(n367), .B(n368), .Z(n365) );
  NANDN U322 ( .A(A[932]), .B(B[932]), .Z(n368) );
  NAND U323 ( .A(n369), .B(n370), .Z(n367) );
  NANDN U324 ( .A(B[932]), .B(A[932]), .Z(n370) );
  AND U325 ( .A(n371), .B(n372), .Z(n369) );
  NAND U326 ( .A(n373), .B(n374), .Z(n372) );
  NANDN U327 ( .A(A[931]), .B(B[931]), .Z(n374) );
  AND U328 ( .A(n375), .B(n376), .Z(n373) );
  NANDN U329 ( .A(A[930]), .B(B[930]), .Z(n376) );
  NAND U330 ( .A(n377), .B(n378), .Z(n375) );
  NANDN U331 ( .A(B[930]), .B(A[930]), .Z(n378) );
  AND U332 ( .A(n379), .B(n380), .Z(n377) );
  NAND U333 ( .A(n381), .B(n382), .Z(n380) );
  NANDN U334 ( .A(A[929]), .B(B[929]), .Z(n382) );
  AND U335 ( .A(n383), .B(n384), .Z(n381) );
  NANDN U336 ( .A(A[928]), .B(B[928]), .Z(n384) );
  NAND U337 ( .A(n385), .B(n386), .Z(n383) );
  NANDN U338 ( .A(B[928]), .B(A[928]), .Z(n386) );
  AND U339 ( .A(n387), .B(n388), .Z(n385) );
  NAND U340 ( .A(n389), .B(n390), .Z(n388) );
  NANDN U341 ( .A(A[927]), .B(B[927]), .Z(n390) );
  AND U342 ( .A(n391), .B(n392), .Z(n389) );
  NANDN U343 ( .A(A[926]), .B(B[926]), .Z(n392) );
  NAND U344 ( .A(n393), .B(n394), .Z(n391) );
  NANDN U345 ( .A(B[926]), .B(A[926]), .Z(n394) );
  AND U346 ( .A(n395), .B(n396), .Z(n393) );
  NAND U347 ( .A(n397), .B(n398), .Z(n396) );
  NANDN U348 ( .A(A[925]), .B(B[925]), .Z(n398) );
  AND U349 ( .A(n399), .B(n400), .Z(n397) );
  NANDN U350 ( .A(A[924]), .B(B[924]), .Z(n400) );
  NAND U351 ( .A(n401), .B(n402), .Z(n399) );
  NANDN U352 ( .A(B[924]), .B(A[924]), .Z(n402) );
  AND U353 ( .A(n403), .B(n404), .Z(n401) );
  NAND U354 ( .A(n405), .B(n406), .Z(n404) );
  NANDN U355 ( .A(A[923]), .B(B[923]), .Z(n406) );
  AND U356 ( .A(n407), .B(n408), .Z(n405) );
  NANDN U357 ( .A(A[922]), .B(B[922]), .Z(n408) );
  NAND U358 ( .A(n409), .B(n410), .Z(n407) );
  NANDN U359 ( .A(B[922]), .B(A[922]), .Z(n410) );
  AND U360 ( .A(n411), .B(n412), .Z(n409) );
  NAND U361 ( .A(n413), .B(n414), .Z(n412) );
  NANDN U362 ( .A(A[921]), .B(B[921]), .Z(n414) );
  AND U363 ( .A(n415), .B(n416), .Z(n413) );
  NANDN U364 ( .A(A[920]), .B(B[920]), .Z(n416) );
  NAND U365 ( .A(n417), .B(n418), .Z(n415) );
  NANDN U366 ( .A(B[920]), .B(A[920]), .Z(n418) );
  AND U367 ( .A(n419), .B(n420), .Z(n417) );
  NAND U368 ( .A(n421), .B(n422), .Z(n420) );
  NANDN U369 ( .A(A[919]), .B(B[919]), .Z(n422) );
  AND U370 ( .A(n423), .B(n424), .Z(n421) );
  NANDN U371 ( .A(A[918]), .B(B[918]), .Z(n424) );
  NAND U372 ( .A(n425), .B(n426), .Z(n423) );
  NANDN U373 ( .A(B[918]), .B(A[918]), .Z(n426) );
  AND U374 ( .A(n427), .B(n428), .Z(n425) );
  NAND U375 ( .A(n429), .B(n430), .Z(n428) );
  NANDN U376 ( .A(A[917]), .B(B[917]), .Z(n430) );
  AND U377 ( .A(n431), .B(n432), .Z(n429) );
  NANDN U378 ( .A(A[916]), .B(B[916]), .Z(n432) );
  NAND U379 ( .A(n433), .B(n434), .Z(n431) );
  NANDN U380 ( .A(B[916]), .B(A[916]), .Z(n434) );
  AND U381 ( .A(n435), .B(n436), .Z(n433) );
  NAND U382 ( .A(n437), .B(n438), .Z(n436) );
  NANDN U383 ( .A(A[915]), .B(B[915]), .Z(n438) );
  AND U384 ( .A(n439), .B(n440), .Z(n437) );
  NANDN U385 ( .A(A[914]), .B(B[914]), .Z(n440) );
  NAND U386 ( .A(n441), .B(n442), .Z(n439) );
  NANDN U387 ( .A(B[914]), .B(A[914]), .Z(n442) );
  AND U388 ( .A(n443), .B(n444), .Z(n441) );
  NAND U389 ( .A(n445), .B(n446), .Z(n444) );
  NANDN U390 ( .A(A[913]), .B(B[913]), .Z(n446) );
  AND U391 ( .A(n447), .B(n448), .Z(n445) );
  NANDN U392 ( .A(A[912]), .B(B[912]), .Z(n448) );
  NAND U393 ( .A(n449), .B(n450), .Z(n447) );
  NANDN U394 ( .A(B[912]), .B(A[912]), .Z(n450) );
  AND U395 ( .A(n451), .B(n452), .Z(n449) );
  NAND U396 ( .A(n453), .B(n454), .Z(n452) );
  NANDN U397 ( .A(A[911]), .B(B[911]), .Z(n454) );
  AND U398 ( .A(n455), .B(n456), .Z(n453) );
  NANDN U399 ( .A(A[910]), .B(B[910]), .Z(n456) );
  NAND U400 ( .A(n457), .B(n458), .Z(n455) );
  NANDN U401 ( .A(B[910]), .B(A[910]), .Z(n458) );
  AND U402 ( .A(n459), .B(n460), .Z(n457) );
  NAND U403 ( .A(n461), .B(n462), .Z(n460) );
  NANDN U404 ( .A(A[909]), .B(B[909]), .Z(n462) );
  AND U405 ( .A(n463), .B(n464), .Z(n461) );
  NANDN U406 ( .A(A[908]), .B(B[908]), .Z(n464) );
  NAND U407 ( .A(n465), .B(n466), .Z(n463) );
  NANDN U408 ( .A(B[908]), .B(A[908]), .Z(n466) );
  AND U409 ( .A(n467), .B(n468), .Z(n465) );
  NAND U410 ( .A(n469), .B(n470), .Z(n468) );
  NANDN U411 ( .A(A[907]), .B(B[907]), .Z(n470) );
  AND U412 ( .A(n471), .B(n472), .Z(n469) );
  NANDN U413 ( .A(A[906]), .B(B[906]), .Z(n472) );
  NAND U414 ( .A(n473), .B(n474), .Z(n471) );
  NANDN U415 ( .A(B[906]), .B(A[906]), .Z(n474) );
  AND U416 ( .A(n475), .B(n476), .Z(n473) );
  NAND U417 ( .A(n477), .B(n478), .Z(n476) );
  NANDN U418 ( .A(A[905]), .B(B[905]), .Z(n478) );
  AND U419 ( .A(n479), .B(n480), .Z(n477) );
  NANDN U420 ( .A(A[904]), .B(B[904]), .Z(n480) );
  NAND U421 ( .A(n481), .B(n482), .Z(n479) );
  NANDN U422 ( .A(B[904]), .B(A[904]), .Z(n482) );
  AND U423 ( .A(n483), .B(n484), .Z(n481) );
  NAND U424 ( .A(n485), .B(n486), .Z(n484) );
  NANDN U425 ( .A(A[903]), .B(B[903]), .Z(n486) );
  AND U426 ( .A(n487), .B(n488), .Z(n485) );
  NANDN U427 ( .A(A[902]), .B(B[902]), .Z(n488) );
  NAND U428 ( .A(n489), .B(n490), .Z(n487) );
  NANDN U429 ( .A(B[902]), .B(A[902]), .Z(n490) );
  AND U430 ( .A(n491), .B(n492), .Z(n489) );
  NAND U431 ( .A(n493), .B(n494), .Z(n492) );
  NANDN U432 ( .A(A[901]), .B(B[901]), .Z(n494) );
  AND U433 ( .A(n495), .B(n496), .Z(n493) );
  NANDN U434 ( .A(A[900]), .B(B[900]), .Z(n496) );
  NAND U435 ( .A(n497), .B(n498), .Z(n495) );
  NANDN U436 ( .A(B[900]), .B(A[900]), .Z(n498) );
  AND U437 ( .A(n499), .B(n500), .Z(n497) );
  NAND U438 ( .A(n501), .B(n502), .Z(n500) );
  NANDN U439 ( .A(A[899]), .B(B[899]), .Z(n502) );
  AND U440 ( .A(n503), .B(n504), .Z(n501) );
  NANDN U441 ( .A(A[898]), .B(B[898]), .Z(n504) );
  NAND U442 ( .A(n505), .B(n506), .Z(n503) );
  NANDN U443 ( .A(B[898]), .B(A[898]), .Z(n506) );
  AND U444 ( .A(n507), .B(n508), .Z(n505) );
  NAND U445 ( .A(n509), .B(n510), .Z(n508) );
  NANDN U446 ( .A(A[897]), .B(B[897]), .Z(n510) );
  AND U447 ( .A(n511), .B(n512), .Z(n509) );
  NANDN U448 ( .A(A[896]), .B(B[896]), .Z(n512) );
  NAND U449 ( .A(n513), .B(n514), .Z(n511) );
  NANDN U450 ( .A(B[896]), .B(A[896]), .Z(n514) );
  AND U451 ( .A(n515), .B(n516), .Z(n513) );
  NAND U452 ( .A(n517), .B(n518), .Z(n516) );
  NANDN U453 ( .A(A[895]), .B(B[895]), .Z(n518) );
  AND U454 ( .A(n519), .B(n520), .Z(n517) );
  NANDN U455 ( .A(A[894]), .B(B[894]), .Z(n520) );
  NAND U456 ( .A(n521), .B(n522), .Z(n519) );
  NANDN U457 ( .A(B[894]), .B(A[894]), .Z(n522) );
  AND U458 ( .A(n523), .B(n524), .Z(n521) );
  NAND U459 ( .A(n525), .B(n526), .Z(n524) );
  NANDN U460 ( .A(A[893]), .B(B[893]), .Z(n526) );
  AND U461 ( .A(n527), .B(n528), .Z(n525) );
  NANDN U462 ( .A(A[892]), .B(B[892]), .Z(n528) );
  NAND U463 ( .A(n529), .B(n530), .Z(n527) );
  NANDN U464 ( .A(B[892]), .B(A[892]), .Z(n530) );
  AND U465 ( .A(n531), .B(n532), .Z(n529) );
  NAND U466 ( .A(n533), .B(n534), .Z(n532) );
  NANDN U467 ( .A(A[891]), .B(B[891]), .Z(n534) );
  AND U468 ( .A(n535), .B(n536), .Z(n533) );
  NANDN U469 ( .A(A[890]), .B(B[890]), .Z(n536) );
  NAND U470 ( .A(n537), .B(n538), .Z(n535) );
  NANDN U471 ( .A(B[890]), .B(A[890]), .Z(n538) );
  AND U472 ( .A(n539), .B(n540), .Z(n537) );
  NAND U473 ( .A(n541), .B(n542), .Z(n540) );
  NANDN U474 ( .A(A[889]), .B(B[889]), .Z(n542) );
  AND U475 ( .A(n543), .B(n544), .Z(n541) );
  NANDN U476 ( .A(A[888]), .B(B[888]), .Z(n544) );
  NAND U477 ( .A(n545), .B(n546), .Z(n543) );
  NANDN U478 ( .A(B[888]), .B(A[888]), .Z(n546) );
  AND U479 ( .A(n547), .B(n548), .Z(n545) );
  NAND U480 ( .A(n549), .B(n550), .Z(n548) );
  NANDN U481 ( .A(A[887]), .B(B[887]), .Z(n550) );
  AND U482 ( .A(n551), .B(n552), .Z(n549) );
  NANDN U483 ( .A(A[886]), .B(B[886]), .Z(n552) );
  NAND U484 ( .A(n553), .B(n554), .Z(n551) );
  NANDN U485 ( .A(B[886]), .B(A[886]), .Z(n554) );
  AND U486 ( .A(n555), .B(n556), .Z(n553) );
  NAND U487 ( .A(n557), .B(n558), .Z(n556) );
  NANDN U488 ( .A(A[885]), .B(B[885]), .Z(n558) );
  AND U489 ( .A(n559), .B(n560), .Z(n557) );
  NANDN U490 ( .A(A[884]), .B(B[884]), .Z(n560) );
  NAND U491 ( .A(n561), .B(n562), .Z(n559) );
  NANDN U492 ( .A(B[884]), .B(A[884]), .Z(n562) );
  AND U493 ( .A(n563), .B(n564), .Z(n561) );
  NAND U494 ( .A(n565), .B(n566), .Z(n564) );
  NANDN U495 ( .A(A[883]), .B(B[883]), .Z(n566) );
  AND U496 ( .A(n567), .B(n568), .Z(n565) );
  NANDN U497 ( .A(A[882]), .B(B[882]), .Z(n568) );
  NAND U498 ( .A(n569), .B(n570), .Z(n567) );
  NANDN U499 ( .A(B[882]), .B(A[882]), .Z(n570) );
  AND U500 ( .A(n571), .B(n572), .Z(n569) );
  NAND U501 ( .A(n573), .B(n574), .Z(n572) );
  NANDN U502 ( .A(A[881]), .B(B[881]), .Z(n574) );
  AND U503 ( .A(n575), .B(n576), .Z(n573) );
  NANDN U504 ( .A(A[880]), .B(B[880]), .Z(n576) );
  NAND U505 ( .A(n577), .B(n578), .Z(n575) );
  NANDN U506 ( .A(B[880]), .B(A[880]), .Z(n578) );
  AND U507 ( .A(n579), .B(n580), .Z(n577) );
  NAND U508 ( .A(n581), .B(n582), .Z(n580) );
  NANDN U509 ( .A(A[879]), .B(B[879]), .Z(n582) );
  AND U510 ( .A(n583), .B(n584), .Z(n581) );
  NANDN U511 ( .A(A[878]), .B(B[878]), .Z(n584) );
  NAND U512 ( .A(n585), .B(n586), .Z(n583) );
  NANDN U513 ( .A(B[878]), .B(A[878]), .Z(n586) );
  AND U514 ( .A(n587), .B(n588), .Z(n585) );
  NAND U515 ( .A(n589), .B(n590), .Z(n588) );
  NANDN U516 ( .A(A[877]), .B(B[877]), .Z(n590) );
  AND U517 ( .A(n591), .B(n592), .Z(n589) );
  NANDN U518 ( .A(A[876]), .B(B[876]), .Z(n592) );
  NAND U519 ( .A(n593), .B(n594), .Z(n591) );
  NANDN U520 ( .A(B[876]), .B(A[876]), .Z(n594) );
  AND U521 ( .A(n595), .B(n596), .Z(n593) );
  NAND U522 ( .A(n597), .B(n598), .Z(n596) );
  NANDN U523 ( .A(A[875]), .B(B[875]), .Z(n598) );
  AND U524 ( .A(n599), .B(n600), .Z(n597) );
  NANDN U525 ( .A(A[874]), .B(B[874]), .Z(n600) );
  NAND U526 ( .A(n601), .B(n602), .Z(n599) );
  NANDN U527 ( .A(B[874]), .B(A[874]), .Z(n602) );
  AND U528 ( .A(n603), .B(n604), .Z(n601) );
  NAND U529 ( .A(n605), .B(n606), .Z(n604) );
  NANDN U530 ( .A(A[873]), .B(B[873]), .Z(n606) );
  AND U531 ( .A(n607), .B(n608), .Z(n605) );
  NANDN U532 ( .A(A[872]), .B(B[872]), .Z(n608) );
  NAND U533 ( .A(n609), .B(n610), .Z(n607) );
  NANDN U534 ( .A(B[872]), .B(A[872]), .Z(n610) );
  AND U535 ( .A(n611), .B(n612), .Z(n609) );
  NAND U536 ( .A(n613), .B(n614), .Z(n612) );
  NANDN U537 ( .A(A[871]), .B(B[871]), .Z(n614) );
  AND U538 ( .A(n615), .B(n616), .Z(n613) );
  NANDN U539 ( .A(A[870]), .B(B[870]), .Z(n616) );
  NAND U540 ( .A(n617), .B(n618), .Z(n615) );
  NANDN U541 ( .A(B[870]), .B(A[870]), .Z(n618) );
  AND U542 ( .A(n619), .B(n620), .Z(n617) );
  NAND U543 ( .A(n621), .B(n622), .Z(n620) );
  NANDN U544 ( .A(A[869]), .B(B[869]), .Z(n622) );
  AND U545 ( .A(n623), .B(n624), .Z(n621) );
  NANDN U546 ( .A(A[868]), .B(B[868]), .Z(n624) );
  NAND U547 ( .A(n625), .B(n626), .Z(n623) );
  NANDN U548 ( .A(B[868]), .B(A[868]), .Z(n626) );
  AND U549 ( .A(n627), .B(n628), .Z(n625) );
  NAND U550 ( .A(n629), .B(n630), .Z(n628) );
  NANDN U551 ( .A(A[867]), .B(B[867]), .Z(n630) );
  AND U552 ( .A(n631), .B(n632), .Z(n629) );
  NANDN U553 ( .A(A[866]), .B(B[866]), .Z(n632) );
  NAND U554 ( .A(n633), .B(n634), .Z(n631) );
  NANDN U555 ( .A(B[866]), .B(A[866]), .Z(n634) );
  AND U556 ( .A(n635), .B(n636), .Z(n633) );
  NAND U557 ( .A(n637), .B(n638), .Z(n636) );
  NANDN U558 ( .A(A[865]), .B(B[865]), .Z(n638) );
  AND U559 ( .A(n639), .B(n640), .Z(n637) );
  NANDN U560 ( .A(A[864]), .B(B[864]), .Z(n640) );
  NAND U561 ( .A(n641), .B(n642), .Z(n639) );
  NANDN U562 ( .A(B[864]), .B(A[864]), .Z(n642) );
  AND U563 ( .A(n643), .B(n644), .Z(n641) );
  NAND U564 ( .A(n645), .B(n646), .Z(n644) );
  NANDN U565 ( .A(A[863]), .B(B[863]), .Z(n646) );
  AND U566 ( .A(n647), .B(n648), .Z(n645) );
  NANDN U567 ( .A(A[862]), .B(B[862]), .Z(n648) );
  NAND U568 ( .A(n649), .B(n650), .Z(n647) );
  NANDN U569 ( .A(B[862]), .B(A[862]), .Z(n650) );
  AND U570 ( .A(n651), .B(n652), .Z(n649) );
  NAND U571 ( .A(n653), .B(n654), .Z(n652) );
  NANDN U572 ( .A(A[861]), .B(B[861]), .Z(n654) );
  AND U573 ( .A(n655), .B(n656), .Z(n653) );
  NANDN U574 ( .A(A[860]), .B(B[860]), .Z(n656) );
  NAND U575 ( .A(n657), .B(n658), .Z(n655) );
  NANDN U576 ( .A(B[860]), .B(A[860]), .Z(n658) );
  AND U577 ( .A(n659), .B(n660), .Z(n657) );
  NAND U578 ( .A(n661), .B(n662), .Z(n660) );
  NANDN U579 ( .A(A[859]), .B(B[859]), .Z(n662) );
  AND U580 ( .A(n663), .B(n664), .Z(n661) );
  NANDN U581 ( .A(A[858]), .B(B[858]), .Z(n664) );
  NAND U582 ( .A(n665), .B(n666), .Z(n663) );
  NANDN U583 ( .A(B[858]), .B(A[858]), .Z(n666) );
  AND U584 ( .A(n667), .B(n668), .Z(n665) );
  NAND U585 ( .A(n669), .B(n670), .Z(n668) );
  NANDN U586 ( .A(A[857]), .B(B[857]), .Z(n670) );
  AND U587 ( .A(n671), .B(n672), .Z(n669) );
  NANDN U588 ( .A(A[856]), .B(B[856]), .Z(n672) );
  NAND U589 ( .A(n673), .B(n674), .Z(n671) );
  NANDN U590 ( .A(B[856]), .B(A[856]), .Z(n674) );
  AND U591 ( .A(n675), .B(n676), .Z(n673) );
  NAND U592 ( .A(n677), .B(n678), .Z(n676) );
  NANDN U593 ( .A(A[855]), .B(B[855]), .Z(n678) );
  AND U594 ( .A(n679), .B(n680), .Z(n677) );
  NANDN U595 ( .A(A[854]), .B(B[854]), .Z(n680) );
  NAND U596 ( .A(n681), .B(n682), .Z(n679) );
  NANDN U597 ( .A(B[854]), .B(A[854]), .Z(n682) );
  AND U598 ( .A(n683), .B(n684), .Z(n681) );
  NAND U599 ( .A(n685), .B(n686), .Z(n684) );
  NANDN U600 ( .A(A[853]), .B(B[853]), .Z(n686) );
  AND U601 ( .A(n687), .B(n688), .Z(n685) );
  NANDN U602 ( .A(A[852]), .B(B[852]), .Z(n688) );
  NAND U603 ( .A(n689), .B(n690), .Z(n687) );
  NANDN U604 ( .A(B[852]), .B(A[852]), .Z(n690) );
  AND U605 ( .A(n691), .B(n692), .Z(n689) );
  NAND U606 ( .A(n693), .B(n694), .Z(n692) );
  NANDN U607 ( .A(A[851]), .B(B[851]), .Z(n694) );
  AND U608 ( .A(n695), .B(n696), .Z(n693) );
  NANDN U609 ( .A(A[850]), .B(B[850]), .Z(n696) );
  NAND U610 ( .A(n697), .B(n698), .Z(n695) );
  NANDN U611 ( .A(B[850]), .B(A[850]), .Z(n698) );
  AND U612 ( .A(n699), .B(n700), .Z(n697) );
  NAND U613 ( .A(n701), .B(n702), .Z(n700) );
  NANDN U614 ( .A(A[849]), .B(B[849]), .Z(n702) );
  AND U615 ( .A(n703), .B(n704), .Z(n701) );
  NANDN U616 ( .A(A[848]), .B(B[848]), .Z(n704) );
  NAND U617 ( .A(n705), .B(n706), .Z(n703) );
  NANDN U618 ( .A(B[848]), .B(A[848]), .Z(n706) );
  AND U619 ( .A(n707), .B(n708), .Z(n705) );
  NAND U620 ( .A(n709), .B(n710), .Z(n708) );
  NANDN U621 ( .A(A[847]), .B(B[847]), .Z(n710) );
  AND U622 ( .A(n711), .B(n712), .Z(n709) );
  NANDN U623 ( .A(A[846]), .B(B[846]), .Z(n712) );
  NAND U624 ( .A(n713), .B(n714), .Z(n711) );
  NANDN U625 ( .A(B[846]), .B(A[846]), .Z(n714) );
  AND U626 ( .A(n715), .B(n716), .Z(n713) );
  NAND U627 ( .A(n717), .B(n718), .Z(n716) );
  NANDN U628 ( .A(A[845]), .B(B[845]), .Z(n718) );
  AND U629 ( .A(n719), .B(n720), .Z(n717) );
  NANDN U630 ( .A(A[844]), .B(B[844]), .Z(n720) );
  NAND U631 ( .A(n721), .B(n722), .Z(n719) );
  NANDN U632 ( .A(B[844]), .B(A[844]), .Z(n722) );
  AND U633 ( .A(n723), .B(n724), .Z(n721) );
  NAND U634 ( .A(n725), .B(n726), .Z(n724) );
  NANDN U635 ( .A(A[843]), .B(B[843]), .Z(n726) );
  AND U636 ( .A(n727), .B(n728), .Z(n725) );
  NANDN U637 ( .A(A[842]), .B(B[842]), .Z(n728) );
  NAND U638 ( .A(n729), .B(n730), .Z(n727) );
  NANDN U639 ( .A(B[842]), .B(A[842]), .Z(n730) );
  AND U640 ( .A(n731), .B(n732), .Z(n729) );
  NAND U641 ( .A(n733), .B(n734), .Z(n732) );
  NANDN U642 ( .A(A[841]), .B(B[841]), .Z(n734) );
  AND U643 ( .A(n735), .B(n736), .Z(n733) );
  NANDN U644 ( .A(A[840]), .B(B[840]), .Z(n736) );
  NAND U645 ( .A(n737), .B(n738), .Z(n735) );
  NANDN U646 ( .A(B[840]), .B(A[840]), .Z(n738) );
  AND U647 ( .A(n739), .B(n740), .Z(n737) );
  NAND U648 ( .A(n741), .B(n742), .Z(n740) );
  NANDN U649 ( .A(A[839]), .B(B[839]), .Z(n742) );
  AND U650 ( .A(n743), .B(n744), .Z(n741) );
  NANDN U651 ( .A(A[838]), .B(B[838]), .Z(n744) );
  NAND U652 ( .A(n745), .B(n746), .Z(n743) );
  NANDN U653 ( .A(B[838]), .B(A[838]), .Z(n746) );
  AND U654 ( .A(n747), .B(n748), .Z(n745) );
  NAND U655 ( .A(n749), .B(n750), .Z(n748) );
  NANDN U656 ( .A(A[837]), .B(B[837]), .Z(n750) );
  AND U657 ( .A(n751), .B(n752), .Z(n749) );
  NANDN U658 ( .A(A[836]), .B(B[836]), .Z(n752) );
  NAND U659 ( .A(n753), .B(n754), .Z(n751) );
  NANDN U660 ( .A(B[836]), .B(A[836]), .Z(n754) );
  AND U661 ( .A(n755), .B(n756), .Z(n753) );
  NAND U662 ( .A(n757), .B(n758), .Z(n756) );
  NANDN U663 ( .A(A[835]), .B(B[835]), .Z(n758) );
  AND U664 ( .A(n759), .B(n760), .Z(n757) );
  NANDN U665 ( .A(A[834]), .B(B[834]), .Z(n760) );
  NAND U666 ( .A(n761), .B(n762), .Z(n759) );
  NANDN U667 ( .A(B[834]), .B(A[834]), .Z(n762) );
  AND U668 ( .A(n763), .B(n764), .Z(n761) );
  NAND U669 ( .A(n765), .B(n766), .Z(n764) );
  NANDN U670 ( .A(A[833]), .B(B[833]), .Z(n766) );
  AND U671 ( .A(n767), .B(n768), .Z(n765) );
  NANDN U672 ( .A(A[832]), .B(B[832]), .Z(n768) );
  NAND U673 ( .A(n769), .B(n770), .Z(n767) );
  NANDN U674 ( .A(B[832]), .B(A[832]), .Z(n770) );
  AND U675 ( .A(n771), .B(n772), .Z(n769) );
  NAND U676 ( .A(n773), .B(n774), .Z(n772) );
  NANDN U677 ( .A(A[831]), .B(B[831]), .Z(n774) );
  AND U678 ( .A(n775), .B(n776), .Z(n773) );
  NANDN U679 ( .A(A[830]), .B(B[830]), .Z(n776) );
  NAND U680 ( .A(n777), .B(n778), .Z(n775) );
  NANDN U681 ( .A(B[830]), .B(A[830]), .Z(n778) );
  AND U682 ( .A(n779), .B(n780), .Z(n777) );
  NAND U683 ( .A(n781), .B(n782), .Z(n780) );
  NANDN U684 ( .A(A[829]), .B(B[829]), .Z(n782) );
  AND U685 ( .A(n783), .B(n784), .Z(n781) );
  NANDN U686 ( .A(A[828]), .B(B[828]), .Z(n784) );
  NAND U687 ( .A(n785), .B(n786), .Z(n783) );
  NANDN U688 ( .A(B[828]), .B(A[828]), .Z(n786) );
  AND U689 ( .A(n787), .B(n788), .Z(n785) );
  NAND U690 ( .A(n789), .B(n790), .Z(n788) );
  NANDN U691 ( .A(A[827]), .B(B[827]), .Z(n790) );
  AND U692 ( .A(n791), .B(n792), .Z(n789) );
  NANDN U693 ( .A(A[826]), .B(B[826]), .Z(n792) );
  NAND U694 ( .A(n793), .B(n794), .Z(n791) );
  NANDN U695 ( .A(B[826]), .B(A[826]), .Z(n794) );
  AND U696 ( .A(n795), .B(n796), .Z(n793) );
  NAND U697 ( .A(n797), .B(n798), .Z(n796) );
  NANDN U698 ( .A(A[825]), .B(B[825]), .Z(n798) );
  AND U699 ( .A(n799), .B(n800), .Z(n797) );
  NANDN U700 ( .A(A[824]), .B(B[824]), .Z(n800) );
  NAND U701 ( .A(n801), .B(n802), .Z(n799) );
  NANDN U702 ( .A(B[824]), .B(A[824]), .Z(n802) );
  AND U703 ( .A(n803), .B(n804), .Z(n801) );
  NAND U704 ( .A(n805), .B(n806), .Z(n804) );
  NANDN U705 ( .A(A[823]), .B(B[823]), .Z(n806) );
  AND U706 ( .A(n807), .B(n808), .Z(n805) );
  NANDN U707 ( .A(A[822]), .B(B[822]), .Z(n808) );
  NAND U708 ( .A(n809), .B(n810), .Z(n807) );
  NANDN U709 ( .A(B[822]), .B(A[822]), .Z(n810) );
  AND U710 ( .A(n811), .B(n812), .Z(n809) );
  NAND U711 ( .A(n813), .B(n814), .Z(n812) );
  NANDN U712 ( .A(A[821]), .B(B[821]), .Z(n814) );
  AND U713 ( .A(n815), .B(n816), .Z(n813) );
  NANDN U714 ( .A(A[820]), .B(B[820]), .Z(n816) );
  NAND U715 ( .A(n817), .B(n818), .Z(n815) );
  NANDN U716 ( .A(B[820]), .B(A[820]), .Z(n818) );
  AND U717 ( .A(n819), .B(n820), .Z(n817) );
  NAND U718 ( .A(n821), .B(n822), .Z(n820) );
  NANDN U719 ( .A(A[819]), .B(B[819]), .Z(n822) );
  AND U720 ( .A(n823), .B(n824), .Z(n821) );
  NANDN U721 ( .A(A[818]), .B(B[818]), .Z(n824) );
  NAND U722 ( .A(n825), .B(n826), .Z(n823) );
  NANDN U723 ( .A(B[818]), .B(A[818]), .Z(n826) );
  AND U724 ( .A(n827), .B(n828), .Z(n825) );
  NAND U725 ( .A(n829), .B(n830), .Z(n828) );
  NANDN U726 ( .A(A[817]), .B(B[817]), .Z(n830) );
  AND U727 ( .A(n831), .B(n832), .Z(n829) );
  NANDN U728 ( .A(A[816]), .B(B[816]), .Z(n832) );
  NAND U729 ( .A(n833), .B(n834), .Z(n831) );
  NANDN U730 ( .A(B[816]), .B(A[816]), .Z(n834) );
  AND U731 ( .A(n835), .B(n836), .Z(n833) );
  NAND U732 ( .A(n837), .B(n838), .Z(n836) );
  NANDN U733 ( .A(A[815]), .B(B[815]), .Z(n838) );
  AND U734 ( .A(n839), .B(n840), .Z(n837) );
  NANDN U735 ( .A(A[814]), .B(B[814]), .Z(n840) );
  NAND U736 ( .A(n841), .B(n842), .Z(n839) );
  NANDN U737 ( .A(B[814]), .B(A[814]), .Z(n842) );
  AND U738 ( .A(n843), .B(n844), .Z(n841) );
  NAND U739 ( .A(n845), .B(n846), .Z(n844) );
  NANDN U740 ( .A(A[813]), .B(B[813]), .Z(n846) );
  AND U741 ( .A(n847), .B(n848), .Z(n845) );
  NANDN U742 ( .A(A[812]), .B(B[812]), .Z(n848) );
  NAND U743 ( .A(n849), .B(n850), .Z(n847) );
  NANDN U744 ( .A(B[812]), .B(A[812]), .Z(n850) );
  AND U745 ( .A(n851), .B(n852), .Z(n849) );
  NAND U746 ( .A(n853), .B(n854), .Z(n852) );
  NANDN U747 ( .A(A[811]), .B(B[811]), .Z(n854) );
  AND U748 ( .A(n855), .B(n856), .Z(n853) );
  NANDN U749 ( .A(A[810]), .B(B[810]), .Z(n856) );
  NAND U750 ( .A(n857), .B(n858), .Z(n855) );
  NANDN U751 ( .A(B[810]), .B(A[810]), .Z(n858) );
  AND U752 ( .A(n859), .B(n860), .Z(n857) );
  NAND U753 ( .A(n861), .B(n862), .Z(n860) );
  NANDN U754 ( .A(A[809]), .B(B[809]), .Z(n862) );
  AND U755 ( .A(n863), .B(n864), .Z(n861) );
  NANDN U756 ( .A(A[808]), .B(B[808]), .Z(n864) );
  NAND U757 ( .A(n865), .B(n866), .Z(n863) );
  NANDN U758 ( .A(B[808]), .B(A[808]), .Z(n866) );
  AND U759 ( .A(n867), .B(n868), .Z(n865) );
  NAND U760 ( .A(n869), .B(n870), .Z(n868) );
  NANDN U761 ( .A(A[807]), .B(B[807]), .Z(n870) );
  AND U762 ( .A(n871), .B(n872), .Z(n869) );
  NANDN U763 ( .A(A[806]), .B(B[806]), .Z(n872) );
  NAND U764 ( .A(n873), .B(n874), .Z(n871) );
  NANDN U765 ( .A(B[806]), .B(A[806]), .Z(n874) );
  AND U766 ( .A(n875), .B(n876), .Z(n873) );
  NAND U767 ( .A(n877), .B(n878), .Z(n876) );
  NANDN U768 ( .A(A[805]), .B(B[805]), .Z(n878) );
  AND U769 ( .A(n879), .B(n880), .Z(n877) );
  NANDN U770 ( .A(A[804]), .B(B[804]), .Z(n880) );
  NAND U771 ( .A(n881), .B(n882), .Z(n879) );
  NANDN U772 ( .A(B[804]), .B(A[804]), .Z(n882) );
  AND U773 ( .A(n883), .B(n884), .Z(n881) );
  NAND U774 ( .A(n885), .B(n886), .Z(n884) );
  NANDN U775 ( .A(A[803]), .B(B[803]), .Z(n886) );
  AND U776 ( .A(n887), .B(n888), .Z(n885) );
  NANDN U777 ( .A(A[802]), .B(B[802]), .Z(n888) );
  NAND U778 ( .A(n889), .B(n890), .Z(n887) );
  NANDN U779 ( .A(B[802]), .B(A[802]), .Z(n890) );
  AND U780 ( .A(n891), .B(n892), .Z(n889) );
  NAND U781 ( .A(n893), .B(n894), .Z(n892) );
  NANDN U782 ( .A(A[801]), .B(B[801]), .Z(n894) );
  AND U783 ( .A(n895), .B(n896), .Z(n893) );
  NANDN U784 ( .A(A[800]), .B(B[800]), .Z(n896) );
  NAND U785 ( .A(n897), .B(n898), .Z(n895) );
  NANDN U786 ( .A(B[800]), .B(A[800]), .Z(n898) );
  AND U787 ( .A(n899), .B(n900), .Z(n897) );
  NAND U788 ( .A(n901), .B(n902), .Z(n900) );
  NANDN U789 ( .A(A[799]), .B(B[799]), .Z(n902) );
  AND U790 ( .A(n903), .B(n904), .Z(n901) );
  NANDN U791 ( .A(A[798]), .B(B[798]), .Z(n904) );
  NAND U792 ( .A(n905), .B(n906), .Z(n903) );
  NANDN U793 ( .A(B[798]), .B(A[798]), .Z(n906) );
  AND U794 ( .A(n907), .B(n908), .Z(n905) );
  NAND U795 ( .A(n909), .B(n910), .Z(n908) );
  NANDN U796 ( .A(A[797]), .B(B[797]), .Z(n910) );
  AND U797 ( .A(n911), .B(n912), .Z(n909) );
  NANDN U798 ( .A(A[796]), .B(B[796]), .Z(n912) );
  NAND U799 ( .A(n913), .B(n914), .Z(n911) );
  NANDN U800 ( .A(B[796]), .B(A[796]), .Z(n914) );
  AND U801 ( .A(n915), .B(n916), .Z(n913) );
  NAND U802 ( .A(n917), .B(n918), .Z(n916) );
  NANDN U803 ( .A(A[795]), .B(B[795]), .Z(n918) );
  AND U804 ( .A(n919), .B(n920), .Z(n917) );
  NANDN U805 ( .A(A[794]), .B(B[794]), .Z(n920) );
  NAND U806 ( .A(n921), .B(n922), .Z(n919) );
  NANDN U807 ( .A(B[794]), .B(A[794]), .Z(n922) );
  AND U808 ( .A(n923), .B(n924), .Z(n921) );
  NAND U809 ( .A(n925), .B(n926), .Z(n924) );
  NANDN U810 ( .A(A[793]), .B(B[793]), .Z(n926) );
  AND U811 ( .A(n927), .B(n928), .Z(n925) );
  NANDN U812 ( .A(A[792]), .B(B[792]), .Z(n928) );
  NAND U813 ( .A(n929), .B(n930), .Z(n927) );
  NANDN U814 ( .A(B[792]), .B(A[792]), .Z(n930) );
  AND U815 ( .A(n931), .B(n932), .Z(n929) );
  NAND U816 ( .A(n933), .B(n934), .Z(n932) );
  NANDN U817 ( .A(A[791]), .B(B[791]), .Z(n934) );
  AND U818 ( .A(n935), .B(n936), .Z(n933) );
  NANDN U819 ( .A(A[790]), .B(B[790]), .Z(n936) );
  NAND U820 ( .A(n937), .B(n938), .Z(n935) );
  NANDN U821 ( .A(B[790]), .B(A[790]), .Z(n938) );
  AND U822 ( .A(n939), .B(n940), .Z(n937) );
  NAND U823 ( .A(n941), .B(n942), .Z(n940) );
  NANDN U824 ( .A(A[789]), .B(B[789]), .Z(n942) );
  AND U825 ( .A(n943), .B(n944), .Z(n941) );
  NANDN U826 ( .A(A[788]), .B(B[788]), .Z(n944) );
  NAND U827 ( .A(n945), .B(n946), .Z(n943) );
  NANDN U828 ( .A(B[788]), .B(A[788]), .Z(n946) );
  AND U829 ( .A(n947), .B(n948), .Z(n945) );
  NAND U830 ( .A(n949), .B(n950), .Z(n948) );
  NANDN U831 ( .A(A[787]), .B(B[787]), .Z(n950) );
  AND U832 ( .A(n951), .B(n952), .Z(n949) );
  NANDN U833 ( .A(A[786]), .B(B[786]), .Z(n952) );
  NAND U834 ( .A(n953), .B(n954), .Z(n951) );
  NANDN U835 ( .A(B[786]), .B(A[786]), .Z(n954) );
  AND U836 ( .A(n955), .B(n956), .Z(n953) );
  NAND U837 ( .A(n957), .B(n958), .Z(n956) );
  NANDN U838 ( .A(A[785]), .B(B[785]), .Z(n958) );
  AND U839 ( .A(n959), .B(n960), .Z(n957) );
  NANDN U840 ( .A(A[784]), .B(B[784]), .Z(n960) );
  NAND U841 ( .A(n961), .B(n962), .Z(n959) );
  NANDN U842 ( .A(B[784]), .B(A[784]), .Z(n962) );
  AND U843 ( .A(n963), .B(n964), .Z(n961) );
  NAND U844 ( .A(n965), .B(n966), .Z(n964) );
  NANDN U845 ( .A(A[783]), .B(B[783]), .Z(n966) );
  AND U846 ( .A(n967), .B(n968), .Z(n965) );
  NANDN U847 ( .A(A[782]), .B(B[782]), .Z(n968) );
  NAND U848 ( .A(n969), .B(n970), .Z(n967) );
  NANDN U849 ( .A(B[782]), .B(A[782]), .Z(n970) );
  AND U850 ( .A(n971), .B(n972), .Z(n969) );
  NAND U851 ( .A(n973), .B(n974), .Z(n972) );
  NANDN U852 ( .A(A[781]), .B(B[781]), .Z(n974) );
  AND U853 ( .A(n975), .B(n976), .Z(n973) );
  NANDN U854 ( .A(A[780]), .B(B[780]), .Z(n976) );
  NAND U855 ( .A(n977), .B(n978), .Z(n975) );
  NANDN U856 ( .A(B[780]), .B(A[780]), .Z(n978) );
  AND U857 ( .A(n979), .B(n980), .Z(n977) );
  NAND U858 ( .A(n981), .B(n982), .Z(n980) );
  NANDN U859 ( .A(A[779]), .B(B[779]), .Z(n982) );
  AND U860 ( .A(n983), .B(n984), .Z(n981) );
  NANDN U861 ( .A(A[778]), .B(B[778]), .Z(n984) );
  NAND U862 ( .A(n985), .B(n986), .Z(n983) );
  NANDN U863 ( .A(B[778]), .B(A[778]), .Z(n986) );
  AND U864 ( .A(n987), .B(n988), .Z(n985) );
  NAND U865 ( .A(n989), .B(n990), .Z(n988) );
  NANDN U866 ( .A(A[777]), .B(B[777]), .Z(n990) );
  AND U867 ( .A(n991), .B(n992), .Z(n989) );
  NANDN U868 ( .A(A[776]), .B(B[776]), .Z(n992) );
  NAND U869 ( .A(n993), .B(n994), .Z(n991) );
  NANDN U870 ( .A(B[776]), .B(A[776]), .Z(n994) );
  AND U871 ( .A(n995), .B(n996), .Z(n993) );
  NAND U872 ( .A(n997), .B(n998), .Z(n996) );
  NANDN U873 ( .A(A[775]), .B(B[775]), .Z(n998) );
  AND U874 ( .A(n999), .B(n1000), .Z(n997) );
  NANDN U875 ( .A(A[774]), .B(B[774]), .Z(n1000) );
  NAND U876 ( .A(n1001), .B(n1002), .Z(n999) );
  NANDN U877 ( .A(B[774]), .B(A[774]), .Z(n1002) );
  AND U878 ( .A(n1003), .B(n1004), .Z(n1001) );
  NAND U879 ( .A(n1005), .B(n1006), .Z(n1004) );
  NANDN U880 ( .A(A[773]), .B(B[773]), .Z(n1006) );
  AND U881 ( .A(n1007), .B(n1008), .Z(n1005) );
  NANDN U882 ( .A(A[772]), .B(B[772]), .Z(n1008) );
  NAND U883 ( .A(n1009), .B(n1010), .Z(n1007) );
  NANDN U884 ( .A(B[772]), .B(A[772]), .Z(n1010) );
  AND U885 ( .A(n1011), .B(n1012), .Z(n1009) );
  NAND U886 ( .A(n1013), .B(n1014), .Z(n1012) );
  NANDN U887 ( .A(A[771]), .B(B[771]), .Z(n1014) );
  AND U888 ( .A(n1015), .B(n1016), .Z(n1013) );
  NANDN U889 ( .A(A[770]), .B(B[770]), .Z(n1016) );
  NAND U890 ( .A(n1017), .B(n1018), .Z(n1015) );
  NANDN U891 ( .A(B[770]), .B(A[770]), .Z(n1018) );
  AND U892 ( .A(n1019), .B(n1020), .Z(n1017) );
  NAND U893 ( .A(n1021), .B(n1022), .Z(n1020) );
  NANDN U894 ( .A(A[769]), .B(B[769]), .Z(n1022) );
  AND U895 ( .A(n1023), .B(n1024), .Z(n1021) );
  NANDN U896 ( .A(A[768]), .B(B[768]), .Z(n1024) );
  NAND U897 ( .A(n1025), .B(n1026), .Z(n1023) );
  NANDN U898 ( .A(B[768]), .B(A[768]), .Z(n1026) );
  AND U899 ( .A(n1027), .B(n1028), .Z(n1025) );
  NAND U900 ( .A(n1029), .B(n1030), .Z(n1028) );
  NANDN U901 ( .A(A[767]), .B(B[767]), .Z(n1030) );
  AND U902 ( .A(n1031), .B(n1032), .Z(n1029) );
  NANDN U903 ( .A(A[766]), .B(B[766]), .Z(n1032) );
  NAND U904 ( .A(n1033), .B(n1034), .Z(n1031) );
  NANDN U905 ( .A(B[766]), .B(A[766]), .Z(n1034) );
  AND U906 ( .A(n1035), .B(n1036), .Z(n1033) );
  NAND U907 ( .A(n1037), .B(n1038), .Z(n1036) );
  NANDN U908 ( .A(A[765]), .B(B[765]), .Z(n1038) );
  AND U909 ( .A(n1039), .B(n1040), .Z(n1037) );
  NANDN U910 ( .A(A[764]), .B(B[764]), .Z(n1040) );
  NAND U911 ( .A(n1041), .B(n1042), .Z(n1039) );
  NANDN U912 ( .A(B[764]), .B(A[764]), .Z(n1042) );
  AND U913 ( .A(n1043), .B(n1044), .Z(n1041) );
  NAND U914 ( .A(n1045), .B(n1046), .Z(n1044) );
  NANDN U915 ( .A(A[763]), .B(B[763]), .Z(n1046) );
  AND U916 ( .A(n1047), .B(n1048), .Z(n1045) );
  NANDN U917 ( .A(A[762]), .B(B[762]), .Z(n1048) );
  NAND U918 ( .A(n1049), .B(n1050), .Z(n1047) );
  NANDN U919 ( .A(B[762]), .B(A[762]), .Z(n1050) );
  AND U920 ( .A(n1051), .B(n1052), .Z(n1049) );
  NAND U921 ( .A(n1053), .B(n1054), .Z(n1052) );
  NANDN U922 ( .A(A[761]), .B(B[761]), .Z(n1054) );
  AND U923 ( .A(n1055), .B(n1056), .Z(n1053) );
  NANDN U924 ( .A(A[760]), .B(B[760]), .Z(n1056) );
  NAND U925 ( .A(n1057), .B(n1058), .Z(n1055) );
  NANDN U926 ( .A(B[760]), .B(A[760]), .Z(n1058) );
  AND U927 ( .A(n1059), .B(n1060), .Z(n1057) );
  NAND U928 ( .A(n1061), .B(n1062), .Z(n1060) );
  NANDN U929 ( .A(A[759]), .B(B[759]), .Z(n1062) );
  AND U930 ( .A(n1063), .B(n1064), .Z(n1061) );
  NANDN U931 ( .A(A[758]), .B(B[758]), .Z(n1064) );
  NAND U932 ( .A(n1065), .B(n1066), .Z(n1063) );
  NANDN U933 ( .A(B[758]), .B(A[758]), .Z(n1066) );
  AND U934 ( .A(n1067), .B(n1068), .Z(n1065) );
  NAND U935 ( .A(n1069), .B(n1070), .Z(n1068) );
  NANDN U936 ( .A(A[757]), .B(B[757]), .Z(n1070) );
  AND U937 ( .A(n1071), .B(n1072), .Z(n1069) );
  NANDN U938 ( .A(A[756]), .B(B[756]), .Z(n1072) );
  NAND U939 ( .A(n1073), .B(n1074), .Z(n1071) );
  NANDN U940 ( .A(B[756]), .B(A[756]), .Z(n1074) );
  AND U941 ( .A(n1075), .B(n1076), .Z(n1073) );
  NAND U942 ( .A(n1077), .B(n1078), .Z(n1076) );
  NANDN U943 ( .A(A[755]), .B(B[755]), .Z(n1078) );
  AND U944 ( .A(n1079), .B(n1080), .Z(n1077) );
  NANDN U945 ( .A(A[754]), .B(B[754]), .Z(n1080) );
  NAND U946 ( .A(n1081), .B(n1082), .Z(n1079) );
  NANDN U947 ( .A(B[754]), .B(A[754]), .Z(n1082) );
  AND U948 ( .A(n1083), .B(n1084), .Z(n1081) );
  NAND U949 ( .A(n1085), .B(n1086), .Z(n1084) );
  NANDN U950 ( .A(A[753]), .B(B[753]), .Z(n1086) );
  AND U951 ( .A(n1087), .B(n1088), .Z(n1085) );
  NANDN U952 ( .A(A[752]), .B(B[752]), .Z(n1088) );
  NAND U953 ( .A(n1089), .B(n1090), .Z(n1087) );
  NANDN U954 ( .A(B[752]), .B(A[752]), .Z(n1090) );
  AND U955 ( .A(n1091), .B(n1092), .Z(n1089) );
  NAND U956 ( .A(n1093), .B(n1094), .Z(n1092) );
  NANDN U957 ( .A(A[751]), .B(B[751]), .Z(n1094) );
  AND U958 ( .A(n1095), .B(n1096), .Z(n1093) );
  NANDN U959 ( .A(A[750]), .B(B[750]), .Z(n1096) );
  NAND U960 ( .A(n1097), .B(n1098), .Z(n1095) );
  NANDN U961 ( .A(B[750]), .B(A[750]), .Z(n1098) );
  AND U962 ( .A(n1099), .B(n1100), .Z(n1097) );
  NAND U963 ( .A(n1101), .B(n1102), .Z(n1100) );
  NANDN U964 ( .A(A[749]), .B(B[749]), .Z(n1102) );
  AND U965 ( .A(n1103), .B(n1104), .Z(n1101) );
  NANDN U966 ( .A(A[748]), .B(B[748]), .Z(n1104) );
  NAND U967 ( .A(n1105), .B(n1106), .Z(n1103) );
  NANDN U968 ( .A(B[748]), .B(A[748]), .Z(n1106) );
  AND U969 ( .A(n1107), .B(n1108), .Z(n1105) );
  NAND U970 ( .A(n1109), .B(n1110), .Z(n1108) );
  NANDN U971 ( .A(A[747]), .B(B[747]), .Z(n1110) );
  AND U972 ( .A(n1111), .B(n1112), .Z(n1109) );
  NANDN U973 ( .A(A[746]), .B(B[746]), .Z(n1112) );
  NAND U974 ( .A(n1113), .B(n1114), .Z(n1111) );
  NANDN U975 ( .A(B[746]), .B(A[746]), .Z(n1114) );
  AND U976 ( .A(n1115), .B(n1116), .Z(n1113) );
  NAND U977 ( .A(n1117), .B(n1118), .Z(n1116) );
  NANDN U978 ( .A(A[745]), .B(B[745]), .Z(n1118) );
  AND U979 ( .A(n1119), .B(n1120), .Z(n1117) );
  NANDN U980 ( .A(A[744]), .B(B[744]), .Z(n1120) );
  NAND U981 ( .A(n1121), .B(n1122), .Z(n1119) );
  NANDN U982 ( .A(B[744]), .B(A[744]), .Z(n1122) );
  AND U983 ( .A(n1123), .B(n1124), .Z(n1121) );
  NAND U984 ( .A(n1125), .B(n1126), .Z(n1124) );
  NANDN U985 ( .A(A[743]), .B(B[743]), .Z(n1126) );
  AND U986 ( .A(n1127), .B(n1128), .Z(n1125) );
  NANDN U987 ( .A(A[742]), .B(B[742]), .Z(n1128) );
  NAND U988 ( .A(n1129), .B(n1130), .Z(n1127) );
  NANDN U989 ( .A(B[742]), .B(A[742]), .Z(n1130) );
  AND U990 ( .A(n1131), .B(n1132), .Z(n1129) );
  NAND U991 ( .A(n1133), .B(n1134), .Z(n1132) );
  NANDN U992 ( .A(A[741]), .B(B[741]), .Z(n1134) );
  AND U993 ( .A(n1135), .B(n1136), .Z(n1133) );
  NANDN U994 ( .A(A[740]), .B(B[740]), .Z(n1136) );
  NAND U995 ( .A(n1137), .B(n1138), .Z(n1135) );
  NANDN U996 ( .A(B[740]), .B(A[740]), .Z(n1138) );
  AND U997 ( .A(n1139), .B(n1140), .Z(n1137) );
  NAND U998 ( .A(n1141), .B(n1142), .Z(n1140) );
  NANDN U999 ( .A(A[739]), .B(B[739]), .Z(n1142) );
  AND U1000 ( .A(n1143), .B(n1144), .Z(n1141) );
  NANDN U1001 ( .A(A[738]), .B(B[738]), .Z(n1144) );
  NAND U1002 ( .A(n1145), .B(n1146), .Z(n1143) );
  NANDN U1003 ( .A(B[738]), .B(A[738]), .Z(n1146) );
  AND U1004 ( .A(n1147), .B(n1148), .Z(n1145) );
  NAND U1005 ( .A(n1149), .B(n1150), .Z(n1148) );
  NANDN U1006 ( .A(A[737]), .B(B[737]), .Z(n1150) );
  AND U1007 ( .A(n1151), .B(n1152), .Z(n1149) );
  NANDN U1008 ( .A(A[736]), .B(B[736]), .Z(n1152) );
  NAND U1009 ( .A(n1153), .B(n1154), .Z(n1151) );
  NANDN U1010 ( .A(B[736]), .B(A[736]), .Z(n1154) );
  AND U1011 ( .A(n1155), .B(n1156), .Z(n1153) );
  NAND U1012 ( .A(n1157), .B(n1158), .Z(n1156) );
  NANDN U1013 ( .A(A[735]), .B(B[735]), .Z(n1158) );
  AND U1014 ( .A(n1159), .B(n1160), .Z(n1157) );
  NANDN U1015 ( .A(A[734]), .B(B[734]), .Z(n1160) );
  NAND U1016 ( .A(n1161), .B(n1162), .Z(n1159) );
  NANDN U1017 ( .A(B[734]), .B(A[734]), .Z(n1162) );
  AND U1018 ( .A(n1163), .B(n1164), .Z(n1161) );
  NAND U1019 ( .A(n1165), .B(n1166), .Z(n1164) );
  NANDN U1020 ( .A(A[733]), .B(B[733]), .Z(n1166) );
  AND U1021 ( .A(n1167), .B(n1168), .Z(n1165) );
  NANDN U1022 ( .A(A[732]), .B(B[732]), .Z(n1168) );
  NAND U1023 ( .A(n1169), .B(n1170), .Z(n1167) );
  NANDN U1024 ( .A(B[732]), .B(A[732]), .Z(n1170) );
  AND U1025 ( .A(n1171), .B(n1172), .Z(n1169) );
  NAND U1026 ( .A(n1173), .B(n1174), .Z(n1172) );
  NANDN U1027 ( .A(A[731]), .B(B[731]), .Z(n1174) );
  AND U1028 ( .A(n1175), .B(n1176), .Z(n1173) );
  NANDN U1029 ( .A(A[730]), .B(B[730]), .Z(n1176) );
  NAND U1030 ( .A(n1177), .B(n1178), .Z(n1175) );
  NANDN U1031 ( .A(B[730]), .B(A[730]), .Z(n1178) );
  AND U1032 ( .A(n1179), .B(n1180), .Z(n1177) );
  NAND U1033 ( .A(n1181), .B(n1182), .Z(n1180) );
  NANDN U1034 ( .A(A[729]), .B(B[729]), .Z(n1182) );
  AND U1035 ( .A(n1183), .B(n1184), .Z(n1181) );
  NANDN U1036 ( .A(A[728]), .B(B[728]), .Z(n1184) );
  NAND U1037 ( .A(n1185), .B(n1186), .Z(n1183) );
  NANDN U1038 ( .A(B[728]), .B(A[728]), .Z(n1186) );
  AND U1039 ( .A(n1187), .B(n1188), .Z(n1185) );
  NAND U1040 ( .A(n1189), .B(n1190), .Z(n1188) );
  NANDN U1041 ( .A(A[727]), .B(B[727]), .Z(n1190) );
  AND U1042 ( .A(n1191), .B(n1192), .Z(n1189) );
  NANDN U1043 ( .A(A[726]), .B(B[726]), .Z(n1192) );
  NAND U1044 ( .A(n1193), .B(n1194), .Z(n1191) );
  NANDN U1045 ( .A(B[726]), .B(A[726]), .Z(n1194) );
  AND U1046 ( .A(n1195), .B(n1196), .Z(n1193) );
  NAND U1047 ( .A(n1197), .B(n1198), .Z(n1196) );
  NANDN U1048 ( .A(A[725]), .B(B[725]), .Z(n1198) );
  AND U1049 ( .A(n1199), .B(n1200), .Z(n1197) );
  NANDN U1050 ( .A(A[724]), .B(B[724]), .Z(n1200) );
  NAND U1051 ( .A(n1201), .B(n1202), .Z(n1199) );
  NANDN U1052 ( .A(B[724]), .B(A[724]), .Z(n1202) );
  AND U1053 ( .A(n1203), .B(n1204), .Z(n1201) );
  NAND U1054 ( .A(n1205), .B(n1206), .Z(n1204) );
  NANDN U1055 ( .A(A[723]), .B(B[723]), .Z(n1206) );
  AND U1056 ( .A(n1207), .B(n1208), .Z(n1205) );
  NANDN U1057 ( .A(A[722]), .B(B[722]), .Z(n1208) );
  NAND U1058 ( .A(n1209), .B(n1210), .Z(n1207) );
  NANDN U1059 ( .A(B[722]), .B(A[722]), .Z(n1210) );
  AND U1060 ( .A(n1211), .B(n1212), .Z(n1209) );
  NAND U1061 ( .A(n1213), .B(n1214), .Z(n1212) );
  NANDN U1062 ( .A(A[721]), .B(B[721]), .Z(n1214) );
  AND U1063 ( .A(n1215), .B(n1216), .Z(n1213) );
  NANDN U1064 ( .A(A[720]), .B(B[720]), .Z(n1216) );
  NAND U1065 ( .A(n1217), .B(n1218), .Z(n1215) );
  NANDN U1066 ( .A(B[720]), .B(A[720]), .Z(n1218) );
  AND U1067 ( .A(n1219), .B(n1220), .Z(n1217) );
  NAND U1068 ( .A(n1221), .B(n1222), .Z(n1220) );
  NANDN U1069 ( .A(A[719]), .B(B[719]), .Z(n1222) );
  AND U1070 ( .A(n1223), .B(n1224), .Z(n1221) );
  NANDN U1071 ( .A(A[718]), .B(B[718]), .Z(n1224) );
  NAND U1072 ( .A(n1225), .B(n1226), .Z(n1223) );
  NANDN U1073 ( .A(B[718]), .B(A[718]), .Z(n1226) );
  AND U1074 ( .A(n1227), .B(n1228), .Z(n1225) );
  NAND U1075 ( .A(n1229), .B(n1230), .Z(n1228) );
  NANDN U1076 ( .A(A[717]), .B(B[717]), .Z(n1230) );
  AND U1077 ( .A(n1231), .B(n1232), .Z(n1229) );
  NANDN U1078 ( .A(A[716]), .B(B[716]), .Z(n1232) );
  NAND U1079 ( .A(n1233), .B(n1234), .Z(n1231) );
  NANDN U1080 ( .A(B[716]), .B(A[716]), .Z(n1234) );
  AND U1081 ( .A(n1235), .B(n1236), .Z(n1233) );
  NAND U1082 ( .A(n1237), .B(n1238), .Z(n1236) );
  NANDN U1083 ( .A(A[715]), .B(B[715]), .Z(n1238) );
  AND U1084 ( .A(n1239), .B(n1240), .Z(n1237) );
  NANDN U1085 ( .A(A[714]), .B(B[714]), .Z(n1240) );
  NAND U1086 ( .A(n1241), .B(n1242), .Z(n1239) );
  NANDN U1087 ( .A(B[714]), .B(A[714]), .Z(n1242) );
  AND U1088 ( .A(n1243), .B(n1244), .Z(n1241) );
  NAND U1089 ( .A(n1245), .B(n1246), .Z(n1244) );
  NANDN U1090 ( .A(A[713]), .B(B[713]), .Z(n1246) );
  AND U1091 ( .A(n1247), .B(n1248), .Z(n1245) );
  NANDN U1092 ( .A(A[712]), .B(B[712]), .Z(n1248) );
  NAND U1093 ( .A(n1249), .B(n1250), .Z(n1247) );
  NANDN U1094 ( .A(B[712]), .B(A[712]), .Z(n1250) );
  AND U1095 ( .A(n1251), .B(n1252), .Z(n1249) );
  NAND U1096 ( .A(n1253), .B(n1254), .Z(n1252) );
  NANDN U1097 ( .A(A[711]), .B(B[711]), .Z(n1254) );
  AND U1098 ( .A(n1255), .B(n1256), .Z(n1253) );
  NANDN U1099 ( .A(A[710]), .B(B[710]), .Z(n1256) );
  NAND U1100 ( .A(n1257), .B(n1258), .Z(n1255) );
  NANDN U1101 ( .A(B[710]), .B(A[710]), .Z(n1258) );
  AND U1102 ( .A(n1259), .B(n1260), .Z(n1257) );
  NAND U1103 ( .A(n1261), .B(n1262), .Z(n1260) );
  NANDN U1104 ( .A(A[709]), .B(B[709]), .Z(n1262) );
  AND U1105 ( .A(n1263), .B(n1264), .Z(n1261) );
  NANDN U1106 ( .A(A[708]), .B(B[708]), .Z(n1264) );
  NAND U1107 ( .A(n1265), .B(n1266), .Z(n1263) );
  NANDN U1108 ( .A(B[708]), .B(A[708]), .Z(n1266) );
  AND U1109 ( .A(n1267), .B(n1268), .Z(n1265) );
  NAND U1110 ( .A(n1269), .B(n1270), .Z(n1268) );
  NANDN U1111 ( .A(A[707]), .B(B[707]), .Z(n1270) );
  AND U1112 ( .A(n1271), .B(n1272), .Z(n1269) );
  NANDN U1113 ( .A(A[706]), .B(B[706]), .Z(n1272) );
  NAND U1114 ( .A(n1273), .B(n1274), .Z(n1271) );
  NANDN U1115 ( .A(B[706]), .B(A[706]), .Z(n1274) );
  AND U1116 ( .A(n1275), .B(n1276), .Z(n1273) );
  NAND U1117 ( .A(n1277), .B(n1278), .Z(n1276) );
  NANDN U1118 ( .A(A[705]), .B(B[705]), .Z(n1278) );
  AND U1119 ( .A(n1279), .B(n1280), .Z(n1277) );
  NANDN U1120 ( .A(A[704]), .B(B[704]), .Z(n1280) );
  NAND U1121 ( .A(n1281), .B(n1282), .Z(n1279) );
  NANDN U1122 ( .A(B[704]), .B(A[704]), .Z(n1282) );
  AND U1123 ( .A(n1283), .B(n1284), .Z(n1281) );
  NAND U1124 ( .A(n1285), .B(n1286), .Z(n1284) );
  NANDN U1125 ( .A(A[703]), .B(B[703]), .Z(n1286) );
  AND U1126 ( .A(n1287), .B(n1288), .Z(n1285) );
  NANDN U1127 ( .A(A[702]), .B(B[702]), .Z(n1288) );
  NAND U1128 ( .A(n1289), .B(n1290), .Z(n1287) );
  NANDN U1129 ( .A(B[702]), .B(A[702]), .Z(n1290) );
  AND U1130 ( .A(n1291), .B(n1292), .Z(n1289) );
  NAND U1131 ( .A(n1293), .B(n1294), .Z(n1292) );
  NANDN U1132 ( .A(A[701]), .B(B[701]), .Z(n1294) );
  AND U1133 ( .A(n1295), .B(n1296), .Z(n1293) );
  NANDN U1134 ( .A(A[700]), .B(B[700]), .Z(n1296) );
  NAND U1135 ( .A(n1297), .B(n1298), .Z(n1295) );
  NANDN U1136 ( .A(B[700]), .B(A[700]), .Z(n1298) );
  AND U1137 ( .A(n1299), .B(n1300), .Z(n1297) );
  NAND U1138 ( .A(n1301), .B(n1302), .Z(n1300) );
  NANDN U1139 ( .A(A[699]), .B(B[699]), .Z(n1302) );
  AND U1140 ( .A(n1303), .B(n1304), .Z(n1301) );
  NANDN U1141 ( .A(A[698]), .B(B[698]), .Z(n1304) );
  NAND U1142 ( .A(n1305), .B(n1306), .Z(n1303) );
  NANDN U1143 ( .A(B[698]), .B(A[698]), .Z(n1306) );
  AND U1144 ( .A(n1307), .B(n1308), .Z(n1305) );
  NAND U1145 ( .A(n1309), .B(n1310), .Z(n1308) );
  NANDN U1146 ( .A(A[697]), .B(B[697]), .Z(n1310) );
  AND U1147 ( .A(n1311), .B(n1312), .Z(n1309) );
  NANDN U1148 ( .A(A[696]), .B(B[696]), .Z(n1312) );
  NAND U1149 ( .A(n1313), .B(n1314), .Z(n1311) );
  NANDN U1150 ( .A(B[696]), .B(A[696]), .Z(n1314) );
  AND U1151 ( .A(n1315), .B(n1316), .Z(n1313) );
  NAND U1152 ( .A(n1317), .B(n1318), .Z(n1316) );
  NANDN U1153 ( .A(A[695]), .B(B[695]), .Z(n1318) );
  AND U1154 ( .A(n1319), .B(n1320), .Z(n1317) );
  NANDN U1155 ( .A(A[694]), .B(B[694]), .Z(n1320) );
  NAND U1156 ( .A(n1321), .B(n1322), .Z(n1319) );
  NANDN U1157 ( .A(B[694]), .B(A[694]), .Z(n1322) );
  AND U1158 ( .A(n1323), .B(n1324), .Z(n1321) );
  NAND U1159 ( .A(n1325), .B(n1326), .Z(n1324) );
  NANDN U1160 ( .A(A[693]), .B(B[693]), .Z(n1326) );
  AND U1161 ( .A(n1327), .B(n1328), .Z(n1325) );
  NANDN U1162 ( .A(A[692]), .B(B[692]), .Z(n1328) );
  NAND U1163 ( .A(n1329), .B(n1330), .Z(n1327) );
  NANDN U1164 ( .A(B[692]), .B(A[692]), .Z(n1330) );
  AND U1165 ( .A(n1331), .B(n1332), .Z(n1329) );
  NAND U1166 ( .A(n1333), .B(n1334), .Z(n1332) );
  NANDN U1167 ( .A(A[691]), .B(B[691]), .Z(n1334) );
  AND U1168 ( .A(n1335), .B(n1336), .Z(n1333) );
  NANDN U1169 ( .A(A[690]), .B(B[690]), .Z(n1336) );
  NAND U1170 ( .A(n1337), .B(n1338), .Z(n1335) );
  NANDN U1171 ( .A(B[690]), .B(A[690]), .Z(n1338) );
  AND U1172 ( .A(n1339), .B(n1340), .Z(n1337) );
  NAND U1173 ( .A(n1341), .B(n1342), .Z(n1340) );
  NANDN U1174 ( .A(A[689]), .B(B[689]), .Z(n1342) );
  AND U1175 ( .A(n1343), .B(n1344), .Z(n1341) );
  NANDN U1176 ( .A(A[688]), .B(B[688]), .Z(n1344) );
  NAND U1177 ( .A(n1345), .B(n1346), .Z(n1343) );
  NANDN U1178 ( .A(B[688]), .B(A[688]), .Z(n1346) );
  AND U1179 ( .A(n1347), .B(n1348), .Z(n1345) );
  NAND U1180 ( .A(n1349), .B(n1350), .Z(n1348) );
  NANDN U1181 ( .A(A[687]), .B(B[687]), .Z(n1350) );
  AND U1182 ( .A(n1351), .B(n1352), .Z(n1349) );
  NANDN U1183 ( .A(A[686]), .B(B[686]), .Z(n1352) );
  NAND U1184 ( .A(n1353), .B(n1354), .Z(n1351) );
  NANDN U1185 ( .A(B[686]), .B(A[686]), .Z(n1354) );
  AND U1186 ( .A(n1355), .B(n1356), .Z(n1353) );
  NAND U1187 ( .A(n1357), .B(n1358), .Z(n1356) );
  NANDN U1188 ( .A(A[685]), .B(B[685]), .Z(n1358) );
  AND U1189 ( .A(n1359), .B(n1360), .Z(n1357) );
  NANDN U1190 ( .A(A[684]), .B(B[684]), .Z(n1360) );
  NAND U1191 ( .A(n1361), .B(n1362), .Z(n1359) );
  NANDN U1192 ( .A(B[684]), .B(A[684]), .Z(n1362) );
  AND U1193 ( .A(n1363), .B(n1364), .Z(n1361) );
  NAND U1194 ( .A(n1365), .B(n1366), .Z(n1364) );
  NANDN U1195 ( .A(A[683]), .B(B[683]), .Z(n1366) );
  AND U1196 ( .A(n1367), .B(n1368), .Z(n1365) );
  NANDN U1197 ( .A(A[682]), .B(B[682]), .Z(n1368) );
  NAND U1198 ( .A(n1369), .B(n1370), .Z(n1367) );
  NANDN U1199 ( .A(B[682]), .B(A[682]), .Z(n1370) );
  AND U1200 ( .A(n1371), .B(n1372), .Z(n1369) );
  NAND U1201 ( .A(n1373), .B(n1374), .Z(n1372) );
  NANDN U1202 ( .A(A[681]), .B(B[681]), .Z(n1374) );
  AND U1203 ( .A(n1375), .B(n1376), .Z(n1373) );
  NANDN U1204 ( .A(A[680]), .B(B[680]), .Z(n1376) );
  NAND U1205 ( .A(n1377), .B(n1378), .Z(n1375) );
  NANDN U1206 ( .A(B[680]), .B(A[680]), .Z(n1378) );
  AND U1207 ( .A(n1379), .B(n1380), .Z(n1377) );
  NAND U1208 ( .A(n1381), .B(n1382), .Z(n1380) );
  NANDN U1209 ( .A(A[679]), .B(B[679]), .Z(n1382) );
  AND U1210 ( .A(n1383), .B(n1384), .Z(n1381) );
  NANDN U1211 ( .A(A[678]), .B(B[678]), .Z(n1384) );
  NAND U1212 ( .A(n1385), .B(n1386), .Z(n1383) );
  NANDN U1213 ( .A(B[678]), .B(A[678]), .Z(n1386) );
  AND U1214 ( .A(n1387), .B(n1388), .Z(n1385) );
  NAND U1215 ( .A(n1389), .B(n1390), .Z(n1388) );
  NANDN U1216 ( .A(A[677]), .B(B[677]), .Z(n1390) );
  AND U1217 ( .A(n1391), .B(n1392), .Z(n1389) );
  NANDN U1218 ( .A(A[676]), .B(B[676]), .Z(n1392) );
  NAND U1219 ( .A(n1393), .B(n1394), .Z(n1391) );
  NANDN U1220 ( .A(B[676]), .B(A[676]), .Z(n1394) );
  AND U1221 ( .A(n1395), .B(n1396), .Z(n1393) );
  NAND U1222 ( .A(n1397), .B(n1398), .Z(n1396) );
  NANDN U1223 ( .A(A[675]), .B(B[675]), .Z(n1398) );
  AND U1224 ( .A(n1399), .B(n1400), .Z(n1397) );
  NANDN U1225 ( .A(A[674]), .B(B[674]), .Z(n1400) );
  NAND U1226 ( .A(n1401), .B(n1402), .Z(n1399) );
  NANDN U1227 ( .A(B[674]), .B(A[674]), .Z(n1402) );
  AND U1228 ( .A(n1403), .B(n1404), .Z(n1401) );
  NAND U1229 ( .A(n1405), .B(n1406), .Z(n1404) );
  NANDN U1230 ( .A(A[673]), .B(B[673]), .Z(n1406) );
  AND U1231 ( .A(n1407), .B(n1408), .Z(n1405) );
  NANDN U1232 ( .A(A[672]), .B(B[672]), .Z(n1408) );
  NAND U1233 ( .A(n1409), .B(n1410), .Z(n1407) );
  NANDN U1234 ( .A(B[672]), .B(A[672]), .Z(n1410) );
  AND U1235 ( .A(n1411), .B(n1412), .Z(n1409) );
  NAND U1236 ( .A(n1413), .B(n1414), .Z(n1412) );
  NANDN U1237 ( .A(A[671]), .B(B[671]), .Z(n1414) );
  AND U1238 ( .A(n1415), .B(n1416), .Z(n1413) );
  NANDN U1239 ( .A(A[670]), .B(B[670]), .Z(n1416) );
  NAND U1240 ( .A(n1417), .B(n1418), .Z(n1415) );
  NANDN U1241 ( .A(B[670]), .B(A[670]), .Z(n1418) );
  AND U1242 ( .A(n1419), .B(n1420), .Z(n1417) );
  NAND U1243 ( .A(n1421), .B(n1422), .Z(n1420) );
  NANDN U1244 ( .A(A[669]), .B(B[669]), .Z(n1422) );
  AND U1245 ( .A(n1423), .B(n1424), .Z(n1421) );
  NANDN U1246 ( .A(A[668]), .B(B[668]), .Z(n1424) );
  NAND U1247 ( .A(n1425), .B(n1426), .Z(n1423) );
  NANDN U1248 ( .A(B[668]), .B(A[668]), .Z(n1426) );
  AND U1249 ( .A(n1427), .B(n1428), .Z(n1425) );
  NAND U1250 ( .A(n1429), .B(n1430), .Z(n1428) );
  NANDN U1251 ( .A(A[667]), .B(B[667]), .Z(n1430) );
  AND U1252 ( .A(n1431), .B(n1432), .Z(n1429) );
  NANDN U1253 ( .A(A[666]), .B(B[666]), .Z(n1432) );
  NAND U1254 ( .A(n1433), .B(n1434), .Z(n1431) );
  NANDN U1255 ( .A(B[666]), .B(A[666]), .Z(n1434) );
  AND U1256 ( .A(n1435), .B(n1436), .Z(n1433) );
  NAND U1257 ( .A(n1437), .B(n1438), .Z(n1436) );
  NANDN U1258 ( .A(A[665]), .B(B[665]), .Z(n1438) );
  AND U1259 ( .A(n1439), .B(n1440), .Z(n1437) );
  NANDN U1260 ( .A(A[664]), .B(B[664]), .Z(n1440) );
  NAND U1261 ( .A(n1441), .B(n1442), .Z(n1439) );
  NANDN U1262 ( .A(B[664]), .B(A[664]), .Z(n1442) );
  AND U1263 ( .A(n1443), .B(n1444), .Z(n1441) );
  NAND U1264 ( .A(n1445), .B(n1446), .Z(n1444) );
  NANDN U1265 ( .A(A[663]), .B(B[663]), .Z(n1446) );
  AND U1266 ( .A(n1447), .B(n1448), .Z(n1445) );
  NANDN U1267 ( .A(A[662]), .B(B[662]), .Z(n1448) );
  NAND U1268 ( .A(n1449), .B(n1450), .Z(n1447) );
  NANDN U1269 ( .A(B[662]), .B(A[662]), .Z(n1450) );
  AND U1270 ( .A(n1451), .B(n1452), .Z(n1449) );
  NAND U1271 ( .A(n1453), .B(n1454), .Z(n1452) );
  NANDN U1272 ( .A(A[661]), .B(B[661]), .Z(n1454) );
  AND U1273 ( .A(n1455), .B(n1456), .Z(n1453) );
  NANDN U1274 ( .A(A[660]), .B(B[660]), .Z(n1456) );
  NAND U1275 ( .A(n1457), .B(n1458), .Z(n1455) );
  NANDN U1276 ( .A(B[660]), .B(A[660]), .Z(n1458) );
  AND U1277 ( .A(n1459), .B(n1460), .Z(n1457) );
  NAND U1278 ( .A(n1461), .B(n1462), .Z(n1460) );
  NANDN U1279 ( .A(A[659]), .B(B[659]), .Z(n1462) );
  AND U1280 ( .A(n1463), .B(n1464), .Z(n1461) );
  NANDN U1281 ( .A(A[658]), .B(B[658]), .Z(n1464) );
  NAND U1282 ( .A(n1465), .B(n1466), .Z(n1463) );
  NANDN U1283 ( .A(B[658]), .B(A[658]), .Z(n1466) );
  AND U1284 ( .A(n1467), .B(n1468), .Z(n1465) );
  NAND U1285 ( .A(n1469), .B(n1470), .Z(n1468) );
  NANDN U1286 ( .A(A[657]), .B(B[657]), .Z(n1470) );
  AND U1287 ( .A(n1471), .B(n1472), .Z(n1469) );
  NANDN U1288 ( .A(A[656]), .B(B[656]), .Z(n1472) );
  NAND U1289 ( .A(n1473), .B(n1474), .Z(n1471) );
  NANDN U1290 ( .A(B[656]), .B(A[656]), .Z(n1474) );
  AND U1291 ( .A(n1475), .B(n1476), .Z(n1473) );
  NAND U1292 ( .A(n1477), .B(n1478), .Z(n1476) );
  NANDN U1293 ( .A(A[655]), .B(B[655]), .Z(n1478) );
  AND U1294 ( .A(n1479), .B(n1480), .Z(n1477) );
  NANDN U1295 ( .A(A[654]), .B(B[654]), .Z(n1480) );
  NAND U1296 ( .A(n1481), .B(n1482), .Z(n1479) );
  NANDN U1297 ( .A(B[654]), .B(A[654]), .Z(n1482) );
  AND U1298 ( .A(n1483), .B(n1484), .Z(n1481) );
  NAND U1299 ( .A(n1485), .B(n1486), .Z(n1484) );
  NANDN U1300 ( .A(A[653]), .B(B[653]), .Z(n1486) );
  AND U1301 ( .A(n1487), .B(n1488), .Z(n1485) );
  NANDN U1302 ( .A(A[652]), .B(B[652]), .Z(n1488) );
  NAND U1303 ( .A(n1489), .B(n1490), .Z(n1487) );
  NANDN U1304 ( .A(B[652]), .B(A[652]), .Z(n1490) );
  AND U1305 ( .A(n1491), .B(n1492), .Z(n1489) );
  NAND U1306 ( .A(n1493), .B(n1494), .Z(n1492) );
  NANDN U1307 ( .A(A[651]), .B(B[651]), .Z(n1494) );
  AND U1308 ( .A(n1495), .B(n1496), .Z(n1493) );
  NANDN U1309 ( .A(A[650]), .B(B[650]), .Z(n1496) );
  NAND U1310 ( .A(n1497), .B(n1498), .Z(n1495) );
  NANDN U1311 ( .A(B[650]), .B(A[650]), .Z(n1498) );
  AND U1312 ( .A(n1499), .B(n1500), .Z(n1497) );
  NAND U1313 ( .A(n1501), .B(n1502), .Z(n1500) );
  NANDN U1314 ( .A(A[649]), .B(B[649]), .Z(n1502) );
  AND U1315 ( .A(n1503), .B(n1504), .Z(n1501) );
  NANDN U1316 ( .A(A[648]), .B(B[648]), .Z(n1504) );
  NAND U1317 ( .A(n1505), .B(n1506), .Z(n1503) );
  NANDN U1318 ( .A(B[648]), .B(A[648]), .Z(n1506) );
  AND U1319 ( .A(n1507), .B(n1508), .Z(n1505) );
  NAND U1320 ( .A(n1509), .B(n1510), .Z(n1508) );
  NANDN U1321 ( .A(A[647]), .B(B[647]), .Z(n1510) );
  AND U1322 ( .A(n1511), .B(n1512), .Z(n1509) );
  NANDN U1323 ( .A(A[646]), .B(B[646]), .Z(n1512) );
  NAND U1324 ( .A(n1513), .B(n1514), .Z(n1511) );
  NANDN U1325 ( .A(B[646]), .B(A[646]), .Z(n1514) );
  AND U1326 ( .A(n1515), .B(n1516), .Z(n1513) );
  NAND U1327 ( .A(n1517), .B(n1518), .Z(n1516) );
  NANDN U1328 ( .A(A[645]), .B(B[645]), .Z(n1518) );
  AND U1329 ( .A(n1519), .B(n1520), .Z(n1517) );
  NANDN U1330 ( .A(A[644]), .B(B[644]), .Z(n1520) );
  NAND U1331 ( .A(n1521), .B(n1522), .Z(n1519) );
  NANDN U1332 ( .A(B[644]), .B(A[644]), .Z(n1522) );
  AND U1333 ( .A(n1523), .B(n1524), .Z(n1521) );
  NAND U1334 ( .A(n1525), .B(n1526), .Z(n1524) );
  NANDN U1335 ( .A(A[643]), .B(B[643]), .Z(n1526) );
  AND U1336 ( .A(n1527), .B(n1528), .Z(n1525) );
  NANDN U1337 ( .A(A[642]), .B(B[642]), .Z(n1528) );
  NAND U1338 ( .A(n1529), .B(n1530), .Z(n1527) );
  NANDN U1339 ( .A(B[642]), .B(A[642]), .Z(n1530) );
  AND U1340 ( .A(n1531), .B(n1532), .Z(n1529) );
  NAND U1341 ( .A(n1533), .B(n1534), .Z(n1532) );
  NANDN U1342 ( .A(A[641]), .B(B[641]), .Z(n1534) );
  AND U1343 ( .A(n1535), .B(n1536), .Z(n1533) );
  NANDN U1344 ( .A(A[640]), .B(B[640]), .Z(n1536) );
  NAND U1345 ( .A(n1537), .B(n1538), .Z(n1535) );
  NANDN U1346 ( .A(B[640]), .B(A[640]), .Z(n1538) );
  AND U1347 ( .A(n1539), .B(n1540), .Z(n1537) );
  NAND U1348 ( .A(n1541), .B(n1542), .Z(n1540) );
  NANDN U1349 ( .A(A[639]), .B(B[639]), .Z(n1542) );
  AND U1350 ( .A(n1543), .B(n1544), .Z(n1541) );
  NANDN U1351 ( .A(A[638]), .B(B[638]), .Z(n1544) );
  NAND U1352 ( .A(n1545), .B(n1546), .Z(n1543) );
  NANDN U1353 ( .A(B[638]), .B(A[638]), .Z(n1546) );
  AND U1354 ( .A(n1547), .B(n1548), .Z(n1545) );
  NAND U1355 ( .A(n1549), .B(n1550), .Z(n1548) );
  NANDN U1356 ( .A(A[637]), .B(B[637]), .Z(n1550) );
  AND U1357 ( .A(n1551), .B(n1552), .Z(n1549) );
  NANDN U1358 ( .A(A[636]), .B(B[636]), .Z(n1552) );
  NAND U1359 ( .A(n1553), .B(n1554), .Z(n1551) );
  NANDN U1360 ( .A(B[636]), .B(A[636]), .Z(n1554) );
  AND U1361 ( .A(n1555), .B(n1556), .Z(n1553) );
  NAND U1362 ( .A(n1557), .B(n1558), .Z(n1556) );
  NANDN U1363 ( .A(A[635]), .B(B[635]), .Z(n1558) );
  AND U1364 ( .A(n1559), .B(n1560), .Z(n1557) );
  NANDN U1365 ( .A(A[634]), .B(B[634]), .Z(n1560) );
  NAND U1366 ( .A(n1561), .B(n1562), .Z(n1559) );
  NANDN U1367 ( .A(B[634]), .B(A[634]), .Z(n1562) );
  AND U1368 ( .A(n1563), .B(n1564), .Z(n1561) );
  NAND U1369 ( .A(n1565), .B(n1566), .Z(n1564) );
  NANDN U1370 ( .A(A[633]), .B(B[633]), .Z(n1566) );
  AND U1371 ( .A(n1567), .B(n1568), .Z(n1565) );
  NANDN U1372 ( .A(A[632]), .B(B[632]), .Z(n1568) );
  NAND U1373 ( .A(n1569), .B(n1570), .Z(n1567) );
  NANDN U1374 ( .A(B[632]), .B(A[632]), .Z(n1570) );
  AND U1375 ( .A(n1571), .B(n1572), .Z(n1569) );
  NAND U1376 ( .A(n1573), .B(n1574), .Z(n1572) );
  NANDN U1377 ( .A(A[631]), .B(B[631]), .Z(n1574) );
  AND U1378 ( .A(n1575), .B(n1576), .Z(n1573) );
  NANDN U1379 ( .A(A[630]), .B(B[630]), .Z(n1576) );
  NAND U1380 ( .A(n1577), .B(n1578), .Z(n1575) );
  NANDN U1381 ( .A(B[630]), .B(A[630]), .Z(n1578) );
  AND U1382 ( .A(n1579), .B(n1580), .Z(n1577) );
  NAND U1383 ( .A(n1581), .B(n1582), .Z(n1580) );
  NANDN U1384 ( .A(A[629]), .B(B[629]), .Z(n1582) );
  AND U1385 ( .A(n1583), .B(n1584), .Z(n1581) );
  NANDN U1386 ( .A(A[628]), .B(B[628]), .Z(n1584) );
  NAND U1387 ( .A(n1585), .B(n1586), .Z(n1583) );
  NANDN U1388 ( .A(B[628]), .B(A[628]), .Z(n1586) );
  AND U1389 ( .A(n1587), .B(n1588), .Z(n1585) );
  NAND U1390 ( .A(n1589), .B(n1590), .Z(n1588) );
  NANDN U1391 ( .A(A[627]), .B(B[627]), .Z(n1590) );
  AND U1392 ( .A(n1591), .B(n1592), .Z(n1589) );
  NANDN U1393 ( .A(A[626]), .B(B[626]), .Z(n1592) );
  NAND U1394 ( .A(n1593), .B(n1594), .Z(n1591) );
  NANDN U1395 ( .A(B[626]), .B(A[626]), .Z(n1594) );
  AND U1396 ( .A(n1595), .B(n1596), .Z(n1593) );
  NAND U1397 ( .A(n1597), .B(n1598), .Z(n1596) );
  NANDN U1398 ( .A(A[625]), .B(B[625]), .Z(n1598) );
  AND U1399 ( .A(n1599), .B(n1600), .Z(n1597) );
  NANDN U1400 ( .A(A[624]), .B(B[624]), .Z(n1600) );
  NAND U1401 ( .A(n1601), .B(n1602), .Z(n1599) );
  NANDN U1402 ( .A(B[624]), .B(A[624]), .Z(n1602) );
  AND U1403 ( .A(n1603), .B(n1604), .Z(n1601) );
  NAND U1404 ( .A(n1605), .B(n1606), .Z(n1604) );
  NANDN U1405 ( .A(A[623]), .B(B[623]), .Z(n1606) );
  AND U1406 ( .A(n1607), .B(n1608), .Z(n1605) );
  NANDN U1407 ( .A(A[622]), .B(B[622]), .Z(n1608) );
  NAND U1408 ( .A(n1609), .B(n1610), .Z(n1607) );
  NANDN U1409 ( .A(B[622]), .B(A[622]), .Z(n1610) );
  AND U1410 ( .A(n1611), .B(n1612), .Z(n1609) );
  NAND U1411 ( .A(n1613), .B(n1614), .Z(n1612) );
  NANDN U1412 ( .A(A[621]), .B(B[621]), .Z(n1614) );
  AND U1413 ( .A(n1615), .B(n1616), .Z(n1613) );
  NANDN U1414 ( .A(A[620]), .B(B[620]), .Z(n1616) );
  NAND U1415 ( .A(n1617), .B(n1618), .Z(n1615) );
  NANDN U1416 ( .A(B[620]), .B(A[620]), .Z(n1618) );
  AND U1417 ( .A(n1619), .B(n1620), .Z(n1617) );
  NAND U1418 ( .A(n1621), .B(n1622), .Z(n1620) );
  NANDN U1419 ( .A(A[619]), .B(B[619]), .Z(n1622) );
  AND U1420 ( .A(n1623), .B(n1624), .Z(n1621) );
  NANDN U1421 ( .A(A[618]), .B(B[618]), .Z(n1624) );
  NAND U1422 ( .A(n1625), .B(n1626), .Z(n1623) );
  NANDN U1423 ( .A(B[618]), .B(A[618]), .Z(n1626) );
  AND U1424 ( .A(n1627), .B(n1628), .Z(n1625) );
  NAND U1425 ( .A(n1629), .B(n1630), .Z(n1628) );
  NANDN U1426 ( .A(A[617]), .B(B[617]), .Z(n1630) );
  AND U1427 ( .A(n1631), .B(n1632), .Z(n1629) );
  NANDN U1428 ( .A(A[616]), .B(B[616]), .Z(n1632) );
  NAND U1429 ( .A(n1633), .B(n1634), .Z(n1631) );
  NANDN U1430 ( .A(B[616]), .B(A[616]), .Z(n1634) );
  AND U1431 ( .A(n1635), .B(n1636), .Z(n1633) );
  NAND U1432 ( .A(n1637), .B(n1638), .Z(n1636) );
  NANDN U1433 ( .A(A[615]), .B(B[615]), .Z(n1638) );
  AND U1434 ( .A(n1639), .B(n1640), .Z(n1637) );
  NANDN U1435 ( .A(A[614]), .B(B[614]), .Z(n1640) );
  NAND U1436 ( .A(n1641), .B(n1642), .Z(n1639) );
  NANDN U1437 ( .A(B[614]), .B(A[614]), .Z(n1642) );
  AND U1438 ( .A(n1643), .B(n1644), .Z(n1641) );
  NAND U1439 ( .A(n1645), .B(n1646), .Z(n1644) );
  NANDN U1440 ( .A(A[613]), .B(B[613]), .Z(n1646) );
  AND U1441 ( .A(n1647), .B(n1648), .Z(n1645) );
  NANDN U1442 ( .A(A[612]), .B(B[612]), .Z(n1648) );
  NAND U1443 ( .A(n1649), .B(n1650), .Z(n1647) );
  NANDN U1444 ( .A(B[612]), .B(A[612]), .Z(n1650) );
  AND U1445 ( .A(n1651), .B(n1652), .Z(n1649) );
  NAND U1446 ( .A(n1653), .B(n1654), .Z(n1652) );
  NANDN U1447 ( .A(A[611]), .B(B[611]), .Z(n1654) );
  AND U1448 ( .A(n1655), .B(n1656), .Z(n1653) );
  NANDN U1449 ( .A(A[610]), .B(B[610]), .Z(n1656) );
  NAND U1450 ( .A(n1657), .B(n1658), .Z(n1655) );
  NANDN U1451 ( .A(B[610]), .B(A[610]), .Z(n1658) );
  AND U1452 ( .A(n1659), .B(n1660), .Z(n1657) );
  NAND U1453 ( .A(n1661), .B(n1662), .Z(n1660) );
  NANDN U1454 ( .A(A[609]), .B(B[609]), .Z(n1662) );
  AND U1455 ( .A(n1663), .B(n1664), .Z(n1661) );
  NANDN U1456 ( .A(A[608]), .B(B[608]), .Z(n1664) );
  NAND U1457 ( .A(n1665), .B(n1666), .Z(n1663) );
  NANDN U1458 ( .A(B[608]), .B(A[608]), .Z(n1666) );
  AND U1459 ( .A(n1667), .B(n1668), .Z(n1665) );
  NAND U1460 ( .A(n1669), .B(n1670), .Z(n1668) );
  NANDN U1461 ( .A(A[607]), .B(B[607]), .Z(n1670) );
  AND U1462 ( .A(n1671), .B(n1672), .Z(n1669) );
  NANDN U1463 ( .A(A[606]), .B(B[606]), .Z(n1672) );
  NAND U1464 ( .A(n1673), .B(n1674), .Z(n1671) );
  NANDN U1465 ( .A(B[606]), .B(A[606]), .Z(n1674) );
  AND U1466 ( .A(n1675), .B(n1676), .Z(n1673) );
  NAND U1467 ( .A(n1677), .B(n1678), .Z(n1676) );
  NANDN U1468 ( .A(A[605]), .B(B[605]), .Z(n1678) );
  AND U1469 ( .A(n1679), .B(n1680), .Z(n1677) );
  NANDN U1470 ( .A(A[604]), .B(B[604]), .Z(n1680) );
  NAND U1471 ( .A(n1681), .B(n1682), .Z(n1679) );
  NANDN U1472 ( .A(B[604]), .B(A[604]), .Z(n1682) );
  AND U1473 ( .A(n1683), .B(n1684), .Z(n1681) );
  NAND U1474 ( .A(n1685), .B(n1686), .Z(n1684) );
  NANDN U1475 ( .A(A[603]), .B(B[603]), .Z(n1686) );
  AND U1476 ( .A(n1687), .B(n1688), .Z(n1685) );
  NANDN U1477 ( .A(A[602]), .B(B[602]), .Z(n1688) );
  NAND U1478 ( .A(n1689), .B(n1690), .Z(n1687) );
  NANDN U1479 ( .A(B[602]), .B(A[602]), .Z(n1690) );
  AND U1480 ( .A(n1691), .B(n1692), .Z(n1689) );
  NAND U1481 ( .A(n1693), .B(n1694), .Z(n1692) );
  NANDN U1482 ( .A(A[601]), .B(B[601]), .Z(n1694) );
  AND U1483 ( .A(n1695), .B(n1696), .Z(n1693) );
  NANDN U1484 ( .A(A[600]), .B(B[600]), .Z(n1696) );
  NAND U1485 ( .A(n1697), .B(n1698), .Z(n1695) );
  NANDN U1486 ( .A(B[600]), .B(A[600]), .Z(n1698) );
  AND U1487 ( .A(n1699), .B(n1700), .Z(n1697) );
  NAND U1488 ( .A(n1701), .B(n1702), .Z(n1700) );
  NANDN U1489 ( .A(A[599]), .B(B[599]), .Z(n1702) );
  AND U1490 ( .A(n1703), .B(n1704), .Z(n1701) );
  NANDN U1491 ( .A(A[598]), .B(B[598]), .Z(n1704) );
  NAND U1492 ( .A(n1705), .B(n1706), .Z(n1703) );
  NANDN U1493 ( .A(B[598]), .B(A[598]), .Z(n1706) );
  AND U1494 ( .A(n1707), .B(n1708), .Z(n1705) );
  NAND U1495 ( .A(n1709), .B(n1710), .Z(n1708) );
  NANDN U1496 ( .A(A[597]), .B(B[597]), .Z(n1710) );
  AND U1497 ( .A(n1711), .B(n1712), .Z(n1709) );
  NANDN U1498 ( .A(A[596]), .B(B[596]), .Z(n1712) );
  NAND U1499 ( .A(n1713), .B(n1714), .Z(n1711) );
  NANDN U1500 ( .A(B[596]), .B(A[596]), .Z(n1714) );
  AND U1501 ( .A(n1715), .B(n1716), .Z(n1713) );
  NAND U1502 ( .A(n1717), .B(n1718), .Z(n1716) );
  NANDN U1503 ( .A(A[595]), .B(B[595]), .Z(n1718) );
  AND U1504 ( .A(n1719), .B(n1720), .Z(n1717) );
  NANDN U1505 ( .A(A[594]), .B(B[594]), .Z(n1720) );
  NAND U1506 ( .A(n1721), .B(n1722), .Z(n1719) );
  NANDN U1507 ( .A(B[594]), .B(A[594]), .Z(n1722) );
  AND U1508 ( .A(n1723), .B(n1724), .Z(n1721) );
  NAND U1509 ( .A(n1725), .B(n1726), .Z(n1724) );
  NANDN U1510 ( .A(A[593]), .B(B[593]), .Z(n1726) );
  AND U1511 ( .A(n1727), .B(n1728), .Z(n1725) );
  NANDN U1512 ( .A(A[592]), .B(B[592]), .Z(n1728) );
  NAND U1513 ( .A(n1729), .B(n1730), .Z(n1727) );
  NANDN U1514 ( .A(B[592]), .B(A[592]), .Z(n1730) );
  AND U1515 ( .A(n1731), .B(n1732), .Z(n1729) );
  NAND U1516 ( .A(n1733), .B(n1734), .Z(n1732) );
  NANDN U1517 ( .A(A[591]), .B(B[591]), .Z(n1734) );
  AND U1518 ( .A(n1735), .B(n1736), .Z(n1733) );
  NANDN U1519 ( .A(A[590]), .B(B[590]), .Z(n1736) );
  NAND U1520 ( .A(n1737), .B(n1738), .Z(n1735) );
  NANDN U1521 ( .A(B[590]), .B(A[590]), .Z(n1738) );
  AND U1522 ( .A(n1739), .B(n1740), .Z(n1737) );
  NAND U1523 ( .A(n1741), .B(n1742), .Z(n1740) );
  NANDN U1524 ( .A(A[589]), .B(B[589]), .Z(n1742) );
  AND U1525 ( .A(n1743), .B(n1744), .Z(n1741) );
  NANDN U1526 ( .A(A[588]), .B(B[588]), .Z(n1744) );
  NAND U1527 ( .A(n1745), .B(n1746), .Z(n1743) );
  NANDN U1528 ( .A(B[588]), .B(A[588]), .Z(n1746) );
  AND U1529 ( .A(n1747), .B(n1748), .Z(n1745) );
  NAND U1530 ( .A(n1749), .B(n1750), .Z(n1748) );
  NANDN U1531 ( .A(A[587]), .B(B[587]), .Z(n1750) );
  AND U1532 ( .A(n1751), .B(n1752), .Z(n1749) );
  NANDN U1533 ( .A(A[586]), .B(B[586]), .Z(n1752) );
  NAND U1534 ( .A(n1753), .B(n1754), .Z(n1751) );
  NANDN U1535 ( .A(B[586]), .B(A[586]), .Z(n1754) );
  AND U1536 ( .A(n1755), .B(n1756), .Z(n1753) );
  NAND U1537 ( .A(n1757), .B(n1758), .Z(n1756) );
  NANDN U1538 ( .A(A[585]), .B(B[585]), .Z(n1758) );
  AND U1539 ( .A(n1759), .B(n1760), .Z(n1757) );
  NANDN U1540 ( .A(A[584]), .B(B[584]), .Z(n1760) );
  NAND U1541 ( .A(n1761), .B(n1762), .Z(n1759) );
  NANDN U1542 ( .A(B[584]), .B(A[584]), .Z(n1762) );
  AND U1543 ( .A(n1763), .B(n1764), .Z(n1761) );
  NAND U1544 ( .A(n1765), .B(n1766), .Z(n1764) );
  NANDN U1545 ( .A(A[583]), .B(B[583]), .Z(n1766) );
  AND U1546 ( .A(n1767), .B(n1768), .Z(n1765) );
  NANDN U1547 ( .A(A[582]), .B(B[582]), .Z(n1768) );
  NAND U1548 ( .A(n1769), .B(n1770), .Z(n1767) );
  NANDN U1549 ( .A(B[582]), .B(A[582]), .Z(n1770) );
  AND U1550 ( .A(n1771), .B(n1772), .Z(n1769) );
  NAND U1551 ( .A(n1773), .B(n1774), .Z(n1772) );
  NANDN U1552 ( .A(A[581]), .B(B[581]), .Z(n1774) );
  AND U1553 ( .A(n1775), .B(n1776), .Z(n1773) );
  NANDN U1554 ( .A(A[580]), .B(B[580]), .Z(n1776) );
  NAND U1555 ( .A(n1777), .B(n1778), .Z(n1775) );
  NANDN U1556 ( .A(B[580]), .B(A[580]), .Z(n1778) );
  AND U1557 ( .A(n1779), .B(n1780), .Z(n1777) );
  NAND U1558 ( .A(n1781), .B(n1782), .Z(n1780) );
  NANDN U1559 ( .A(A[579]), .B(B[579]), .Z(n1782) );
  AND U1560 ( .A(n1783), .B(n1784), .Z(n1781) );
  NANDN U1561 ( .A(A[578]), .B(B[578]), .Z(n1784) );
  NAND U1562 ( .A(n1785), .B(n1786), .Z(n1783) );
  NANDN U1563 ( .A(B[578]), .B(A[578]), .Z(n1786) );
  AND U1564 ( .A(n1787), .B(n1788), .Z(n1785) );
  NAND U1565 ( .A(n1789), .B(n1790), .Z(n1788) );
  NANDN U1566 ( .A(A[577]), .B(B[577]), .Z(n1790) );
  AND U1567 ( .A(n1791), .B(n1792), .Z(n1789) );
  NANDN U1568 ( .A(A[576]), .B(B[576]), .Z(n1792) );
  NAND U1569 ( .A(n1793), .B(n1794), .Z(n1791) );
  NANDN U1570 ( .A(B[576]), .B(A[576]), .Z(n1794) );
  AND U1571 ( .A(n1795), .B(n1796), .Z(n1793) );
  NAND U1572 ( .A(n1797), .B(n1798), .Z(n1796) );
  NANDN U1573 ( .A(A[575]), .B(B[575]), .Z(n1798) );
  AND U1574 ( .A(n1799), .B(n1800), .Z(n1797) );
  NANDN U1575 ( .A(A[574]), .B(B[574]), .Z(n1800) );
  NAND U1576 ( .A(n1801), .B(n1802), .Z(n1799) );
  NANDN U1577 ( .A(B[574]), .B(A[574]), .Z(n1802) );
  AND U1578 ( .A(n1803), .B(n1804), .Z(n1801) );
  NAND U1579 ( .A(n1805), .B(n1806), .Z(n1804) );
  NANDN U1580 ( .A(A[573]), .B(B[573]), .Z(n1806) );
  AND U1581 ( .A(n1807), .B(n1808), .Z(n1805) );
  NANDN U1582 ( .A(A[572]), .B(B[572]), .Z(n1808) );
  NAND U1583 ( .A(n1809), .B(n1810), .Z(n1807) );
  NANDN U1584 ( .A(B[572]), .B(A[572]), .Z(n1810) );
  AND U1585 ( .A(n1811), .B(n1812), .Z(n1809) );
  NAND U1586 ( .A(n1813), .B(n1814), .Z(n1812) );
  NANDN U1587 ( .A(A[571]), .B(B[571]), .Z(n1814) );
  AND U1588 ( .A(n1815), .B(n1816), .Z(n1813) );
  NANDN U1589 ( .A(A[570]), .B(B[570]), .Z(n1816) );
  NAND U1590 ( .A(n1817), .B(n1818), .Z(n1815) );
  NANDN U1591 ( .A(B[570]), .B(A[570]), .Z(n1818) );
  AND U1592 ( .A(n1819), .B(n1820), .Z(n1817) );
  NAND U1593 ( .A(n1821), .B(n1822), .Z(n1820) );
  NANDN U1594 ( .A(A[569]), .B(B[569]), .Z(n1822) );
  AND U1595 ( .A(n1823), .B(n1824), .Z(n1821) );
  NANDN U1596 ( .A(A[568]), .B(B[568]), .Z(n1824) );
  NAND U1597 ( .A(n1825), .B(n1826), .Z(n1823) );
  NANDN U1598 ( .A(B[568]), .B(A[568]), .Z(n1826) );
  AND U1599 ( .A(n1827), .B(n1828), .Z(n1825) );
  NAND U1600 ( .A(n1829), .B(n1830), .Z(n1828) );
  NANDN U1601 ( .A(A[567]), .B(B[567]), .Z(n1830) );
  AND U1602 ( .A(n1831), .B(n1832), .Z(n1829) );
  NANDN U1603 ( .A(A[566]), .B(B[566]), .Z(n1832) );
  NAND U1604 ( .A(n1833), .B(n1834), .Z(n1831) );
  NANDN U1605 ( .A(B[566]), .B(A[566]), .Z(n1834) );
  AND U1606 ( .A(n1835), .B(n1836), .Z(n1833) );
  NAND U1607 ( .A(n1837), .B(n1838), .Z(n1836) );
  NANDN U1608 ( .A(A[565]), .B(B[565]), .Z(n1838) );
  AND U1609 ( .A(n1839), .B(n1840), .Z(n1837) );
  NANDN U1610 ( .A(A[564]), .B(B[564]), .Z(n1840) );
  NAND U1611 ( .A(n1841), .B(n1842), .Z(n1839) );
  NANDN U1612 ( .A(B[564]), .B(A[564]), .Z(n1842) );
  AND U1613 ( .A(n1843), .B(n1844), .Z(n1841) );
  NAND U1614 ( .A(n1845), .B(n1846), .Z(n1844) );
  NANDN U1615 ( .A(A[563]), .B(B[563]), .Z(n1846) );
  AND U1616 ( .A(n1847), .B(n1848), .Z(n1845) );
  NANDN U1617 ( .A(A[562]), .B(B[562]), .Z(n1848) );
  NAND U1618 ( .A(n1849), .B(n1850), .Z(n1847) );
  NANDN U1619 ( .A(B[562]), .B(A[562]), .Z(n1850) );
  AND U1620 ( .A(n1851), .B(n1852), .Z(n1849) );
  NAND U1621 ( .A(n1853), .B(n1854), .Z(n1852) );
  NANDN U1622 ( .A(A[561]), .B(B[561]), .Z(n1854) );
  AND U1623 ( .A(n1855), .B(n1856), .Z(n1853) );
  NANDN U1624 ( .A(A[560]), .B(B[560]), .Z(n1856) );
  NAND U1625 ( .A(n1857), .B(n1858), .Z(n1855) );
  NANDN U1626 ( .A(B[560]), .B(A[560]), .Z(n1858) );
  AND U1627 ( .A(n1859), .B(n1860), .Z(n1857) );
  NAND U1628 ( .A(n1861), .B(n1862), .Z(n1860) );
  NANDN U1629 ( .A(A[559]), .B(B[559]), .Z(n1862) );
  AND U1630 ( .A(n1863), .B(n1864), .Z(n1861) );
  NANDN U1631 ( .A(A[558]), .B(B[558]), .Z(n1864) );
  NAND U1632 ( .A(n1865), .B(n1866), .Z(n1863) );
  NANDN U1633 ( .A(B[558]), .B(A[558]), .Z(n1866) );
  AND U1634 ( .A(n1867), .B(n1868), .Z(n1865) );
  NAND U1635 ( .A(n1869), .B(n1870), .Z(n1868) );
  NANDN U1636 ( .A(A[557]), .B(B[557]), .Z(n1870) );
  AND U1637 ( .A(n1871), .B(n1872), .Z(n1869) );
  NANDN U1638 ( .A(A[556]), .B(B[556]), .Z(n1872) );
  NAND U1639 ( .A(n1873), .B(n1874), .Z(n1871) );
  NANDN U1640 ( .A(B[556]), .B(A[556]), .Z(n1874) );
  AND U1641 ( .A(n1875), .B(n1876), .Z(n1873) );
  NAND U1642 ( .A(n1877), .B(n1878), .Z(n1876) );
  NANDN U1643 ( .A(A[555]), .B(B[555]), .Z(n1878) );
  AND U1644 ( .A(n1879), .B(n1880), .Z(n1877) );
  NANDN U1645 ( .A(A[554]), .B(B[554]), .Z(n1880) );
  NAND U1646 ( .A(n1881), .B(n1882), .Z(n1879) );
  NANDN U1647 ( .A(B[554]), .B(A[554]), .Z(n1882) );
  AND U1648 ( .A(n1883), .B(n1884), .Z(n1881) );
  NAND U1649 ( .A(n1885), .B(n1886), .Z(n1884) );
  NANDN U1650 ( .A(A[553]), .B(B[553]), .Z(n1886) );
  AND U1651 ( .A(n1887), .B(n1888), .Z(n1885) );
  NANDN U1652 ( .A(A[552]), .B(B[552]), .Z(n1888) );
  NAND U1653 ( .A(n1889), .B(n1890), .Z(n1887) );
  NANDN U1654 ( .A(B[552]), .B(A[552]), .Z(n1890) );
  AND U1655 ( .A(n1891), .B(n1892), .Z(n1889) );
  NAND U1656 ( .A(n1893), .B(n1894), .Z(n1892) );
  NANDN U1657 ( .A(A[551]), .B(B[551]), .Z(n1894) );
  AND U1658 ( .A(n1895), .B(n1896), .Z(n1893) );
  NANDN U1659 ( .A(A[550]), .B(B[550]), .Z(n1896) );
  NAND U1660 ( .A(n1897), .B(n1898), .Z(n1895) );
  NANDN U1661 ( .A(B[550]), .B(A[550]), .Z(n1898) );
  AND U1662 ( .A(n1899), .B(n1900), .Z(n1897) );
  NAND U1663 ( .A(n1901), .B(n1902), .Z(n1900) );
  NANDN U1664 ( .A(A[549]), .B(B[549]), .Z(n1902) );
  AND U1665 ( .A(n1903), .B(n1904), .Z(n1901) );
  NANDN U1666 ( .A(A[548]), .B(B[548]), .Z(n1904) );
  NAND U1667 ( .A(n1905), .B(n1906), .Z(n1903) );
  NANDN U1668 ( .A(B[548]), .B(A[548]), .Z(n1906) );
  AND U1669 ( .A(n1907), .B(n1908), .Z(n1905) );
  NAND U1670 ( .A(n1909), .B(n1910), .Z(n1908) );
  NANDN U1671 ( .A(A[547]), .B(B[547]), .Z(n1910) );
  AND U1672 ( .A(n1911), .B(n1912), .Z(n1909) );
  NANDN U1673 ( .A(A[546]), .B(B[546]), .Z(n1912) );
  NAND U1674 ( .A(n1913), .B(n1914), .Z(n1911) );
  NANDN U1675 ( .A(B[546]), .B(A[546]), .Z(n1914) );
  AND U1676 ( .A(n1915), .B(n1916), .Z(n1913) );
  NAND U1677 ( .A(n1917), .B(n1918), .Z(n1916) );
  NANDN U1678 ( .A(A[545]), .B(B[545]), .Z(n1918) );
  AND U1679 ( .A(n1919), .B(n1920), .Z(n1917) );
  NANDN U1680 ( .A(A[544]), .B(B[544]), .Z(n1920) );
  NAND U1681 ( .A(n1921), .B(n1922), .Z(n1919) );
  NANDN U1682 ( .A(B[544]), .B(A[544]), .Z(n1922) );
  AND U1683 ( .A(n1923), .B(n1924), .Z(n1921) );
  NAND U1684 ( .A(n1925), .B(n1926), .Z(n1924) );
  NANDN U1685 ( .A(A[543]), .B(B[543]), .Z(n1926) );
  AND U1686 ( .A(n1927), .B(n1928), .Z(n1925) );
  NANDN U1687 ( .A(A[542]), .B(B[542]), .Z(n1928) );
  NAND U1688 ( .A(n1929), .B(n1930), .Z(n1927) );
  NANDN U1689 ( .A(B[542]), .B(A[542]), .Z(n1930) );
  AND U1690 ( .A(n1931), .B(n1932), .Z(n1929) );
  NAND U1691 ( .A(n1933), .B(n1934), .Z(n1932) );
  NANDN U1692 ( .A(A[541]), .B(B[541]), .Z(n1934) );
  AND U1693 ( .A(n1935), .B(n1936), .Z(n1933) );
  NANDN U1694 ( .A(A[540]), .B(B[540]), .Z(n1936) );
  NAND U1695 ( .A(n1937), .B(n1938), .Z(n1935) );
  NANDN U1696 ( .A(B[540]), .B(A[540]), .Z(n1938) );
  AND U1697 ( .A(n1939), .B(n1940), .Z(n1937) );
  NAND U1698 ( .A(n1941), .B(n1942), .Z(n1940) );
  NANDN U1699 ( .A(A[539]), .B(B[539]), .Z(n1942) );
  AND U1700 ( .A(n1943), .B(n1944), .Z(n1941) );
  NANDN U1701 ( .A(A[538]), .B(B[538]), .Z(n1944) );
  NAND U1702 ( .A(n1945), .B(n1946), .Z(n1943) );
  NANDN U1703 ( .A(B[538]), .B(A[538]), .Z(n1946) );
  AND U1704 ( .A(n1947), .B(n1948), .Z(n1945) );
  NAND U1705 ( .A(n1949), .B(n1950), .Z(n1948) );
  NANDN U1706 ( .A(A[537]), .B(B[537]), .Z(n1950) );
  AND U1707 ( .A(n1951), .B(n1952), .Z(n1949) );
  NANDN U1708 ( .A(A[536]), .B(B[536]), .Z(n1952) );
  NAND U1709 ( .A(n1953), .B(n1954), .Z(n1951) );
  NANDN U1710 ( .A(B[536]), .B(A[536]), .Z(n1954) );
  AND U1711 ( .A(n1955), .B(n1956), .Z(n1953) );
  NAND U1712 ( .A(n1957), .B(n1958), .Z(n1956) );
  NANDN U1713 ( .A(A[535]), .B(B[535]), .Z(n1958) );
  AND U1714 ( .A(n1959), .B(n1960), .Z(n1957) );
  NANDN U1715 ( .A(A[534]), .B(B[534]), .Z(n1960) );
  NAND U1716 ( .A(n1961), .B(n1962), .Z(n1959) );
  NANDN U1717 ( .A(B[534]), .B(A[534]), .Z(n1962) );
  AND U1718 ( .A(n1963), .B(n1964), .Z(n1961) );
  NAND U1719 ( .A(n1965), .B(n1966), .Z(n1964) );
  NANDN U1720 ( .A(A[533]), .B(B[533]), .Z(n1966) );
  AND U1721 ( .A(n1967), .B(n1968), .Z(n1965) );
  NANDN U1722 ( .A(A[532]), .B(B[532]), .Z(n1968) );
  NAND U1723 ( .A(n1969), .B(n1970), .Z(n1967) );
  NANDN U1724 ( .A(B[532]), .B(A[532]), .Z(n1970) );
  AND U1725 ( .A(n1971), .B(n1972), .Z(n1969) );
  NAND U1726 ( .A(n1973), .B(n1974), .Z(n1972) );
  NANDN U1727 ( .A(A[531]), .B(B[531]), .Z(n1974) );
  AND U1728 ( .A(n1975), .B(n1976), .Z(n1973) );
  NANDN U1729 ( .A(A[530]), .B(B[530]), .Z(n1976) );
  NAND U1730 ( .A(n1977), .B(n1978), .Z(n1975) );
  NANDN U1731 ( .A(B[530]), .B(A[530]), .Z(n1978) );
  AND U1732 ( .A(n1979), .B(n1980), .Z(n1977) );
  NAND U1733 ( .A(n1981), .B(n1982), .Z(n1980) );
  NANDN U1734 ( .A(A[529]), .B(B[529]), .Z(n1982) );
  AND U1735 ( .A(n1983), .B(n1984), .Z(n1981) );
  NANDN U1736 ( .A(A[528]), .B(B[528]), .Z(n1984) );
  NAND U1737 ( .A(n1985), .B(n1986), .Z(n1983) );
  NANDN U1738 ( .A(B[528]), .B(A[528]), .Z(n1986) );
  AND U1739 ( .A(n1987), .B(n1988), .Z(n1985) );
  NAND U1740 ( .A(n1989), .B(n1990), .Z(n1988) );
  NANDN U1741 ( .A(A[527]), .B(B[527]), .Z(n1990) );
  AND U1742 ( .A(n1991), .B(n1992), .Z(n1989) );
  NANDN U1743 ( .A(A[526]), .B(B[526]), .Z(n1992) );
  NAND U1744 ( .A(n1993), .B(n1994), .Z(n1991) );
  NANDN U1745 ( .A(B[526]), .B(A[526]), .Z(n1994) );
  AND U1746 ( .A(n1995), .B(n1996), .Z(n1993) );
  NAND U1747 ( .A(n1997), .B(n1998), .Z(n1996) );
  NANDN U1748 ( .A(A[525]), .B(B[525]), .Z(n1998) );
  AND U1749 ( .A(n1999), .B(n2000), .Z(n1997) );
  NANDN U1750 ( .A(A[524]), .B(B[524]), .Z(n2000) );
  NAND U1751 ( .A(n2001), .B(n2002), .Z(n1999) );
  NANDN U1752 ( .A(B[524]), .B(A[524]), .Z(n2002) );
  AND U1753 ( .A(n2003), .B(n2004), .Z(n2001) );
  NAND U1754 ( .A(n2005), .B(n2006), .Z(n2004) );
  NANDN U1755 ( .A(A[523]), .B(B[523]), .Z(n2006) );
  AND U1756 ( .A(n2007), .B(n2008), .Z(n2005) );
  NANDN U1757 ( .A(A[522]), .B(B[522]), .Z(n2008) );
  NAND U1758 ( .A(n2009), .B(n2010), .Z(n2007) );
  NANDN U1759 ( .A(B[522]), .B(A[522]), .Z(n2010) );
  AND U1760 ( .A(n2011), .B(n2012), .Z(n2009) );
  NAND U1761 ( .A(n2013), .B(n2014), .Z(n2012) );
  NANDN U1762 ( .A(A[521]), .B(B[521]), .Z(n2014) );
  AND U1763 ( .A(n2015), .B(n2016), .Z(n2013) );
  NANDN U1764 ( .A(A[520]), .B(B[520]), .Z(n2016) );
  NAND U1765 ( .A(n2017), .B(n2018), .Z(n2015) );
  NANDN U1766 ( .A(B[520]), .B(A[520]), .Z(n2018) );
  AND U1767 ( .A(n2019), .B(n2020), .Z(n2017) );
  NAND U1768 ( .A(n2021), .B(n2022), .Z(n2020) );
  NANDN U1769 ( .A(A[519]), .B(B[519]), .Z(n2022) );
  AND U1770 ( .A(n2023), .B(n2024), .Z(n2021) );
  NANDN U1771 ( .A(A[518]), .B(B[518]), .Z(n2024) );
  NAND U1772 ( .A(n2025), .B(n2026), .Z(n2023) );
  NANDN U1773 ( .A(B[518]), .B(A[518]), .Z(n2026) );
  AND U1774 ( .A(n2027), .B(n2028), .Z(n2025) );
  NAND U1775 ( .A(n2029), .B(n2030), .Z(n2028) );
  NANDN U1776 ( .A(A[517]), .B(B[517]), .Z(n2030) );
  AND U1777 ( .A(n2031), .B(n2032), .Z(n2029) );
  NANDN U1778 ( .A(A[516]), .B(B[516]), .Z(n2032) );
  NAND U1779 ( .A(n2033), .B(n2034), .Z(n2031) );
  NANDN U1780 ( .A(B[516]), .B(A[516]), .Z(n2034) );
  AND U1781 ( .A(n2035), .B(n2036), .Z(n2033) );
  NAND U1782 ( .A(n2037), .B(n2038), .Z(n2036) );
  NANDN U1783 ( .A(A[515]), .B(B[515]), .Z(n2038) );
  AND U1784 ( .A(n2039), .B(n2040), .Z(n2037) );
  NANDN U1785 ( .A(A[514]), .B(B[514]), .Z(n2040) );
  NAND U1786 ( .A(n2041), .B(n2042), .Z(n2039) );
  NANDN U1787 ( .A(B[514]), .B(A[514]), .Z(n2042) );
  AND U1788 ( .A(n2043), .B(n2044), .Z(n2041) );
  NAND U1789 ( .A(n2045), .B(n2046), .Z(n2044) );
  NANDN U1790 ( .A(A[513]), .B(B[513]), .Z(n2046) );
  AND U1791 ( .A(n2047), .B(n2048), .Z(n2045) );
  NANDN U1792 ( .A(A[512]), .B(B[512]), .Z(n2048) );
  NAND U1793 ( .A(n2049), .B(n2050), .Z(n2047) );
  NANDN U1794 ( .A(B[512]), .B(A[512]), .Z(n2050) );
  AND U1795 ( .A(n2051), .B(n2052), .Z(n2049) );
  NAND U1796 ( .A(n2053), .B(n2054), .Z(n2052) );
  NANDN U1797 ( .A(A[511]), .B(B[511]), .Z(n2054) );
  AND U1798 ( .A(n2055), .B(n2056), .Z(n2053) );
  NANDN U1799 ( .A(A[510]), .B(B[510]), .Z(n2056) );
  NAND U1800 ( .A(n2057), .B(n2058), .Z(n2055) );
  NANDN U1801 ( .A(B[510]), .B(A[510]), .Z(n2058) );
  AND U1802 ( .A(n2059), .B(n2060), .Z(n2057) );
  NAND U1803 ( .A(n2061), .B(n2062), .Z(n2060) );
  NANDN U1804 ( .A(A[509]), .B(B[509]), .Z(n2062) );
  AND U1805 ( .A(n2063), .B(n2064), .Z(n2061) );
  NANDN U1806 ( .A(A[508]), .B(B[508]), .Z(n2064) );
  NAND U1807 ( .A(n2065), .B(n2066), .Z(n2063) );
  NANDN U1808 ( .A(B[508]), .B(A[508]), .Z(n2066) );
  AND U1809 ( .A(n2067), .B(n2068), .Z(n2065) );
  NAND U1810 ( .A(n2069), .B(n2070), .Z(n2068) );
  NANDN U1811 ( .A(A[507]), .B(B[507]), .Z(n2070) );
  AND U1812 ( .A(n2071), .B(n2072), .Z(n2069) );
  NANDN U1813 ( .A(A[506]), .B(B[506]), .Z(n2072) );
  NAND U1814 ( .A(n2073), .B(n2074), .Z(n2071) );
  NANDN U1815 ( .A(B[506]), .B(A[506]), .Z(n2074) );
  AND U1816 ( .A(n2075), .B(n2076), .Z(n2073) );
  NAND U1817 ( .A(n2077), .B(n2078), .Z(n2076) );
  NANDN U1818 ( .A(A[505]), .B(B[505]), .Z(n2078) );
  AND U1819 ( .A(n2079), .B(n2080), .Z(n2077) );
  NANDN U1820 ( .A(A[504]), .B(B[504]), .Z(n2080) );
  NAND U1821 ( .A(n2081), .B(n2082), .Z(n2079) );
  NANDN U1822 ( .A(B[504]), .B(A[504]), .Z(n2082) );
  AND U1823 ( .A(n2083), .B(n2084), .Z(n2081) );
  NAND U1824 ( .A(n2085), .B(n2086), .Z(n2084) );
  NANDN U1825 ( .A(A[503]), .B(B[503]), .Z(n2086) );
  AND U1826 ( .A(n2087), .B(n2088), .Z(n2085) );
  NANDN U1827 ( .A(A[502]), .B(B[502]), .Z(n2088) );
  NAND U1828 ( .A(n2089), .B(n2090), .Z(n2087) );
  NANDN U1829 ( .A(B[502]), .B(A[502]), .Z(n2090) );
  AND U1830 ( .A(n2091), .B(n2092), .Z(n2089) );
  NAND U1831 ( .A(n2093), .B(n2094), .Z(n2092) );
  NANDN U1832 ( .A(A[501]), .B(B[501]), .Z(n2094) );
  AND U1833 ( .A(n2095), .B(n2096), .Z(n2093) );
  NANDN U1834 ( .A(A[500]), .B(B[500]), .Z(n2096) );
  NAND U1835 ( .A(n2097), .B(n2098), .Z(n2095) );
  NANDN U1836 ( .A(B[500]), .B(A[500]), .Z(n2098) );
  AND U1837 ( .A(n2099), .B(n2100), .Z(n2097) );
  NAND U1838 ( .A(n2101), .B(n2102), .Z(n2100) );
  NANDN U1839 ( .A(A[499]), .B(B[499]), .Z(n2102) );
  AND U1840 ( .A(n2103), .B(n2104), .Z(n2101) );
  NANDN U1841 ( .A(A[498]), .B(B[498]), .Z(n2104) );
  NAND U1842 ( .A(n2105), .B(n2106), .Z(n2103) );
  NANDN U1843 ( .A(B[498]), .B(A[498]), .Z(n2106) );
  AND U1844 ( .A(n2107), .B(n2108), .Z(n2105) );
  NAND U1845 ( .A(n2109), .B(n2110), .Z(n2108) );
  NANDN U1846 ( .A(A[497]), .B(B[497]), .Z(n2110) );
  AND U1847 ( .A(n2111), .B(n2112), .Z(n2109) );
  NANDN U1848 ( .A(A[496]), .B(B[496]), .Z(n2112) );
  NAND U1849 ( .A(n2113), .B(n2114), .Z(n2111) );
  NANDN U1850 ( .A(B[496]), .B(A[496]), .Z(n2114) );
  AND U1851 ( .A(n2115), .B(n2116), .Z(n2113) );
  NAND U1852 ( .A(n2117), .B(n2118), .Z(n2116) );
  NANDN U1853 ( .A(A[495]), .B(B[495]), .Z(n2118) );
  AND U1854 ( .A(n2119), .B(n2120), .Z(n2117) );
  NANDN U1855 ( .A(A[494]), .B(B[494]), .Z(n2120) );
  NAND U1856 ( .A(n2121), .B(n2122), .Z(n2119) );
  NANDN U1857 ( .A(B[494]), .B(A[494]), .Z(n2122) );
  AND U1858 ( .A(n2123), .B(n2124), .Z(n2121) );
  NAND U1859 ( .A(n2125), .B(n2126), .Z(n2124) );
  NANDN U1860 ( .A(A[493]), .B(B[493]), .Z(n2126) );
  AND U1861 ( .A(n2127), .B(n2128), .Z(n2125) );
  NANDN U1862 ( .A(A[492]), .B(B[492]), .Z(n2128) );
  NAND U1863 ( .A(n2129), .B(n2130), .Z(n2127) );
  NANDN U1864 ( .A(B[492]), .B(A[492]), .Z(n2130) );
  AND U1865 ( .A(n2131), .B(n2132), .Z(n2129) );
  NAND U1866 ( .A(n2133), .B(n2134), .Z(n2132) );
  NANDN U1867 ( .A(A[491]), .B(B[491]), .Z(n2134) );
  AND U1868 ( .A(n2135), .B(n2136), .Z(n2133) );
  NANDN U1869 ( .A(A[490]), .B(B[490]), .Z(n2136) );
  NAND U1870 ( .A(n2137), .B(n2138), .Z(n2135) );
  NANDN U1871 ( .A(B[490]), .B(A[490]), .Z(n2138) );
  AND U1872 ( .A(n2139), .B(n2140), .Z(n2137) );
  NAND U1873 ( .A(n2141), .B(n2142), .Z(n2140) );
  NANDN U1874 ( .A(A[489]), .B(B[489]), .Z(n2142) );
  AND U1875 ( .A(n2143), .B(n2144), .Z(n2141) );
  NANDN U1876 ( .A(A[488]), .B(B[488]), .Z(n2144) );
  NAND U1877 ( .A(n2145), .B(n2146), .Z(n2143) );
  NANDN U1878 ( .A(B[488]), .B(A[488]), .Z(n2146) );
  AND U1879 ( .A(n2147), .B(n2148), .Z(n2145) );
  NAND U1880 ( .A(n2149), .B(n2150), .Z(n2148) );
  NANDN U1881 ( .A(A[487]), .B(B[487]), .Z(n2150) );
  AND U1882 ( .A(n2151), .B(n2152), .Z(n2149) );
  NANDN U1883 ( .A(A[486]), .B(B[486]), .Z(n2152) );
  NAND U1884 ( .A(n2153), .B(n2154), .Z(n2151) );
  NANDN U1885 ( .A(B[486]), .B(A[486]), .Z(n2154) );
  AND U1886 ( .A(n2155), .B(n2156), .Z(n2153) );
  NAND U1887 ( .A(n2157), .B(n2158), .Z(n2156) );
  NANDN U1888 ( .A(A[485]), .B(B[485]), .Z(n2158) );
  AND U1889 ( .A(n2159), .B(n2160), .Z(n2157) );
  NANDN U1890 ( .A(A[484]), .B(B[484]), .Z(n2160) );
  NAND U1891 ( .A(n2161), .B(n2162), .Z(n2159) );
  NANDN U1892 ( .A(B[484]), .B(A[484]), .Z(n2162) );
  AND U1893 ( .A(n2163), .B(n2164), .Z(n2161) );
  NAND U1894 ( .A(n2165), .B(n2166), .Z(n2164) );
  NANDN U1895 ( .A(A[483]), .B(B[483]), .Z(n2166) );
  AND U1896 ( .A(n2167), .B(n2168), .Z(n2165) );
  NANDN U1897 ( .A(A[482]), .B(B[482]), .Z(n2168) );
  NAND U1898 ( .A(n2169), .B(n2170), .Z(n2167) );
  NANDN U1899 ( .A(B[482]), .B(A[482]), .Z(n2170) );
  AND U1900 ( .A(n2171), .B(n2172), .Z(n2169) );
  NAND U1901 ( .A(n2173), .B(n2174), .Z(n2172) );
  NANDN U1902 ( .A(A[481]), .B(B[481]), .Z(n2174) );
  AND U1903 ( .A(n2175), .B(n2176), .Z(n2173) );
  NANDN U1904 ( .A(A[480]), .B(B[480]), .Z(n2176) );
  NAND U1905 ( .A(n2177), .B(n2178), .Z(n2175) );
  NANDN U1906 ( .A(B[480]), .B(A[480]), .Z(n2178) );
  AND U1907 ( .A(n2179), .B(n2180), .Z(n2177) );
  NAND U1908 ( .A(n2181), .B(n2182), .Z(n2180) );
  NANDN U1909 ( .A(A[479]), .B(B[479]), .Z(n2182) );
  AND U1910 ( .A(n2183), .B(n2184), .Z(n2181) );
  NANDN U1911 ( .A(A[478]), .B(B[478]), .Z(n2184) );
  NAND U1912 ( .A(n2185), .B(n2186), .Z(n2183) );
  NANDN U1913 ( .A(B[478]), .B(A[478]), .Z(n2186) );
  AND U1914 ( .A(n2187), .B(n2188), .Z(n2185) );
  NAND U1915 ( .A(n2189), .B(n2190), .Z(n2188) );
  NANDN U1916 ( .A(A[477]), .B(B[477]), .Z(n2190) );
  AND U1917 ( .A(n2191), .B(n2192), .Z(n2189) );
  NANDN U1918 ( .A(A[476]), .B(B[476]), .Z(n2192) );
  NAND U1919 ( .A(n2193), .B(n2194), .Z(n2191) );
  NANDN U1920 ( .A(B[476]), .B(A[476]), .Z(n2194) );
  AND U1921 ( .A(n2195), .B(n2196), .Z(n2193) );
  NAND U1922 ( .A(n2197), .B(n2198), .Z(n2196) );
  NANDN U1923 ( .A(A[475]), .B(B[475]), .Z(n2198) );
  AND U1924 ( .A(n2199), .B(n2200), .Z(n2197) );
  NANDN U1925 ( .A(A[474]), .B(B[474]), .Z(n2200) );
  NAND U1926 ( .A(n2201), .B(n2202), .Z(n2199) );
  NANDN U1927 ( .A(B[474]), .B(A[474]), .Z(n2202) );
  AND U1928 ( .A(n2203), .B(n2204), .Z(n2201) );
  NAND U1929 ( .A(n2205), .B(n2206), .Z(n2204) );
  NANDN U1930 ( .A(A[473]), .B(B[473]), .Z(n2206) );
  AND U1931 ( .A(n2207), .B(n2208), .Z(n2205) );
  NANDN U1932 ( .A(A[472]), .B(B[472]), .Z(n2208) );
  NAND U1933 ( .A(n2209), .B(n2210), .Z(n2207) );
  NANDN U1934 ( .A(B[472]), .B(A[472]), .Z(n2210) );
  AND U1935 ( .A(n2211), .B(n2212), .Z(n2209) );
  NAND U1936 ( .A(n2213), .B(n2214), .Z(n2212) );
  NANDN U1937 ( .A(A[471]), .B(B[471]), .Z(n2214) );
  AND U1938 ( .A(n2215), .B(n2216), .Z(n2213) );
  NANDN U1939 ( .A(A[470]), .B(B[470]), .Z(n2216) );
  NAND U1940 ( .A(n2217), .B(n2218), .Z(n2215) );
  NANDN U1941 ( .A(B[470]), .B(A[470]), .Z(n2218) );
  AND U1942 ( .A(n2219), .B(n2220), .Z(n2217) );
  NAND U1943 ( .A(n2221), .B(n2222), .Z(n2220) );
  NANDN U1944 ( .A(A[469]), .B(B[469]), .Z(n2222) );
  AND U1945 ( .A(n2223), .B(n2224), .Z(n2221) );
  NANDN U1946 ( .A(A[468]), .B(B[468]), .Z(n2224) );
  NAND U1947 ( .A(n2225), .B(n2226), .Z(n2223) );
  NANDN U1948 ( .A(B[468]), .B(A[468]), .Z(n2226) );
  AND U1949 ( .A(n2227), .B(n2228), .Z(n2225) );
  NAND U1950 ( .A(n2229), .B(n2230), .Z(n2228) );
  NANDN U1951 ( .A(A[467]), .B(B[467]), .Z(n2230) );
  AND U1952 ( .A(n2231), .B(n2232), .Z(n2229) );
  NANDN U1953 ( .A(A[466]), .B(B[466]), .Z(n2232) );
  NAND U1954 ( .A(n2233), .B(n2234), .Z(n2231) );
  NANDN U1955 ( .A(B[466]), .B(A[466]), .Z(n2234) );
  AND U1956 ( .A(n2235), .B(n2236), .Z(n2233) );
  NAND U1957 ( .A(n2237), .B(n2238), .Z(n2236) );
  NANDN U1958 ( .A(A[465]), .B(B[465]), .Z(n2238) );
  AND U1959 ( .A(n2239), .B(n2240), .Z(n2237) );
  NANDN U1960 ( .A(A[464]), .B(B[464]), .Z(n2240) );
  NAND U1961 ( .A(n2241), .B(n2242), .Z(n2239) );
  NANDN U1962 ( .A(B[464]), .B(A[464]), .Z(n2242) );
  AND U1963 ( .A(n2243), .B(n2244), .Z(n2241) );
  NAND U1964 ( .A(n2245), .B(n2246), .Z(n2244) );
  NANDN U1965 ( .A(A[463]), .B(B[463]), .Z(n2246) );
  AND U1966 ( .A(n2247), .B(n2248), .Z(n2245) );
  NANDN U1967 ( .A(A[462]), .B(B[462]), .Z(n2248) );
  NAND U1968 ( .A(n2249), .B(n2250), .Z(n2247) );
  NANDN U1969 ( .A(B[462]), .B(A[462]), .Z(n2250) );
  AND U1970 ( .A(n2251), .B(n2252), .Z(n2249) );
  NAND U1971 ( .A(n2253), .B(n2254), .Z(n2252) );
  NANDN U1972 ( .A(A[461]), .B(B[461]), .Z(n2254) );
  AND U1973 ( .A(n2255), .B(n2256), .Z(n2253) );
  NANDN U1974 ( .A(A[460]), .B(B[460]), .Z(n2256) );
  NAND U1975 ( .A(n2257), .B(n2258), .Z(n2255) );
  NANDN U1976 ( .A(B[460]), .B(A[460]), .Z(n2258) );
  AND U1977 ( .A(n2259), .B(n2260), .Z(n2257) );
  NAND U1978 ( .A(n2261), .B(n2262), .Z(n2260) );
  NANDN U1979 ( .A(A[459]), .B(B[459]), .Z(n2262) );
  AND U1980 ( .A(n2263), .B(n2264), .Z(n2261) );
  NANDN U1981 ( .A(A[458]), .B(B[458]), .Z(n2264) );
  NAND U1982 ( .A(n2265), .B(n2266), .Z(n2263) );
  NANDN U1983 ( .A(B[458]), .B(A[458]), .Z(n2266) );
  AND U1984 ( .A(n2267), .B(n2268), .Z(n2265) );
  NAND U1985 ( .A(n2269), .B(n2270), .Z(n2268) );
  NANDN U1986 ( .A(A[457]), .B(B[457]), .Z(n2270) );
  AND U1987 ( .A(n2271), .B(n2272), .Z(n2269) );
  NANDN U1988 ( .A(A[456]), .B(B[456]), .Z(n2272) );
  NAND U1989 ( .A(n2273), .B(n2274), .Z(n2271) );
  NANDN U1990 ( .A(B[456]), .B(A[456]), .Z(n2274) );
  AND U1991 ( .A(n2275), .B(n2276), .Z(n2273) );
  NAND U1992 ( .A(n2277), .B(n2278), .Z(n2276) );
  NANDN U1993 ( .A(A[455]), .B(B[455]), .Z(n2278) );
  AND U1994 ( .A(n2279), .B(n2280), .Z(n2277) );
  NANDN U1995 ( .A(A[454]), .B(B[454]), .Z(n2280) );
  NAND U1996 ( .A(n2281), .B(n2282), .Z(n2279) );
  NANDN U1997 ( .A(B[454]), .B(A[454]), .Z(n2282) );
  AND U1998 ( .A(n2283), .B(n2284), .Z(n2281) );
  NAND U1999 ( .A(n2285), .B(n2286), .Z(n2284) );
  NANDN U2000 ( .A(A[453]), .B(B[453]), .Z(n2286) );
  AND U2001 ( .A(n2287), .B(n2288), .Z(n2285) );
  NANDN U2002 ( .A(A[452]), .B(B[452]), .Z(n2288) );
  NAND U2003 ( .A(n2289), .B(n2290), .Z(n2287) );
  NANDN U2004 ( .A(B[452]), .B(A[452]), .Z(n2290) );
  AND U2005 ( .A(n2291), .B(n2292), .Z(n2289) );
  NAND U2006 ( .A(n2293), .B(n2294), .Z(n2292) );
  NANDN U2007 ( .A(A[451]), .B(B[451]), .Z(n2294) );
  AND U2008 ( .A(n2295), .B(n2296), .Z(n2293) );
  NANDN U2009 ( .A(A[450]), .B(B[450]), .Z(n2296) );
  NAND U2010 ( .A(n2297), .B(n2298), .Z(n2295) );
  NANDN U2011 ( .A(B[450]), .B(A[450]), .Z(n2298) );
  AND U2012 ( .A(n2299), .B(n2300), .Z(n2297) );
  NAND U2013 ( .A(n2301), .B(n2302), .Z(n2300) );
  NANDN U2014 ( .A(A[449]), .B(B[449]), .Z(n2302) );
  AND U2015 ( .A(n2303), .B(n2304), .Z(n2301) );
  NANDN U2016 ( .A(A[448]), .B(B[448]), .Z(n2304) );
  NAND U2017 ( .A(n2305), .B(n2306), .Z(n2303) );
  NANDN U2018 ( .A(B[448]), .B(A[448]), .Z(n2306) );
  AND U2019 ( .A(n2307), .B(n2308), .Z(n2305) );
  NAND U2020 ( .A(n2309), .B(n2310), .Z(n2308) );
  NANDN U2021 ( .A(A[447]), .B(B[447]), .Z(n2310) );
  AND U2022 ( .A(n2311), .B(n2312), .Z(n2309) );
  NANDN U2023 ( .A(A[446]), .B(B[446]), .Z(n2312) );
  NAND U2024 ( .A(n2313), .B(n2314), .Z(n2311) );
  NANDN U2025 ( .A(B[446]), .B(A[446]), .Z(n2314) );
  AND U2026 ( .A(n2315), .B(n2316), .Z(n2313) );
  NAND U2027 ( .A(n2317), .B(n2318), .Z(n2316) );
  NANDN U2028 ( .A(A[445]), .B(B[445]), .Z(n2318) );
  AND U2029 ( .A(n2319), .B(n2320), .Z(n2317) );
  NANDN U2030 ( .A(A[444]), .B(B[444]), .Z(n2320) );
  NAND U2031 ( .A(n2321), .B(n2322), .Z(n2319) );
  NANDN U2032 ( .A(B[444]), .B(A[444]), .Z(n2322) );
  AND U2033 ( .A(n2323), .B(n2324), .Z(n2321) );
  NAND U2034 ( .A(n2325), .B(n2326), .Z(n2324) );
  NANDN U2035 ( .A(A[443]), .B(B[443]), .Z(n2326) );
  AND U2036 ( .A(n2327), .B(n2328), .Z(n2325) );
  NANDN U2037 ( .A(A[442]), .B(B[442]), .Z(n2328) );
  NAND U2038 ( .A(n2329), .B(n2330), .Z(n2327) );
  NANDN U2039 ( .A(B[442]), .B(A[442]), .Z(n2330) );
  AND U2040 ( .A(n2331), .B(n2332), .Z(n2329) );
  NAND U2041 ( .A(n2333), .B(n2334), .Z(n2332) );
  NANDN U2042 ( .A(A[441]), .B(B[441]), .Z(n2334) );
  AND U2043 ( .A(n2335), .B(n2336), .Z(n2333) );
  NANDN U2044 ( .A(A[440]), .B(B[440]), .Z(n2336) );
  NAND U2045 ( .A(n2337), .B(n2338), .Z(n2335) );
  NANDN U2046 ( .A(B[440]), .B(A[440]), .Z(n2338) );
  AND U2047 ( .A(n2339), .B(n2340), .Z(n2337) );
  NAND U2048 ( .A(n2341), .B(n2342), .Z(n2340) );
  NANDN U2049 ( .A(A[439]), .B(B[439]), .Z(n2342) );
  AND U2050 ( .A(n2343), .B(n2344), .Z(n2341) );
  NANDN U2051 ( .A(A[438]), .B(B[438]), .Z(n2344) );
  NAND U2052 ( .A(n2345), .B(n2346), .Z(n2343) );
  NANDN U2053 ( .A(B[438]), .B(A[438]), .Z(n2346) );
  AND U2054 ( .A(n2347), .B(n2348), .Z(n2345) );
  NAND U2055 ( .A(n2349), .B(n2350), .Z(n2348) );
  NANDN U2056 ( .A(A[437]), .B(B[437]), .Z(n2350) );
  AND U2057 ( .A(n2351), .B(n2352), .Z(n2349) );
  NANDN U2058 ( .A(A[436]), .B(B[436]), .Z(n2352) );
  NAND U2059 ( .A(n2353), .B(n2354), .Z(n2351) );
  NANDN U2060 ( .A(B[436]), .B(A[436]), .Z(n2354) );
  AND U2061 ( .A(n2355), .B(n2356), .Z(n2353) );
  NAND U2062 ( .A(n2357), .B(n2358), .Z(n2356) );
  NANDN U2063 ( .A(A[435]), .B(B[435]), .Z(n2358) );
  AND U2064 ( .A(n2359), .B(n2360), .Z(n2357) );
  NANDN U2065 ( .A(A[434]), .B(B[434]), .Z(n2360) );
  NAND U2066 ( .A(n2361), .B(n2362), .Z(n2359) );
  NANDN U2067 ( .A(B[434]), .B(A[434]), .Z(n2362) );
  AND U2068 ( .A(n2363), .B(n2364), .Z(n2361) );
  NAND U2069 ( .A(n2365), .B(n2366), .Z(n2364) );
  NANDN U2070 ( .A(A[433]), .B(B[433]), .Z(n2366) );
  AND U2071 ( .A(n2367), .B(n2368), .Z(n2365) );
  NANDN U2072 ( .A(A[432]), .B(B[432]), .Z(n2368) );
  NAND U2073 ( .A(n2369), .B(n2370), .Z(n2367) );
  NANDN U2074 ( .A(B[432]), .B(A[432]), .Z(n2370) );
  AND U2075 ( .A(n2371), .B(n2372), .Z(n2369) );
  NAND U2076 ( .A(n2373), .B(n2374), .Z(n2372) );
  NANDN U2077 ( .A(A[431]), .B(B[431]), .Z(n2374) );
  AND U2078 ( .A(n2375), .B(n2376), .Z(n2373) );
  NANDN U2079 ( .A(A[430]), .B(B[430]), .Z(n2376) );
  NAND U2080 ( .A(n2377), .B(n2378), .Z(n2375) );
  NANDN U2081 ( .A(B[430]), .B(A[430]), .Z(n2378) );
  AND U2082 ( .A(n2379), .B(n2380), .Z(n2377) );
  NAND U2083 ( .A(n2381), .B(n2382), .Z(n2380) );
  NANDN U2084 ( .A(A[429]), .B(B[429]), .Z(n2382) );
  AND U2085 ( .A(n2383), .B(n2384), .Z(n2381) );
  NANDN U2086 ( .A(A[428]), .B(B[428]), .Z(n2384) );
  NAND U2087 ( .A(n2385), .B(n2386), .Z(n2383) );
  NANDN U2088 ( .A(B[428]), .B(A[428]), .Z(n2386) );
  AND U2089 ( .A(n2387), .B(n2388), .Z(n2385) );
  NAND U2090 ( .A(n2389), .B(n2390), .Z(n2388) );
  NANDN U2091 ( .A(A[427]), .B(B[427]), .Z(n2390) );
  AND U2092 ( .A(n2391), .B(n2392), .Z(n2389) );
  NANDN U2093 ( .A(A[426]), .B(B[426]), .Z(n2392) );
  NAND U2094 ( .A(n2393), .B(n2394), .Z(n2391) );
  NANDN U2095 ( .A(B[426]), .B(A[426]), .Z(n2394) );
  AND U2096 ( .A(n2395), .B(n2396), .Z(n2393) );
  NAND U2097 ( .A(n2397), .B(n2398), .Z(n2396) );
  NANDN U2098 ( .A(A[425]), .B(B[425]), .Z(n2398) );
  AND U2099 ( .A(n2399), .B(n2400), .Z(n2397) );
  NANDN U2100 ( .A(A[424]), .B(B[424]), .Z(n2400) );
  NAND U2101 ( .A(n2401), .B(n2402), .Z(n2399) );
  NANDN U2102 ( .A(B[424]), .B(A[424]), .Z(n2402) );
  AND U2103 ( .A(n2403), .B(n2404), .Z(n2401) );
  NAND U2104 ( .A(n2405), .B(n2406), .Z(n2404) );
  NANDN U2105 ( .A(A[423]), .B(B[423]), .Z(n2406) );
  AND U2106 ( .A(n2407), .B(n2408), .Z(n2405) );
  NANDN U2107 ( .A(A[422]), .B(B[422]), .Z(n2408) );
  NAND U2108 ( .A(n2409), .B(n2410), .Z(n2407) );
  NANDN U2109 ( .A(B[422]), .B(A[422]), .Z(n2410) );
  AND U2110 ( .A(n2411), .B(n2412), .Z(n2409) );
  NAND U2111 ( .A(n2413), .B(n2414), .Z(n2412) );
  NANDN U2112 ( .A(A[421]), .B(B[421]), .Z(n2414) );
  AND U2113 ( .A(n2415), .B(n2416), .Z(n2413) );
  NANDN U2114 ( .A(A[420]), .B(B[420]), .Z(n2416) );
  NAND U2115 ( .A(n2417), .B(n2418), .Z(n2415) );
  NANDN U2116 ( .A(B[420]), .B(A[420]), .Z(n2418) );
  AND U2117 ( .A(n2419), .B(n2420), .Z(n2417) );
  NAND U2118 ( .A(n2421), .B(n2422), .Z(n2420) );
  NANDN U2119 ( .A(A[419]), .B(B[419]), .Z(n2422) );
  AND U2120 ( .A(n2423), .B(n2424), .Z(n2421) );
  NANDN U2121 ( .A(A[418]), .B(B[418]), .Z(n2424) );
  NAND U2122 ( .A(n2425), .B(n2426), .Z(n2423) );
  NANDN U2123 ( .A(B[418]), .B(A[418]), .Z(n2426) );
  AND U2124 ( .A(n2427), .B(n2428), .Z(n2425) );
  NAND U2125 ( .A(n2429), .B(n2430), .Z(n2428) );
  NANDN U2126 ( .A(A[417]), .B(B[417]), .Z(n2430) );
  AND U2127 ( .A(n2431), .B(n2432), .Z(n2429) );
  NANDN U2128 ( .A(A[416]), .B(B[416]), .Z(n2432) );
  NAND U2129 ( .A(n2433), .B(n2434), .Z(n2431) );
  NANDN U2130 ( .A(B[416]), .B(A[416]), .Z(n2434) );
  AND U2131 ( .A(n2435), .B(n2436), .Z(n2433) );
  NAND U2132 ( .A(n2437), .B(n2438), .Z(n2436) );
  NANDN U2133 ( .A(A[415]), .B(B[415]), .Z(n2438) );
  AND U2134 ( .A(n2439), .B(n2440), .Z(n2437) );
  NANDN U2135 ( .A(A[414]), .B(B[414]), .Z(n2440) );
  NAND U2136 ( .A(n2441), .B(n2442), .Z(n2439) );
  NANDN U2137 ( .A(B[414]), .B(A[414]), .Z(n2442) );
  AND U2138 ( .A(n2443), .B(n2444), .Z(n2441) );
  NAND U2139 ( .A(n2445), .B(n2446), .Z(n2444) );
  NANDN U2140 ( .A(A[413]), .B(B[413]), .Z(n2446) );
  AND U2141 ( .A(n2447), .B(n2448), .Z(n2445) );
  NANDN U2142 ( .A(A[412]), .B(B[412]), .Z(n2448) );
  NAND U2143 ( .A(n2449), .B(n2450), .Z(n2447) );
  NANDN U2144 ( .A(B[412]), .B(A[412]), .Z(n2450) );
  AND U2145 ( .A(n2451), .B(n2452), .Z(n2449) );
  NAND U2146 ( .A(n2453), .B(n2454), .Z(n2452) );
  NANDN U2147 ( .A(A[411]), .B(B[411]), .Z(n2454) );
  AND U2148 ( .A(n2455), .B(n2456), .Z(n2453) );
  NANDN U2149 ( .A(A[410]), .B(B[410]), .Z(n2456) );
  NAND U2150 ( .A(n2457), .B(n2458), .Z(n2455) );
  NANDN U2151 ( .A(B[410]), .B(A[410]), .Z(n2458) );
  AND U2152 ( .A(n2459), .B(n2460), .Z(n2457) );
  NAND U2153 ( .A(n2461), .B(n2462), .Z(n2460) );
  NANDN U2154 ( .A(A[409]), .B(B[409]), .Z(n2462) );
  AND U2155 ( .A(n2463), .B(n2464), .Z(n2461) );
  NANDN U2156 ( .A(A[408]), .B(B[408]), .Z(n2464) );
  NAND U2157 ( .A(n2465), .B(n2466), .Z(n2463) );
  NANDN U2158 ( .A(B[408]), .B(A[408]), .Z(n2466) );
  AND U2159 ( .A(n2467), .B(n2468), .Z(n2465) );
  NAND U2160 ( .A(n2469), .B(n2470), .Z(n2468) );
  NANDN U2161 ( .A(A[407]), .B(B[407]), .Z(n2470) );
  AND U2162 ( .A(n2471), .B(n2472), .Z(n2469) );
  NANDN U2163 ( .A(A[406]), .B(B[406]), .Z(n2472) );
  NAND U2164 ( .A(n2473), .B(n2474), .Z(n2471) );
  NANDN U2165 ( .A(B[406]), .B(A[406]), .Z(n2474) );
  AND U2166 ( .A(n2475), .B(n2476), .Z(n2473) );
  NAND U2167 ( .A(n2477), .B(n2478), .Z(n2476) );
  NANDN U2168 ( .A(A[405]), .B(B[405]), .Z(n2478) );
  AND U2169 ( .A(n2479), .B(n2480), .Z(n2477) );
  NANDN U2170 ( .A(A[404]), .B(B[404]), .Z(n2480) );
  NAND U2171 ( .A(n2481), .B(n2482), .Z(n2479) );
  NANDN U2172 ( .A(B[404]), .B(A[404]), .Z(n2482) );
  AND U2173 ( .A(n2483), .B(n2484), .Z(n2481) );
  NAND U2174 ( .A(n2485), .B(n2486), .Z(n2484) );
  NANDN U2175 ( .A(A[403]), .B(B[403]), .Z(n2486) );
  AND U2176 ( .A(n2487), .B(n2488), .Z(n2485) );
  NANDN U2177 ( .A(A[402]), .B(B[402]), .Z(n2488) );
  NAND U2178 ( .A(n2489), .B(n2490), .Z(n2487) );
  NANDN U2179 ( .A(B[402]), .B(A[402]), .Z(n2490) );
  AND U2180 ( .A(n2491), .B(n2492), .Z(n2489) );
  NAND U2181 ( .A(n2493), .B(n2494), .Z(n2492) );
  NANDN U2182 ( .A(A[401]), .B(B[401]), .Z(n2494) );
  AND U2183 ( .A(n2495), .B(n2496), .Z(n2493) );
  NANDN U2184 ( .A(A[400]), .B(B[400]), .Z(n2496) );
  NAND U2185 ( .A(n2497), .B(n2498), .Z(n2495) );
  NANDN U2186 ( .A(B[400]), .B(A[400]), .Z(n2498) );
  AND U2187 ( .A(n2499), .B(n2500), .Z(n2497) );
  NAND U2188 ( .A(n2501), .B(n2502), .Z(n2500) );
  NANDN U2189 ( .A(A[399]), .B(B[399]), .Z(n2502) );
  AND U2190 ( .A(n2503), .B(n2504), .Z(n2501) );
  NANDN U2191 ( .A(A[398]), .B(B[398]), .Z(n2504) );
  NAND U2192 ( .A(n2505), .B(n2506), .Z(n2503) );
  NANDN U2193 ( .A(B[398]), .B(A[398]), .Z(n2506) );
  AND U2194 ( .A(n2507), .B(n2508), .Z(n2505) );
  NAND U2195 ( .A(n2509), .B(n2510), .Z(n2508) );
  NANDN U2196 ( .A(A[397]), .B(B[397]), .Z(n2510) );
  AND U2197 ( .A(n2511), .B(n2512), .Z(n2509) );
  NANDN U2198 ( .A(A[396]), .B(B[396]), .Z(n2512) );
  NAND U2199 ( .A(n2513), .B(n2514), .Z(n2511) );
  NANDN U2200 ( .A(B[396]), .B(A[396]), .Z(n2514) );
  AND U2201 ( .A(n2515), .B(n2516), .Z(n2513) );
  NAND U2202 ( .A(n2517), .B(n2518), .Z(n2516) );
  NANDN U2203 ( .A(A[395]), .B(B[395]), .Z(n2518) );
  AND U2204 ( .A(n2519), .B(n2520), .Z(n2517) );
  NANDN U2205 ( .A(A[394]), .B(B[394]), .Z(n2520) );
  NAND U2206 ( .A(n2521), .B(n2522), .Z(n2519) );
  NANDN U2207 ( .A(B[394]), .B(A[394]), .Z(n2522) );
  AND U2208 ( .A(n2523), .B(n2524), .Z(n2521) );
  NAND U2209 ( .A(n2525), .B(n2526), .Z(n2524) );
  NANDN U2210 ( .A(A[393]), .B(B[393]), .Z(n2526) );
  AND U2211 ( .A(n2527), .B(n2528), .Z(n2525) );
  NANDN U2212 ( .A(A[392]), .B(B[392]), .Z(n2528) );
  NAND U2213 ( .A(n2529), .B(n2530), .Z(n2527) );
  NANDN U2214 ( .A(B[392]), .B(A[392]), .Z(n2530) );
  AND U2215 ( .A(n2531), .B(n2532), .Z(n2529) );
  NAND U2216 ( .A(n2533), .B(n2534), .Z(n2532) );
  NANDN U2217 ( .A(A[391]), .B(B[391]), .Z(n2534) );
  AND U2218 ( .A(n2535), .B(n2536), .Z(n2533) );
  NANDN U2219 ( .A(A[390]), .B(B[390]), .Z(n2536) );
  NAND U2220 ( .A(n2537), .B(n2538), .Z(n2535) );
  NANDN U2221 ( .A(B[390]), .B(A[390]), .Z(n2538) );
  AND U2222 ( .A(n2539), .B(n2540), .Z(n2537) );
  NAND U2223 ( .A(n2541), .B(n2542), .Z(n2540) );
  NANDN U2224 ( .A(A[389]), .B(B[389]), .Z(n2542) );
  AND U2225 ( .A(n2543), .B(n2544), .Z(n2541) );
  NANDN U2226 ( .A(A[388]), .B(B[388]), .Z(n2544) );
  NAND U2227 ( .A(n2545), .B(n2546), .Z(n2543) );
  NANDN U2228 ( .A(B[388]), .B(A[388]), .Z(n2546) );
  AND U2229 ( .A(n2547), .B(n2548), .Z(n2545) );
  NAND U2230 ( .A(n2549), .B(n2550), .Z(n2548) );
  NANDN U2231 ( .A(A[387]), .B(B[387]), .Z(n2550) );
  AND U2232 ( .A(n2551), .B(n2552), .Z(n2549) );
  NANDN U2233 ( .A(A[386]), .B(B[386]), .Z(n2552) );
  NAND U2234 ( .A(n2553), .B(n2554), .Z(n2551) );
  NANDN U2235 ( .A(B[386]), .B(A[386]), .Z(n2554) );
  AND U2236 ( .A(n2555), .B(n2556), .Z(n2553) );
  NAND U2237 ( .A(n2557), .B(n2558), .Z(n2556) );
  NANDN U2238 ( .A(A[385]), .B(B[385]), .Z(n2558) );
  AND U2239 ( .A(n2559), .B(n2560), .Z(n2557) );
  NANDN U2240 ( .A(A[384]), .B(B[384]), .Z(n2560) );
  NAND U2241 ( .A(n2561), .B(n2562), .Z(n2559) );
  NANDN U2242 ( .A(B[384]), .B(A[384]), .Z(n2562) );
  AND U2243 ( .A(n2563), .B(n2564), .Z(n2561) );
  NAND U2244 ( .A(n2565), .B(n2566), .Z(n2564) );
  NANDN U2245 ( .A(A[383]), .B(B[383]), .Z(n2566) );
  AND U2246 ( .A(n2567), .B(n2568), .Z(n2565) );
  NANDN U2247 ( .A(A[382]), .B(B[382]), .Z(n2568) );
  NAND U2248 ( .A(n2569), .B(n2570), .Z(n2567) );
  NANDN U2249 ( .A(B[382]), .B(A[382]), .Z(n2570) );
  AND U2250 ( .A(n2571), .B(n2572), .Z(n2569) );
  NAND U2251 ( .A(n2573), .B(n2574), .Z(n2572) );
  NANDN U2252 ( .A(A[381]), .B(B[381]), .Z(n2574) );
  AND U2253 ( .A(n2575), .B(n2576), .Z(n2573) );
  NANDN U2254 ( .A(A[380]), .B(B[380]), .Z(n2576) );
  NAND U2255 ( .A(n2577), .B(n2578), .Z(n2575) );
  NANDN U2256 ( .A(B[380]), .B(A[380]), .Z(n2578) );
  AND U2257 ( .A(n2579), .B(n2580), .Z(n2577) );
  NAND U2258 ( .A(n2581), .B(n2582), .Z(n2580) );
  NANDN U2259 ( .A(A[379]), .B(B[379]), .Z(n2582) );
  AND U2260 ( .A(n2583), .B(n2584), .Z(n2581) );
  NANDN U2261 ( .A(A[378]), .B(B[378]), .Z(n2584) );
  NAND U2262 ( .A(n2585), .B(n2586), .Z(n2583) );
  NANDN U2263 ( .A(B[378]), .B(A[378]), .Z(n2586) );
  AND U2264 ( .A(n2587), .B(n2588), .Z(n2585) );
  NAND U2265 ( .A(n2589), .B(n2590), .Z(n2588) );
  NANDN U2266 ( .A(A[377]), .B(B[377]), .Z(n2590) );
  AND U2267 ( .A(n2591), .B(n2592), .Z(n2589) );
  NANDN U2268 ( .A(A[376]), .B(B[376]), .Z(n2592) );
  NAND U2269 ( .A(n2593), .B(n2594), .Z(n2591) );
  NANDN U2270 ( .A(B[376]), .B(A[376]), .Z(n2594) );
  AND U2271 ( .A(n2595), .B(n2596), .Z(n2593) );
  NAND U2272 ( .A(n2597), .B(n2598), .Z(n2596) );
  NANDN U2273 ( .A(A[375]), .B(B[375]), .Z(n2598) );
  AND U2274 ( .A(n2599), .B(n2600), .Z(n2597) );
  NANDN U2275 ( .A(A[374]), .B(B[374]), .Z(n2600) );
  NAND U2276 ( .A(n2601), .B(n2602), .Z(n2599) );
  NANDN U2277 ( .A(B[374]), .B(A[374]), .Z(n2602) );
  AND U2278 ( .A(n2603), .B(n2604), .Z(n2601) );
  NAND U2279 ( .A(n2605), .B(n2606), .Z(n2604) );
  NANDN U2280 ( .A(A[373]), .B(B[373]), .Z(n2606) );
  AND U2281 ( .A(n2607), .B(n2608), .Z(n2605) );
  NANDN U2282 ( .A(A[372]), .B(B[372]), .Z(n2608) );
  NAND U2283 ( .A(n2609), .B(n2610), .Z(n2607) );
  NANDN U2284 ( .A(B[372]), .B(A[372]), .Z(n2610) );
  AND U2285 ( .A(n2611), .B(n2612), .Z(n2609) );
  NAND U2286 ( .A(n2613), .B(n2614), .Z(n2612) );
  NANDN U2287 ( .A(A[371]), .B(B[371]), .Z(n2614) );
  AND U2288 ( .A(n2615), .B(n2616), .Z(n2613) );
  NANDN U2289 ( .A(A[370]), .B(B[370]), .Z(n2616) );
  NAND U2290 ( .A(n2617), .B(n2618), .Z(n2615) );
  NANDN U2291 ( .A(B[370]), .B(A[370]), .Z(n2618) );
  AND U2292 ( .A(n2619), .B(n2620), .Z(n2617) );
  NAND U2293 ( .A(n2621), .B(n2622), .Z(n2620) );
  NANDN U2294 ( .A(A[369]), .B(B[369]), .Z(n2622) );
  AND U2295 ( .A(n2623), .B(n2624), .Z(n2621) );
  NANDN U2296 ( .A(A[368]), .B(B[368]), .Z(n2624) );
  NAND U2297 ( .A(n2625), .B(n2626), .Z(n2623) );
  NANDN U2298 ( .A(B[368]), .B(A[368]), .Z(n2626) );
  AND U2299 ( .A(n2627), .B(n2628), .Z(n2625) );
  NAND U2300 ( .A(n2629), .B(n2630), .Z(n2628) );
  NANDN U2301 ( .A(A[367]), .B(B[367]), .Z(n2630) );
  AND U2302 ( .A(n2631), .B(n2632), .Z(n2629) );
  NANDN U2303 ( .A(A[366]), .B(B[366]), .Z(n2632) );
  NAND U2304 ( .A(n2633), .B(n2634), .Z(n2631) );
  NANDN U2305 ( .A(B[366]), .B(A[366]), .Z(n2634) );
  AND U2306 ( .A(n2635), .B(n2636), .Z(n2633) );
  NAND U2307 ( .A(n2637), .B(n2638), .Z(n2636) );
  NANDN U2308 ( .A(A[365]), .B(B[365]), .Z(n2638) );
  AND U2309 ( .A(n2639), .B(n2640), .Z(n2637) );
  NANDN U2310 ( .A(A[364]), .B(B[364]), .Z(n2640) );
  NAND U2311 ( .A(n2641), .B(n2642), .Z(n2639) );
  NANDN U2312 ( .A(B[364]), .B(A[364]), .Z(n2642) );
  AND U2313 ( .A(n2643), .B(n2644), .Z(n2641) );
  NAND U2314 ( .A(n2645), .B(n2646), .Z(n2644) );
  NANDN U2315 ( .A(A[363]), .B(B[363]), .Z(n2646) );
  AND U2316 ( .A(n2647), .B(n2648), .Z(n2645) );
  NANDN U2317 ( .A(A[362]), .B(B[362]), .Z(n2648) );
  NAND U2318 ( .A(n2649), .B(n2650), .Z(n2647) );
  NANDN U2319 ( .A(B[362]), .B(A[362]), .Z(n2650) );
  AND U2320 ( .A(n2651), .B(n2652), .Z(n2649) );
  NAND U2321 ( .A(n2653), .B(n2654), .Z(n2652) );
  NANDN U2322 ( .A(A[361]), .B(B[361]), .Z(n2654) );
  AND U2323 ( .A(n2655), .B(n2656), .Z(n2653) );
  NANDN U2324 ( .A(A[360]), .B(B[360]), .Z(n2656) );
  NAND U2325 ( .A(n2657), .B(n2658), .Z(n2655) );
  NANDN U2326 ( .A(B[360]), .B(A[360]), .Z(n2658) );
  AND U2327 ( .A(n2659), .B(n2660), .Z(n2657) );
  NAND U2328 ( .A(n2661), .B(n2662), .Z(n2660) );
  NANDN U2329 ( .A(A[359]), .B(B[359]), .Z(n2662) );
  AND U2330 ( .A(n2663), .B(n2664), .Z(n2661) );
  NANDN U2331 ( .A(A[358]), .B(B[358]), .Z(n2664) );
  NAND U2332 ( .A(n2665), .B(n2666), .Z(n2663) );
  NANDN U2333 ( .A(B[358]), .B(A[358]), .Z(n2666) );
  AND U2334 ( .A(n2667), .B(n2668), .Z(n2665) );
  NAND U2335 ( .A(n2669), .B(n2670), .Z(n2668) );
  NANDN U2336 ( .A(A[357]), .B(B[357]), .Z(n2670) );
  AND U2337 ( .A(n2671), .B(n2672), .Z(n2669) );
  NANDN U2338 ( .A(A[356]), .B(B[356]), .Z(n2672) );
  NAND U2339 ( .A(n2673), .B(n2674), .Z(n2671) );
  NANDN U2340 ( .A(B[356]), .B(A[356]), .Z(n2674) );
  AND U2341 ( .A(n2675), .B(n2676), .Z(n2673) );
  NAND U2342 ( .A(n2677), .B(n2678), .Z(n2676) );
  NANDN U2343 ( .A(A[355]), .B(B[355]), .Z(n2678) );
  AND U2344 ( .A(n2679), .B(n2680), .Z(n2677) );
  NANDN U2345 ( .A(A[354]), .B(B[354]), .Z(n2680) );
  NAND U2346 ( .A(n2681), .B(n2682), .Z(n2679) );
  NANDN U2347 ( .A(B[354]), .B(A[354]), .Z(n2682) );
  AND U2348 ( .A(n2683), .B(n2684), .Z(n2681) );
  NAND U2349 ( .A(n2685), .B(n2686), .Z(n2684) );
  NANDN U2350 ( .A(A[353]), .B(B[353]), .Z(n2686) );
  AND U2351 ( .A(n2687), .B(n2688), .Z(n2685) );
  NANDN U2352 ( .A(A[352]), .B(B[352]), .Z(n2688) );
  NAND U2353 ( .A(n2689), .B(n2690), .Z(n2687) );
  NANDN U2354 ( .A(B[352]), .B(A[352]), .Z(n2690) );
  AND U2355 ( .A(n2691), .B(n2692), .Z(n2689) );
  NAND U2356 ( .A(n2693), .B(n2694), .Z(n2692) );
  NANDN U2357 ( .A(A[351]), .B(B[351]), .Z(n2694) );
  AND U2358 ( .A(n2695), .B(n2696), .Z(n2693) );
  NANDN U2359 ( .A(A[350]), .B(B[350]), .Z(n2696) );
  NAND U2360 ( .A(n2697), .B(n2698), .Z(n2695) );
  NANDN U2361 ( .A(B[350]), .B(A[350]), .Z(n2698) );
  AND U2362 ( .A(n2699), .B(n2700), .Z(n2697) );
  NAND U2363 ( .A(n2701), .B(n2702), .Z(n2700) );
  NANDN U2364 ( .A(A[349]), .B(B[349]), .Z(n2702) );
  AND U2365 ( .A(n2703), .B(n2704), .Z(n2701) );
  NANDN U2366 ( .A(A[348]), .B(B[348]), .Z(n2704) );
  NAND U2367 ( .A(n2705), .B(n2706), .Z(n2703) );
  NANDN U2368 ( .A(B[348]), .B(A[348]), .Z(n2706) );
  AND U2369 ( .A(n2707), .B(n2708), .Z(n2705) );
  NAND U2370 ( .A(n2709), .B(n2710), .Z(n2708) );
  NANDN U2371 ( .A(A[347]), .B(B[347]), .Z(n2710) );
  AND U2372 ( .A(n2711), .B(n2712), .Z(n2709) );
  NANDN U2373 ( .A(A[346]), .B(B[346]), .Z(n2712) );
  NAND U2374 ( .A(n2713), .B(n2714), .Z(n2711) );
  NANDN U2375 ( .A(B[346]), .B(A[346]), .Z(n2714) );
  AND U2376 ( .A(n2715), .B(n2716), .Z(n2713) );
  NAND U2377 ( .A(n2717), .B(n2718), .Z(n2716) );
  NANDN U2378 ( .A(A[345]), .B(B[345]), .Z(n2718) );
  AND U2379 ( .A(n2719), .B(n2720), .Z(n2717) );
  NANDN U2380 ( .A(A[344]), .B(B[344]), .Z(n2720) );
  NAND U2381 ( .A(n2721), .B(n2722), .Z(n2719) );
  NANDN U2382 ( .A(B[344]), .B(A[344]), .Z(n2722) );
  AND U2383 ( .A(n2723), .B(n2724), .Z(n2721) );
  NAND U2384 ( .A(n2725), .B(n2726), .Z(n2724) );
  NANDN U2385 ( .A(A[343]), .B(B[343]), .Z(n2726) );
  AND U2386 ( .A(n2727), .B(n2728), .Z(n2725) );
  NANDN U2387 ( .A(A[342]), .B(B[342]), .Z(n2728) );
  NAND U2388 ( .A(n2729), .B(n2730), .Z(n2727) );
  NANDN U2389 ( .A(B[342]), .B(A[342]), .Z(n2730) );
  AND U2390 ( .A(n2731), .B(n2732), .Z(n2729) );
  NAND U2391 ( .A(n2733), .B(n2734), .Z(n2732) );
  NANDN U2392 ( .A(A[341]), .B(B[341]), .Z(n2734) );
  AND U2393 ( .A(n2735), .B(n2736), .Z(n2733) );
  NANDN U2394 ( .A(A[340]), .B(B[340]), .Z(n2736) );
  NAND U2395 ( .A(n2737), .B(n2738), .Z(n2735) );
  NANDN U2396 ( .A(B[340]), .B(A[340]), .Z(n2738) );
  AND U2397 ( .A(n2739), .B(n2740), .Z(n2737) );
  NAND U2398 ( .A(n2741), .B(n2742), .Z(n2740) );
  NANDN U2399 ( .A(A[339]), .B(B[339]), .Z(n2742) );
  AND U2400 ( .A(n2743), .B(n2744), .Z(n2741) );
  NANDN U2401 ( .A(A[338]), .B(B[338]), .Z(n2744) );
  NAND U2402 ( .A(n2745), .B(n2746), .Z(n2743) );
  NANDN U2403 ( .A(B[338]), .B(A[338]), .Z(n2746) );
  AND U2404 ( .A(n2747), .B(n2748), .Z(n2745) );
  NAND U2405 ( .A(n2749), .B(n2750), .Z(n2748) );
  NANDN U2406 ( .A(A[337]), .B(B[337]), .Z(n2750) );
  AND U2407 ( .A(n2751), .B(n2752), .Z(n2749) );
  NANDN U2408 ( .A(A[336]), .B(B[336]), .Z(n2752) );
  NAND U2409 ( .A(n2753), .B(n2754), .Z(n2751) );
  NANDN U2410 ( .A(B[336]), .B(A[336]), .Z(n2754) );
  AND U2411 ( .A(n2755), .B(n2756), .Z(n2753) );
  NAND U2412 ( .A(n2757), .B(n2758), .Z(n2756) );
  NANDN U2413 ( .A(A[335]), .B(B[335]), .Z(n2758) );
  AND U2414 ( .A(n2759), .B(n2760), .Z(n2757) );
  NANDN U2415 ( .A(A[334]), .B(B[334]), .Z(n2760) );
  NAND U2416 ( .A(n2761), .B(n2762), .Z(n2759) );
  NANDN U2417 ( .A(B[334]), .B(A[334]), .Z(n2762) );
  AND U2418 ( .A(n2763), .B(n2764), .Z(n2761) );
  NAND U2419 ( .A(n2765), .B(n2766), .Z(n2764) );
  NANDN U2420 ( .A(A[333]), .B(B[333]), .Z(n2766) );
  AND U2421 ( .A(n2767), .B(n2768), .Z(n2765) );
  NANDN U2422 ( .A(A[332]), .B(B[332]), .Z(n2768) );
  NAND U2423 ( .A(n2769), .B(n2770), .Z(n2767) );
  NANDN U2424 ( .A(B[332]), .B(A[332]), .Z(n2770) );
  AND U2425 ( .A(n2771), .B(n2772), .Z(n2769) );
  NAND U2426 ( .A(n2773), .B(n2774), .Z(n2772) );
  NANDN U2427 ( .A(A[331]), .B(B[331]), .Z(n2774) );
  AND U2428 ( .A(n2775), .B(n2776), .Z(n2773) );
  NANDN U2429 ( .A(A[330]), .B(B[330]), .Z(n2776) );
  NAND U2430 ( .A(n2777), .B(n2778), .Z(n2775) );
  NANDN U2431 ( .A(B[330]), .B(A[330]), .Z(n2778) );
  AND U2432 ( .A(n2779), .B(n2780), .Z(n2777) );
  NAND U2433 ( .A(n2781), .B(n2782), .Z(n2780) );
  NANDN U2434 ( .A(A[329]), .B(B[329]), .Z(n2782) );
  AND U2435 ( .A(n2783), .B(n2784), .Z(n2781) );
  NANDN U2436 ( .A(A[328]), .B(B[328]), .Z(n2784) );
  NAND U2437 ( .A(n2785), .B(n2786), .Z(n2783) );
  NANDN U2438 ( .A(B[328]), .B(A[328]), .Z(n2786) );
  AND U2439 ( .A(n2787), .B(n2788), .Z(n2785) );
  NAND U2440 ( .A(n2789), .B(n2790), .Z(n2788) );
  NANDN U2441 ( .A(A[327]), .B(B[327]), .Z(n2790) );
  AND U2442 ( .A(n2791), .B(n2792), .Z(n2789) );
  NANDN U2443 ( .A(A[326]), .B(B[326]), .Z(n2792) );
  NAND U2444 ( .A(n2793), .B(n2794), .Z(n2791) );
  NANDN U2445 ( .A(B[326]), .B(A[326]), .Z(n2794) );
  AND U2446 ( .A(n2795), .B(n2796), .Z(n2793) );
  NAND U2447 ( .A(n2797), .B(n2798), .Z(n2796) );
  NANDN U2448 ( .A(A[325]), .B(B[325]), .Z(n2798) );
  AND U2449 ( .A(n2799), .B(n2800), .Z(n2797) );
  NANDN U2450 ( .A(A[324]), .B(B[324]), .Z(n2800) );
  NAND U2451 ( .A(n2801), .B(n2802), .Z(n2799) );
  NANDN U2452 ( .A(B[324]), .B(A[324]), .Z(n2802) );
  AND U2453 ( .A(n2803), .B(n2804), .Z(n2801) );
  NAND U2454 ( .A(n2805), .B(n2806), .Z(n2804) );
  NANDN U2455 ( .A(A[323]), .B(B[323]), .Z(n2806) );
  AND U2456 ( .A(n2807), .B(n2808), .Z(n2805) );
  NANDN U2457 ( .A(A[322]), .B(B[322]), .Z(n2808) );
  NAND U2458 ( .A(n2809), .B(n2810), .Z(n2807) );
  NANDN U2459 ( .A(B[322]), .B(A[322]), .Z(n2810) );
  AND U2460 ( .A(n2811), .B(n2812), .Z(n2809) );
  NAND U2461 ( .A(n2813), .B(n2814), .Z(n2812) );
  NANDN U2462 ( .A(A[321]), .B(B[321]), .Z(n2814) );
  AND U2463 ( .A(n2815), .B(n2816), .Z(n2813) );
  NANDN U2464 ( .A(A[320]), .B(B[320]), .Z(n2816) );
  NAND U2465 ( .A(n2817), .B(n2818), .Z(n2815) );
  NANDN U2466 ( .A(B[320]), .B(A[320]), .Z(n2818) );
  AND U2467 ( .A(n2819), .B(n2820), .Z(n2817) );
  NAND U2468 ( .A(n2821), .B(n2822), .Z(n2820) );
  NANDN U2469 ( .A(A[319]), .B(B[319]), .Z(n2822) );
  AND U2470 ( .A(n2823), .B(n2824), .Z(n2821) );
  NANDN U2471 ( .A(A[318]), .B(B[318]), .Z(n2824) );
  NAND U2472 ( .A(n2825), .B(n2826), .Z(n2823) );
  NANDN U2473 ( .A(B[318]), .B(A[318]), .Z(n2826) );
  AND U2474 ( .A(n2827), .B(n2828), .Z(n2825) );
  NAND U2475 ( .A(n2829), .B(n2830), .Z(n2828) );
  NANDN U2476 ( .A(A[317]), .B(B[317]), .Z(n2830) );
  AND U2477 ( .A(n2831), .B(n2832), .Z(n2829) );
  NANDN U2478 ( .A(A[316]), .B(B[316]), .Z(n2832) );
  NAND U2479 ( .A(n2833), .B(n2834), .Z(n2831) );
  NANDN U2480 ( .A(B[316]), .B(A[316]), .Z(n2834) );
  AND U2481 ( .A(n2835), .B(n2836), .Z(n2833) );
  NAND U2482 ( .A(n2837), .B(n2838), .Z(n2836) );
  NANDN U2483 ( .A(A[315]), .B(B[315]), .Z(n2838) );
  AND U2484 ( .A(n2839), .B(n2840), .Z(n2837) );
  NANDN U2485 ( .A(A[314]), .B(B[314]), .Z(n2840) );
  NAND U2486 ( .A(n2841), .B(n2842), .Z(n2839) );
  NANDN U2487 ( .A(B[314]), .B(A[314]), .Z(n2842) );
  AND U2488 ( .A(n2843), .B(n2844), .Z(n2841) );
  NAND U2489 ( .A(n2845), .B(n2846), .Z(n2844) );
  NANDN U2490 ( .A(A[313]), .B(B[313]), .Z(n2846) );
  AND U2491 ( .A(n2847), .B(n2848), .Z(n2845) );
  NANDN U2492 ( .A(A[312]), .B(B[312]), .Z(n2848) );
  NAND U2493 ( .A(n2849), .B(n2850), .Z(n2847) );
  NANDN U2494 ( .A(B[312]), .B(A[312]), .Z(n2850) );
  AND U2495 ( .A(n2851), .B(n2852), .Z(n2849) );
  NAND U2496 ( .A(n2853), .B(n2854), .Z(n2852) );
  NANDN U2497 ( .A(A[311]), .B(B[311]), .Z(n2854) );
  AND U2498 ( .A(n2855), .B(n2856), .Z(n2853) );
  NANDN U2499 ( .A(A[310]), .B(B[310]), .Z(n2856) );
  NAND U2500 ( .A(n2857), .B(n2858), .Z(n2855) );
  NANDN U2501 ( .A(B[310]), .B(A[310]), .Z(n2858) );
  AND U2502 ( .A(n2859), .B(n2860), .Z(n2857) );
  NAND U2503 ( .A(n2861), .B(n2862), .Z(n2860) );
  NANDN U2504 ( .A(A[309]), .B(B[309]), .Z(n2862) );
  AND U2505 ( .A(n2863), .B(n2864), .Z(n2861) );
  NANDN U2506 ( .A(A[308]), .B(B[308]), .Z(n2864) );
  NAND U2507 ( .A(n2865), .B(n2866), .Z(n2863) );
  NANDN U2508 ( .A(B[308]), .B(A[308]), .Z(n2866) );
  AND U2509 ( .A(n2867), .B(n2868), .Z(n2865) );
  NAND U2510 ( .A(n2869), .B(n2870), .Z(n2868) );
  NANDN U2511 ( .A(A[307]), .B(B[307]), .Z(n2870) );
  AND U2512 ( .A(n2871), .B(n2872), .Z(n2869) );
  NANDN U2513 ( .A(A[306]), .B(B[306]), .Z(n2872) );
  NAND U2514 ( .A(n2873), .B(n2874), .Z(n2871) );
  NANDN U2515 ( .A(B[306]), .B(A[306]), .Z(n2874) );
  AND U2516 ( .A(n2875), .B(n2876), .Z(n2873) );
  NAND U2517 ( .A(n2877), .B(n2878), .Z(n2876) );
  NANDN U2518 ( .A(A[305]), .B(B[305]), .Z(n2878) );
  AND U2519 ( .A(n2879), .B(n2880), .Z(n2877) );
  NANDN U2520 ( .A(A[304]), .B(B[304]), .Z(n2880) );
  NAND U2521 ( .A(n2881), .B(n2882), .Z(n2879) );
  NANDN U2522 ( .A(B[304]), .B(A[304]), .Z(n2882) );
  AND U2523 ( .A(n2883), .B(n2884), .Z(n2881) );
  NAND U2524 ( .A(n2885), .B(n2886), .Z(n2884) );
  NANDN U2525 ( .A(A[303]), .B(B[303]), .Z(n2886) );
  AND U2526 ( .A(n2887), .B(n2888), .Z(n2885) );
  NANDN U2527 ( .A(A[302]), .B(B[302]), .Z(n2888) );
  NAND U2528 ( .A(n2889), .B(n2890), .Z(n2887) );
  NANDN U2529 ( .A(B[302]), .B(A[302]), .Z(n2890) );
  AND U2530 ( .A(n2891), .B(n2892), .Z(n2889) );
  NAND U2531 ( .A(n2893), .B(n2894), .Z(n2892) );
  NANDN U2532 ( .A(A[301]), .B(B[301]), .Z(n2894) );
  AND U2533 ( .A(n2895), .B(n2896), .Z(n2893) );
  NANDN U2534 ( .A(A[300]), .B(B[300]), .Z(n2896) );
  NAND U2535 ( .A(n2897), .B(n2898), .Z(n2895) );
  NANDN U2536 ( .A(B[300]), .B(A[300]), .Z(n2898) );
  AND U2537 ( .A(n2899), .B(n2900), .Z(n2897) );
  NAND U2538 ( .A(n2901), .B(n2902), .Z(n2900) );
  NANDN U2539 ( .A(A[299]), .B(B[299]), .Z(n2902) );
  AND U2540 ( .A(n2903), .B(n2904), .Z(n2901) );
  NANDN U2541 ( .A(A[298]), .B(B[298]), .Z(n2904) );
  NAND U2542 ( .A(n2905), .B(n2906), .Z(n2903) );
  NANDN U2543 ( .A(B[298]), .B(A[298]), .Z(n2906) );
  AND U2544 ( .A(n2907), .B(n2908), .Z(n2905) );
  NAND U2545 ( .A(n2909), .B(n2910), .Z(n2908) );
  NANDN U2546 ( .A(A[297]), .B(B[297]), .Z(n2910) );
  AND U2547 ( .A(n2911), .B(n2912), .Z(n2909) );
  NANDN U2548 ( .A(A[296]), .B(B[296]), .Z(n2912) );
  NAND U2549 ( .A(n2913), .B(n2914), .Z(n2911) );
  NANDN U2550 ( .A(B[296]), .B(A[296]), .Z(n2914) );
  AND U2551 ( .A(n2915), .B(n2916), .Z(n2913) );
  NAND U2552 ( .A(n2917), .B(n2918), .Z(n2916) );
  NANDN U2553 ( .A(A[295]), .B(B[295]), .Z(n2918) );
  AND U2554 ( .A(n2919), .B(n2920), .Z(n2917) );
  NANDN U2555 ( .A(A[294]), .B(B[294]), .Z(n2920) );
  NAND U2556 ( .A(n2921), .B(n2922), .Z(n2919) );
  NANDN U2557 ( .A(B[294]), .B(A[294]), .Z(n2922) );
  AND U2558 ( .A(n2923), .B(n2924), .Z(n2921) );
  NAND U2559 ( .A(n2925), .B(n2926), .Z(n2924) );
  NANDN U2560 ( .A(A[293]), .B(B[293]), .Z(n2926) );
  AND U2561 ( .A(n2927), .B(n2928), .Z(n2925) );
  NANDN U2562 ( .A(A[292]), .B(B[292]), .Z(n2928) );
  NAND U2563 ( .A(n2929), .B(n2930), .Z(n2927) );
  NANDN U2564 ( .A(B[292]), .B(A[292]), .Z(n2930) );
  AND U2565 ( .A(n2931), .B(n2932), .Z(n2929) );
  NAND U2566 ( .A(n2933), .B(n2934), .Z(n2932) );
  NANDN U2567 ( .A(A[291]), .B(B[291]), .Z(n2934) );
  AND U2568 ( .A(n2935), .B(n2936), .Z(n2933) );
  NANDN U2569 ( .A(A[290]), .B(B[290]), .Z(n2936) );
  NAND U2570 ( .A(n2937), .B(n2938), .Z(n2935) );
  NANDN U2571 ( .A(B[290]), .B(A[290]), .Z(n2938) );
  AND U2572 ( .A(n2939), .B(n2940), .Z(n2937) );
  NAND U2573 ( .A(n2941), .B(n2942), .Z(n2940) );
  NANDN U2574 ( .A(A[289]), .B(B[289]), .Z(n2942) );
  AND U2575 ( .A(n2943), .B(n2944), .Z(n2941) );
  NANDN U2576 ( .A(A[288]), .B(B[288]), .Z(n2944) );
  NAND U2577 ( .A(n2945), .B(n2946), .Z(n2943) );
  NANDN U2578 ( .A(B[288]), .B(A[288]), .Z(n2946) );
  AND U2579 ( .A(n2947), .B(n2948), .Z(n2945) );
  NAND U2580 ( .A(n2949), .B(n2950), .Z(n2948) );
  NANDN U2581 ( .A(A[287]), .B(B[287]), .Z(n2950) );
  AND U2582 ( .A(n2951), .B(n2952), .Z(n2949) );
  NANDN U2583 ( .A(A[286]), .B(B[286]), .Z(n2952) );
  NAND U2584 ( .A(n2953), .B(n2954), .Z(n2951) );
  NANDN U2585 ( .A(B[286]), .B(A[286]), .Z(n2954) );
  AND U2586 ( .A(n2955), .B(n2956), .Z(n2953) );
  NAND U2587 ( .A(n2957), .B(n2958), .Z(n2956) );
  NANDN U2588 ( .A(A[285]), .B(B[285]), .Z(n2958) );
  AND U2589 ( .A(n2959), .B(n2960), .Z(n2957) );
  NANDN U2590 ( .A(A[284]), .B(B[284]), .Z(n2960) );
  NAND U2591 ( .A(n2961), .B(n2962), .Z(n2959) );
  NANDN U2592 ( .A(B[284]), .B(A[284]), .Z(n2962) );
  AND U2593 ( .A(n2963), .B(n2964), .Z(n2961) );
  NAND U2594 ( .A(n2965), .B(n2966), .Z(n2964) );
  NANDN U2595 ( .A(A[283]), .B(B[283]), .Z(n2966) );
  AND U2596 ( .A(n2967), .B(n2968), .Z(n2965) );
  NANDN U2597 ( .A(A[282]), .B(B[282]), .Z(n2968) );
  NAND U2598 ( .A(n2969), .B(n2970), .Z(n2967) );
  NANDN U2599 ( .A(B[282]), .B(A[282]), .Z(n2970) );
  AND U2600 ( .A(n2971), .B(n2972), .Z(n2969) );
  NAND U2601 ( .A(n2973), .B(n2974), .Z(n2972) );
  NANDN U2602 ( .A(A[281]), .B(B[281]), .Z(n2974) );
  AND U2603 ( .A(n2975), .B(n2976), .Z(n2973) );
  NANDN U2604 ( .A(A[280]), .B(B[280]), .Z(n2976) );
  NAND U2605 ( .A(n2977), .B(n2978), .Z(n2975) );
  NANDN U2606 ( .A(B[280]), .B(A[280]), .Z(n2978) );
  AND U2607 ( .A(n2979), .B(n2980), .Z(n2977) );
  NAND U2608 ( .A(n2981), .B(n2982), .Z(n2980) );
  NANDN U2609 ( .A(A[279]), .B(B[279]), .Z(n2982) );
  AND U2610 ( .A(n2983), .B(n2984), .Z(n2981) );
  NANDN U2611 ( .A(A[278]), .B(B[278]), .Z(n2984) );
  NAND U2612 ( .A(n2985), .B(n2986), .Z(n2983) );
  NANDN U2613 ( .A(B[278]), .B(A[278]), .Z(n2986) );
  AND U2614 ( .A(n2987), .B(n2988), .Z(n2985) );
  NAND U2615 ( .A(n2989), .B(n2990), .Z(n2988) );
  NANDN U2616 ( .A(A[277]), .B(B[277]), .Z(n2990) );
  AND U2617 ( .A(n2991), .B(n2992), .Z(n2989) );
  NANDN U2618 ( .A(A[276]), .B(B[276]), .Z(n2992) );
  NAND U2619 ( .A(n2993), .B(n2994), .Z(n2991) );
  NANDN U2620 ( .A(B[276]), .B(A[276]), .Z(n2994) );
  AND U2621 ( .A(n2995), .B(n2996), .Z(n2993) );
  NAND U2622 ( .A(n2997), .B(n2998), .Z(n2996) );
  NANDN U2623 ( .A(A[275]), .B(B[275]), .Z(n2998) );
  AND U2624 ( .A(n2999), .B(n3000), .Z(n2997) );
  NANDN U2625 ( .A(A[274]), .B(B[274]), .Z(n3000) );
  NAND U2626 ( .A(n3001), .B(n3002), .Z(n2999) );
  NANDN U2627 ( .A(B[274]), .B(A[274]), .Z(n3002) );
  AND U2628 ( .A(n3003), .B(n3004), .Z(n3001) );
  NAND U2629 ( .A(n3005), .B(n3006), .Z(n3004) );
  NANDN U2630 ( .A(A[273]), .B(B[273]), .Z(n3006) );
  AND U2631 ( .A(n3007), .B(n3008), .Z(n3005) );
  NANDN U2632 ( .A(A[272]), .B(B[272]), .Z(n3008) );
  NAND U2633 ( .A(n3009), .B(n3010), .Z(n3007) );
  NANDN U2634 ( .A(B[272]), .B(A[272]), .Z(n3010) );
  AND U2635 ( .A(n3011), .B(n3012), .Z(n3009) );
  NAND U2636 ( .A(n3013), .B(n3014), .Z(n3012) );
  NANDN U2637 ( .A(A[271]), .B(B[271]), .Z(n3014) );
  AND U2638 ( .A(n3015), .B(n3016), .Z(n3013) );
  NANDN U2639 ( .A(A[270]), .B(B[270]), .Z(n3016) );
  NAND U2640 ( .A(n3017), .B(n3018), .Z(n3015) );
  NANDN U2641 ( .A(B[270]), .B(A[270]), .Z(n3018) );
  AND U2642 ( .A(n3019), .B(n3020), .Z(n3017) );
  NAND U2643 ( .A(n3021), .B(n3022), .Z(n3020) );
  NANDN U2644 ( .A(A[269]), .B(B[269]), .Z(n3022) );
  AND U2645 ( .A(n3023), .B(n3024), .Z(n3021) );
  NANDN U2646 ( .A(A[268]), .B(B[268]), .Z(n3024) );
  NAND U2647 ( .A(n3025), .B(n3026), .Z(n3023) );
  NANDN U2648 ( .A(B[268]), .B(A[268]), .Z(n3026) );
  AND U2649 ( .A(n3027), .B(n3028), .Z(n3025) );
  NAND U2650 ( .A(n3029), .B(n3030), .Z(n3028) );
  NANDN U2651 ( .A(A[267]), .B(B[267]), .Z(n3030) );
  AND U2652 ( .A(n3031), .B(n3032), .Z(n3029) );
  NANDN U2653 ( .A(A[266]), .B(B[266]), .Z(n3032) );
  NAND U2654 ( .A(n3033), .B(n3034), .Z(n3031) );
  NANDN U2655 ( .A(B[266]), .B(A[266]), .Z(n3034) );
  AND U2656 ( .A(n3035), .B(n3036), .Z(n3033) );
  NAND U2657 ( .A(n3037), .B(n3038), .Z(n3036) );
  NANDN U2658 ( .A(A[265]), .B(B[265]), .Z(n3038) );
  AND U2659 ( .A(n3039), .B(n3040), .Z(n3037) );
  NANDN U2660 ( .A(A[264]), .B(B[264]), .Z(n3040) );
  NAND U2661 ( .A(n3041), .B(n3042), .Z(n3039) );
  NANDN U2662 ( .A(B[264]), .B(A[264]), .Z(n3042) );
  AND U2663 ( .A(n3043), .B(n3044), .Z(n3041) );
  NAND U2664 ( .A(n3045), .B(n3046), .Z(n3044) );
  NANDN U2665 ( .A(A[263]), .B(B[263]), .Z(n3046) );
  AND U2666 ( .A(n3047), .B(n3048), .Z(n3045) );
  NANDN U2667 ( .A(A[262]), .B(B[262]), .Z(n3048) );
  NAND U2668 ( .A(n3049), .B(n3050), .Z(n3047) );
  NANDN U2669 ( .A(B[262]), .B(A[262]), .Z(n3050) );
  AND U2670 ( .A(n3051), .B(n3052), .Z(n3049) );
  NAND U2671 ( .A(n3053), .B(n3054), .Z(n3052) );
  NANDN U2672 ( .A(A[261]), .B(B[261]), .Z(n3054) );
  AND U2673 ( .A(n3055), .B(n3056), .Z(n3053) );
  NANDN U2674 ( .A(A[260]), .B(B[260]), .Z(n3056) );
  NAND U2675 ( .A(n3057), .B(n3058), .Z(n3055) );
  NANDN U2676 ( .A(B[260]), .B(A[260]), .Z(n3058) );
  AND U2677 ( .A(n3059), .B(n3060), .Z(n3057) );
  NAND U2678 ( .A(n3061), .B(n3062), .Z(n3060) );
  NANDN U2679 ( .A(A[259]), .B(B[259]), .Z(n3062) );
  AND U2680 ( .A(n3063), .B(n3064), .Z(n3061) );
  NANDN U2681 ( .A(A[258]), .B(B[258]), .Z(n3064) );
  NAND U2682 ( .A(n3065), .B(n3066), .Z(n3063) );
  NANDN U2683 ( .A(B[258]), .B(A[258]), .Z(n3066) );
  AND U2684 ( .A(n3067), .B(n3068), .Z(n3065) );
  NAND U2685 ( .A(n3069), .B(n3070), .Z(n3068) );
  NANDN U2686 ( .A(A[257]), .B(B[257]), .Z(n3070) );
  AND U2687 ( .A(n3071), .B(n3072), .Z(n3069) );
  NANDN U2688 ( .A(A[256]), .B(B[256]), .Z(n3072) );
  NAND U2689 ( .A(n3073), .B(n3074), .Z(n3071) );
  NANDN U2690 ( .A(B[256]), .B(A[256]), .Z(n3074) );
  AND U2691 ( .A(n3075), .B(n3076), .Z(n3073) );
  NAND U2692 ( .A(n3077), .B(n3078), .Z(n3076) );
  NANDN U2693 ( .A(A[255]), .B(B[255]), .Z(n3078) );
  AND U2694 ( .A(n3079), .B(n3080), .Z(n3077) );
  NANDN U2695 ( .A(A[254]), .B(B[254]), .Z(n3080) );
  NAND U2696 ( .A(n3081), .B(n3082), .Z(n3079) );
  NANDN U2697 ( .A(B[254]), .B(A[254]), .Z(n3082) );
  AND U2698 ( .A(n3083), .B(n3084), .Z(n3081) );
  NAND U2699 ( .A(n3085), .B(n3086), .Z(n3084) );
  NANDN U2700 ( .A(A[253]), .B(B[253]), .Z(n3086) );
  AND U2701 ( .A(n3087), .B(n3088), .Z(n3085) );
  NANDN U2702 ( .A(A[252]), .B(B[252]), .Z(n3088) );
  NAND U2703 ( .A(n3089), .B(n3090), .Z(n3087) );
  NANDN U2704 ( .A(B[252]), .B(A[252]), .Z(n3090) );
  AND U2705 ( .A(n3091), .B(n3092), .Z(n3089) );
  NAND U2706 ( .A(n3093), .B(n3094), .Z(n3092) );
  NANDN U2707 ( .A(A[251]), .B(B[251]), .Z(n3094) );
  AND U2708 ( .A(n3095), .B(n3096), .Z(n3093) );
  NANDN U2709 ( .A(A[250]), .B(B[250]), .Z(n3096) );
  NAND U2710 ( .A(n3097), .B(n3098), .Z(n3095) );
  NANDN U2711 ( .A(B[250]), .B(A[250]), .Z(n3098) );
  AND U2712 ( .A(n3099), .B(n3100), .Z(n3097) );
  NAND U2713 ( .A(n3101), .B(n3102), .Z(n3100) );
  NANDN U2714 ( .A(A[249]), .B(B[249]), .Z(n3102) );
  AND U2715 ( .A(n3103), .B(n3104), .Z(n3101) );
  NANDN U2716 ( .A(A[248]), .B(B[248]), .Z(n3104) );
  NAND U2717 ( .A(n3105), .B(n3106), .Z(n3103) );
  NANDN U2718 ( .A(B[248]), .B(A[248]), .Z(n3106) );
  AND U2719 ( .A(n3107), .B(n3108), .Z(n3105) );
  NAND U2720 ( .A(n3109), .B(n3110), .Z(n3108) );
  NANDN U2721 ( .A(A[247]), .B(B[247]), .Z(n3110) );
  AND U2722 ( .A(n3111), .B(n3112), .Z(n3109) );
  NANDN U2723 ( .A(A[246]), .B(B[246]), .Z(n3112) );
  NAND U2724 ( .A(n3113), .B(n3114), .Z(n3111) );
  NANDN U2725 ( .A(B[246]), .B(A[246]), .Z(n3114) );
  AND U2726 ( .A(n3115), .B(n3116), .Z(n3113) );
  NAND U2727 ( .A(n3117), .B(n3118), .Z(n3116) );
  NANDN U2728 ( .A(A[245]), .B(B[245]), .Z(n3118) );
  AND U2729 ( .A(n3119), .B(n3120), .Z(n3117) );
  NANDN U2730 ( .A(A[244]), .B(B[244]), .Z(n3120) );
  NAND U2731 ( .A(n3121), .B(n3122), .Z(n3119) );
  NANDN U2732 ( .A(B[244]), .B(A[244]), .Z(n3122) );
  AND U2733 ( .A(n3123), .B(n3124), .Z(n3121) );
  NAND U2734 ( .A(n3125), .B(n3126), .Z(n3124) );
  NANDN U2735 ( .A(A[243]), .B(B[243]), .Z(n3126) );
  AND U2736 ( .A(n3127), .B(n3128), .Z(n3125) );
  NANDN U2737 ( .A(A[242]), .B(B[242]), .Z(n3128) );
  NAND U2738 ( .A(n3129), .B(n3130), .Z(n3127) );
  NANDN U2739 ( .A(B[242]), .B(A[242]), .Z(n3130) );
  AND U2740 ( .A(n3131), .B(n3132), .Z(n3129) );
  NAND U2741 ( .A(n3133), .B(n3134), .Z(n3132) );
  NANDN U2742 ( .A(A[241]), .B(B[241]), .Z(n3134) );
  AND U2743 ( .A(n3135), .B(n3136), .Z(n3133) );
  NANDN U2744 ( .A(A[240]), .B(B[240]), .Z(n3136) );
  NAND U2745 ( .A(n3137), .B(n3138), .Z(n3135) );
  NANDN U2746 ( .A(B[240]), .B(A[240]), .Z(n3138) );
  AND U2747 ( .A(n3139), .B(n3140), .Z(n3137) );
  NAND U2748 ( .A(n3141), .B(n3142), .Z(n3140) );
  NANDN U2749 ( .A(A[239]), .B(B[239]), .Z(n3142) );
  AND U2750 ( .A(n3143), .B(n3144), .Z(n3141) );
  NANDN U2751 ( .A(A[238]), .B(B[238]), .Z(n3144) );
  NAND U2752 ( .A(n3145), .B(n3146), .Z(n3143) );
  NANDN U2753 ( .A(B[238]), .B(A[238]), .Z(n3146) );
  AND U2754 ( .A(n3147), .B(n3148), .Z(n3145) );
  NAND U2755 ( .A(n3149), .B(n3150), .Z(n3148) );
  NANDN U2756 ( .A(A[237]), .B(B[237]), .Z(n3150) );
  AND U2757 ( .A(n3151), .B(n3152), .Z(n3149) );
  NANDN U2758 ( .A(A[236]), .B(B[236]), .Z(n3152) );
  NAND U2759 ( .A(n3153), .B(n3154), .Z(n3151) );
  NANDN U2760 ( .A(B[236]), .B(A[236]), .Z(n3154) );
  AND U2761 ( .A(n3155), .B(n3156), .Z(n3153) );
  NAND U2762 ( .A(n3157), .B(n3158), .Z(n3156) );
  NANDN U2763 ( .A(A[235]), .B(B[235]), .Z(n3158) );
  AND U2764 ( .A(n3159), .B(n3160), .Z(n3157) );
  NANDN U2765 ( .A(A[234]), .B(B[234]), .Z(n3160) );
  NAND U2766 ( .A(n3161), .B(n3162), .Z(n3159) );
  NANDN U2767 ( .A(B[234]), .B(A[234]), .Z(n3162) );
  AND U2768 ( .A(n3163), .B(n3164), .Z(n3161) );
  NAND U2769 ( .A(n3165), .B(n3166), .Z(n3164) );
  NANDN U2770 ( .A(A[233]), .B(B[233]), .Z(n3166) );
  AND U2771 ( .A(n3167), .B(n3168), .Z(n3165) );
  NANDN U2772 ( .A(A[232]), .B(B[232]), .Z(n3168) );
  NAND U2773 ( .A(n3169), .B(n3170), .Z(n3167) );
  NANDN U2774 ( .A(B[232]), .B(A[232]), .Z(n3170) );
  AND U2775 ( .A(n3171), .B(n3172), .Z(n3169) );
  NAND U2776 ( .A(n3173), .B(n3174), .Z(n3172) );
  NANDN U2777 ( .A(A[231]), .B(B[231]), .Z(n3174) );
  AND U2778 ( .A(n3175), .B(n3176), .Z(n3173) );
  NANDN U2779 ( .A(A[230]), .B(B[230]), .Z(n3176) );
  NAND U2780 ( .A(n3177), .B(n3178), .Z(n3175) );
  NANDN U2781 ( .A(B[230]), .B(A[230]), .Z(n3178) );
  AND U2782 ( .A(n3179), .B(n3180), .Z(n3177) );
  NAND U2783 ( .A(n3181), .B(n3182), .Z(n3180) );
  NANDN U2784 ( .A(A[229]), .B(B[229]), .Z(n3182) );
  AND U2785 ( .A(n3183), .B(n3184), .Z(n3181) );
  NANDN U2786 ( .A(A[228]), .B(B[228]), .Z(n3184) );
  NAND U2787 ( .A(n3185), .B(n3186), .Z(n3183) );
  NANDN U2788 ( .A(B[228]), .B(A[228]), .Z(n3186) );
  AND U2789 ( .A(n3187), .B(n3188), .Z(n3185) );
  NAND U2790 ( .A(n3189), .B(n3190), .Z(n3188) );
  NANDN U2791 ( .A(A[227]), .B(B[227]), .Z(n3190) );
  AND U2792 ( .A(n3191), .B(n3192), .Z(n3189) );
  NANDN U2793 ( .A(A[226]), .B(B[226]), .Z(n3192) );
  NAND U2794 ( .A(n3193), .B(n3194), .Z(n3191) );
  NANDN U2795 ( .A(B[226]), .B(A[226]), .Z(n3194) );
  AND U2796 ( .A(n3195), .B(n3196), .Z(n3193) );
  NAND U2797 ( .A(n3197), .B(n3198), .Z(n3196) );
  NANDN U2798 ( .A(A[225]), .B(B[225]), .Z(n3198) );
  AND U2799 ( .A(n3199), .B(n3200), .Z(n3197) );
  NANDN U2800 ( .A(A[224]), .B(B[224]), .Z(n3200) );
  NAND U2801 ( .A(n3201), .B(n3202), .Z(n3199) );
  NANDN U2802 ( .A(B[224]), .B(A[224]), .Z(n3202) );
  AND U2803 ( .A(n3203), .B(n3204), .Z(n3201) );
  NAND U2804 ( .A(n3205), .B(n3206), .Z(n3204) );
  NANDN U2805 ( .A(A[223]), .B(B[223]), .Z(n3206) );
  AND U2806 ( .A(n3207), .B(n3208), .Z(n3205) );
  NANDN U2807 ( .A(A[222]), .B(B[222]), .Z(n3208) );
  NAND U2808 ( .A(n3209), .B(n3210), .Z(n3207) );
  NANDN U2809 ( .A(B[222]), .B(A[222]), .Z(n3210) );
  AND U2810 ( .A(n3211), .B(n3212), .Z(n3209) );
  NAND U2811 ( .A(n3213), .B(n3214), .Z(n3212) );
  NANDN U2812 ( .A(A[221]), .B(B[221]), .Z(n3214) );
  AND U2813 ( .A(n3215), .B(n3216), .Z(n3213) );
  NANDN U2814 ( .A(A[220]), .B(B[220]), .Z(n3216) );
  NAND U2815 ( .A(n3217), .B(n3218), .Z(n3215) );
  NANDN U2816 ( .A(B[220]), .B(A[220]), .Z(n3218) );
  AND U2817 ( .A(n3219), .B(n3220), .Z(n3217) );
  NAND U2818 ( .A(n3221), .B(n3222), .Z(n3220) );
  NANDN U2819 ( .A(A[219]), .B(B[219]), .Z(n3222) );
  AND U2820 ( .A(n3223), .B(n3224), .Z(n3221) );
  NANDN U2821 ( .A(A[218]), .B(B[218]), .Z(n3224) );
  NAND U2822 ( .A(n3225), .B(n3226), .Z(n3223) );
  NANDN U2823 ( .A(B[218]), .B(A[218]), .Z(n3226) );
  AND U2824 ( .A(n3227), .B(n3228), .Z(n3225) );
  NAND U2825 ( .A(n3229), .B(n3230), .Z(n3228) );
  NANDN U2826 ( .A(A[217]), .B(B[217]), .Z(n3230) );
  AND U2827 ( .A(n3231), .B(n3232), .Z(n3229) );
  NANDN U2828 ( .A(A[216]), .B(B[216]), .Z(n3232) );
  NAND U2829 ( .A(n3233), .B(n3234), .Z(n3231) );
  NANDN U2830 ( .A(B[216]), .B(A[216]), .Z(n3234) );
  AND U2831 ( .A(n3235), .B(n3236), .Z(n3233) );
  NAND U2832 ( .A(n3237), .B(n3238), .Z(n3236) );
  NANDN U2833 ( .A(A[215]), .B(B[215]), .Z(n3238) );
  AND U2834 ( .A(n3239), .B(n3240), .Z(n3237) );
  NANDN U2835 ( .A(A[214]), .B(B[214]), .Z(n3240) );
  NAND U2836 ( .A(n3241), .B(n3242), .Z(n3239) );
  NANDN U2837 ( .A(B[214]), .B(A[214]), .Z(n3242) );
  AND U2838 ( .A(n3243), .B(n3244), .Z(n3241) );
  NAND U2839 ( .A(n3245), .B(n3246), .Z(n3244) );
  NANDN U2840 ( .A(A[213]), .B(B[213]), .Z(n3246) );
  AND U2841 ( .A(n3247), .B(n3248), .Z(n3245) );
  NANDN U2842 ( .A(A[212]), .B(B[212]), .Z(n3248) );
  NAND U2843 ( .A(n3249), .B(n3250), .Z(n3247) );
  NANDN U2844 ( .A(B[212]), .B(A[212]), .Z(n3250) );
  AND U2845 ( .A(n3251), .B(n3252), .Z(n3249) );
  NAND U2846 ( .A(n3253), .B(n3254), .Z(n3252) );
  NANDN U2847 ( .A(A[211]), .B(B[211]), .Z(n3254) );
  AND U2848 ( .A(n3255), .B(n3256), .Z(n3253) );
  NANDN U2849 ( .A(A[210]), .B(B[210]), .Z(n3256) );
  NAND U2850 ( .A(n3257), .B(n3258), .Z(n3255) );
  NANDN U2851 ( .A(B[210]), .B(A[210]), .Z(n3258) );
  AND U2852 ( .A(n3259), .B(n3260), .Z(n3257) );
  NAND U2853 ( .A(n3261), .B(n3262), .Z(n3260) );
  NANDN U2854 ( .A(A[209]), .B(B[209]), .Z(n3262) );
  AND U2855 ( .A(n3263), .B(n3264), .Z(n3261) );
  NANDN U2856 ( .A(A[208]), .B(B[208]), .Z(n3264) );
  NAND U2857 ( .A(n3265), .B(n3266), .Z(n3263) );
  NANDN U2858 ( .A(B[208]), .B(A[208]), .Z(n3266) );
  AND U2859 ( .A(n3267), .B(n3268), .Z(n3265) );
  NAND U2860 ( .A(n3269), .B(n3270), .Z(n3268) );
  NANDN U2861 ( .A(A[207]), .B(B[207]), .Z(n3270) );
  AND U2862 ( .A(n3271), .B(n3272), .Z(n3269) );
  NANDN U2863 ( .A(A[206]), .B(B[206]), .Z(n3272) );
  NAND U2864 ( .A(n3273), .B(n3274), .Z(n3271) );
  NANDN U2865 ( .A(B[206]), .B(A[206]), .Z(n3274) );
  AND U2866 ( .A(n3275), .B(n3276), .Z(n3273) );
  NAND U2867 ( .A(n3277), .B(n3278), .Z(n3276) );
  NANDN U2868 ( .A(A[205]), .B(B[205]), .Z(n3278) );
  AND U2869 ( .A(n3279), .B(n3280), .Z(n3277) );
  NANDN U2870 ( .A(A[204]), .B(B[204]), .Z(n3280) );
  NAND U2871 ( .A(n3281), .B(n3282), .Z(n3279) );
  NANDN U2872 ( .A(B[204]), .B(A[204]), .Z(n3282) );
  AND U2873 ( .A(n3283), .B(n3284), .Z(n3281) );
  NAND U2874 ( .A(n3285), .B(n3286), .Z(n3284) );
  NANDN U2875 ( .A(A[203]), .B(B[203]), .Z(n3286) );
  AND U2876 ( .A(n3287), .B(n3288), .Z(n3285) );
  NANDN U2877 ( .A(A[202]), .B(B[202]), .Z(n3288) );
  NAND U2878 ( .A(n3289), .B(n3290), .Z(n3287) );
  NANDN U2879 ( .A(B[202]), .B(A[202]), .Z(n3290) );
  AND U2880 ( .A(n3291), .B(n3292), .Z(n3289) );
  NAND U2881 ( .A(n3293), .B(n3294), .Z(n3292) );
  NANDN U2882 ( .A(A[201]), .B(B[201]), .Z(n3294) );
  AND U2883 ( .A(n3295), .B(n3296), .Z(n3293) );
  NANDN U2884 ( .A(A[200]), .B(B[200]), .Z(n3296) );
  NAND U2885 ( .A(n3297), .B(n3298), .Z(n3295) );
  NANDN U2886 ( .A(B[200]), .B(A[200]), .Z(n3298) );
  AND U2887 ( .A(n3299), .B(n3300), .Z(n3297) );
  NAND U2888 ( .A(n3301), .B(n3302), .Z(n3300) );
  NANDN U2889 ( .A(A[199]), .B(B[199]), .Z(n3302) );
  AND U2890 ( .A(n3303), .B(n3304), .Z(n3301) );
  NANDN U2891 ( .A(A[198]), .B(B[198]), .Z(n3304) );
  NAND U2892 ( .A(n3305), .B(n3306), .Z(n3303) );
  NANDN U2893 ( .A(B[198]), .B(A[198]), .Z(n3306) );
  AND U2894 ( .A(n3307), .B(n3308), .Z(n3305) );
  NAND U2895 ( .A(n3309), .B(n3310), .Z(n3308) );
  NANDN U2896 ( .A(A[197]), .B(B[197]), .Z(n3310) );
  AND U2897 ( .A(n3311), .B(n3312), .Z(n3309) );
  NANDN U2898 ( .A(A[196]), .B(B[196]), .Z(n3312) );
  NAND U2899 ( .A(n3313), .B(n3314), .Z(n3311) );
  NANDN U2900 ( .A(B[196]), .B(A[196]), .Z(n3314) );
  AND U2901 ( .A(n3315), .B(n3316), .Z(n3313) );
  NAND U2902 ( .A(n3317), .B(n3318), .Z(n3316) );
  NANDN U2903 ( .A(A[195]), .B(B[195]), .Z(n3318) );
  AND U2904 ( .A(n3319), .B(n3320), .Z(n3317) );
  NANDN U2905 ( .A(A[194]), .B(B[194]), .Z(n3320) );
  NAND U2906 ( .A(n3321), .B(n3322), .Z(n3319) );
  NANDN U2907 ( .A(B[194]), .B(A[194]), .Z(n3322) );
  AND U2908 ( .A(n3323), .B(n3324), .Z(n3321) );
  NAND U2909 ( .A(n3325), .B(n3326), .Z(n3324) );
  NANDN U2910 ( .A(A[193]), .B(B[193]), .Z(n3326) );
  AND U2911 ( .A(n3327), .B(n3328), .Z(n3325) );
  NANDN U2912 ( .A(A[192]), .B(B[192]), .Z(n3328) );
  NAND U2913 ( .A(n3329), .B(n3330), .Z(n3327) );
  NANDN U2914 ( .A(B[192]), .B(A[192]), .Z(n3330) );
  AND U2915 ( .A(n3331), .B(n3332), .Z(n3329) );
  NAND U2916 ( .A(n3333), .B(n3334), .Z(n3332) );
  NANDN U2917 ( .A(A[191]), .B(B[191]), .Z(n3334) );
  AND U2918 ( .A(n3335), .B(n3336), .Z(n3333) );
  NANDN U2919 ( .A(A[190]), .B(B[190]), .Z(n3336) );
  NAND U2920 ( .A(n3337), .B(n3338), .Z(n3335) );
  NANDN U2921 ( .A(B[190]), .B(A[190]), .Z(n3338) );
  AND U2922 ( .A(n3339), .B(n3340), .Z(n3337) );
  NAND U2923 ( .A(n3341), .B(n3342), .Z(n3340) );
  NANDN U2924 ( .A(A[189]), .B(B[189]), .Z(n3342) );
  AND U2925 ( .A(n3343), .B(n3344), .Z(n3341) );
  NANDN U2926 ( .A(A[188]), .B(B[188]), .Z(n3344) );
  NAND U2927 ( .A(n3345), .B(n3346), .Z(n3343) );
  NANDN U2928 ( .A(B[188]), .B(A[188]), .Z(n3346) );
  AND U2929 ( .A(n3347), .B(n3348), .Z(n3345) );
  NAND U2930 ( .A(n3349), .B(n3350), .Z(n3348) );
  NANDN U2931 ( .A(A[187]), .B(B[187]), .Z(n3350) );
  AND U2932 ( .A(n3351), .B(n3352), .Z(n3349) );
  NANDN U2933 ( .A(A[186]), .B(B[186]), .Z(n3352) );
  NAND U2934 ( .A(n3353), .B(n3354), .Z(n3351) );
  NANDN U2935 ( .A(B[186]), .B(A[186]), .Z(n3354) );
  AND U2936 ( .A(n3355), .B(n3356), .Z(n3353) );
  NAND U2937 ( .A(n3357), .B(n3358), .Z(n3356) );
  NANDN U2938 ( .A(A[185]), .B(B[185]), .Z(n3358) );
  AND U2939 ( .A(n3359), .B(n3360), .Z(n3357) );
  NANDN U2940 ( .A(A[184]), .B(B[184]), .Z(n3360) );
  NAND U2941 ( .A(n3361), .B(n3362), .Z(n3359) );
  NANDN U2942 ( .A(B[184]), .B(A[184]), .Z(n3362) );
  AND U2943 ( .A(n3363), .B(n3364), .Z(n3361) );
  NAND U2944 ( .A(n3365), .B(n3366), .Z(n3364) );
  NANDN U2945 ( .A(A[183]), .B(B[183]), .Z(n3366) );
  AND U2946 ( .A(n3367), .B(n3368), .Z(n3365) );
  NANDN U2947 ( .A(A[182]), .B(B[182]), .Z(n3368) );
  NAND U2948 ( .A(n3369), .B(n3370), .Z(n3367) );
  NANDN U2949 ( .A(B[182]), .B(A[182]), .Z(n3370) );
  AND U2950 ( .A(n3371), .B(n3372), .Z(n3369) );
  NAND U2951 ( .A(n3373), .B(n3374), .Z(n3372) );
  NANDN U2952 ( .A(A[181]), .B(B[181]), .Z(n3374) );
  AND U2953 ( .A(n3375), .B(n3376), .Z(n3373) );
  NANDN U2954 ( .A(A[180]), .B(B[180]), .Z(n3376) );
  NAND U2955 ( .A(n3377), .B(n3378), .Z(n3375) );
  NANDN U2956 ( .A(B[180]), .B(A[180]), .Z(n3378) );
  AND U2957 ( .A(n3379), .B(n3380), .Z(n3377) );
  NAND U2958 ( .A(n3381), .B(n3382), .Z(n3380) );
  NANDN U2959 ( .A(A[179]), .B(B[179]), .Z(n3382) );
  AND U2960 ( .A(n3383), .B(n3384), .Z(n3381) );
  NANDN U2961 ( .A(A[178]), .B(B[178]), .Z(n3384) );
  NAND U2962 ( .A(n3385), .B(n3386), .Z(n3383) );
  NANDN U2963 ( .A(B[178]), .B(A[178]), .Z(n3386) );
  AND U2964 ( .A(n3387), .B(n3388), .Z(n3385) );
  NAND U2965 ( .A(n3389), .B(n3390), .Z(n3388) );
  NANDN U2966 ( .A(A[177]), .B(B[177]), .Z(n3390) );
  AND U2967 ( .A(n3391), .B(n3392), .Z(n3389) );
  NANDN U2968 ( .A(A[176]), .B(B[176]), .Z(n3392) );
  NAND U2969 ( .A(n3393), .B(n3394), .Z(n3391) );
  NANDN U2970 ( .A(B[176]), .B(A[176]), .Z(n3394) );
  AND U2971 ( .A(n3395), .B(n3396), .Z(n3393) );
  NAND U2972 ( .A(n3397), .B(n3398), .Z(n3396) );
  NANDN U2973 ( .A(A[175]), .B(B[175]), .Z(n3398) );
  AND U2974 ( .A(n3399), .B(n3400), .Z(n3397) );
  NANDN U2975 ( .A(A[174]), .B(B[174]), .Z(n3400) );
  NAND U2976 ( .A(n3401), .B(n3402), .Z(n3399) );
  NANDN U2977 ( .A(B[174]), .B(A[174]), .Z(n3402) );
  AND U2978 ( .A(n3403), .B(n3404), .Z(n3401) );
  NAND U2979 ( .A(n3405), .B(n3406), .Z(n3404) );
  NANDN U2980 ( .A(A[173]), .B(B[173]), .Z(n3406) );
  AND U2981 ( .A(n3407), .B(n3408), .Z(n3405) );
  NANDN U2982 ( .A(A[172]), .B(B[172]), .Z(n3408) );
  NAND U2983 ( .A(n3409), .B(n3410), .Z(n3407) );
  NANDN U2984 ( .A(B[172]), .B(A[172]), .Z(n3410) );
  AND U2985 ( .A(n3411), .B(n3412), .Z(n3409) );
  NAND U2986 ( .A(n3413), .B(n3414), .Z(n3412) );
  NANDN U2987 ( .A(A[171]), .B(B[171]), .Z(n3414) );
  AND U2988 ( .A(n3415), .B(n3416), .Z(n3413) );
  NANDN U2989 ( .A(A[170]), .B(B[170]), .Z(n3416) );
  NAND U2990 ( .A(n3417), .B(n3418), .Z(n3415) );
  NANDN U2991 ( .A(B[170]), .B(A[170]), .Z(n3418) );
  AND U2992 ( .A(n3419), .B(n3420), .Z(n3417) );
  NAND U2993 ( .A(n3421), .B(n3422), .Z(n3420) );
  NANDN U2994 ( .A(A[169]), .B(B[169]), .Z(n3422) );
  AND U2995 ( .A(n3423), .B(n3424), .Z(n3421) );
  NANDN U2996 ( .A(A[168]), .B(B[168]), .Z(n3424) );
  NAND U2997 ( .A(n3425), .B(n3426), .Z(n3423) );
  NANDN U2998 ( .A(B[168]), .B(A[168]), .Z(n3426) );
  AND U2999 ( .A(n3427), .B(n3428), .Z(n3425) );
  NAND U3000 ( .A(n3429), .B(n3430), .Z(n3428) );
  NANDN U3001 ( .A(A[167]), .B(B[167]), .Z(n3430) );
  AND U3002 ( .A(n3431), .B(n3432), .Z(n3429) );
  NANDN U3003 ( .A(A[166]), .B(B[166]), .Z(n3432) );
  NAND U3004 ( .A(n3433), .B(n3434), .Z(n3431) );
  NANDN U3005 ( .A(B[166]), .B(A[166]), .Z(n3434) );
  AND U3006 ( .A(n3435), .B(n3436), .Z(n3433) );
  NAND U3007 ( .A(n3437), .B(n3438), .Z(n3436) );
  NANDN U3008 ( .A(A[165]), .B(B[165]), .Z(n3438) );
  AND U3009 ( .A(n3439), .B(n3440), .Z(n3437) );
  NANDN U3010 ( .A(A[164]), .B(B[164]), .Z(n3440) );
  NAND U3011 ( .A(n3441), .B(n3442), .Z(n3439) );
  NANDN U3012 ( .A(B[164]), .B(A[164]), .Z(n3442) );
  AND U3013 ( .A(n3443), .B(n3444), .Z(n3441) );
  NAND U3014 ( .A(n3445), .B(n3446), .Z(n3444) );
  NANDN U3015 ( .A(A[163]), .B(B[163]), .Z(n3446) );
  AND U3016 ( .A(n3447), .B(n3448), .Z(n3445) );
  NANDN U3017 ( .A(A[162]), .B(B[162]), .Z(n3448) );
  NAND U3018 ( .A(n3449), .B(n3450), .Z(n3447) );
  NANDN U3019 ( .A(B[162]), .B(A[162]), .Z(n3450) );
  AND U3020 ( .A(n3451), .B(n3452), .Z(n3449) );
  NAND U3021 ( .A(n3453), .B(n3454), .Z(n3452) );
  NANDN U3022 ( .A(A[161]), .B(B[161]), .Z(n3454) );
  AND U3023 ( .A(n3455), .B(n3456), .Z(n3453) );
  NANDN U3024 ( .A(A[160]), .B(B[160]), .Z(n3456) );
  NAND U3025 ( .A(n3457), .B(n3458), .Z(n3455) );
  NANDN U3026 ( .A(B[160]), .B(A[160]), .Z(n3458) );
  AND U3027 ( .A(n3459), .B(n3460), .Z(n3457) );
  NAND U3028 ( .A(n3461), .B(n3462), .Z(n3460) );
  NANDN U3029 ( .A(A[159]), .B(B[159]), .Z(n3462) );
  AND U3030 ( .A(n3463), .B(n3464), .Z(n3461) );
  NANDN U3031 ( .A(A[158]), .B(B[158]), .Z(n3464) );
  NAND U3032 ( .A(n3465), .B(n3466), .Z(n3463) );
  NANDN U3033 ( .A(B[158]), .B(A[158]), .Z(n3466) );
  AND U3034 ( .A(n3467), .B(n3468), .Z(n3465) );
  NAND U3035 ( .A(n3469), .B(n3470), .Z(n3468) );
  NANDN U3036 ( .A(A[157]), .B(B[157]), .Z(n3470) );
  AND U3037 ( .A(n3471), .B(n3472), .Z(n3469) );
  NANDN U3038 ( .A(A[156]), .B(B[156]), .Z(n3472) );
  NAND U3039 ( .A(n3473), .B(n3474), .Z(n3471) );
  NANDN U3040 ( .A(B[156]), .B(A[156]), .Z(n3474) );
  AND U3041 ( .A(n3475), .B(n3476), .Z(n3473) );
  NAND U3042 ( .A(n3477), .B(n3478), .Z(n3476) );
  NANDN U3043 ( .A(A[155]), .B(B[155]), .Z(n3478) );
  AND U3044 ( .A(n3479), .B(n3480), .Z(n3477) );
  NANDN U3045 ( .A(A[154]), .B(B[154]), .Z(n3480) );
  NAND U3046 ( .A(n3481), .B(n3482), .Z(n3479) );
  NANDN U3047 ( .A(B[154]), .B(A[154]), .Z(n3482) );
  AND U3048 ( .A(n3483), .B(n3484), .Z(n3481) );
  NAND U3049 ( .A(n3485), .B(n3486), .Z(n3484) );
  NANDN U3050 ( .A(A[153]), .B(B[153]), .Z(n3486) );
  AND U3051 ( .A(n3487), .B(n3488), .Z(n3485) );
  NANDN U3052 ( .A(A[152]), .B(B[152]), .Z(n3488) );
  NAND U3053 ( .A(n3489), .B(n3490), .Z(n3487) );
  NANDN U3054 ( .A(B[152]), .B(A[152]), .Z(n3490) );
  AND U3055 ( .A(n3491), .B(n3492), .Z(n3489) );
  NAND U3056 ( .A(n3493), .B(n3494), .Z(n3492) );
  NANDN U3057 ( .A(A[151]), .B(B[151]), .Z(n3494) );
  AND U3058 ( .A(n3495), .B(n3496), .Z(n3493) );
  NANDN U3059 ( .A(A[150]), .B(B[150]), .Z(n3496) );
  NAND U3060 ( .A(n3497), .B(n3498), .Z(n3495) );
  NANDN U3061 ( .A(B[150]), .B(A[150]), .Z(n3498) );
  AND U3062 ( .A(n3499), .B(n3500), .Z(n3497) );
  NAND U3063 ( .A(n3501), .B(n3502), .Z(n3500) );
  NANDN U3064 ( .A(A[149]), .B(B[149]), .Z(n3502) );
  AND U3065 ( .A(n3503), .B(n3504), .Z(n3501) );
  NANDN U3066 ( .A(A[148]), .B(B[148]), .Z(n3504) );
  NAND U3067 ( .A(n3505), .B(n3506), .Z(n3503) );
  NANDN U3068 ( .A(B[148]), .B(A[148]), .Z(n3506) );
  AND U3069 ( .A(n3507), .B(n3508), .Z(n3505) );
  NAND U3070 ( .A(n3509), .B(n3510), .Z(n3508) );
  NANDN U3071 ( .A(A[147]), .B(B[147]), .Z(n3510) );
  AND U3072 ( .A(n3511), .B(n3512), .Z(n3509) );
  NANDN U3073 ( .A(A[146]), .B(B[146]), .Z(n3512) );
  NAND U3074 ( .A(n3513), .B(n3514), .Z(n3511) );
  NANDN U3075 ( .A(B[146]), .B(A[146]), .Z(n3514) );
  AND U3076 ( .A(n3515), .B(n3516), .Z(n3513) );
  NAND U3077 ( .A(n3517), .B(n3518), .Z(n3516) );
  NANDN U3078 ( .A(A[145]), .B(B[145]), .Z(n3518) );
  AND U3079 ( .A(n3519), .B(n3520), .Z(n3517) );
  NANDN U3080 ( .A(A[144]), .B(B[144]), .Z(n3520) );
  NAND U3081 ( .A(n3521), .B(n3522), .Z(n3519) );
  NANDN U3082 ( .A(B[144]), .B(A[144]), .Z(n3522) );
  AND U3083 ( .A(n3523), .B(n3524), .Z(n3521) );
  NAND U3084 ( .A(n3525), .B(n3526), .Z(n3524) );
  NANDN U3085 ( .A(A[143]), .B(B[143]), .Z(n3526) );
  AND U3086 ( .A(n3527), .B(n3528), .Z(n3525) );
  NANDN U3087 ( .A(A[142]), .B(B[142]), .Z(n3528) );
  NAND U3088 ( .A(n3529), .B(n3530), .Z(n3527) );
  NANDN U3089 ( .A(B[142]), .B(A[142]), .Z(n3530) );
  AND U3090 ( .A(n3531), .B(n3532), .Z(n3529) );
  NAND U3091 ( .A(n3533), .B(n3534), .Z(n3532) );
  NANDN U3092 ( .A(A[141]), .B(B[141]), .Z(n3534) );
  AND U3093 ( .A(n3535), .B(n3536), .Z(n3533) );
  NANDN U3094 ( .A(A[140]), .B(B[140]), .Z(n3536) );
  NAND U3095 ( .A(n3537), .B(n3538), .Z(n3535) );
  NANDN U3096 ( .A(B[140]), .B(A[140]), .Z(n3538) );
  AND U3097 ( .A(n3539), .B(n3540), .Z(n3537) );
  NAND U3098 ( .A(n3541), .B(n3542), .Z(n3540) );
  NANDN U3099 ( .A(A[139]), .B(B[139]), .Z(n3542) );
  AND U3100 ( .A(n3543), .B(n3544), .Z(n3541) );
  NANDN U3101 ( .A(A[138]), .B(B[138]), .Z(n3544) );
  NAND U3102 ( .A(n3545), .B(n3546), .Z(n3543) );
  NANDN U3103 ( .A(B[138]), .B(A[138]), .Z(n3546) );
  AND U3104 ( .A(n3547), .B(n3548), .Z(n3545) );
  NAND U3105 ( .A(n3549), .B(n3550), .Z(n3548) );
  NANDN U3106 ( .A(A[137]), .B(B[137]), .Z(n3550) );
  AND U3107 ( .A(n3551), .B(n3552), .Z(n3549) );
  NANDN U3108 ( .A(A[136]), .B(B[136]), .Z(n3552) );
  NAND U3109 ( .A(n3553), .B(n3554), .Z(n3551) );
  NANDN U3110 ( .A(B[136]), .B(A[136]), .Z(n3554) );
  AND U3111 ( .A(n3555), .B(n3556), .Z(n3553) );
  NAND U3112 ( .A(n3557), .B(n3558), .Z(n3556) );
  NANDN U3113 ( .A(A[135]), .B(B[135]), .Z(n3558) );
  AND U3114 ( .A(n3559), .B(n3560), .Z(n3557) );
  NANDN U3115 ( .A(A[134]), .B(B[134]), .Z(n3560) );
  NAND U3116 ( .A(n3561), .B(n3562), .Z(n3559) );
  NANDN U3117 ( .A(B[134]), .B(A[134]), .Z(n3562) );
  AND U3118 ( .A(n3563), .B(n3564), .Z(n3561) );
  NAND U3119 ( .A(n3565), .B(n3566), .Z(n3564) );
  NANDN U3120 ( .A(A[133]), .B(B[133]), .Z(n3566) );
  AND U3121 ( .A(n3567), .B(n3568), .Z(n3565) );
  NANDN U3122 ( .A(A[132]), .B(B[132]), .Z(n3568) );
  NAND U3123 ( .A(n3569), .B(n3570), .Z(n3567) );
  NANDN U3124 ( .A(B[132]), .B(A[132]), .Z(n3570) );
  AND U3125 ( .A(n3571), .B(n3572), .Z(n3569) );
  NAND U3126 ( .A(n3573), .B(n3574), .Z(n3572) );
  NANDN U3127 ( .A(A[131]), .B(B[131]), .Z(n3574) );
  AND U3128 ( .A(n3575), .B(n3576), .Z(n3573) );
  NANDN U3129 ( .A(A[130]), .B(B[130]), .Z(n3576) );
  NAND U3130 ( .A(n3577), .B(n3578), .Z(n3575) );
  NANDN U3131 ( .A(B[130]), .B(A[130]), .Z(n3578) );
  AND U3132 ( .A(n3579), .B(n3580), .Z(n3577) );
  NAND U3133 ( .A(n3581), .B(n3582), .Z(n3580) );
  NANDN U3134 ( .A(A[129]), .B(B[129]), .Z(n3582) );
  AND U3135 ( .A(n3583), .B(n3584), .Z(n3581) );
  NANDN U3136 ( .A(A[128]), .B(B[128]), .Z(n3584) );
  NAND U3137 ( .A(n3585), .B(n3586), .Z(n3583) );
  NANDN U3138 ( .A(B[128]), .B(A[128]), .Z(n3586) );
  AND U3139 ( .A(n3587), .B(n3588), .Z(n3585) );
  NAND U3140 ( .A(n3589), .B(n3590), .Z(n3588) );
  NANDN U3141 ( .A(A[127]), .B(B[127]), .Z(n3590) );
  AND U3142 ( .A(n3591), .B(n3592), .Z(n3589) );
  NANDN U3143 ( .A(A[126]), .B(B[126]), .Z(n3592) );
  NAND U3144 ( .A(n3593), .B(n3594), .Z(n3591) );
  NANDN U3145 ( .A(B[126]), .B(A[126]), .Z(n3594) );
  AND U3146 ( .A(n3595), .B(n3596), .Z(n3593) );
  NAND U3147 ( .A(n3597), .B(n3598), .Z(n3596) );
  NANDN U3148 ( .A(A[125]), .B(B[125]), .Z(n3598) );
  AND U3149 ( .A(n3599), .B(n3600), .Z(n3597) );
  NANDN U3150 ( .A(A[124]), .B(B[124]), .Z(n3600) );
  NAND U3151 ( .A(n3601), .B(n3602), .Z(n3599) );
  NANDN U3152 ( .A(B[124]), .B(A[124]), .Z(n3602) );
  AND U3153 ( .A(n3603), .B(n3604), .Z(n3601) );
  NAND U3154 ( .A(n3605), .B(n3606), .Z(n3604) );
  NANDN U3155 ( .A(A[123]), .B(B[123]), .Z(n3606) );
  AND U3156 ( .A(n3607), .B(n3608), .Z(n3605) );
  NANDN U3157 ( .A(A[122]), .B(B[122]), .Z(n3608) );
  NAND U3158 ( .A(n3609), .B(n3610), .Z(n3607) );
  NANDN U3159 ( .A(B[122]), .B(A[122]), .Z(n3610) );
  AND U3160 ( .A(n3611), .B(n3612), .Z(n3609) );
  NAND U3161 ( .A(n3613), .B(n3614), .Z(n3612) );
  NANDN U3162 ( .A(A[121]), .B(B[121]), .Z(n3614) );
  AND U3163 ( .A(n3615), .B(n3616), .Z(n3613) );
  NANDN U3164 ( .A(A[120]), .B(B[120]), .Z(n3616) );
  NAND U3165 ( .A(n3617), .B(n3618), .Z(n3615) );
  NANDN U3166 ( .A(B[120]), .B(A[120]), .Z(n3618) );
  AND U3167 ( .A(n3619), .B(n3620), .Z(n3617) );
  NAND U3168 ( .A(n3621), .B(n3622), .Z(n3620) );
  NANDN U3169 ( .A(A[119]), .B(B[119]), .Z(n3622) );
  AND U3170 ( .A(n3623), .B(n3624), .Z(n3621) );
  NANDN U3171 ( .A(A[118]), .B(B[118]), .Z(n3624) );
  NAND U3172 ( .A(n3625), .B(n3626), .Z(n3623) );
  NANDN U3173 ( .A(B[118]), .B(A[118]), .Z(n3626) );
  AND U3174 ( .A(n3627), .B(n3628), .Z(n3625) );
  NAND U3175 ( .A(n3629), .B(n3630), .Z(n3628) );
  NANDN U3176 ( .A(A[117]), .B(B[117]), .Z(n3630) );
  AND U3177 ( .A(n3631), .B(n3632), .Z(n3629) );
  NANDN U3178 ( .A(A[116]), .B(B[116]), .Z(n3632) );
  NAND U3179 ( .A(n3633), .B(n3634), .Z(n3631) );
  NANDN U3180 ( .A(B[116]), .B(A[116]), .Z(n3634) );
  AND U3181 ( .A(n3635), .B(n3636), .Z(n3633) );
  NAND U3182 ( .A(n3637), .B(n3638), .Z(n3636) );
  NANDN U3183 ( .A(A[115]), .B(B[115]), .Z(n3638) );
  AND U3184 ( .A(n3639), .B(n3640), .Z(n3637) );
  NANDN U3185 ( .A(A[114]), .B(B[114]), .Z(n3640) );
  NAND U3186 ( .A(n3641), .B(n3642), .Z(n3639) );
  NANDN U3187 ( .A(B[114]), .B(A[114]), .Z(n3642) );
  AND U3188 ( .A(n3643), .B(n3644), .Z(n3641) );
  NAND U3189 ( .A(n3645), .B(n3646), .Z(n3644) );
  NANDN U3190 ( .A(A[113]), .B(B[113]), .Z(n3646) );
  AND U3191 ( .A(n3647), .B(n3648), .Z(n3645) );
  NANDN U3192 ( .A(A[112]), .B(B[112]), .Z(n3648) );
  NAND U3193 ( .A(n3649), .B(n3650), .Z(n3647) );
  NANDN U3194 ( .A(B[112]), .B(A[112]), .Z(n3650) );
  AND U3195 ( .A(n3651), .B(n3652), .Z(n3649) );
  NAND U3196 ( .A(n3653), .B(n3654), .Z(n3652) );
  NANDN U3197 ( .A(A[111]), .B(B[111]), .Z(n3654) );
  AND U3198 ( .A(n3655), .B(n3656), .Z(n3653) );
  NANDN U3199 ( .A(A[110]), .B(B[110]), .Z(n3656) );
  NAND U3200 ( .A(n3657), .B(n3658), .Z(n3655) );
  NANDN U3201 ( .A(B[110]), .B(A[110]), .Z(n3658) );
  AND U3202 ( .A(n3659), .B(n3660), .Z(n3657) );
  NAND U3203 ( .A(n3661), .B(n3662), .Z(n3660) );
  NANDN U3204 ( .A(A[109]), .B(B[109]), .Z(n3662) );
  AND U3205 ( .A(n3663), .B(n3664), .Z(n3661) );
  NANDN U3206 ( .A(A[108]), .B(B[108]), .Z(n3664) );
  NAND U3207 ( .A(n3665), .B(n3666), .Z(n3663) );
  NANDN U3208 ( .A(B[108]), .B(A[108]), .Z(n3666) );
  AND U3209 ( .A(n3667), .B(n3668), .Z(n3665) );
  NAND U3210 ( .A(n3669), .B(n3670), .Z(n3668) );
  NANDN U3211 ( .A(A[107]), .B(B[107]), .Z(n3670) );
  AND U3212 ( .A(n3671), .B(n3672), .Z(n3669) );
  NANDN U3213 ( .A(A[106]), .B(B[106]), .Z(n3672) );
  NAND U3214 ( .A(n3673), .B(n3674), .Z(n3671) );
  NANDN U3215 ( .A(B[106]), .B(A[106]), .Z(n3674) );
  AND U3216 ( .A(n3675), .B(n3676), .Z(n3673) );
  NAND U3217 ( .A(n3677), .B(n3678), .Z(n3676) );
  NANDN U3218 ( .A(A[105]), .B(B[105]), .Z(n3678) );
  AND U3219 ( .A(n3679), .B(n3680), .Z(n3677) );
  NANDN U3220 ( .A(A[104]), .B(B[104]), .Z(n3680) );
  NAND U3221 ( .A(n3681), .B(n3682), .Z(n3679) );
  NANDN U3222 ( .A(B[104]), .B(A[104]), .Z(n3682) );
  AND U3223 ( .A(n3683), .B(n3684), .Z(n3681) );
  NAND U3224 ( .A(n3685), .B(n3686), .Z(n3684) );
  NANDN U3225 ( .A(A[103]), .B(B[103]), .Z(n3686) );
  AND U3226 ( .A(n3687), .B(n3688), .Z(n3685) );
  NANDN U3227 ( .A(A[102]), .B(B[102]), .Z(n3688) );
  NAND U3228 ( .A(n3689), .B(n3690), .Z(n3687) );
  NANDN U3229 ( .A(B[102]), .B(A[102]), .Z(n3690) );
  AND U3230 ( .A(n3691), .B(n3692), .Z(n3689) );
  NAND U3231 ( .A(n3693), .B(n3694), .Z(n3692) );
  NANDN U3232 ( .A(A[101]), .B(B[101]), .Z(n3694) );
  AND U3233 ( .A(n3695), .B(n3696), .Z(n3693) );
  NANDN U3234 ( .A(A[100]), .B(B[100]), .Z(n3696) );
  NAND U3235 ( .A(n3697), .B(n3698), .Z(n3695) );
  NANDN U3236 ( .A(B[99]), .B(A[99]), .Z(n3698) );
  AND U3237 ( .A(n3699), .B(n3700), .Z(n3697) );
  NAND U3238 ( .A(n3701), .B(n3702), .Z(n3700) );
  NANDN U3239 ( .A(A[99]), .B(B[99]), .Z(n3702) );
  AND U3240 ( .A(n3703), .B(n3704), .Z(n3701) );
  NANDN U3241 ( .A(A[98]), .B(B[98]), .Z(n3704) );
  NAND U3242 ( .A(n3705), .B(n3706), .Z(n3703) );
  NANDN U3243 ( .A(B[98]), .B(A[98]), .Z(n3706) );
  AND U3244 ( .A(n3707), .B(n3708), .Z(n3705) );
  NAND U3245 ( .A(n3709), .B(n3710), .Z(n3708) );
  NANDN U3246 ( .A(A[97]), .B(B[97]), .Z(n3710) );
  AND U3247 ( .A(n3711), .B(n3712), .Z(n3709) );
  NANDN U3248 ( .A(A[96]), .B(B[96]), .Z(n3712) );
  NAND U3249 ( .A(n3713), .B(n3714), .Z(n3711) );
  NANDN U3250 ( .A(B[96]), .B(A[96]), .Z(n3714) );
  AND U3251 ( .A(n3715), .B(n3716), .Z(n3713) );
  NAND U3252 ( .A(n3717), .B(n3718), .Z(n3716) );
  NANDN U3253 ( .A(A[95]), .B(B[95]), .Z(n3718) );
  AND U3254 ( .A(n3719), .B(n3720), .Z(n3717) );
  NANDN U3255 ( .A(A[94]), .B(B[94]), .Z(n3720) );
  NAND U3256 ( .A(n3721), .B(n3722), .Z(n3719) );
  NANDN U3257 ( .A(B[94]), .B(A[94]), .Z(n3722) );
  AND U3258 ( .A(n3723), .B(n3724), .Z(n3721) );
  NAND U3259 ( .A(n3725), .B(n3726), .Z(n3724) );
  NANDN U3260 ( .A(A[93]), .B(B[93]), .Z(n3726) );
  AND U3261 ( .A(n3727), .B(n3728), .Z(n3725) );
  NANDN U3262 ( .A(A[92]), .B(B[92]), .Z(n3728) );
  NAND U3263 ( .A(n3729), .B(n3730), .Z(n3727) );
  NANDN U3264 ( .A(B[92]), .B(A[92]), .Z(n3730) );
  AND U3265 ( .A(n3731), .B(n3732), .Z(n3729) );
  NAND U3266 ( .A(n3733), .B(n3734), .Z(n3732) );
  NANDN U3267 ( .A(A[91]), .B(B[91]), .Z(n3734) );
  AND U3268 ( .A(n3735), .B(n3736), .Z(n3733) );
  NANDN U3269 ( .A(A[90]), .B(B[90]), .Z(n3736) );
  NAND U3270 ( .A(n3737), .B(n3738), .Z(n3735) );
  NANDN U3271 ( .A(B[90]), .B(A[90]), .Z(n3738) );
  AND U3272 ( .A(n3739), .B(n3740), .Z(n3737) );
  NAND U3273 ( .A(n3741), .B(n3742), .Z(n3740) );
  NANDN U3274 ( .A(A[89]), .B(B[89]), .Z(n3742) );
  AND U3275 ( .A(n3743), .B(n3744), .Z(n3741) );
  NANDN U3276 ( .A(A[88]), .B(B[88]), .Z(n3744) );
  NAND U3277 ( .A(n3745), .B(n3746), .Z(n3743) );
  NANDN U3278 ( .A(B[88]), .B(A[88]), .Z(n3746) );
  AND U3279 ( .A(n3747), .B(n3748), .Z(n3745) );
  NAND U3280 ( .A(n3749), .B(n3750), .Z(n3748) );
  NANDN U3281 ( .A(A[87]), .B(B[87]), .Z(n3750) );
  AND U3282 ( .A(n3751), .B(n3752), .Z(n3749) );
  NANDN U3283 ( .A(A[86]), .B(B[86]), .Z(n3752) );
  NAND U3284 ( .A(n3753), .B(n3754), .Z(n3751) );
  NANDN U3285 ( .A(B[86]), .B(A[86]), .Z(n3754) );
  AND U3286 ( .A(n3755), .B(n3756), .Z(n3753) );
  NAND U3287 ( .A(n3757), .B(n3758), .Z(n3756) );
  NANDN U3288 ( .A(A[85]), .B(B[85]), .Z(n3758) );
  AND U3289 ( .A(n3759), .B(n3760), .Z(n3757) );
  NANDN U3290 ( .A(A[84]), .B(B[84]), .Z(n3760) );
  NAND U3291 ( .A(n3761), .B(n3762), .Z(n3759) );
  NANDN U3292 ( .A(B[84]), .B(A[84]), .Z(n3762) );
  AND U3293 ( .A(n3763), .B(n3764), .Z(n3761) );
  NAND U3294 ( .A(n3765), .B(n3766), .Z(n3764) );
  NANDN U3295 ( .A(A[83]), .B(B[83]), .Z(n3766) );
  AND U3296 ( .A(n3767), .B(n3768), .Z(n3765) );
  NANDN U3297 ( .A(A[82]), .B(B[82]), .Z(n3768) );
  NAND U3298 ( .A(n3769), .B(n3770), .Z(n3767) );
  NANDN U3299 ( .A(B[82]), .B(A[82]), .Z(n3770) );
  AND U3300 ( .A(n3771), .B(n3772), .Z(n3769) );
  NAND U3301 ( .A(n3773), .B(n3774), .Z(n3772) );
  NANDN U3302 ( .A(A[81]), .B(B[81]), .Z(n3774) );
  AND U3303 ( .A(n3775), .B(n3776), .Z(n3773) );
  NANDN U3304 ( .A(A[80]), .B(B[80]), .Z(n3776) );
  NAND U3305 ( .A(n3777), .B(n3778), .Z(n3775) );
  NANDN U3306 ( .A(B[80]), .B(A[80]), .Z(n3778) );
  AND U3307 ( .A(n3779), .B(n3780), .Z(n3777) );
  NAND U3308 ( .A(n3781), .B(n3782), .Z(n3780) );
  NANDN U3309 ( .A(A[79]), .B(B[79]), .Z(n3782) );
  AND U3310 ( .A(n3783), .B(n3784), .Z(n3781) );
  NANDN U3311 ( .A(A[78]), .B(B[78]), .Z(n3784) );
  NAND U3312 ( .A(n3785), .B(n3786), .Z(n3783) );
  NANDN U3313 ( .A(B[78]), .B(A[78]), .Z(n3786) );
  AND U3314 ( .A(n3787), .B(n3788), .Z(n3785) );
  NAND U3315 ( .A(n3789), .B(n3790), .Z(n3788) );
  NANDN U3316 ( .A(A[77]), .B(B[77]), .Z(n3790) );
  AND U3317 ( .A(n3791), .B(n3792), .Z(n3789) );
  NANDN U3318 ( .A(A[76]), .B(B[76]), .Z(n3792) );
  NAND U3319 ( .A(n3793), .B(n3794), .Z(n3791) );
  NANDN U3320 ( .A(B[76]), .B(A[76]), .Z(n3794) );
  AND U3321 ( .A(n3795), .B(n3796), .Z(n3793) );
  NAND U3322 ( .A(n3797), .B(n3798), .Z(n3796) );
  NANDN U3323 ( .A(A[75]), .B(B[75]), .Z(n3798) );
  AND U3324 ( .A(n3799), .B(n3800), .Z(n3797) );
  NANDN U3325 ( .A(A[74]), .B(B[74]), .Z(n3800) );
  NAND U3326 ( .A(n3801), .B(n3802), .Z(n3799) );
  NANDN U3327 ( .A(B[74]), .B(A[74]), .Z(n3802) );
  AND U3328 ( .A(n3803), .B(n3804), .Z(n3801) );
  NAND U3329 ( .A(n3805), .B(n3806), .Z(n3804) );
  NANDN U3330 ( .A(A[73]), .B(B[73]), .Z(n3806) );
  AND U3331 ( .A(n3807), .B(n3808), .Z(n3805) );
  NANDN U3332 ( .A(A[72]), .B(B[72]), .Z(n3808) );
  NAND U3333 ( .A(n3809), .B(n3810), .Z(n3807) );
  NANDN U3334 ( .A(B[72]), .B(A[72]), .Z(n3810) );
  AND U3335 ( .A(n3811), .B(n3812), .Z(n3809) );
  NAND U3336 ( .A(n3813), .B(n3814), .Z(n3812) );
  NANDN U3337 ( .A(A[71]), .B(B[71]), .Z(n3814) );
  AND U3338 ( .A(n3815), .B(n3816), .Z(n3813) );
  NANDN U3339 ( .A(A[70]), .B(B[70]), .Z(n3816) );
  NAND U3340 ( .A(n3817), .B(n3818), .Z(n3815) );
  NANDN U3341 ( .A(B[70]), .B(A[70]), .Z(n3818) );
  AND U3342 ( .A(n3819), .B(n3820), .Z(n3817) );
  NAND U3343 ( .A(n3821), .B(n3822), .Z(n3820) );
  NANDN U3344 ( .A(A[69]), .B(B[69]), .Z(n3822) );
  AND U3345 ( .A(n3823), .B(n3824), .Z(n3821) );
  NANDN U3346 ( .A(A[68]), .B(B[68]), .Z(n3824) );
  NAND U3347 ( .A(n3825), .B(n3826), .Z(n3823) );
  NANDN U3348 ( .A(B[68]), .B(A[68]), .Z(n3826) );
  AND U3349 ( .A(n3827), .B(n3828), .Z(n3825) );
  NAND U3350 ( .A(n3829), .B(n3830), .Z(n3828) );
  NANDN U3351 ( .A(A[67]), .B(B[67]), .Z(n3830) );
  AND U3352 ( .A(n3831), .B(n3832), .Z(n3829) );
  NANDN U3353 ( .A(A[66]), .B(B[66]), .Z(n3832) );
  NAND U3354 ( .A(n3833), .B(n3834), .Z(n3831) );
  NANDN U3355 ( .A(B[66]), .B(A[66]), .Z(n3834) );
  AND U3356 ( .A(n3835), .B(n3836), .Z(n3833) );
  NAND U3357 ( .A(n3837), .B(n3838), .Z(n3836) );
  NANDN U3358 ( .A(A[65]), .B(B[65]), .Z(n3838) );
  AND U3359 ( .A(n3839), .B(n3840), .Z(n3837) );
  NANDN U3360 ( .A(A[64]), .B(B[64]), .Z(n3840) );
  NAND U3361 ( .A(n3841), .B(n3842), .Z(n3839) );
  NANDN U3362 ( .A(B[64]), .B(A[64]), .Z(n3842) );
  AND U3363 ( .A(n3843), .B(n3844), .Z(n3841) );
  NAND U3364 ( .A(n3845), .B(n3846), .Z(n3844) );
  NANDN U3365 ( .A(A[63]), .B(B[63]), .Z(n3846) );
  AND U3366 ( .A(n3847), .B(n3848), .Z(n3845) );
  NANDN U3367 ( .A(A[62]), .B(B[62]), .Z(n3848) );
  NAND U3368 ( .A(n3849), .B(n3850), .Z(n3847) );
  NANDN U3369 ( .A(B[62]), .B(A[62]), .Z(n3850) );
  AND U3370 ( .A(n3851), .B(n3852), .Z(n3849) );
  NAND U3371 ( .A(n3853), .B(n3854), .Z(n3852) );
  NANDN U3372 ( .A(A[61]), .B(B[61]), .Z(n3854) );
  AND U3373 ( .A(n3855), .B(n3856), .Z(n3853) );
  NANDN U3374 ( .A(A[60]), .B(B[60]), .Z(n3856) );
  NAND U3375 ( .A(n3857), .B(n3858), .Z(n3855) );
  NANDN U3376 ( .A(B[60]), .B(A[60]), .Z(n3858) );
  AND U3377 ( .A(n3859), .B(n3860), .Z(n3857) );
  NAND U3378 ( .A(n3861), .B(n3862), .Z(n3860) );
  NANDN U3379 ( .A(A[59]), .B(B[59]), .Z(n3862) );
  AND U3380 ( .A(n3863), .B(n3864), .Z(n3861) );
  NANDN U3381 ( .A(A[58]), .B(B[58]), .Z(n3864) );
  NAND U3382 ( .A(n3865), .B(n3866), .Z(n3863) );
  NANDN U3383 ( .A(B[58]), .B(A[58]), .Z(n3866) );
  AND U3384 ( .A(n3867), .B(n3868), .Z(n3865) );
  NAND U3385 ( .A(n3869), .B(n3870), .Z(n3868) );
  NANDN U3386 ( .A(A[57]), .B(B[57]), .Z(n3870) );
  AND U3387 ( .A(n3871), .B(n3872), .Z(n3869) );
  NANDN U3388 ( .A(A[56]), .B(B[56]), .Z(n3872) );
  NAND U3389 ( .A(n3873), .B(n3874), .Z(n3871) );
  NANDN U3390 ( .A(B[56]), .B(A[56]), .Z(n3874) );
  AND U3391 ( .A(n3875), .B(n3876), .Z(n3873) );
  NAND U3392 ( .A(n3877), .B(n3878), .Z(n3876) );
  NANDN U3393 ( .A(A[55]), .B(B[55]), .Z(n3878) );
  AND U3394 ( .A(n3879), .B(n3880), .Z(n3877) );
  NANDN U3395 ( .A(A[54]), .B(B[54]), .Z(n3880) );
  NAND U3396 ( .A(n3881), .B(n3882), .Z(n3879) );
  NANDN U3397 ( .A(B[54]), .B(A[54]), .Z(n3882) );
  AND U3398 ( .A(n3883), .B(n3884), .Z(n3881) );
  NAND U3399 ( .A(n3885), .B(n3886), .Z(n3884) );
  NANDN U3400 ( .A(A[53]), .B(B[53]), .Z(n3886) );
  AND U3401 ( .A(n3887), .B(n3888), .Z(n3885) );
  NANDN U3402 ( .A(A[52]), .B(B[52]), .Z(n3888) );
  NAND U3403 ( .A(n3889), .B(n3890), .Z(n3887) );
  NANDN U3404 ( .A(B[52]), .B(A[52]), .Z(n3890) );
  AND U3405 ( .A(n3891), .B(n3892), .Z(n3889) );
  NAND U3406 ( .A(n3893), .B(n3894), .Z(n3892) );
  NANDN U3407 ( .A(A[51]), .B(B[51]), .Z(n3894) );
  AND U3408 ( .A(n3895), .B(n3896), .Z(n3893) );
  NANDN U3409 ( .A(A[50]), .B(B[50]), .Z(n3896) );
  NAND U3410 ( .A(n3897), .B(n3898), .Z(n3895) );
  NANDN U3411 ( .A(B[50]), .B(A[50]), .Z(n3898) );
  AND U3412 ( .A(n3899), .B(n3900), .Z(n3897) );
  NAND U3413 ( .A(n3901), .B(n3902), .Z(n3900) );
  NANDN U3414 ( .A(A[49]), .B(B[49]), .Z(n3902) );
  AND U3415 ( .A(n3903), .B(n3904), .Z(n3901) );
  NANDN U3416 ( .A(A[48]), .B(B[48]), .Z(n3904) );
  NAND U3417 ( .A(n3905), .B(n3906), .Z(n3903) );
  NANDN U3418 ( .A(B[48]), .B(A[48]), .Z(n3906) );
  AND U3419 ( .A(n3907), .B(n3908), .Z(n3905) );
  NAND U3420 ( .A(n3909), .B(n3910), .Z(n3908) );
  NANDN U3421 ( .A(A[47]), .B(B[47]), .Z(n3910) );
  AND U3422 ( .A(n3911), .B(n3912), .Z(n3909) );
  NANDN U3423 ( .A(A[46]), .B(B[46]), .Z(n3912) );
  NAND U3424 ( .A(n3913), .B(n3914), .Z(n3911) );
  NANDN U3425 ( .A(B[46]), .B(A[46]), .Z(n3914) );
  AND U3426 ( .A(n3915), .B(n3916), .Z(n3913) );
  NAND U3427 ( .A(n3917), .B(n3918), .Z(n3916) );
  NANDN U3428 ( .A(A[45]), .B(B[45]), .Z(n3918) );
  AND U3429 ( .A(n3919), .B(n3920), .Z(n3917) );
  NANDN U3430 ( .A(A[44]), .B(B[44]), .Z(n3920) );
  NAND U3431 ( .A(n3921), .B(n3922), .Z(n3919) );
  NANDN U3432 ( .A(B[44]), .B(A[44]), .Z(n3922) );
  AND U3433 ( .A(n3923), .B(n3924), .Z(n3921) );
  NAND U3434 ( .A(n3925), .B(n3926), .Z(n3924) );
  NANDN U3435 ( .A(A[43]), .B(B[43]), .Z(n3926) );
  AND U3436 ( .A(n3927), .B(n3928), .Z(n3925) );
  NANDN U3437 ( .A(A[42]), .B(B[42]), .Z(n3928) );
  NAND U3438 ( .A(n3929), .B(n3930), .Z(n3927) );
  NANDN U3439 ( .A(B[42]), .B(A[42]), .Z(n3930) );
  AND U3440 ( .A(n3931), .B(n3932), .Z(n3929) );
  NAND U3441 ( .A(n3933), .B(n3934), .Z(n3932) );
  NANDN U3442 ( .A(A[41]), .B(B[41]), .Z(n3934) );
  AND U3443 ( .A(n3935), .B(n3936), .Z(n3933) );
  NANDN U3444 ( .A(A[40]), .B(B[40]), .Z(n3936) );
  NAND U3445 ( .A(n3937), .B(n3938), .Z(n3935) );
  NANDN U3446 ( .A(B[40]), .B(A[40]), .Z(n3938) );
  AND U3447 ( .A(n3939), .B(n3940), .Z(n3937) );
  NAND U3448 ( .A(n3941), .B(n3942), .Z(n3940) );
  NANDN U3449 ( .A(A[39]), .B(B[39]), .Z(n3942) );
  AND U3450 ( .A(n3943), .B(n3944), .Z(n3941) );
  NANDN U3451 ( .A(A[38]), .B(B[38]), .Z(n3944) );
  NAND U3452 ( .A(n3945), .B(n3946), .Z(n3943) );
  NANDN U3453 ( .A(B[38]), .B(A[38]), .Z(n3946) );
  AND U3454 ( .A(n3947), .B(n3948), .Z(n3945) );
  NAND U3455 ( .A(n3949), .B(n3950), .Z(n3948) );
  NANDN U3456 ( .A(A[37]), .B(B[37]), .Z(n3950) );
  AND U3457 ( .A(n3951), .B(n3952), .Z(n3949) );
  NANDN U3458 ( .A(A[36]), .B(B[36]), .Z(n3952) );
  NAND U3459 ( .A(n3953), .B(n3954), .Z(n3951) );
  NANDN U3460 ( .A(B[36]), .B(A[36]), .Z(n3954) );
  AND U3461 ( .A(n3955), .B(n3956), .Z(n3953) );
  NAND U3462 ( .A(n3957), .B(n3958), .Z(n3956) );
  NANDN U3463 ( .A(A[35]), .B(B[35]), .Z(n3958) );
  AND U3464 ( .A(n3959), .B(n3960), .Z(n3957) );
  NANDN U3465 ( .A(A[34]), .B(B[34]), .Z(n3960) );
  NAND U3466 ( .A(n3961), .B(n3962), .Z(n3959) );
  NANDN U3467 ( .A(B[34]), .B(A[34]), .Z(n3962) );
  AND U3468 ( .A(n3963), .B(n3964), .Z(n3961) );
  NAND U3469 ( .A(n3965), .B(n3966), .Z(n3964) );
  NANDN U3470 ( .A(A[33]), .B(B[33]), .Z(n3966) );
  AND U3471 ( .A(n3967), .B(n3968), .Z(n3965) );
  NANDN U3472 ( .A(A[32]), .B(B[32]), .Z(n3968) );
  NAND U3473 ( .A(n3969), .B(n3970), .Z(n3967) );
  NANDN U3474 ( .A(B[32]), .B(A[32]), .Z(n3970) );
  AND U3475 ( .A(n3971), .B(n3972), .Z(n3969) );
  NAND U3476 ( .A(n3973), .B(n3974), .Z(n3972) );
  NANDN U3477 ( .A(A[31]), .B(B[31]), .Z(n3974) );
  AND U3478 ( .A(n3975), .B(n3976), .Z(n3973) );
  NANDN U3479 ( .A(A[30]), .B(B[30]), .Z(n3976) );
  NAND U3480 ( .A(n3977), .B(n3978), .Z(n3975) );
  NANDN U3481 ( .A(B[30]), .B(A[30]), .Z(n3978) );
  AND U3482 ( .A(n3979), .B(n3980), .Z(n3977) );
  NAND U3483 ( .A(n3981), .B(n3982), .Z(n3980) );
  NANDN U3484 ( .A(A[29]), .B(B[29]), .Z(n3982) );
  AND U3485 ( .A(n3983), .B(n3984), .Z(n3981) );
  NANDN U3486 ( .A(A[28]), .B(B[28]), .Z(n3984) );
  NAND U3487 ( .A(n3985), .B(n3986), .Z(n3983) );
  NANDN U3488 ( .A(B[28]), .B(A[28]), .Z(n3986) );
  AND U3489 ( .A(n3987), .B(n3988), .Z(n3985) );
  NAND U3490 ( .A(n3989), .B(n3990), .Z(n3988) );
  NANDN U3491 ( .A(A[27]), .B(B[27]), .Z(n3990) );
  AND U3492 ( .A(n3991), .B(n3992), .Z(n3989) );
  NANDN U3493 ( .A(A[26]), .B(B[26]), .Z(n3992) );
  NAND U3494 ( .A(n3993), .B(n3994), .Z(n3991) );
  NANDN U3495 ( .A(B[26]), .B(A[26]), .Z(n3994) );
  AND U3496 ( .A(n3995), .B(n3996), .Z(n3993) );
  NAND U3497 ( .A(n3997), .B(n3998), .Z(n3996) );
  NANDN U3498 ( .A(A[25]), .B(B[25]), .Z(n3998) );
  AND U3499 ( .A(n3999), .B(n4000), .Z(n3997) );
  NANDN U3500 ( .A(A[24]), .B(B[24]), .Z(n4000) );
  NAND U3501 ( .A(n4001), .B(n4002), .Z(n3999) );
  NANDN U3502 ( .A(B[24]), .B(A[24]), .Z(n4002) );
  AND U3503 ( .A(n4003), .B(n4004), .Z(n4001) );
  NAND U3504 ( .A(n4005), .B(n4006), .Z(n4004) );
  NANDN U3505 ( .A(A[23]), .B(B[23]), .Z(n4006) );
  AND U3506 ( .A(n4007), .B(n4008), .Z(n4005) );
  NANDN U3507 ( .A(A[22]), .B(B[22]), .Z(n4008) );
  NAND U3508 ( .A(n4009), .B(n4010), .Z(n4007) );
  NANDN U3509 ( .A(B[22]), .B(A[22]), .Z(n4010) );
  AND U3510 ( .A(n4011), .B(n4012), .Z(n4009) );
  NAND U3511 ( .A(n4013), .B(n4014), .Z(n4012) );
  NANDN U3512 ( .A(A[21]), .B(B[21]), .Z(n4014) );
  AND U3513 ( .A(n4015), .B(n4016), .Z(n4013) );
  NANDN U3514 ( .A(A[20]), .B(B[20]), .Z(n4016) );
  NAND U3515 ( .A(n4017), .B(n4018), .Z(n4015) );
  NANDN U3516 ( .A(B[20]), .B(A[20]), .Z(n4018) );
  AND U3517 ( .A(n4019), .B(n4020), .Z(n4017) );
  NAND U3518 ( .A(n4021), .B(n4022), .Z(n4020) );
  NANDN U3519 ( .A(A[19]), .B(B[19]), .Z(n4022) );
  AND U3520 ( .A(n4023), .B(n4024), .Z(n4021) );
  NANDN U3521 ( .A(A[18]), .B(B[18]), .Z(n4024) );
  NAND U3522 ( .A(n4025), .B(n4026), .Z(n4023) );
  NANDN U3523 ( .A(B[18]), .B(A[18]), .Z(n4026) );
  AND U3524 ( .A(n4027), .B(n4028), .Z(n4025) );
  NAND U3525 ( .A(n4029), .B(n4030), .Z(n4028) );
  NANDN U3526 ( .A(A[17]), .B(B[17]), .Z(n4030) );
  AND U3527 ( .A(n4031), .B(n4032), .Z(n4029) );
  NANDN U3528 ( .A(A[16]), .B(B[16]), .Z(n4032) );
  NAND U3529 ( .A(n4033), .B(n4034), .Z(n4031) );
  NANDN U3530 ( .A(B[16]), .B(A[16]), .Z(n4034) );
  AND U3531 ( .A(n4035), .B(n4036), .Z(n4033) );
  NAND U3532 ( .A(n4037), .B(n4038), .Z(n4036) );
  NANDN U3533 ( .A(A[15]), .B(B[15]), .Z(n4038) );
  AND U3534 ( .A(n4039), .B(n4040), .Z(n4037) );
  NANDN U3535 ( .A(A[14]), .B(B[14]), .Z(n4040) );
  NAND U3536 ( .A(n4041), .B(n4042), .Z(n4039) );
  NANDN U3537 ( .A(B[14]), .B(A[14]), .Z(n4042) );
  AND U3538 ( .A(n4043), .B(n4044), .Z(n4041) );
  NAND U3539 ( .A(n4045), .B(n4046), .Z(n4044) );
  NANDN U3540 ( .A(A[13]), .B(B[13]), .Z(n4046) );
  AND U3541 ( .A(n4047), .B(n4048), .Z(n4045) );
  NANDN U3542 ( .A(A[12]), .B(B[12]), .Z(n4048) );
  NAND U3543 ( .A(n4049), .B(n4050), .Z(n4047) );
  NANDN U3544 ( .A(B[12]), .B(A[12]), .Z(n4050) );
  AND U3545 ( .A(n4051), .B(n4052), .Z(n4049) );
  NAND U3546 ( .A(n4053), .B(n4054), .Z(n4052) );
  NANDN U3547 ( .A(A[11]), .B(B[11]), .Z(n4054) );
  AND U3548 ( .A(n4055), .B(n4056), .Z(n4053) );
  NANDN U3549 ( .A(A[10]), .B(B[10]), .Z(n4056) );
  NAND U3550 ( .A(n4057), .B(n4058), .Z(n4055) );
  NANDN U3551 ( .A(B[9]), .B(A[9]), .Z(n4058) );
  AND U3552 ( .A(n4059), .B(n4060), .Z(n4057) );
  NAND U3553 ( .A(n4061), .B(n4062), .Z(n4060) );
  NANDN U3554 ( .A(A[9]), .B(B[9]), .Z(n4062) );
  AND U3555 ( .A(n4063), .B(n4064), .Z(n4061) );
  NANDN U3556 ( .A(A[8]), .B(B[8]), .Z(n4064) );
  NAND U3557 ( .A(n4065), .B(n4066), .Z(n4063) );
  NANDN U3558 ( .A(B[8]), .B(A[8]), .Z(n4066) );
  AND U3559 ( .A(n4067), .B(n4068), .Z(n4065) );
  NAND U3560 ( .A(n4069), .B(n4070), .Z(n4068) );
  NANDN U3561 ( .A(A[7]), .B(B[7]), .Z(n4070) );
  AND U3562 ( .A(n4071), .B(n4072), .Z(n4069) );
  NANDN U3563 ( .A(A[6]), .B(B[6]), .Z(n4072) );
  NAND U3564 ( .A(n4073), .B(n4074), .Z(n4071) );
  NANDN U3565 ( .A(B[6]), .B(A[6]), .Z(n4074) );
  AND U3566 ( .A(n4075), .B(n4076), .Z(n4073) );
  NAND U3567 ( .A(n4077), .B(n4078), .Z(n4076) );
  NANDN U3568 ( .A(A[5]), .B(B[5]), .Z(n4078) );
  AND U3569 ( .A(n4079), .B(n4080), .Z(n4077) );
  NANDN U3570 ( .A(A[4]), .B(B[4]), .Z(n4080) );
  NAND U3571 ( .A(n4081), .B(n4082), .Z(n4079) );
  NANDN U3572 ( .A(B[4]), .B(A[4]), .Z(n4082) );
  AND U3573 ( .A(n4083), .B(n4084), .Z(n4081) );
  NAND U3574 ( .A(n4085), .B(n4086), .Z(n4084) );
  NANDN U3575 ( .A(A[3]), .B(B[3]), .Z(n4086) );
  AND U3576 ( .A(n4087), .B(n4088), .Z(n4085) );
  NANDN U3577 ( .A(A[2]), .B(B[2]), .Z(n4088) );
  NAND U3578 ( .A(n4089), .B(n4090), .Z(n4087) );
  NANDN U3579 ( .A(B[2]), .B(A[2]), .Z(n4090) );
  AND U3580 ( .A(n4091), .B(n4092), .Z(n4089) );
  NAND U3581 ( .A(n4093), .B(A[0]), .Z(n4092) );
  ANDN U3582 ( .B(n4094), .A(B[0]), .Z(n4093) );
  NANDN U3583 ( .A(A[1]), .B(B[1]), .Z(n4094) );
  NANDN U3584 ( .A(B[1]), .B(A[1]), .Z(n4091) );
  NANDN U3585 ( .A(B[3]), .B(A[3]), .Z(n4083) );
  NANDN U3586 ( .A(B[5]), .B(A[5]), .Z(n4075) );
  NANDN U3587 ( .A(B[7]), .B(A[7]), .Z(n4067) );
  NANDN U3588 ( .A(B[10]), .B(A[10]), .Z(n4059) );
  NANDN U3589 ( .A(B[11]), .B(A[11]), .Z(n4051) );
  NANDN U3590 ( .A(B[13]), .B(A[13]), .Z(n4043) );
  NANDN U3591 ( .A(B[15]), .B(A[15]), .Z(n4035) );
  NANDN U3592 ( .A(B[17]), .B(A[17]), .Z(n4027) );
  NANDN U3593 ( .A(B[19]), .B(A[19]), .Z(n4019) );
  NANDN U3594 ( .A(B[21]), .B(A[21]), .Z(n4011) );
  NANDN U3595 ( .A(B[23]), .B(A[23]), .Z(n4003) );
  NANDN U3596 ( .A(B[25]), .B(A[25]), .Z(n3995) );
  NANDN U3597 ( .A(B[27]), .B(A[27]), .Z(n3987) );
  NANDN U3598 ( .A(B[29]), .B(A[29]), .Z(n3979) );
  NANDN U3599 ( .A(B[31]), .B(A[31]), .Z(n3971) );
  NANDN U3600 ( .A(B[33]), .B(A[33]), .Z(n3963) );
  NANDN U3601 ( .A(B[35]), .B(A[35]), .Z(n3955) );
  NANDN U3602 ( .A(B[37]), .B(A[37]), .Z(n3947) );
  NANDN U3603 ( .A(B[39]), .B(A[39]), .Z(n3939) );
  NANDN U3604 ( .A(B[41]), .B(A[41]), .Z(n3931) );
  NANDN U3605 ( .A(B[43]), .B(A[43]), .Z(n3923) );
  NANDN U3606 ( .A(B[45]), .B(A[45]), .Z(n3915) );
  NANDN U3607 ( .A(B[47]), .B(A[47]), .Z(n3907) );
  NANDN U3608 ( .A(B[49]), .B(A[49]), .Z(n3899) );
  NANDN U3609 ( .A(B[51]), .B(A[51]), .Z(n3891) );
  NANDN U3610 ( .A(B[53]), .B(A[53]), .Z(n3883) );
  NANDN U3611 ( .A(B[55]), .B(A[55]), .Z(n3875) );
  NANDN U3612 ( .A(B[57]), .B(A[57]), .Z(n3867) );
  NANDN U3613 ( .A(B[59]), .B(A[59]), .Z(n3859) );
  NANDN U3614 ( .A(B[61]), .B(A[61]), .Z(n3851) );
  NANDN U3615 ( .A(B[63]), .B(A[63]), .Z(n3843) );
  NANDN U3616 ( .A(B[65]), .B(A[65]), .Z(n3835) );
  NANDN U3617 ( .A(B[67]), .B(A[67]), .Z(n3827) );
  NANDN U3618 ( .A(B[69]), .B(A[69]), .Z(n3819) );
  NANDN U3619 ( .A(B[71]), .B(A[71]), .Z(n3811) );
  NANDN U3620 ( .A(B[73]), .B(A[73]), .Z(n3803) );
  NANDN U3621 ( .A(B[75]), .B(A[75]), .Z(n3795) );
  NANDN U3622 ( .A(B[77]), .B(A[77]), .Z(n3787) );
  NANDN U3623 ( .A(B[79]), .B(A[79]), .Z(n3779) );
  NANDN U3624 ( .A(B[81]), .B(A[81]), .Z(n3771) );
  NANDN U3625 ( .A(B[83]), .B(A[83]), .Z(n3763) );
  NANDN U3626 ( .A(B[85]), .B(A[85]), .Z(n3755) );
  NANDN U3627 ( .A(B[87]), .B(A[87]), .Z(n3747) );
  NANDN U3628 ( .A(B[89]), .B(A[89]), .Z(n3739) );
  NANDN U3629 ( .A(B[91]), .B(A[91]), .Z(n3731) );
  NANDN U3630 ( .A(B[93]), .B(A[93]), .Z(n3723) );
  NANDN U3631 ( .A(B[95]), .B(A[95]), .Z(n3715) );
  NANDN U3632 ( .A(B[97]), .B(A[97]), .Z(n3707) );
  NANDN U3633 ( .A(B[100]), .B(A[100]), .Z(n3699) );
  NANDN U3634 ( .A(B[101]), .B(A[101]), .Z(n3691) );
  NANDN U3635 ( .A(B[103]), .B(A[103]), .Z(n3683) );
  NANDN U3636 ( .A(B[105]), .B(A[105]), .Z(n3675) );
  NANDN U3637 ( .A(B[107]), .B(A[107]), .Z(n3667) );
  NANDN U3638 ( .A(B[109]), .B(A[109]), .Z(n3659) );
  NANDN U3639 ( .A(B[111]), .B(A[111]), .Z(n3651) );
  NANDN U3640 ( .A(B[113]), .B(A[113]), .Z(n3643) );
  NANDN U3641 ( .A(B[115]), .B(A[115]), .Z(n3635) );
  NANDN U3642 ( .A(B[117]), .B(A[117]), .Z(n3627) );
  NANDN U3643 ( .A(B[119]), .B(A[119]), .Z(n3619) );
  NANDN U3644 ( .A(B[121]), .B(A[121]), .Z(n3611) );
  NANDN U3645 ( .A(B[123]), .B(A[123]), .Z(n3603) );
  NANDN U3646 ( .A(B[125]), .B(A[125]), .Z(n3595) );
  NANDN U3647 ( .A(B[127]), .B(A[127]), .Z(n3587) );
  NANDN U3648 ( .A(B[129]), .B(A[129]), .Z(n3579) );
  NANDN U3649 ( .A(B[131]), .B(A[131]), .Z(n3571) );
  NANDN U3650 ( .A(B[133]), .B(A[133]), .Z(n3563) );
  NANDN U3651 ( .A(B[135]), .B(A[135]), .Z(n3555) );
  NANDN U3652 ( .A(B[137]), .B(A[137]), .Z(n3547) );
  NANDN U3653 ( .A(B[139]), .B(A[139]), .Z(n3539) );
  NANDN U3654 ( .A(B[141]), .B(A[141]), .Z(n3531) );
  NANDN U3655 ( .A(B[143]), .B(A[143]), .Z(n3523) );
  NANDN U3656 ( .A(B[145]), .B(A[145]), .Z(n3515) );
  NANDN U3657 ( .A(B[147]), .B(A[147]), .Z(n3507) );
  NANDN U3658 ( .A(B[149]), .B(A[149]), .Z(n3499) );
  NANDN U3659 ( .A(B[151]), .B(A[151]), .Z(n3491) );
  NANDN U3660 ( .A(B[153]), .B(A[153]), .Z(n3483) );
  NANDN U3661 ( .A(B[155]), .B(A[155]), .Z(n3475) );
  NANDN U3662 ( .A(B[157]), .B(A[157]), .Z(n3467) );
  NANDN U3663 ( .A(B[159]), .B(A[159]), .Z(n3459) );
  NANDN U3664 ( .A(B[161]), .B(A[161]), .Z(n3451) );
  NANDN U3665 ( .A(B[163]), .B(A[163]), .Z(n3443) );
  NANDN U3666 ( .A(B[165]), .B(A[165]), .Z(n3435) );
  NANDN U3667 ( .A(B[167]), .B(A[167]), .Z(n3427) );
  NANDN U3668 ( .A(B[169]), .B(A[169]), .Z(n3419) );
  NANDN U3669 ( .A(B[171]), .B(A[171]), .Z(n3411) );
  NANDN U3670 ( .A(B[173]), .B(A[173]), .Z(n3403) );
  NANDN U3671 ( .A(B[175]), .B(A[175]), .Z(n3395) );
  NANDN U3672 ( .A(B[177]), .B(A[177]), .Z(n3387) );
  NANDN U3673 ( .A(B[179]), .B(A[179]), .Z(n3379) );
  NANDN U3674 ( .A(B[181]), .B(A[181]), .Z(n3371) );
  NANDN U3675 ( .A(B[183]), .B(A[183]), .Z(n3363) );
  NANDN U3676 ( .A(B[185]), .B(A[185]), .Z(n3355) );
  NANDN U3677 ( .A(B[187]), .B(A[187]), .Z(n3347) );
  NANDN U3678 ( .A(B[189]), .B(A[189]), .Z(n3339) );
  NANDN U3679 ( .A(B[191]), .B(A[191]), .Z(n3331) );
  NANDN U3680 ( .A(B[193]), .B(A[193]), .Z(n3323) );
  NANDN U3681 ( .A(B[195]), .B(A[195]), .Z(n3315) );
  NANDN U3682 ( .A(B[197]), .B(A[197]), .Z(n3307) );
  NANDN U3683 ( .A(B[199]), .B(A[199]), .Z(n3299) );
  NANDN U3684 ( .A(B[201]), .B(A[201]), .Z(n3291) );
  NANDN U3685 ( .A(B[203]), .B(A[203]), .Z(n3283) );
  NANDN U3686 ( .A(B[205]), .B(A[205]), .Z(n3275) );
  NANDN U3687 ( .A(B[207]), .B(A[207]), .Z(n3267) );
  NANDN U3688 ( .A(B[209]), .B(A[209]), .Z(n3259) );
  NANDN U3689 ( .A(B[211]), .B(A[211]), .Z(n3251) );
  NANDN U3690 ( .A(B[213]), .B(A[213]), .Z(n3243) );
  NANDN U3691 ( .A(B[215]), .B(A[215]), .Z(n3235) );
  NANDN U3692 ( .A(B[217]), .B(A[217]), .Z(n3227) );
  NANDN U3693 ( .A(B[219]), .B(A[219]), .Z(n3219) );
  NANDN U3694 ( .A(B[221]), .B(A[221]), .Z(n3211) );
  NANDN U3695 ( .A(B[223]), .B(A[223]), .Z(n3203) );
  NANDN U3696 ( .A(B[225]), .B(A[225]), .Z(n3195) );
  NANDN U3697 ( .A(B[227]), .B(A[227]), .Z(n3187) );
  NANDN U3698 ( .A(B[229]), .B(A[229]), .Z(n3179) );
  NANDN U3699 ( .A(B[231]), .B(A[231]), .Z(n3171) );
  NANDN U3700 ( .A(B[233]), .B(A[233]), .Z(n3163) );
  NANDN U3701 ( .A(B[235]), .B(A[235]), .Z(n3155) );
  NANDN U3702 ( .A(B[237]), .B(A[237]), .Z(n3147) );
  NANDN U3703 ( .A(B[239]), .B(A[239]), .Z(n3139) );
  NANDN U3704 ( .A(B[241]), .B(A[241]), .Z(n3131) );
  NANDN U3705 ( .A(B[243]), .B(A[243]), .Z(n3123) );
  NANDN U3706 ( .A(B[245]), .B(A[245]), .Z(n3115) );
  NANDN U3707 ( .A(B[247]), .B(A[247]), .Z(n3107) );
  NANDN U3708 ( .A(B[249]), .B(A[249]), .Z(n3099) );
  NANDN U3709 ( .A(B[251]), .B(A[251]), .Z(n3091) );
  NANDN U3710 ( .A(B[253]), .B(A[253]), .Z(n3083) );
  NANDN U3711 ( .A(B[255]), .B(A[255]), .Z(n3075) );
  NANDN U3712 ( .A(B[257]), .B(A[257]), .Z(n3067) );
  NANDN U3713 ( .A(B[259]), .B(A[259]), .Z(n3059) );
  NANDN U3714 ( .A(B[261]), .B(A[261]), .Z(n3051) );
  NANDN U3715 ( .A(B[263]), .B(A[263]), .Z(n3043) );
  NANDN U3716 ( .A(B[265]), .B(A[265]), .Z(n3035) );
  NANDN U3717 ( .A(B[267]), .B(A[267]), .Z(n3027) );
  NANDN U3718 ( .A(B[269]), .B(A[269]), .Z(n3019) );
  NANDN U3719 ( .A(B[271]), .B(A[271]), .Z(n3011) );
  NANDN U3720 ( .A(B[273]), .B(A[273]), .Z(n3003) );
  NANDN U3721 ( .A(B[275]), .B(A[275]), .Z(n2995) );
  NANDN U3722 ( .A(B[277]), .B(A[277]), .Z(n2987) );
  NANDN U3723 ( .A(B[279]), .B(A[279]), .Z(n2979) );
  NANDN U3724 ( .A(B[281]), .B(A[281]), .Z(n2971) );
  NANDN U3725 ( .A(B[283]), .B(A[283]), .Z(n2963) );
  NANDN U3726 ( .A(B[285]), .B(A[285]), .Z(n2955) );
  NANDN U3727 ( .A(B[287]), .B(A[287]), .Z(n2947) );
  NANDN U3728 ( .A(B[289]), .B(A[289]), .Z(n2939) );
  NANDN U3729 ( .A(B[291]), .B(A[291]), .Z(n2931) );
  NANDN U3730 ( .A(B[293]), .B(A[293]), .Z(n2923) );
  NANDN U3731 ( .A(B[295]), .B(A[295]), .Z(n2915) );
  NANDN U3732 ( .A(B[297]), .B(A[297]), .Z(n2907) );
  NANDN U3733 ( .A(B[299]), .B(A[299]), .Z(n2899) );
  NANDN U3734 ( .A(B[301]), .B(A[301]), .Z(n2891) );
  NANDN U3735 ( .A(B[303]), .B(A[303]), .Z(n2883) );
  NANDN U3736 ( .A(B[305]), .B(A[305]), .Z(n2875) );
  NANDN U3737 ( .A(B[307]), .B(A[307]), .Z(n2867) );
  NANDN U3738 ( .A(B[309]), .B(A[309]), .Z(n2859) );
  NANDN U3739 ( .A(B[311]), .B(A[311]), .Z(n2851) );
  NANDN U3740 ( .A(B[313]), .B(A[313]), .Z(n2843) );
  NANDN U3741 ( .A(B[315]), .B(A[315]), .Z(n2835) );
  NANDN U3742 ( .A(B[317]), .B(A[317]), .Z(n2827) );
  NANDN U3743 ( .A(B[319]), .B(A[319]), .Z(n2819) );
  NANDN U3744 ( .A(B[321]), .B(A[321]), .Z(n2811) );
  NANDN U3745 ( .A(B[323]), .B(A[323]), .Z(n2803) );
  NANDN U3746 ( .A(B[325]), .B(A[325]), .Z(n2795) );
  NANDN U3747 ( .A(B[327]), .B(A[327]), .Z(n2787) );
  NANDN U3748 ( .A(B[329]), .B(A[329]), .Z(n2779) );
  NANDN U3749 ( .A(B[331]), .B(A[331]), .Z(n2771) );
  NANDN U3750 ( .A(B[333]), .B(A[333]), .Z(n2763) );
  NANDN U3751 ( .A(B[335]), .B(A[335]), .Z(n2755) );
  NANDN U3752 ( .A(B[337]), .B(A[337]), .Z(n2747) );
  NANDN U3753 ( .A(B[339]), .B(A[339]), .Z(n2739) );
  NANDN U3754 ( .A(B[341]), .B(A[341]), .Z(n2731) );
  NANDN U3755 ( .A(B[343]), .B(A[343]), .Z(n2723) );
  NANDN U3756 ( .A(B[345]), .B(A[345]), .Z(n2715) );
  NANDN U3757 ( .A(B[347]), .B(A[347]), .Z(n2707) );
  NANDN U3758 ( .A(B[349]), .B(A[349]), .Z(n2699) );
  NANDN U3759 ( .A(B[351]), .B(A[351]), .Z(n2691) );
  NANDN U3760 ( .A(B[353]), .B(A[353]), .Z(n2683) );
  NANDN U3761 ( .A(B[355]), .B(A[355]), .Z(n2675) );
  NANDN U3762 ( .A(B[357]), .B(A[357]), .Z(n2667) );
  NANDN U3763 ( .A(B[359]), .B(A[359]), .Z(n2659) );
  NANDN U3764 ( .A(B[361]), .B(A[361]), .Z(n2651) );
  NANDN U3765 ( .A(B[363]), .B(A[363]), .Z(n2643) );
  NANDN U3766 ( .A(B[365]), .B(A[365]), .Z(n2635) );
  NANDN U3767 ( .A(B[367]), .B(A[367]), .Z(n2627) );
  NANDN U3768 ( .A(B[369]), .B(A[369]), .Z(n2619) );
  NANDN U3769 ( .A(B[371]), .B(A[371]), .Z(n2611) );
  NANDN U3770 ( .A(B[373]), .B(A[373]), .Z(n2603) );
  NANDN U3771 ( .A(B[375]), .B(A[375]), .Z(n2595) );
  NANDN U3772 ( .A(B[377]), .B(A[377]), .Z(n2587) );
  NANDN U3773 ( .A(B[379]), .B(A[379]), .Z(n2579) );
  NANDN U3774 ( .A(B[381]), .B(A[381]), .Z(n2571) );
  NANDN U3775 ( .A(B[383]), .B(A[383]), .Z(n2563) );
  NANDN U3776 ( .A(B[385]), .B(A[385]), .Z(n2555) );
  NANDN U3777 ( .A(B[387]), .B(A[387]), .Z(n2547) );
  NANDN U3778 ( .A(B[389]), .B(A[389]), .Z(n2539) );
  NANDN U3779 ( .A(B[391]), .B(A[391]), .Z(n2531) );
  NANDN U3780 ( .A(B[393]), .B(A[393]), .Z(n2523) );
  NANDN U3781 ( .A(B[395]), .B(A[395]), .Z(n2515) );
  NANDN U3782 ( .A(B[397]), .B(A[397]), .Z(n2507) );
  NANDN U3783 ( .A(B[399]), .B(A[399]), .Z(n2499) );
  NANDN U3784 ( .A(B[401]), .B(A[401]), .Z(n2491) );
  NANDN U3785 ( .A(B[403]), .B(A[403]), .Z(n2483) );
  NANDN U3786 ( .A(B[405]), .B(A[405]), .Z(n2475) );
  NANDN U3787 ( .A(B[407]), .B(A[407]), .Z(n2467) );
  NANDN U3788 ( .A(B[409]), .B(A[409]), .Z(n2459) );
  NANDN U3789 ( .A(B[411]), .B(A[411]), .Z(n2451) );
  NANDN U3790 ( .A(B[413]), .B(A[413]), .Z(n2443) );
  NANDN U3791 ( .A(B[415]), .B(A[415]), .Z(n2435) );
  NANDN U3792 ( .A(B[417]), .B(A[417]), .Z(n2427) );
  NANDN U3793 ( .A(B[419]), .B(A[419]), .Z(n2419) );
  NANDN U3794 ( .A(B[421]), .B(A[421]), .Z(n2411) );
  NANDN U3795 ( .A(B[423]), .B(A[423]), .Z(n2403) );
  NANDN U3796 ( .A(B[425]), .B(A[425]), .Z(n2395) );
  NANDN U3797 ( .A(B[427]), .B(A[427]), .Z(n2387) );
  NANDN U3798 ( .A(B[429]), .B(A[429]), .Z(n2379) );
  NANDN U3799 ( .A(B[431]), .B(A[431]), .Z(n2371) );
  NANDN U3800 ( .A(B[433]), .B(A[433]), .Z(n2363) );
  NANDN U3801 ( .A(B[435]), .B(A[435]), .Z(n2355) );
  NANDN U3802 ( .A(B[437]), .B(A[437]), .Z(n2347) );
  NANDN U3803 ( .A(B[439]), .B(A[439]), .Z(n2339) );
  NANDN U3804 ( .A(B[441]), .B(A[441]), .Z(n2331) );
  NANDN U3805 ( .A(B[443]), .B(A[443]), .Z(n2323) );
  NANDN U3806 ( .A(B[445]), .B(A[445]), .Z(n2315) );
  NANDN U3807 ( .A(B[447]), .B(A[447]), .Z(n2307) );
  NANDN U3808 ( .A(B[449]), .B(A[449]), .Z(n2299) );
  NANDN U3809 ( .A(B[451]), .B(A[451]), .Z(n2291) );
  NANDN U3810 ( .A(B[453]), .B(A[453]), .Z(n2283) );
  NANDN U3811 ( .A(B[455]), .B(A[455]), .Z(n2275) );
  NANDN U3812 ( .A(B[457]), .B(A[457]), .Z(n2267) );
  NANDN U3813 ( .A(B[459]), .B(A[459]), .Z(n2259) );
  NANDN U3814 ( .A(B[461]), .B(A[461]), .Z(n2251) );
  NANDN U3815 ( .A(B[463]), .B(A[463]), .Z(n2243) );
  NANDN U3816 ( .A(B[465]), .B(A[465]), .Z(n2235) );
  NANDN U3817 ( .A(B[467]), .B(A[467]), .Z(n2227) );
  NANDN U3818 ( .A(B[469]), .B(A[469]), .Z(n2219) );
  NANDN U3819 ( .A(B[471]), .B(A[471]), .Z(n2211) );
  NANDN U3820 ( .A(B[473]), .B(A[473]), .Z(n2203) );
  NANDN U3821 ( .A(B[475]), .B(A[475]), .Z(n2195) );
  NANDN U3822 ( .A(B[477]), .B(A[477]), .Z(n2187) );
  NANDN U3823 ( .A(B[479]), .B(A[479]), .Z(n2179) );
  NANDN U3824 ( .A(B[481]), .B(A[481]), .Z(n2171) );
  NANDN U3825 ( .A(B[483]), .B(A[483]), .Z(n2163) );
  NANDN U3826 ( .A(B[485]), .B(A[485]), .Z(n2155) );
  NANDN U3827 ( .A(B[487]), .B(A[487]), .Z(n2147) );
  NANDN U3828 ( .A(B[489]), .B(A[489]), .Z(n2139) );
  NANDN U3829 ( .A(B[491]), .B(A[491]), .Z(n2131) );
  NANDN U3830 ( .A(B[493]), .B(A[493]), .Z(n2123) );
  NANDN U3831 ( .A(B[495]), .B(A[495]), .Z(n2115) );
  NANDN U3832 ( .A(B[497]), .B(A[497]), .Z(n2107) );
  NANDN U3833 ( .A(B[499]), .B(A[499]), .Z(n2099) );
  NANDN U3834 ( .A(B[501]), .B(A[501]), .Z(n2091) );
  NANDN U3835 ( .A(B[503]), .B(A[503]), .Z(n2083) );
  NANDN U3836 ( .A(B[505]), .B(A[505]), .Z(n2075) );
  NANDN U3837 ( .A(B[507]), .B(A[507]), .Z(n2067) );
  NANDN U3838 ( .A(B[509]), .B(A[509]), .Z(n2059) );
  NANDN U3839 ( .A(B[511]), .B(A[511]), .Z(n2051) );
  NANDN U3840 ( .A(B[513]), .B(A[513]), .Z(n2043) );
  NANDN U3841 ( .A(B[515]), .B(A[515]), .Z(n2035) );
  NANDN U3842 ( .A(B[517]), .B(A[517]), .Z(n2027) );
  NANDN U3843 ( .A(B[519]), .B(A[519]), .Z(n2019) );
  NANDN U3844 ( .A(B[521]), .B(A[521]), .Z(n2011) );
  NANDN U3845 ( .A(B[523]), .B(A[523]), .Z(n2003) );
  NANDN U3846 ( .A(B[525]), .B(A[525]), .Z(n1995) );
  NANDN U3847 ( .A(B[527]), .B(A[527]), .Z(n1987) );
  NANDN U3848 ( .A(B[529]), .B(A[529]), .Z(n1979) );
  NANDN U3849 ( .A(B[531]), .B(A[531]), .Z(n1971) );
  NANDN U3850 ( .A(B[533]), .B(A[533]), .Z(n1963) );
  NANDN U3851 ( .A(B[535]), .B(A[535]), .Z(n1955) );
  NANDN U3852 ( .A(B[537]), .B(A[537]), .Z(n1947) );
  NANDN U3853 ( .A(B[539]), .B(A[539]), .Z(n1939) );
  NANDN U3854 ( .A(B[541]), .B(A[541]), .Z(n1931) );
  NANDN U3855 ( .A(B[543]), .B(A[543]), .Z(n1923) );
  NANDN U3856 ( .A(B[545]), .B(A[545]), .Z(n1915) );
  NANDN U3857 ( .A(B[547]), .B(A[547]), .Z(n1907) );
  NANDN U3858 ( .A(B[549]), .B(A[549]), .Z(n1899) );
  NANDN U3859 ( .A(B[551]), .B(A[551]), .Z(n1891) );
  NANDN U3860 ( .A(B[553]), .B(A[553]), .Z(n1883) );
  NANDN U3861 ( .A(B[555]), .B(A[555]), .Z(n1875) );
  NANDN U3862 ( .A(B[557]), .B(A[557]), .Z(n1867) );
  NANDN U3863 ( .A(B[559]), .B(A[559]), .Z(n1859) );
  NANDN U3864 ( .A(B[561]), .B(A[561]), .Z(n1851) );
  NANDN U3865 ( .A(B[563]), .B(A[563]), .Z(n1843) );
  NANDN U3866 ( .A(B[565]), .B(A[565]), .Z(n1835) );
  NANDN U3867 ( .A(B[567]), .B(A[567]), .Z(n1827) );
  NANDN U3868 ( .A(B[569]), .B(A[569]), .Z(n1819) );
  NANDN U3869 ( .A(B[571]), .B(A[571]), .Z(n1811) );
  NANDN U3870 ( .A(B[573]), .B(A[573]), .Z(n1803) );
  NANDN U3871 ( .A(B[575]), .B(A[575]), .Z(n1795) );
  NANDN U3872 ( .A(B[577]), .B(A[577]), .Z(n1787) );
  NANDN U3873 ( .A(B[579]), .B(A[579]), .Z(n1779) );
  NANDN U3874 ( .A(B[581]), .B(A[581]), .Z(n1771) );
  NANDN U3875 ( .A(B[583]), .B(A[583]), .Z(n1763) );
  NANDN U3876 ( .A(B[585]), .B(A[585]), .Z(n1755) );
  NANDN U3877 ( .A(B[587]), .B(A[587]), .Z(n1747) );
  NANDN U3878 ( .A(B[589]), .B(A[589]), .Z(n1739) );
  NANDN U3879 ( .A(B[591]), .B(A[591]), .Z(n1731) );
  NANDN U3880 ( .A(B[593]), .B(A[593]), .Z(n1723) );
  NANDN U3881 ( .A(B[595]), .B(A[595]), .Z(n1715) );
  NANDN U3882 ( .A(B[597]), .B(A[597]), .Z(n1707) );
  NANDN U3883 ( .A(B[599]), .B(A[599]), .Z(n1699) );
  NANDN U3884 ( .A(B[601]), .B(A[601]), .Z(n1691) );
  NANDN U3885 ( .A(B[603]), .B(A[603]), .Z(n1683) );
  NANDN U3886 ( .A(B[605]), .B(A[605]), .Z(n1675) );
  NANDN U3887 ( .A(B[607]), .B(A[607]), .Z(n1667) );
  NANDN U3888 ( .A(B[609]), .B(A[609]), .Z(n1659) );
  NANDN U3889 ( .A(B[611]), .B(A[611]), .Z(n1651) );
  NANDN U3890 ( .A(B[613]), .B(A[613]), .Z(n1643) );
  NANDN U3891 ( .A(B[615]), .B(A[615]), .Z(n1635) );
  NANDN U3892 ( .A(B[617]), .B(A[617]), .Z(n1627) );
  NANDN U3893 ( .A(B[619]), .B(A[619]), .Z(n1619) );
  NANDN U3894 ( .A(B[621]), .B(A[621]), .Z(n1611) );
  NANDN U3895 ( .A(B[623]), .B(A[623]), .Z(n1603) );
  NANDN U3896 ( .A(B[625]), .B(A[625]), .Z(n1595) );
  NANDN U3897 ( .A(B[627]), .B(A[627]), .Z(n1587) );
  NANDN U3898 ( .A(B[629]), .B(A[629]), .Z(n1579) );
  NANDN U3899 ( .A(B[631]), .B(A[631]), .Z(n1571) );
  NANDN U3900 ( .A(B[633]), .B(A[633]), .Z(n1563) );
  NANDN U3901 ( .A(B[635]), .B(A[635]), .Z(n1555) );
  NANDN U3902 ( .A(B[637]), .B(A[637]), .Z(n1547) );
  NANDN U3903 ( .A(B[639]), .B(A[639]), .Z(n1539) );
  NANDN U3904 ( .A(B[641]), .B(A[641]), .Z(n1531) );
  NANDN U3905 ( .A(B[643]), .B(A[643]), .Z(n1523) );
  NANDN U3906 ( .A(B[645]), .B(A[645]), .Z(n1515) );
  NANDN U3907 ( .A(B[647]), .B(A[647]), .Z(n1507) );
  NANDN U3908 ( .A(B[649]), .B(A[649]), .Z(n1499) );
  NANDN U3909 ( .A(B[651]), .B(A[651]), .Z(n1491) );
  NANDN U3910 ( .A(B[653]), .B(A[653]), .Z(n1483) );
  NANDN U3911 ( .A(B[655]), .B(A[655]), .Z(n1475) );
  NANDN U3912 ( .A(B[657]), .B(A[657]), .Z(n1467) );
  NANDN U3913 ( .A(B[659]), .B(A[659]), .Z(n1459) );
  NANDN U3914 ( .A(B[661]), .B(A[661]), .Z(n1451) );
  NANDN U3915 ( .A(B[663]), .B(A[663]), .Z(n1443) );
  NANDN U3916 ( .A(B[665]), .B(A[665]), .Z(n1435) );
  NANDN U3917 ( .A(B[667]), .B(A[667]), .Z(n1427) );
  NANDN U3918 ( .A(B[669]), .B(A[669]), .Z(n1419) );
  NANDN U3919 ( .A(B[671]), .B(A[671]), .Z(n1411) );
  NANDN U3920 ( .A(B[673]), .B(A[673]), .Z(n1403) );
  NANDN U3921 ( .A(B[675]), .B(A[675]), .Z(n1395) );
  NANDN U3922 ( .A(B[677]), .B(A[677]), .Z(n1387) );
  NANDN U3923 ( .A(B[679]), .B(A[679]), .Z(n1379) );
  NANDN U3924 ( .A(B[681]), .B(A[681]), .Z(n1371) );
  NANDN U3925 ( .A(B[683]), .B(A[683]), .Z(n1363) );
  NANDN U3926 ( .A(B[685]), .B(A[685]), .Z(n1355) );
  NANDN U3927 ( .A(B[687]), .B(A[687]), .Z(n1347) );
  NANDN U3928 ( .A(B[689]), .B(A[689]), .Z(n1339) );
  NANDN U3929 ( .A(B[691]), .B(A[691]), .Z(n1331) );
  NANDN U3930 ( .A(B[693]), .B(A[693]), .Z(n1323) );
  NANDN U3931 ( .A(B[695]), .B(A[695]), .Z(n1315) );
  NANDN U3932 ( .A(B[697]), .B(A[697]), .Z(n1307) );
  NANDN U3933 ( .A(B[699]), .B(A[699]), .Z(n1299) );
  NANDN U3934 ( .A(B[701]), .B(A[701]), .Z(n1291) );
  NANDN U3935 ( .A(B[703]), .B(A[703]), .Z(n1283) );
  NANDN U3936 ( .A(B[705]), .B(A[705]), .Z(n1275) );
  NANDN U3937 ( .A(B[707]), .B(A[707]), .Z(n1267) );
  NANDN U3938 ( .A(B[709]), .B(A[709]), .Z(n1259) );
  NANDN U3939 ( .A(B[711]), .B(A[711]), .Z(n1251) );
  NANDN U3940 ( .A(B[713]), .B(A[713]), .Z(n1243) );
  NANDN U3941 ( .A(B[715]), .B(A[715]), .Z(n1235) );
  NANDN U3942 ( .A(B[717]), .B(A[717]), .Z(n1227) );
  NANDN U3943 ( .A(B[719]), .B(A[719]), .Z(n1219) );
  NANDN U3944 ( .A(B[721]), .B(A[721]), .Z(n1211) );
  NANDN U3945 ( .A(B[723]), .B(A[723]), .Z(n1203) );
  NANDN U3946 ( .A(B[725]), .B(A[725]), .Z(n1195) );
  NANDN U3947 ( .A(B[727]), .B(A[727]), .Z(n1187) );
  NANDN U3948 ( .A(B[729]), .B(A[729]), .Z(n1179) );
  NANDN U3949 ( .A(B[731]), .B(A[731]), .Z(n1171) );
  NANDN U3950 ( .A(B[733]), .B(A[733]), .Z(n1163) );
  NANDN U3951 ( .A(B[735]), .B(A[735]), .Z(n1155) );
  NANDN U3952 ( .A(B[737]), .B(A[737]), .Z(n1147) );
  NANDN U3953 ( .A(B[739]), .B(A[739]), .Z(n1139) );
  NANDN U3954 ( .A(B[741]), .B(A[741]), .Z(n1131) );
  NANDN U3955 ( .A(B[743]), .B(A[743]), .Z(n1123) );
  NANDN U3956 ( .A(B[745]), .B(A[745]), .Z(n1115) );
  NANDN U3957 ( .A(B[747]), .B(A[747]), .Z(n1107) );
  NANDN U3958 ( .A(B[749]), .B(A[749]), .Z(n1099) );
  NANDN U3959 ( .A(B[751]), .B(A[751]), .Z(n1091) );
  NANDN U3960 ( .A(B[753]), .B(A[753]), .Z(n1083) );
  NANDN U3961 ( .A(B[755]), .B(A[755]), .Z(n1075) );
  NANDN U3962 ( .A(B[757]), .B(A[757]), .Z(n1067) );
  NANDN U3963 ( .A(B[759]), .B(A[759]), .Z(n1059) );
  NANDN U3964 ( .A(B[761]), .B(A[761]), .Z(n1051) );
  NANDN U3965 ( .A(B[763]), .B(A[763]), .Z(n1043) );
  NANDN U3966 ( .A(B[765]), .B(A[765]), .Z(n1035) );
  NANDN U3967 ( .A(B[767]), .B(A[767]), .Z(n1027) );
  NANDN U3968 ( .A(B[769]), .B(A[769]), .Z(n1019) );
  NANDN U3969 ( .A(B[771]), .B(A[771]), .Z(n1011) );
  NANDN U3970 ( .A(B[773]), .B(A[773]), .Z(n1003) );
  NANDN U3971 ( .A(B[775]), .B(A[775]), .Z(n995) );
  NANDN U3972 ( .A(B[777]), .B(A[777]), .Z(n987) );
  NANDN U3973 ( .A(B[779]), .B(A[779]), .Z(n979) );
  NANDN U3974 ( .A(B[781]), .B(A[781]), .Z(n971) );
  NANDN U3975 ( .A(B[783]), .B(A[783]), .Z(n963) );
  NANDN U3976 ( .A(B[785]), .B(A[785]), .Z(n955) );
  NANDN U3977 ( .A(B[787]), .B(A[787]), .Z(n947) );
  NANDN U3978 ( .A(B[789]), .B(A[789]), .Z(n939) );
  NANDN U3979 ( .A(B[791]), .B(A[791]), .Z(n931) );
  NANDN U3980 ( .A(B[793]), .B(A[793]), .Z(n923) );
  NANDN U3981 ( .A(B[795]), .B(A[795]), .Z(n915) );
  NANDN U3982 ( .A(B[797]), .B(A[797]), .Z(n907) );
  NANDN U3983 ( .A(B[799]), .B(A[799]), .Z(n899) );
  NANDN U3984 ( .A(B[801]), .B(A[801]), .Z(n891) );
  NANDN U3985 ( .A(B[803]), .B(A[803]), .Z(n883) );
  NANDN U3986 ( .A(B[805]), .B(A[805]), .Z(n875) );
  NANDN U3987 ( .A(B[807]), .B(A[807]), .Z(n867) );
  NANDN U3988 ( .A(B[809]), .B(A[809]), .Z(n859) );
  NANDN U3989 ( .A(B[811]), .B(A[811]), .Z(n851) );
  NANDN U3990 ( .A(B[813]), .B(A[813]), .Z(n843) );
  NANDN U3991 ( .A(B[815]), .B(A[815]), .Z(n835) );
  NANDN U3992 ( .A(B[817]), .B(A[817]), .Z(n827) );
  NANDN U3993 ( .A(B[819]), .B(A[819]), .Z(n819) );
  NANDN U3994 ( .A(B[821]), .B(A[821]), .Z(n811) );
  NANDN U3995 ( .A(B[823]), .B(A[823]), .Z(n803) );
  NANDN U3996 ( .A(B[825]), .B(A[825]), .Z(n795) );
  NANDN U3997 ( .A(B[827]), .B(A[827]), .Z(n787) );
  NANDN U3998 ( .A(B[829]), .B(A[829]), .Z(n779) );
  NANDN U3999 ( .A(B[831]), .B(A[831]), .Z(n771) );
  NANDN U4000 ( .A(B[833]), .B(A[833]), .Z(n763) );
  NANDN U4001 ( .A(B[835]), .B(A[835]), .Z(n755) );
  NANDN U4002 ( .A(B[837]), .B(A[837]), .Z(n747) );
  NANDN U4003 ( .A(B[839]), .B(A[839]), .Z(n739) );
  NANDN U4004 ( .A(B[841]), .B(A[841]), .Z(n731) );
  NANDN U4005 ( .A(B[843]), .B(A[843]), .Z(n723) );
  NANDN U4006 ( .A(B[845]), .B(A[845]), .Z(n715) );
  NANDN U4007 ( .A(B[847]), .B(A[847]), .Z(n707) );
  NANDN U4008 ( .A(B[849]), .B(A[849]), .Z(n699) );
  NANDN U4009 ( .A(B[851]), .B(A[851]), .Z(n691) );
  NANDN U4010 ( .A(B[853]), .B(A[853]), .Z(n683) );
  NANDN U4011 ( .A(B[855]), .B(A[855]), .Z(n675) );
  NANDN U4012 ( .A(B[857]), .B(A[857]), .Z(n667) );
  NANDN U4013 ( .A(B[859]), .B(A[859]), .Z(n659) );
  NANDN U4014 ( .A(B[861]), .B(A[861]), .Z(n651) );
  NANDN U4015 ( .A(B[863]), .B(A[863]), .Z(n643) );
  NANDN U4016 ( .A(B[865]), .B(A[865]), .Z(n635) );
  NANDN U4017 ( .A(B[867]), .B(A[867]), .Z(n627) );
  NANDN U4018 ( .A(B[869]), .B(A[869]), .Z(n619) );
  NANDN U4019 ( .A(B[871]), .B(A[871]), .Z(n611) );
  NANDN U4020 ( .A(B[873]), .B(A[873]), .Z(n603) );
  NANDN U4021 ( .A(B[875]), .B(A[875]), .Z(n595) );
  NANDN U4022 ( .A(B[877]), .B(A[877]), .Z(n587) );
  NANDN U4023 ( .A(B[879]), .B(A[879]), .Z(n579) );
  NANDN U4024 ( .A(B[881]), .B(A[881]), .Z(n571) );
  NANDN U4025 ( .A(B[883]), .B(A[883]), .Z(n563) );
  NANDN U4026 ( .A(B[885]), .B(A[885]), .Z(n555) );
  NANDN U4027 ( .A(B[887]), .B(A[887]), .Z(n547) );
  NANDN U4028 ( .A(B[889]), .B(A[889]), .Z(n539) );
  NANDN U4029 ( .A(B[891]), .B(A[891]), .Z(n531) );
  NANDN U4030 ( .A(B[893]), .B(A[893]), .Z(n523) );
  NANDN U4031 ( .A(B[895]), .B(A[895]), .Z(n515) );
  NANDN U4032 ( .A(B[897]), .B(A[897]), .Z(n507) );
  NANDN U4033 ( .A(B[899]), .B(A[899]), .Z(n499) );
  NANDN U4034 ( .A(B[901]), .B(A[901]), .Z(n491) );
  NANDN U4035 ( .A(B[903]), .B(A[903]), .Z(n483) );
  NANDN U4036 ( .A(B[905]), .B(A[905]), .Z(n475) );
  NANDN U4037 ( .A(B[907]), .B(A[907]), .Z(n467) );
  NANDN U4038 ( .A(B[909]), .B(A[909]), .Z(n459) );
  NANDN U4039 ( .A(B[911]), .B(A[911]), .Z(n451) );
  NANDN U4040 ( .A(B[913]), .B(A[913]), .Z(n443) );
  NANDN U4041 ( .A(B[915]), .B(A[915]), .Z(n435) );
  NANDN U4042 ( .A(B[917]), .B(A[917]), .Z(n427) );
  NANDN U4043 ( .A(B[919]), .B(A[919]), .Z(n419) );
  NANDN U4044 ( .A(B[921]), .B(A[921]), .Z(n411) );
  NANDN U4045 ( .A(B[923]), .B(A[923]), .Z(n403) );
  NANDN U4046 ( .A(B[925]), .B(A[925]), .Z(n395) );
  NANDN U4047 ( .A(B[927]), .B(A[927]), .Z(n387) );
  NANDN U4048 ( .A(B[929]), .B(A[929]), .Z(n379) );
  NANDN U4049 ( .A(B[931]), .B(A[931]), .Z(n371) );
  NANDN U4050 ( .A(B[933]), .B(A[933]), .Z(n363) );
  NANDN U4051 ( .A(B[935]), .B(A[935]), .Z(n355) );
  NANDN U4052 ( .A(B[937]), .B(A[937]), .Z(n347) );
  NANDN U4053 ( .A(B[939]), .B(A[939]), .Z(n339) );
  NANDN U4054 ( .A(B[941]), .B(A[941]), .Z(n331) );
  NANDN U4055 ( .A(B[943]), .B(A[943]), .Z(n323) );
  NANDN U4056 ( .A(B[945]), .B(A[945]), .Z(n315) );
  NANDN U4057 ( .A(B[947]), .B(A[947]), .Z(n307) );
  NANDN U4058 ( .A(B[949]), .B(A[949]), .Z(n299) );
  NANDN U4059 ( .A(B[951]), .B(A[951]), .Z(n291) );
  NANDN U4060 ( .A(B[953]), .B(A[953]), .Z(n283) );
  NANDN U4061 ( .A(B[955]), .B(A[955]), .Z(n275) );
  NANDN U4062 ( .A(B[957]), .B(A[957]), .Z(n267) );
  NANDN U4063 ( .A(B[959]), .B(A[959]), .Z(n259) );
  NANDN U4064 ( .A(B[961]), .B(A[961]), .Z(n251) );
  NANDN U4065 ( .A(B[963]), .B(A[963]), .Z(n243) );
  NANDN U4066 ( .A(B[965]), .B(A[965]), .Z(n235) );
  NANDN U4067 ( .A(B[967]), .B(A[967]), .Z(n227) );
  NANDN U4068 ( .A(B[969]), .B(A[969]), .Z(n219) );
  NANDN U4069 ( .A(B[971]), .B(A[971]), .Z(n211) );
  NANDN U4070 ( .A(B[973]), .B(A[973]), .Z(n203) );
  NANDN U4071 ( .A(B[975]), .B(A[975]), .Z(n195) );
  NANDN U4072 ( .A(B[977]), .B(A[977]), .Z(n187) );
  NANDN U4073 ( .A(B[979]), .B(A[979]), .Z(n179) );
  NANDN U4074 ( .A(B[981]), .B(A[981]), .Z(n171) );
  NANDN U4075 ( .A(B[983]), .B(A[983]), .Z(n163) );
  NANDN U4076 ( .A(B[985]), .B(A[985]), .Z(n155) );
  NANDN U4077 ( .A(B[987]), .B(A[987]), .Z(n147) );
  NANDN U4078 ( .A(B[989]), .B(A[989]), .Z(n139) );
  NANDN U4079 ( .A(B[991]), .B(A[991]), .Z(n131) );
  NANDN U4080 ( .A(B[993]), .B(A[993]), .Z(n123) );
  NANDN U4081 ( .A(B[995]), .B(A[995]), .Z(n115) );
  NANDN U4082 ( .A(B[997]), .B(A[997]), .Z(n107) );
  NANDN U4083 ( .A(B[1000]), .B(A[1000]), .Z(n99) );
  NANDN U4084 ( .A(B[1001]), .B(A[1001]), .Z(n91) );
  NANDN U4085 ( .A(B[1003]), .B(A[1003]), .Z(n83) );
  NANDN U4086 ( .A(B[1005]), .B(A[1005]), .Z(n75) );
  NANDN U4087 ( .A(B[1007]), .B(A[1007]), .Z(n67) );
  NANDN U4088 ( .A(B[1009]), .B(A[1009]), .Z(n59) );
  NANDN U4089 ( .A(B[1011]), .B(A[1011]), .Z(n51) );
  NANDN U4090 ( .A(B[1013]), .B(A[1013]), .Z(n43) );
  NANDN U4091 ( .A(B[1015]), .B(A[1015]), .Z(n35) );
  NANDN U4092 ( .A(B[1017]), .B(A[1017]), .Z(n27) );
  NANDN U4093 ( .A(B[1019]), .B(A[1019]), .Z(n19) );
  NANDN U4094 ( .A(B[1021]), .B(A[1021]), .Z(n11) );
  NANDN U4095 ( .A(A[1023]), .B(B[1023]), .Z(n3) );
endmodule


module modmult_step_N1024_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [1025:0] A;
  input [1025:0] B;
  output [1025:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120;

  IV U1 ( .A(A[1]), .Z(n1) );
  IV U2 ( .A(n5119), .Z(n2) );
  XNOR U3 ( .A(n3), .B(n4), .Z(DIFF[9]) );
  XOR U4 ( .A(B[9]), .B(A[9]), .Z(n4) );
  XNOR U5 ( .A(n5), .B(n6), .Z(DIFF[99]) );
  XOR U6 ( .A(B[99]), .B(A[99]), .Z(n6) );
  XNOR U7 ( .A(n7), .B(n8), .Z(DIFF[999]) );
  XOR U8 ( .A(B[999]), .B(A[999]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(DIFF[998]) );
  XOR U10 ( .A(B[998]), .B(A[998]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(DIFF[997]) );
  XOR U12 ( .A(B[997]), .B(A[997]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(DIFF[996]) );
  XOR U14 ( .A(B[996]), .B(A[996]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(DIFF[995]) );
  XOR U16 ( .A(B[995]), .B(A[995]), .Z(n16) );
  XOR U17 ( .A(n17), .B(n18), .Z(DIFF[994]) );
  XOR U18 ( .A(B[994]), .B(A[994]), .Z(n18) );
  XOR U19 ( .A(n19), .B(n20), .Z(DIFF[993]) );
  XOR U20 ( .A(B[993]), .B(A[993]), .Z(n20) );
  XOR U21 ( .A(n21), .B(n22), .Z(DIFF[992]) );
  XOR U22 ( .A(B[992]), .B(A[992]), .Z(n22) );
  XOR U23 ( .A(n23), .B(n24), .Z(DIFF[991]) );
  XOR U24 ( .A(B[991]), .B(A[991]), .Z(n24) );
  XOR U25 ( .A(n25), .B(n26), .Z(DIFF[990]) );
  XOR U26 ( .A(B[990]), .B(A[990]), .Z(n26) );
  XOR U27 ( .A(n27), .B(n28), .Z(DIFF[98]) );
  XOR U28 ( .A(B[98]), .B(A[98]), .Z(n28) );
  XOR U29 ( .A(n29), .B(n30), .Z(DIFF[989]) );
  XOR U30 ( .A(B[989]), .B(A[989]), .Z(n30) );
  XOR U31 ( .A(n31), .B(n32), .Z(DIFF[988]) );
  XOR U32 ( .A(B[988]), .B(A[988]), .Z(n32) );
  XOR U33 ( .A(n33), .B(n34), .Z(DIFF[987]) );
  XOR U34 ( .A(B[987]), .B(A[987]), .Z(n34) );
  XOR U35 ( .A(n35), .B(n36), .Z(DIFF[986]) );
  XOR U36 ( .A(B[986]), .B(A[986]), .Z(n36) );
  XOR U37 ( .A(n37), .B(n38), .Z(DIFF[985]) );
  XOR U38 ( .A(B[985]), .B(A[985]), .Z(n38) );
  XOR U39 ( .A(n39), .B(n40), .Z(DIFF[984]) );
  XOR U40 ( .A(B[984]), .B(A[984]), .Z(n40) );
  XOR U41 ( .A(n41), .B(n42), .Z(DIFF[983]) );
  XOR U42 ( .A(B[983]), .B(A[983]), .Z(n42) );
  XOR U43 ( .A(n43), .B(n44), .Z(DIFF[982]) );
  XOR U44 ( .A(B[982]), .B(A[982]), .Z(n44) );
  XOR U45 ( .A(n45), .B(n46), .Z(DIFF[981]) );
  XOR U46 ( .A(B[981]), .B(A[981]), .Z(n46) );
  XOR U47 ( .A(n47), .B(n48), .Z(DIFF[980]) );
  XOR U48 ( .A(B[980]), .B(A[980]), .Z(n48) );
  XOR U49 ( .A(n49), .B(n50), .Z(DIFF[97]) );
  XOR U50 ( .A(B[97]), .B(A[97]), .Z(n50) );
  XOR U51 ( .A(n51), .B(n52), .Z(DIFF[979]) );
  XOR U52 ( .A(B[979]), .B(A[979]), .Z(n52) );
  XOR U53 ( .A(n53), .B(n54), .Z(DIFF[978]) );
  XOR U54 ( .A(B[978]), .B(A[978]), .Z(n54) );
  XOR U55 ( .A(n55), .B(n56), .Z(DIFF[977]) );
  XOR U56 ( .A(B[977]), .B(A[977]), .Z(n56) );
  XOR U57 ( .A(n57), .B(n58), .Z(DIFF[976]) );
  XOR U58 ( .A(B[976]), .B(A[976]), .Z(n58) );
  XOR U59 ( .A(n59), .B(n60), .Z(DIFF[975]) );
  XOR U60 ( .A(B[975]), .B(A[975]), .Z(n60) );
  XOR U61 ( .A(n61), .B(n62), .Z(DIFF[974]) );
  XOR U62 ( .A(B[974]), .B(A[974]), .Z(n62) );
  XOR U63 ( .A(n63), .B(n64), .Z(DIFF[973]) );
  XOR U64 ( .A(B[973]), .B(A[973]), .Z(n64) );
  XOR U65 ( .A(n65), .B(n66), .Z(DIFF[972]) );
  XOR U66 ( .A(B[972]), .B(A[972]), .Z(n66) );
  XOR U67 ( .A(n67), .B(n68), .Z(DIFF[971]) );
  XOR U68 ( .A(B[971]), .B(A[971]), .Z(n68) );
  XOR U69 ( .A(n69), .B(n70), .Z(DIFF[970]) );
  XOR U70 ( .A(B[970]), .B(A[970]), .Z(n70) );
  XOR U71 ( .A(n71), .B(n72), .Z(DIFF[96]) );
  XOR U72 ( .A(B[96]), .B(A[96]), .Z(n72) );
  XOR U73 ( .A(n73), .B(n74), .Z(DIFF[969]) );
  XOR U74 ( .A(B[969]), .B(A[969]), .Z(n74) );
  XOR U75 ( .A(n75), .B(n76), .Z(DIFF[968]) );
  XOR U76 ( .A(B[968]), .B(A[968]), .Z(n76) );
  XOR U77 ( .A(n77), .B(n78), .Z(DIFF[967]) );
  XOR U78 ( .A(B[967]), .B(A[967]), .Z(n78) );
  XOR U79 ( .A(n79), .B(n80), .Z(DIFF[966]) );
  XOR U80 ( .A(B[966]), .B(A[966]), .Z(n80) );
  XOR U81 ( .A(n81), .B(n82), .Z(DIFF[965]) );
  XOR U82 ( .A(B[965]), .B(A[965]), .Z(n82) );
  XOR U83 ( .A(n83), .B(n84), .Z(DIFF[964]) );
  XOR U84 ( .A(B[964]), .B(A[964]), .Z(n84) );
  XOR U85 ( .A(n85), .B(n86), .Z(DIFF[963]) );
  XOR U86 ( .A(B[963]), .B(A[963]), .Z(n86) );
  XOR U87 ( .A(n87), .B(n88), .Z(DIFF[962]) );
  XOR U88 ( .A(B[962]), .B(A[962]), .Z(n88) );
  XOR U89 ( .A(n89), .B(n90), .Z(DIFF[961]) );
  XOR U90 ( .A(B[961]), .B(A[961]), .Z(n90) );
  XOR U91 ( .A(n91), .B(n92), .Z(DIFF[960]) );
  XOR U92 ( .A(B[960]), .B(A[960]), .Z(n92) );
  XOR U93 ( .A(n93), .B(n94), .Z(DIFF[95]) );
  XOR U94 ( .A(B[95]), .B(A[95]), .Z(n94) );
  XOR U95 ( .A(n95), .B(n96), .Z(DIFF[959]) );
  XOR U96 ( .A(B[959]), .B(A[959]), .Z(n96) );
  XOR U97 ( .A(n97), .B(n98), .Z(DIFF[958]) );
  XOR U98 ( .A(B[958]), .B(A[958]), .Z(n98) );
  XOR U99 ( .A(n99), .B(n100), .Z(DIFF[957]) );
  XOR U100 ( .A(B[957]), .B(A[957]), .Z(n100) );
  XOR U101 ( .A(n101), .B(n102), .Z(DIFF[956]) );
  XOR U102 ( .A(B[956]), .B(A[956]), .Z(n102) );
  XOR U103 ( .A(n103), .B(n104), .Z(DIFF[955]) );
  XOR U104 ( .A(B[955]), .B(A[955]), .Z(n104) );
  XOR U105 ( .A(n105), .B(n106), .Z(DIFF[954]) );
  XOR U106 ( .A(B[954]), .B(A[954]), .Z(n106) );
  XOR U107 ( .A(n107), .B(n108), .Z(DIFF[953]) );
  XOR U108 ( .A(B[953]), .B(A[953]), .Z(n108) );
  XOR U109 ( .A(n109), .B(n110), .Z(DIFF[952]) );
  XOR U110 ( .A(B[952]), .B(A[952]), .Z(n110) );
  XOR U111 ( .A(n111), .B(n112), .Z(DIFF[951]) );
  XOR U112 ( .A(B[951]), .B(A[951]), .Z(n112) );
  XOR U113 ( .A(n113), .B(n114), .Z(DIFF[950]) );
  XOR U114 ( .A(B[950]), .B(A[950]), .Z(n114) );
  XOR U115 ( .A(n115), .B(n116), .Z(DIFF[94]) );
  XOR U116 ( .A(B[94]), .B(A[94]), .Z(n116) );
  XOR U117 ( .A(n117), .B(n118), .Z(DIFF[949]) );
  XOR U118 ( .A(B[949]), .B(A[949]), .Z(n118) );
  XOR U119 ( .A(n119), .B(n120), .Z(DIFF[948]) );
  XOR U120 ( .A(B[948]), .B(A[948]), .Z(n120) );
  XOR U121 ( .A(n121), .B(n122), .Z(DIFF[947]) );
  XOR U122 ( .A(B[947]), .B(A[947]), .Z(n122) );
  XOR U123 ( .A(n123), .B(n124), .Z(DIFF[946]) );
  XOR U124 ( .A(B[946]), .B(A[946]), .Z(n124) );
  XOR U125 ( .A(n125), .B(n126), .Z(DIFF[945]) );
  XOR U126 ( .A(B[945]), .B(A[945]), .Z(n126) );
  XOR U127 ( .A(n127), .B(n128), .Z(DIFF[944]) );
  XOR U128 ( .A(B[944]), .B(A[944]), .Z(n128) );
  XOR U129 ( .A(n129), .B(n130), .Z(DIFF[943]) );
  XOR U130 ( .A(B[943]), .B(A[943]), .Z(n130) );
  XOR U131 ( .A(n131), .B(n132), .Z(DIFF[942]) );
  XOR U132 ( .A(B[942]), .B(A[942]), .Z(n132) );
  XOR U133 ( .A(n133), .B(n134), .Z(DIFF[941]) );
  XOR U134 ( .A(B[941]), .B(A[941]), .Z(n134) );
  XOR U135 ( .A(n135), .B(n136), .Z(DIFF[940]) );
  XOR U136 ( .A(B[940]), .B(A[940]), .Z(n136) );
  XOR U137 ( .A(n137), .B(n138), .Z(DIFF[93]) );
  XOR U138 ( .A(B[93]), .B(A[93]), .Z(n138) );
  XOR U139 ( .A(n139), .B(n140), .Z(DIFF[939]) );
  XOR U140 ( .A(B[939]), .B(A[939]), .Z(n140) );
  XOR U141 ( .A(n141), .B(n142), .Z(DIFF[938]) );
  XOR U142 ( .A(B[938]), .B(A[938]), .Z(n142) );
  XOR U143 ( .A(n143), .B(n144), .Z(DIFF[937]) );
  XOR U144 ( .A(B[937]), .B(A[937]), .Z(n144) );
  XOR U145 ( .A(n145), .B(n146), .Z(DIFF[936]) );
  XOR U146 ( .A(B[936]), .B(A[936]), .Z(n146) );
  XOR U147 ( .A(n147), .B(n148), .Z(DIFF[935]) );
  XOR U148 ( .A(B[935]), .B(A[935]), .Z(n148) );
  XOR U149 ( .A(n149), .B(n150), .Z(DIFF[934]) );
  XOR U150 ( .A(B[934]), .B(A[934]), .Z(n150) );
  XOR U151 ( .A(n151), .B(n152), .Z(DIFF[933]) );
  XOR U152 ( .A(B[933]), .B(A[933]), .Z(n152) );
  XOR U153 ( .A(n153), .B(n154), .Z(DIFF[932]) );
  XOR U154 ( .A(B[932]), .B(A[932]), .Z(n154) );
  XOR U155 ( .A(n155), .B(n156), .Z(DIFF[931]) );
  XOR U156 ( .A(B[931]), .B(A[931]), .Z(n156) );
  XOR U157 ( .A(n157), .B(n158), .Z(DIFF[930]) );
  XOR U158 ( .A(B[930]), .B(A[930]), .Z(n158) );
  XOR U159 ( .A(n159), .B(n160), .Z(DIFF[92]) );
  XOR U160 ( .A(B[92]), .B(A[92]), .Z(n160) );
  XOR U161 ( .A(n161), .B(n162), .Z(DIFF[929]) );
  XOR U162 ( .A(B[929]), .B(A[929]), .Z(n162) );
  XOR U163 ( .A(n163), .B(n164), .Z(DIFF[928]) );
  XOR U164 ( .A(B[928]), .B(A[928]), .Z(n164) );
  XOR U165 ( .A(n165), .B(n166), .Z(DIFF[927]) );
  XOR U166 ( .A(B[927]), .B(A[927]), .Z(n166) );
  XOR U167 ( .A(n167), .B(n168), .Z(DIFF[926]) );
  XOR U168 ( .A(B[926]), .B(A[926]), .Z(n168) );
  XOR U169 ( .A(n169), .B(n170), .Z(DIFF[925]) );
  XOR U170 ( .A(B[925]), .B(A[925]), .Z(n170) );
  XOR U171 ( .A(n171), .B(n172), .Z(DIFF[924]) );
  XOR U172 ( .A(B[924]), .B(A[924]), .Z(n172) );
  XOR U173 ( .A(n173), .B(n174), .Z(DIFF[923]) );
  XOR U174 ( .A(B[923]), .B(A[923]), .Z(n174) );
  XOR U175 ( .A(n175), .B(n176), .Z(DIFF[922]) );
  XOR U176 ( .A(B[922]), .B(A[922]), .Z(n176) );
  XOR U177 ( .A(n177), .B(n178), .Z(DIFF[921]) );
  XOR U178 ( .A(B[921]), .B(A[921]), .Z(n178) );
  XOR U179 ( .A(n179), .B(n180), .Z(DIFF[920]) );
  XOR U180 ( .A(B[920]), .B(A[920]), .Z(n180) );
  XOR U181 ( .A(n181), .B(n182), .Z(DIFF[91]) );
  XOR U182 ( .A(B[91]), .B(A[91]), .Z(n182) );
  XOR U183 ( .A(n183), .B(n184), .Z(DIFF[919]) );
  XOR U184 ( .A(B[919]), .B(A[919]), .Z(n184) );
  XOR U185 ( .A(n185), .B(n186), .Z(DIFF[918]) );
  XOR U186 ( .A(B[918]), .B(A[918]), .Z(n186) );
  XOR U187 ( .A(n187), .B(n188), .Z(DIFF[917]) );
  XOR U188 ( .A(B[917]), .B(A[917]), .Z(n188) );
  XOR U189 ( .A(n189), .B(n190), .Z(DIFF[916]) );
  XOR U190 ( .A(B[916]), .B(A[916]), .Z(n190) );
  XOR U191 ( .A(n191), .B(n192), .Z(DIFF[915]) );
  XOR U192 ( .A(B[915]), .B(A[915]), .Z(n192) );
  XOR U193 ( .A(n193), .B(n194), .Z(DIFF[914]) );
  XOR U194 ( .A(B[914]), .B(A[914]), .Z(n194) );
  XOR U195 ( .A(n195), .B(n196), .Z(DIFF[913]) );
  XOR U196 ( .A(B[913]), .B(A[913]), .Z(n196) );
  XOR U197 ( .A(n197), .B(n198), .Z(DIFF[912]) );
  XOR U198 ( .A(B[912]), .B(A[912]), .Z(n198) );
  XOR U199 ( .A(n199), .B(n200), .Z(DIFF[911]) );
  XOR U200 ( .A(B[911]), .B(A[911]), .Z(n200) );
  XOR U201 ( .A(n201), .B(n202), .Z(DIFF[910]) );
  XOR U202 ( .A(B[910]), .B(A[910]), .Z(n202) );
  XOR U203 ( .A(n203), .B(n204), .Z(DIFF[90]) );
  XOR U204 ( .A(B[90]), .B(A[90]), .Z(n204) );
  XOR U205 ( .A(n205), .B(n206), .Z(DIFF[909]) );
  XOR U206 ( .A(B[909]), .B(A[909]), .Z(n206) );
  XOR U207 ( .A(n207), .B(n208), .Z(DIFF[908]) );
  XOR U208 ( .A(B[908]), .B(A[908]), .Z(n208) );
  XOR U209 ( .A(n209), .B(n210), .Z(DIFF[907]) );
  XOR U210 ( .A(B[907]), .B(A[907]), .Z(n210) );
  XOR U211 ( .A(n211), .B(n212), .Z(DIFF[906]) );
  XOR U212 ( .A(B[906]), .B(A[906]), .Z(n212) );
  XOR U213 ( .A(n213), .B(n214), .Z(DIFF[905]) );
  XOR U214 ( .A(B[905]), .B(A[905]), .Z(n214) );
  XOR U215 ( .A(n215), .B(n216), .Z(DIFF[904]) );
  XOR U216 ( .A(B[904]), .B(A[904]), .Z(n216) );
  XOR U217 ( .A(n217), .B(n218), .Z(DIFF[903]) );
  XOR U218 ( .A(B[903]), .B(A[903]), .Z(n218) );
  XOR U219 ( .A(n219), .B(n220), .Z(DIFF[902]) );
  XOR U220 ( .A(B[902]), .B(A[902]), .Z(n220) );
  XOR U221 ( .A(n221), .B(n222), .Z(DIFF[901]) );
  XOR U222 ( .A(B[901]), .B(A[901]), .Z(n222) );
  XOR U223 ( .A(n223), .B(n224), .Z(DIFF[900]) );
  XOR U224 ( .A(B[900]), .B(A[900]), .Z(n224) );
  XOR U225 ( .A(n225), .B(n226), .Z(DIFF[8]) );
  XOR U226 ( .A(B[8]), .B(A[8]), .Z(n226) );
  XOR U227 ( .A(n227), .B(n228), .Z(DIFF[89]) );
  XOR U228 ( .A(B[89]), .B(A[89]), .Z(n228) );
  XOR U229 ( .A(n229), .B(n230), .Z(DIFF[899]) );
  XOR U230 ( .A(B[899]), .B(A[899]), .Z(n230) );
  XOR U231 ( .A(n231), .B(n232), .Z(DIFF[898]) );
  XOR U232 ( .A(B[898]), .B(A[898]), .Z(n232) );
  XOR U233 ( .A(n233), .B(n234), .Z(DIFF[897]) );
  XOR U234 ( .A(B[897]), .B(A[897]), .Z(n234) );
  XOR U235 ( .A(n235), .B(n236), .Z(DIFF[896]) );
  XOR U236 ( .A(B[896]), .B(A[896]), .Z(n236) );
  XOR U237 ( .A(n237), .B(n238), .Z(DIFF[895]) );
  XOR U238 ( .A(B[895]), .B(A[895]), .Z(n238) );
  XOR U239 ( .A(n239), .B(n240), .Z(DIFF[894]) );
  XOR U240 ( .A(B[894]), .B(A[894]), .Z(n240) );
  XOR U241 ( .A(n241), .B(n242), .Z(DIFF[893]) );
  XOR U242 ( .A(B[893]), .B(A[893]), .Z(n242) );
  XOR U243 ( .A(n243), .B(n244), .Z(DIFF[892]) );
  XOR U244 ( .A(B[892]), .B(A[892]), .Z(n244) );
  XOR U245 ( .A(n245), .B(n246), .Z(DIFF[891]) );
  XOR U246 ( .A(B[891]), .B(A[891]), .Z(n246) );
  XOR U247 ( .A(n247), .B(n248), .Z(DIFF[890]) );
  XOR U248 ( .A(B[890]), .B(A[890]), .Z(n248) );
  XOR U249 ( .A(n249), .B(n250), .Z(DIFF[88]) );
  XOR U250 ( .A(B[88]), .B(A[88]), .Z(n250) );
  XOR U251 ( .A(n251), .B(n252), .Z(DIFF[889]) );
  XOR U252 ( .A(B[889]), .B(A[889]), .Z(n252) );
  XOR U253 ( .A(n253), .B(n254), .Z(DIFF[888]) );
  XOR U254 ( .A(B[888]), .B(A[888]), .Z(n254) );
  XOR U255 ( .A(n255), .B(n256), .Z(DIFF[887]) );
  XOR U256 ( .A(B[887]), .B(A[887]), .Z(n256) );
  XOR U257 ( .A(n257), .B(n258), .Z(DIFF[886]) );
  XOR U258 ( .A(B[886]), .B(A[886]), .Z(n258) );
  XOR U259 ( .A(n259), .B(n260), .Z(DIFF[885]) );
  XOR U260 ( .A(B[885]), .B(A[885]), .Z(n260) );
  XOR U261 ( .A(n261), .B(n262), .Z(DIFF[884]) );
  XOR U262 ( .A(B[884]), .B(A[884]), .Z(n262) );
  XOR U263 ( .A(n263), .B(n264), .Z(DIFF[883]) );
  XOR U264 ( .A(B[883]), .B(A[883]), .Z(n264) );
  XOR U265 ( .A(n265), .B(n266), .Z(DIFF[882]) );
  XOR U266 ( .A(B[882]), .B(A[882]), .Z(n266) );
  XOR U267 ( .A(n267), .B(n268), .Z(DIFF[881]) );
  XOR U268 ( .A(B[881]), .B(A[881]), .Z(n268) );
  XOR U269 ( .A(n269), .B(n270), .Z(DIFF[880]) );
  XOR U270 ( .A(B[880]), .B(A[880]), .Z(n270) );
  XOR U271 ( .A(n271), .B(n272), .Z(DIFF[87]) );
  XOR U272 ( .A(B[87]), .B(A[87]), .Z(n272) );
  XOR U273 ( .A(n273), .B(n274), .Z(DIFF[879]) );
  XOR U274 ( .A(B[879]), .B(A[879]), .Z(n274) );
  XOR U275 ( .A(n275), .B(n276), .Z(DIFF[878]) );
  XOR U276 ( .A(B[878]), .B(A[878]), .Z(n276) );
  XOR U277 ( .A(n277), .B(n278), .Z(DIFF[877]) );
  XOR U278 ( .A(B[877]), .B(A[877]), .Z(n278) );
  XOR U279 ( .A(n279), .B(n280), .Z(DIFF[876]) );
  XOR U280 ( .A(B[876]), .B(A[876]), .Z(n280) );
  XOR U281 ( .A(n281), .B(n282), .Z(DIFF[875]) );
  XOR U282 ( .A(B[875]), .B(A[875]), .Z(n282) );
  XOR U283 ( .A(n283), .B(n284), .Z(DIFF[874]) );
  XOR U284 ( .A(B[874]), .B(A[874]), .Z(n284) );
  XOR U285 ( .A(n285), .B(n286), .Z(DIFF[873]) );
  XOR U286 ( .A(B[873]), .B(A[873]), .Z(n286) );
  XOR U287 ( .A(n287), .B(n288), .Z(DIFF[872]) );
  XOR U288 ( .A(B[872]), .B(A[872]), .Z(n288) );
  XOR U289 ( .A(n289), .B(n290), .Z(DIFF[871]) );
  XOR U290 ( .A(B[871]), .B(A[871]), .Z(n290) );
  XOR U291 ( .A(n291), .B(n292), .Z(DIFF[870]) );
  XOR U292 ( .A(B[870]), .B(A[870]), .Z(n292) );
  XOR U293 ( .A(n293), .B(n294), .Z(DIFF[86]) );
  XOR U294 ( .A(B[86]), .B(A[86]), .Z(n294) );
  XOR U295 ( .A(n295), .B(n296), .Z(DIFF[869]) );
  XOR U296 ( .A(B[869]), .B(A[869]), .Z(n296) );
  XOR U297 ( .A(n297), .B(n298), .Z(DIFF[868]) );
  XOR U298 ( .A(B[868]), .B(A[868]), .Z(n298) );
  XOR U299 ( .A(n299), .B(n300), .Z(DIFF[867]) );
  XOR U300 ( .A(B[867]), .B(A[867]), .Z(n300) );
  XOR U301 ( .A(n301), .B(n302), .Z(DIFF[866]) );
  XOR U302 ( .A(B[866]), .B(A[866]), .Z(n302) );
  XOR U303 ( .A(n303), .B(n304), .Z(DIFF[865]) );
  XOR U304 ( .A(B[865]), .B(A[865]), .Z(n304) );
  XOR U305 ( .A(n305), .B(n306), .Z(DIFF[864]) );
  XOR U306 ( .A(B[864]), .B(A[864]), .Z(n306) );
  XOR U307 ( .A(n307), .B(n308), .Z(DIFF[863]) );
  XOR U308 ( .A(B[863]), .B(A[863]), .Z(n308) );
  XOR U309 ( .A(n309), .B(n310), .Z(DIFF[862]) );
  XOR U310 ( .A(B[862]), .B(A[862]), .Z(n310) );
  XOR U311 ( .A(n311), .B(n312), .Z(DIFF[861]) );
  XOR U312 ( .A(B[861]), .B(A[861]), .Z(n312) );
  XOR U313 ( .A(n313), .B(n314), .Z(DIFF[860]) );
  XOR U314 ( .A(B[860]), .B(A[860]), .Z(n314) );
  XOR U315 ( .A(n315), .B(n316), .Z(DIFF[85]) );
  XOR U316 ( .A(B[85]), .B(A[85]), .Z(n316) );
  XOR U317 ( .A(n317), .B(n318), .Z(DIFF[859]) );
  XOR U318 ( .A(B[859]), .B(A[859]), .Z(n318) );
  XOR U319 ( .A(n319), .B(n320), .Z(DIFF[858]) );
  XOR U320 ( .A(B[858]), .B(A[858]), .Z(n320) );
  XOR U321 ( .A(n321), .B(n322), .Z(DIFF[857]) );
  XOR U322 ( .A(B[857]), .B(A[857]), .Z(n322) );
  XOR U323 ( .A(n323), .B(n324), .Z(DIFF[856]) );
  XOR U324 ( .A(B[856]), .B(A[856]), .Z(n324) );
  XOR U325 ( .A(n325), .B(n326), .Z(DIFF[855]) );
  XOR U326 ( .A(B[855]), .B(A[855]), .Z(n326) );
  XOR U327 ( .A(n327), .B(n328), .Z(DIFF[854]) );
  XOR U328 ( .A(B[854]), .B(A[854]), .Z(n328) );
  XOR U329 ( .A(n329), .B(n330), .Z(DIFF[853]) );
  XOR U330 ( .A(B[853]), .B(A[853]), .Z(n330) );
  XOR U331 ( .A(n331), .B(n332), .Z(DIFF[852]) );
  XOR U332 ( .A(B[852]), .B(A[852]), .Z(n332) );
  XOR U333 ( .A(n333), .B(n334), .Z(DIFF[851]) );
  XOR U334 ( .A(B[851]), .B(A[851]), .Z(n334) );
  XOR U335 ( .A(n335), .B(n336), .Z(DIFF[850]) );
  XOR U336 ( .A(B[850]), .B(A[850]), .Z(n336) );
  XOR U337 ( .A(n337), .B(n338), .Z(DIFF[84]) );
  XOR U338 ( .A(B[84]), .B(A[84]), .Z(n338) );
  XOR U339 ( .A(n339), .B(n340), .Z(DIFF[849]) );
  XOR U340 ( .A(B[849]), .B(A[849]), .Z(n340) );
  XOR U341 ( .A(n341), .B(n342), .Z(DIFF[848]) );
  XOR U342 ( .A(B[848]), .B(A[848]), .Z(n342) );
  XOR U343 ( .A(n343), .B(n344), .Z(DIFF[847]) );
  XOR U344 ( .A(B[847]), .B(A[847]), .Z(n344) );
  XOR U345 ( .A(n345), .B(n346), .Z(DIFF[846]) );
  XOR U346 ( .A(B[846]), .B(A[846]), .Z(n346) );
  XOR U347 ( .A(n347), .B(n348), .Z(DIFF[845]) );
  XOR U348 ( .A(B[845]), .B(A[845]), .Z(n348) );
  XOR U349 ( .A(n349), .B(n350), .Z(DIFF[844]) );
  XOR U350 ( .A(B[844]), .B(A[844]), .Z(n350) );
  XOR U351 ( .A(n351), .B(n352), .Z(DIFF[843]) );
  XOR U352 ( .A(B[843]), .B(A[843]), .Z(n352) );
  XOR U353 ( .A(n353), .B(n354), .Z(DIFF[842]) );
  XOR U354 ( .A(B[842]), .B(A[842]), .Z(n354) );
  XOR U355 ( .A(n355), .B(n356), .Z(DIFF[841]) );
  XOR U356 ( .A(B[841]), .B(A[841]), .Z(n356) );
  XOR U357 ( .A(n357), .B(n358), .Z(DIFF[840]) );
  XOR U358 ( .A(B[840]), .B(A[840]), .Z(n358) );
  XOR U359 ( .A(n359), .B(n360), .Z(DIFF[83]) );
  XOR U360 ( .A(B[83]), .B(A[83]), .Z(n360) );
  XOR U361 ( .A(n361), .B(n362), .Z(DIFF[839]) );
  XOR U362 ( .A(B[839]), .B(A[839]), .Z(n362) );
  XOR U363 ( .A(n363), .B(n364), .Z(DIFF[838]) );
  XOR U364 ( .A(B[838]), .B(A[838]), .Z(n364) );
  XOR U365 ( .A(n365), .B(n366), .Z(DIFF[837]) );
  XOR U366 ( .A(B[837]), .B(A[837]), .Z(n366) );
  XOR U367 ( .A(n367), .B(n368), .Z(DIFF[836]) );
  XOR U368 ( .A(B[836]), .B(A[836]), .Z(n368) );
  XOR U369 ( .A(n369), .B(n370), .Z(DIFF[835]) );
  XOR U370 ( .A(B[835]), .B(A[835]), .Z(n370) );
  XOR U371 ( .A(n371), .B(n372), .Z(DIFF[834]) );
  XOR U372 ( .A(B[834]), .B(A[834]), .Z(n372) );
  XOR U373 ( .A(n373), .B(n374), .Z(DIFF[833]) );
  XOR U374 ( .A(B[833]), .B(A[833]), .Z(n374) );
  XOR U375 ( .A(n375), .B(n376), .Z(DIFF[832]) );
  XOR U376 ( .A(B[832]), .B(A[832]), .Z(n376) );
  XOR U377 ( .A(n377), .B(n378), .Z(DIFF[831]) );
  XOR U378 ( .A(B[831]), .B(A[831]), .Z(n378) );
  XOR U379 ( .A(n379), .B(n380), .Z(DIFF[830]) );
  XOR U380 ( .A(B[830]), .B(A[830]), .Z(n380) );
  XOR U381 ( .A(n381), .B(n382), .Z(DIFF[82]) );
  XOR U382 ( .A(B[82]), .B(A[82]), .Z(n382) );
  XOR U383 ( .A(n383), .B(n384), .Z(DIFF[829]) );
  XOR U384 ( .A(B[829]), .B(A[829]), .Z(n384) );
  XOR U385 ( .A(n385), .B(n386), .Z(DIFF[828]) );
  XOR U386 ( .A(B[828]), .B(A[828]), .Z(n386) );
  XOR U387 ( .A(n387), .B(n388), .Z(DIFF[827]) );
  XOR U388 ( .A(B[827]), .B(A[827]), .Z(n388) );
  XOR U389 ( .A(n389), .B(n390), .Z(DIFF[826]) );
  XOR U390 ( .A(B[826]), .B(A[826]), .Z(n390) );
  XOR U391 ( .A(n391), .B(n392), .Z(DIFF[825]) );
  XOR U392 ( .A(B[825]), .B(A[825]), .Z(n392) );
  XOR U393 ( .A(n393), .B(n394), .Z(DIFF[824]) );
  XOR U394 ( .A(B[824]), .B(A[824]), .Z(n394) );
  XOR U395 ( .A(n395), .B(n396), .Z(DIFF[823]) );
  XOR U396 ( .A(B[823]), .B(A[823]), .Z(n396) );
  XOR U397 ( .A(n397), .B(n398), .Z(DIFF[822]) );
  XOR U398 ( .A(B[822]), .B(A[822]), .Z(n398) );
  XOR U399 ( .A(n399), .B(n400), .Z(DIFF[821]) );
  XOR U400 ( .A(B[821]), .B(A[821]), .Z(n400) );
  XOR U401 ( .A(n401), .B(n402), .Z(DIFF[820]) );
  XOR U402 ( .A(B[820]), .B(A[820]), .Z(n402) );
  XOR U403 ( .A(n403), .B(n404), .Z(DIFF[81]) );
  XOR U404 ( .A(B[81]), .B(A[81]), .Z(n404) );
  XOR U405 ( .A(n405), .B(n406), .Z(DIFF[819]) );
  XOR U406 ( .A(B[819]), .B(A[819]), .Z(n406) );
  XOR U407 ( .A(n407), .B(n408), .Z(DIFF[818]) );
  XOR U408 ( .A(B[818]), .B(A[818]), .Z(n408) );
  XOR U409 ( .A(n409), .B(n410), .Z(DIFF[817]) );
  XOR U410 ( .A(B[817]), .B(A[817]), .Z(n410) );
  XOR U411 ( .A(n411), .B(n412), .Z(DIFF[816]) );
  XOR U412 ( .A(B[816]), .B(A[816]), .Z(n412) );
  XOR U413 ( .A(n413), .B(n414), .Z(DIFF[815]) );
  XOR U414 ( .A(B[815]), .B(A[815]), .Z(n414) );
  XOR U415 ( .A(n415), .B(n416), .Z(DIFF[814]) );
  XOR U416 ( .A(B[814]), .B(A[814]), .Z(n416) );
  XOR U417 ( .A(n417), .B(n418), .Z(DIFF[813]) );
  XOR U418 ( .A(B[813]), .B(A[813]), .Z(n418) );
  XOR U419 ( .A(n419), .B(n420), .Z(DIFF[812]) );
  XOR U420 ( .A(B[812]), .B(A[812]), .Z(n420) );
  XOR U421 ( .A(n421), .B(n422), .Z(DIFF[811]) );
  XOR U422 ( .A(B[811]), .B(A[811]), .Z(n422) );
  XOR U423 ( .A(n423), .B(n424), .Z(DIFF[810]) );
  XOR U424 ( .A(B[810]), .B(A[810]), .Z(n424) );
  XOR U425 ( .A(n425), .B(n426), .Z(DIFF[80]) );
  XOR U426 ( .A(B[80]), .B(A[80]), .Z(n426) );
  XOR U427 ( .A(n427), .B(n428), .Z(DIFF[809]) );
  XOR U428 ( .A(B[809]), .B(A[809]), .Z(n428) );
  XOR U429 ( .A(n429), .B(n430), .Z(DIFF[808]) );
  XOR U430 ( .A(B[808]), .B(A[808]), .Z(n430) );
  XOR U431 ( .A(n431), .B(n432), .Z(DIFF[807]) );
  XOR U432 ( .A(B[807]), .B(A[807]), .Z(n432) );
  XOR U433 ( .A(n433), .B(n434), .Z(DIFF[806]) );
  XOR U434 ( .A(B[806]), .B(A[806]), .Z(n434) );
  XOR U435 ( .A(n435), .B(n436), .Z(DIFF[805]) );
  XOR U436 ( .A(B[805]), .B(A[805]), .Z(n436) );
  XOR U437 ( .A(n437), .B(n438), .Z(DIFF[804]) );
  XOR U438 ( .A(B[804]), .B(A[804]), .Z(n438) );
  XOR U439 ( .A(n439), .B(n440), .Z(DIFF[803]) );
  XOR U440 ( .A(B[803]), .B(A[803]), .Z(n440) );
  XOR U441 ( .A(n441), .B(n442), .Z(DIFF[802]) );
  XOR U442 ( .A(B[802]), .B(A[802]), .Z(n442) );
  XOR U443 ( .A(n443), .B(n444), .Z(DIFF[801]) );
  XOR U444 ( .A(B[801]), .B(A[801]), .Z(n444) );
  XOR U445 ( .A(n445), .B(n446), .Z(DIFF[800]) );
  XOR U446 ( .A(B[800]), .B(A[800]), .Z(n446) );
  XOR U447 ( .A(n447), .B(n448), .Z(DIFF[7]) );
  XOR U448 ( .A(B[7]), .B(A[7]), .Z(n448) );
  XOR U449 ( .A(n449), .B(n450), .Z(DIFF[79]) );
  XOR U450 ( .A(B[79]), .B(A[79]), .Z(n450) );
  XOR U451 ( .A(n451), .B(n452), .Z(DIFF[799]) );
  XOR U452 ( .A(B[799]), .B(A[799]), .Z(n452) );
  XOR U453 ( .A(n453), .B(n454), .Z(DIFF[798]) );
  XOR U454 ( .A(B[798]), .B(A[798]), .Z(n454) );
  XOR U455 ( .A(n455), .B(n456), .Z(DIFF[797]) );
  XOR U456 ( .A(B[797]), .B(A[797]), .Z(n456) );
  XOR U457 ( .A(n457), .B(n458), .Z(DIFF[796]) );
  XOR U458 ( .A(B[796]), .B(A[796]), .Z(n458) );
  XOR U459 ( .A(n459), .B(n460), .Z(DIFF[795]) );
  XOR U460 ( .A(B[795]), .B(A[795]), .Z(n460) );
  XOR U461 ( .A(n461), .B(n462), .Z(DIFF[794]) );
  XOR U462 ( .A(B[794]), .B(A[794]), .Z(n462) );
  XOR U463 ( .A(n463), .B(n464), .Z(DIFF[793]) );
  XOR U464 ( .A(B[793]), .B(A[793]), .Z(n464) );
  XOR U465 ( .A(n465), .B(n466), .Z(DIFF[792]) );
  XOR U466 ( .A(B[792]), .B(A[792]), .Z(n466) );
  XOR U467 ( .A(n467), .B(n468), .Z(DIFF[791]) );
  XOR U468 ( .A(B[791]), .B(A[791]), .Z(n468) );
  XOR U469 ( .A(n469), .B(n470), .Z(DIFF[790]) );
  XOR U470 ( .A(B[790]), .B(A[790]), .Z(n470) );
  XOR U471 ( .A(n471), .B(n472), .Z(DIFF[78]) );
  XOR U472 ( .A(B[78]), .B(A[78]), .Z(n472) );
  XOR U473 ( .A(n473), .B(n474), .Z(DIFF[789]) );
  XOR U474 ( .A(B[789]), .B(A[789]), .Z(n474) );
  XOR U475 ( .A(n475), .B(n476), .Z(DIFF[788]) );
  XOR U476 ( .A(B[788]), .B(A[788]), .Z(n476) );
  XOR U477 ( .A(n477), .B(n478), .Z(DIFF[787]) );
  XOR U478 ( .A(B[787]), .B(A[787]), .Z(n478) );
  XOR U479 ( .A(n479), .B(n480), .Z(DIFF[786]) );
  XOR U480 ( .A(B[786]), .B(A[786]), .Z(n480) );
  XOR U481 ( .A(n481), .B(n482), .Z(DIFF[785]) );
  XOR U482 ( .A(B[785]), .B(A[785]), .Z(n482) );
  XOR U483 ( .A(n483), .B(n484), .Z(DIFF[784]) );
  XOR U484 ( .A(B[784]), .B(A[784]), .Z(n484) );
  XOR U485 ( .A(n485), .B(n486), .Z(DIFF[783]) );
  XOR U486 ( .A(B[783]), .B(A[783]), .Z(n486) );
  XOR U487 ( .A(n487), .B(n488), .Z(DIFF[782]) );
  XOR U488 ( .A(B[782]), .B(A[782]), .Z(n488) );
  XOR U489 ( .A(n489), .B(n490), .Z(DIFF[781]) );
  XOR U490 ( .A(B[781]), .B(A[781]), .Z(n490) );
  XOR U491 ( .A(n491), .B(n492), .Z(DIFF[780]) );
  XOR U492 ( .A(B[780]), .B(A[780]), .Z(n492) );
  XOR U493 ( .A(n493), .B(n494), .Z(DIFF[77]) );
  XOR U494 ( .A(B[77]), .B(A[77]), .Z(n494) );
  XOR U495 ( .A(n495), .B(n496), .Z(DIFF[779]) );
  XOR U496 ( .A(B[779]), .B(A[779]), .Z(n496) );
  XOR U497 ( .A(n497), .B(n498), .Z(DIFF[778]) );
  XOR U498 ( .A(B[778]), .B(A[778]), .Z(n498) );
  XOR U499 ( .A(n499), .B(n500), .Z(DIFF[777]) );
  XOR U500 ( .A(B[777]), .B(A[777]), .Z(n500) );
  XOR U501 ( .A(n501), .B(n502), .Z(DIFF[776]) );
  XOR U502 ( .A(B[776]), .B(A[776]), .Z(n502) );
  XOR U503 ( .A(n503), .B(n504), .Z(DIFF[775]) );
  XOR U504 ( .A(B[775]), .B(A[775]), .Z(n504) );
  XOR U505 ( .A(n505), .B(n506), .Z(DIFF[774]) );
  XOR U506 ( .A(B[774]), .B(A[774]), .Z(n506) );
  XOR U507 ( .A(n507), .B(n508), .Z(DIFF[773]) );
  XOR U508 ( .A(B[773]), .B(A[773]), .Z(n508) );
  XOR U509 ( .A(n509), .B(n510), .Z(DIFF[772]) );
  XOR U510 ( .A(B[772]), .B(A[772]), .Z(n510) );
  XOR U511 ( .A(n511), .B(n512), .Z(DIFF[771]) );
  XOR U512 ( .A(B[771]), .B(A[771]), .Z(n512) );
  XOR U513 ( .A(n513), .B(n514), .Z(DIFF[770]) );
  XOR U514 ( .A(B[770]), .B(A[770]), .Z(n514) );
  XOR U515 ( .A(n515), .B(n516), .Z(DIFF[76]) );
  XOR U516 ( .A(B[76]), .B(A[76]), .Z(n516) );
  XOR U517 ( .A(n517), .B(n518), .Z(DIFF[769]) );
  XOR U518 ( .A(B[769]), .B(A[769]), .Z(n518) );
  XOR U519 ( .A(n519), .B(n520), .Z(DIFF[768]) );
  XOR U520 ( .A(B[768]), .B(A[768]), .Z(n520) );
  XOR U521 ( .A(n521), .B(n522), .Z(DIFF[767]) );
  XOR U522 ( .A(B[767]), .B(A[767]), .Z(n522) );
  XOR U523 ( .A(n523), .B(n524), .Z(DIFF[766]) );
  XOR U524 ( .A(B[766]), .B(A[766]), .Z(n524) );
  XOR U525 ( .A(n525), .B(n526), .Z(DIFF[765]) );
  XOR U526 ( .A(B[765]), .B(A[765]), .Z(n526) );
  XOR U527 ( .A(n527), .B(n528), .Z(DIFF[764]) );
  XOR U528 ( .A(B[764]), .B(A[764]), .Z(n528) );
  XOR U529 ( .A(n529), .B(n530), .Z(DIFF[763]) );
  XOR U530 ( .A(B[763]), .B(A[763]), .Z(n530) );
  XOR U531 ( .A(n531), .B(n532), .Z(DIFF[762]) );
  XOR U532 ( .A(B[762]), .B(A[762]), .Z(n532) );
  XOR U533 ( .A(n533), .B(n534), .Z(DIFF[761]) );
  XOR U534 ( .A(B[761]), .B(A[761]), .Z(n534) );
  XOR U535 ( .A(n535), .B(n536), .Z(DIFF[760]) );
  XOR U536 ( .A(B[760]), .B(A[760]), .Z(n536) );
  XOR U537 ( .A(n537), .B(n538), .Z(DIFF[75]) );
  XOR U538 ( .A(B[75]), .B(A[75]), .Z(n538) );
  XOR U539 ( .A(n539), .B(n540), .Z(DIFF[759]) );
  XOR U540 ( .A(B[759]), .B(A[759]), .Z(n540) );
  XOR U541 ( .A(n541), .B(n542), .Z(DIFF[758]) );
  XOR U542 ( .A(B[758]), .B(A[758]), .Z(n542) );
  XOR U543 ( .A(n543), .B(n544), .Z(DIFF[757]) );
  XOR U544 ( .A(B[757]), .B(A[757]), .Z(n544) );
  XOR U545 ( .A(n545), .B(n546), .Z(DIFF[756]) );
  XOR U546 ( .A(B[756]), .B(A[756]), .Z(n546) );
  XOR U547 ( .A(n547), .B(n548), .Z(DIFF[755]) );
  XOR U548 ( .A(B[755]), .B(A[755]), .Z(n548) );
  XOR U549 ( .A(n549), .B(n550), .Z(DIFF[754]) );
  XOR U550 ( .A(B[754]), .B(A[754]), .Z(n550) );
  XOR U551 ( .A(n551), .B(n552), .Z(DIFF[753]) );
  XOR U552 ( .A(B[753]), .B(A[753]), .Z(n552) );
  XOR U553 ( .A(n553), .B(n554), .Z(DIFF[752]) );
  XOR U554 ( .A(B[752]), .B(A[752]), .Z(n554) );
  XOR U555 ( .A(n555), .B(n556), .Z(DIFF[751]) );
  XOR U556 ( .A(B[751]), .B(A[751]), .Z(n556) );
  XOR U557 ( .A(n557), .B(n558), .Z(DIFF[750]) );
  XOR U558 ( .A(B[750]), .B(A[750]), .Z(n558) );
  XOR U559 ( .A(n559), .B(n560), .Z(DIFF[74]) );
  XOR U560 ( .A(B[74]), .B(A[74]), .Z(n560) );
  XOR U561 ( .A(n561), .B(n562), .Z(DIFF[749]) );
  XOR U562 ( .A(B[749]), .B(A[749]), .Z(n562) );
  XOR U563 ( .A(n563), .B(n564), .Z(DIFF[748]) );
  XOR U564 ( .A(B[748]), .B(A[748]), .Z(n564) );
  XOR U565 ( .A(n565), .B(n566), .Z(DIFF[747]) );
  XOR U566 ( .A(B[747]), .B(A[747]), .Z(n566) );
  XOR U567 ( .A(n567), .B(n568), .Z(DIFF[746]) );
  XOR U568 ( .A(B[746]), .B(A[746]), .Z(n568) );
  XOR U569 ( .A(n569), .B(n570), .Z(DIFF[745]) );
  XOR U570 ( .A(B[745]), .B(A[745]), .Z(n570) );
  XOR U571 ( .A(n571), .B(n572), .Z(DIFF[744]) );
  XOR U572 ( .A(B[744]), .B(A[744]), .Z(n572) );
  XOR U573 ( .A(n573), .B(n574), .Z(DIFF[743]) );
  XOR U574 ( .A(B[743]), .B(A[743]), .Z(n574) );
  XOR U575 ( .A(n575), .B(n576), .Z(DIFF[742]) );
  XOR U576 ( .A(B[742]), .B(A[742]), .Z(n576) );
  XOR U577 ( .A(n577), .B(n578), .Z(DIFF[741]) );
  XOR U578 ( .A(B[741]), .B(A[741]), .Z(n578) );
  XOR U579 ( .A(n579), .B(n580), .Z(DIFF[740]) );
  XOR U580 ( .A(B[740]), .B(A[740]), .Z(n580) );
  XOR U581 ( .A(n581), .B(n582), .Z(DIFF[73]) );
  XOR U582 ( .A(B[73]), .B(A[73]), .Z(n582) );
  XOR U583 ( .A(n583), .B(n584), .Z(DIFF[739]) );
  XOR U584 ( .A(B[739]), .B(A[739]), .Z(n584) );
  XOR U585 ( .A(n585), .B(n586), .Z(DIFF[738]) );
  XOR U586 ( .A(B[738]), .B(A[738]), .Z(n586) );
  XOR U587 ( .A(n587), .B(n588), .Z(DIFF[737]) );
  XOR U588 ( .A(B[737]), .B(A[737]), .Z(n588) );
  XOR U589 ( .A(n589), .B(n590), .Z(DIFF[736]) );
  XOR U590 ( .A(B[736]), .B(A[736]), .Z(n590) );
  XOR U591 ( .A(n591), .B(n592), .Z(DIFF[735]) );
  XOR U592 ( .A(B[735]), .B(A[735]), .Z(n592) );
  XOR U593 ( .A(n593), .B(n594), .Z(DIFF[734]) );
  XOR U594 ( .A(B[734]), .B(A[734]), .Z(n594) );
  XOR U595 ( .A(n595), .B(n596), .Z(DIFF[733]) );
  XOR U596 ( .A(B[733]), .B(A[733]), .Z(n596) );
  XOR U597 ( .A(n597), .B(n598), .Z(DIFF[732]) );
  XOR U598 ( .A(B[732]), .B(A[732]), .Z(n598) );
  XOR U599 ( .A(n599), .B(n600), .Z(DIFF[731]) );
  XOR U600 ( .A(B[731]), .B(A[731]), .Z(n600) );
  XOR U601 ( .A(n601), .B(n602), .Z(DIFF[730]) );
  XOR U602 ( .A(B[730]), .B(A[730]), .Z(n602) );
  XOR U603 ( .A(n603), .B(n604), .Z(DIFF[72]) );
  XOR U604 ( .A(B[72]), .B(A[72]), .Z(n604) );
  XOR U605 ( .A(n605), .B(n606), .Z(DIFF[729]) );
  XOR U606 ( .A(B[729]), .B(A[729]), .Z(n606) );
  XOR U607 ( .A(n607), .B(n608), .Z(DIFF[728]) );
  XOR U608 ( .A(B[728]), .B(A[728]), .Z(n608) );
  XOR U609 ( .A(n609), .B(n610), .Z(DIFF[727]) );
  XOR U610 ( .A(B[727]), .B(A[727]), .Z(n610) );
  XOR U611 ( .A(n611), .B(n612), .Z(DIFF[726]) );
  XOR U612 ( .A(B[726]), .B(A[726]), .Z(n612) );
  XOR U613 ( .A(n613), .B(n614), .Z(DIFF[725]) );
  XOR U614 ( .A(B[725]), .B(A[725]), .Z(n614) );
  XOR U615 ( .A(n615), .B(n616), .Z(DIFF[724]) );
  XOR U616 ( .A(B[724]), .B(A[724]), .Z(n616) );
  XOR U617 ( .A(n617), .B(n618), .Z(DIFF[723]) );
  XOR U618 ( .A(B[723]), .B(A[723]), .Z(n618) );
  XOR U619 ( .A(n619), .B(n620), .Z(DIFF[722]) );
  XOR U620 ( .A(B[722]), .B(A[722]), .Z(n620) );
  XOR U621 ( .A(n621), .B(n622), .Z(DIFF[721]) );
  XOR U622 ( .A(B[721]), .B(A[721]), .Z(n622) );
  XOR U623 ( .A(n623), .B(n624), .Z(DIFF[720]) );
  XOR U624 ( .A(B[720]), .B(A[720]), .Z(n624) );
  XOR U625 ( .A(n625), .B(n626), .Z(DIFF[71]) );
  XOR U626 ( .A(B[71]), .B(A[71]), .Z(n626) );
  XOR U627 ( .A(n627), .B(n628), .Z(DIFF[719]) );
  XOR U628 ( .A(B[719]), .B(A[719]), .Z(n628) );
  XOR U629 ( .A(n629), .B(n630), .Z(DIFF[718]) );
  XOR U630 ( .A(B[718]), .B(A[718]), .Z(n630) );
  XOR U631 ( .A(n631), .B(n632), .Z(DIFF[717]) );
  XOR U632 ( .A(B[717]), .B(A[717]), .Z(n632) );
  XOR U633 ( .A(n633), .B(n634), .Z(DIFF[716]) );
  XOR U634 ( .A(B[716]), .B(A[716]), .Z(n634) );
  XOR U635 ( .A(n635), .B(n636), .Z(DIFF[715]) );
  XOR U636 ( .A(B[715]), .B(A[715]), .Z(n636) );
  XOR U637 ( .A(n637), .B(n638), .Z(DIFF[714]) );
  XOR U638 ( .A(B[714]), .B(A[714]), .Z(n638) );
  XOR U639 ( .A(n639), .B(n640), .Z(DIFF[713]) );
  XOR U640 ( .A(B[713]), .B(A[713]), .Z(n640) );
  XOR U641 ( .A(n641), .B(n642), .Z(DIFF[712]) );
  XOR U642 ( .A(B[712]), .B(A[712]), .Z(n642) );
  XOR U643 ( .A(n643), .B(n644), .Z(DIFF[711]) );
  XOR U644 ( .A(B[711]), .B(A[711]), .Z(n644) );
  XOR U645 ( .A(n645), .B(n646), .Z(DIFF[710]) );
  XOR U646 ( .A(B[710]), .B(A[710]), .Z(n646) );
  XOR U647 ( .A(n647), .B(n648), .Z(DIFF[70]) );
  XOR U648 ( .A(B[70]), .B(A[70]), .Z(n648) );
  XOR U649 ( .A(n649), .B(n650), .Z(DIFF[709]) );
  XOR U650 ( .A(B[709]), .B(A[709]), .Z(n650) );
  XOR U651 ( .A(n651), .B(n652), .Z(DIFF[708]) );
  XOR U652 ( .A(B[708]), .B(A[708]), .Z(n652) );
  XOR U653 ( .A(n653), .B(n654), .Z(DIFF[707]) );
  XOR U654 ( .A(B[707]), .B(A[707]), .Z(n654) );
  XOR U655 ( .A(n655), .B(n656), .Z(DIFF[706]) );
  XOR U656 ( .A(B[706]), .B(A[706]), .Z(n656) );
  XOR U657 ( .A(n657), .B(n658), .Z(DIFF[705]) );
  XOR U658 ( .A(B[705]), .B(A[705]), .Z(n658) );
  XOR U659 ( .A(n659), .B(n660), .Z(DIFF[704]) );
  XOR U660 ( .A(B[704]), .B(A[704]), .Z(n660) );
  XOR U661 ( .A(n661), .B(n662), .Z(DIFF[703]) );
  XOR U662 ( .A(B[703]), .B(A[703]), .Z(n662) );
  XOR U663 ( .A(n663), .B(n664), .Z(DIFF[702]) );
  XOR U664 ( .A(B[702]), .B(A[702]), .Z(n664) );
  XOR U665 ( .A(n665), .B(n666), .Z(DIFF[701]) );
  XOR U666 ( .A(B[701]), .B(A[701]), .Z(n666) );
  XOR U667 ( .A(n667), .B(n668), .Z(DIFF[700]) );
  XOR U668 ( .A(B[700]), .B(A[700]), .Z(n668) );
  XOR U669 ( .A(n669), .B(n670), .Z(DIFF[6]) );
  XOR U670 ( .A(B[6]), .B(A[6]), .Z(n670) );
  XOR U671 ( .A(n671), .B(n672), .Z(DIFF[69]) );
  XOR U672 ( .A(B[69]), .B(A[69]), .Z(n672) );
  XOR U673 ( .A(n673), .B(n674), .Z(DIFF[699]) );
  XOR U674 ( .A(B[699]), .B(A[699]), .Z(n674) );
  XOR U675 ( .A(n675), .B(n676), .Z(DIFF[698]) );
  XOR U676 ( .A(B[698]), .B(A[698]), .Z(n676) );
  XOR U677 ( .A(n677), .B(n678), .Z(DIFF[697]) );
  XOR U678 ( .A(B[697]), .B(A[697]), .Z(n678) );
  XOR U679 ( .A(n679), .B(n680), .Z(DIFF[696]) );
  XOR U680 ( .A(B[696]), .B(A[696]), .Z(n680) );
  XOR U681 ( .A(n681), .B(n682), .Z(DIFF[695]) );
  XOR U682 ( .A(B[695]), .B(A[695]), .Z(n682) );
  XOR U683 ( .A(n683), .B(n684), .Z(DIFF[694]) );
  XOR U684 ( .A(B[694]), .B(A[694]), .Z(n684) );
  XOR U685 ( .A(n685), .B(n686), .Z(DIFF[693]) );
  XOR U686 ( .A(B[693]), .B(A[693]), .Z(n686) );
  XOR U687 ( .A(n687), .B(n688), .Z(DIFF[692]) );
  XOR U688 ( .A(B[692]), .B(A[692]), .Z(n688) );
  XOR U689 ( .A(n689), .B(n690), .Z(DIFF[691]) );
  XOR U690 ( .A(B[691]), .B(A[691]), .Z(n690) );
  XOR U691 ( .A(n691), .B(n692), .Z(DIFF[690]) );
  XOR U692 ( .A(B[690]), .B(A[690]), .Z(n692) );
  XOR U693 ( .A(n693), .B(n694), .Z(DIFF[68]) );
  XOR U694 ( .A(B[68]), .B(A[68]), .Z(n694) );
  XOR U695 ( .A(n695), .B(n696), .Z(DIFF[689]) );
  XOR U696 ( .A(B[689]), .B(A[689]), .Z(n696) );
  XOR U697 ( .A(n697), .B(n698), .Z(DIFF[688]) );
  XOR U698 ( .A(B[688]), .B(A[688]), .Z(n698) );
  XOR U699 ( .A(n699), .B(n700), .Z(DIFF[687]) );
  XOR U700 ( .A(B[687]), .B(A[687]), .Z(n700) );
  XOR U701 ( .A(n701), .B(n702), .Z(DIFF[686]) );
  XOR U702 ( .A(B[686]), .B(A[686]), .Z(n702) );
  XOR U703 ( .A(n703), .B(n704), .Z(DIFF[685]) );
  XOR U704 ( .A(B[685]), .B(A[685]), .Z(n704) );
  XOR U705 ( .A(n705), .B(n706), .Z(DIFF[684]) );
  XOR U706 ( .A(B[684]), .B(A[684]), .Z(n706) );
  XOR U707 ( .A(n707), .B(n708), .Z(DIFF[683]) );
  XOR U708 ( .A(B[683]), .B(A[683]), .Z(n708) );
  XOR U709 ( .A(n709), .B(n710), .Z(DIFF[682]) );
  XOR U710 ( .A(B[682]), .B(A[682]), .Z(n710) );
  XOR U711 ( .A(n711), .B(n712), .Z(DIFF[681]) );
  XOR U712 ( .A(B[681]), .B(A[681]), .Z(n712) );
  XOR U713 ( .A(n713), .B(n714), .Z(DIFF[680]) );
  XOR U714 ( .A(B[680]), .B(A[680]), .Z(n714) );
  XOR U715 ( .A(n715), .B(n716), .Z(DIFF[67]) );
  XOR U716 ( .A(B[67]), .B(A[67]), .Z(n716) );
  XOR U717 ( .A(n717), .B(n718), .Z(DIFF[679]) );
  XOR U718 ( .A(B[679]), .B(A[679]), .Z(n718) );
  XOR U719 ( .A(n719), .B(n720), .Z(DIFF[678]) );
  XOR U720 ( .A(B[678]), .B(A[678]), .Z(n720) );
  XOR U721 ( .A(n721), .B(n722), .Z(DIFF[677]) );
  XOR U722 ( .A(B[677]), .B(A[677]), .Z(n722) );
  XOR U723 ( .A(n723), .B(n724), .Z(DIFF[676]) );
  XOR U724 ( .A(B[676]), .B(A[676]), .Z(n724) );
  XOR U725 ( .A(n725), .B(n726), .Z(DIFF[675]) );
  XOR U726 ( .A(B[675]), .B(A[675]), .Z(n726) );
  XOR U727 ( .A(n727), .B(n728), .Z(DIFF[674]) );
  XOR U728 ( .A(B[674]), .B(A[674]), .Z(n728) );
  XOR U729 ( .A(n729), .B(n730), .Z(DIFF[673]) );
  XOR U730 ( .A(B[673]), .B(A[673]), .Z(n730) );
  XOR U731 ( .A(n731), .B(n732), .Z(DIFF[672]) );
  XOR U732 ( .A(B[672]), .B(A[672]), .Z(n732) );
  XOR U733 ( .A(n733), .B(n734), .Z(DIFF[671]) );
  XOR U734 ( .A(B[671]), .B(A[671]), .Z(n734) );
  XOR U735 ( .A(n735), .B(n736), .Z(DIFF[670]) );
  XOR U736 ( .A(B[670]), .B(A[670]), .Z(n736) );
  XOR U737 ( .A(n737), .B(n738), .Z(DIFF[66]) );
  XOR U738 ( .A(B[66]), .B(A[66]), .Z(n738) );
  XOR U739 ( .A(n739), .B(n740), .Z(DIFF[669]) );
  XOR U740 ( .A(B[669]), .B(A[669]), .Z(n740) );
  XOR U741 ( .A(n741), .B(n742), .Z(DIFF[668]) );
  XOR U742 ( .A(B[668]), .B(A[668]), .Z(n742) );
  XOR U743 ( .A(n743), .B(n744), .Z(DIFF[667]) );
  XOR U744 ( .A(B[667]), .B(A[667]), .Z(n744) );
  XOR U745 ( .A(n745), .B(n746), .Z(DIFF[666]) );
  XOR U746 ( .A(B[666]), .B(A[666]), .Z(n746) );
  XOR U747 ( .A(n747), .B(n748), .Z(DIFF[665]) );
  XOR U748 ( .A(B[665]), .B(A[665]), .Z(n748) );
  XOR U749 ( .A(n749), .B(n750), .Z(DIFF[664]) );
  XOR U750 ( .A(B[664]), .B(A[664]), .Z(n750) );
  XOR U751 ( .A(n751), .B(n752), .Z(DIFF[663]) );
  XOR U752 ( .A(B[663]), .B(A[663]), .Z(n752) );
  XOR U753 ( .A(n753), .B(n754), .Z(DIFF[662]) );
  XOR U754 ( .A(B[662]), .B(A[662]), .Z(n754) );
  XOR U755 ( .A(n755), .B(n756), .Z(DIFF[661]) );
  XOR U756 ( .A(B[661]), .B(A[661]), .Z(n756) );
  XOR U757 ( .A(n757), .B(n758), .Z(DIFF[660]) );
  XOR U758 ( .A(B[660]), .B(A[660]), .Z(n758) );
  XOR U759 ( .A(n759), .B(n760), .Z(DIFF[65]) );
  XOR U760 ( .A(B[65]), .B(A[65]), .Z(n760) );
  XOR U761 ( .A(n761), .B(n762), .Z(DIFF[659]) );
  XOR U762 ( .A(B[659]), .B(A[659]), .Z(n762) );
  XOR U763 ( .A(n763), .B(n764), .Z(DIFF[658]) );
  XOR U764 ( .A(B[658]), .B(A[658]), .Z(n764) );
  XOR U765 ( .A(n765), .B(n766), .Z(DIFF[657]) );
  XOR U766 ( .A(B[657]), .B(A[657]), .Z(n766) );
  XOR U767 ( .A(n767), .B(n768), .Z(DIFF[656]) );
  XOR U768 ( .A(B[656]), .B(A[656]), .Z(n768) );
  XOR U769 ( .A(n769), .B(n770), .Z(DIFF[655]) );
  XOR U770 ( .A(B[655]), .B(A[655]), .Z(n770) );
  XOR U771 ( .A(n771), .B(n772), .Z(DIFF[654]) );
  XOR U772 ( .A(B[654]), .B(A[654]), .Z(n772) );
  XOR U773 ( .A(n773), .B(n774), .Z(DIFF[653]) );
  XOR U774 ( .A(B[653]), .B(A[653]), .Z(n774) );
  XOR U775 ( .A(n775), .B(n776), .Z(DIFF[652]) );
  XOR U776 ( .A(B[652]), .B(A[652]), .Z(n776) );
  XOR U777 ( .A(n777), .B(n778), .Z(DIFF[651]) );
  XOR U778 ( .A(B[651]), .B(A[651]), .Z(n778) );
  XOR U779 ( .A(n779), .B(n780), .Z(DIFF[650]) );
  XOR U780 ( .A(B[650]), .B(A[650]), .Z(n780) );
  XOR U781 ( .A(n781), .B(n782), .Z(DIFF[64]) );
  XOR U782 ( .A(B[64]), .B(A[64]), .Z(n782) );
  XOR U783 ( .A(n783), .B(n784), .Z(DIFF[649]) );
  XOR U784 ( .A(B[649]), .B(A[649]), .Z(n784) );
  XOR U785 ( .A(n785), .B(n786), .Z(DIFF[648]) );
  XOR U786 ( .A(B[648]), .B(A[648]), .Z(n786) );
  XOR U787 ( .A(n787), .B(n788), .Z(DIFF[647]) );
  XOR U788 ( .A(B[647]), .B(A[647]), .Z(n788) );
  XOR U789 ( .A(n789), .B(n790), .Z(DIFF[646]) );
  XOR U790 ( .A(B[646]), .B(A[646]), .Z(n790) );
  XOR U791 ( .A(n791), .B(n792), .Z(DIFF[645]) );
  XOR U792 ( .A(B[645]), .B(A[645]), .Z(n792) );
  XOR U793 ( .A(n793), .B(n794), .Z(DIFF[644]) );
  XOR U794 ( .A(B[644]), .B(A[644]), .Z(n794) );
  XOR U795 ( .A(n795), .B(n796), .Z(DIFF[643]) );
  XOR U796 ( .A(B[643]), .B(A[643]), .Z(n796) );
  XOR U797 ( .A(n797), .B(n798), .Z(DIFF[642]) );
  XOR U798 ( .A(B[642]), .B(A[642]), .Z(n798) );
  XOR U799 ( .A(n799), .B(n800), .Z(DIFF[641]) );
  XOR U800 ( .A(B[641]), .B(A[641]), .Z(n800) );
  XOR U801 ( .A(n801), .B(n802), .Z(DIFF[640]) );
  XOR U802 ( .A(B[640]), .B(A[640]), .Z(n802) );
  XOR U803 ( .A(n803), .B(n804), .Z(DIFF[63]) );
  XOR U804 ( .A(B[63]), .B(A[63]), .Z(n804) );
  XOR U805 ( .A(n805), .B(n806), .Z(DIFF[639]) );
  XOR U806 ( .A(B[639]), .B(A[639]), .Z(n806) );
  XOR U807 ( .A(n807), .B(n808), .Z(DIFF[638]) );
  XOR U808 ( .A(B[638]), .B(A[638]), .Z(n808) );
  XOR U809 ( .A(n809), .B(n810), .Z(DIFF[637]) );
  XOR U810 ( .A(B[637]), .B(A[637]), .Z(n810) );
  XOR U811 ( .A(n811), .B(n812), .Z(DIFF[636]) );
  XOR U812 ( .A(B[636]), .B(A[636]), .Z(n812) );
  XOR U813 ( .A(n813), .B(n814), .Z(DIFF[635]) );
  XOR U814 ( .A(B[635]), .B(A[635]), .Z(n814) );
  XOR U815 ( .A(n815), .B(n816), .Z(DIFF[634]) );
  XOR U816 ( .A(B[634]), .B(A[634]), .Z(n816) );
  XOR U817 ( .A(n817), .B(n818), .Z(DIFF[633]) );
  XOR U818 ( .A(B[633]), .B(A[633]), .Z(n818) );
  XOR U819 ( .A(n819), .B(n820), .Z(DIFF[632]) );
  XOR U820 ( .A(B[632]), .B(A[632]), .Z(n820) );
  XOR U821 ( .A(n821), .B(n822), .Z(DIFF[631]) );
  XOR U822 ( .A(B[631]), .B(A[631]), .Z(n822) );
  XOR U823 ( .A(n823), .B(n824), .Z(DIFF[630]) );
  XOR U824 ( .A(B[630]), .B(A[630]), .Z(n824) );
  XOR U825 ( .A(n825), .B(n826), .Z(DIFF[62]) );
  XOR U826 ( .A(B[62]), .B(A[62]), .Z(n826) );
  XOR U827 ( .A(n827), .B(n828), .Z(DIFF[629]) );
  XOR U828 ( .A(B[629]), .B(A[629]), .Z(n828) );
  XOR U829 ( .A(n829), .B(n830), .Z(DIFF[628]) );
  XOR U830 ( .A(B[628]), .B(A[628]), .Z(n830) );
  XOR U831 ( .A(n831), .B(n832), .Z(DIFF[627]) );
  XOR U832 ( .A(B[627]), .B(A[627]), .Z(n832) );
  XOR U833 ( .A(n833), .B(n834), .Z(DIFF[626]) );
  XOR U834 ( .A(B[626]), .B(A[626]), .Z(n834) );
  XOR U835 ( .A(n835), .B(n836), .Z(DIFF[625]) );
  XOR U836 ( .A(B[625]), .B(A[625]), .Z(n836) );
  XOR U837 ( .A(n837), .B(n838), .Z(DIFF[624]) );
  XOR U838 ( .A(B[624]), .B(A[624]), .Z(n838) );
  XOR U839 ( .A(n839), .B(n840), .Z(DIFF[623]) );
  XOR U840 ( .A(B[623]), .B(A[623]), .Z(n840) );
  XOR U841 ( .A(n841), .B(n842), .Z(DIFF[622]) );
  XOR U842 ( .A(B[622]), .B(A[622]), .Z(n842) );
  XOR U843 ( .A(n843), .B(n844), .Z(DIFF[621]) );
  XOR U844 ( .A(B[621]), .B(A[621]), .Z(n844) );
  XOR U845 ( .A(n845), .B(n846), .Z(DIFF[620]) );
  XOR U846 ( .A(B[620]), .B(A[620]), .Z(n846) );
  XOR U847 ( .A(n847), .B(n848), .Z(DIFF[61]) );
  XOR U848 ( .A(B[61]), .B(A[61]), .Z(n848) );
  XOR U849 ( .A(n849), .B(n850), .Z(DIFF[619]) );
  XOR U850 ( .A(B[619]), .B(A[619]), .Z(n850) );
  XOR U851 ( .A(n851), .B(n852), .Z(DIFF[618]) );
  XOR U852 ( .A(B[618]), .B(A[618]), .Z(n852) );
  XOR U853 ( .A(n853), .B(n854), .Z(DIFF[617]) );
  XOR U854 ( .A(B[617]), .B(A[617]), .Z(n854) );
  XOR U855 ( .A(n855), .B(n856), .Z(DIFF[616]) );
  XOR U856 ( .A(B[616]), .B(A[616]), .Z(n856) );
  XOR U857 ( .A(n857), .B(n858), .Z(DIFF[615]) );
  XOR U858 ( .A(B[615]), .B(A[615]), .Z(n858) );
  XOR U859 ( .A(n859), .B(n860), .Z(DIFF[614]) );
  XOR U860 ( .A(B[614]), .B(A[614]), .Z(n860) );
  XOR U861 ( .A(n861), .B(n862), .Z(DIFF[613]) );
  XOR U862 ( .A(B[613]), .B(A[613]), .Z(n862) );
  XOR U863 ( .A(n863), .B(n864), .Z(DIFF[612]) );
  XOR U864 ( .A(B[612]), .B(A[612]), .Z(n864) );
  XOR U865 ( .A(n865), .B(n866), .Z(DIFF[611]) );
  XOR U866 ( .A(B[611]), .B(A[611]), .Z(n866) );
  XOR U867 ( .A(n867), .B(n868), .Z(DIFF[610]) );
  XOR U868 ( .A(B[610]), .B(A[610]), .Z(n868) );
  XOR U869 ( .A(n869), .B(n870), .Z(DIFF[60]) );
  XOR U870 ( .A(B[60]), .B(A[60]), .Z(n870) );
  XOR U871 ( .A(n871), .B(n872), .Z(DIFF[609]) );
  XOR U872 ( .A(B[609]), .B(A[609]), .Z(n872) );
  XOR U873 ( .A(n873), .B(n874), .Z(DIFF[608]) );
  XOR U874 ( .A(B[608]), .B(A[608]), .Z(n874) );
  XOR U875 ( .A(n875), .B(n876), .Z(DIFF[607]) );
  XOR U876 ( .A(B[607]), .B(A[607]), .Z(n876) );
  XOR U877 ( .A(n877), .B(n878), .Z(DIFF[606]) );
  XOR U878 ( .A(B[606]), .B(A[606]), .Z(n878) );
  XOR U879 ( .A(n879), .B(n880), .Z(DIFF[605]) );
  XOR U880 ( .A(B[605]), .B(A[605]), .Z(n880) );
  XOR U881 ( .A(n881), .B(n882), .Z(DIFF[604]) );
  XOR U882 ( .A(B[604]), .B(A[604]), .Z(n882) );
  XOR U883 ( .A(n883), .B(n884), .Z(DIFF[603]) );
  XOR U884 ( .A(B[603]), .B(A[603]), .Z(n884) );
  XOR U885 ( .A(n885), .B(n886), .Z(DIFF[602]) );
  XOR U886 ( .A(B[602]), .B(A[602]), .Z(n886) );
  XOR U887 ( .A(n887), .B(n888), .Z(DIFF[601]) );
  XOR U888 ( .A(B[601]), .B(A[601]), .Z(n888) );
  XOR U889 ( .A(n889), .B(n890), .Z(DIFF[600]) );
  XOR U890 ( .A(B[600]), .B(A[600]), .Z(n890) );
  XOR U891 ( .A(n891), .B(n892), .Z(DIFF[5]) );
  XOR U892 ( .A(B[5]), .B(A[5]), .Z(n892) );
  XOR U893 ( .A(n893), .B(n894), .Z(DIFF[59]) );
  XOR U894 ( .A(B[59]), .B(A[59]), .Z(n894) );
  XOR U895 ( .A(n895), .B(n896), .Z(DIFF[599]) );
  XOR U896 ( .A(B[599]), .B(A[599]), .Z(n896) );
  XOR U897 ( .A(n897), .B(n898), .Z(DIFF[598]) );
  XOR U898 ( .A(B[598]), .B(A[598]), .Z(n898) );
  XOR U899 ( .A(n899), .B(n900), .Z(DIFF[597]) );
  XOR U900 ( .A(B[597]), .B(A[597]), .Z(n900) );
  XOR U901 ( .A(n901), .B(n902), .Z(DIFF[596]) );
  XOR U902 ( .A(B[596]), .B(A[596]), .Z(n902) );
  XOR U903 ( .A(n903), .B(n904), .Z(DIFF[595]) );
  XOR U904 ( .A(B[595]), .B(A[595]), .Z(n904) );
  XOR U905 ( .A(n905), .B(n906), .Z(DIFF[594]) );
  XOR U906 ( .A(B[594]), .B(A[594]), .Z(n906) );
  XOR U907 ( .A(n907), .B(n908), .Z(DIFF[593]) );
  XOR U908 ( .A(B[593]), .B(A[593]), .Z(n908) );
  XOR U909 ( .A(n909), .B(n910), .Z(DIFF[592]) );
  XOR U910 ( .A(B[592]), .B(A[592]), .Z(n910) );
  XOR U911 ( .A(n911), .B(n912), .Z(DIFF[591]) );
  XOR U912 ( .A(B[591]), .B(A[591]), .Z(n912) );
  XOR U913 ( .A(n913), .B(n914), .Z(DIFF[590]) );
  XOR U914 ( .A(B[590]), .B(A[590]), .Z(n914) );
  XOR U915 ( .A(n915), .B(n916), .Z(DIFF[58]) );
  XOR U916 ( .A(B[58]), .B(A[58]), .Z(n916) );
  XOR U917 ( .A(n917), .B(n918), .Z(DIFF[589]) );
  XOR U918 ( .A(B[589]), .B(A[589]), .Z(n918) );
  XOR U919 ( .A(n919), .B(n920), .Z(DIFF[588]) );
  XOR U920 ( .A(B[588]), .B(A[588]), .Z(n920) );
  XOR U921 ( .A(n921), .B(n922), .Z(DIFF[587]) );
  XOR U922 ( .A(B[587]), .B(A[587]), .Z(n922) );
  XOR U923 ( .A(n923), .B(n924), .Z(DIFF[586]) );
  XOR U924 ( .A(B[586]), .B(A[586]), .Z(n924) );
  XOR U925 ( .A(n925), .B(n926), .Z(DIFF[585]) );
  XOR U926 ( .A(B[585]), .B(A[585]), .Z(n926) );
  XOR U927 ( .A(n927), .B(n928), .Z(DIFF[584]) );
  XOR U928 ( .A(B[584]), .B(A[584]), .Z(n928) );
  XOR U929 ( .A(n929), .B(n930), .Z(DIFF[583]) );
  XOR U930 ( .A(B[583]), .B(A[583]), .Z(n930) );
  XOR U931 ( .A(n931), .B(n932), .Z(DIFF[582]) );
  XOR U932 ( .A(B[582]), .B(A[582]), .Z(n932) );
  XOR U933 ( .A(n933), .B(n934), .Z(DIFF[581]) );
  XOR U934 ( .A(B[581]), .B(A[581]), .Z(n934) );
  XOR U935 ( .A(n935), .B(n936), .Z(DIFF[580]) );
  XOR U936 ( .A(B[580]), .B(A[580]), .Z(n936) );
  XOR U937 ( .A(n937), .B(n938), .Z(DIFF[57]) );
  XOR U938 ( .A(B[57]), .B(A[57]), .Z(n938) );
  XOR U939 ( .A(n939), .B(n940), .Z(DIFF[579]) );
  XOR U940 ( .A(B[579]), .B(A[579]), .Z(n940) );
  XOR U941 ( .A(n941), .B(n942), .Z(DIFF[578]) );
  XOR U942 ( .A(B[578]), .B(A[578]), .Z(n942) );
  XOR U943 ( .A(n943), .B(n944), .Z(DIFF[577]) );
  XOR U944 ( .A(B[577]), .B(A[577]), .Z(n944) );
  XOR U945 ( .A(n945), .B(n946), .Z(DIFF[576]) );
  XOR U946 ( .A(B[576]), .B(A[576]), .Z(n946) );
  XOR U947 ( .A(n947), .B(n948), .Z(DIFF[575]) );
  XOR U948 ( .A(B[575]), .B(A[575]), .Z(n948) );
  XOR U949 ( .A(n949), .B(n950), .Z(DIFF[574]) );
  XOR U950 ( .A(B[574]), .B(A[574]), .Z(n950) );
  XOR U951 ( .A(n951), .B(n952), .Z(DIFF[573]) );
  XOR U952 ( .A(B[573]), .B(A[573]), .Z(n952) );
  XOR U953 ( .A(n953), .B(n954), .Z(DIFF[572]) );
  XOR U954 ( .A(B[572]), .B(A[572]), .Z(n954) );
  XOR U955 ( .A(n955), .B(n956), .Z(DIFF[571]) );
  XOR U956 ( .A(B[571]), .B(A[571]), .Z(n956) );
  XOR U957 ( .A(n957), .B(n958), .Z(DIFF[570]) );
  XOR U958 ( .A(B[570]), .B(A[570]), .Z(n958) );
  XOR U959 ( .A(n959), .B(n960), .Z(DIFF[56]) );
  XOR U960 ( .A(B[56]), .B(A[56]), .Z(n960) );
  XOR U961 ( .A(n961), .B(n962), .Z(DIFF[569]) );
  XOR U962 ( .A(B[569]), .B(A[569]), .Z(n962) );
  XOR U963 ( .A(n963), .B(n964), .Z(DIFF[568]) );
  XOR U964 ( .A(B[568]), .B(A[568]), .Z(n964) );
  XOR U965 ( .A(n965), .B(n966), .Z(DIFF[567]) );
  XOR U966 ( .A(B[567]), .B(A[567]), .Z(n966) );
  XOR U967 ( .A(n967), .B(n968), .Z(DIFF[566]) );
  XOR U968 ( .A(B[566]), .B(A[566]), .Z(n968) );
  XOR U969 ( .A(n969), .B(n970), .Z(DIFF[565]) );
  XOR U970 ( .A(B[565]), .B(A[565]), .Z(n970) );
  XOR U971 ( .A(n971), .B(n972), .Z(DIFF[564]) );
  XOR U972 ( .A(B[564]), .B(A[564]), .Z(n972) );
  XOR U973 ( .A(n973), .B(n974), .Z(DIFF[563]) );
  XOR U974 ( .A(B[563]), .B(A[563]), .Z(n974) );
  XOR U975 ( .A(n975), .B(n976), .Z(DIFF[562]) );
  XOR U976 ( .A(B[562]), .B(A[562]), .Z(n976) );
  XOR U977 ( .A(n977), .B(n978), .Z(DIFF[561]) );
  XOR U978 ( .A(B[561]), .B(A[561]), .Z(n978) );
  XOR U979 ( .A(n979), .B(n980), .Z(DIFF[560]) );
  XOR U980 ( .A(B[560]), .B(A[560]), .Z(n980) );
  XOR U981 ( .A(n981), .B(n982), .Z(DIFF[55]) );
  XOR U982 ( .A(B[55]), .B(A[55]), .Z(n982) );
  XOR U983 ( .A(n983), .B(n984), .Z(DIFF[559]) );
  XOR U984 ( .A(B[559]), .B(A[559]), .Z(n984) );
  XOR U985 ( .A(n985), .B(n986), .Z(DIFF[558]) );
  XOR U986 ( .A(B[558]), .B(A[558]), .Z(n986) );
  XOR U987 ( .A(n987), .B(n988), .Z(DIFF[557]) );
  XOR U988 ( .A(B[557]), .B(A[557]), .Z(n988) );
  XOR U989 ( .A(n989), .B(n990), .Z(DIFF[556]) );
  XOR U990 ( .A(B[556]), .B(A[556]), .Z(n990) );
  XOR U991 ( .A(n991), .B(n992), .Z(DIFF[555]) );
  XOR U992 ( .A(B[555]), .B(A[555]), .Z(n992) );
  XOR U993 ( .A(n993), .B(n994), .Z(DIFF[554]) );
  XOR U994 ( .A(B[554]), .B(A[554]), .Z(n994) );
  XOR U995 ( .A(n995), .B(n996), .Z(DIFF[553]) );
  XOR U996 ( .A(B[553]), .B(A[553]), .Z(n996) );
  XOR U997 ( .A(n997), .B(n998), .Z(DIFF[552]) );
  XOR U998 ( .A(B[552]), .B(A[552]), .Z(n998) );
  XOR U999 ( .A(n999), .B(n1000), .Z(DIFF[551]) );
  XOR U1000 ( .A(B[551]), .B(A[551]), .Z(n1000) );
  XOR U1001 ( .A(n1001), .B(n1002), .Z(DIFF[550]) );
  XOR U1002 ( .A(B[550]), .B(A[550]), .Z(n1002) );
  XOR U1003 ( .A(n1003), .B(n1004), .Z(DIFF[54]) );
  XOR U1004 ( .A(B[54]), .B(A[54]), .Z(n1004) );
  XOR U1005 ( .A(n1005), .B(n1006), .Z(DIFF[549]) );
  XOR U1006 ( .A(B[549]), .B(A[549]), .Z(n1006) );
  XOR U1007 ( .A(n1007), .B(n1008), .Z(DIFF[548]) );
  XOR U1008 ( .A(B[548]), .B(A[548]), .Z(n1008) );
  XOR U1009 ( .A(n1009), .B(n1010), .Z(DIFF[547]) );
  XOR U1010 ( .A(B[547]), .B(A[547]), .Z(n1010) );
  XOR U1011 ( .A(n1011), .B(n1012), .Z(DIFF[546]) );
  XOR U1012 ( .A(B[546]), .B(A[546]), .Z(n1012) );
  XOR U1013 ( .A(n1013), .B(n1014), .Z(DIFF[545]) );
  XOR U1014 ( .A(B[545]), .B(A[545]), .Z(n1014) );
  XOR U1015 ( .A(n1015), .B(n1016), .Z(DIFF[544]) );
  XOR U1016 ( .A(B[544]), .B(A[544]), .Z(n1016) );
  XOR U1017 ( .A(n1017), .B(n1018), .Z(DIFF[543]) );
  XOR U1018 ( .A(B[543]), .B(A[543]), .Z(n1018) );
  XOR U1019 ( .A(n1019), .B(n1020), .Z(DIFF[542]) );
  XOR U1020 ( .A(B[542]), .B(A[542]), .Z(n1020) );
  XOR U1021 ( .A(n1021), .B(n1022), .Z(DIFF[541]) );
  XOR U1022 ( .A(B[541]), .B(A[541]), .Z(n1022) );
  XOR U1023 ( .A(n1023), .B(n1024), .Z(DIFF[540]) );
  XOR U1024 ( .A(B[540]), .B(A[540]), .Z(n1024) );
  XOR U1025 ( .A(n1025), .B(n1026), .Z(DIFF[53]) );
  XOR U1026 ( .A(B[53]), .B(A[53]), .Z(n1026) );
  XOR U1027 ( .A(n1027), .B(n1028), .Z(DIFF[539]) );
  XOR U1028 ( .A(B[539]), .B(A[539]), .Z(n1028) );
  XOR U1029 ( .A(n1029), .B(n1030), .Z(DIFF[538]) );
  XOR U1030 ( .A(B[538]), .B(A[538]), .Z(n1030) );
  XOR U1031 ( .A(n1031), .B(n1032), .Z(DIFF[537]) );
  XOR U1032 ( .A(B[537]), .B(A[537]), .Z(n1032) );
  XOR U1033 ( .A(n1033), .B(n1034), .Z(DIFF[536]) );
  XOR U1034 ( .A(B[536]), .B(A[536]), .Z(n1034) );
  XOR U1035 ( .A(n1035), .B(n1036), .Z(DIFF[535]) );
  XOR U1036 ( .A(B[535]), .B(A[535]), .Z(n1036) );
  XOR U1037 ( .A(n1037), .B(n1038), .Z(DIFF[534]) );
  XOR U1038 ( .A(B[534]), .B(A[534]), .Z(n1038) );
  XOR U1039 ( .A(n1039), .B(n1040), .Z(DIFF[533]) );
  XOR U1040 ( .A(B[533]), .B(A[533]), .Z(n1040) );
  XOR U1041 ( .A(n1041), .B(n1042), .Z(DIFF[532]) );
  XOR U1042 ( .A(B[532]), .B(A[532]), .Z(n1042) );
  XOR U1043 ( .A(n1043), .B(n1044), .Z(DIFF[531]) );
  XOR U1044 ( .A(B[531]), .B(A[531]), .Z(n1044) );
  XOR U1045 ( .A(n1045), .B(n1046), .Z(DIFF[530]) );
  XOR U1046 ( .A(B[530]), .B(A[530]), .Z(n1046) );
  XOR U1047 ( .A(n1047), .B(n1048), .Z(DIFF[52]) );
  XOR U1048 ( .A(B[52]), .B(A[52]), .Z(n1048) );
  XOR U1049 ( .A(n1049), .B(n1050), .Z(DIFF[529]) );
  XOR U1050 ( .A(B[529]), .B(A[529]), .Z(n1050) );
  XOR U1051 ( .A(n1051), .B(n1052), .Z(DIFF[528]) );
  XOR U1052 ( .A(B[528]), .B(A[528]), .Z(n1052) );
  XOR U1053 ( .A(n1053), .B(n1054), .Z(DIFF[527]) );
  XOR U1054 ( .A(B[527]), .B(A[527]), .Z(n1054) );
  XOR U1055 ( .A(n1055), .B(n1056), .Z(DIFF[526]) );
  XOR U1056 ( .A(B[526]), .B(A[526]), .Z(n1056) );
  XOR U1057 ( .A(n1057), .B(n1058), .Z(DIFF[525]) );
  XOR U1058 ( .A(B[525]), .B(A[525]), .Z(n1058) );
  XOR U1059 ( .A(n1059), .B(n1060), .Z(DIFF[524]) );
  XOR U1060 ( .A(B[524]), .B(A[524]), .Z(n1060) );
  XOR U1061 ( .A(n1061), .B(n1062), .Z(DIFF[523]) );
  XOR U1062 ( .A(B[523]), .B(A[523]), .Z(n1062) );
  XOR U1063 ( .A(n1063), .B(n1064), .Z(DIFF[522]) );
  XOR U1064 ( .A(B[522]), .B(A[522]), .Z(n1064) );
  XOR U1065 ( .A(n1065), .B(n1066), .Z(DIFF[521]) );
  XOR U1066 ( .A(B[521]), .B(A[521]), .Z(n1066) );
  XOR U1067 ( .A(n1067), .B(n1068), .Z(DIFF[520]) );
  XOR U1068 ( .A(B[520]), .B(A[520]), .Z(n1068) );
  XOR U1069 ( .A(n1069), .B(n1070), .Z(DIFF[51]) );
  XOR U1070 ( .A(B[51]), .B(A[51]), .Z(n1070) );
  XOR U1071 ( .A(n1071), .B(n1072), .Z(DIFF[519]) );
  XOR U1072 ( .A(B[519]), .B(A[519]), .Z(n1072) );
  XOR U1073 ( .A(n1073), .B(n1074), .Z(DIFF[518]) );
  XOR U1074 ( .A(B[518]), .B(A[518]), .Z(n1074) );
  XOR U1075 ( .A(n1075), .B(n1076), .Z(DIFF[517]) );
  XOR U1076 ( .A(B[517]), .B(A[517]), .Z(n1076) );
  XOR U1077 ( .A(n1077), .B(n1078), .Z(DIFF[516]) );
  XOR U1078 ( .A(B[516]), .B(A[516]), .Z(n1078) );
  XOR U1079 ( .A(n1079), .B(n1080), .Z(DIFF[515]) );
  XOR U1080 ( .A(B[515]), .B(A[515]), .Z(n1080) );
  XOR U1081 ( .A(n1081), .B(n1082), .Z(DIFF[514]) );
  XOR U1082 ( .A(B[514]), .B(A[514]), .Z(n1082) );
  XOR U1083 ( .A(n1083), .B(n1084), .Z(DIFF[513]) );
  XOR U1084 ( .A(B[513]), .B(A[513]), .Z(n1084) );
  XOR U1085 ( .A(n1085), .B(n1086), .Z(DIFF[512]) );
  XOR U1086 ( .A(B[512]), .B(A[512]), .Z(n1086) );
  XOR U1087 ( .A(n1087), .B(n1088), .Z(DIFF[511]) );
  XOR U1088 ( .A(B[511]), .B(A[511]), .Z(n1088) );
  XOR U1089 ( .A(n1089), .B(n1090), .Z(DIFF[510]) );
  XOR U1090 ( .A(B[510]), .B(A[510]), .Z(n1090) );
  XOR U1091 ( .A(n1091), .B(n1092), .Z(DIFF[50]) );
  XOR U1092 ( .A(B[50]), .B(A[50]), .Z(n1092) );
  XOR U1093 ( .A(n1093), .B(n1094), .Z(DIFF[509]) );
  XOR U1094 ( .A(B[509]), .B(A[509]), .Z(n1094) );
  XOR U1095 ( .A(n1095), .B(n1096), .Z(DIFF[508]) );
  XOR U1096 ( .A(B[508]), .B(A[508]), .Z(n1096) );
  XOR U1097 ( .A(n1097), .B(n1098), .Z(DIFF[507]) );
  XOR U1098 ( .A(B[507]), .B(A[507]), .Z(n1098) );
  XOR U1099 ( .A(n1099), .B(n1100), .Z(DIFF[506]) );
  XOR U1100 ( .A(B[506]), .B(A[506]), .Z(n1100) );
  XOR U1101 ( .A(n1101), .B(n1102), .Z(DIFF[505]) );
  XOR U1102 ( .A(B[505]), .B(A[505]), .Z(n1102) );
  XOR U1103 ( .A(n1103), .B(n1104), .Z(DIFF[504]) );
  XOR U1104 ( .A(B[504]), .B(A[504]), .Z(n1104) );
  XOR U1105 ( .A(n1105), .B(n1106), .Z(DIFF[503]) );
  XOR U1106 ( .A(B[503]), .B(A[503]), .Z(n1106) );
  XOR U1107 ( .A(n1107), .B(n1108), .Z(DIFF[502]) );
  XOR U1108 ( .A(B[502]), .B(A[502]), .Z(n1108) );
  XOR U1109 ( .A(n1109), .B(n1110), .Z(DIFF[501]) );
  XOR U1110 ( .A(B[501]), .B(A[501]), .Z(n1110) );
  XOR U1111 ( .A(n1111), .B(n1112), .Z(DIFF[500]) );
  XOR U1112 ( .A(B[500]), .B(A[500]), .Z(n1112) );
  XOR U1113 ( .A(n1113), .B(n1114), .Z(DIFF[4]) );
  XOR U1114 ( .A(B[4]), .B(A[4]), .Z(n1114) );
  XOR U1115 ( .A(n1115), .B(n1116), .Z(DIFF[49]) );
  XOR U1116 ( .A(B[49]), .B(A[49]), .Z(n1116) );
  XOR U1117 ( .A(n1117), .B(n1118), .Z(DIFF[499]) );
  XOR U1118 ( .A(B[499]), .B(A[499]), .Z(n1118) );
  XOR U1119 ( .A(n1119), .B(n1120), .Z(DIFF[498]) );
  XOR U1120 ( .A(B[498]), .B(A[498]), .Z(n1120) );
  XOR U1121 ( .A(n1121), .B(n1122), .Z(DIFF[497]) );
  XOR U1122 ( .A(B[497]), .B(A[497]), .Z(n1122) );
  XOR U1123 ( .A(n1123), .B(n1124), .Z(DIFF[496]) );
  XOR U1124 ( .A(B[496]), .B(A[496]), .Z(n1124) );
  XOR U1125 ( .A(n1125), .B(n1126), .Z(DIFF[495]) );
  XOR U1126 ( .A(B[495]), .B(A[495]), .Z(n1126) );
  XOR U1127 ( .A(n1127), .B(n1128), .Z(DIFF[494]) );
  XOR U1128 ( .A(B[494]), .B(A[494]), .Z(n1128) );
  XOR U1129 ( .A(n1129), .B(n1130), .Z(DIFF[493]) );
  XOR U1130 ( .A(B[493]), .B(A[493]), .Z(n1130) );
  XOR U1131 ( .A(n1131), .B(n1132), .Z(DIFF[492]) );
  XOR U1132 ( .A(B[492]), .B(A[492]), .Z(n1132) );
  XOR U1133 ( .A(n1133), .B(n1134), .Z(DIFF[491]) );
  XOR U1134 ( .A(B[491]), .B(A[491]), .Z(n1134) );
  XOR U1135 ( .A(n1135), .B(n1136), .Z(DIFF[490]) );
  XOR U1136 ( .A(B[490]), .B(A[490]), .Z(n1136) );
  XOR U1137 ( .A(n1137), .B(n1138), .Z(DIFF[48]) );
  XOR U1138 ( .A(B[48]), .B(A[48]), .Z(n1138) );
  XOR U1139 ( .A(n1139), .B(n1140), .Z(DIFF[489]) );
  XOR U1140 ( .A(B[489]), .B(A[489]), .Z(n1140) );
  XOR U1141 ( .A(n1141), .B(n1142), .Z(DIFF[488]) );
  XOR U1142 ( .A(B[488]), .B(A[488]), .Z(n1142) );
  XOR U1143 ( .A(n1143), .B(n1144), .Z(DIFF[487]) );
  XOR U1144 ( .A(B[487]), .B(A[487]), .Z(n1144) );
  XOR U1145 ( .A(n1145), .B(n1146), .Z(DIFF[486]) );
  XOR U1146 ( .A(B[486]), .B(A[486]), .Z(n1146) );
  XOR U1147 ( .A(n1147), .B(n1148), .Z(DIFF[485]) );
  XOR U1148 ( .A(B[485]), .B(A[485]), .Z(n1148) );
  XOR U1149 ( .A(n1149), .B(n1150), .Z(DIFF[484]) );
  XOR U1150 ( .A(B[484]), .B(A[484]), .Z(n1150) );
  XOR U1151 ( .A(n1151), .B(n1152), .Z(DIFF[483]) );
  XOR U1152 ( .A(B[483]), .B(A[483]), .Z(n1152) );
  XOR U1153 ( .A(n1153), .B(n1154), .Z(DIFF[482]) );
  XOR U1154 ( .A(B[482]), .B(A[482]), .Z(n1154) );
  XOR U1155 ( .A(n1155), .B(n1156), .Z(DIFF[481]) );
  XOR U1156 ( .A(B[481]), .B(A[481]), .Z(n1156) );
  XOR U1157 ( .A(n1157), .B(n1158), .Z(DIFF[480]) );
  XOR U1158 ( .A(B[480]), .B(A[480]), .Z(n1158) );
  XOR U1159 ( .A(n1159), .B(n1160), .Z(DIFF[47]) );
  XOR U1160 ( .A(B[47]), .B(A[47]), .Z(n1160) );
  XOR U1161 ( .A(n1161), .B(n1162), .Z(DIFF[479]) );
  XOR U1162 ( .A(B[479]), .B(A[479]), .Z(n1162) );
  XOR U1163 ( .A(n1163), .B(n1164), .Z(DIFF[478]) );
  XOR U1164 ( .A(B[478]), .B(A[478]), .Z(n1164) );
  XOR U1165 ( .A(n1165), .B(n1166), .Z(DIFF[477]) );
  XOR U1166 ( .A(B[477]), .B(A[477]), .Z(n1166) );
  XOR U1167 ( .A(n1167), .B(n1168), .Z(DIFF[476]) );
  XOR U1168 ( .A(B[476]), .B(A[476]), .Z(n1168) );
  XOR U1169 ( .A(n1169), .B(n1170), .Z(DIFF[475]) );
  XOR U1170 ( .A(B[475]), .B(A[475]), .Z(n1170) );
  XOR U1171 ( .A(n1171), .B(n1172), .Z(DIFF[474]) );
  XOR U1172 ( .A(B[474]), .B(A[474]), .Z(n1172) );
  XOR U1173 ( .A(n1173), .B(n1174), .Z(DIFF[473]) );
  XOR U1174 ( .A(B[473]), .B(A[473]), .Z(n1174) );
  XOR U1175 ( .A(n1175), .B(n1176), .Z(DIFF[472]) );
  XOR U1176 ( .A(B[472]), .B(A[472]), .Z(n1176) );
  XOR U1177 ( .A(n1177), .B(n1178), .Z(DIFF[471]) );
  XOR U1178 ( .A(B[471]), .B(A[471]), .Z(n1178) );
  XOR U1179 ( .A(n1179), .B(n1180), .Z(DIFF[470]) );
  XOR U1180 ( .A(B[470]), .B(A[470]), .Z(n1180) );
  XOR U1181 ( .A(n1181), .B(n1182), .Z(DIFF[46]) );
  XOR U1182 ( .A(B[46]), .B(A[46]), .Z(n1182) );
  XOR U1183 ( .A(n1183), .B(n1184), .Z(DIFF[469]) );
  XOR U1184 ( .A(B[469]), .B(A[469]), .Z(n1184) );
  XOR U1185 ( .A(n1185), .B(n1186), .Z(DIFF[468]) );
  XOR U1186 ( .A(B[468]), .B(A[468]), .Z(n1186) );
  XOR U1187 ( .A(n1187), .B(n1188), .Z(DIFF[467]) );
  XOR U1188 ( .A(B[467]), .B(A[467]), .Z(n1188) );
  XOR U1189 ( .A(n1189), .B(n1190), .Z(DIFF[466]) );
  XOR U1190 ( .A(B[466]), .B(A[466]), .Z(n1190) );
  XOR U1191 ( .A(n1191), .B(n1192), .Z(DIFF[465]) );
  XOR U1192 ( .A(B[465]), .B(A[465]), .Z(n1192) );
  XOR U1193 ( .A(n1193), .B(n1194), .Z(DIFF[464]) );
  XOR U1194 ( .A(B[464]), .B(A[464]), .Z(n1194) );
  XOR U1195 ( .A(n1195), .B(n1196), .Z(DIFF[463]) );
  XOR U1196 ( .A(B[463]), .B(A[463]), .Z(n1196) );
  XOR U1197 ( .A(n1197), .B(n1198), .Z(DIFF[462]) );
  XOR U1198 ( .A(B[462]), .B(A[462]), .Z(n1198) );
  XOR U1199 ( .A(n1199), .B(n1200), .Z(DIFF[461]) );
  XOR U1200 ( .A(B[461]), .B(A[461]), .Z(n1200) );
  XOR U1201 ( .A(n1201), .B(n1202), .Z(DIFF[460]) );
  XOR U1202 ( .A(B[460]), .B(A[460]), .Z(n1202) );
  XOR U1203 ( .A(n1203), .B(n1204), .Z(DIFF[45]) );
  XOR U1204 ( .A(B[45]), .B(A[45]), .Z(n1204) );
  XOR U1205 ( .A(n1205), .B(n1206), .Z(DIFF[459]) );
  XOR U1206 ( .A(B[459]), .B(A[459]), .Z(n1206) );
  XOR U1207 ( .A(n1207), .B(n1208), .Z(DIFF[458]) );
  XOR U1208 ( .A(B[458]), .B(A[458]), .Z(n1208) );
  XOR U1209 ( .A(n1209), .B(n1210), .Z(DIFF[457]) );
  XOR U1210 ( .A(B[457]), .B(A[457]), .Z(n1210) );
  XOR U1211 ( .A(n1211), .B(n1212), .Z(DIFF[456]) );
  XOR U1212 ( .A(B[456]), .B(A[456]), .Z(n1212) );
  XOR U1213 ( .A(n1213), .B(n1214), .Z(DIFF[455]) );
  XOR U1214 ( .A(B[455]), .B(A[455]), .Z(n1214) );
  XOR U1215 ( .A(n1215), .B(n1216), .Z(DIFF[454]) );
  XOR U1216 ( .A(B[454]), .B(A[454]), .Z(n1216) );
  XOR U1217 ( .A(n1217), .B(n1218), .Z(DIFF[453]) );
  XOR U1218 ( .A(B[453]), .B(A[453]), .Z(n1218) );
  XOR U1219 ( .A(n1219), .B(n1220), .Z(DIFF[452]) );
  XOR U1220 ( .A(B[452]), .B(A[452]), .Z(n1220) );
  XOR U1221 ( .A(n1221), .B(n1222), .Z(DIFF[451]) );
  XOR U1222 ( .A(B[451]), .B(A[451]), .Z(n1222) );
  XOR U1223 ( .A(n1223), .B(n1224), .Z(DIFF[450]) );
  XOR U1224 ( .A(B[450]), .B(A[450]), .Z(n1224) );
  XOR U1225 ( .A(n1225), .B(n1226), .Z(DIFF[44]) );
  XOR U1226 ( .A(B[44]), .B(A[44]), .Z(n1226) );
  XOR U1227 ( .A(n1227), .B(n1228), .Z(DIFF[449]) );
  XOR U1228 ( .A(B[449]), .B(A[449]), .Z(n1228) );
  XOR U1229 ( .A(n1229), .B(n1230), .Z(DIFF[448]) );
  XOR U1230 ( .A(B[448]), .B(A[448]), .Z(n1230) );
  XOR U1231 ( .A(n1231), .B(n1232), .Z(DIFF[447]) );
  XOR U1232 ( .A(B[447]), .B(A[447]), .Z(n1232) );
  XOR U1233 ( .A(n1233), .B(n1234), .Z(DIFF[446]) );
  XOR U1234 ( .A(B[446]), .B(A[446]), .Z(n1234) );
  XOR U1235 ( .A(n1235), .B(n1236), .Z(DIFF[445]) );
  XOR U1236 ( .A(B[445]), .B(A[445]), .Z(n1236) );
  XOR U1237 ( .A(n1237), .B(n1238), .Z(DIFF[444]) );
  XOR U1238 ( .A(B[444]), .B(A[444]), .Z(n1238) );
  XOR U1239 ( .A(n1239), .B(n1240), .Z(DIFF[443]) );
  XOR U1240 ( .A(B[443]), .B(A[443]), .Z(n1240) );
  XOR U1241 ( .A(n1241), .B(n1242), .Z(DIFF[442]) );
  XOR U1242 ( .A(B[442]), .B(A[442]), .Z(n1242) );
  XOR U1243 ( .A(n1243), .B(n1244), .Z(DIFF[441]) );
  XOR U1244 ( .A(B[441]), .B(A[441]), .Z(n1244) );
  XOR U1245 ( .A(n1245), .B(n1246), .Z(DIFF[440]) );
  XOR U1246 ( .A(B[440]), .B(A[440]), .Z(n1246) );
  XOR U1247 ( .A(n1247), .B(n1248), .Z(DIFF[43]) );
  XOR U1248 ( .A(B[43]), .B(A[43]), .Z(n1248) );
  XOR U1249 ( .A(n1249), .B(n1250), .Z(DIFF[439]) );
  XOR U1250 ( .A(B[439]), .B(A[439]), .Z(n1250) );
  XOR U1251 ( .A(n1251), .B(n1252), .Z(DIFF[438]) );
  XOR U1252 ( .A(B[438]), .B(A[438]), .Z(n1252) );
  XOR U1253 ( .A(n1253), .B(n1254), .Z(DIFF[437]) );
  XOR U1254 ( .A(B[437]), .B(A[437]), .Z(n1254) );
  XOR U1255 ( .A(n1255), .B(n1256), .Z(DIFF[436]) );
  XOR U1256 ( .A(B[436]), .B(A[436]), .Z(n1256) );
  XOR U1257 ( .A(n1257), .B(n1258), .Z(DIFF[435]) );
  XOR U1258 ( .A(B[435]), .B(A[435]), .Z(n1258) );
  XOR U1259 ( .A(n1259), .B(n1260), .Z(DIFF[434]) );
  XOR U1260 ( .A(B[434]), .B(A[434]), .Z(n1260) );
  XOR U1261 ( .A(n1261), .B(n1262), .Z(DIFF[433]) );
  XOR U1262 ( .A(B[433]), .B(A[433]), .Z(n1262) );
  XOR U1263 ( .A(n1263), .B(n1264), .Z(DIFF[432]) );
  XOR U1264 ( .A(B[432]), .B(A[432]), .Z(n1264) );
  XOR U1265 ( .A(n1265), .B(n1266), .Z(DIFF[431]) );
  XOR U1266 ( .A(B[431]), .B(A[431]), .Z(n1266) );
  XOR U1267 ( .A(n1267), .B(n1268), .Z(DIFF[430]) );
  XOR U1268 ( .A(B[430]), .B(A[430]), .Z(n1268) );
  XOR U1269 ( .A(n1269), .B(n1270), .Z(DIFF[42]) );
  XOR U1270 ( .A(B[42]), .B(A[42]), .Z(n1270) );
  XOR U1271 ( .A(n1271), .B(n1272), .Z(DIFF[429]) );
  XOR U1272 ( .A(B[429]), .B(A[429]), .Z(n1272) );
  XOR U1273 ( .A(n1273), .B(n1274), .Z(DIFF[428]) );
  XOR U1274 ( .A(B[428]), .B(A[428]), .Z(n1274) );
  XOR U1275 ( .A(n1275), .B(n1276), .Z(DIFF[427]) );
  XOR U1276 ( .A(B[427]), .B(A[427]), .Z(n1276) );
  XOR U1277 ( .A(n1277), .B(n1278), .Z(DIFF[426]) );
  XOR U1278 ( .A(B[426]), .B(A[426]), .Z(n1278) );
  XOR U1279 ( .A(n1279), .B(n1280), .Z(DIFF[425]) );
  XOR U1280 ( .A(B[425]), .B(A[425]), .Z(n1280) );
  XOR U1281 ( .A(n1281), .B(n1282), .Z(DIFF[424]) );
  XOR U1282 ( .A(B[424]), .B(A[424]), .Z(n1282) );
  XOR U1283 ( .A(n1283), .B(n1284), .Z(DIFF[423]) );
  XOR U1284 ( .A(B[423]), .B(A[423]), .Z(n1284) );
  XOR U1285 ( .A(n1285), .B(n1286), .Z(DIFF[422]) );
  XOR U1286 ( .A(B[422]), .B(A[422]), .Z(n1286) );
  XOR U1287 ( .A(n1287), .B(n1288), .Z(DIFF[421]) );
  XOR U1288 ( .A(B[421]), .B(A[421]), .Z(n1288) );
  XOR U1289 ( .A(n1289), .B(n1290), .Z(DIFF[420]) );
  XOR U1290 ( .A(B[420]), .B(A[420]), .Z(n1290) );
  XOR U1291 ( .A(n1291), .B(n1292), .Z(DIFF[41]) );
  XOR U1292 ( .A(B[41]), .B(A[41]), .Z(n1292) );
  XOR U1293 ( .A(n1293), .B(n1294), .Z(DIFF[419]) );
  XOR U1294 ( .A(B[419]), .B(A[419]), .Z(n1294) );
  XOR U1295 ( .A(n1295), .B(n1296), .Z(DIFF[418]) );
  XOR U1296 ( .A(B[418]), .B(A[418]), .Z(n1296) );
  XOR U1297 ( .A(n1297), .B(n1298), .Z(DIFF[417]) );
  XOR U1298 ( .A(B[417]), .B(A[417]), .Z(n1298) );
  XOR U1299 ( .A(n1299), .B(n1300), .Z(DIFF[416]) );
  XOR U1300 ( .A(B[416]), .B(A[416]), .Z(n1300) );
  XOR U1301 ( .A(n1301), .B(n1302), .Z(DIFF[415]) );
  XOR U1302 ( .A(B[415]), .B(A[415]), .Z(n1302) );
  XOR U1303 ( .A(n1303), .B(n1304), .Z(DIFF[414]) );
  XOR U1304 ( .A(B[414]), .B(A[414]), .Z(n1304) );
  XOR U1305 ( .A(n1305), .B(n1306), .Z(DIFF[413]) );
  XOR U1306 ( .A(B[413]), .B(A[413]), .Z(n1306) );
  XOR U1307 ( .A(n1307), .B(n1308), .Z(DIFF[412]) );
  XOR U1308 ( .A(B[412]), .B(A[412]), .Z(n1308) );
  XOR U1309 ( .A(n1309), .B(n1310), .Z(DIFF[411]) );
  XOR U1310 ( .A(B[411]), .B(A[411]), .Z(n1310) );
  XOR U1311 ( .A(n1311), .B(n1312), .Z(DIFF[410]) );
  XOR U1312 ( .A(B[410]), .B(A[410]), .Z(n1312) );
  XOR U1313 ( .A(n1313), .B(n1314), .Z(DIFF[40]) );
  XOR U1314 ( .A(B[40]), .B(A[40]), .Z(n1314) );
  XOR U1315 ( .A(n1315), .B(n1316), .Z(DIFF[409]) );
  XOR U1316 ( .A(B[409]), .B(A[409]), .Z(n1316) );
  XOR U1317 ( .A(n1317), .B(n1318), .Z(DIFF[408]) );
  XOR U1318 ( .A(B[408]), .B(A[408]), .Z(n1318) );
  XOR U1319 ( .A(n1319), .B(n1320), .Z(DIFF[407]) );
  XOR U1320 ( .A(B[407]), .B(A[407]), .Z(n1320) );
  XOR U1321 ( .A(n1321), .B(n1322), .Z(DIFF[406]) );
  XOR U1322 ( .A(B[406]), .B(A[406]), .Z(n1322) );
  XOR U1323 ( .A(n1323), .B(n1324), .Z(DIFF[405]) );
  XOR U1324 ( .A(B[405]), .B(A[405]), .Z(n1324) );
  XOR U1325 ( .A(n1325), .B(n1326), .Z(DIFF[404]) );
  XOR U1326 ( .A(B[404]), .B(A[404]), .Z(n1326) );
  XOR U1327 ( .A(n1327), .B(n1328), .Z(DIFF[403]) );
  XOR U1328 ( .A(B[403]), .B(A[403]), .Z(n1328) );
  XOR U1329 ( .A(n1329), .B(n1330), .Z(DIFF[402]) );
  XOR U1330 ( .A(B[402]), .B(A[402]), .Z(n1330) );
  XOR U1331 ( .A(n1331), .B(n1332), .Z(DIFF[401]) );
  XOR U1332 ( .A(B[401]), .B(A[401]), .Z(n1332) );
  XOR U1333 ( .A(n1333), .B(n1334), .Z(DIFF[400]) );
  XOR U1334 ( .A(B[400]), .B(A[400]), .Z(n1334) );
  XOR U1335 ( .A(n1335), .B(n1336), .Z(DIFF[3]) );
  XOR U1336 ( .A(B[3]), .B(A[3]), .Z(n1336) );
  XOR U1337 ( .A(n1337), .B(n1338), .Z(DIFF[39]) );
  XOR U1338 ( .A(B[39]), .B(A[39]), .Z(n1338) );
  XOR U1339 ( .A(n1339), .B(n1340), .Z(DIFF[399]) );
  XOR U1340 ( .A(B[399]), .B(A[399]), .Z(n1340) );
  XOR U1341 ( .A(n1341), .B(n1342), .Z(DIFF[398]) );
  XOR U1342 ( .A(B[398]), .B(A[398]), .Z(n1342) );
  XOR U1343 ( .A(n1343), .B(n1344), .Z(DIFF[397]) );
  XOR U1344 ( .A(B[397]), .B(A[397]), .Z(n1344) );
  XOR U1345 ( .A(n1345), .B(n1346), .Z(DIFF[396]) );
  XOR U1346 ( .A(B[396]), .B(A[396]), .Z(n1346) );
  XOR U1347 ( .A(n1347), .B(n1348), .Z(DIFF[395]) );
  XOR U1348 ( .A(B[395]), .B(A[395]), .Z(n1348) );
  XOR U1349 ( .A(n1349), .B(n1350), .Z(DIFF[394]) );
  XOR U1350 ( .A(B[394]), .B(A[394]), .Z(n1350) );
  XOR U1351 ( .A(n1351), .B(n1352), .Z(DIFF[393]) );
  XOR U1352 ( .A(B[393]), .B(A[393]), .Z(n1352) );
  XOR U1353 ( .A(n1353), .B(n1354), .Z(DIFF[392]) );
  XOR U1354 ( .A(B[392]), .B(A[392]), .Z(n1354) );
  XOR U1355 ( .A(n1355), .B(n1356), .Z(DIFF[391]) );
  XOR U1356 ( .A(B[391]), .B(A[391]), .Z(n1356) );
  XOR U1357 ( .A(n1357), .B(n1358), .Z(DIFF[390]) );
  XOR U1358 ( .A(B[390]), .B(A[390]), .Z(n1358) );
  XOR U1359 ( .A(n1359), .B(n1360), .Z(DIFF[38]) );
  XOR U1360 ( .A(B[38]), .B(A[38]), .Z(n1360) );
  XOR U1361 ( .A(n1361), .B(n1362), .Z(DIFF[389]) );
  XOR U1362 ( .A(B[389]), .B(A[389]), .Z(n1362) );
  XOR U1363 ( .A(n1363), .B(n1364), .Z(DIFF[388]) );
  XOR U1364 ( .A(B[388]), .B(A[388]), .Z(n1364) );
  XOR U1365 ( .A(n1365), .B(n1366), .Z(DIFF[387]) );
  XOR U1366 ( .A(B[387]), .B(A[387]), .Z(n1366) );
  XOR U1367 ( .A(n1367), .B(n1368), .Z(DIFF[386]) );
  XOR U1368 ( .A(B[386]), .B(A[386]), .Z(n1368) );
  XOR U1369 ( .A(n1369), .B(n1370), .Z(DIFF[385]) );
  XOR U1370 ( .A(B[385]), .B(A[385]), .Z(n1370) );
  XOR U1371 ( .A(n1371), .B(n1372), .Z(DIFF[384]) );
  XOR U1372 ( .A(B[384]), .B(A[384]), .Z(n1372) );
  XOR U1373 ( .A(n1373), .B(n1374), .Z(DIFF[383]) );
  XOR U1374 ( .A(B[383]), .B(A[383]), .Z(n1374) );
  XOR U1375 ( .A(n1375), .B(n1376), .Z(DIFF[382]) );
  XOR U1376 ( .A(B[382]), .B(A[382]), .Z(n1376) );
  XOR U1377 ( .A(n1377), .B(n1378), .Z(DIFF[381]) );
  XOR U1378 ( .A(B[381]), .B(A[381]), .Z(n1378) );
  XOR U1379 ( .A(n1379), .B(n1380), .Z(DIFF[380]) );
  XOR U1380 ( .A(B[380]), .B(A[380]), .Z(n1380) );
  XOR U1381 ( .A(n1381), .B(n1382), .Z(DIFF[37]) );
  XOR U1382 ( .A(B[37]), .B(A[37]), .Z(n1382) );
  XOR U1383 ( .A(n1383), .B(n1384), .Z(DIFF[379]) );
  XOR U1384 ( .A(B[379]), .B(A[379]), .Z(n1384) );
  XOR U1385 ( .A(n1385), .B(n1386), .Z(DIFF[378]) );
  XOR U1386 ( .A(B[378]), .B(A[378]), .Z(n1386) );
  XOR U1387 ( .A(n1387), .B(n1388), .Z(DIFF[377]) );
  XOR U1388 ( .A(B[377]), .B(A[377]), .Z(n1388) );
  XOR U1389 ( .A(n1389), .B(n1390), .Z(DIFF[376]) );
  XOR U1390 ( .A(B[376]), .B(A[376]), .Z(n1390) );
  XOR U1391 ( .A(n1391), .B(n1392), .Z(DIFF[375]) );
  XOR U1392 ( .A(B[375]), .B(A[375]), .Z(n1392) );
  XOR U1393 ( .A(n1393), .B(n1394), .Z(DIFF[374]) );
  XOR U1394 ( .A(B[374]), .B(A[374]), .Z(n1394) );
  XOR U1395 ( .A(n1395), .B(n1396), .Z(DIFF[373]) );
  XOR U1396 ( .A(B[373]), .B(A[373]), .Z(n1396) );
  XOR U1397 ( .A(n1397), .B(n1398), .Z(DIFF[372]) );
  XOR U1398 ( .A(B[372]), .B(A[372]), .Z(n1398) );
  XOR U1399 ( .A(n1399), .B(n1400), .Z(DIFF[371]) );
  XOR U1400 ( .A(B[371]), .B(A[371]), .Z(n1400) );
  XOR U1401 ( .A(n1401), .B(n1402), .Z(DIFF[370]) );
  XOR U1402 ( .A(B[370]), .B(A[370]), .Z(n1402) );
  XOR U1403 ( .A(n1403), .B(n1404), .Z(DIFF[36]) );
  XOR U1404 ( .A(B[36]), .B(A[36]), .Z(n1404) );
  XOR U1405 ( .A(n1405), .B(n1406), .Z(DIFF[369]) );
  XOR U1406 ( .A(B[369]), .B(A[369]), .Z(n1406) );
  XOR U1407 ( .A(n1407), .B(n1408), .Z(DIFF[368]) );
  XOR U1408 ( .A(B[368]), .B(A[368]), .Z(n1408) );
  XOR U1409 ( .A(n1409), .B(n1410), .Z(DIFF[367]) );
  XOR U1410 ( .A(B[367]), .B(A[367]), .Z(n1410) );
  XOR U1411 ( .A(n1411), .B(n1412), .Z(DIFF[366]) );
  XOR U1412 ( .A(B[366]), .B(A[366]), .Z(n1412) );
  XOR U1413 ( .A(n1413), .B(n1414), .Z(DIFF[365]) );
  XOR U1414 ( .A(B[365]), .B(A[365]), .Z(n1414) );
  XOR U1415 ( .A(n1415), .B(n1416), .Z(DIFF[364]) );
  XOR U1416 ( .A(B[364]), .B(A[364]), .Z(n1416) );
  XOR U1417 ( .A(n1417), .B(n1418), .Z(DIFF[363]) );
  XOR U1418 ( .A(B[363]), .B(A[363]), .Z(n1418) );
  XOR U1419 ( .A(n1419), .B(n1420), .Z(DIFF[362]) );
  XOR U1420 ( .A(B[362]), .B(A[362]), .Z(n1420) );
  XOR U1421 ( .A(n1421), .B(n1422), .Z(DIFF[361]) );
  XOR U1422 ( .A(B[361]), .B(A[361]), .Z(n1422) );
  XOR U1423 ( .A(n1423), .B(n1424), .Z(DIFF[360]) );
  XOR U1424 ( .A(B[360]), .B(A[360]), .Z(n1424) );
  XOR U1425 ( .A(n1425), .B(n1426), .Z(DIFF[35]) );
  XOR U1426 ( .A(B[35]), .B(A[35]), .Z(n1426) );
  XOR U1427 ( .A(n1427), .B(n1428), .Z(DIFF[359]) );
  XOR U1428 ( .A(B[359]), .B(A[359]), .Z(n1428) );
  XOR U1429 ( .A(n1429), .B(n1430), .Z(DIFF[358]) );
  XOR U1430 ( .A(B[358]), .B(A[358]), .Z(n1430) );
  XOR U1431 ( .A(n1431), .B(n1432), .Z(DIFF[357]) );
  XOR U1432 ( .A(B[357]), .B(A[357]), .Z(n1432) );
  XOR U1433 ( .A(n1433), .B(n1434), .Z(DIFF[356]) );
  XOR U1434 ( .A(B[356]), .B(A[356]), .Z(n1434) );
  XOR U1435 ( .A(n1435), .B(n1436), .Z(DIFF[355]) );
  XOR U1436 ( .A(B[355]), .B(A[355]), .Z(n1436) );
  XOR U1437 ( .A(n1437), .B(n1438), .Z(DIFF[354]) );
  XOR U1438 ( .A(B[354]), .B(A[354]), .Z(n1438) );
  XOR U1439 ( .A(n1439), .B(n1440), .Z(DIFF[353]) );
  XOR U1440 ( .A(B[353]), .B(A[353]), .Z(n1440) );
  XOR U1441 ( .A(n1441), .B(n1442), .Z(DIFF[352]) );
  XOR U1442 ( .A(B[352]), .B(A[352]), .Z(n1442) );
  XOR U1443 ( .A(n1443), .B(n1444), .Z(DIFF[351]) );
  XOR U1444 ( .A(B[351]), .B(A[351]), .Z(n1444) );
  XOR U1445 ( .A(n1445), .B(n1446), .Z(DIFF[350]) );
  XOR U1446 ( .A(B[350]), .B(A[350]), .Z(n1446) );
  XOR U1447 ( .A(n1447), .B(n1448), .Z(DIFF[34]) );
  XOR U1448 ( .A(B[34]), .B(A[34]), .Z(n1448) );
  XOR U1449 ( .A(n1449), .B(n1450), .Z(DIFF[349]) );
  XOR U1450 ( .A(B[349]), .B(A[349]), .Z(n1450) );
  XOR U1451 ( .A(n1451), .B(n1452), .Z(DIFF[348]) );
  XOR U1452 ( .A(B[348]), .B(A[348]), .Z(n1452) );
  XOR U1453 ( .A(n1453), .B(n1454), .Z(DIFF[347]) );
  XOR U1454 ( .A(B[347]), .B(A[347]), .Z(n1454) );
  XOR U1455 ( .A(n1455), .B(n1456), .Z(DIFF[346]) );
  XOR U1456 ( .A(B[346]), .B(A[346]), .Z(n1456) );
  XOR U1457 ( .A(n1457), .B(n1458), .Z(DIFF[345]) );
  XOR U1458 ( .A(B[345]), .B(A[345]), .Z(n1458) );
  XOR U1459 ( .A(n1459), .B(n1460), .Z(DIFF[344]) );
  XOR U1460 ( .A(B[344]), .B(A[344]), .Z(n1460) );
  XOR U1461 ( .A(n1461), .B(n1462), .Z(DIFF[343]) );
  XOR U1462 ( .A(B[343]), .B(A[343]), .Z(n1462) );
  XOR U1463 ( .A(n1463), .B(n1464), .Z(DIFF[342]) );
  XOR U1464 ( .A(B[342]), .B(A[342]), .Z(n1464) );
  XOR U1465 ( .A(n1465), .B(n1466), .Z(DIFF[341]) );
  XOR U1466 ( .A(B[341]), .B(A[341]), .Z(n1466) );
  XOR U1467 ( .A(n1467), .B(n1468), .Z(DIFF[340]) );
  XOR U1468 ( .A(B[340]), .B(A[340]), .Z(n1468) );
  XOR U1469 ( .A(n1469), .B(n1470), .Z(DIFF[33]) );
  XOR U1470 ( .A(B[33]), .B(A[33]), .Z(n1470) );
  XOR U1471 ( .A(n1471), .B(n1472), .Z(DIFF[339]) );
  XOR U1472 ( .A(B[339]), .B(A[339]), .Z(n1472) );
  XOR U1473 ( .A(n1473), .B(n1474), .Z(DIFF[338]) );
  XOR U1474 ( .A(B[338]), .B(A[338]), .Z(n1474) );
  XOR U1475 ( .A(n1475), .B(n1476), .Z(DIFF[337]) );
  XOR U1476 ( .A(B[337]), .B(A[337]), .Z(n1476) );
  XOR U1477 ( .A(n1477), .B(n1478), .Z(DIFF[336]) );
  XOR U1478 ( .A(B[336]), .B(A[336]), .Z(n1478) );
  XOR U1479 ( .A(n1479), .B(n1480), .Z(DIFF[335]) );
  XOR U1480 ( .A(B[335]), .B(A[335]), .Z(n1480) );
  XOR U1481 ( .A(n1481), .B(n1482), .Z(DIFF[334]) );
  XOR U1482 ( .A(B[334]), .B(A[334]), .Z(n1482) );
  XOR U1483 ( .A(n1483), .B(n1484), .Z(DIFF[333]) );
  XOR U1484 ( .A(B[333]), .B(A[333]), .Z(n1484) );
  XOR U1485 ( .A(n1485), .B(n1486), .Z(DIFF[332]) );
  XOR U1486 ( .A(B[332]), .B(A[332]), .Z(n1486) );
  XOR U1487 ( .A(n1487), .B(n1488), .Z(DIFF[331]) );
  XOR U1488 ( .A(B[331]), .B(A[331]), .Z(n1488) );
  XOR U1489 ( .A(n1489), .B(n1490), .Z(DIFF[330]) );
  XOR U1490 ( .A(B[330]), .B(A[330]), .Z(n1490) );
  XOR U1491 ( .A(n1491), .B(n1492), .Z(DIFF[32]) );
  XOR U1492 ( .A(B[32]), .B(A[32]), .Z(n1492) );
  XOR U1493 ( .A(n1493), .B(n1494), .Z(DIFF[329]) );
  XOR U1494 ( .A(B[329]), .B(A[329]), .Z(n1494) );
  XOR U1495 ( .A(n1495), .B(n1496), .Z(DIFF[328]) );
  XOR U1496 ( .A(B[328]), .B(A[328]), .Z(n1496) );
  XOR U1497 ( .A(n1497), .B(n1498), .Z(DIFF[327]) );
  XOR U1498 ( .A(B[327]), .B(A[327]), .Z(n1498) );
  XOR U1499 ( .A(n1499), .B(n1500), .Z(DIFF[326]) );
  XOR U1500 ( .A(B[326]), .B(A[326]), .Z(n1500) );
  XOR U1501 ( .A(n1501), .B(n1502), .Z(DIFF[325]) );
  XOR U1502 ( .A(B[325]), .B(A[325]), .Z(n1502) );
  XOR U1503 ( .A(n1503), .B(n1504), .Z(DIFF[324]) );
  XOR U1504 ( .A(B[324]), .B(A[324]), .Z(n1504) );
  XOR U1505 ( .A(n1505), .B(n1506), .Z(DIFF[323]) );
  XOR U1506 ( .A(B[323]), .B(A[323]), .Z(n1506) );
  XOR U1507 ( .A(n1507), .B(n1508), .Z(DIFF[322]) );
  XOR U1508 ( .A(B[322]), .B(A[322]), .Z(n1508) );
  XOR U1509 ( .A(n1509), .B(n1510), .Z(DIFF[321]) );
  XOR U1510 ( .A(B[321]), .B(A[321]), .Z(n1510) );
  XOR U1511 ( .A(n1511), .B(n1512), .Z(DIFF[320]) );
  XOR U1512 ( .A(B[320]), .B(A[320]), .Z(n1512) );
  XOR U1513 ( .A(n1513), .B(n1514), .Z(DIFF[31]) );
  XOR U1514 ( .A(B[31]), .B(A[31]), .Z(n1514) );
  XOR U1515 ( .A(n1515), .B(n1516), .Z(DIFF[319]) );
  XOR U1516 ( .A(B[319]), .B(A[319]), .Z(n1516) );
  XOR U1517 ( .A(n1517), .B(n1518), .Z(DIFF[318]) );
  XOR U1518 ( .A(B[318]), .B(A[318]), .Z(n1518) );
  XOR U1519 ( .A(n1519), .B(n1520), .Z(DIFF[317]) );
  XOR U1520 ( .A(B[317]), .B(A[317]), .Z(n1520) );
  XOR U1521 ( .A(n1521), .B(n1522), .Z(DIFF[316]) );
  XOR U1522 ( .A(B[316]), .B(A[316]), .Z(n1522) );
  XOR U1523 ( .A(n1523), .B(n1524), .Z(DIFF[315]) );
  XOR U1524 ( .A(B[315]), .B(A[315]), .Z(n1524) );
  XOR U1525 ( .A(n1525), .B(n1526), .Z(DIFF[314]) );
  XOR U1526 ( .A(B[314]), .B(A[314]), .Z(n1526) );
  XOR U1527 ( .A(n1527), .B(n1528), .Z(DIFF[313]) );
  XOR U1528 ( .A(B[313]), .B(A[313]), .Z(n1528) );
  XOR U1529 ( .A(n1529), .B(n1530), .Z(DIFF[312]) );
  XOR U1530 ( .A(B[312]), .B(A[312]), .Z(n1530) );
  XOR U1531 ( .A(n1531), .B(n1532), .Z(DIFF[311]) );
  XOR U1532 ( .A(B[311]), .B(A[311]), .Z(n1532) );
  XOR U1533 ( .A(n1533), .B(n1534), .Z(DIFF[310]) );
  XOR U1534 ( .A(B[310]), .B(A[310]), .Z(n1534) );
  XOR U1535 ( .A(n1535), .B(n1536), .Z(DIFF[30]) );
  XOR U1536 ( .A(B[30]), .B(A[30]), .Z(n1536) );
  XOR U1537 ( .A(n1537), .B(n1538), .Z(DIFF[309]) );
  XOR U1538 ( .A(B[309]), .B(A[309]), .Z(n1538) );
  XOR U1539 ( .A(n1539), .B(n1540), .Z(DIFF[308]) );
  XOR U1540 ( .A(B[308]), .B(A[308]), .Z(n1540) );
  XOR U1541 ( .A(n1541), .B(n1542), .Z(DIFF[307]) );
  XOR U1542 ( .A(B[307]), .B(A[307]), .Z(n1542) );
  XOR U1543 ( .A(n1543), .B(n1544), .Z(DIFF[306]) );
  XOR U1544 ( .A(B[306]), .B(A[306]), .Z(n1544) );
  XOR U1545 ( .A(n1545), .B(n1546), .Z(DIFF[305]) );
  XOR U1546 ( .A(B[305]), .B(A[305]), .Z(n1546) );
  XOR U1547 ( .A(n1547), .B(n1548), .Z(DIFF[304]) );
  XOR U1548 ( .A(B[304]), .B(A[304]), .Z(n1548) );
  XOR U1549 ( .A(n1549), .B(n1550), .Z(DIFF[303]) );
  XOR U1550 ( .A(B[303]), .B(A[303]), .Z(n1550) );
  XOR U1551 ( .A(n1551), .B(n1552), .Z(DIFF[302]) );
  XOR U1552 ( .A(B[302]), .B(A[302]), .Z(n1552) );
  XOR U1553 ( .A(n1553), .B(n1554), .Z(DIFF[301]) );
  XOR U1554 ( .A(B[301]), .B(A[301]), .Z(n1554) );
  XOR U1555 ( .A(n1555), .B(n1556), .Z(DIFF[300]) );
  XOR U1556 ( .A(B[300]), .B(A[300]), .Z(n1556) );
  XOR U1557 ( .A(n1557), .B(n1558), .Z(DIFF[2]) );
  XOR U1558 ( .A(B[2]), .B(A[2]), .Z(n1558) );
  XOR U1559 ( .A(n1559), .B(n1560), .Z(DIFF[29]) );
  XOR U1560 ( .A(B[29]), .B(A[29]), .Z(n1560) );
  XOR U1561 ( .A(n1561), .B(n1562), .Z(DIFF[299]) );
  XOR U1562 ( .A(B[299]), .B(A[299]), .Z(n1562) );
  XOR U1563 ( .A(n1563), .B(n1564), .Z(DIFF[298]) );
  XOR U1564 ( .A(B[298]), .B(A[298]), .Z(n1564) );
  XOR U1565 ( .A(n1565), .B(n1566), .Z(DIFF[297]) );
  XOR U1566 ( .A(B[297]), .B(A[297]), .Z(n1566) );
  XOR U1567 ( .A(n1567), .B(n1568), .Z(DIFF[296]) );
  XOR U1568 ( .A(B[296]), .B(A[296]), .Z(n1568) );
  XOR U1569 ( .A(n1569), .B(n1570), .Z(DIFF[295]) );
  XOR U1570 ( .A(B[295]), .B(A[295]), .Z(n1570) );
  XOR U1571 ( .A(n1571), .B(n1572), .Z(DIFF[294]) );
  XOR U1572 ( .A(B[294]), .B(A[294]), .Z(n1572) );
  XOR U1573 ( .A(n1573), .B(n1574), .Z(DIFF[293]) );
  XOR U1574 ( .A(B[293]), .B(A[293]), .Z(n1574) );
  XOR U1575 ( .A(n1575), .B(n1576), .Z(DIFF[292]) );
  XOR U1576 ( .A(B[292]), .B(A[292]), .Z(n1576) );
  XOR U1577 ( .A(n1577), .B(n1578), .Z(DIFF[291]) );
  XOR U1578 ( .A(B[291]), .B(A[291]), .Z(n1578) );
  XOR U1579 ( .A(n1579), .B(n1580), .Z(DIFF[290]) );
  XOR U1580 ( .A(B[290]), .B(A[290]), .Z(n1580) );
  XOR U1581 ( .A(n1581), .B(n1582), .Z(DIFF[28]) );
  XOR U1582 ( .A(B[28]), .B(A[28]), .Z(n1582) );
  XOR U1583 ( .A(n1583), .B(n1584), .Z(DIFF[289]) );
  XOR U1584 ( .A(B[289]), .B(A[289]), .Z(n1584) );
  XOR U1585 ( .A(n1585), .B(n1586), .Z(DIFF[288]) );
  XOR U1586 ( .A(B[288]), .B(A[288]), .Z(n1586) );
  XOR U1587 ( .A(n1587), .B(n1588), .Z(DIFF[287]) );
  XOR U1588 ( .A(B[287]), .B(A[287]), .Z(n1588) );
  XOR U1589 ( .A(n1589), .B(n1590), .Z(DIFF[286]) );
  XOR U1590 ( .A(B[286]), .B(A[286]), .Z(n1590) );
  XOR U1591 ( .A(n1591), .B(n1592), .Z(DIFF[285]) );
  XOR U1592 ( .A(B[285]), .B(A[285]), .Z(n1592) );
  XOR U1593 ( .A(n1593), .B(n1594), .Z(DIFF[284]) );
  XOR U1594 ( .A(B[284]), .B(A[284]), .Z(n1594) );
  XOR U1595 ( .A(n1595), .B(n1596), .Z(DIFF[283]) );
  XOR U1596 ( .A(B[283]), .B(A[283]), .Z(n1596) );
  XOR U1597 ( .A(n1597), .B(n1598), .Z(DIFF[282]) );
  XOR U1598 ( .A(B[282]), .B(A[282]), .Z(n1598) );
  XOR U1599 ( .A(n1599), .B(n1600), .Z(DIFF[281]) );
  XOR U1600 ( .A(B[281]), .B(A[281]), .Z(n1600) );
  XOR U1601 ( .A(n1601), .B(n1602), .Z(DIFF[280]) );
  XOR U1602 ( .A(B[280]), .B(A[280]), .Z(n1602) );
  XOR U1603 ( .A(n1603), .B(n1604), .Z(DIFF[27]) );
  XOR U1604 ( .A(B[27]), .B(A[27]), .Z(n1604) );
  XOR U1605 ( .A(n1605), .B(n1606), .Z(DIFF[279]) );
  XOR U1606 ( .A(B[279]), .B(A[279]), .Z(n1606) );
  XOR U1607 ( .A(n1607), .B(n1608), .Z(DIFF[278]) );
  XOR U1608 ( .A(B[278]), .B(A[278]), .Z(n1608) );
  XOR U1609 ( .A(n1609), .B(n1610), .Z(DIFF[277]) );
  XOR U1610 ( .A(B[277]), .B(A[277]), .Z(n1610) );
  XOR U1611 ( .A(n1611), .B(n1612), .Z(DIFF[276]) );
  XOR U1612 ( .A(B[276]), .B(A[276]), .Z(n1612) );
  XOR U1613 ( .A(n1613), .B(n1614), .Z(DIFF[275]) );
  XOR U1614 ( .A(B[275]), .B(A[275]), .Z(n1614) );
  XOR U1615 ( .A(n1615), .B(n1616), .Z(DIFF[274]) );
  XOR U1616 ( .A(B[274]), .B(A[274]), .Z(n1616) );
  XOR U1617 ( .A(n1617), .B(n1618), .Z(DIFF[273]) );
  XOR U1618 ( .A(B[273]), .B(A[273]), .Z(n1618) );
  XOR U1619 ( .A(n1619), .B(n1620), .Z(DIFF[272]) );
  XOR U1620 ( .A(B[272]), .B(A[272]), .Z(n1620) );
  XOR U1621 ( .A(n1621), .B(n1622), .Z(DIFF[271]) );
  XOR U1622 ( .A(B[271]), .B(A[271]), .Z(n1622) );
  XOR U1623 ( .A(n1623), .B(n1624), .Z(DIFF[270]) );
  XOR U1624 ( .A(B[270]), .B(A[270]), .Z(n1624) );
  XOR U1625 ( .A(n1625), .B(n1626), .Z(DIFF[26]) );
  XOR U1626 ( .A(B[26]), .B(A[26]), .Z(n1626) );
  XOR U1627 ( .A(n1627), .B(n1628), .Z(DIFF[269]) );
  XOR U1628 ( .A(B[269]), .B(A[269]), .Z(n1628) );
  XOR U1629 ( .A(n1629), .B(n1630), .Z(DIFF[268]) );
  XOR U1630 ( .A(B[268]), .B(A[268]), .Z(n1630) );
  XOR U1631 ( .A(n1631), .B(n1632), .Z(DIFF[267]) );
  XOR U1632 ( .A(B[267]), .B(A[267]), .Z(n1632) );
  XOR U1633 ( .A(n1633), .B(n1634), .Z(DIFF[266]) );
  XOR U1634 ( .A(B[266]), .B(A[266]), .Z(n1634) );
  XOR U1635 ( .A(n1635), .B(n1636), .Z(DIFF[265]) );
  XOR U1636 ( .A(B[265]), .B(A[265]), .Z(n1636) );
  XOR U1637 ( .A(n1637), .B(n1638), .Z(DIFF[264]) );
  XOR U1638 ( .A(B[264]), .B(A[264]), .Z(n1638) );
  XOR U1639 ( .A(n1639), .B(n1640), .Z(DIFF[263]) );
  XOR U1640 ( .A(B[263]), .B(A[263]), .Z(n1640) );
  XOR U1641 ( .A(n1641), .B(n1642), .Z(DIFF[262]) );
  XOR U1642 ( .A(B[262]), .B(A[262]), .Z(n1642) );
  XOR U1643 ( .A(n1643), .B(n1644), .Z(DIFF[261]) );
  XOR U1644 ( .A(B[261]), .B(A[261]), .Z(n1644) );
  XOR U1645 ( .A(n1645), .B(n1646), .Z(DIFF[260]) );
  XOR U1646 ( .A(B[260]), .B(A[260]), .Z(n1646) );
  XOR U1647 ( .A(n1647), .B(n1648), .Z(DIFF[25]) );
  XOR U1648 ( .A(B[25]), .B(A[25]), .Z(n1648) );
  XOR U1649 ( .A(n1649), .B(n1650), .Z(DIFF[259]) );
  XOR U1650 ( .A(B[259]), .B(A[259]), .Z(n1650) );
  XOR U1651 ( .A(n1651), .B(n1652), .Z(DIFF[258]) );
  XOR U1652 ( .A(B[258]), .B(A[258]), .Z(n1652) );
  XOR U1653 ( .A(n1653), .B(n1654), .Z(DIFF[257]) );
  XOR U1654 ( .A(B[257]), .B(A[257]), .Z(n1654) );
  XOR U1655 ( .A(n1655), .B(n1656), .Z(DIFF[256]) );
  XOR U1656 ( .A(B[256]), .B(A[256]), .Z(n1656) );
  XOR U1657 ( .A(n1657), .B(n1658), .Z(DIFF[255]) );
  XOR U1658 ( .A(B[255]), .B(A[255]), .Z(n1658) );
  XOR U1659 ( .A(n1659), .B(n1660), .Z(DIFF[254]) );
  XOR U1660 ( .A(B[254]), .B(A[254]), .Z(n1660) );
  XOR U1661 ( .A(n1661), .B(n1662), .Z(DIFF[253]) );
  XOR U1662 ( .A(B[253]), .B(A[253]), .Z(n1662) );
  XOR U1663 ( .A(n1663), .B(n1664), .Z(DIFF[252]) );
  XOR U1664 ( .A(B[252]), .B(A[252]), .Z(n1664) );
  XOR U1665 ( .A(n1665), .B(n1666), .Z(DIFF[251]) );
  XOR U1666 ( .A(B[251]), .B(A[251]), .Z(n1666) );
  XOR U1667 ( .A(n1667), .B(n1668), .Z(DIFF[250]) );
  XOR U1668 ( .A(B[250]), .B(A[250]), .Z(n1668) );
  XOR U1669 ( .A(n1669), .B(n1670), .Z(DIFF[24]) );
  XOR U1670 ( .A(B[24]), .B(A[24]), .Z(n1670) );
  XOR U1671 ( .A(n1671), .B(n1672), .Z(DIFF[249]) );
  XOR U1672 ( .A(B[249]), .B(A[249]), .Z(n1672) );
  XOR U1673 ( .A(n1673), .B(n1674), .Z(DIFF[248]) );
  XOR U1674 ( .A(B[248]), .B(A[248]), .Z(n1674) );
  XOR U1675 ( .A(n1675), .B(n1676), .Z(DIFF[247]) );
  XOR U1676 ( .A(B[247]), .B(A[247]), .Z(n1676) );
  XOR U1677 ( .A(n1677), .B(n1678), .Z(DIFF[246]) );
  XOR U1678 ( .A(B[246]), .B(A[246]), .Z(n1678) );
  XOR U1679 ( .A(n1679), .B(n1680), .Z(DIFF[245]) );
  XOR U1680 ( .A(B[245]), .B(A[245]), .Z(n1680) );
  XOR U1681 ( .A(n1681), .B(n1682), .Z(DIFF[244]) );
  XOR U1682 ( .A(B[244]), .B(A[244]), .Z(n1682) );
  XOR U1683 ( .A(n1683), .B(n1684), .Z(DIFF[243]) );
  XOR U1684 ( .A(B[243]), .B(A[243]), .Z(n1684) );
  XOR U1685 ( .A(n1685), .B(n1686), .Z(DIFF[242]) );
  XOR U1686 ( .A(B[242]), .B(A[242]), .Z(n1686) );
  XOR U1687 ( .A(n1687), .B(n1688), .Z(DIFF[241]) );
  XOR U1688 ( .A(B[241]), .B(A[241]), .Z(n1688) );
  XOR U1689 ( .A(n1689), .B(n1690), .Z(DIFF[240]) );
  XOR U1690 ( .A(B[240]), .B(A[240]), .Z(n1690) );
  XOR U1691 ( .A(n1691), .B(n1692), .Z(DIFF[23]) );
  XOR U1692 ( .A(B[23]), .B(A[23]), .Z(n1692) );
  XOR U1693 ( .A(n1693), .B(n1694), .Z(DIFF[239]) );
  XOR U1694 ( .A(B[239]), .B(A[239]), .Z(n1694) );
  XOR U1695 ( .A(n1695), .B(n1696), .Z(DIFF[238]) );
  XOR U1696 ( .A(B[238]), .B(A[238]), .Z(n1696) );
  XOR U1697 ( .A(n1697), .B(n1698), .Z(DIFF[237]) );
  XOR U1698 ( .A(B[237]), .B(A[237]), .Z(n1698) );
  XOR U1699 ( .A(n1699), .B(n1700), .Z(DIFF[236]) );
  XOR U1700 ( .A(B[236]), .B(A[236]), .Z(n1700) );
  XOR U1701 ( .A(n1701), .B(n1702), .Z(DIFF[235]) );
  XOR U1702 ( .A(B[235]), .B(A[235]), .Z(n1702) );
  XOR U1703 ( .A(n1703), .B(n1704), .Z(DIFF[234]) );
  XOR U1704 ( .A(B[234]), .B(A[234]), .Z(n1704) );
  XOR U1705 ( .A(n1705), .B(n1706), .Z(DIFF[233]) );
  XOR U1706 ( .A(B[233]), .B(A[233]), .Z(n1706) );
  XOR U1707 ( .A(n1707), .B(n1708), .Z(DIFF[232]) );
  XOR U1708 ( .A(B[232]), .B(A[232]), .Z(n1708) );
  XOR U1709 ( .A(n1709), .B(n1710), .Z(DIFF[231]) );
  XOR U1710 ( .A(B[231]), .B(A[231]), .Z(n1710) );
  XOR U1711 ( .A(n1711), .B(n1712), .Z(DIFF[230]) );
  XOR U1712 ( .A(B[230]), .B(A[230]), .Z(n1712) );
  XOR U1713 ( .A(n1713), .B(n1714), .Z(DIFF[22]) );
  XOR U1714 ( .A(B[22]), .B(A[22]), .Z(n1714) );
  XOR U1715 ( .A(n1715), .B(n1716), .Z(DIFF[229]) );
  XOR U1716 ( .A(B[229]), .B(A[229]), .Z(n1716) );
  XOR U1717 ( .A(n1717), .B(n1718), .Z(DIFF[228]) );
  XOR U1718 ( .A(B[228]), .B(A[228]), .Z(n1718) );
  XOR U1719 ( .A(n1719), .B(n1720), .Z(DIFF[227]) );
  XOR U1720 ( .A(B[227]), .B(A[227]), .Z(n1720) );
  XOR U1721 ( .A(n1721), .B(n1722), .Z(DIFF[226]) );
  XOR U1722 ( .A(B[226]), .B(A[226]), .Z(n1722) );
  XOR U1723 ( .A(n1723), .B(n1724), .Z(DIFF[225]) );
  XOR U1724 ( .A(B[225]), .B(A[225]), .Z(n1724) );
  XOR U1725 ( .A(n1725), .B(n1726), .Z(DIFF[224]) );
  XOR U1726 ( .A(B[224]), .B(A[224]), .Z(n1726) );
  XOR U1727 ( .A(n1727), .B(n1728), .Z(DIFF[223]) );
  XOR U1728 ( .A(B[223]), .B(A[223]), .Z(n1728) );
  XOR U1729 ( .A(n1729), .B(n1730), .Z(DIFF[222]) );
  XOR U1730 ( .A(B[222]), .B(A[222]), .Z(n1730) );
  XOR U1731 ( .A(n1731), .B(n1732), .Z(DIFF[221]) );
  XOR U1732 ( .A(B[221]), .B(A[221]), .Z(n1732) );
  XOR U1733 ( .A(n1733), .B(n1734), .Z(DIFF[220]) );
  XOR U1734 ( .A(B[220]), .B(A[220]), .Z(n1734) );
  XOR U1735 ( .A(n1735), .B(n1736), .Z(DIFF[21]) );
  XOR U1736 ( .A(B[21]), .B(A[21]), .Z(n1736) );
  XOR U1737 ( .A(n1737), .B(n1738), .Z(DIFF[219]) );
  XOR U1738 ( .A(B[219]), .B(A[219]), .Z(n1738) );
  XOR U1739 ( .A(n1739), .B(n1740), .Z(DIFF[218]) );
  XOR U1740 ( .A(B[218]), .B(A[218]), .Z(n1740) );
  XOR U1741 ( .A(n1741), .B(n1742), .Z(DIFF[217]) );
  XOR U1742 ( .A(B[217]), .B(A[217]), .Z(n1742) );
  XOR U1743 ( .A(n1743), .B(n1744), .Z(DIFF[216]) );
  XOR U1744 ( .A(B[216]), .B(A[216]), .Z(n1744) );
  XOR U1745 ( .A(n1745), .B(n1746), .Z(DIFF[215]) );
  XOR U1746 ( .A(B[215]), .B(A[215]), .Z(n1746) );
  XOR U1747 ( .A(n1747), .B(n1748), .Z(DIFF[214]) );
  XOR U1748 ( .A(B[214]), .B(A[214]), .Z(n1748) );
  XOR U1749 ( .A(n1749), .B(n1750), .Z(DIFF[213]) );
  XOR U1750 ( .A(B[213]), .B(A[213]), .Z(n1750) );
  XOR U1751 ( .A(n1751), .B(n1752), .Z(DIFF[212]) );
  XOR U1752 ( .A(B[212]), .B(A[212]), .Z(n1752) );
  XOR U1753 ( .A(n1753), .B(n1754), .Z(DIFF[211]) );
  XOR U1754 ( .A(B[211]), .B(A[211]), .Z(n1754) );
  XOR U1755 ( .A(n1755), .B(n1756), .Z(DIFF[210]) );
  XOR U1756 ( .A(B[210]), .B(A[210]), .Z(n1756) );
  XOR U1757 ( .A(n1757), .B(n1758), .Z(DIFF[20]) );
  XOR U1758 ( .A(B[20]), .B(A[20]), .Z(n1758) );
  XOR U1759 ( .A(n1759), .B(n1760), .Z(DIFF[209]) );
  XOR U1760 ( .A(B[209]), .B(A[209]), .Z(n1760) );
  XOR U1761 ( .A(n1761), .B(n1762), .Z(DIFF[208]) );
  XOR U1762 ( .A(B[208]), .B(A[208]), .Z(n1762) );
  XOR U1763 ( .A(n1763), .B(n1764), .Z(DIFF[207]) );
  XOR U1764 ( .A(B[207]), .B(A[207]), .Z(n1764) );
  XOR U1765 ( .A(n1765), .B(n1766), .Z(DIFF[206]) );
  XOR U1766 ( .A(B[206]), .B(A[206]), .Z(n1766) );
  XOR U1767 ( .A(n1767), .B(n1768), .Z(DIFF[205]) );
  XOR U1768 ( .A(B[205]), .B(A[205]), .Z(n1768) );
  XOR U1769 ( .A(n1769), .B(n1770), .Z(DIFF[204]) );
  XOR U1770 ( .A(B[204]), .B(A[204]), .Z(n1770) );
  XOR U1771 ( .A(n1771), .B(n1772), .Z(DIFF[203]) );
  XOR U1772 ( .A(B[203]), .B(A[203]), .Z(n1772) );
  XOR U1773 ( .A(n1773), .B(n1774), .Z(DIFF[202]) );
  XOR U1774 ( .A(B[202]), .B(A[202]), .Z(n1774) );
  XOR U1775 ( .A(n1775), .B(n1776), .Z(DIFF[201]) );
  XOR U1776 ( .A(B[201]), .B(A[201]), .Z(n1776) );
  XOR U1777 ( .A(n1777), .B(n1778), .Z(DIFF[200]) );
  XOR U1778 ( .A(B[200]), .B(A[200]), .Z(n1778) );
  XOR U1779 ( .A(n2), .B(n1779), .Z(DIFF[1]) );
  XOR U1780 ( .A(B[1]), .B(A[1]), .Z(n1779) );
  XOR U1781 ( .A(n1780), .B(n1781), .Z(DIFF[19]) );
  XOR U1782 ( .A(B[19]), .B(A[19]), .Z(n1781) );
  XOR U1783 ( .A(n1782), .B(n1783), .Z(DIFF[199]) );
  XOR U1784 ( .A(B[199]), .B(A[199]), .Z(n1783) );
  XOR U1785 ( .A(n1784), .B(n1785), .Z(DIFF[198]) );
  XOR U1786 ( .A(B[198]), .B(A[198]), .Z(n1785) );
  XOR U1787 ( .A(n1786), .B(n1787), .Z(DIFF[197]) );
  XOR U1788 ( .A(B[197]), .B(A[197]), .Z(n1787) );
  XOR U1789 ( .A(n1788), .B(n1789), .Z(DIFF[196]) );
  XOR U1790 ( .A(B[196]), .B(A[196]), .Z(n1789) );
  XOR U1791 ( .A(n1790), .B(n1791), .Z(DIFF[195]) );
  XOR U1792 ( .A(B[195]), .B(A[195]), .Z(n1791) );
  XOR U1793 ( .A(n1792), .B(n1793), .Z(DIFF[194]) );
  XOR U1794 ( .A(B[194]), .B(A[194]), .Z(n1793) );
  XOR U1795 ( .A(n1794), .B(n1795), .Z(DIFF[193]) );
  XOR U1796 ( .A(B[193]), .B(A[193]), .Z(n1795) );
  XOR U1797 ( .A(n1796), .B(n1797), .Z(DIFF[192]) );
  XOR U1798 ( .A(B[192]), .B(A[192]), .Z(n1797) );
  XOR U1799 ( .A(n1798), .B(n1799), .Z(DIFF[191]) );
  XOR U1800 ( .A(B[191]), .B(A[191]), .Z(n1799) );
  XOR U1801 ( .A(n1800), .B(n1801), .Z(DIFF[190]) );
  XOR U1802 ( .A(B[190]), .B(A[190]), .Z(n1801) );
  XOR U1803 ( .A(n1802), .B(n1803), .Z(DIFF[18]) );
  XOR U1804 ( .A(B[18]), .B(A[18]), .Z(n1803) );
  XOR U1805 ( .A(n1804), .B(n1805), .Z(DIFF[189]) );
  XOR U1806 ( .A(B[189]), .B(A[189]), .Z(n1805) );
  XOR U1807 ( .A(n1806), .B(n1807), .Z(DIFF[188]) );
  XOR U1808 ( .A(B[188]), .B(A[188]), .Z(n1807) );
  XOR U1809 ( .A(n1808), .B(n1809), .Z(DIFF[187]) );
  XOR U1810 ( .A(B[187]), .B(A[187]), .Z(n1809) );
  XOR U1811 ( .A(n1810), .B(n1811), .Z(DIFF[186]) );
  XOR U1812 ( .A(B[186]), .B(A[186]), .Z(n1811) );
  XOR U1813 ( .A(n1812), .B(n1813), .Z(DIFF[185]) );
  XOR U1814 ( .A(B[185]), .B(A[185]), .Z(n1813) );
  XOR U1815 ( .A(n1814), .B(n1815), .Z(DIFF[184]) );
  XOR U1816 ( .A(B[184]), .B(A[184]), .Z(n1815) );
  XOR U1817 ( .A(n1816), .B(n1817), .Z(DIFF[183]) );
  XOR U1818 ( .A(B[183]), .B(A[183]), .Z(n1817) );
  XOR U1819 ( .A(n1818), .B(n1819), .Z(DIFF[182]) );
  XOR U1820 ( .A(B[182]), .B(A[182]), .Z(n1819) );
  XOR U1821 ( .A(n1820), .B(n1821), .Z(DIFF[181]) );
  XOR U1822 ( .A(B[181]), .B(A[181]), .Z(n1821) );
  XOR U1823 ( .A(n1822), .B(n1823), .Z(DIFF[180]) );
  XOR U1824 ( .A(B[180]), .B(A[180]), .Z(n1823) );
  XOR U1825 ( .A(n1824), .B(n1825), .Z(DIFF[17]) );
  XOR U1826 ( .A(B[17]), .B(A[17]), .Z(n1825) );
  XOR U1827 ( .A(n1826), .B(n1827), .Z(DIFF[179]) );
  XOR U1828 ( .A(B[179]), .B(A[179]), .Z(n1827) );
  XOR U1829 ( .A(n1828), .B(n1829), .Z(DIFF[178]) );
  XOR U1830 ( .A(B[178]), .B(A[178]), .Z(n1829) );
  XOR U1831 ( .A(n1830), .B(n1831), .Z(DIFF[177]) );
  XOR U1832 ( .A(B[177]), .B(A[177]), .Z(n1831) );
  XOR U1833 ( .A(n1832), .B(n1833), .Z(DIFF[176]) );
  XOR U1834 ( .A(B[176]), .B(A[176]), .Z(n1833) );
  XOR U1835 ( .A(n1834), .B(n1835), .Z(DIFF[175]) );
  XOR U1836 ( .A(B[175]), .B(A[175]), .Z(n1835) );
  XOR U1837 ( .A(n1836), .B(n1837), .Z(DIFF[174]) );
  XOR U1838 ( .A(B[174]), .B(A[174]), .Z(n1837) );
  XOR U1839 ( .A(n1838), .B(n1839), .Z(DIFF[173]) );
  XOR U1840 ( .A(B[173]), .B(A[173]), .Z(n1839) );
  XOR U1841 ( .A(n1840), .B(n1841), .Z(DIFF[172]) );
  XOR U1842 ( .A(B[172]), .B(A[172]), .Z(n1841) );
  XOR U1843 ( .A(n1842), .B(n1843), .Z(DIFF[171]) );
  XOR U1844 ( .A(B[171]), .B(A[171]), .Z(n1843) );
  XOR U1845 ( .A(n1844), .B(n1845), .Z(DIFF[170]) );
  XOR U1846 ( .A(B[170]), .B(A[170]), .Z(n1845) );
  XOR U1847 ( .A(n1846), .B(n1847), .Z(DIFF[16]) );
  XOR U1848 ( .A(B[16]), .B(A[16]), .Z(n1847) );
  XOR U1849 ( .A(n1848), .B(n1849), .Z(DIFF[169]) );
  XOR U1850 ( .A(B[169]), .B(A[169]), .Z(n1849) );
  XOR U1851 ( .A(n1850), .B(n1851), .Z(DIFF[168]) );
  XOR U1852 ( .A(B[168]), .B(A[168]), .Z(n1851) );
  XOR U1853 ( .A(n1852), .B(n1853), .Z(DIFF[167]) );
  XOR U1854 ( .A(B[167]), .B(A[167]), .Z(n1853) );
  XOR U1855 ( .A(n1854), .B(n1855), .Z(DIFF[166]) );
  XOR U1856 ( .A(B[166]), .B(A[166]), .Z(n1855) );
  XOR U1857 ( .A(n1856), .B(n1857), .Z(DIFF[165]) );
  XOR U1858 ( .A(B[165]), .B(A[165]), .Z(n1857) );
  XOR U1859 ( .A(n1858), .B(n1859), .Z(DIFF[164]) );
  XOR U1860 ( .A(B[164]), .B(A[164]), .Z(n1859) );
  XOR U1861 ( .A(n1860), .B(n1861), .Z(DIFF[163]) );
  XOR U1862 ( .A(B[163]), .B(A[163]), .Z(n1861) );
  XOR U1863 ( .A(n1862), .B(n1863), .Z(DIFF[162]) );
  XOR U1864 ( .A(B[162]), .B(A[162]), .Z(n1863) );
  XOR U1865 ( .A(n1864), .B(n1865), .Z(DIFF[161]) );
  XOR U1866 ( .A(B[161]), .B(A[161]), .Z(n1865) );
  XOR U1867 ( .A(n1866), .B(n1867), .Z(DIFF[160]) );
  XOR U1868 ( .A(B[160]), .B(A[160]), .Z(n1867) );
  XOR U1869 ( .A(n1868), .B(n1869), .Z(DIFF[15]) );
  XOR U1870 ( .A(B[15]), .B(A[15]), .Z(n1869) );
  XOR U1871 ( .A(n1870), .B(n1871), .Z(DIFF[159]) );
  XOR U1872 ( .A(B[159]), .B(A[159]), .Z(n1871) );
  XOR U1873 ( .A(n1872), .B(n1873), .Z(DIFF[158]) );
  XOR U1874 ( .A(B[158]), .B(A[158]), .Z(n1873) );
  XOR U1875 ( .A(n1874), .B(n1875), .Z(DIFF[157]) );
  XOR U1876 ( .A(B[157]), .B(A[157]), .Z(n1875) );
  XOR U1877 ( .A(n1876), .B(n1877), .Z(DIFF[156]) );
  XOR U1878 ( .A(B[156]), .B(A[156]), .Z(n1877) );
  XOR U1879 ( .A(n1878), .B(n1879), .Z(DIFF[155]) );
  XOR U1880 ( .A(B[155]), .B(A[155]), .Z(n1879) );
  XOR U1881 ( .A(n1880), .B(n1881), .Z(DIFF[154]) );
  XOR U1882 ( .A(B[154]), .B(A[154]), .Z(n1881) );
  XOR U1883 ( .A(n1882), .B(n1883), .Z(DIFF[153]) );
  XOR U1884 ( .A(B[153]), .B(A[153]), .Z(n1883) );
  XOR U1885 ( .A(n1884), .B(n1885), .Z(DIFF[152]) );
  XOR U1886 ( .A(B[152]), .B(A[152]), .Z(n1885) );
  XOR U1887 ( .A(n1886), .B(n1887), .Z(DIFF[151]) );
  XOR U1888 ( .A(B[151]), .B(A[151]), .Z(n1887) );
  XOR U1889 ( .A(n1888), .B(n1889), .Z(DIFF[150]) );
  XOR U1890 ( .A(B[150]), .B(A[150]), .Z(n1889) );
  XOR U1891 ( .A(n1890), .B(n1891), .Z(DIFF[14]) );
  XOR U1892 ( .A(B[14]), .B(A[14]), .Z(n1891) );
  XOR U1893 ( .A(n1892), .B(n1893), .Z(DIFF[149]) );
  XOR U1894 ( .A(B[149]), .B(A[149]), .Z(n1893) );
  XOR U1895 ( .A(n1894), .B(n1895), .Z(DIFF[148]) );
  XOR U1896 ( .A(B[148]), .B(A[148]), .Z(n1895) );
  XOR U1897 ( .A(n1896), .B(n1897), .Z(DIFF[147]) );
  XOR U1898 ( .A(B[147]), .B(A[147]), .Z(n1897) );
  XOR U1899 ( .A(n1898), .B(n1899), .Z(DIFF[146]) );
  XOR U1900 ( .A(B[146]), .B(A[146]), .Z(n1899) );
  XOR U1901 ( .A(n1900), .B(n1901), .Z(DIFF[145]) );
  XOR U1902 ( .A(B[145]), .B(A[145]), .Z(n1901) );
  XOR U1903 ( .A(n1902), .B(n1903), .Z(DIFF[144]) );
  XOR U1904 ( .A(B[144]), .B(A[144]), .Z(n1903) );
  XOR U1905 ( .A(n1904), .B(n1905), .Z(DIFF[143]) );
  XOR U1906 ( .A(B[143]), .B(A[143]), .Z(n1905) );
  XOR U1907 ( .A(n1906), .B(n1907), .Z(DIFF[142]) );
  XOR U1908 ( .A(B[142]), .B(A[142]), .Z(n1907) );
  XOR U1909 ( .A(n1908), .B(n1909), .Z(DIFF[141]) );
  XOR U1910 ( .A(B[141]), .B(A[141]), .Z(n1909) );
  XOR U1911 ( .A(n1910), .B(n1911), .Z(DIFF[140]) );
  XOR U1912 ( .A(B[140]), .B(A[140]), .Z(n1911) );
  XOR U1913 ( .A(n1912), .B(n1913), .Z(DIFF[13]) );
  XOR U1914 ( .A(B[13]), .B(A[13]), .Z(n1913) );
  XOR U1915 ( .A(n1914), .B(n1915), .Z(DIFF[139]) );
  XOR U1916 ( .A(B[139]), .B(A[139]), .Z(n1915) );
  XOR U1917 ( .A(n1916), .B(n1917), .Z(DIFF[138]) );
  XOR U1918 ( .A(B[138]), .B(A[138]), .Z(n1917) );
  XOR U1919 ( .A(n1918), .B(n1919), .Z(DIFF[137]) );
  XOR U1920 ( .A(B[137]), .B(A[137]), .Z(n1919) );
  XOR U1921 ( .A(n1920), .B(n1921), .Z(DIFF[136]) );
  XOR U1922 ( .A(B[136]), .B(A[136]), .Z(n1921) );
  XOR U1923 ( .A(n1922), .B(n1923), .Z(DIFF[135]) );
  XOR U1924 ( .A(B[135]), .B(A[135]), .Z(n1923) );
  XOR U1925 ( .A(n1924), .B(n1925), .Z(DIFF[134]) );
  XOR U1926 ( .A(B[134]), .B(A[134]), .Z(n1925) );
  XOR U1927 ( .A(n1926), .B(n1927), .Z(DIFF[133]) );
  XOR U1928 ( .A(B[133]), .B(A[133]), .Z(n1927) );
  XOR U1929 ( .A(n1928), .B(n1929), .Z(DIFF[132]) );
  XOR U1930 ( .A(B[132]), .B(A[132]), .Z(n1929) );
  XOR U1931 ( .A(n1930), .B(n1931), .Z(DIFF[131]) );
  XOR U1932 ( .A(B[131]), .B(A[131]), .Z(n1931) );
  XOR U1933 ( .A(n1932), .B(n1933), .Z(DIFF[130]) );
  XOR U1934 ( .A(B[130]), .B(A[130]), .Z(n1933) );
  XOR U1935 ( .A(n1934), .B(n1935), .Z(DIFF[12]) );
  XOR U1936 ( .A(B[12]), .B(A[12]), .Z(n1935) );
  XOR U1937 ( .A(n1936), .B(n1937), .Z(DIFF[129]) );
  XOR U1938 ( .A(B[129]), .B(A[129]), .Z(n1937) );
  XOR U1939 ( .A(n1938), .B(n1939), .Z(DIFF[128]) );
  XOR U1940 ( .A(B[128]), .B(A[128]), .Z(n1939) );
  XOR U1941 ( .A(n1940), .B(n1941), .Z(DIFF[127]) );
  XOR U1942 ( .A(B[127]), .B(A[127]), .Z(n1941) );
  XOR U1943 ( .A(n1942), .B(n1943), .Z(DIFF[126]) );
  XOR U1944 ( .A(B[126]), .B(A[126]), .Z(n1943) );
  XOR U1945 ( .A(n1944), .B(n1945), .Z(DIFF[125]) );
  XOR U1946 ( .A(B[125]), .B(A[125]), .Z(n1945) );
  XOR U1947 ( .A(n1946), .B(n1947), .Z(DIFF[124]) );
  XOR U1948 ( .A(B[124]), .B(A[124]), .Z(n1947) );
  XOR U1949 ( .A(n1948), .B(n1949), .Z(DIFF[123]) );
  XOR U1950 ( .A(B[123]), .B(A[123]), .Z(n1949) );
  XOR U1951 ( .A(n1950), .B(n1951), .Z(DIFF[122]) );
  XOR U1952 ( .A(B[122]), .B(A[122]), .Z(n1951) );
  XOR U1953 ( .A(n1952), .B(n1953), .Z(DIFF[121]) );
  XOR U1954 ( .A(B[121]), .B(A[121]), .Z(n1953) );
  XOR U1955 ( .A(n1954), .B(n1955), .Z(DIFF[120]) );
  XOR U1956 ( .A(B[120]), .B(A[120]), .Z(n1955) );
  XOR U1957 ( .A(n1956), .B(n1957), .Z(DIFF[11]) );
  XOR U1958 ( .A(B[11]), .B(A[11]), .Z(n1957) );
  XOR U1959 ( .A(n1958), .B(n1959), .Z(DIFF[119]) );
  XOR U1960 ( .A(B[119]), .B(A[119]), .Z(n1959) );
  XOR U1961 ( .A(n1960), .B(n1961), .Z(DIFF[118]) );
  XOR U1962 ( .A(B[118]), .B(A[118]), .Z(n1961) );
  XOR U1963 ( .A(n1962), .B(n1963), .Z(DIFF[117]) );
  XOR U1964 ( .A(B[117]), .B(A[117]), .Z(n1963) );
  XOR U1965 ( .A(n1964), .B(n1965), .Z(DIFF[116]) );
  XOR U1966 ( .A(B[116]), .B(A[116]), .Z(n1965) );
  XOR U1967 ( .A(n1966), .B(n1967), .Z(DIFF[115]) );
  XOR U1968 ( .A(B[115]), .B(A[115]), .Z(n1967) );
  XOR U1969 ( .A(n1968), .B(n1969), .Z(DIFF[114]) );
  XOR U1970 ( .A(B[114]), .B(A[114]), .Z(n1969) );
  XOR U1971 ( .A(n1970), .B(n1971), .Z(DIFF[113]) );
  XOR U1972 ( .A(B[113]), .B(A[113]), .Z(n1971) );
  XOR U1973 ( .A(n1972), .B(n1973), .Z(DIFF[112]) );
  XOR U1974 ( .A(B[112]), .B(A[112]), .Z(n1973) );
  XOR U1975 ( .A(n1974), .B(n1975), .Z(DIFF[111]) );
  XOR U1976 ( .A(B[111]), .B(A[111]), .Z(n1975) );
  XOR U1977 ( .A(n1976), .B(n1977), .Z(DIFF[110]) );
  XOR U1978 ( .A(B[110]), .B(A[110]), .Z(n1977) );
  XOR U1979 ( .A(n1978), .B(n1979), .Z(DIFF[10]) );
  XOR U1980 ( .A(B[10]), .B(A[10]), .Z(n1979) );
  XOR U1981 ( .A(n1980), .B(n1981), .Z(DIFF[109]) );
  XOR U1982 ( .A(B[109]), .B(A[109]), .Z(n1981) );
  XOR U1983 ( .A(n1982), .B(n1983), .Z(DIFF[108]) );
  XOR U1984 ( .A(B[108]), .B(A[108]), .Z(n1983) );
  XOR U1985 ( .A(n1984), .B(n1985), .Z(DIFF[107]) );
  XOR U1986 ( .A(B[107]), .B(A[107]), .Z(n1985) );
  XOR U1987 ( .A(n1986), .B(n1987), .Z(DIFF[106]) );
  XOR U1988 ( .A(B[106]), .B(A[106]), .Z(n1987) );
  XOR U1989 ( .A(n1988), .B(n1989), .Z(DIFF[105]) );
  XOR U1990 ( .A(B[105]), .B(A[105]), .Z(n1989) );
  XOR U1991 ( .A(n1990), .B(n1991), .Z(DIFF[104]) );
  XOR U1992 ( .A(B[104]), .B(A[104]), .Z(n1991) );
  XOR U1993 ( .A(n1992), .B(n1993), .Z(DIFF[103]) );
  XOR U1994 ( .A(B[103]), .B(A[103]), .Z(n1993) );
  XOR U1995 ( .A(n1994), .B(n1995), .Z(DIFF[102]) );
  XOR U1996 ( .A(B[102]), .B(A[102]), .Z(n1995) );
  XOR U1997 ( .A(A[1025]), .B(n1996), .Z(DIFF[1025]) );
  ANDN U1998 ( .B(n1997), .A(A[1024]), .Z(n1996) );
  XOR U1999 ( .A(A[1024]), .B(n1997), .Z(DIFF[1024]) );
  AND U2000 ( .A(n1998), .B(n1999), .Z(n1997) );
  NANDN U2001 ( .A(B[1023]), .B(n2000), .Z(n1999) );
  NANDN U2002 ( .A(A[1023]), .B(n2001), .Z(n2000) );
  NANDN U2003 ( .A(n2001), .B(A[1023]), .Z(n1998) );
  XOR U2004 ( .A(n2001), .B(n2002), .Z(DIFF[1023]) );
  XOR U2005 ( .A(B[1023]), .B(A[1023]), .Z(n2002) );
  AND U2006 ( .A(n2003), .B(n2004), .Z(n2001) );
  NANDN U2007 ( .A(B[1022]), .B(n2005), .Z(n2004) );
  NANDN U2008 ( .A(A[1022]), .B(n2006), .Z(n2005) );
  NANDN U2009 ( .A(n2006), .B(A[1022]), .Z(n2003) );
  XOR U2010 ( .A(n2006), .B(n2007), .Z(DIFF[1022]) );
  XOR U2011 ( .A(B[1022]), .B(A[1022]), .Z(n2007) );
  AND U2012 ( .A(n2008), .B(n2009), .Z(n2006) );
  NANDN U2013 ( .A(B[1021]), .B(n2010), .Z(n2009) );
  NANDN U2014 ( .A(A[1021]), .B(n2011), .Z(n2010) );
  NANDN U2015 ( .A(n2011), .B(A[1021]), .Z(n2008) );
  XOR U2016 ( .A(n2011), .B(n2012), .Z(DIFF[1021]) );
  XOR U2017 ( .A(B[1021]), .B(A[1021]), .Z(n2012) );
  AND U2018 ( .A(n2013), .B(n2014), .Z(n2011) );
  NANDN U2019 ( .A(B[1020]), .B(n2015), .Z(n2014) );
  NANDN U2020 ( .A(A[1020]), .B(n2016), .Z(n2015) );
  NANDN U2021 ( .A(n2016), .B(A[1020]), .Z(n2013) );
  XOR U2022 ( .A(n2016), .B(n2017), .Z(DIFF[1020]) );
  XOR U2023 ( .A(B[1020]), .B(A[1020]), .Z(n2017) );
  AND U2024 ( .A(n2018), .B(n2019), .Z(n2016) );
  NANDN U2025 ( .A(B[1019]), .B(n2020), .Z(n2019) );
  NANDN U2026 ( .A(A[1019]), .B(n2021), .Z(n2020) );
  NANDN U2027 ( .A(n2021), .B(A[1019]), .Z(n2018) );
  XOR U2028 ( .A(n2022), .B(n2023), .Z(DIFF[101]) );
  XOR U2029 ( .A(B[101]), .B(A[101]), .Z(n2023) );
  XOR U2030 ( .A(n2021), .B(n2024), .Z(DIFF[1019]) );
  XOR U2031 ( .A(B[1019]), .B(A[1019]), .Z(n2024) );
  AND U2032 ( .A(n2025), .B(n2026), .Z(n2021) );
  NANDN U2033 ( .A(B[1018]), .B(n2027), .Z(n2026) );
  NANDN U2034 ( .A(A[1018]), .B(n2028), .Z(n2027) );
  NANDN U2035 ( .A(n2028), .B(A[1018]), .Z(n2025) );
  XOR U2036 ( .A(n2028), .B(n2029), .Z(DIFF[1018]) );
  XOR U2037 ( .A(B[1018]), .B(A[1018]), .Z(n2029) );
  AND U2038 ( .A(n2030), .B(n2031), .Z(n2028) );
  NANDN U2039 ( .A(B[1017]), .B(n2032), .Z(n2031) );
  NANDN U2040 ( .A(A[1017]), .B(n2033), .Z(n2032) );
  NANDN U2041 ( .A(n2033), .B(A[1017]), .Z(n2030) );
  XOR U2042 ( .A(n2033), .B(n2034), .Z(DIFF[1017]) );
  XOR U2043 ( .A(B[1017]), .B(A[1017]), .Z(n2034) );
  AND U2044 ( .A(n2035), .B(n2036), .Z(n2033) );
  NANDN U2045 ( .A(B[1016]), .B(n2037), .Z(n2036) );
  NANDN U2046 ( .A(A[1016]), .B(n2038), .Z(n2037) );
  NANDN U2047 ( .A(n2038), .B(A[1016]), .Z(n2035) );
  XOR U2048 ( .A(n2038), .B(n2039), .Z(DIFF[1016]) );
  XOR U2049 ( .A(B[1016]), .B(A[1016]), .Z(n2039) );
  AND U2050 ( .A(n2040), .B(n2041), .Z(n2038) );
  NANDN U2051 ( .A(B[1015]), .B(n2042), .Z(n2041) );
  NANDN U2052 ( .A(A[1015]), .B(n2043), .Z(n2042) );
  NANDN U2053 ( .A(n2043), .B(A[1015]), .Z(n2040) );
  XOR U2054 ( .A(n2043), .B(n2044), .Z(DIFF[1015]) );
  XOR U2055 ( .A(B[1015]), .B(A[1015]), .Z(n2044) );
  AND U2056 ( .A(n2045), .B(n2046), .Z(n2043) );
  NANDN U2057 ( .A(B[1014]), .B(n2047), .Z(n2046) );
  NANDN U2058 ( .A(A[1014]), .B(n2048), .Z(n2047) );
  NANDN U2059 ( .A(n2048), .B(A[1014]), .Z(n2045) );
  XOR U2060 ( .A(n2048), .B(n2049), .Z(DIFF[1014]) );
  XOR U2061 ( .A(B[1014]), .B(A[1014]), .Z(n2049) );
  AND U2062 ( .A(n2050), .B(n2051), .Z(n2048) );
  NANDN U2063 ( .A(B[1013]), .B(n2052), .Z(n2051) );
  NANDN U2064 ( .A(A[1013]), .B(n2053), .Z(n2052) );
  NANDN U2065 ( .A(n2053), .B(A[1013]), .Z(n2050) );
  XOR U2066 ( .A(n2053), .B(n2054), .Z(DIFF[1013]) );
  XOR U2067 ( .A(B[1013]), .B(A[1013]), .Z(n2054) );
  AND U2068 ( .A(n2055), .B(n2056), .Z(n2053) );
  NANDN U2069 ( .A(B[1012]), .B(n2057), .Z(n2056) );
  NANDN U2070 ( .A(A[1012]), .B(n2058), .Z(n2057) );
  NANDN U2071 ( .A(n2058), .B(A[1012]), .Z(n2055) );
  XOR U2072 ( .A(n2058), .B(n2059), .Z(DIFF[1012]) );
  XOR U2073 ( .A(B[1012]), .B(A[1012]), .Z(n2059) );
  AND U2074 ( .A(n2060), .B(n2061), .Z(n2058) );
  NANDN U2075 ( .A(B[1011]), .B(n2062), .Z(n2061) );
  NANDN U2076 ( .A(A[1011]), .B(n2063), .Z(n2062) );
  NANDN U2077 ( .A(n2063), .B(A[1011]), .Z(n2060) );
  XOR U2078 ( .A(n2063), .B(n2064), .Z(DIFF[1011]) );
  XOR U2079 ( .A(B[1011]), .B(A[1011]), .Z(n2064) );
  AND U2080 ( .A(n2065), .B(n2066), .Z(n2063) );
  NANDN U2081 ( .A(B[1010]), .B(n2067), .Z(n2066) );
  NANDN U2082 ( .A(A[1010]), .B(n2068), .Z(n2067) );
  NANDN U2083 ( .A(n2068), .B(A[1010]), .Z(n2065) );
  XOR U2084 ( .A(n2068), .B(n2069), .Z(DIFF[1010]) );
  XOR U2085 ( .A(B[1010]), .B(A[1010]), .Z(n2069) );
  AND U2086 ( .A(n2070), .B(n2071), .Z(n2068) );
  NANDN U2087 ( .A(B[1009]), .B(n2072), .Z(n2071) );
  NANDN U2088 ( .A(A[1009]), .B(n2073), .Z(n2072) );
  NANDN U2089 ( .A(n2073), .B(A[1009]), .Z(n2070) );
  XOR U2090 ( .A(n2074), .B(n2075), .Z(DIFF[100]) );
  XOR U2091 ( .A(B[100]), .B(A[100]), .Z(n2075) );
  XOR U2092 ( .A(n2073), .B(n2076), .Z(DIFF[1009]) );
  XOR U2093 ( .A(B[1009]), .B(A[1009]), .Z(n2076) );
  AND U2094 ( .A(n2077), .B(n2078), .Z(n2073) );
  NANDN U2095 ( .A(B[1008]), .B(n2079), .Z(n2078) );
  NANDN U2096 ( .A(A[1008]), .B(n2080), .Z(n2079) );
  NANDN U2097 ( .A(n2080), .B(A[1008]), .Z(n2077) );
  XOR U2098 ( .A(n2080), .B(n2081), .Z(DIFF[1008]) );
  XOR U2099 ( .A(B[1008]), .B(A[1008]), .Z(n2081) );
  AND U2100 ( .A(n2082), .B(n2083), .Z(n2080) );
  NANDN U2101 ( .A(B[1007]), .B(n2084), .Z(n2083) );
  NANDN U2102 ( .A(A[1007]), .B(n2085), .Z(n2084) );
  NANDN U2103 ( .A(n2085), .B(A[1007]), .Z(n2082) );
  XOR U2104 ( .A(n2085), .B(n2086), .Z(DIFF[1007]) );
  XOR U2105 ( .A(B[1007]), .B(A[1007]), .Z(n2086) );
  AND U2106 ( .A(n2087), .B(n2088), .Z(n2085) );
  NANDN U2107 ( .A(B[1006]), .B(n2089), .Z(n2088) );
  NANDN U2108 ( .A(A[1006]), .B(n2090), .Z(n2089) );
  NANDN U2109 ( .A(n2090), .B(A[1006]), .Z(n2087) );
  XOR U2110 ( .A(n2090), .B(n2091), .Z(DIFF[1006]) );
  XOR U2111 ( .A(B[1006]), .B(A[1006]), .Z(n2091) );
  AND U2112 ( .A(n2092), .B(n2093), .Z(n2090) );
  NANDN U2113 ( .A(B[1005]), .B(n2094), .Z(n2093) );
  NANDN U2114 ( .A(A[1005]), .B(n2095), .Z(n2094) );
  NANDN U2115 ( .A(n2095), .B(A[1005]), .Z(n2092) );
  XOR U2116 ( .A(n2095), .B(n2096), .Z(DIFF[1005]) );
  XOR U2117 ( .A(B[1005]), .B(A[1005]), .Z(n2096) );
  AND U2118 ( .A(n2097), .B(n2098), .Z(n2095) );
  NANDN U2119 ( .A(B[1004]), .B(n2099), .Z(n2098) );
  NANDN U2120 ( .A(A[1004]), .B(n2100), .Z(n2099) );
  NANDN U2121 ( .A(n2100), .B(A[1004]), .Z(n2097) );
  XOR U2122 ( .A(n2100), .B(n2101), .Z(DIFF[1004]) );
  XOR U2123 ( .A(B[1004]), .B(A[1004]), .Z(n2101) );
  AND U2124 ( .A(n2102), .B(n2103), .Z(n2100) );
  NANDN U2125 ( .A(B[1003]), .B(n2104), .Z(n2103) );
  NANDN U2126 ( .A(A[1003]), .B(n2105), .Z(n2104) );
  NANDN U2127 ( .A(n2105), .B(A[1003]), .Z(n2102) );
  XOR U2128 ( .A(n2105), .B(n2106), .Z(DIFF[1003]) );
  XOR U2129 ( .A(B[1003]), .B(A[1003]), .Z(n2106) );
  AND U2130 ( .A(n2107), .B(n2108), .Z(n2105) );
  NANDN U2131 ( .A(B[1002]), .B(n2109), .Z(n2108) );
  NANDN U2132 ( .A(A[1002]), .B(n2110), .Z(n2109) );
  NANDN U2133 ( .A(n2110), .B(A[1002]), .Z(n2107) );
  XOR U2134 ( .A(n2110), .B(n2111), .Z(DIFF[1002]) );
  XOR U2135 ( .A(B[1002]), .B(A[1002]), .Z(n2111) );
  AND U2136 ( .A(n2112), .B(n2113), .Z(n2110) );
  NANDN U2137 ( .A(B[1001]), .B(n2114), .Z(n2113) );
  NANDN U2138 ( .A(A[1001]), .B(n2115), .Z(n2114) );
  NANDN U2139 ( .A(n2115), .B(A[1001]), .Z(n2112) );
  XOR U2140 ( .A(n2115), .B(n2116), .Z(DIFF[1001]) );
  XOR U2141 ( .A(B[1001]), .B(A[1001]), .Z(n2116) );
  AND U2142 ( .A(n2117), .B(n2118), .Z(n2115) );
  NANDN U2143 ( .A(B[1000]), .B(n2119), .Z(n2118) );
  NANDN U2144 ( .A(A[1000]), .B(n2120), .Z(n2119) );
  NANDN U2145 ( .A(n2120), .B(A[1000]), .Z(n2117) );
  XOR U2146 ( .A(n2120), .B(n2121), .Z(DIFF[1000]) );
  XOR U2147 ( .A(B[1000]), .B(A[1000]), .Z(n2121) );
  AND U2148 ( .A(n2122), .B(n2123), .Z(n2120) );
  NANDN U2149 ( .A(B[999]), .B(n2124), .Z(n2123) );
  OR U2150 ( .A(n7), .B(A[999]), .Z(n2124) );
  NAND U2151 ( .A(A[999]), .B(n7), .Z(n2122) );
  NAND U2152 ( .A(n2125), .B(n2126), .Z(n7) );
  NANDN U2153 ( .A(B[998]), .B(n2127), .Z(n2126) );
  NANDN U2154 ( .A(A[998]), .B(n9), .Z(n2127) );
  NANDN U2155 ( .A(n9), .B(A[998]), .Z(n2125) );
  AND U2156 ( .A(n2128), .B(n2129), .Z(n9) );
  NANDN U2157 ( .A(B[997]), .B(n2130), .Z(n2129) );
  NANDN U2158 ( .A(A[997]), .B(n11), .Z(n2130) );
  NANDN U2159 ( .A(n11), .B(A[997]), .Z(n2128) );
  AND U2160 ( .A(n2131), .B(n2132), .Z(n11) );
  NANDN U2161 ( .A(B[996]), .B(n2133), .Z(n2132) );
  NANDN U2162 ( .A(A[996]), .B(n13), .Z(n2133) );
  NANDN U2163 ( .A(n13), .B(A[996]), .Z(n2131) );
  AND U2164 ( .A(n2134), .B(n2135), .Z(n13) );
  NANDN U2165 ( .A(B[995]), .B(n2136), .Z(n2135) );
  NANDN U2166 ( .A(A[995]), .B(n15), .Z(n2136) );
  NANDN U2167 ( .A(n15), .B(A[995]), .Z(n2134) );
  AND U2168 ( .A(n2137), .B(n2138), .Z(n15) );
  NANDN U2169 ( .A(B[994]), .B(n2139), .Z(n2138) );
  NANDN U2170 ( .A(A[994]), .B(n17), .Z(n2139) );
  NANDN U2171 ( .A(n17), .B(A[994]), .Z(n2137) );
  AND U2172 ( .A(n2140), .B(n2141), .Z(n17) );
  NANDN U2173 ( .A(B[993]), .B(n2142), .Z(n2141) );
  NANDN U2174 ( .A(A[993]), .B(n19), .Z(n2142) );
  NANDN U2175 ( .A(n19), .B(A[993]), .Z(n2140) );
  AND U2176 ( .A(n2143), .B(n2144), .Z(n19) );
  NANDN U2177 ( .A(B[992]), .B(n2145), .Z(n2144) );
  NANDN U2178 ( .A(A[992]), .B(n21), .Z(n2145) );
  NANDN U2179 ( .A(n21), .B(A[992]), .Z(n2143) );
  AND U2180 ( .A(n2146), .B(n2147), .Z(n21) );
  NANDN U2181 ( .A(B[991]), .B(n2148), .Z(n2147) );
  NANDN U2182 ( .A(A[991]), .B(n23), .Z(n2148) );
  NANDN U2183 ( .A(n23), .B(A[991]), .Z(n2146) );
  AND U2184 ( .A(n2149), .B(n2150), .Z(n23) );
  NANDN U2185 ( .A(B[990]), .B(n2151), .Z(n2150) );
  NANDN U2186 ( .A(A[990]), .B(n25), .Z(n2151) );
  NANDN U2187 ( .A(n25), .B(A[990]), .Z(n2149) );
  AND U2188 ( .A(n2152), .B(n2153), .Z(n25) );
  NANDN U2189 ( .A(B[989]), .B(n2154), .Z(n2153) );
  NANDN U2190 ( .A(A[989]), .B(n29), .Z(n2154) );
  NANDN U2191 ( .A(n29), .B(A[989]), .Z(n2152) );
  AND U2192 ( .A(n2155), .B(n2156), .Z(n29) );
  NANDN U2193 ( .A(B[988]), .B(n2157), .Z(n2156) );
  NANDN U2194 ( .A(A[988]), .B(n31), .Z(n2157) );
  NANDN U2195 ( .A(n31), .B(A[988]), .Z(n2155) );
  AND U2196 ( .A(n2158), .B(n2159), .Z(n31) );
  NANDN U2197 ( .A(B[987]), .B(n2160), .Z(n2159) );
  NANDN U2198 ( .A(A[987]), .B(n33), .Z(n2160) );
  NANDN U2199 ( .A(n33), .B(A[987]), .Z(n2158) );
  AND U2200 ( .A(n2161), .B(n2162), .Z(n33) );
  NANDN U2201 ( .A(B[986]), .B(n2163), .Z(n2162) );
  NANDN U2202 ( .A(A[986]), .B(n35), .Z(n2163) );
  NANDN U2203 ( .A(n35), .B(A[986]), .Z(n2161) );
  AND U2204 ( .A(n2164), .B(n2165), .Z(n35) );
  NANDN U2205 ( .A(B[985]), .B(n2166), .Z(n2165) );
  NANDN U2206 ( .A(A[985]), .B(n37), .Z(n2166) );
  NANDN U2207 ( .A(n37), .B(A[985]), .Z(n2164) );
  AND U2208 ( .A(n2167), .B(n2168), .Z(n37) );
  NANDN U2209 ( .A(B[984]), .B(n2169), .Z(n2168) );
  NANDN U2210 ( .A(A[984]), .B(n39), .Z(n2169) );
  NANDN U2211 ( .A(n39), .B(A[984]), .Z(n2167) );
  AND U2212 ( .A(n2170), .B(n2171), .Z(n39) );
  NANDN U2213 ( .A(B[983]), .B(n2172), .Z(n2171) );
  NANDN U2214 ( .A(A[983]), .B(n41), .Z(n2172) );
  NANDN U2215 ( .A(n41), .B(A[983]), .Z(n2170) );
  AND U2216 ( .A(n2173), .B(n2174), .Z(n41) );
  NANDN U2217 ( .A(B[982]), .B(n2175), .Z(n2174) );
  NANDN U2218 ( .A(A[982]), .B(n43), .Z(n2175) );
  NANDN U2219 ( .A(n43), .B(A[982]), .Z(n2173) );
  AND U2220 ( .A(n2176), .B(n2177), .Z(n43) );
  NANDN U2221 ( .A(B[981]), .B(n2178), .Z(n2177) );
  NANDN U2222 ( .A(A[981]), .B(n45), .Z(n2178) );
  NANDN U2223 ( .A(n45), .B(A[981]), .Z(n2176) );
  AND U2224 ( .A(n2179), .B(n2180), .Z(n45) );
  NANDN U2225 ( .A(B[980]), .B(n2181), .Z(n2180) );
  NANDN U2226 ( .A(A[980]), .B(n47), .Z(n2181) );
  NANDN U2227 ( .A(n47), .B(A[980]), .Z(n2179) );
  AND U2228 ( .A(n2182), .B(n2183), .Z(n47) );
  NANDN U2229 ( .A(B[979]), .B(n2184), .Z(n2183) );
  NANDN U2230 ( .A(A[979]), .B(n51), .Z(n2184) );
  NANDN U2231 ( .A(n51), .B(A[979]), .Z(n2182) );
  AND U2232 ( .A(n2185), .B(n2186), .Z(n51) );
  NANDN U2233 ( .A(B[978]), .B(n2187), .Z(n2186) );
  NANDN U2234 ( .A(A[978]), .B(n53), .Z(n2187) );
  NANDN U2235 ( .A(n53), .B(A[978]), .Z(n2185) );
  AND U2236 ( .A(n2188), .B(n2189), .Z(n53) );
  NANDN U2237 ( .A(B[977]), .B(n2190), .Z(n2189) );
  NANDN U2238 ( .A(A[977]), .B(n55), .Z(n2190) );
  NANDN U2239 ( .A(n55), .B(A[977]), .Z(n2188) );
  AND U2240 ( .A(n2191), .B(n2192), .Z(n55) );
  NANDN U2241 ( .A(B[976]), .B(n2193), .Z(n2192) );
  NANDN U2242 ( .A(A[976]), .B(n57), .Z(n2193) );
  NANDN U2243 ( .A(n57), .B(A[976]), .Z(n2191) );
  AND U2244 ( .A(n2194), .B(n2195), .Z(n57) );
  NANDN U2245 ( .A(B[975]), .B(n2196), .Z(n2195) );
  NANDN U2246 ( .A(A[975]), .B(n59), .Z(n2196) );
  NANDN U2247 ( .A(n59), .B(A[975]), .Z(n2194) );
  AND U2248 ( .A(n2197), .B(n2198), .Z(n59) );
  NANDN U2249 ( .A(B[974]), .B(n2199), .Z(n2198) );
  NANDN U2250 ( .A(A[974]), .B(n61), .Z(n2199) );
  NANDN U2251 ( .A(n61), .B(A[974]), .Z(n2197) );
  AND U2252 ( .A(n2200), .B(n2201), .Z(n61) );
  NANDN U2253 ( .A(B[973]), .B(n2202), .Z(n2201) );
  NANDN U2254 ( .A(A[973]), .B(n63), .Z(n2202) );
  NANDN U2255 ( .A(n63), .B(A[973]), .Z(n2200) );
  AND U2256 ( .A(n2203), .B(n2204), .Z(n63) );
  NANDN U2257 ( .A(B[972]), .B(n2205), .Z(n2204) );
  NANDN U2258 ( .A(A[972]), .B(n65), .Z(n2205) );
  NANDN U2259 ( .A(n65), .B(A[972]), .Z(n2203) );
  AND U2260 ( .A(n2206), .B(n2207), .Z(n65) );
  NANDN U2261 ( .A(B[971]), .B(n2208), .Z(n2207) );
  NANDN U2262 ( .A(A[971]), .B(n67), .Z(n2208) );
  NANDN U2263 ( .A(n67), .B(A[971]), .Z(n2206) );
  AND U2264 ( .A(n2209), .B(n2210), .Z(n67) );
  NANDN U2265 ( .A(B[970]), .B(n2211), .Z(n2210) );
  NANDN U2266 ( .A(A[970]), .B(n69), .Z(n2211) );
  NANDN U2267 ( .A(n69), .B(A[970]), .Z(n2209) );
  AND U2268 ( .A(n2212), .B(n2213), .Z(n69) );
  NANDN U2269 ( .A(B[969]), .B(n2214), .Z(n2213) );
  NANDN U2270 ( .A(A[969]), .B(n73), .Z(n2214) );
  NANDN U2271 ( .A(n73), .B(A[969]), .Z(n2212) );
  AND U2272 ( .A(n2215), .B(n2216), .Z(n73) );
  NANDN U2273 ( .A(B[968]), .B(n2217), .Z(n2216) );
  NANDN U2274 ( .A(A[968]), .B(n75), .Z(n2217) );
  NANDN U2275 ( .A(n75), .B(A[968]), .Z(n2215) );
  AND U2276 ( .A(n2218), .B(n2219), .Z(n75) );
  NANDN U2277 ( .A(B[967]), .B(n2220), .Z(n2219) );
  NANDN U2278 ( .A(A[967]), .B(n77), .Z(n2220) );
  NANDN U2279 ( .A(n77), .B(A[967]), .Z(n2218) );
  AND U2280 ( .A(n2221), .B(n2222), .Z(n77) );
  NANDN U2281 ( .A(B[966]), .B(n2223), .Z(n2222) );
  NANDN U2282 ( .A(A[966]), .B(n79), .Z(n2223) );
  NANDN U2283 ( .A(n79), .B(A[966]), .Z(n2221) );
  AND U2284 ( .A(n2224), .B(n2225), .Z(n79) );
  NANDN U2285 ( .A(B[965]), .B(n2226), .Z(n2225) );
  NANDN U2286 ( .A(A[965]), .B(n81), .Z(n2226) );
  NANDN U2287 ( .A(n81), .B(A[965]), .Z(n2224) );
  AND U2288 ( .A(n2227), .B(n2228), .Z(n81) );
  NANDN U2289 ( .A(B[964]), .B(n2229), .Z(n2228) );
  NANDN U2290 ( .A(A[964]), .B(n83), .Z(n2229) );
  NANDN U2291 ( .A(n83), .B(A[964]), .Z(n2227) );
  AND U2292 ( .A(n2230), .B(n2231), .Z(n83) );
  NANDN U2293 ( .A(B[963]), .B(n2232), .Z(n2231) );
  NANDN U2294 ( .A(A[963]), .B(n85), .Z(n2232) );
  NANDN U2295 ( .A(n85), .B(A[963]), .Z(n2230) );
  AND U2296 ( .A(n2233), .B(n2234), .Z(n85) );
  NANDN U2297 ( .A(B[962]), .B(n2235), .Z(n2234) );
  NANDN U2298 ( .A(A[962]), .B(n87), .Z(n2235) );
  NANDN U2299 ( .A(n87), .B(A[962]), .Z(n2233) );
  AND U2300 ( .A(n2236), .B(n2237), .Z(n87) );
  NANDN U2301 ( .A(B[961]), .B(n2238), .Z(n2237) );
  NANDN U2302 ( .A(A[961]), .B(n89), .Z(n2238) );
  NANDN U2303 ( .A(n89), .B(A[961]), .Z(n2236) );
  AND U2304 ( .A(n2239), .B(n2240), .Z(n89) );
  NANDN U2305 ( .A(B[960]), .B(n2241), .Z(n2240) );
  NANDN U2306 ( .A(A[960]), .B(n91), .Z(n2241) );
  NANDN U2307 ( .A(n91), .B(A[960]), .Z(n2239) );
  AND U2308 ( .A(n2242), .B(n2243), .Z(n91) );
  NANDN U2309 ( .A(B[959]), .B(n2244), .Z(n2243) );
  NANDN U2310 ( .A(A[959]), .B(n95), .Z(n2244) );
  NANDN U2311 ( .A(n95), .B(A[959]), .Z(n2242) );
  AND U2312 ( .A(n2245), .B(n2246), .Z(n95) );
  NANDN U2313 ( .A(B[958]), .B(n2247), .Z(n2246) );
  NANDN U2314 ( .A(A[958]), .B(n97), .Z(n2247) );
  NANDN U2315 ( .A(n97), .B(A[958]), .Z(n2245) );
  AND U2316 ( .A(n2248), .B(n2249), .Z(n97) );
  NANDN U2317 ( .A(B[957]), .B(n2250), .Z(n2249) );
  NANDN U2318 ( .A(A[957]), .B(n99), .Z(n2250) );
  NANDN U2319 ( .A(n99), .B(A[957]), .Z(n2248) );
  AND U2320 ( .A(n2251), .B(n2252), .Z(n99) );
  NANDN U2321 ( .A(B[956]), .B(n2253), .Z(n2252) );
  NANDN U2322 ( .A(A[956]), .B(n101), .Z(n2253) );
  NANDN U2323 ( .A(n101), .B(A[956]), .Z(n2251) );
  AND U2324 ( .A(n2254), .B(n2255), .Z(n101) );
  NANDN U2325 ( .A(B[955]), .B(n2256), .Z(n2255) );
  NANDN U2326 ( .A(A[955]), .B(n103), .Z(n2256) );
  NANDN U2327 ( .A(n103), .B(A[955]), .Z(n2254) );
  AND U2328 ( .A(n2257), .B(n2258), .Z(n103) );
  NANDN U2329 ( .A(B[954]), .B(n2259), .Z(n2258) );
  NANDN U2330 ( .A(A[954]), .B(n105), .Z(n2259) );
  NANDN U2331 ( .A(n105), .B(A[954]), .Z(n2257) );
  AND U2332 ( .A(n2260), .B(n2261), .Z(n105) );
  NANDN U2333 ( .A(B[953]), .B(n2262), .Z(n2261) );
  NANDN U2334 ( .A(A[953]), .B(n107), .Z(n2262) );
  NANDN U2335 ( .A(n107), .B(A[953]), .Z(n2260) );
  AND U2336 ( .A(n2263), .B(n2264), .Z(n107) );
  NANDN U2337 ( .A(B[952]), .B(n2265), .Z(n2264) );
  NANDN U2338 ( .A(A[952]), .B(n109), .Z(n2265) );
  NANDN U2339 ( .A(n109), .B(A[952]), .Z(n2263) );
  AND U2340 ( .A(n2266), .B(n2267), .Z(n109) );
  NANDN U2341 ( .A(B[951]), .B(n2268), .Z(n2267) );
  NANDN U2342 ( .A(A[951]), .B(n111), .Z(n2268) );
  NANDN U2343 ( .A(n111), .B(A[951]), .Z(n2266) );
  AND U2344 ( .A(n2269), .B(n2270), .Z(n111) );
  NANDN U2345 ( .A(B[950]), .B(n2271), .Z(n2270) );
  NANDN U2346 ( .A(A[950]), .B(n113), .Z(n2271) );
  NANDN U2347 ( .A(n113), .B(A[950]), .Z(n2269) );
  AND U2348 ( .A(n2272), .B(n2273), .Z(n113) );
  NANDN U2349 ( .A(B[949]), .B(n2274), .Z(n2273) );
  NANDN U2350 ( .A(A[949]), .B(n117), .Z(n2274) );
  NANDN U2351 ( .A(n117), .B(A[949]), .Z(n2272) );
  AND U2352 ( .A(n2275), .B(n2276), .Z(n117) );
  NANDN U2353 ( .A(B[948]), .B(n2277), .Z(n2276) );
  NANDN U2354 ( .A(A[948]), .B(n119), .Z(n2277) );
  NANDN U2355 ( .A(n119), .B(A[948]), .Z(n2275) );
  AND U2356 ( .A(n2278), .B(n2279), .Z(n119) );
  NANDN U2357 ( .A(B[947]), .B(n2280), .Z(n2279) );
  NANDN U2358 ( .A(A[947]), .B(n121), .Z(n2280) );
  NANDN U2359 ( .A(n121), .B(A[947]), .Z(n2278) );
  AND U2360 ( .A(n2281), .B(n2282), .Z(n121) );
  NANDN U2361 ( .A(B[946]), .B(n2283), .Z(n2282) );
  NANDN U2362 ( .A(A[946]), .B(n123), .Z(n2283) );
  NANDN U2363 ( .A(n123), .B(A[946]), .Z(n2281) );
  AND U2364 ( .A(n2284), .B(n2285), .Z(n123) );
  NANDN U2365 ( .A(B[945]), .B(n2286), .Z(n2285) );
  NANDN U2366 ( .A(A[945]), .B(n125), .Z(n2286) );
  NANDN U2367 ( .A(n125), .B(A[945]), .Z(n2284) );
  AND U2368 ( .A(n2287), .B(n2288), .Z(n125) );
  NANDN U2369 ( .A(B[944]), .B(n2289), .Z(n2288) );
  NANDN U2370 ( .A(A[944]), .B(n127), .Z(n2289) );
  NANDN U2371 ( .A(n127), .B(A[944]), .Z(n2287) );
  AND U2372 ( .A(n2290), .B(n2291), .Z(n127) );
  NANDN U2373 ( .A(B[943]), .B(n2292), .Z(n2291) );
  NANDN U2374 ( .A(A[943]), .B(n129), .Z(n2292) );
  NANDN U2375 ( .A(n129), .B(A[943]), .Z(n2290) );
  AND U2376 ( .A(n2293), .B(n2294), .Z(n129) );
  NANDN U2377 ( .A(B[942]), .B(n2295), .Z(n2294) );
  NANDN U2378 ( .A(A[942]), .B(n131), .Z(n2295) );
  NANDN U2379 ( .A(n131), .B(A[942]), .Z(n2293) );
  AND U2380 ( .A(n2296), .B(n2297), .Z(n131) );
  NANDN U2381 ( .A(B[941]), .B(n2298), .Z(n2297) );
  NANDN U2382 ( .A(A[941]), .B(n133), .Z(n2298) );
  NANDN U2383 ( .A(n133), .B(A[941]), .Z(n2296) );
  AND U2384 ( .A(n2299), .B(n2300), .Z(n133) );
  NANDN U2385 ( .A(B[940]), .B(n2301), .Z(n2300) );
  NANDN U2386 ( .A(A[940]), .B(n135), .Z(n2301) );
  NANDN U2387 ( .A(n135), .B(A[940]), .Z(n2299) );
  AND U2388 ( .A(n2302), .B(n2303), .Z(n135) );
  NANDN U2389 ( .A(B[939]), .B(n2304), .Z(n2303) );
  NANDN U2390 ( .A(A[939]), .B(n139), .Z(n2304) );
  NANDN U2391 ( .A(n139), .B(A[939]), .Z(n2302) );
  AND U2392 ( .A(n2305), .B(n2306), .Z(n139) );
  NANDN U2393 ( .A(B[938]), .B(n2307), .Z(n2306) );
  NANDN U2394 ( .A(A[938]), .B(n141), .Z(n2307) );
  NANDN U2395 ( .A(n141), .B(A[938]), .Z(n2305) );
  AND U2396 ( .A(n2308), .B(n2309), .Z(n141) );
  NANDN U2397 ( .A(B[937]), .B(n2310), .Z(n2309) );
  NANDN U2398 ( .A(A[937]), .B(n143), .Z(n2310) );
  NANDN U2399 ( .A(n143), .B(A[937]), .Z(n2308) );
  AND U2400 ( .A(n2311), .B(n2312), .Z(n143) );
  NANDN U2401 ( .A(B[936]), .B(n2313), .Z(n2312) );
  NANDN U2402 ( .A(A[936]), .B(n145), .Z(n2313) );
  NANDN U2403 ( .A(n145), .B(A[936]), .Z(n2311) );
  AND U2404 ( .A(n2314), .B(n2315), .Z(n145) );
  NANDN U2405 ( .A(B[935]), .B(n2316), .Z(n2315) );
  NANDN U2406 ( .A(A[935]), .B(n147), .Z(n2316) );
  NANDN U2407 ( .A(n147), .B(A[935]), .Z(n2314) );
  AND U2408 ( .A(n2317), .B(n2318), .Z(n147) );
  NANDN U2409 ( .A(B[934]), .B(n2319), .Z(n2318) );
  NANDN U2410 ( .A(A[934]), .B(n149), .Z(n2319) );
  NANDN U2411 ( .A(n149), .B(A[934]), .Z(n2317) );
  AND U2412 ( .A(n2320), .B(n2321), .Z(n149) );
  NANDN U2413 ( .A(B[933]), .B(n2322), .Z(n2321) );
  NANDN U2414 ( .A(A[933]), .B(n151), .Z(n2322) );
  NANDN U2415 ( .A(n151), .B(A[933]), .Z(n2320) );
  AND U2416 ( .A(n2323), .B(n2324), .Z(n151) );
  NANDN U2417 ( .A(B[932]), .B(n2325), .Z(n2324) );
  NANDN U2418 ( .A(A[932]), .B(n153), .Z(n2325) );
  NANDN U2419 ( .A(n153), .B(A[932]), .Z(n2323) );
  AND U2420 ( .A(n2326), .B(n2327), .Z(n153) );
  NANDN U2421 ( .A(B[931]), .B(n2328), .Z(n2327) );
  NANDN U2422 ( .A(A[931]), .B(n155), .Z(n2328) );
  NANDN U2423 ( .A(n155), .B(A[931]), .Z(n2326) );
  AND U2424 ( .A(n2329), .B(n2330), .Z(n155) );
  NANDN U2425 ( .A(B[930]), .B(n2331), .Z(n2330) );
  NANDN U2426 ( .A(A[930]), .B(n157), .Z(n2331) );
  NANDN U2427 ( .A(n157), .B(A[930]), .Z(n2329) );
  AND U2428 ( .A(n2332), .B(n2333), .Z(n157) );
  NANDN U2429 ( .A(B[929]), .B(n2334), .Z(n2333) );
  NANDN U2430 ( .A(A[929]), .B(n161), .Z(n2334) );
  NANDN U2431 ( .A(n161), .B(A[929]), .Z(n2332) );
  AND U2432 ( .A(n2335), .B(n2336), .Z(n161) );
  NANDN U2433 ( .A(B[928]), .B(n2337), .Z(n2336) );
  NANDN U2434 ( .A(A[928]), .B(n163), .Z(n2337) );
  NANDN U2435 ( .A(n163), .B(A[928]), .Z(n2335) );
  AND U2436 ( .A(n2338), .B(n2339), .Z(n163) );
  NANDN U2437 ( .A(B[927]), .B(n2340), .Z(n2339) );
  NANDN U2438 ( .A(A[927]), .B(n165), .Z(n2340) );
  NANDN U2439 ( .A(n165), .B(A[927]), .Z(n2338) );
  AND U2440 ( .A(n2341), .B(n2342), .Z(n165) );
  NANDN U2441 ( .A(B[926]), .B(n2343), .Z(n2342) );
  NANDN U2442 ( .A(A[926]), .B(n167), .Z(n2343) );
  NANDN U2443 ( .A(n167), .B(A[926]), .Z(n2341) );
  AND U2444 ( .A(n2344), .B(n2345), .Z(n167) );
  NANDN U2445 ( .A(B[925]), .B(n2346), .Z(n2345) );
  NANDN U2446 ( .A(A[925]), .B(n169), .Z(n2346) );
  NANDN U2447 ( .A(n169), .B(A[925]), .Z(n2344) );
  AND U2448 ( .A(n2347), .B(n2348), .Z(n169) );
  NANDN U2449 ( .A(B[924]), .B(n2349), .Z(n2348) );
  NANDN U2450 ( .A(A[924]), .B(n171), .Z(n2349) );
  NANDN U2451 ( .A(n171), .B(A[924]), .Z(n2347) );
  AND U2452 ( .A(n2350), .B(n2351), .Z(n171) );
  NANDN U2453 ( .A(B[923]), .B(n2352), .Z(n2351) );
  NANDN U2454 ( .A(A[923]), .B(n173), .Z(n2352) );
  NANDN U2455 ( .A(n173), .B(A[923]), .Z(n2350) );
  AND U2456 ( .A(n2353), .B(n2354), .Z(n173) );
  NANDN U2457 ( .A(B[922]), .B(n2355), .Z(n2354) );
  NANDN U2458 ( .A(A[922]), .B(n175), .Z(n2355) );
  NANDN U2459 ( .A(n175), .B(A[922]), .Z(n2353) );
  AND U2460 ( .A(n2356), .B(n2357), .Z(n175) );
  NANDN U2461 ( .A(B[921]), .B(n2358), .Z(n2357) );
  NANDN U2462 ( .A(A[921]), .B(n177), .Z(n2358) );
  NANDN U2463 ( .A(n177), .B(A[921]), .Z(n2356) );
  AND U2464 ( .A(n2359), .B(n2360), .Z(n177) );
  NANDN U2465 ( .A(B[920]), .B(n2361), .Z(n2360) );
  NANDN U2466 ( .A(A[920]), .B(n179), .Z(n2361) );
  NANDN U2467 ( .A(n179), .B(A[920]), .Z(n2359) );
  AND U2468 ( .A(n2362), .B(n2363), .Z(n179) );
  NANDN U2469 ( .A(B[919]), .B(n2364), .Z(n2363) );
  NANDN U2470 ( .A(A[919]), .B(n183), .Z(n2364) );
  NANDN U2471 ( .A(n183), .B(A[919]), .Z(n2362) );
  AND U2472 ( .A(n2365), .B(n2366), .Z(n183) );
  NANDN U2473 ( .A(B[918]), .B(n2367), .Z(n2366) );
  NANDN U2474 ( .A(A[918]), .B(n185), .Z(n2367) );
  NANDN U2475 ( .A(n185), .B(A[918]), .Z(n2365) );
  AND U2476 ( .A(n2368), .B(n2369), .Z(n185) );
  NANDN U2477 ( .A(B[917]), .B(n2370), .Z(n2369) );
  NANDN U2478 ( .A(A[917]), .B(n187), .Z(n2370) );
  NANDN U2479 ( .A(n187), .B(A[917]), .Z(n2368) );
  AND U2480 ( .A(n2371), .B(n2372), .Z(n187) );
  NANDN U2481 ( .A(B[916]), .B(n2373), .Z(n2372) );
  NANDN U2482 ( .A(A[916]), .B(n189), .Z(n2373) );
  NANDN U2483 ( .A(n189), .B(A[916]), .Z(n2371) );
  AND U2484 ( .A(n2374), .B(n2375), .Z(n189) );
  NANDN U2485 ( .A(B[915]), .B(n2376), .Z(n2375) );
  NANDN U2486 ( .A(A[915]), .B(n191), .Z(n2376) );
  NANDN U2487 ( .A(n191), .B(A[915]), .Z(n2374) );
  AND U2488 ( .A(n2377), .B(n2378), .Z(n191) );
  NANDN U2489 ( .A(B[914]), .B(n2379), .Z(n2378) );
  NANDN U2490 ( .A(A[914]), .B(n193), .Z(n2379) );
  NANDN U2491 ( .A(n193), .B(A[914]), .Z(n2377) );
  AND U2492 ( .A(n2380), .B(n2381), .Z(n193) );
  NANDN U2493 ( .A(B[913]), .B(n2382), .Z(n2381) );
  NANDN U2494 ( .A(A[913]), .B(n195), .Z(n2382) );
  NANDN U2495 ( .A(n195), .B(A[913]), .Z(n2380) );
  AND U2496 ( .A(n2383), .B(n2384), .Z(n195) );
  NANDN U2497 ( .A(B[912]), .B(n2385), .Z(n2384) );
  NANDN U2498 ( .A(A[912]), .B(n197), .Z(n2385) );
  NANDN U2499 ( .A(n197), .B(A[912]), .Z(n2383) );
  AND U2500 ( .A(n2386), .B(n2387), .Z(n197) );
  NANDN U2501 ( .A(B[911]), .B(n2388), .Z(n2387) );
  NANDN U2502 ( .A(A[911]), .B(n199), .Z(n2388) );
  NANDN U2503 ( .A(n199), .B(A[911]), .Z(n2386) );
  AND U2504 ( .A(n2389), .B(n2390), .Z(n199) );
  NANDN U2505 ( .A(B[910]), .B(n2391), .Z(n2390) );
  NANDN U2506 ( .A(A[910]), .B(n201), .Z(n2391) );
  NANDN U2507 ( .A(n201), .B(A[910]), .Z(n2389) );
  AND U2508 ( .A(n2392), .B(n2393), .Z(n201) );
  NANDN U2509 ( .A(B[909]), .B(n2394), .Z(n2393) );
  NANDN U2510 ( .A(A[909]), .B(n205), .Z(n2394) );
  NANDN U2511 ( .A(n205), .B(A[909]), .Z(n2392) );
  AND U2512 ( .A(n2395), .B(n2396), .Z(n205) );
  NANDN U2513 ( .A(B[908]), .B(n2397), .Z(n2396) );
  NANDN U2514 ( .A(A[908]), .B(n207), .Z(n2397) );
  NANDN U2515 ( .A(n207), .B(A[908]), .Z(n2395) );
  AND U2516 ( .A(n2398), .B(n2399), .Z(n207) );
  NANDN U2517 ( .A(B[907]), .B(n2400), .Z(n2399) );
  NANDN U2518 ( .A(A[907]), .B(n209), .Z(n2400) );
  NANDN U2519 ( .A(n209), .B(A[907]), .Z(n2398) );
  AND U2520 ( .A(n2401), .B(n2402), .Z(n209) );
  NANDN U2521 ( .A(B[906]), .B(n2403), .Z(n2402) );
  NANDN U2522 ( .A(A[906]), .B(n211), .Z(n2403) );
  NANDN U2523 ( .A(n211), .B(A[906]), .Z(n2401) );
  AND U2524 ( .A(n2404), .B(n2405), .Z(n211) );
  NANDN U2525 ( .A(B[905]), .B(n2406), .Z(n2405) );
  NANDN U2526 ( .A(A[905]), .B(n213), .Z(n2406) );
  NANDN U2527 ( .A(n213), .B(A[905]), .Z(n2404) );
  AND U2528 ( .A(n2407), .B(n2408), .Z(n213) );
  NANDN U2529 ( .A(B[904]), .B(n2409), .Z(n2408) );
  NANDN U2530 ( .A(A[904]), .B(n215), .Z(n2409) );
  NANDN U2531 ( .A(n215), .B(A[904]), .Z(n2407) );
  AND U2532 ( .A(n2410), .B(n2411), .Z(n215) );
  NANDN U2533 ( .A(B[903]), .B(n2412), .Z(n2411) );
  NANDN U2534 ( .A(A[903]), .B(n217), .Z(n2412) );
  NANDN U2535 ( .A(n217), .B(A[903]), .Z(n2410) );
  AND U2536 ( .A(n2413), .B(n2414), .Z(n217) );
  NANDN U2537 ( .A(B[902]), .B(n2415), .Z(n2414) );
  NANDN U2538 ( .A(A[902]), .B(n219), .Z(n2415) );
  NANDN U2539 ( .A(n219), .B(A[902]), .Z(n2413) );
  AND U2540 ( .A(n2416), .B(n2417), .Z(n219) );
  NANDN U2541 ( .A(B[901]), .B(n2418), .Z(n2417) );
  NANDN U2542 ( .A(A[901]), .B(n221), .Z(n2418) );
  NANDN U2543 ( .A(n221), .B(A[901]), .Z(n2416) );
  AND U2544 ( .A(n2419), .B(n2420), .Z(n221) );
  NANDN U2545 ( .A(B[900]), .B(n2421), .Z(n2420) );
  NANDN U2546 ( .A(A[900]), .B(n223), .Z(n2421) );
  NANDN U2547 ( .A(n223), .B(A[900]), .Z(n2419) );
  AND U2548 ( .A(n2422), .B(n2423), .Z(n223) );
  NANDN U2549 ( .A(B[899]), .B(n2424), .Z(n2423) );
  NANDN U2550 ( .A(A[899]), .B(n229), .Z(n2424) );
  NANDN U2551 ( .A(n229), .B(A[899]), .Z(n2422) );
  AND U2552 ( .A(n2425), .B(n2426), .Z(n229) );
  NANDN U2553 ( .A(B[898]), .B(n2427), .Z(n2426) );
  NANDN U2554 ( .A(A[898]), .B(n231), .Z(n2427) );
  NANDN U2555 ( .A(n231), .B(A[898]), .Z(n2425) );
  AND U2556 ( .A(n2428), .B(n2429), .Z(n231) );
  NANDN U2557 ( .A(B[897]), .B(n2430), .Z(n2429) );
  NANDN U2558 ( .A(A[897]), .B(n233), .Z(n2430) );
  NANDN U2559 ( .A(n233), .B(A[897]), .Z(n2428) );
  AND U2560 ( .A(n2431), .B(n2432), .Z(n233) );
  NANDN U2561 ( .A(B[896]), .B(n2433), .Z(n2432) );
  NANDN U2562 ( .A(A[896]), .B(n235), .Z(n2433) );
  NANDN U2563 ( .A(n235), .B(A[896]), .Z(n2431) );
  AND U2564 ( .A(n2434), .B(n2435), .Z(n235) );
  NANDN U2565 ( .A(B[895]), .B(n2436), .Z(n2435) );
  NANDN U2566 ( .A(A[895]), .B(n237), .Z(n2436) );
  NANDN U2567 ( .A(n237), .B(A[895]), .Z(n2434) );
  AND U2568 ( .A(n2437), .B(n2438), .Z(n237) );
  NANDN U2569 ( .A(B[894]), .B(n2439), .Z(n2438) );
  NANDN U2570 ( .A(A[894]), .B(n239), .Z(n2439) );
  NANDN U2571 ( .A(n239), .B(A[894]), .Z(n2437) );
  AND U2572 ( .A(n2440), .B(n2441), .Z(n239) );
  NANDN U2573 ( .A(B[893]), .B(n2442), .Z(n2441) );
  NANDN U2574 ( .A(A[893]), .B(n241), .Z(n2442) );
  NANDN U2575 ( .A(n241), .B(A[893]), .Z(n2440) );
  AND U2576 ( .A(n2443), .B(n2444), .Z(n241) );
  NANDN U2577 ( .A(B[892]), .B(n2445), .Z(n2444) );
  NANDN U2578 ( .A(A[892]), .B(n243), .Z(n2445) );
  NANDN U2579 ( .A(n243), .B(A[892]), .Z(n2443) );
  AND U2580 ( .A(n2446), .B(n2447), .Z(n243) );
  NANDN U2581 ( .A(B[891]), .B(n2448), .Z(n2447) );
  NANDN U2582 ( .A(A[891]), .B(n245), .Z(n2448) );
  NANDN U2583 ( .A(n245), .B(A[891]), .Z(n2446) );
  AND U2584 ( .A(n2449), .B(n2450), .Z(n245) );
  NANDN U2585 ( .A(B[890]), .B(n2451), .Z(n2450) );
  NANDN U2586 ( .A(A[890]), .B(n247), .Z(n2451) );
  NANDN U2587 ( .A(n247), .B(A[890]), .Z(n2449) );
  AND U2588 ( .A(n2452), .B(n2453), .Z(n247) );
  NANDN U2589 ( .A(B[889]), .B(n2454), .Z(n2453) );
  NANDN U2590 ( .A(A[889]), .B(n251), .Z(n2454) );
  NANDN U2591 ( .A(n251), .B(A[889]), .Z(n2452) );
  AND U2592 ( .A(n2455), .B(n2456), .Z(n251) );
  NANDN U2593 ( .A(B[888]), .B(n2457), .Z(n2456) );
  NANDN U2594 ( .A(A[888]), .B(n253), .Z(n2457) );
  NANDN U2595 ( .A(n253), .B(A[888]), .Z(n2455) );
  AND U2596 ( .A(n2458), .B(n2459), .Z(n253) );
  NANDN U2597 ( .A(B[887]), .B(n2460), .Z(n2459) );
  NANDN U2598 ( .A(A[887]), .B(n255), .Z(n2460) );
  NANDN U2599 ( .A(n255), .B(A[887]), .Z(n2458) );
  AND U2600 ( .A(n2461), .B(n2462), .Z(n255) );
  NANDN U2601 ( .A(B[886]), .B(n2463), .Z(n2462) );
  NANDN U2602 ( .A(A[886]), .B(n257), .Z(n2463) );
  NANDN U2603 ( .A(n257), .B(A[886]), .Z(n2461) );
  AND U2604 ( .A(n2464), .B(n2465), .Z(n257) );
  NANDN U2605 ( .A(B[885]), .B(n2466), .Z(n2465) );
  NANDN U2606 ( .A(A[885]), .B(n259), .Z(n2466) );
  NANDN U2607 ( .A(n259), .B(A[885]), .Z(n2464) );
  AND U2608 ( .A(n2467), .B(n2468), .Z(n259) );
  NANDN U2609 ( .A(B[884]), .B(n2469), .Z(n2468) );
  NANDN U2610 ( .A(A[884]), .B(n261), .Z(n2469) );
  NANDN U2611 ( .A(n261), .B(A[884]), .Z(n2467) );
  AND U2612 ( .A(n2470), .B(n2471), .Z(n261) );
  NANDN U2613 ( .A(B[883]), .B(n2472), .Z(n2471) );
  NANDN U2614 ( .A(A[883]), .B(n263), .Z(n2472) );
  NANDN U2615 ( .A(n263), .B(A[883]), .Z(n2470) );
  AND U2616 ( .A(n2473), .B(n2474), .Z(n263) );
  NANDN U2617 ( .A(B[882]), .B(n2475), .Z(n2474) );
  NANDN U2618 ( .A(A[882]), .B(n265), .Z(n2475) );
  NANDN U2619 ( .A(n265), .B(A[882]), .Z(n2473) );
  AND U2620 ( .A(n2476), .B(n2477), .Z(n265) );
  NANDN U2621 ( .A(B[881]), .B(n2478), .Z(n2477) );
  NANDN U2622 ( .A(A[881]), .B(n267), .Z(n2478) );
  NANDN U2623 ( .A(n267), .B(A[881]), .Z(n2476) );
  AND U2624 ( .A(n2479), .B(n2480), .Z(n267) );
  NANDN U2625 ( .A(B[880]), .B(n2481), .Z(n2480) );
  NANDN U2626 ( .A(A[880]), .B(n269), .Z(n2481) );
  NANDN U2627 ( .A(n269), .B(A[880]), .Z(n2479) );
  AND U2628 ( .A(n2482), .B(n2483), .Z(n269) );
  NANDN U2629 ( .A(B[879]), .B(n2484), .Z(n2483) );
  NANDN U2630 ( .A(A[879]), .B(n273), .Z(n2484) );
  NANDN U2631 ( .A(n273), .B(A[879]), .Z(n2482) );
  AND U2632 ( .A(n2485), .B(n2486), .Z(n273) );
  NANDN U2633 ( .A(B[878]), .B(n2487), .Z(n2486) );
  NANDN U2634 ( .A(A[878]), .B(n275), .Z(n2487) );
  NANDN U2635 ( .A(n275), .B(A[878]), .Z(n2485) );
  AND U2636 ( .A(n2488), .B(n2489), .Z(n275) );
  NANDN U2637 ( .A(B[877]), .B(n2490), .Z(n2489) );
  NANDN U2638 ( .A(A[877]), .B(n277), .Z(n2490) );
  NANDN U2639 ( .A(n277), .B(A[877]), .Z(n2488) );
  AND U2640 ( .A(n2491), .B(n2492), .Z(n277) );
  NANDN U2641 ( .A(B[876]), .B(n2493), .Z(n2492) );
  NANDN U2642 ( .A(A[876]), .B(n279), .Z(n2493) );
  NANDN U2643 ( .A(n279), .B(A[876]), .Z(n2491) );
  AND U2644 ( .A(n2494), .B(n2495), .Z(n279) );
  NANDN U2645 ( .A(B[875]), .B(n2496), .Z(n2495) );
  NANDN U2646 ( .A(A[875]), .B(n281), .Z(n2496) );
  NANDN U2647 ( .A(n281), .B(A[875]), .Z(n2494) );
  AND U2648 ( .A(n2497), .B(n2498), .Z(n281) );
  NANDN U2649 ( .A(B[874]), .B(n2499), .Z(n2498) );
  NANDN U2650 ( .A(A[874]), .B(n283), .Z(n2499) );
  NANDN U2651 ( .A(n283), .B(A[874]), .Z(n2497) );
  AND U2652 ( .A(n2500), .B(n2501), .Z(n283) );
  NANDN U2653 ( .A(B[873]), .B(n2502), .Z(n2501) );
  NANDN U2654 ( .A(A[873]), .B(n285), .Z(n2502) );
  NANDN U2655 ( .A(n285), .B(A[873]), .Z(n2500) );
  AND U2656 ( .A(n2503), .B(n2504), .Z(n285) );
  NANDN U2657 ( .A(B[872]), .B(n2505), .Z(n2504) );
  NANDN U2658 ( .A(A[872]), .B(n287), .Z(n2505) );
  NANDN U2659 ( .A(n287), .B(A[872]), .Z(n2503) );
  AND U2660 ( .A(n2506), .B(n2507), .Z(n287) );
  NANDN U2661 ( .A(B[871]), .B(n2508), .Z(n2507) );
  NANDN U2662 ( .A(A[871]), .B(n289), .Z(n2508) );
  NANDN U2663 ( .A(n289), .B(A[871]), .Z(n2506) );
  AND U2664 ( .A(n2509), .B(n2510), .Z(n289) );
  NANDN U2665 ( .A(B[870]), .B(n2511), .Z(n2510) );
  NANDN U2666 ( .A(A[870]), .B(n291), .Z(n2511) );
  NANDN U2667 ( .A(n291), .B(A[870]), .Z(n2509) );
  AND U2668 ( .A(n2512), .B(n2513), .Z(n291) );
  NANDN U2669 ( .A(B[869]), .B(n2514), .Z(n2513) );
  NANDN U2670 ( .A(A[869]), .B(n295), .Z(n2514) );
  NANDN U2671 ( .A(n295), .B(A[869]), .Z(n2512) );
  AND U2672 ( .A(n2515), .B(n2516), .Z(n295) );
  NANDN U2673 ( .A(B[868]), .B(n2517), .Z(n2516) );
  NANDN U2674 ( .A(A[868]), .B(n297), .Z(n2517) );
  NANDN U2675 ( .A(n297), .B(A[868]), .Z(n2515) );
  AND U2676 ( .A(n2518), .B(n2519), .Z(n297) );
  NANDN U2677 ( .A(B[867]), .B(n2520), .Z(n2519) );
  NANDN U2678 ( .A(A[867]), .B(n299), .Z(n2520) );
  NANDN U2679 ( .A(n299), .B(A[867]), .Z(n2518) );
  AND U2680 ( .A(n2521), .B(n2522), .Z(n299) );
  NANDN U2681 ( .A(B[866]), .B(n2523), .Z(n2522) );
  NANDN U2682 ( .A(A[866]), .B(n301), .Z(n2523) );
  NANDN U2683 ( .A(n301), .B(A[866]), .Z(n2521) );
  AND U2684 ( .A(n2524), .B(n2525), .Z(n301) );
  NANDN U2685 ( .A(B[865]), .B(n2526), .Z(n2525) );
  NANDN U2686 ( .A(A[865]), .B(n303), .Z(n2526) );
  NANDN U2687 ( .A(n303), .B(A[865]), .Z(n2524) );
  AND U2688 ( .A(n2527), .B(n2528), .Z(n303) );
  NANDN U2689 ( .A(B[864]), .B(n2529), .Z(n2528) );
  NANDN U2690 ( .A(A[864]), .B(n305), .Z(n2529) );
  NANDN U2691 ( .A(n305), .B(A[864]), .Z(n2527) );
  AND U2692 ( .A(n2530), .B(n2531), .Z(n305) );
  NANDN U2693 ( .A(B[863]), .B(n2532), .Z(n2531) );
  NANDN U2694 ( .A(A[863]), .B(n307), .Z(n2532) );
  NANDN U2695 ( .A(n307), .B(A[863]), .Z(n2530) );
  AND U2696 ( .A(n2533), .B(n2534), .Z(n307) );
  NANDN U2697 ( .A(B[862]), .B(n2535), .Z(n2534) );
  NANDN U2698 ( .A(A[862]), .B(n309), .Z(n2535) );
  NANDN U2699 ( .A(n309), .B(A[862]), .Z(n2533) );
  AND U2700 ( .A(n2536), .B(n2537), .Z(n309) );
  NANDN U2701 ( .A(B[861]), .B(n2538), .Z(n2537) );
  NANDN U2702 ( .A(A[861]), .B(n311), .Z(n2538) );
  NANDN U2703 ( .A(n311), .B(A[861]), .Z(n2536) );
  AND U2704 ( .A(n2539), .B(n2540), .Z(n311) );
  NANDN U2705 ( .A(B[860]), .B(n2541), .Z(n2540) );
  NANDN U2706 ( .A(A[860]), .B(n313), .Z(n2541) );
  NANDN U2707 ( .A(n313), .B(A[860]), .Z(n2539) );
  AND U2708 ( .A(n2542), .B(n2543), .Z(n313) );
  NANDN U2709 ( .A(B[859]), .B(n2544), .Z(n2543) );
  NANDN U2710 ( .A(A[859]), .B(n317), .Z(n2544) );
  NANDN U2711 ( .A(n317), .B(A[859]), .Z(n2542) );
  AND U2712 ( .A(n2545), .B(n2546), .Z(n317) );
  NANDN U2713 ( .A(B[858]), .B(n2547), .Z(n2546) );
  NANDN U2714 ( .A(A[858]), .B(n319), .Z(n2547) );
  NANDN U2715 ( .A(n319), .B(A[858]), .Z(n2545) );
  AND U2716 ( .A(n2548), .B(n2549), .Z(n319) );
  NANDN U2717 ( .A(B[857]), .B(n2550), .Z(n2549) );
  NANDN U2718 ( .A(A[857]), .B(n321), .Z(n2550) );
  NANDN U2719 ( .A(n321), .B(A[857]), .Z(n2548) );
  AND U2720 ( .A(n2551), .B(n2552), .Z(n321) );
  NANDN U2721 ( .A(B[856]), .B(n2553), .Z(n2552) );
  NANDN U2722 ( .A(A[856]), .B(n323), .Z(n2553) );
  NANDN U2723 ( .A(n323), .B(A[856]), .Z(n2551) );
  AND U2724 ( .A(n2554), .B(n2555), .Z(n323) );
  NANDN U2725 ( .A(B[855]), .B(n2556), .Z(n2555) );
  NANDN U2726 ( .A(A[855]), .B(n325), .Z(n2556) );
  NANDN U2727 ( .A(n325), .B(A[855]), .Z(n2554) );
  AND U2728 ( .A(n2557), .B(n2558), .Z(n325) );
  NANDN U2729 ( .A(B[854]), .B(n2559), .Z(n2558) );
  NANDN U2730 ( .A(A[854]), .B(n327), .Z(n2559) );
  NANDN U2731 ( .A(n327), .B(A[854]), .Z(n2557) );
  AND U2732 ( .A(n2560), .B(n2561), .Z(n327) );
  NANDN U2733 ( .A(B[853]), .B(n2562), .Z(n2561) );
  NANDN U2734 ( .A(A[853]), .B(n329), .Z(n2562) );
  NANDN U2735 ( .A(n329), .B(A[853]), .Z(n2560) );
  AND U2736 ( .A(n2563), .B(n2564), .Z(n329) );
  NANDN U2737 ( .A(B[852]), .B(n2565), .Z(n2564) );
  NANDN U2738 ( .A(A[852]), .B(n331), .Z(n2565) );
  NANDN U2739 ( .A(n331), .B(A[852]), .Z(n2563) );
  AND U2740 ( .A(n2566), .B(n2567), .Z(n331) );
  NANDN U2741 ( .A(B[851]), .B(n2568), .Z(n2567) );
  NANDN U2742 ( .A(A[851]), .B(n333), .Z(n2568) );
  NANDN U2743 ( .A(n333), .B(A[851]), .Z(n2566) );
  AND U2744 ( .A(n2569), .B(n2570), .Z(n333) );
  NANDN U2745 ( .A(B[850]), .B(n2571), .Z(n2570) );
  NANDN U2746 ( .A(A[850]), .B(n335), .Z(n2571) );
  NANDN U2747 ( .A(n335), .B(A[850]), .Z(n2569) );
  AND U2748 ( .A(n2572), .B(n2573), .Z(n335) );
  NANDN U2749 ( .A(B[849]), .B(n2574), .Z(n2573) );
  NANDN U2750 ( .A(A[849]), .B(n339), .Z(n2574) );
  NANDN U2751 ( .A(n339), .B(A[849]), .Z(n2572) );
  AND U2752 ( .A(n2575), .B(n2576), .Z(n339) );
  NANDN U2753 ( .A(B[848]), .B(n2577), .Z(n2576) );
  NANDN U2754 ( .A(A[848]), .B(n341), .Z(n2577) );
  NANDN U2755 ( .A(n341), .B(A[848]), .Z(n2575) );
  AND U2756 ( .A(n2578), .B(n2579), .Z(n341) );
  NANDN U2757 ( .A(B[847]), .B(n2580), .Z(n2579) );
  NANDN U2758 ( .A(A[847]), .B(n343), .Z(n2580) );
  NANDN U2759 ( .A(n343), .B(A[847]), .Z(n2578) );
  AND U2760 ( .A(n2581), .B(n2582), .Z(n343) );
  NANDN U2761 ( .A(B[846]), .B(n2583), .Z(n2582) );
  NANDN U2762 ( .A(A[846]), .B(n345), .Z(n2583) );
  NANDN U2763 ( .A(n345), .B(A[846]), .Z(n2581) );
  AND U2764 ( .A(n2584), .B(n2585), .Z(n345) );
  NANDN U2765 ( .A(B[845]), .B(n2586), .Z(n2585) );
  NANDN U2766 ( .A(A[845]), .B(n347), .Z(n2586) );
  NANDN U2767 ( .A(n347), .B(A[845]), .Z(n2584) );
  AND U2768 ( .A(n2587), .B(n2588), .Z(n347) );
  NANDN U2769 ( .A(B[844]), .B(n2589), .Z(n2588) );
  NANDN U2770 ( .A(A[844]), .B(n349), .Z(n2589) );
  NANDN U2771 ( .A(n349), .B(A[844]), .Z(n2587) );
  AND U2772 ( .A(n2590), .B(n2591), .Z(n349) );
  NANDN U2773 ( .A(B[843]), .B(n2592), .Z(n2591) );
  NANDN U2774 ( .A(A[843]), .B(n351), .Z(n2592) );
  NANDN U2775 ( .A(n351), .B(A[843]), .Z(n2590) );
  AND U2776 ( .A(n2593), .B(n2594), .Z(n351) );
  NANDN U2777 ( .A(B[842]), .B(n2595), .Z(n2594) );
  NANDN U2778 ( .A(A[842]), .B(n353), .Z(n2595) );
  NANDN U2779 ( .A(n353), .B(A[842]), .Z(n2593) );
  AND U2780 ( .A(n2596), .B(n2597), .Z(n353) );
  NANDN U2781 ( .A(B[841]), .B(n2598), .Z(n2597) );
  NANDN U2782 ( .A(A[841]), .B(n355), .Z(n2598) );
  NANDN U2783 ( .A(n355), .B(A[841]), .Z(n2596) );
  AND U2784 ( .A(n2599), .B(n2600), .Z(n355) );
  NANDN U2785 ( .A(B[840]), .B(n2601), .Z(n2600) );
  NANDN U2786 ( .A(A[840]), .B(n357), .Z(n2601) );
  NANDN U2787 ( .A(n357), .B(A[840]), .Z(n2599) );
  AND U2788 ( .A(n2602), .B(n2603), .Z(n357) );
  NANDN U2789 ( .A(B[839]), .B(n2604), .Z(n2603) );
  NANDN U2790 ( .A(A[839]), .B(n361), .Z(n2604) );
  NANDN U2791 ( .A(n361), .B(A[839]), .Z(n2602) );
  AND U2792 ( .A(n2605), .B(n2606), .Z(n361) );
  NANDN U2793 ( .A(B[838]), .B(n2607), .Z(n2606) );
  NANDN U2794 ( .A(A[838]), .B(n363), .Z(n2607) );
  NANDN U2795 ( .A(n363), .B(A[838]), .Z(n2605) );
  AND U2796 ( .A(n2608), .B(n2609), .Z(n363) );
  NANDN U2797 ( .A(B[837]), .B(n2610), .Z(n2609) );
  NANDN U2798 ( .A(A[837]), .B(n365), .Z(n2610) );
  NANDN U2799 ( .A(n365), .B(A[837]), .Z(n2608) );
  AND U2800 ( .A(n2611), .B(n2612), .Z(n365) );
  NANDN U2801 ( .A(B[836]), .B(n2613), .Z(n2612) );
  NANDN U2802 ( .A(A[836]), .B(n367), .Z(n2613) );
  NANDN U2803 ( .A(n367), .B(A[836]), .Z(n2611) );
  AND U2804 ( .A(n2614), .B(n2615), .Z(n367) );
  NANDN U2805 ( .A(B[835]), .B(n2616), .Z(n2615) );
  NANDN U2806 ( .A(A[835]), .B(n369), .Z(n2616) );
  NANDN U2807 ( .A(n369), .B(A[835]), .Z(n2614) );
  AND U2808 ( .A(n2617), .B(n2618), .Z(n369) );
  NANDN U2809 ( .A(B[834]), .B(n2619), .Z(n2618) );
  NANDN U2810 ( .A(A[834]), .B(n371), .Z(n2619) );
  NANDN U2811 ( .A(n371), .B(A[834]), .Z(n2617) );
  AND U2812 ( .A(n2620), .B(n2621), .Z(n371) );
  NANDN U2813 ( .A(B[833]), .B(n2622), .Z(n2621) );
  NANDN U2814 ( .A(A[833]), .B(n373), .Z(n2622) );
  NANDN U2815 ( .A(n373), .B(A[833]), .Z(n2620) );
  AND U2816 ( .A(n2623), .B(n2624), .Z(n373) );
  NANDN U2817 ( .A(B[832]), .B(n2625), .Z(n2624) );
  NANDN U2818 ( .A(A[832]), .B(n375), .Z(n2625) );
  NANDN U2819 ( .A(n375), .B(A[832]), .Z(n2623) );
  AND U2820 ( .A(n2626), .B(n2627), .Z(n375) );
  NANDN U2821 ( .A(B[831]), .B(n2628), .Z(n2627) );
  NANDN U2822 ( .A(A[831]), .B(n377), .Z(n2628) );
  NANDN U2823 ( .A(n377), .B(A[831]), .Z(n2626) );
  AND U2824 ( .A(n2629), .B(n2630), .Z(n377) );
  NANDN U2825 ( .A(B[830]), .B(n2631), .Z(n2630) );
  NANDN U2826 ( .A(A[830]), .B(n379), .Z(n2631) );
  NANDN U2827 ( .A(n379), .B(A[830]), .Z(n2629) );
  AND U2828 ( .A(n2632), .B(n2633), .Z(n379) );
  NANDN U2829 ( .A(B[829]), .B(n2634), .Z(n2633) );
  NANDN U2830 ( .A(A[829]), .B(n383), .Z(n2634) );
  NANDN U2831 ( .A(n383), .B(A[829]), .Z(n2632) );
  AND U2832 ( .A(n2635), .B(n2636), .Z(n383) );
  NANDN U2833 ( .A(B[828]), .B(n2637), .Z(n2636) );
  NANDN U2834 ( .A(A[828]), .B(n385), .Z(n2637) );
  NANDN U2835 ( .A(n385), .B(A[828]), .Z(n2635) );
  AND U2836 ( .A(n2638), .B(n2639), .Z(n385) );
  NANDN U2837 ( .A(B[827]), .B(n2640), .Z(n2639) );
  NANDN U2838 ( .A(A[827]), .B(n387), .Z(n2640) );
  NANDN U2839 ( .A(n387), .B(A[827]), .Z(n2638) );
  AND U2840 ( .A(n2641), .B(n2642), .Z(n387) );
  NANDN U2841 ( .A(B[826]), .B(n2643), .Z(n2642) );
  NANDN U2842 ( .A(A[826]), .B(n389), .Z(n2643) );
  NANDN U2843 ( .A(n389), .B(A[826]), .Z(n2641) );
  AND U2844 ( .A(n2644), .B(n2645), .Z(n389) );
  NANDN U2845 ( .A(B[825]), .B(n2646), .Z(n2645) );
  NANDN U2846 ( .A(A[825]), .B(n391), .Z(n2646) );
  NANDN U2847 ( .A(n391), .B(A[825]), .Z(n2644) );
  AND U2848 ( .A(n2647), .B(n2648), .Z(n391) );
  NANDN U2849 ( .A(B[824]), .B(n2649), .Z(n2648) );
  NANDN U2850 ( .A(A[824]), .B(n393), .Z(n2649) );
  NANDN U2851 ( .A(n393), .B(A[824]), .Z(n2647) );
  AND U2852 ( .A(n2650), .B(n2651), .Z(n393) );
  NANDN U2853 ( .A(B[823]), .B(n2652), .Z(n2651) );
  NANDN U2854 ( .A(A[823]), .B(n395), .Z(n2652) );
  NANDN U2855 ( .A(n395), .B(A[823]), .Z(n2650) );
  AND U2856 ( .A(n2653), .B(n2654), .Z(n395) );
  NANDN U2857 ( .A(B[822]), .B(n2655), .Z(n2654) );
  NANDN U2858 ( .A(A[822]), .B(n397), .Z(n2655) );
  NANDN U2859 ( .A(n397), .B(A[822]), .Z(n2653) );
  AND U2860 ( .A(n2656), .B(n2657), .Z(n397) );
  NANDN U2861 ( .A(B[821]), .B(n2658), .Z(n2657) );
  NANDN U2862 ( .A(A[821]), .B(n399), .Z(n2658) );
  NANDN U2863 ( .A(n399), .B(A[821]), .Z(n2656) );
  AND U2864 ( .A(n2659), .B(n2660), .Z(n399) );
  NANDN U2865 ( .A(B[820]), .B(n2661), .Z(n2660) );
  NANDN U2866 ( .A(A[820]), .B(n401), .Z(n2661) );
  NANDN U2867 ( .A(n401), .B(A[820]), .Z(n2659) );
  AND U2868 ( .A(n2662), .B(n2663), .Z(n401) );
  NANDN U2869 ( .A(B[819]), .B(n2664), .Z(n2663) );
  NANDN U2870 ( .A(A[819]), .B(n405), .Z(n2664) );
  NANDN U2871 ( .A(n405), .B(A[819]), .Z(n2662) );
  AND U2872 ( .A(n2665), .B(n2666), .Z(n405) );
  NANDN U2873 ( .A(B[818]), .B(n2667), .Z(n2666) );
  NANDN U2874 ( .A(A[818]), .B(n407), .Z(n2667) );
  NANDN U2875 ( .A(n407), .B(A[818]), .Z(n2665) );
  AND U2876 ( .A(n2668), .B(n2669), .Z(n407) );
  NANDN U2877 ( .A(B[817]), .B(n2670), .Z(n2669) );
  NANDN U2878 ( .A(A[817]), .B(n409), .Z(n2670) );
  NANDN U2879 ( .A(n409), .B(A[817]), .Z(n2668) );
  AND U2880 ( .A(n2671), .B(n2672), .Z(n409) );
  NANDN U2881 ( .A(B[816]), .B(n2673), .Z(n2672) );
  NANDN U2882 ( .A(A[816]), .B(n411), .Z(n2673) );
  NANDN U2883 ( .A(n411), .B(A[816]), .Z(n2671) );
  AND U2884 ( .A(n2674), .B(n2675), .Z(n411) );
  NANDN U2885 ( .A(B[815]), .B(n2676), .Z(n2675) );
  NANDN U2886 ( .A(A[815]), .B(n413), .Z(n2676) );
  NANDN U2887 ( .A(n413), .B(A[815]), .Z(n2674) );
  AND U2888 ( .A(n2677), .B(n2678), .Z(n413) );
  NANDN U2889 ( .A(B[814]), .B(n2679), .Z(n2678) );
  NANDN U2890 ( .A(A[814]), .B(n415), .Z(n2679) );
  NANDN U2891 ( .A(n415), .B(A[814]), .Z(n2677) );
  AND U2892 ( .A(n2680), .B(n2681), .Z(n415) );
  NANDN U2893 ( .A(B[813]), .B(n2682), .Z(n2681) );
  NANDN U2894 ( .A(A[813]), .B(n417), .Z(n2682) );
  NANDN U2895 ( .A(n417), .B(A[813]), .Z(n2680) );
  AND U2896 ( .A(n2683), .B(n2684), .Z(n417) );
  NANDN U2897 ( .A(B[812]), .B(n2685), .Z(n2684) );
  NANDN U2898 ( .A(A[812]), .B(n419), .Z(n2685) );
  NANDN U2899 ( .A(n419), .B(A[812]), .Z(n2683) );
  AND U2900 ( .A(n2686), .B(n2687), .Z(n419) );
  NANDN U2901 ( .A(B[811]), .B(n2688), .Z(n2687) );
  NANDN U2902 ( .A(A[811]), .B(n421), .Z(n2688) );
  NANDN U2903 ( .A(n421), .B(A[811]), .Z(n2686) );
  AND U2904 ( .A(n2689), .B(n2690), .Z(n421) );
  NANDN U2905 ( .A(B[810]), .B(n2691), .Z(n2690) );
  NANDN U2906 ( .A(A[810]), .B(n423), .Z(n2691) );
  NANDN U2907 ( .A(n423), .B(A[810]), .Z(n2689) );
  AND U2908 ( .A(n2692), .B(n2693), .Z(n423) );
  NANDN U2909 ( .A(B[809]), .B(n2694), .Z(n2693) );
  NANDN U2910 ( .A(A[809]), .B(n427), .Z(n2694) );
  NANDN U2911 ( .A(n427), .B(A[809]), .Z(n2692) );
  AND U2912 ( .A(n2695), .B(n2696), .Z(n427) );
  NANDN U2913 ( .A(B[808]), .B(n2697), .Z(n2696) );
  NANDN U2914 ( .A(A[808]), .B(n429), .Z(n2697) );
  NANDN U2915 ( .A(n429), .B(A[808]), .Z(n2695) );
  AND U2916 ( .A(n2698), .B(n2699), .Z(n429) );
  NANDN U2917 ( .A(B[807]), .B(n2700), .Z(n2699) );
  NANDN U2918 ( .A(A[807]), .B(n431), .Z(n2700) );
  NANDN U2919 ( .A(n431), .B(A[807]), .Z(n2698) );
  AND U2920 ( .A(n2701), .B(n2702), .Z(n431) );
  NANDN U2921 ( .A(B[806]), .B(n2703), .Z(n2702) );
  NANDN U2922 ( .A(A[806]), .B(n433), .Z(n2703) );
  NANDN U2923 ( .A(n433), .B(A[806]), .Z(n2701) );
  AND U2924 ( .A(n2704), .B(n2705), .Z(n433) );
  NANDN U2925 ( .A(B[805]), .B(n2706), .Z(n2705) );
  NANDN U2926 ( .A(A[805]), .B(n435), .Z(n2706) );
  NANDN U2927 ( .A(n435), .B(A[805]), .Z(n2704) );
  AND U2928 ( .A(n2707), .B(n2708), .Z(n435) );
  NANDN U2929 ( .A(B[804]), .B(n2709), .Z(n2708) );
  NANDN U2930 ( .A(A[804]), .B(n437), .Z(n2709) );
  NANDN U2931 ( .A(n437), .B(A[804]), .Z(n2707) );
  AND U2932 ( .A(n2710), .B(n2711), .Z(n437) );
  NANDN U2933 ( .A(B[803]), .B(n2712), .Z(n2711) );
  NANDN U2934 ( .A(A[803]), .B(n439), .Z(n2712) );
  NANDN U2935 ( .A(n439), .B(A[803]), .Z(n2710) );
  AND U2936 ( .A(n2713), .B(n2714), .Z(n439) );
  NANDN U2937 ( .A(B[802]), .B(n2715), .Z(n2714) );
  NANDN U2938 ( .A(A[802]), .B(n441), .Z(n2715) );
  NANDN U2939 ( .A(n441), .B(A[802]), .Z(n2713) );
  AND U2940 ( .A(n2716), .B(n2717), .Z(n441) );
  NANDN U2941 ( .A(B[801]), .B(n2718), .Z(n2717) );
  NANDN U2942 ( .A(A[801]), .B(n443), .Z(n2718) );
  NANDN U2943 ( .A(n443), .B(A[801]), .Z(n2716) );
  AND U2944 ( .A(n2719), .B(n2720), .Z(n443) );
  NANDN U2945 ( .A(B[800]), .B(n2721), .Z(n2720) );
  NANDN U2946 ( .A(A[800]), .B(n445), .Z(n2721) );
  NANDN U2947 ( .A(n445), .B(A[800]), .Z(n2719) );
  AND U2948 ( .A(n2722), .B(n2723), .Z(n445) );
  NANDN U2949 ( .A(B[799]), .B(n2724), .Z(n2723) );
  NANDN U2950 ( .A(A[799]), .B(n451), .Z(n2724) );
  NANDN U2951 ( .A(n451), .B(A[799]), .Z(n2722) );
  AND U2952 ( .A(n2725), .B(n2726), .Z(n451) );
  NANDN U2953 ( .A(B[798]), .B(n2727), .Z(n2726) );
  NANDN U2954 ( .A(A[798]), .B(n453), .Z(n2727) );
  NANDN U2955 ( .A(n453), .B(A[798]), .Z(n2725) );
  AND U2956 ( .A(n2728), .B(n2729), .Z(n453) );
  NANDN U2957 ( .A(B[797]), .B(n2730), .Z(n2729) );
  NANDN U2958 ( .A(A[797]), .B(n455), .Z(n2730) );
  NANDN U2959 ( .A(n455), .B(A[797]), .Z(n2728) );
  AND U2960 ( .A(n2731), .B(n2732), .Z(n455) );
  NANDN U2961 ( .A(B[796]), .B(n2733), .Z(n2732) );
  NANDN U2962 ( .A(A[796]), .B(n457), .Z(n2733) );
  NANDN U2963 ( .A(n457), .B(A[796]), .Z(n2731) );
  AND U2964 ( .A(n2734), .B(n2735), .Z(n457) );
  NANDN U2965 ( .A(B[795]), .B(n2736), .Z(n2735) );
  NANDN U2966 ( .A(A[795]), .B(n459), .Z(n2736) );
  NANDN U2967 ( .A(n459), .B(A[795]), .Z(n2734) );
  AND U2968 ( .A(n2737), .B(n2738), .Z(n459) );
  NANDN U2969 ( .A(B[794]), .B(n2739), .Z(n2738) );
  NANDN U2970 ( .A(A[794]), .B(n461), .Z(n2739) );
  NANDN U2971 ( .A(n461), .B(A[794]), .Z(n2737) );
  AND U2972 ( .A(n2740), .B(n2741), .Z(n461) );
  NANDN U2973 ( .A(B[793]), .B(n2742), .Z(n2741) );
  NANDN U2974 ( .A(A[793]), .B(n463), .Z(n2742) );
  NANDN U2975 ( .A(n463), .B(A[793]), .Z(n2740) );
  AND U2976 ( .A(n2743), .B(n2744), .Z(n463) );
  NANDN U2977 ( .A(B[792]), .B(n2745), .Z(n2744) );
  NANDN U2978 ( .A(A[792]), .B(n465), .Z(n2745) );
  NANDN U2979 ( .A(n465), .B(A[792]), .Z(n2743) );
  AND U2980 ( .A(n2746), .B(n2747), .Z(n465) );
  NANDN U2981 ( .A(B[791]), .B(n2748), .Z(n2747) );
  NANDN U2982 ( .A(A[791]), .B(n467), .Z(n2748) );
  NANDN U2983 ( .A(n467), .B(A[791]), .Z(n2746) );
  AND U2984 ( .A(n2749), .B(n2750), .Z(n467) );
  NANDN U2985 ( .A(B[790]), .B(n2751), .Z(n2750) );
  NANDN U2986 ( .A(A[790]), .B(n469), .Z(n2751) );
  NANDN U2987 ( .A(n469), .B(A[790]), .Z(n2749) );
  AND U2988 ( .A(n2752), .B(n2753), .Z(n469) );
  NANDN U2989 ( .A(B[789]), .B(n2754), .Z(n2753) );
  NANDN U2990 ( .A(A[789]), .B(n473), .Z(n2754) );
  NANDN U2991 ( .A(n473), .B(A[789]), .Z(n2752) );
  AND U2992 ( .A(n2755), .B(n2756), .Z(n473) );
  NANDN U2993 ( .A(B[788]), .B(n2757), .Z(n2756) );
  NANDN U2994 ( .A(A[788]), .B(n475), .Z(n2757) );
  NANDN U2995 ( .A(n475), .B(A[788]), .Z(n2755) );
  AND U2996 ( .A(n2758), .B(n2759), .Z(n475) );
  NANDN U2997 ( .A(B[787]), .B(n2760), .Z(n2759) );
  NANDN U2998 ( .A(A[787]), .B(n477), .Z(n2760) );
  NANDN U2999 ( .A(n477), .B(A[787]), .Z(n2758) );
  AND U3000 ( .A(n2761), .B(n2762), .Z(n477) );
  NANDN U3001 ( .A(B[786]), .B(n2763), .Z(n2762) );
  NANDN U3002 ( .A(A[786]), .B(n479), .Z(n2763) );
  NANDN U3003 ( .A(n479), .B(A[786]), .Z(n2761) );
  AND U3004 ( .A(n2764), .B(n2765), .Z(n479) );
  NANDN U3005 ( .A(B[785]), .B(n2766), .Z(n2765) );
  NANDN U3006 ( .A(A[785]), .B(n481), .Z(n2766) );
  NANDN U3007 ( .A(n481), .B(A[785]), .Z(n2764) );
  AND U3008 ( .A(n2767), .B(n2768), .Z(n481) );
  NANDN U3009 ( .A(B[784]), .B(n2769), .Z(n2768) );
  NANDN U3010 ( .A(A[784]), .B(n483), .Z(n2769) );
  NANDN U3011 ( .A(n483), .B(A[784]), .Z(n2767) );
  AND U3012 ( .A(n2770), .B(n2771), .Z(n483) );
  NANDN U3013 ( .A(B[783]), .B(n2772), .Z(n2771) );
  NANDN U3014 ( .A(A[783]), .B(n485), .Z(n2772) );
  NANDN U3015 ( .A(n485), .B(A[783]), .Z(n2770) );
  AND U3016 ( .A(n2773), .B(n2774), .Z(n485) );
  NANDN U3017 ( .A(B[782]), .B(n2775), .Z(n2774) );
  NANDN U3018 ( .A(A[782]), .B(n487), .Z(n2775) );
  NANDN U3019 ( .A(n487), .B(A[782]), .Z(n2773) );
  AND U3020 ( .A(n2776), .B(n2777), .Z(n487) );
  NANDN U3021 ( .A(B[781]), .B(n2778), .Z(n2777) );
  NANDN U3022 ( .A(A[781]), .B(n489), .Z(n2778) );
  NANDN U3023 ( .A(n489), .B(A[781]), .Z(n2776) );
  AND U3024 ( .A(n2779), .B(n2780), .Z(n489) );
  NANDN U3025 ( .A(B[780]), .B(n2781), .Z(n2780) );
  NANDN U3026 ( .A(A[780]), .B(n491), .Z(n2781) );
  NANDN U3027 ( .A(n491), .B(A[780]), .Z(n2779) );
  AND U3028 ( .A(n2782), .B(n2783), .Z(n491) );
  NANDN U3029 ( .A(B[779]), .B(n2784), .Z(n2783) );
  NANDN U3030 ( .A(A[779]), .B(n495), .Z(n2784) );
  NANDN U3031 ( .A(n495), .B(A[779]), .Z(n2782) );
  AND U3032 ( .A(n2785), .B(n2786), .Z(n495) );
  NANDN U3033 ( .A(B[778]), .B(n2787), .Z(n2786) );
  NANDN U3034 ( .A(A[778]), .B(n497), .Z(n2787) );
  NANDN U3035 ( .A(n497), .B(A[778]), .Z(n2785) );
  AND U3036 ( .A(n2788), .B(n2789), .Z(n497) );
  NANDN U3037 ( .A(B[777]), .B(n2790), .Z(n2789) );
  NANDN U3038 ( .A(A[777]), .B(n499), .Z(n2790) );
  NANDN U3039 ( .A(n499), .B(A[777]), .Z(n2788) );
  AND U3040 ( .A(n2791), .B(n2792), .Z(n499) );
  NANDN U3041 ( .A(B[776]), .B(n2793), .Z(n2792) );
  NANDN U3042 ( .A(A[776]), .B(n501), .Z(n2793) );
  NANDN U3043 ( .A(n501), .B(A[776]), .Z(n2791) );
  AND U3044 ( .A(n2794), .B(n2795), .Z(n501) );
  NANDN U3045 ( .A(B[775]), .B(n2796), .Z(n2795) );
  NANDN U3046 ( .A(A[775]), .B(n503), .Z(n2796) );
  NANDN U3047 ( .A(n503), .B(A[775]), .Z(n2794) );
  AND U3048 ( .A(n2797), .B(n2798), .Z(n503) );
  NANDN U3049 ( .A(B[774]), .B(n2799), .Z(n2798) );
  NANDN U3050 ( .A(A[774]), .B(n505), .Z(n2799) );
  NANDN U3051 ( .A(n505), .B(A[774]), .Z(n2797) );
  AND U3052 ( .A(n2800), .B(n2801), .Z(n505) );
  NANDN U3053 ( .A(B[773]), .B(n2802), .Z(n2801) );
  NANDN U3054 ( .A(A[773]), .B(n507), .Z(n2802) );
  NANDN U3055 ( .A(n507), .B(A[773]), .Z(n2800) );
  AND U3056 ( .A(n2803), .B(n2804), .Z(n507) );
  NANDN U3057 ( .A(B[772]), .B(n2805), .Z(n2804) );
  NANDN U3058 ( .A(A[772]), .B(n509), .Z(n2805) );
  NANDN U3059 ( .A(n509), .B(A[772]), .Z(n2803) );
  AND U3060 ( .A(n2806), .B(n2807), .Z(n509) );
  NANDN U3061 ( .A(B[771]), .B(n2808), .Z(n2807) );
  NANDN U3062 ( .A(A[771]), .B(n511), .Z(n2808) );
  NANDN U3063 ( .A(n511), .B(A[771]), .Z(n2806) );
  AND U3064 ( .A(n2809), .B(n2810), .Z(n511) );
  NANDN U3065 ( .A(B[770]), .B(n2811), .Z(n2810) );
  NANDN U3066 ( .A(A[770]), .B(n513), .Z(n2811) );
  NANDN U3067 ( .A(n513), .B(A[770]), .Z(n2809) );
  AND U3068 ( .A(n2812), .B(n2813), .Z(n513) );
  NANDN U3069 ( .A(B[769]), .B(n2814), .Z(n2813) );
  NANDN U3070 ( .A(A[769]), .B(n517), .Z(n2814) );
  NANDN U3071 ( .A(n517), .B(A[769]), .Z(n2812) );
  AND U3072 ( .A(n2815), .B(n2816), .Z(n517) );
  NANDN U3073 ( .A(B[768]), .B(n2817), .Z(n2816) );
  NANDN U3074 ( .A(A[768]), .B(n519), .Z(n2817) );
  NANDN U3075 ( .A(n519), .B(A[768]), .Z(n2815) );
  AND U3076 ( .A(n2818), .B(n2819), .Z(n519) );
  NANDN U3077 ( .A(B[767]), .B(n2820), .Z(n2819) );
  NANDN U3078 ( .A(A[767]), .B(n521), .Z(n2820) );
  NANDN U3079 ( .A(n521), .B(A[767]), .Z(n2818) );
  AND U3080 ( .A(n2821), .B(n2822), .Z(n521) );
  NANDN U3081 ( .A(B[766]), .B(n2823), .Z(n2822) );
  NANDN U3082 ( .A(A[766]), .B(n523), .Z(n2823) );
  NANDN U3083 ( .A(n523), .B(A[766]), .Z(n2821) );
  AND U3084 ( .A(n2824), .B(n2825), .Z(n523) );
  NANDN U3085 ( .A(B[765]), .B(n2826), .Z(n2825) );
  NANDN U3086 ( .A(A[765]), .B(n525), .Z(n2826) );
  NANDN U3087 ( .A(n525), .B(A[765]), .Z(n2824) );
  AND U3088 ( .A(n2827), .B(n2828), .Z(n525) );
  NANDN U3089 ( .A(B[764]), .B(n2829), .Z(n2828) );
  NANDN U3090 ( .A(A[764]), .B(n527), .Z(n2829) );
  NANDN U3091 ( .A(n527), .B(A[764]), .Z(n2827) );
  AND U3092 ( .A(n2830), .B(n2831), .Z(n527) );
  NANDN U3093 ( .A(B[763]), .B(n2832), .Z(n2831) );
  NANDN U3094 ( .A(A[763]), .B(n529), .Z(n2832) );
  NANDN U3095 ( .A(n529), .B(A[763]), .Z(n2830) );
  AND U3096 ( .A(n2833), .B(n2834), .Z(n529) );
  NANDN U3097 ( .A(B[762]), .B(n2835), .Z(n2834) );
  NANDN U3098 ( .A(A[762]), .B(n531), .Z(n2835) );
  NANDN U3099 ( .A(n531), .B(A[762]), .Z(n2833) );
  AND U3100 ( .A(n2836), .B(n2837), .Z(n531) );
  NANDN U3101 ( .A(B[761]), .B(n2838), .Z(n2837) );
  NANDN U3102 ( .A(A[761]), .B(n533), .Z(n2838) );
  NANDN U3103 ( .A(n533), .B(A[761]), .Z(n2836) );
  AND U3104 ( .A(n2839), .B(n2840), .Z(n533) );
  NANDN U3105 ( .A(B[760]), .B(n2841), .Z(n2840) );
  NANDN U3106 ( .A(A[760]), .B(n535), .Z(n2841) );
  NANDN U3107 ( .A(n535), .B(A[760]), .Z(n2839) );
  AND U3108 ( .A(n2842), .B(n2843), .Z(n535) );
  NANDN U3109 ( .A(B[759]), .B(n2844), .Z(n2843) );
  NANDN U3110 ( .A(A[759]), .B(n539), .Z(n2844) );
  NANDN U3111 ( .A(n539), .B(A[759]), .Z(n2842) );
  AND U3112 ( .A(n2845), .B(n2846), .Z(n539) );
  NANDN U3113 ( .A(B[758]), .B(n2847), .Z(n2846) );
  NANDN U3114 ( .A(A[758]), .B(n541), .Z(n2847) );
  NANDN U3115 ( .A(n541), .B(A[758]), .Z(n2845) );
  AND U3116 ( .A(n2848), .B(n2849), .Z(n541) );
  NANDN U3117 ( .A(B[757]), .B(n2850), .Z(n2849) );
  NANDN U3118 ( .A(A[757]), .B(n543), .Z(n2850) );
  NANDN U3119 ( .A(n543), .B(A[757]), .Z(n2848) );
  AND U3120 ( .A(n2851), .B(n2852), .Z(n543) );
  NANDN U3121 ( .A(B[756]), .B(n2853), .Z(n2852) );
  NANDN U3122 ( .A(A[756]), .B(n545), .Z(n2853) );
  NANDN U3123 ( .A(n545), .B(A[756]), .Z(n2851) );
  AND U3124 ( .A(n2854), .B(n2855), .Z(n545) );
  NANDN U3125 ( .A(B[755]), .B(n2856), .Z(n2855) );
  NANDN U3126 ( .A(A[755]), .B(n547), .Z(n2856) );
  NANDN U3127 ( .A(n547), .B(A[755]), .Z(n2854) );
  AND U3128 ( .A(n2857), .B(n2858), .Z(n547) );
  NANDN U3129 ( .A(B[754]), .B(n2859), .Z(n2858) );
  NANDN U3130 ( .A(A[754]), .B(n549), .Z(n2859) );
  NANDN U3131 ( .A(n549), .B(A[754]), .Z(n2857) );
  AND U3132 ( .A(n2860), .B(n2861), .Z(n549) );
  NANDN U3133 ( .A(B[753]), .B(n2862), .Z(n2861) );
  NANDN U3134 ( .A(A[753]), .B(n551), .Z(n2862) );
  NANDN U3135 ( .A(n551), .B(A[753]), .Z(n2860) );
  AND U3136 ( .A(n2863), .B(n2864), .Z(n551) );
  NANDN U3137 ( .A(B[752]), .B(n2865), .Z(n2864) );
  NANDN U3138 ( .A(A[752]), .B(n553), .Z(n2865) );
  NANDN U3139 ( .A(n553), .B(A[752]), .Z(n2863) );
  AND U3140 ( .A(n2866), .B(n2867), .Z(n553) );
  NANDN U3141 ( .A(B[751]), .B(n2868), .Z(n2867) );
  NANDN U3142 ( .A(A[751]), .B(n555), .Z(n2868) );
  NANDN U3143 ( .A(n555), .B(A[751]), .Z(n2866) );
  AND U3144 ( .A(n2869), .B(n2870), .Z(n555) );
  NANDN U3145 ( .A(B[750]), .B(n2871), .Z(n2870) );
  NANDN U3146 ( .A(A[750]), .B(n557), .Z(n2871) );
  NANDN U3147 ( .A(n557), .B(A[750]), .Z(n2869) );
  AND U3148 ( .A(n2872), .B(n2873), .Z(n557) );
  NANDN U3149 ( .A(B[749]), .B(n2874), .Z(n2873) );
  NANDN U3150 ( .A(A[749]), .B(n561), .Z(n2874) );
  NANDN U3151 ( .A(n561), .B(A[749]), .Z(n2872) );
  AND U3152 ( .A(n2875), .B(n2876), .Z(n561) );
  NANDN U3153 ( .A(B[748]), .B(n2877), .Z(n2876) );
  NANDN U3154 ( .A(A[748]), .B(n563), .Z(n2877) );
  NANDN U3155 ( .A(n563), .B(A[748]), .Z(n2875) );
  AND U3156 ( .A(n2878), .B(n2879), .Z(n563) );
  NANDN U3157 ( .A(B[747]), .B(n2880), .Z(n2879) );
  NANDN U3158 ( .A(A[747]), .B(n565), .Z(n2880) );
  NANDN U3159 ( .A(n565), .B(A[747]), .Z(n2878) );
  AND U3160 ( .A(n2881), .B(n2882), .Z(n565) );
  NANDN U3161 ( .A(B[746]), .B(n2883), .Z(n2882) );
  NANDN U3162 ( .A(A[746]), .B(n567), .Z(n2883) );
  NANDN U3163 ( .A(n567), .B(A[746]), .Z(n2881) );
  AND U3164 ( .A(n2884), .B(n2885), .Z(n567) );
  NANDN U3165 ( .A(B[745]), .B(n2886), .Z(n2885) );
  NANDN U3166 ( .A(A[745]), .B(n569), .Z(n2886) );
  NANDN U3167 ( .A(n569), .B(A[745]), .Z(n2884) );
  AND U3168 ( .A(n2887), .B(n2888), .Z(n569) );
  NANDN U3169 ( .A(B[744]), .B(n2889), .Z(n2888) );
  NANDN U3170 ( .A(A[744]), .B(n571), .Z(n2889) );
  NANDN U3171 ( .A(n571), .B(A[744]), .Z(n2887) );
  AND U3172 ( .A(n2890), .B(n2891), .Z(n571) );
  NANDN U3173 ( .A(B[743]), .B(n2892), .Z(n2891) );
  NANDN U3174 ( .A(A[743]), .B(n573), .Z(n2892) );
  NANDN U3175 ( .A(n573), .B(A[743]), .Z(n2890) );
  AND U3176 ( .A(n2893), .B(n2894), .Z(n573) );
  NANDN U3177 ( .A(B[742]), .B(n2895), .Z(n2894) );
  NANDN U3178 ( .A(A[742]), .B(n575), .Z(n2895) );
  NANDN U3179 ( .A(n575), .B(A[742]), .Z(n2893) );
  AND U3180 ( .A(n2896), .B(n2897), .Z(n575) );
  NANDN U3181 ( .A(B[741]), .B(n2898), .Z(n2897) );
  NANDN U3182 ( .A(A[741]), .B(n577), .Z(n2898) );
  NANDN U3183 ( .A(n577), .B(A[741]), .Z(n2896) );
  AND U3184 ( .A(n2899), .B(n2900), .Z(n577) );
  NANDN U3185 ( .A(B[740]), .B(n2901), .Z(n2900) );
  NANDN U3186 ( .A(A[740]), .B(n579), .Z(n2901) );
  NANDN U3187 ( .A(n579), .B(A[740]), .Z(n2899) );
  AND U3188 ( .A(n2902), .B(n2903), .Z(n579) );
  NANDN U3189 ( .A(B[739]), .B(n2904), .Z(n2903) );
  NANDN U3190 ( .A(A[739]), .B(n583), .Z(n2904) );
  NANDN U3191 ( .A(n583), .B(A[739]), .Z(n2902) );
  AND U3192 ( .A(n2905), .B(n2906), .Z(n583) );
  NANDN U3193 ( .A(B[738]), .B(n2907), .Z(n2906) );
  NANDN U3194 ( .A(A[738]), .B(n585), .Z(n2907) );
  NANDN U3195 ( .A(n585), .B(A[738]), .Z(n2905) );
  AND U3196 ( .A(n2908), .B(n2909), .Z(n585) );
  NANDN U3197 ( .A(B[737]), .B(n2910), .Z(n2909) );
  NANDN U3198 ( .A(A[737]), .B(n587), .Z(n2910) );
  NANDN U3199 ( .A(n587), .B(A[737]), .Z(n2908) );
  AND U3200 ( .A(n2911), .B(n2912), .Z(n587) );
  NANDN U3201 ( .A(B[736]), .B(n2913), .Z(n2912) );
  NANDN U3202 ( .A(A[736]), .B(n589), .Z(n2913) );
  NANDN U3203 ( .A(n589), .B(A[736]), .Z(n2911) );
  AND U3204 ( .A(n2914), .B(n2915), .Z(n589) );
  NANDN U3205 ( .A(B[735]), .B(n2916), .Z(n2915) );
  NANDN U3206 ( .A(A[735]), .B(n591), .Z(n2916) );
  NANDN U3207 ( .A(n591), .B(A[735]), .Z(n2914) );
  AND U3208 ( .A(n2917), .B(n2918), .Z(n591) );
  NANDN U3209 ( .A(B[734]), .B(n2919), .Z(n2918) );
  NANDN U3210 ( .A(A[734]), .B(n593), .Z(n2919) );
  NANDN U3211 ( .A(n593), .B(A[734]), .Z(n2917) );
  AND U3212 ( .A(n2920), .B(n2921), .Z(n593) );
  NANDN U3213 ( .A(B[733]), .B(n2922), .Z(n2921) );
  NANDN U3214 ( .A(A[733]), .B(n595), .Z(n2922) );
  NANDN U3215 ( .A(n595), .B(A[733]), .Z(n2920) );
  AND U3216 ( .A(n2923), .B(n2924), .Z(n595) );
  NANDN U3217 ( .A(B[732]), .B(n2925), .Z(n2924) );
  NANDN U3218 ( .A(A[732]), .B(n597), .Z(n2925) );
  NANDN U3219 ( .A(n597), .B(A[732]), .Z(n2923) );
  AND U3220 ( .A(n2926), .B(n2927), .Z(n597) );
  NANDN U3221 ( .A(B[731]), .B(n2928), .Z(n2927) );
  NANDN U3222 ( .A(A[731]), .B(n599), .Z(n2928) );
  NANDN U3223 ( .A(n599), .B(A[731]), .Z(n2926) );
  AND U3224 ( .A(n2929), .B(n2930), .Z(n599) );
  NANDN U3225 ( .A(B[730]), .B(n2931), .Z(n2930) );
  NANDN U3226 ( .A(A[730]), .B(n601), .Z(n2931) );
  NANDN U3227 ( .A(n601), .B(A[730]), .Z(n2929) );
  AND U3228 ( .A(n2932), .B(n2933), .Z(n601) );
  NANDN U3229 ( .A(B[729]), .B(n2934), .Z(n2933) );
  NANDN U3230 ( .A(A[729]), .B(n605), .Z(n2934) );
  NANDN U3231 ( .A(n605), .B(A[729]), .Z(n2932) );
  AND U3232 ( .A(n2935), .B(n2936), .Z(n605) );
  NANDN U3233 ( .A(B[728]), .B(n2937), .Z(n2936) );
  NANDN U3234 ( .A(A[728]), .B(n607), .Z(n2937) );
  NANDN U3235 ( .A(n607), .B(A[728]), .Z(n2935) );
  AND U3236 ( .A(n2938), .B(n2939), .Z(n607) );
  NANDN U3237 ( .A(B[727]), .B(n2940), .Z(n2939) );
  NANDN U3238 ( .A(A[727]), .B(n609), .Z(n2940) );
  NANDN U3239 ( .A(n609), .B(A[727]), .Z(n2938) );
  AND U3240 ( .A(n2941), .B(n2942), .Z(n609) );
  NANDN U3241 ( .A(B[726]), .B(n2943), .Z(n2942) );
  NANDN U3242 ( .A(A[726]), .B(n611), .Z(n2943) );
  NANDN U3243 ( .A(n611), .B(A[726]), .Z(n2941) );
  AND U3244 ( .A(n2944), .B(n2945), .Z(n611) );
  NANDN U3245 ( .A(B[725]), .B(n2946), .Z(n2945) );
  NANDN U3246 ( .A(A[725]), .B(n613), .Z(n2946) );
  NANDN U3247 ( .A(n613), .B(A[725]), .Z(n2944) );
  AND U3248 ( .A(n2947), .B(n2948), .Z(n613) );
  NANDN U3249 ( .A(B[724]), .B(n2949), .Z(n2948) );
  NANDN U3250 ( .A(A[724]), .B(n615), .Z(n2949) );
  NANDN U3251 ( .A(n615), .B(A[724]), .Z(n2947) );
  AND U3252 ( .A(n2950), .B(n2951), .Z(n615) );
  NANDN U3253 ( .A(B[723]), .B(n2952), .Z(n2951) );
  NANDN U3254 ( .A(A[723]), .B(n617), .Z(n2952) );
  NANDN U3255 ( .A(n617), .B(A[723]), .Z(n2950) );
  AND U3256 ( .A(n2953), .B(n2954), .Z(n617) );
  NANDN U3257 ( .A(B[722]), .B(n2955), .Z(n2954) );
  NANDN U3258 ( .A(A[722]), .B(n619), .Z(n2955) );
  NANDN U3259 ( .A(n619), .B(A[722]), .Z(n2953) );
  AND U3260 ( .A(n2956), .B(n2957), .Z(n619) );
  NANDN U3261 ( .A(B[721]), .B(n2958), .Z(n2957) );
  NANDN U3262 ( .A(A[721]), .B(n621), .Z(n2958) );
  NANDN U3263 ( .A(n621), .B(A[721]), .Z(n2956) );
  AND U3264 ( .A(n2959), .B(n2960), .Z(n621) );
  NANDN U3265 ( .A(B[720]), .B(n2961), .Z(n2960) );
  NANDN U3266 ( .A(A[720]), .B(n623), .Z(n2961) );
  NANDN U3267 ( .A(n623), .B(A[720]), .Z(n2959) );
  AND U3268 ( .A(n2962), .B(n2963), .Z(n623) );
  NANDN U3269 ( .A(B[719]), .B(n2964), .Z(n2963) );
  NANDN U3270 ( .A(A[719]), .B(n627), .Z(n2964) );
  NANDN U3271 ( .A(n627), .B(A[719]), .Z(n2962) );
  AND U3272 ( .A(n2965), .B(n2966), .Z(n627) );
  NANDN U3273 ( .A(B[718]), .B(n2967), .Z(n2966) );
  NANDN U3274 ( .A(A[718]), .B(n629), .Z(n2967) );
  NANDN U3275 ( .A(n629), .B(A[718]), .Z(n2965) );
  AND U3276 ( .A(n2968), .B(n2969), .Z(n629) );
  NANDN U3277 ( .A(B[717]), .B(n2970), .Z(n2969) );
  NANDN U3278 ( .A(A[717]), .B(n631), .Z(n2970) );
  NANDN U3279 ( .A(n631), .B(A[717]), .Z(n2968) );
  AND U3280 ( .A(n2971), .B(n2972), .Z(n631) );
  NANDN U3281 ( .A(B[716]), .B(n2973), .Z(n2972) );
  NANDN U3282 ( .A(A[716]), .B(n633), .Z(n2973) );
  NANDN U3283 ( .A(n633), .B(A[716]), .Z(n2971) );
  AND U3284 ( .A(n2974), .B(n2975), .Z(n633) );
  NANDN U3285 ( .A(B[715]), .B(n2976), .Z(n2975) );
  NANDN U3286 ( .A(A[715]), .B(n635), .Z(n2976) );
  NANDN U3287 ( .A(n635), .B(A[715]), .Z(n2974) );
  AND U3288 ( .A(n2977), .B(n2978), .Z(n635) );
  NANDN U3289 ( .A(B[714]), .B(n2979), .Z(n2978) );
  NANDN U3290 ( .A(A[714]), .B(n637), .Z(n2979) );
  NANDN U3291 ( .A(n637), .B(A[714]), .Z(n2977) );
  AND U3292 ( .A(n2980), .B(n2981), .Z(n637) );
  NANDN U3293 ( .A(B[713]), .B(n2982), .Z(n2981) );
  NANDN U3294 ( .A(A[713]), .B(n639), .Z(n2982) );
  NANDN U3295 ( .A(n639), .B(A[713]), .Z(n2980) );
  AND U3296 ( .A(n2983), .B(n2984), .Z(n639) );
  NANDN U3297 ( .A(B[712]), .B(n2985), .Z(n2984) );
  NANDN U3298 ( .A(A[712]), .B(n641), .Z(n2985) );
  NANDN U3299 ( .A(n641), .B(A[712]), .Z(n2983) );
  AND U3300 ( .A(n2986), .B(n2987), .Z(n641) );
  NANDN U3301 ( .A(B[711]), .B(n2988), .Z(n2987) );
  NANDN U3302 ( .A(A[711]), .B(n643), .Z(n2988) );
  NANDN U3303 ( .A(n643), .B(A[711]), .Z(n2986) );
  AND U3304 ( .A(n2989), .B(n2990), .Z(n643) );
  NANDN U3305 ( .A(B[710]), .B(n2991), .Z(n2990) );
  NANDN U3306 ( .A(A[710]), .B(n645), .Z(n2991) );
  NANDN U3307 ( .A(n645), .B(A[710]), .Z(n2989) );
  AND U3308 ( .A(n2992), .B(n2993), .Z(n645) );
  NANDN U3309 ( .A(B[709]), .B(n2994), .Z(n2993) );
  NANDN U3310 ( .A(A[709]), .B(n649), .Z(n2994) );
  NANDN U3311 ( .A(n649), .B(A[709]), .Z(n2992) );
  AND U3312 ( .A(n2995), .B(n2996), .Z(n649) );
  NANDN U3313 ( .A(B[708]), .B(n2997), .Z(n2996) );
  NANDN U3314 ( .A(A[708]), .B(n651), .Z(n2997) );
  NANDN U3315 ( .A(n651), .B(A[708]), .Z(n2995) );
  AND U3316 ( .A(n2998), .B(n2999), .Z(n651) );
  NANDN U3317 ( .A(B[707]), .B(n3000), .Z(n2999) );
  NANDN U3318 ( .A(A[707]), .B(n653), .Z(n3000) );
  NANDN U3319 ( .A(n653), .B(A[707]), .Z(n2998) );
  AND U3320 ( .A(n3001), .B(n3002), .Z(n653) );
  NANDN U3321 ( .A(B[706]), .B(n3003), .Z(n3002) );
  NANDN U3322 ( .A(A[706]), .B(n655), .Z(n3003) );
  NANDN U3323 ( .A(n655), .B(A[706]), .Z(n3001) );
  AND U3324 ( .A(n3004), .B(n3005), .Z(n655) );
  NANDN U3325 ( .A(B[705]), .B(n3006), .Z(n3005) );
  NANDN U3326 ( .A(A[705]), .B(n657), .Z(n3006) );
  NANDN U3327 ( .A(n657), .B(A[705]), .Z(n3004) );
  AND U3328 ( .A(n3007), .B(n3008), .Z(n657) );
  NANDN U3329 ( .A(B[704]), .B(n3009), .Z(n3008) );
  NANDN U3330 ( .A(A[704]), .B(n659), .Z(n3009) );
  NANDN U3331 ( .A(n659), .B(A[704]), .Z(n3007) );
  AND U3332 ( .A(n3010), .B(n3011), .Z(n659) );
  NANDN U3333 ( .A(B[703]), .B(n3012), .Z(n3011) );
  NANDN U3334 ( .A(A[703]), .B(n661), .Z(n3012) );
  NANDN U3335 ( .A(n661), .B(A[703]), .Z(n3010) );
  AND U3336 ( .A(n3013), .B(n3014), .Z(n661) );
  NANDN U3337 ( .A(B[702]), .B(n3015), .Z(n3014) );
  NANDN U3338 ( .A(A[702]), .B(n663), .Z(n3015) );
  NANDN U3339 ( .A(n663), .B(A[702]), .Z(n3013) );
  AND U3340 ( .A(n3016), .B(n3017), .Z(n663) );
  NANDN U3341 ( .A(B[701]), .B(n3018), .Z(n3017) );
  NANDN U3342 ( .A(A[701]), .B(n665), .Z(n3018) );
  NANDN U3343 ( .A(n665), .B(A[701]), .Z(n3016) );
  AND U3344 ( .A(n3019), .B(n3020), .Z(n665) );
  NANDN U3345 ( .A(B[700]), .B(n3021), .Z(n3020) );
  NANDN U3346 ( .A(A[700]), .B(n667), .Z(n3021) );
  NANDN U3347 ( .A(n667), .B(A[700]), .Z(n3019) );
  AND U3348 ( .A(n3022), .B(n3023), .Z(n667) );
  NANDN U3349 ( .A(B[699]), .B(n3024), .Z(n3023) );
  NANDN U3350 ( .A(A[699]), .B(n673), .Z(n3024) );
  NANDN U3351 ( .A(n673), .B(A[699]), .Z(n3022) );
  AND U3352 ( .A(n3025), .B(n3026), .Z(n673) );
  NANDN U3353 ( .A(B[698]), .B(n3027), .Z(n3026) );
  NANDN U3354 ( .A(A[698]), .B(n675), .Z(n3027) );
  NANDN U3355 ( .A(n675), .B(A[698]), .Z(n3025) );
  AND U3356 ( .A(n3028), .B(n3029), .Z(n675) );
  NANDN U3357 ( .A(B[697]), .B(n3030), .Z(n3029) );
  NANDN U3358 ( .A(A[697]), .B(n677), .Z(n3030) );
  NANDN U3359 ( .A(n677), .B(A[697]), .Z(n3028) );
  AND U3360 ( .A(n3031), .B(n3032), .Z(n677) );
  NANDN U3361 ( .A(B[696]), .B(n3033), .Z(n3032) );
  NANDN U3362 ( .A(A[696]), .B(n679), .Z(n3033) );
  NANDN U3363 ( .A(n679), .B(A[696]), .Z(n3031) );
  AND U3364 ( .A(n3034), .B(n3035), .Z(n679) );
  NANDN U3365 ( .A(B[695]), .B(n3036), .Z(n3035) );
  NANDN U3366 ( .A(A[695]), .B(n681), .Z(n3036) );
  NANDN U3367 ( .A(n681), .B(A[695]), .Z(n3034) );
  AND U3368 ( .A(n3037), .B(n3038), .Z(n681) );
  NANDN U3369 ( .A(B[694]), .B(n3039), .Z(n3038) );
  NANDN U3370 ( .A(A[694]), .B(n683), .Z(n3039) );
  NANDN U3371 ( .A(n683), .B(A[694]), .Z(n3037) );
  AND U3372 ( .A(n3040), .B(n3041), .Z(n683) );
  NANDN U3373 ( .A(B[693]), .B(n3042), .Z(n3041) );
  NANDN U3374 ( .A(A[693]), .B(n685), .Z(n3042) );
  NANDN U3375 ( .A(n685), .B(A[693]), .Z(n3040) );
  AND U3376 ( .A(n3043), .B(n3044), .Z(n685) );
  NANDN U3377 ( .A(B[692]), .B(n3045), .Z(n3044) );
  NANDN U3378 ( .A(A[692]), .B(n687), .Z(n3045) );
  NANDN U3379 ( .A(n687), .B(A[692]), .Z(n3043) );
  AND U3380 ( .A(n3046), .B(n3047), .Z(n687) );
  NANDN U3381 ( .A(B[691]), .B(n3048), .Z(n3047) );
  NANDN U3382 ( .A(A[691]), .B(n689), .Z(n3048) );
  NANDN U3383 ( .A(n689), .B(A[691]), .Z(n3046) );
  AND U3384 ( .A(n3049), .B(n3050), .Z(n689) );
  NANDN U3385 ( .A(B[690]), .B(n3051), .Z(n3050) );
  NANDN U3386 ( .A(A[690]), .B(n691), .Z(n3051) );
  NANDN U3387 ( .A(n691), .B(A[690]), .Z(n3049) );
  AND U3388 ( .A(n3052), .B(n3053), .Z(n691) );
  NANDN U3389 ( .A(B[689]), .B(n3054), .Z(n3053) );
  NANDN U3390 ( .A(A[689]), .B(n695), .Z(n3054) );
  NANDN U3391 ( .A(n695), .B(A[689]), .Z(n3052) );
  AND U3392 ( .A(n3055), .B(n3056), .Z(n695) );
  NANDN U3393 ( .A(B[688]), .B(n3057), .Z(n3056) );
  NANDN U3394 ( .A(A[688]), .B(n697), .Z(n3057) );
  NANDN U3395 ( .A(n697), .B(A[688]), .Z(n3055) );
  AND U3396 ( .A(n3058), .B(n3059), .Z(n697) );
  NANDN U3397 ( .A(B[687]), .B(n3060), .Z(n3059) );
  NANDN U3398 ( .A(A[687]), .B(n699), .Z(n3060) );
  NANDN U3399 ( .A(n699), .B(A[687]), .Z(n3058) );
  AND U3400 ( .A(n3061), .B(n3062), .Z(n699) );
  NANDN U3401 ( .A(B[686]), .B(n3063), .Z(n3062) );
  NANDN U3402 ( .A(A[686]), .B(n701), .Z(n3063) );
  NANDN U3403 ( .A(n701), .B(A[686]), .Z(n3061) );
  AND U3404 ( .A(n3064), .B(n3065), .Z(n701) );
  NANDN U3405 ( .A(B[685]), .B(n3066), .Z(n3065) );
  NANDN U3406 ( .A(A[685]), .B(n703), .Z(n3066) );
  NANDN U3407 ( .A(n703), .B(A[685]), .Z(n3064) );
  AND U3408 ( .A(n3067), .B(n3068), .Z(n703) );
  NANDN U3409 ( .A(B[684]), .B(n3069), .Z(n3068) );
  NANDN U3410 ( .A(A[684]), .B(n705), .Z(n3069) );
  NANDN U3411 ( .A(n705), .B(A[684]), .Z(n3067) );
  AND U3412 ( .A(n3070), .B(n3071), .Z(n705) );
  NANDN U3413 ( .A(B[683]), .B(n3072), .Z(n3071) );
  NANDN U3414 ( .A(A[683]), .B(n707), .Z(n3072) );
  NANDN U3415 ( .A(n707), .B(A[683]), .Z(n3070) );
  AND U3416 ( .A(n3073), .B(n3074), .Z(n707) );
  NANDN U3417 ( .A(B[682]), .B(n3075), .Z(n3074) );
  NANDN U3418 ( .A(A[682]), .B(n709), .Z(n3075) );
  NANDN U3419 ( .A(n709), .B(A[682]), .Z(n3073) );
  AND U3420 ( .A(n3076), .B(n3077), .Z(n709) );
  NANDN U3421 ( .A(B[681]), .B(n3078), .Z(n3077) );
  NANDN U3422 ( .A(A[681]), .B(n711), .Z(n3078) );
  NANDN U3423 ( .A(n711), .B(A[681]), .Z(n3076) );
  AND U3424 ( .A(n3079), .B(n3080), .Z(n711) );
  NANDN U3425 ( .A(B[680]), .B(n3081), .Z(n3080) );
  NANDN U3426 ( .A(A[680]), .B(n713), .Z(n3081) );
  NANDN U3427 ( .A(n713), .B(A[680]), .Z(n3079) );
  AND U3428 ( .A(n3082), .B(n3083), .Z(n713) );
  NANDN U3429 ( .A(B[679]), .B(n3084), .Z(n3083) );
  NANDN U3430 ( .A(A[679]), .B(n717), .Z(n3084) );
  NANDN U3431 ( .A(n717), .B(A[679]), .Z(n3082) );
  AND U3432 ( .A(n3085), .B(n3086), .Z(n717) );
  NANDN U3433 ( .A(B[678]), .B(n3087), .Z(n3086) );
  NANDN U3434 ( .A(A[678]), .B(n719), .Z(n3087) );
  NANDN U3435 ( .A(n719), .B(A[678]), .Z(n3085) );
  AND U3436 ( .A(n3088), .B(n3089), .Z(n719) );
  NANDN U3437 ( .A(B[677]), .B(n3090), .Z(n3089) );
  NANDN U3438 ( .A(A[677]), .B(n721), .Z(n3090) );
  NANDN U3439 ( .A(n721), .B(A[677]), .Z(n3088) );
  AND U3440 ( .A(n3091), .B(n3092), .Z(n721) );
  NANDN U3441 ( .A(B[676]), .B(n3093), .Z(n3092) );
  NANDN U3442 ( .A(A[676]), .B(n723), .Z(n3093) );
  NANDN U3443 ( .A(n723), .B(A[676]), .Z(n3091) );
  AND U3444 ( .A(n3094), .B(n3095), .Z(n723) );
  NANDN U3445 ( .A(B[675]), .B(n3096), .Z(n3095) );
  NANDN U3446 ( .A(A[675]), .B(n725), .Z(n3096) );
  NANDN U3447 ( .A(n725), .B(A[675]), .Z(n3094) );
  AND U3448 ( .A(n3097), .B(n3098), .Z(n725) );
  NANDN U3449 ( .A(B[674]), .B(n3099), .Z(n3098) );
  NANDN U3450 ( .A(A[674]), .B(n727), .Z(n3099) );
  NANDN U3451 ( .A(n727), .B(A[674]), .Z(n3097) );
  AND U3452 ( .A(n3100), .B(n3101), .Z(n727) );
  NANDN U3453 ( .A(B[673]), .B(n3102), .Z(n3101) );
  NANDN U3454 ( .A(A[673]), .B(n729), .Z(n3102) );
  NANDN U3455 ( .A(n729), .B(A[673]), .Z(n3100) );
  AND U3456 ( .A(n3103), .B(n3104), .Z(n729) );
  NANDN U3457 ( .A(B[672]), .B(n3105), .Z(n3104) );
  NANDN U3458 ( .A(A[672]), .B(n731), .Z(n3105) );
  NANDN U3459 ( .A(n731), .B(A[672]), .Z(n3103) );
  AND U3460 ( .A(n3106), .B(n3107), .Z(n731) );
  NANDN U3461 ( .A(B[671]), .B(n3108), .Z(n3107) );
  NANDN U3462 ( .A(A[671]), .B(n733), .Z(n3108) );
  NANDN U3463 ( .A(n733), .B(A[671]), .Z(n3106) );
  AND U3464 ( .A(n3109), .B(n3110), .Z(n733) );
  NANDN U3465 ( .A(B[670]), .B(n3111), .Z(n3110) );
  NANDN U3466 ( .A(A[670]), .B(n735), .Z(n3111) );
  NANDN U3467 ( .A(n735), .B(A[670]), .Z(n3109) );
  AND U3468 ( .A(n3112), .B(n3113), .Z(n735) );
  NANDN U3469 ( .A(B[669]), .B(n3114), .Z(n3113) );
  NANDN U3470 ( .A(A[669]), .B(n739), .Z(n3114) );
  NANDN U3471 ( .A(n739), .B(A[669]), .Z(n3112) );
  AND U3472 ( .A(n3115), .B(n3116), .Z(n739) );
  NANDN U3473 ( .A(B[668]), .B(n3117), .Z(n3116) );
  NANDN U3474 ( .A(A[668]), .B(n741), .Z(n3117) );
  NANDN U3475 ( .A(n741), .B(A[668]), .Z(n3115) );
  AND U3476 ( .A(n3118), .B(n3119), .Z(n741) );
  NANDN U3477 ( .A(B[667]), .B(n3120), .Z(n3119) );
  NANDN U3478 ( .A(A[667]), .B(n743), .Z(n3120) );
  NANDN U3479 ( .A(n743), .B(A[667]), .Z(n3118) );
  AND U3480 ( .A(n3121), .B(n3122), .Z(n743) );
  NANDN U3481 ( .A(B[666]), .B(n3123), .Z(n3122) );
  NANDN U3482 ( .A(A[666]), .B(n745), .Z(n3123) );
  NANDN U3483 ( .A(n745), .B(A[666]), .Z(n3121) );
  AND U3484 ( .A(n3124), .B(n3125), .Z(n745) );
  NANDN U3485 ( .A(B[665]), .B(n3126), .Z(n3125) );
  NANDN U3486 ( .A(A[665]), .B(n747), .Z(n3126) );
  NANDN U3487 ( .A(n747), .B(A[665]), .Z(n3124) );
  AND U3488 ( .A(n3127), .B(n3128), .Z(n747) );
  NANDN U3489 ( .A(B[664]), .B(n3129), .Z(n3128) );
  NANDN U3490 ( .A(A[664]), .B(n749), .Z(n3129) );
  NANDN U3491 ( .A(n749), .B(A[664]), .Z(n3127) );
  AND U3492 ( .A(n3130), .B(n3131), .Z(n749) );
  NANDN U3493 ( .A(B[663]), .B(n3132), .Z(n3131) );
  NANDN U3494 ( .A(A[663]), .B(n751), .Z(n3132) );
  NANDN U3495 ( .A(n751), .B(A[663]), .Z(n3130) );
  AND U3496 ( .A(n3133), .B(n3134), .Z(n751) );
  NANDN U3497 ( .A(B[662]), .B(n3135), .Z(n3134) );
  NANDN U3498 ( .A(A[662]), .B(n753), .Z(n3135) );
  NANDN U3499 ( .A(n753), .B(A[662]), .Z(n3133) );
  AND U3500 ( .A(n3136), .B(n3137), .Z(n753) );
  NANDN U3501 ( .A(B[661]), .B(n3138), .Z(n3137) );
  NANDN U3502 ( .A(A[661]), .B(n755), .Z(n3138) );
  NANDN U3503 ( .A(n755), .B(A[661]), .Z(n3136) );
  AND U3504 ( .A(n3139), .B(n3140), .Z(n755) );
  NANDN U3505 ( .A(B[660]), .B(n3141), .Z(n3140) );
  NANDN U3506 ( .A(A[660]), .B(n757), .Z(n3141) );
  NANDN U3507 ( .A(n757), .B(A[660]), .Z(n3139) );
  AND U3508 ( .A(n3142), .B(n3143), .Z(n757) );
  NANDN U3509 ( .A(B[659]), .B(n3144), .Z(n3143) );
  NANDN U3510 ( .A(A[659]), .B(n761), .Z(n3144) );
  NANDN U3511 ( .A(n761), .B(A[659]), .Z(n3142) );
  AND U3512 ( .A(n3145), .B(n3146), .Z(n761) );
  NANDN U3513 ( .A(B[658]), .B(n3147), .Z(n3146) );
  NANDN U3514 ( .A(A[658]), .B(n763), .Z(n3147) );
  NANDN U3515 ( .A(n763), .B(A[658]), .Z(n3145) );
  AND U3516 ( .A(n3148), .B(n3149), .Z(n763) );
  NANDN U3517 ( .A(B[657]), .B(n3150), .Z(n3149) );
  NANDN U3518 ( .A(A[657]), .B(n765), .Z(n3150) );
  NANDN U3519 ( .A(n765), .B(A[657]), .Z(n3148) );
  AND U3520 ( .A(n3151), .B(n3152), .Z(n765) );
  NANDN U3521 ( .A(B[656]), .B(n3153), .Z(n3152) );
  NANDN U3522 ( .A(A[656]), .B(n767), .Z(n3153) );
  NANDN U3523 ( .A(n767), .B(A[656]), .Z(n3151) );
  AND U3524 ( .A(n3154), .B(n3155), .Z(n767) );
  NANDN U3525 ( .A(B[655]), .B(n3156), .Z(n3155) );
  NANDN U3526 ( .A(A[655]), .B(n769), .Z(n3156) );
  NANDN U3527 ( .A(n769), .B(A[655]), .Z(n3154) );
  AND U3528 ( .A(n3157), .B(n3158), .Z(n769) );
  NANDN U3529 ( .A(B[654]), .B(n3159), .Z(n3158) );
  NANDN U3530 ( .A(A[654]), .B(n771), .Z(n3159) );
  NANDN U3531 ( .A(n771), .B(A[654]), .Z(n3157) );
  AND U3532 ( .A(n3160), .B(n3161), .Z(n771) );
  NANDN U3533 ( .A(B[653]), .B(n3162), .Z(n3161) );
  NANDN U3534 ( .A(A[653]), .B(n773), .Z(n3162) );
  NANDN U3535 ( .A(n773), .B(A[653]), .Z(n3160) );
  AND U3536 ( .A(n3163), .B(n3164), .Z(n773) );
  NANDN U3537 ( .A(B[652]), .B(n3165), .Z(n3164) );
  NANDN U3538 ( .A(A[652]), .B(n775), .Z(n3165) );
  NANDN U3539 ( .A(n775), .B(A[652]), .Z(n3163) );
  AND U3540 ( .A(n3166), .B(n3167), .Z(n775) );
  NANDN U3541 ( .A(B[651]), .B(n3168), .Z(n3167) );
  NANDN U3542 ( .A(A[651]), .B(n777), .Z(n3168) );
  NANDN U3543 ( .A(n777), .B(A[651]), .Z(n3166) );
  AND U3544 ( .A(n3169), .B(n3170), .Z(n777) );
  NANDN U3545 ( .A(B[650]), .B(n3171), .Z(n3170) );
  NANDN U3546 ( .A(A[650]), .B(n779), .Z(n3171) );
  NANDN U3547 ( .A(n779), .B(A[650]), .Z(n3169) );
  AND U3548 ( .A(n3172), .B(n3173), .Z(n779) );
  NANDN U3549 ( .A(B[649]), .B(n3174), .Z(n3173) );
  NANDN U3550 ( .A(A[649]), .B(n783), .Z(n3174) );
  NANDN U3551 ( .A(n783), .B(A[649]), .Z(n3172) );
  AND U3552 ( .A(n3175), .B(n3176), .Z(n783) );
  NANDN U3553 ( .A(B[648]), .B(n3177), .Z(n3176) );
  NANDN U3554 ( .A(A[648]), .B(n785), .Z(n3177) );
  NANDN U3555 ( .A(n785), .B(A[648]), .Z(n3175) );
  AND U3556 ( .A(n3178), .B(n3179), .Z(n785) );
  NANDN U3557 ( .A(B[647]), .B(n3180), .Z(n3179) );
  NANDN U3558 ( .A(A[647]), .B(n787), .Z(n3180) );
  NANDN U3559 ( .A(n787), .B(A[647]), .Z(n3178) );
  AND U3560 ( .A(n3181), .B(n3182), .Z(n787) );
  NANDN U3561 ( .A(B[646]), .B(n3183), .Z(n3182) );
  NANDN U3562 ( .A(A[646]), .B(n789), .Z(n3183) );
  NANDN U3563 ( .A(n789), .B(A[646]), .Z(n3181) );
  AND U3564 ( .A(n3184), .B(n3185), .Z(n789) );
  NANDN U3565 ( .A(B[645]), .B(n3186), .Z(n3185) );
  NANDN U3566 ( .A(A[645]), .B(n791), .Z(n3186) );
  NANDN U3567 ( .A(n791), .B(A[645]), .Z(n3184) );
  AND U3568 ( .A(n3187), .B(n3188), .Z(n791) );
  NANDN U3569 ( .A(B[644]), .B(n3189), .Z(n3188) );
  NANDN U3570 ( .A(A[644]), .B(n793), .Z(n3189) );
  NANDN U3571 ( .A(n793), .B(A[644]), .Z(n3187) );
  AND U3572 ( .A(n3190), .B(n3191), .Z(n793) );
  NANDN U3573 ( .A(B[643]), .B(n3192), .Z(n3191) );
  NANDN U3574 ( .A(A[643]), .B(n795), .Z(n3192) );
  NANDN U3575 ( .A(n795), .B(A[643]), .Z(n3190) );
  AND U3576 ( .A(n3193), .B(n3194), .Z(n795) );
  NANDN U3577 ( .A(B[642]), .B(n3195), .Z(n3194) );
  NANDN U3578 ( .A(A[642]), .B(n797), .Z(n3195) );
  NANDN U3579 ( .A(n797), .B(A[642]), .Z(n3193) );
  AND U3580 ( .A(n3196), .B(n3197), .Z(n797) );
  NANDN U3581 ( .A(B[641]), .B(n3198), .Z(n3197) );
  NANDN U3582 ( .A(A[641]), .B(n799), .Z(n3198) );
  NANDN U3583 ( .A(n799), .B(A[641]), .Z(n3196) );
  AND U3584 ( .A(n3199), .B(n3200), .Z(n799) );
  NANDN U3585 ( .A(B[640]), .B(n3201), .Z(n3200) );
  NANDN U3586 ( .A(A[640]), .B(n801), .Z(n3201) );
  NANDN U3587 ( .A(n801), .B(A[640]), .Z(n3199) );
  AND U3588 ( .A(n3202), .B(n3203), .Z(n801) );
  NANDN U3589 ( .A(B[639]), .B(n3204), .Z(n3203) );
  NANDN U3590 ( .A(A[639]), .B(n805), .Z(n3204) );
  NANDN U3591 ( .A(n805), .B(A[639]), .Z(n3202) );
  AND U3592 ( .A(n3205), .B(n3206), .Z(n805) );
  NANDN U3593 ( .A(B[638]), .B(n3207), .Z(n3206) );
  NANDN U3594 ( .A(A[638]), .B(n807), .Z(n3207) );
  NANDN U3595 ( .A(n807), .B(A[638]), .Z(n3205) );
  AND U3596 ( .A(n3208), .B(n3209), .Z(n807) );
  NANDN U3597 ( .A(B[637]), .B(n3210), .Z(n3209) );
  NANDN U3598 ( .A(A[637]), .B(n809), .Z(n3210) );
  NANDN U3599 ( .A(n809), .B(A[637]), .Z(n3208) );
  AND U3600 ( .A(n3211), .B(n3212), .Z(n809) );
  NANDN U3601 ( .A(B[636]), .B(n3213), .Z(n3212) );
  NANDN U3602 ( .A(A[636]), .B(n811), .Z(n3213) );
  NANDN U3603 ( .A(n811), .B(A[636]), .Z(n3211) );
  AND U3604 ( .A(n3214), .B(n3215), .Z(n811) );
  NANDN U3605 ( .A(B[635]), .B(n3216), .Z(n3215) );
  NANDN U3606 ( .A(A[635]), .B(n813), .Z(n3216) );
  NANDN U3607 ( .A(n813), .B(A[635]), .Z(n3214) );
  AND U3608 ( .A(n3217), .B(n3218), .Z(n813) );
  NANDN U3609 ( .A(B[634]), .B(n3219), .Z(n3218) );
  NANDN U3610 ( .A(A[634]), .B(n815), .Z(n3219) );
  NANDN U3611 ( .A(n815), .B(A[634]), .Z(n3217) );
  AND U3612 ( .A(n3220), .B(n3221), .Z(n815) );
  NANDN U3613 ( .A(B[633]), .B(n3222), .Z(n3221) );
  NANDN U3614 ( .A(A[633]), .B(n817), .Z(n3222) );
  NANDN U3615 ( .A(n817), .B(A[633]), .Z(n3220) );
  AND U3616 ( .A(n3223), .B(n3224), .Z(n817) );
  NANDN U3617 ( .A(B[632]), .B(n3225), .Z(n3224) );
  NANDN U3618 ( .A(A[632]), .B(n819), .Z(n3225) );
  NANDN U3619 ( .A(n819), .B(A[632]), .Z(n3223) );
  AND U3620 ( .A(n3226), .B(n3227), .Z(n819) );
  NANDN U3621 ( .A(B[631]), .B(n3228), .Z(n3227) );
  NANDN U3622 ( .A(A[631]), .B(n821), .Z(n3228) );
  NANDN U3623 ( .A(n821), .B(A[631]), .Z(n3226) );
  AND U3624 ( .A(n3229), .B(n3230), .Z(n821) );
  NANDN U3625 ( .A(B[630]), .B(n3231), .Z(n3230) );
  NANDN U3626 ( .A(A[630]), .B(n823), .Z(n3231) );
  NANDN U3627 ( .A(n823), .B(A[630]), .Z(n3229) );
  AND U3628 ( .A(n3232), .B(n3233), .Z(n823) );
  NANDN U3629 ( .A(B[629]), .B(n3234), .Z(n3233) );
  NANDN U3630 ( .A(A[629]), .B(n827), .Z(n3234) );
  NANDN U3631 ( .A(n827), .B(A[629]), .Z(n3232) );
  AND U3632 ( .A(n3235), .B(n3236), .Z(n827) );
  NANDN U3633 ( .A(B[628]), .B(n3237), .Z(n3236) );
  NANDN U3634 ( .A(A[628]), .B(n829), .Z(n3237) );
  NANDN U3635 ( .A(n829), .B(A[628]), .Z(n3235) );
  AND U3636 ( .A(n3238), .B(n3239), .Z(n829) );
  NANDN U3637 ( .A(B[627]), .B(n3240), .Z(n3239) );
  NANDN U3638 ( .A(A[627]), .B(n831), .Z(n3240) );
  NANDN U3639 ( .A(n831), .B(A[627]), .Z(n3238) );
  AND U3640 ( .A(n3241), .B(n3242), .Z(n831) );
  NANDN U3641 ( .A(B[626]), .B(n3243), .Z(n3242) );
  NANDN U3642 ( .A(A[626]), .B(n833), .Z(n3243) );
  NANDN U3643 ( .A(n833), .B(A[626]), .Z(n3241) );
  AND U3644 ( .A(n3244), .B(n3245), .Z(n833) );
  NANDN U3645 ( .A(B[625]), .B(n3246), .Z(n3245) );
  NANDN U3646 ( .A(A[625]), .B(n835), .Z(n3246) );
  NANDN U3647 ( .A(n835), .B(A[625]), .Z(n3244) );
  AND U3648 ( .A(n3247), .B(n3248), .Z(n835) );
  NANDN U3649 ( .A(B[624]), .B(n3249), .Z(n3248) );
  NANDN U3650 ( .A(A[624]), .B(n837), .Z(n3249) );
  NANDN U3651 ( .A(n837), .B(A[624]), .Z(n3247) );
  AND U3652 ( .A(n3250), .B(n3251), .Z(n837) );
  NANDN U3653 ( .A(B[623]), .B(n3252), .Z(n3251) );
  NANDN U3654 ( .A(A[623]), .B(n839), .Z(n3252) );
  NANDN U3655 ( .A(n839), .B(A[623]), .Z(n3250) );
  AND U3656 ( .A(n3253), .B(n3254), .Z(n839) );
  NANDN U3657 ( .A(B[622]), .B(n3255), .Z(n3254) );
  NANDN U3658 ( .A(A[622]), .B(n841), .Z(n3255) );
  NANDN U3659 ( .A(n841), .B(A[622]), .Z(n3253) );
  AND U3660 ( .A(n3256), .B(n3257), .Z(n841) );
  NANDN U3661 ( .A(B[621]), .B(n3258), .Z(n3257) );
  NANDN U3662 ( .A(A[621]), .B(n843), .Z(n3258) );
  NANDN U3663 ( .A(n843), .B(A[621]), .Z(n3256) );
  AND U3664 ( .A(n3259), .B(n3260), .Z(n843) );
  NANDN U3665 ( .A(B[620]), .B(n3261), .Z(n3260) );
  NANDN U3666 ( .A(A[620]), .B(n845), .Z(n3261) );
  NANDN U3667 ( .A(n845), .B(A[620]), .Z(n3259) );
  AND U3668 ( .A(n3262), .B(n3263), .Z(n845) );
  NANDN U3669 ( .A(B[619]), .B(n3264), .Z(n3263) );
  NANDN U3670 ( .A(A[619]), .B(n849), .Z(n3264) );
  NANDN U3671 ( .A(n849), .B(A[619]), .Z(n3262) );
  AND U3672 ( .A(n3265), .B(n3266), .Z(n849) );
  NANDN U3673 ( .A(B[618]), .B(n3267), .Z(n3266) );
  NANDN U3674 ( .A(A[618]), .B(n851), .Z(n3267) );
  NANDN U3675 ( .A(n851), .B(A[618]), .Z(n3265) );
  AND U3676 ( .A(n3268), .B(n3269), .Z(n851) );
  NANDN U3677 ( .A(B[617]), .B(n3270), .Z(n3269) );
  NANDN U3678 ( .A(A[617]), .B(n853), .Z(n3270) );
  NANDN U3679 ( .A(n853), .B(A[617]), .Z(n3268) );
  AND U3680 ( .A(n3271), .B(n3272), .Z(n853) );
  NANDN U3681 ( .A(B[616]), .B(n3273), .Z(n3272) );
  NANDN U3682 ( .A(A[616]), .B(n855), .Z(n3273) );
  NANDN U3683 ( .A(n855), .B(A[616]), .Z(n3271) );
  AND U3684 ( .A(n3274), .B(n3275), .Z(n855) );
  NANDN U3685 ( .A(B[615]), .B(n3276), .Z(n3275) );
  NANDN U3686 ( .A(A[615]), .B(n857), .Z(n3276) );
  NANDN U3687 ( .A(n857), .B(A[615]), .Z(n3274) );
  AND U3688 ( .A(n3277), .B(n3278), .Z(n857) );
  NANDN U3689 ( .A(B[614]), .B(n3279), .Z(n3278) );
  NANDN U3690 ( .A(A[614]), .B(n859), .Z(n3279) );
  NANDN U3691 ( .A(n859), .B(A[614]), .Z(n3277) );
  AND U3692 ( .A(n3280), .B(n3281), .Z(n859) );
  NANDN U3693 ( .A(B[613]), .B(n3282), .Z(n3281) );
  NANDN U3694 ( .A(A[613]), .B(n861), .Z(n3282) );
  NANDN U3695 ( .A(n861), .B(A[613]), .Z(n3280) );
  AND U3696 ( .A(n3283), .B(n3284), .Z(n861) );
  NANDN U3697 ( .A(B[612]), .B(n3285), .Z(n3284) );
  NANDN U3698 ( .A(A[612]), .B(n863), .Z(n3285) );
  NANDN U3699 ( .A(n863), .B(A[612]), .Z(n3283) );
  AND U3700 ( .A(n3286), .B(n3287), .Z(n863) );
  NANDN U3701 ( .A(B[611]), .B(n3288), .Z(n3287) );
  NANDN U3702 ( .A(A[611]), .B(n865), .Z(n3288) );
  NANDN U3703 ( .A(n865), .B(A[611]), .Z(n3286) );
  AND U3704 ( .A(n3289), .B(n3290), .Z(n865) );
  NANDN U3705 ( .A(B[610]), .B(n3291), .Z(n3290) );
  NANDN U3706 ( .A(A[610]), .B(n867), .Z(n3291) );
  NANDN U3707 ( .A(n867), .B(A[610]), .Z(n3289) );
  AND U3708 ( .A(n3292), .B(n3293), .Z(n867) );
  NANDN U3709 ( .A(B[609]), .B(n3294), .Z(n3293) );
  NANDN U3710 ( .A(A[609]), .B(n871), .Z(n3294) );
  NANDN U3711 ( .A(n871), .B(A[609]), .Z(n3292) );
  AND U3712 ( .A(n3295), .B(n3296), .Z(n871) );
  NANDN U3713 ( .A(B[608]), .B(n3297), .Z(n3296) );
  NANDN U3714 ( .A(A[608]), .B(n873), .Z(n3297) );
  NANDN U3715 ( .A(n873), .B(A[608]), .Z(n3295) );
  AND U3716 ( .A(n3298), .B(n3299), .Z(n873) );
  NANDN U3717 ( .A(B[607]), .B(n3300), .Z(n3299) );
  NANDN U3718 ( .A(A[607]), .B(n875), .Z(n3300) );
  NANDN U3719 ( .A(n875), .B(A[607]), .Z(n3298) );
  AND U3720 ( .A(n3301), .B(n3302), .Z(n875) );
  NANDN U3721 ( .A(B[606]), .B(n3303), .Z(n3302) );
  NANDN U3722 ( .A(A[606]), .B(n877), .Z(n3303) );
  NANDN U3723 ( .A(n877), .B(A[606]), .Z(n3301) );
  AND U3724 ( .A(n3304), .B(n3305), .Z(n877) );
  NANDN U3725 ( .A(B[605]), .B(n3306), .Z(n3305) );
  NANDN U3726 ( .A(A[605]), .B(n879), .Z(n3306) );
  NANDN U3727 ( .A(n879), .B(A[605]), .Z(n3304) );
  AND U3728 ( .A(n3307), .B(n3308), .Z(n879) );
  NANDN U3729 ( .A(B[604]), .B(n3309), .Z(n3308) );
  NANDN U3730 ( .A(A[604]), .B(n881), .Z(n3309) );
  NANDN U3731 ( .A(n881), .B(A[604]), .Z(n3307) );
  AND U3732 ( .A(n3310), .B(n3311), .Z(n881) );
  NANDN U3733 ( .A(B[603]), .B(n3312), .Z(n3311) );
  NANDN U3734 ( .A(A[603]), .B(n883), .Z(n3312) );
  NANDN U3735 ( .A(n883), .B(A[603]), .Z(n3310) );
  AND U3736 ( .A(n3313), .B(n3314), .Z(n883) );
  NANDN U3737 ( .A(B[602]), .B(n3315), .Z(n3314) );
  NANDN U3738 ( .A(A[602]), .B(n885), .Z(n3315) );
  NANDN U3739 ( .A(n885), .B(A[602]), .Z(n3313) );
  AND U3740 ( .A(n3316), .B(n3317), .Z(n885) );
  NANDN U3741 ( .A(B[601]), .B(n3318), .Z(n3317) );
  NANDN U3742 ( .A(A[601]), .B(n887), .Z(n3318) );
  NANDN U3743 ( .A(n887), .B(A[601]), .Z(n3316) );
  AND U3744 ( .A(n3319), .B(n3320), .Z(n887) );
  NANDN U3745 ( .A(B[600]), .B(n3321), .Z(n3320) );
  NANDN U3746 ( .A(A[600]), .B(n889), .Z(n3321) );
  NANDN U3747 ( .A(n889), .B(A[600]), .Z(n3319) );
  AND U3748 ( .A(n3322), .B(n3323), .Z(n889) );
  NANDN U3749 ( .A(B[599]), .B(n3324), .Z(n3323) );
  NANDN U3750 ( .A(A[599]), .B(n895), .Z(n3324) );
  NANDN U3751 ( .A(n895), .B(A[599]), .Z(n3322) );
  AND U3752 ( .A(n3325), .B(n3326), .Z(n895) );
  NANDN U3753 ( .A(B[598]), .B(n3327), .Z(n3326) );
  NANDN U3754 ( .A(A[598]), .B(n897), .Z(n3327) );
  NANDN U3755 ( .A(n897), .B(A[598]), .Z(n3325) );
  AND U3756 ( .A(n3328), .B(n3329), .Z(n897) );
  NANDN U3757 ( .A(B[597]), .B(n3330), .Z(n3329) );
  NANDN U3758 ( .A(A[597]), .B(n899), .Z(n3330) );
  NANDN U3759 ( .A(n899), .B(A[597]), .Z(n3328) );
  AND U3760 ( .A(n3331), .B(n3332), .Z(n899) );
  NANDN U3761 ( .A(B[596]), .B(n3333), .Z(n3332) );
  NANDN U3762 ( .A(A[596]), .B(n901), .Z(n3333) );
  NANDN U3763 ( .A(n901), .B(A[596]), .Z(n3331) );
  AND U3764 ( .A(n3334), .B(n3335), .Z(n901) );
  NANDN U3765 ( .A(B[595]), .B(n3336), .Z(n3335) );
  NANDN U3766 ( .A(A[595]), .B(n903), .Z(n3336) );
  NANDN U3767 ( .A(n903), .B(A[595]), .Z(n3334) );
  AND U3768 ( .A(n3337), .B(n3338), .Z(n903) );
  NANDN U3769 ( .A(B[594]), .B(n3339), .Z(n3338) );
  NANDN U3770 ( .A(A[594]), .B(n905), .Z(n3339) );
  NANDN U3771 ( .A(n905), .B(A[594]), .Z(n3337) );
  AND U3772 ( .A(n3340), .B(n3341), .Z(n905) );
  NANDN U3773 ( .A(B[593]), .B(n3342), .Z(n3341) );
  NANDN U3774 ( .A(A[593]), .B(n907), .Z(n3342) );
  NANDN U3775 ( .A(n907), .B(A[593]), .Z(n3340) );
  AND U3776 ( .A(n3343), .B(n3344), .Z(n907) );
  NANDN U3777 ( .A(B[592]), .B(n3345), .Z(n3344) );
  NANDN U3778 ( .A(A[592]), .B(n909), .Z(n3345) );
  NANDN U3779 ( .A(n909), .B(A[592]), .Z(n3343) );
  AND U3780 ( .A(n3346), .B(n3347), .Z(n909) );
  NANDN U3781 ( .A(B[591]), .B(n3348), .Z(n3347) );
  NANDN U3782 ( .A(A[591]), .B(n911), .Z(n3348) );
  NANDN U3783 ( .A(n911), .B(A[591]), .Z(n3346) );
  AND U3784 ( .A(n3349), .B(n3350), .Z(n911) );
  NANDN U3785 ( .A(B[590]), .B(n3351), .Z(n3350) );
  NANDN U3786 ( .A(A[590]), .B(n913), .Z(n3351) );
  NANDN U3787 ( .A(n913), .B(A[590]), .Z(n3349) );
  AND U3788 ( .A(n3352), .B(n3353), .Z(n913) );
  NANDN U3789 ( .A(B[589]), .B(n3354), .Z(n3353) );
  NANDN U3790 ( .A(A[589]), .B(n917), .Z(n3354) );
  NANDN U3791 ( .A(n917), .B(A[589]), .Z(n3352) );
  AND U3792 ( .A(n3355), .B(n3356), .Z(n917) );
  NANDN U3793 ( .A(B[588]), .B(n3357), .Z(n3356) );
  NANDN U3794 ( .A(A[588]), .B(n919), .Z(n3357) );
  NANDN U3795 ( .A(n919), .B(A[588]), .Z(n3355) );
  AND U3796 ( .A(n3358), .B(n3359), .Z(n919) );
  NANDN U3797 ( .A(B[587]), .B(n3360), .Z(n3359) );
  NANDN U3798 ( .A(A[587]), .B(n921), .Z(n3360) );
  NANDN U3799 ( .A(n921), .B(A[587]), .Z(n3358) );
  AND U3800 ( .A(n3361), .B(n3362), .Z(n921) );
  NANDN U3801 ( .A(B[586]), .B(n3363), .Z(n3362) );
  NANDN U3802 ( .A(A[586]), .B(n923), .Z(n3363) );
  NANDN U3803 ( .A(n923), .B(A[586]), .Z(n3361) );
  AND U3804 ( .A(n3364), .B(n3365), .Z(n923) );
  NANDN U3805 ( .A(B[585]), .B(n3366), .Z(n3365) );
  NANDN U3806 ( .A(A[585]), .B(n925), .Z(n3366) );
  NANDN U3807 ( .A(n925), .B(A[585]), .Z(n3364) );
  AND U3808 ( .A(n3367), .B(n3368), .Z(n925) );
  NANDN U3809 ( .A(B[584]), .B(n3369), .Z(n3368) );
  NANDN U3810 ( .A(A[584]), .B(n927), .Z(n3369) );
  NANDN U3811 ( .A(n927), .B(A[584]), .Z(n3367) );
  AND U3812 ( .A(n3370), .B(n3371), .Z(n927) );
  NANDN U3813 ( .A(B[583]), .B(n3372), .Z(n3371) );
  NANDN U3814 ( .A(A[583]), .B(n929), .Z(n3372) );
  NANDN U3815 ( .A(n929), .B(A[583]), .Z(n3370) );
  AND U3816 ( .A(n3373), .B(n3374), .Z(n929) );
  NANDN U3817 ( .A(B[582]), .B(n3375), .Z(n3374) );
  NANDN U3818 ( .A(A[582]), .B(n931), .Z(n3375) );
  NANDN U3819 ( .A(n931), .B(A[582]), .Z(n3373) );
  AND U3820 ( .A(n3376), .B(n3377), .Z(n931) );
  NANDN U3821 ( .A(B[581]), .B(n3378), .Z(n3377) );
  NANDN U3822 ( .A(A[581]), .B(n933), .Z(n3378) );
  NANDN U3823 ( .A(n933), .B(A[581]), .Z(n3376) );
  AND U3824 ( .A(n3379), .B(n3380), .Z(n933) );
  NANDN U3825 ( .A(B[580]), .B(n3381), .Z(n3380) );
  NANDN U3826 ( .A(A[580]), .B(n935), .Z(n3381) );
  NANDN U3827 ( .A(n935), .B(A[580]), .Z(n3379) );
  AND U3828 ( .A(n3382), .B(n3383), .Z(n935) );
  NANDN U3829 ( .A(B[579]), .B(n3384), .Z(n3383) );
  NANDN U3830 ( .A(A[579]), .B(n939), .Z(n3384) );
  NANDN U3831 ( .A(n939), .B(A[579]), .Z(n3382) );
  AND U3832 ( .A(n3385), .B(n3386), .Z(n939) );
  NANDN U3833 ( .A(B[578]), .B(n3387), .Z(n3386) );
  NANDN U3834 ( .A(A[578]), .B(n941), .Z(n3387) );
  NANDN U3835 ( .A(n941), .B(A[578]), .Z(n3385) );
  AND U3836 ( .A(n3388), .B(n3389), .Z(n941) );
  NANDN U3837 ( .A(B[577]), .B(n3390), .Z(n3389) );
  NANDN U3838 ( .A(A[577]), .B(n943), .Z(n3390) );
  NANDN U3839 ( .A(n943), .B(A[577]), .Z(n3388) );
  AND U3840 ( .A(n3391), .B(n3392), .Z(n943) );
  NANDN U3841 ( .A(B[576]), .B(n3393), .Z(n3392) );
  NANDN U3842 ( .A(A[576]), .B(n945), .Z(n3393) );
  NANDN U3843 ( .A(n945), .B(A[576]), .Z(n3391) );
  AND U3844 ( .A(n3394), .B(n3395), .Z(n945) );
  NANDN U3845 ( .A(B[575]), .B(n3396), .Z(n3395) );
  NANDN U3846 ( .A(A[575]), .B(n947), .Z(n3396) );
  NANDN U3847 ( .A(n947), .B(A[575]), .Z(n3394) );
  AND U3848 ( .A(n3397), .B(n3398), .Z(n947) );
  NANDN U3849 ( .A(B[574]), .B(n3399), .Z(n3398) );
  NANDN U3850 ( .A(A[574]), .B(n949), .Z(n3399) );
  NANDN U3851 ( .A(n949), .B(A[574]), .Z(n3397) );
  AND U3852 ( .A(n3400), .B(n3401), .Z(n949) );
  NANDN U3853 ( .A(B[573]), .B(n3402), .Z(n3401) );
  NANDN U3854 ( .A(A[573]), .B(n951), .Z(n3402) );
  NANDN U3855 ( .A(n951), .B(A[573]), .Z(n3400) );
  AND U3856 ( .A(n3403), .B(n3404), .Z(n951) );
  NANDN U3857 ( .A(B[572]), .B(n3405), .Z(n3404) );
  NANDN U3858 ( .A(A[572]), .B(n953), .Z(n3405) );
  NANDN U3859 ( .A(n953), .B(A[572]), .Z(n3403) );
  AND U3860 ( .A(n3406), .B(n3407), .Z(n953) );
  NANDN U3861 ( .A(B[571]), .B(n3408), .Z(n3407) );
  NANDN U3862 ( .A(A[571]), .B(n955), .Z(n3408) );
  NANDN U3863 ( .A(n955), .B(A[571]), .Z(n3406) );
  AND U3864 ( .A(n3409), .B(n3410), .Z(n955) );
  NANDN U3865 ( .A(B[570]), .B(n3411), .Z(n3410) );
  NANDN U3866 ( .A(A[570]), .B(n957), .Z(n3411) );
  NANDN U3867 ( .A(n957), .B(A[570]), .Z(n3409) );
  AND U3868 ( .A(n3412), .B(n3413), .Z(n957) );
  NANDN U3869 ( .A(B[569]), .B(n3414), .Z(n3413) );
  NANDN U3870 ( .A(A[569]), .B(n961), .Z(n3414) );
  NANDN U3871 ( .A(n961), .B(A[569]), .Z(n3412) );
  AND U3872 ( .A(n3415), .B(n3416), .Z(n961) );
  NANDN U3873 ( .A(B[568]), .B(n3417), .Z(n3416) );
  NANDN U3874 ( .A(A[568]), .B(n963), .Z(n3417) );
  NANDN U3875 ( .A(n963), .B(A[568]), .Z(n3415) );
  AND U3876 ( .A(n3418), .B(n3419), .Z(n963) );
  NANDN U3877 ( .A(B[567]), .B(n3420), .Z(n3419) );
  NANDN U3878 ( .A(A[567]), .B(n965), .Z(n3420) );
  NANDN U3879 ( .A(n965), .B(A[567]), .Z(n3418) );
  AND U3880 ( .A(n3421), .B(n3422), .Z(n965) );
  NANDN U3881 ( .A(B[566]), .B(n3423), .Z(n3422) );
  NANDN U3882 ( .A(A[566]), .B(n967), .Z(n3423) );
  NANDN U3883 ( .A(n967), .B(A[566]), .Z(n3421) );
  AND U3884 ( .A(n3424), .B(n3425), .Z(n967) );
  NANDN U3885 ( .A(B[565]), .B(n3426), .Z(n3425) );
  NANDN U3886 ( .A(A[565]), .B(n969), .Z(n3426) );
  NANDN U3887 ( .A(n969), .B(A[565]), .Z(n3424) );
  AND U3888 ( .A(n3427), .B(n3428), .Z(n969) );
  NANDN U3889 ( .A(B[564]), .B(n3429), .Z(n3428) );
  NANDN U3890 ( .A(A[564]), .B(n971), .Z(n3429) );
  NANDN U3891 ( .A(n971), .B(A[564]), .Z(n3427) );
  AND U3892 ( .A(n3430), .B(n3431), .Z(n971) );
  NANDN U3893 ( .A(B[563]), .B(n3432), .Z(n3431) );
  NANDN U3894 ( .A(A[563]), .B(n973), .Z(n3432) );
  NANDN U3895 ( .A(n973), .B(A[563]), .Z(n3430) );
  AND U3896 ( .A(n3433), .B(n3434), .Z(n973) );
  NANDN U3897 ( .A(B[562]), .B(n3435), .Z(n3434) );
  NANDN U3898 ( .A(A[562]), .B(n975), .Z(n3435) );
  NANDN U3899 ( .A(n975), .B(A[562]), .Z(n3433) );
  AND U3900 ( .A(n3436), .B(n3437), .Z(n975) );
  NANDN U3901 ( .A(B[561]), .B(n3438), .Z(n3437) );
  NANDN U3902 ( .A(A[561]), .B(n977), .Z(n3438) );
  NANDN U3903 ( .A(n977), .B(A[561]), .Z(n3436) );
  AND U3904 ( .A(n3439), .B(n3440), .Z(n977) );
  NANDN U3905 ( .A(B[560]), .B(n3441), .Z(n3440) );
  NANDN U3906 ( .A(A[560]), .B(n979), .Z(n3441) );
  NANDN U3907 ( .A(n979), .B(A[560]), .Z(n3439) );
  AND U3908 ( .A(n3442), .B(n3443), .Z(n979) );
  NANDN U3909 ( .A(B[559]), .B(n3444), .Z(n3443) );
  NANDN U3910 ( .A(A[559]), .B(n983), .Z(n3444) );
  NANDN U3911 ( .A(n983), .B(A[559]), .Z(n3442) );
  AND U3912 ( .A(n3445), .B(n3446), .Z(n983) );
  NANDN U3913 ( .A(B[558]), .B(n3447), .Z(n3446) );
  NANDN U3914 ( .A(A[558]), .B(n985), .Z(n3447) );
  NANDN U3915 ( .A(n985), .B(A[558]), .Z(n3445) );
  AND U3916 ( .A(n3448), .B(n3449), .Z(n985) );
  NANDN U3917 ( .A(B[557]), .B(n3450), .Z(n3449) );
  NANDN U3918 ( .A(A[557]), .B(n987), .Z(n3450) );
  NANDN U3919 ( .A(n987), .B(A[557]), .Z(n3448) );
  AND U3920 ( .A(n3451), .B(n3452), .Z(n987) );
  NANDN U3921 ( .A(B[556]), .B(n3453), .Z(n3452) );
  NANDN U3922 ( .A(A[556]), .B(n989), .Z(n3453) );
  NANDN U3923 ( .A(n989), .B(A[556]), .Z(n3451) );
  AND U3924 ( .A(n3454), .B(n3455), .Z(n989) );
  NANDN U3925 ( .A(B[555]), .B(n3456), .Z(n3455) );
  NANDN U3926 ( .A(A[555]), .B(n991), .Z(n3456) );
  NANDN U3927 ( .A(n991), .B(A[555]), .Z(n3454) );
  AND U3928 ( .A(n3457), .B(n3458), .Z(n991) );
  NANDN U3929 ( .A(B[554]), .B(n3459), .Z(n3458) );
  NANDN U3930 ( .A(A[554]), .B(n993), .Z(n3459) );
  NANDN U3931 ( .A(n993), .B(A[554]), .Z(n3457) );
  AND U3932 ( .A(n3460), .B(n3461), .Z(n993) );
  NANDN U3933 ( .A(B[553]), .B(n3462), .Z(n3461) );
  NANDN U3934 ( .A(A[553]), .B(n995), .Z(n3462) );
  NANDN U3935 ( .A(n995), .B(A[553]), .Z(n3460) );
  AND U3936 ( .A(n3463), .B(n3464), .Z(n995) );
  NANDN U3937 ( .A(B[552]), .B(n3465), .Z(n3464) );
  NANDN U3938 ( .A(A[552]), .B(n997), .Z(n3465) );
  NANDN U3939 ( .A(n997), .B(A[552]), .Z(n3463) );
  AND U3940 ( .A(n3466), .B(n3467), .Z(n997) );
  NANDN U3941 ( .A(B[551]), .B(n3468), .Z(n3467) );
  NANDN U3942 ( .A(A[551]), .B(n999), .Z(n3468) );
  NANDN U3943 ( .A(n999), .B(A[551]), .Z(n3466) );
  AND U3944 ( .A(n3469), .B(n3470), .Z(n999) );
  NANDN U3945 ( .A(B[550]), .B(n3471), .Z(n3470) );
  NANDN U3946 ( .A(A[550]), .B(n1001), .Z(n3471) );
  NANDN U3947 ( .A(n1001), .B(A[550]), .Z(n3469) );
  AND U3948 ( .A(n3472), .B(n3473), .Z(n1001) );
  NANDN U3949 ( .A(B[549]), .B(n3474), .Z(n3473) );
  NANDN U3950 ( .A(A[549]), .B(n1005), .Z(n3474) );
  NANDN U3951 ( .A(n1005), .B(A[549]), .Z(n3472) );
  AND U3952 ( .A(n3475), .B(n3476), .Z(n1005) );
  NANDN U3953 ( .A(B[548]), .B(n3477), .Z(n3476) );
  NANDN U3954 ( .A(A[548]), .B(n1007), .Z(n3477) );
  NANDN U3955 ( .A(n1007), .B(A[548]), .Z(n3475) );
  AND U3956 ( .A(n3478), .B(n3479), .Z(n1007) );
  NANDN U3957 ( .A(B[547]), .B(n3480), .Z(n3479) );
  NANDN U3958 ( .A(A[547]), .B(n1009), .Z(n3480) );
  NANDN U3959 ( .A(n1009), .B(A[547]), .Z(n3478) );
  AND U3960 ( .A(n3481), .B(n3482), .Z(n1009) );
  NANDN U3961 ( .A(B[546]), .B(n3483), .Z(n3482) );
  NANDN U3962 ( .A(A[546]), .B(n1011), .Z(n3483) );
  NANDN U3963 ( .A(n1011), .B(A[546]), .Z(n3481) );
  AND U3964 ( .A(n3484), .B(n3485), .Z(n1011) );
  NANDN U3965 ( .A(B[545]), .B(n3486), .Z(n3485) );
  NANDN U3966 ( .A(A[545]), .B(n1013), .Z(n3486) );
  NANDN U3967 ( .A(n1013), .B(A[545]), .Z(n3484) );
  AND U3968 ( .A(n3487), .B(n3488), .Z(n1013) );
  NANDN U3969 ( .A(B[544]), .B(n3489), .Z(n3488) );
  NANDN U3970 ( .A(A[544]), .B(n1015), .Z(n3489) );
  NANDN U3971 ( .A(n1015), .B(A[544]), .Z(n3487) );
  AND U3972 ( .A(n3490), .B(n3491), .Z(n1015) );
  NANDN U3973 ( .A(B[543]), .B(n3492), .Z(n3491) );
  NANDN U3974 ( .A(A[543]), .B(n1017), .Z(n3492) );
  NANDN U3975 ( .A(n1017), .B(A[543]), .Z(n3490) );
  AND U3976 ( .A(n3493), .B(n3494), .Z(n1017) );
  NANDN U3977 ( .A(B[542]), .B(n3495), .Z(n3494) );
  NANDN U3978 ( .A(A[542]), .B(n1019), .Z(n3495) );
  NANDN U3979 ( .A(n1019), .B(A[542]), .Z(n3493) );
  AND U3980 ( .A(n3496), .B(n3497), .Z(n1019) );
  NANDN U3981 ( .A(B[541]), .B(n3498), .Z(n3497) );
  NANDN U3982 ( .A(A[541]), .B(n1021), .Z(n3498) );
  NANDN U3983 ( .A(n1021), .B(A[541]), .Z(n3496) );
  AND U3984 ( .A(n3499), .B(n3500), .Z(n1021) );
  NANDN U3985 ( .A(B[540]), .B(n3501), .Z(n3500) );
  NANDN U3986 ( .A(A[540]), .B(n1023), .Z(n3501) );
  NANDN U3987 ( .A(n1023), .B(A[540]), .Z(n3499) );
  AND U3988 ( .A(n3502), .B(n3503), .Z(n1023) );
  NANDN U3989 ( .A(B[539]), .B(n3504), .Z(n3503) );
  NANDN U3990 ( .A(A[539]), .B(n1027), .Z(n3504) );
  NANDN U3991 ( .A(n1027), .B(A[539]), .Z(n3502) );
  AND U3992 ( .A(n3505), .B(n3506), .Z(n1027) );
  NANDN U3993 ( .A(B[538]), .B(n3507), .Z(n3506) );
  NANDN U3994 ( .A(A[538]), .B(n1029), .Z(n3507) );
  NANDN U3995 ( .A(n1029), .B(A[538]), .Z(n3505) );
  AND U3996 ( .A(n3508), .B(n3509), .Z(n1029) );
  NANDN U3997 ( .A(B[537]), .B(n3510), .Z(n3509) );
  NANDN U3998 ( .A(A[537]), .B(n1031), .Z(n3510) );
  NANDN U3999 ( .A(n1031), .B(A[537]), .Z(n3508) );
  AND U4000 ( .A(n3511), .B(n3512), .Z(n1031) );
  NANDN U4001 ( .A(B[536]), .B(n3513), .Z(n3512) );
  NANDN U4002 ( .A(A[536]), .B(n1033), .Z(n3513) );
  NANDN U4003 ( .A(n1033), .B(A[536]), .Z(n3511) );
  AND U4004 ( .A(n3514), .B(n3515), .Z(n1033) );
  NANDN U4005 ( .A(B[535]), .B(n3516), .Z(n3515) );
  NANDN U4006 ( .A(A[535]), .B(n1035), .Z(n3516) );
  NANDN U4007 ( .A(n1035), .B(A[535]), .Z(n3514) );
  AND U4008 ( .A(n3517), .B(n3518), .Z(n1035) );
  NANDN U4009 ( .A(B[534]), .B(n3519), .Z(n3518) );
  NANDN U4010 ( .A(A[534]), .B(n1037), .Z(n3519) );
  NANDN U4011 ( .A(n1037), .B(A[534]), .Z(n3517) );
  AND U4012 ( .A(n3520), .B(n3521), .Z(n1037) );
  NANDN U4013 ( .A(B[533]), .B(n3522), .Z(n3521) );
  NANDN U4014 ( .A(A[533]), .B(n1039), .Z(n3522) );
  NANDN U4015 ( .A(n1039), .B(A[533]), .Z(n3520) );
  AND U4016 ( .A(n3523), .B(n3524), .Z(n1039) );
  NANDN U4017 ( .A(B[532]), .B(n3525), .Z(n3524) );
  NANDN U4018 ( .A(A[532]), .B(n1041), .Z(n3525) );
  NANDN U4019 ( .A(n1041), .B(A[532]), .Z(n3523) );
  AND U4020 ( .A(n3526), .B(n3527), .Z(n1041) );
  NANDN U4021 ( .A(B[531]), .B(n3528), .Z(n3527) );
  NANDN U4022 ( .A(A[531]), .B(n1043), .Z(n3528) );
  NANDN U4023 ( .A(n1043), .B(A[531]), .Z(n3526) );
  AND U4024 ( .A(n3529), .B(n3530), .Z(n1043) );
  NANDN U4025 ( .A(B[530]), .B(n3531), .Z(n3530) );
  NANDN U4026 ( .A(A[530]), .B(n1045), .Z(n3531) );
  NANDN U4027 ( .A(n1045), .B(A[530]), .Z(n3529) );
  AND U4028 ( .A(n3532), .B(n3533), .Z(n1045) );
  NANDN U4029 ( .A(B[529]), .B(n3534), .Z(n3533) );
  NANDN U4030 ( .A(A[529]), .B(n1049), .Z(n3534) );
  NANDN U4031 ( .A(n1049), .B(A[529]), .Z(n3532) );
  AND U4032 ( .A(n3535), .B(n3536), .Z(n1049) );
  NANDN U4033 ( .A(B[528]), .B(n3537), .Z(n3536) );
  NANDN U4034 ( .A(A[528]), .B(n1051), .Z(n3537) );
  NANDN U4035 ( .A(n1051), .B(A[528]), .Z(n3535) );
  AND U4036 ( .A(n3538), .B(n3539), .Z(n1051) );
  NANDN U4037 ( .A(B[527]), .B(n3540), .Z(n3539) );
  NANDN U4038 ( .A(A[527]), .B(n1053), .Z(n3540) );
  NANDN U4039 ( .A(n1053), .B(A[527]), .Z(n3538) );
  AND U4040 ( .A(n3541), .B(n3542), .Z(n1053) );
  NANDN U4041 ( .A(B[526]), .B(n3543), .Z(n3542) );
  NANDN U4042 ( .A(A[526]), .B(n1055), .Z(n3543) );
  NANDN U4043 ( .A(n1055), .B(A[526]), .Z(n3541) );
  AND U4044 ( .A(n3544), .B(n3545), .Z(n1055) );
  NANDN U4045 ( .A(B[525]), .B(n3546), .Z(n3545) );
  NANDN U4046 ( .A(A[525]), .B(n1057), .Z(n3546) );
  NANDN U4047 ( .A(n1057), .B(A[525]), .Z(n3544) );
  AND U4048 ( .A(n3547), .B(n3548), .Z(n1057) );
  NANDN U4049 ( .A(B[524]), .B(n3549), .Z(n3548) );
  NANDN U4050 ( .A(A[524]), .B(n1059), .Z(n3549) );
  NANDN U4051 ( .A(n1059), .B(A[524]), .Z(n3547) );
  AND U4052 ( .A(n3550), .B(n3551), .Z(n1059) );
  NANDN U4053 ( .A(B[523]), .B(n3552), .Z(n3551) );
  NANDN U4054 ( .A(A[523]), .B(n1061), .Z(n3552) );
  NANDN U4055 ( .A(n1061), .B(A[523]), .Z(n3550) );
  AND U4056 ( .A(n3553), .B(n3554), .Z(n1061) );
  NANDN U4057 ( .A(B[522]), .B(n3555), .Z(n3554) );
  NANDN U4058 ( .A(A[522]), .B(n1063), .Z(n3555) );
  NANDN U4059 ( .A(n1063), .B(A[522]), .Z(n3553) );
  AND U4060 ( .A(n3556), .B(n3557), .Z(n1063) );
  NANDN U4061 ( .A(B[521]), .B(n3558), .Z(n3557) );
  NANDN U4062 ( .A(A[521]), .B(n1065), .Z(n3558) );
  NANDN U4063 ( .A(n1065), .B(A[521]), .Z(n3556) );
  AND U4064 ( .A(n3559), .B(n3560), .Z(n1065) );
  NANDN U4065 ( .A(B[520]), .B(n3561), .Z(n3560) );
  NANDN U4066 ( .A(A[520]), .B(n1067), .Z(n3561) );
  NANDN U4067 ( .A(n1067), .B(A[520]), .Z(n3559) );
  AND U4068 ( .A(n3562), .B(n3563), .Z(n1067) );
  NANDN U4069 ( .A(B[519]), .B(n3564), .Z(n3563) );
  NANDN U4070 ( .A(A[519]), .B(n1071), .Z(n3564) );
  NANDN U4071 ( .A(n1071), .B(A[519]), .Z(n3562) );
  AND U4072 ( .A(n3565), .B(n3566), .Z(n1071) );
  NANDN U4073 ( .A(B[518]), .B(n3567), .Z(n3566) );
  NANDN U4074 ( .A(A[518]), .B(n1073), .Z(n3567) );
  NANDN U4075 ( .A(n1073), .B(A[518]), .Z(n3565) );
  AND U4076 ( .A(n3568), .B(n3569), .Z(n1073) );
  NANDN U4077 ( .A(B[517]), .B(n3570), .Z(n3569) );
  NANDN U4078 ( .A(A[517]), .B(n1075), .Z(n3570) );
  NANDN U4079 ( .A(n1075), .B(A[517]), .Z(n3568) );
  AND U4080 ( .A(n3571), .B(n3572), .Z(n1075) );
  NANDN U4081 ( .A(B[516]), .B(n3573), .Z(n3572) );
  NANDN U4082 ( .A(A[516]), .B(n1077), .Z(n3573) );
  NANDN U4083 ( .A(n1077), .B(A[516]), .Z(n3571) );
  AND U4084 ( .A(n3574), .B(n3575), .Z(n1077) );
  NANDN U4085 ( .A(B[515]), .B(n3576), .Z(n3575) );
  NANDN U4086 ( .A(A[515]), .B(n1079), .Z(n3576) );
  NANDN U4087 ( .A(n1079), .B(A[515]), .Z(n3574) );
  AND U4088 ( .A(n3577), .B(n3578), .Z(n1079) );
  NANDN U4089 ( .A(B[514]), .B(n3579), .Z(n3578) );
  NANDN U4090 ( .A(A[514]), .B(n1081), .Z(n3579) );
  NANDN U4091 ( .A(n1081), .B(A[514]), .Z(n3577) );
  AND U4092 ( .A(n3580), .B(n3581), .Z(n1081) );
  NANDN U4093 ( .A(B[513]), .B(n3582), .Z(n3581) );
  NANDN U4094 ( .A(A[513]), .B(n1083), .Z(n3582) );
  NANDN U4095 ( .A(n1083), .B(A[513]), .Z(n3580) );
  AND U4096 ( .A(n3583), .B(n3584), .Z(n1083) );
  NANDN U4097 ( .A(B[512]), .B(n3585), .Z(n3584) );
  NANDN U4098 ( .A(A[512]), .B(n1085), .Z(n3585) );
  NANDN U4099 ( .A(n1085), .B(A[512]), .Z(n3583) );
  AND U4100 ( .A(n3586), .B(n3587), .Z(n1085) );
  NANDN U4101 ( .A(B[511]), .B(n3588), .Z(n3587) );
  NANDN U4102 ( .A(A[511]), .B(n1087), .Z(n3588) );
  NANDN U4103 ( .A(n1087), .B(A[511]), .Z(n3586) );
  AND U4104 ( .A(n3589), .B(n3590), .Z(n1087) );
  NANDN U4105 ( .A(B[510]), .B(n3591), .Z(n3590) );
  NANDN U4106 ( .A(A[510]), .B(n1089), .Z(n3591) );
  NANDN U4107 ( .A(n1089), .B(A[510]), .Z(n3589) );
  AND U4108 ( .A(n3592), .B(n3593), .Z(n1089) );
  NANDN U4109 ( .A(B[509]), .B(n3594), .Z(n3593) );
  NANDN U4110 ( .A(A[509]), .B(n1093), .Z(n3594) );
  NANDN U4111 ( .A(n1093), .B(A[509]), .Z(n3592) );
  AND U4112 ( .A(n3595), .B(n3596), .Z(n1093) );
  NANDN U4113 ( .A(B[508]), .B(n3597), .Z(n3596) );
  NANDN U4114 ( .A(A[508]), .B(n1095), .Z(n3597) );
  NANDN U4115 ( .A(n1095), .B(A[508]), .Z(n3595) );
  AND U4116 ( .A(n3598), .B(n3599), .Z(n1095) );
  NANDN U4117 ( .A(B[507]), .B(n3600), .Z(n3599) );
  NANDN U4118 ( .A(A[507]), .B(n1097), .Z(n3600) );
  NANDN U4119 ( .A(n1097), .B(A[507]), .Z(n3598) );
  AND U4120 ( .A(n3601), .B(n3602), .Z(n1097) );
  NANDN U4121 ( .A(B[506]), .B(n3603), .Z(n3602) );
  NANDN U4122 ( .A(A[506]), .B(n1099), .Z(n3603) );
  NANDN U4123 ( .A(n1099), .B(A[506]), .Z(n3601) );
  AND U4124 ( .A(n3604), .B(n3605), .Z(n1099) );
  NANDN U4125 ( .A(B[505]), .B(n3606), .Z(n3605) );
  NANDN U4126 ( .A(A[505]), .B(n1101), .Z(n3606) );
  NANDN U4127 ( .A(n1101), .B(A[505]), .Z(n3604) );
  AND U4128 ( .A(n3607), .B(n3608), .Z(n1101) );
  NANDN U4129 ( .A(B[504]), .B(n3609), .Z(n3608) );
  NANDN U4130 ( .A(A[504]), .B(n1103), .Z(n3609) );
  NANDN U4131 ( .A(n1103), .B(A[504]), .Z(n3607) );
  AND U4132 ( .A(n3610), .B(n3611), .Z(n1103) );
  NANDN U4133 ( .A(B[503]), .B(n3612), .Z(n3611) );
  NANDN U4134 ( .A(A[503]), .B(n1105), .Z(n3612) );
  NANDN U4135 ( .A(n1105), .B(A[503]), .Z(n3610) );
  AND U4136 ( .A(n3613), .B(n3614), .Z(n1105) );
  NANDN U4137 ( .A(B[502]), .B(n3615), .Z(n3614) );
  NANDN U4138 ( .A(A[502]), .B(n1107), .Z(n3615) );
  NANDN U4139 ( .A(n1107), .B(A[502]), .Z(n3613) );
  AND U4140 ( .A(n3616), .B(n3617), .Z(n1107) );
  NANDN U4141 ( .A(B[501]), .B(n3618), .Z(n3617) );
  NANDN U4142 ( .A(A[501]), .B(n1109), .Z(n3618) );
  NANDN U4143 ( .A(n1109), .B(A[501]), .Z(n3616) );
  AND U4144 ( .A(n3619), .B(n3620), .Z(n1109) );
  NANDN U4145 ( .A(B[500]), .B(n3621), .Z(n3620) );
  NANDN U4146 ( .A(A[500]), .B(n1111), .Z(n3621) );
  NANDN U4147 ( .A(n1111), .B(A[500]), .Z(n3619) );
  AND U4148 ( .A(n3622), .B(n3623), .Z(n1111) );
  NANDN U4149 ( .A(B[499]), .B(n3624), .Z(n3623) );
  NANDN U4150 ( .A(A[499]), .B(n1117), .Z(n3624) );
  NANDN U4151 ( .A(n1117), .B(A[499]), .Z(n3622) );
  AND U4152 ( .A(n3625), .B(n3626), .Z(n1117) );
  NANDN U4153 ( .A(B[498]), .B(n3627), .Z(n3626) );
  NANDN U4154 ( .A(A[498]), .B(n1119), .Z(n3627) );
  NANDN U4155 ( .A(n1119), .B(A[498]), .Z(n3625) );
  AND U4156 ( .A(n3628), .B(n3629), .Z(n1119) );
  NANDN U4157 ( .A(B[497]), .B(n3630), .Z(n3629) );
  NANDN U4158 ( .A(A[497]), .B(n1121), .Z(n3630) );
  NANDN U4159 ( .A(n1121), .B(A[497]), .Z(n3628) );
  AND U4160 ( .A(n3631), .B(n3632), .Z(n1121) );
  NANDN U4161 ( .A(B[496]), .B(n3633), .Z(n3632) );
  NANDN U4162 ( .A(A[496]), .B(n1123), .Z(n3633) );
  NANDN U4163 ( .A(n1123), .B(A[496]), .Z(n3631) );
  AND U4164 ( .A(n3634), .B(n3635), .Z(n1123) );
  NANDN U4165 ( .A(B[495]), .B(n3636), .Z(n3635) );
  NANDN U4166 ( .A(A[495]), .B(n1125), .Z(n3636) );
  NANDN U4167 ( .A(n1125), .B(A[495]), .Z(n3634) );
  AND U4168 ( .A(n3637), .B(n3638), .Z(n1125) );
  NANDN U4169 ( .A(B[494]), .B(n3639), .Z(n3638) );
  NANDN U4170 ( .A(A[494]), .B(n1127), .Z(n3639) );
  NANDN U4171 ( .A(n1127), .B(A[494]), .Z(n3637) );
  AND U4172 ( .A(n3640), .B(n3641), .Z(n1127) );
  NANDN U4173 ( .A(B[493]), .B(n3642), .Z(n3641) );
  NANDN U4174 ( .A(A[493]), .B(n1129), .Z(n3642) );
  NANDN U4175 ( .A(n1129), .B(A[493]), .Z(n3640) );
  AND U4176 ( .A(n3643), .B(n3644), .Z(n1129) );
  NANDN U4177 ( .A(B[492]), .B(n3645), .Z(n3644) );
  NANDN U4178 ( .A(A[492]), .B(n1131), .Z(n3645) );
  NANDN U4179 ( .A(n1131), .B(A[492]), .Z(n3643) );
  AND U4180 ( .A(n3646), .B(n3647), .Z(n1131) );
  NANDN U4181 ( .A(B[491]), .B(n3648), .Z(n3647) );
  NANDN U4182 ( .A(A[491]), .B(n1133), .Z(n3648) );
  NANDN U4183 ( .A(n1133), .B(A[491]), .Z(n3646) );
  AND U4184 ( .A(n3649), .B(n3650), .Z(n1133) );
  NANDN U4185 ( .A(B[490]), .B(n3651), .Z(n3650) );
  NANDN U4186 ( .A(A[490]), .B(n1135), .Z(n3651) );
  NANDN U4187 ( .A(n1135), .B(A[490]), .Z(n3649) );
  AND U4188 ( .A(n3652), .B(n3653), .Z(n1135) );
  NANDN U4189 ( .A(B[489]), .B(n3654), .Z(n3653) );
  NANDN U4190 ( .A(A[489]), .B(n1139), .Z(n3654) );
  NANDN U4191 ( .A(n1139), .B(A[489]), .Z(n3652) );
  AND U4192 ( .A(n3655), .B(n3656), .Z(n1139) );
  NANDN U4193 ( .A(B[488]), .B(n3657), .Z(n3656) );
  NANDN U4194 ( .A(A[488]), .B(n1141), .Z(n3657) );
  NANDN U4195 ( .A(n1141), .B(A[488]), .Z(n3655) );
  AND U4196 ( .A(n3658), .B(n3659), .Z(n1141) );
  NANDN U4197 ( .A(B[487]), .B(n3660), .Z(n3659) );
  NANDN U4198 ( .A(A[487]), .B(n1143), .Z(n3660) );
  NANDN U4199 ( .A(n1143), .B(A[487]), .Z(n3658) );
  AND U4200 ( .A(n3661), .B(n3662), .Z(n1143) );
  NANDN U4201 ( .A(B[486]), .B(n3663), .Z(n3662) );
  NANDN U4202 ( .A(A[486]), .B(n1145), .Z(n3663) );
  NANDN U4203 ( .A(n1145), .B(A[486]), .Z(n3661) );
  AND U4204 ( .A(n3664), .B(n3665), .Z(n1145) );
  NANDN U4205 ( .A(B[485]), .B(n3666), .Z(n3665) );
  NANDN U4206 ( .A(A[485]), .B(n1147), .Z(n3666) );
  NANDN U4207 ( .A(n1147), .B(A[485]), .Z(n3664) );
  AND U4208 ( .A(n3667), .B(n3668), .Z(n1147) );
  NANDN U4209 ( .A(B[484]), .B(n3669), .Z(n3668) );
  NANDN U4210 ( .A(A[484]), .B(n1149), .Z(n3669) );
  NANDN U4211 ( .A(n1149), .B(A[484]), .Z(n3667) );
  AND U4212 ( .A(n3670), .B(n3671), .Z(n1149) );
  NANDN U4213 ( .A(B[483]), .B(n3672), .Z(n3671) );
  NANDN U4214 ( .A(A[483]), .B(n1151), .Z(n3672) );
  NANDN U4215 ( .A(n1151), .B(A[483]), .Z(n3670) );
  AND U4216 ( .A(n3673), .B(n3674), .Z(n1151) );
  NANDN U4217 ( .A(B[482]), .B(n3675), .Z(n3674) );
  NANDN U4218 ( .A(A[482]), .B(n1153), .Z(n3675) );
  NANDN U4219 ( .A(n1153), .B(A[482]), .Z(n3673) );
  AND U4220 ( .A(n3676), .B(n3677), .Z(n1153) );
  NANDN U4221 ( .A(B[481]), .B(n3678), .Z(n3677) );
  NANDN U4222 ( .A(A[481]), .B(n1155), .Z(n3678) );
  NANDN U4223 ( .A(n1155), .B(A[481]), .Z(n3676) );
  AND U4224 ( .A(n3679), .B(n3680), .Z(n1155) );
  NANDN U4225 ( .A(B[480]), .B(n3681), .Z(n3680) );
  NANDN U4226 ( .A(A[480]), .B(n1157), .Z(n3681) );
  NANDN U4227 ( .A(n1157), .B(A[480]), .Z(n3679) );
  AND U4228 ( .A(n3682), .B(n3683), .Z(n1157) );
  NANDN U4229 ( .A(B[479]), .B(n3684), .Z(n3683) );
  NANDN U4230 ( .A(A[479]), .B(n1161), .Z(n3684) );
  NANDN U4231 ( .A(n1161), .B(A[479]), .Z(n3682) );
  AND U4232 ( .A(n3685), .B(n3686), .Z(n1161) );
  NANDN U4233 ( .A(B[478]), .B(n3687), .Z(n3686) );
  NANDN U4234 ( .A(A[478]), .B(n1163), .Z(n3687) );
  NANDN U4235 ( .A(n1163), .B(A[478]), .Z(n3685) );
  AND U4236 ( .A(n3688), .B(n3689), .Z(n1163) );
  NANDN U4237 ( .A(B[477]), .B(n3690), .Z(n3689) );
  NANDN U4238 ( .A(A[477]), .B(n1165), .Z(n3690) );
  NANDN U4239 ( .A(n1165), .B(A[477]), .Z(n3688) );
  AND U4240 ( .A(n3691), .B(n3692), .Z(n1165) );
  NANDN U4241 ( .A(B[476]), .B(n3693), .Z(n3692) );
  NANDN U4242 ( .A(A[476]), .B(n1167), .Z(n3693) );
  NANDN U4243 ( .A(n1167), .B(A[476]), .Z(n3691) );
  AND U4244 ( .A(n3694), .B(n3695), .Z(n1167) );
  NANDN U4245 ( .A(B[475]), .B(n3696), .Z(n3695) );
  NANDN U4246 ( .A(A[475]), .B(n1169), .Z(n3696) );
  NANDN U4247 ( .A(n1169), .B(A[475]), .Z(n3694) );
  AND U4248 ( .A(n3697), .B(n3698), .Z(n1169) );
  NANDN U4249 ( .A(B[474]), .B(n3699), .Z(n3698) );
  NANDN U4250 ( .A(A[474]), .B(n1171), .Z(n3699) );
  NANDN U4251 ( .A(n1171), .B(A[474]), .Z(n3697) );
  AND U4252 ( .A(n3700), .B(n3701), .Z(n1171) );
  NANDN U4253 ( .A(B[473]), .B(n3702), .Z(n3701) );
  NANDN U4254 ( .A(A[473]), .B(n1173), .Z(n3702) );
  NANDN U4255 ( .A(n1173), .B(A[473]), .Z(n3700) );
  AND U4256 ( .A(n3703), .B(n3704), .Z(n1173) );
  NANDN U4257 ( .A(B[472]), .B(n3705), .Z(n3704) );
  NANDN U4258 ( .A(A[472]), .B(n1175), .Z(n3705) );
  NANDN U4259 ( .A(n1175), .B(A[472]), .Z(n3703) );
  AND U4260 ( .A(n3706), .B(n3707), .Z(n1175) );
  NANDN U4261 ( .A(B[471]), .B(n3708), .Z(n3707) );
  NANDN U4262 ( .A(A[471]), .B(n1177), .Z(n3708) );
  NANDN U4263 ( .A(n1177), .B(A[471]), .Z(n3706) );
  AND U4264 ( .A(n3709), .B(n3710), .Z(n1177) );
  NANDN U4265 ( .A(B[470]), .B(n3711), .Z(n3710) );
  NANDN U4266 ( .A(A[470]), .B(n1179), .Z(n3711) );
  NANDN U4267 ( .A(n1179), .B(A[470]), .Z(n3709) );
  AND U4268 ( .A(n3712), .B(n3713), .Z(n1179) );
  NANDN U4269 ( .A(B[469]), .B(n3714), .Z(n3713) );
  NANDN U4270 ( .A(A[469]), .B(n1183), .Z(n3714) );
  NANDN U4271 ( .A(n1183), .B(A[469]), .Z(n3712) );
  AND U4272 ( .A(n3715), .B(n3716), .Z(n1183) );
  NANDN U4273 ( .A(B[468]), .B(n3717), .Z(n3716) );
  NANDN U4274 ( .A(A[468]), .B(n1185), .Z(n3717) );
  NANDN U4275 ( .A(n1185), .B(A[468]), .Z(n3715) );
  AND U4276 ( .A(n3718), .B(n3719), .Z(n1185) );
  NANDN U4277 ( .A(B[467]), .B(n3720), .Z(n3719) );
  NANDN U4278 ( .A(A[467]), .B(n1187), .Z(n3720) );
  NANDN U4279 ( .A(n1187), .B(A[467]), .Z(n3718) );
  AND U4280 ( .A(n3721), .B(n3722), .Z(n1187) );
  NANDN U4281 ( .A(B[466]), .B(n3723), .Z(n3722) );
  NANDN U4282 ( .A(A[466]), .B(n1189), .Z(n3723) );
  NANDN U4283 ( .A(n1189), .B(A[466]), .Z(n3721) );
  AND U4284 ( .A(n3724), .B(n3725), .Z(n1189) );
  NANDN U4285 ( .A(B[465]), .B(n3726), .Z(n3725) );
  NANDN U4286 ( .A(A[465]), .B(n1191), .Z(n3726) );
  NANDN U4287 ( .A(n1191), .B(A[465]), .Z(n3724) );
  AND U4288 ( .A(n3727), .B(n3728), .Z(n1191) );
  NANDN U4289 ( .A(B[464]), .B(n3729), .Z(n3728) );
  NANDN U4290 ( .A(A[464]), .B(n1193), .Z(n3729) );
  NANDN U4291 ( .A(n1193), .B(A[464]), .Z(n3727) );
  AND U4292 ( .A(n3730), .B(n3731), .Z(n1193) );
  NANDN U4293 ( .A(B[463]), .B(n3732), .Z(n3731) );
  NANDN U4294 ( .A(A[463]), .B(n1195), .Z(n3732) );
  NANDN U4295 ( .A(n1195), .B(A[463]), .Z(n3730) );
  AND U4296 ( .A(n3733), .B(n3734), .Z(n1195) );
  NANDN U4297 ( .A(B[462]), .B(n3735), .Z(n3734) );
  NANDN U4298 ( .A(A[462]), .B(n1197), .Z(n3735) );
  NANDN U4299 ( .A(n1197), .B(A[462]), .Z(n3733) );
  AND U4300 ( .A(n3736), .B(n3737), .Z(n1197) );
  NANDN U4301 ( .A(B[461]), .B(n3738), .Z(n3737) );
  NANDN U4302 ( .A(A[461]), .B(n1199), .Z(n3738) );
  NANDN U4303 ( .A(n1199), .B(A[461]), .Z(n3736) );
  AND U4304 ( .A(n3739), .B(n3740), .Z(n1199) );
  NANDN U4305 ( .A(B[460]), .B(n3741), .Z(n3740) );
  NANDN U4306 ( .A(A[460]), .B(n1201), .Z(n3741) );
  NANDN U4307 ( .A(n1201), .B(A[460]), .Z(n3739) );
  AND U4308 ( .A(n3742), .B(n3743), .Z(n1201) );
  NANDN U4309 ( .A(B[459]), .B(n3744), .Z(n3743) );
  NANDN U4310 ( .A(A[459]), .B(n1205), .Z(n3744) );
  NANDN U4311 ( .A(n1205), .B(A[459]), .Z(n3742) );
  AND U4312 ( .A(n3745), .B(n3746), .Z(n1205) );
  NANDN U4313 ( .A(B[458]), .B(n3747), .Z(n3746) );
  NANDN U4314 ( .A(A[458]), .B(n1207), .Z(n3747) );
  NANDN U4315 ( .A(n1207), .B(A[458]), .Z(n3745) );
  AND U4316 ( .A(n3748), .B(n3749), .Z(n1207) );
  NANDN U4317 ( .A(B[457]), .B(n3750), .Z(n3749) );
  NANDN U4318 ( .A(A[457]), .B(n1209), .Z(n3750) );
  NANDN U4319 ( .A(n1209), .B(A[457]), .Z(n3748) );
  AND U4320 ( .A(n3751), .B(n3752), .Z(n1209) );
  NANDN U4321 ( .A(B[456]), .B(n3753), .Z(n3752) );
  NANDN U4322 ( .A(A[456]), .B(n1211), .Z(n3753) );
  NANDN U4323 ( .A(n1211), .B(A[456]), .Z(n3751) );
  AND U4324 ( .A(n3754), .B(n3755), .Z(n1211) );
  NANDN U4325 ( .A(B[455]), .B(n3756), .Z(n3755) );
  NANDN U4326 ( .A(A[455]), .B(n1213), .Z(n3756) );
  NANDN U4327 ( .A(n1213), .B(A[455]), .Z(n3754) );
  AND U4328 ( .A(n3757), .B(n3758), .Z(n1213) );
  NANDN U4329 ( .A(B[454]), .B(n3759), .Z(n3758) );
  NANDN U4330 ( .A(A[454]), .B(n1215), .Z(n3759) );
  NANDN U4331 ( .A(n1215), .B(A[454]), .Z(n3757) );
  AND U4332 ( .A(n3760), .B(n3761), .Z(n1215) );
  NANDN U4333 ( .A(B[453]), .B(n3762), .Z(n3761) );
  NANDN U4334 ( .A(A[453]), .B(n1217), .Z(n3762) );
  NANDN U4335 ( .A(n1217), .B(A[453]), .Z(n3760) );
  AND U4336 ( .A(n3763), .B(n3764), .Z(n1217) );
  NANDN U4337 ( .A(B[452]), .B(n3765), .Z(n3764) );
  NANDN U4338 ( .A(A[452]), .B(n1219), .Z(n3765) );
  NANDN U4339 ( .A(n1219), .B(A[452]), .Z(n3763) );
  AND U4340 ( .A(n3766), .B(n3767), .Z(n1219) );
  NANDN U4341 ( .A(B[451]), .B(n3768), .Z(n3767) );
  NANDN U4342 ( .A(A[451]), .B(n1221), .Z(n3768) );
  NANDN U4343 ( .A(n1221), .B(A[451]), .Z(n3766) );
  AND U4344 ( .A(n3769), .B(n3770), .Z(n1221) );
  NANDN U4345 ( .A(B[450]), .B(n3771), .Z(n3770) );
  NANDN U4346 ( .A(A[450]), .B(n1223), .Z(n3771) );
  NANDN U4347 ( .A(n1223), .B(A[450]), .Z(n3769) );
  AND U4348 ( .A(n3772), .B(n3773), .Z(n1223) );
  NANDN U4349 ( .A(B[449]), .B(n3774), .Z(n3773) );
  NANDN U4350 ( .A(A[449]), .B(n1227), .Z(n3774) );
  NANDN U4351 ( .A(n1227), .B(A[449]), .Z(n3772) );
  AND U4352 ( .A(n3775), .B(n3776), .Z(n1227) );
  NANDN U4353 ( .A(B[448]), .B(n3777), .Z(n3776) );
  NANDN U4354 ( .A(A[448]), .B(n1229), .Z(n3777) );
  NANDN U4355 ( .A(n1229), .B(A[448]), .Z(n3775) );
  AND U4356 ( .A(n3778), .B(n3779), .Z(n1229) );
  NANDN U4357 ( .A(B[447]), .B(n3780), .Z(n3779) );
  NANDN U4358 ( .A(A[447]), .B(n1231), .Z(n3780) );
  NANDN U4359 ( .A(n1231), .B(A[447]), .Z(n3778) );
  AND U4360 ( .A(n3781), .B(n3782), .Z(n1231) );
  NANDN U4361 ( .A(B[446]), .B(n3783), .Z(n3782) );
  NANDN U4362 ( .A(A[446]), .B(n1233), .Z(n3783) );
  NANDN U4363 ( .A(n1233), .B(A[446]), .Z(n3781) );
  AND U4364 ( .A(n3784), .B(n3785), .Z(n1233) );
  NANDN U4365 ( .A(B[445]), .B(n3786), .Z(n3785) );
  NANDN U4366 ( .A(A[445]), .B(n1235), .Z(n3786) );
  NANDN U4367 ( .A(n1235), .B(A[445]), .Z(n3784) );
  AND U4368 ( .A(n3787), .B(n3788), .Z(n1235) );
  NANDN U4369 ( .A(B[444]), .B(n3789), .Z(n3788) );
  NANDN U4370 ( .A(A[444]), .B(n1237), .Z(n3789) );
  NANDN U4371 ( .A(n1237), .B(A[444]), .Z(n3787) );
  AND U4372 ( .A(n3790), .B(n3791), .Z(n1237) );
  NANDN U4373 ( .A(B[443]), .B(n3792), .Z(n3791) );
  NANDN U4374 ( .A(A[443]), .B(n1239), .Z(n3792) );
  NANDN U4375 ( .A(n1239), .B(A[443]), .Z(n3790) );
  AND U4376 ( .A(n3793), .B(n3794), .Z(n1239) );
  NANDN U4377 ( .A(B[442]), .B(n3795), .Z(n3794) );
  NANDN U4378 ( .A(A[442]), .B(n1241), .Z(n3795) );
  NANDN U4379 ( .A(n1241), .B(A[442]), .Z(n3793) );
  AND U4380 ( .A(n3796), .B(n3797), .Z(n1241) );
  NANDN U4381 ( .A(B[441]), .B(n3798), .Z(n3797) );
  NANDN U4382 ( .A(A[441]), .B(n1243), .Z(n3798) );
  NANDN U4383 ( .A(n1243), .B(A[441]), .Z(n3796) );
  AND U4384 ( .A(n3799), .B(n3800), .Z(n1243) );
  NANDN U4385 ( .A(B[440]), .B(n3801), .Z(n3800) );
  NANDN U4386 ( .A(A[440]), .B(n1245), .Z(n3801) );
  NANDN U4387 ( .A(n1245), .B(A[440]), .Z(n3799) );
  AND U4388 ( .A(n3802), .B(n3803), .Z(n1245) );
  NANDN U4389 ( .A(B[439]), .B(n3804), .Z(n3803) );
  NANDN U4390 ( .A(A[439]), .B(n1249), .Z(n3804) );
  NANDN U4391 ( .A(n1249), .B(A[439]), .Z(n3802) );
  AND U4392 ( .A(n3805), .B(n3806), .Z(n1249) );
  NANDN U4393 ( .A(B[438]), .B(n3807), .Z(n3806) );
  NANDN U4394 ( .A(A[438]), .B(n1251), .Z(n3807) );
  NANDN U4395 ( .A(n1251), .B(A[438]), .Z(n3805) );
  AND U4396 ( .A(n3808), .B(n3809), .Z(n1251) );
  NANDN U4397 ( .A(B[437]), .B(n3810), .Z(n3809) );
  NANDN U4398 ( .A(A[437]), .B(n1253), .Z(n3810) );
  NANDN U4399 ( .A(n1253), .B(A[437]), .Z(n3808) );
  AND U4400 ( .A(n3811), .B(n3812), .Z(n1253) );
  NANDN U4401 ( .A(B[436]), .B(n3813), .Z(n3812) );
  NANDN U4402 ( .A(A[436]), .B(n1255), .Z(n3813) );
  NANDN U4403 ( .A(n1255), .B(A[436]), .Z(n3811) );
  AND U4404 ( .A(n3814), .B(n3815), .Z(n1255) );
  NANDN U4405 ( .A(B[435]), .B(n3816), .Z(n3815) );
  NANDN U4406 ( .A(A[435]), .B(n1257), .Z(n3816) );
  NANDN U4407 ( .A(n1257), .B(A[435]), .Z(n3814) );
  AND U4408 ( .A(n3817), .B(n3818), .Z(n1257) );
  NANDN U4409 ( .A(B[434]), .B(n3819), .Z(n3818) );
  NANDN U4410 ( .A(A[434]), .B(n1259), .Z(n3819) );
  NANDN U4411 ( .A(n1259), .B(A[434]), .Z(n3817) );
  AND U4412 ( .A(n3820), .B(n3821), .Z(n1259) );
  NANDN U4413 ( .A(B[433]), .B(n3822), .Z(n3821) );
  NANDN U4414 ( .A(A[433]), .B(n1261), .Z(n3822) );
  NANDN U4415 ( .A(n1261), .B(A[433]), .Z(n3820) );
  AND U4416 ( .A(n3823), .B(n3824), .Z(n1261) );
  NANDN U4417 ( .A(B[432]), .B(n3825), .Z(n3824) );
  NANDN U4418 ( .A(A[432]), .B(n1263), .Z(n3825) );
  NANDN U4419 ( .A(n1263), .B(A[432]), .Z(n3823) );
  AND U4420 ( .A(n3826), .B(n3827), .Z(n1263) );
  NANDN U4421 ( .A(B[431]), .B(n3828), .Z(n3827) );
  NANDN U4422 ( .A(A[431]), .B(n1265), .Z(n3828) );
  NANDN U4423 ( .A(n1265), .B(A[431]), .Z(n3826) );
  AND U4424 ( .A(n3829), .B(n3830), .Z(n1265) );
  NANDN U4425 ( .A(B[430]), .B(n3831), .Z(n3830) );
  NANDN U4426 ( .A(A[430]), .B(n1267), .Z(n3831) );
  NANDN U4427 ( .A(n1267), .B(A[430]), .Z(n3829) );
  AND U4428 ( .A(n3832), .B(n3833), .Z(n1267) );
  NANDN U4429 ( .A(B[429]), .B(n3834), .Z(n3833) );
  NANDN U4430 ( .A(A[429]), .B(n1271), .Z(n3834) );
  NANDN U4431 ( .A(n1271), .B(A[429]), .Z(n3832) );
  AND U4432 ( .A(n3835), .B(n3836), .Z(n1271) );
  NANDN U4433 ( .A(B[428]), .B(n3837), .Z(n3836) );
  NANDN U4434 ( .A(A[428]), .B(n1273), .Z(n3837) );
  NANDN U4435 ( .A(n1273), .B(A[428]), .Z(n3835) );
  AND U4436 ( .A(n3838), .B(n3839), .Z(n1273) );
  NANDN U4437 ( .A(B[427]), .B(n3840), .Z(n3839) );
  NANDN U4438 ( .A(A[427]), .B(n1275), .Z(n3840) );
  NANDN U4439 ( .A(n1275), .B(A[427]), .Z(n3838) );
  AND U4440 ( .A(n3841), .B(n3842), .Z(n1275) );
  NANDN U4441 ( .A(B[426]), .B(n3843), .Z(n3842) );
  NANDN U4442 ( .A(A[426]), .B(n1277), .Z(n3843) );
  NANDN U4443 ( .A(n1277), .B(A[426]), .Z(n3841) );
  AND U4444 ( .A(n3844), .B(n3845), .Z(n1277) );
  NANDN U4445 ( .A(B[425]), .B(n3846), .Z(n3845) );
  NANDN U4446 ( .A(A[425]), .B(n1279), .Z(n3846) );
  NANDN U4447 ( .A(n1279), .B(A[425]), .Z(n3844) );
  AND U4448 ( .A(n3847), .B(n3848), .Z(n1279) );
  NANDN U4449 ( .A(B[424]), .B(n3849), .Z(n3848) );
  NANDN U4450 ( .A(A[424]), .B(n1281), .Z(n3849) );
  NANDN U4451 ( .A(n1281), .B(A[424]), .Z(n3847) );
  AND U4452 ( .A(n3850), .B(n3851), .Z(n1281) );
  NANDN U4453 ( .A(B[423]), .B(n3852), .Z(n3851) );
  NANDN U4454 ( .A(A[423]), .B(n1283), .Z(n3852) );
  NANDN U4455 ( .A(n1283), .B(A[423]), .Z(n3850) );
  AND U4456 ( .A(n3853), .B(n3854), .Z(n1283) );
  NANDN U4457 ( .A(B[422]), .B(n3855), .Z(n3854) );
  NANDN U4458 ( .A(A[422]), .B(n1285), .Z(n3855) );
  NANDN U4459 ( .A(n1285), .B(A[422]), .Z(n3853) );
  AND U4460 ( .A(n3856), .B(n3857), .Z(n1285) );
  NANDN U4461 ( .A(B[421]), .B(n3858), .Z(n3857) );
  NANDN U4462 ( .A(A[421]), .B(n1287), .Z(n3858) );
  NANDN U4463 ( .A(n1287), .B(A[421]), .Z(n3856) );
  AND U4464 ( .A(n3859), .B(n3860), .Z(n1287) );
  NANDN U4465 ( .A(B[420]), .B(n3861), .Z(n3860) );
  NANDN U4466 ( .A(A[420]), .B(n1289), .Z(n3861) );
  NANDN U4467 ( .A(n1289), .B(A[420]), .Z(n3859) );
  AND U4468 ( .A(n3862), .B(n3863), .Z(n1289) );
  NANDN U4469 ( .A(B[419]), .B(n3864), .Z(n3863) );
  NANDN U4470 ( .A(A[419]), .B(n1293), .Z(n3864) );
  NANDN U4471 ( .A(n1293), .B(A[419]), .Z(n3862) );
  AND U4472 ( .A(n3865), .B(n3866), .Z(n1293) );
  NANDN U4473 ( .A(B[418]), .B(n3867), .Z(n3866) );
  NANDN U4474 ( .A(A[418]), .B(n1295), .Z(n3867) );
  NANDN U4475 ( .A(n1295), .B(A[418]), .Z(n3865) );
  AND U4476 ( .A(n3868), .B(n3869), .Z(n1295) );
  NANDN U4477 ( .A(B[417]), .B(n3870), .Z(n3869) );
  NANDN U4478 ( .A(A[417]), .B(n1297), .Z(n3870) );
  NANDN U4479 ( .A(n1297), .B(A[417]), .Z(n3868) );
  AND U4480 ( .A(n3871), .B(n3872), .Z(n1297) );
  NANDN U4481 ( .A(B[416]), .B(n3873), .Z(n3872) );
  NANDN U4482 ( .A(A[416]), .B(n1299), .Z(n3873) );
  NANDN U4483 ( .A(n1299), .B(A[416]), .Z(n3871) );
  AND U4484 ( .A(n3874), .B(n3875), .Z(n1299) );
  NANDN U4485 ( .A(B[415]), .B(n3876), .Z(n3875) );
  NANDN U4486 ( .A(A[415]), .B(n1301), .Z(n3876) );
  NANDN U4487 ( .A(n1301), .B(A[415]), .Z(n3874) );
  AND U4488 ( .A(n3877), .B(n3878), .Z(n1301) );
  NANDN U4489 ( .A(B[414]), .B(n3879), .Z(n3878) );
  NANDN U4490 ( .A(A[414]), .B(n1303), .Z(n3879) );
  NANDN U4491 ( .A(n1303), .B(A[414]), .Z(n3877) );
  AND U4492 ( .A(n3880), .B(n3881), .Z(n1303) );
  NANDN U4493 ( .A(B[413]), .B(n3882), .Z(n3881) );
  NANDN U4494 ( .A(A[413]), .B(n1305), .Z(n3882) );
  NANDN U4495 ( .A(n1305), .B(A[413]), .Z(n3880) );
  AND U4496 ( .A(n3883), .B(n3884), .Z(n1305) );
  NANDN U4497 ( .A(B[412]), .B(n3885), .Z(n3884) );
  NANDN U4498 ( .A(A[412]), .B(n1307), .Z(n3885) );
  NANDN U4499 ( .A(n1307), .B(A[412]), .Z(n3883) );
  AND U4500 ( .A(n3886), .B(n3887), .Z(n1307) );
  NANDN U4501 ( .A(B[411]), .B(n3888), .Z(n3887) );
  NANDN U4502 ( .A(A[411]), .B(n1309), .Z(n3888) );
  NANDN U4503 ( .A(n1309), .B(A[411]), .Z(n3886) );
  AND U4504 ( .A(n3889), .B(n3890), .Z(n1309) );
  NANDN U4505 ( .A(B[410]), .B(n3891), .Z(n3890) );
  NANDN U4506 ( .A(A[410]), .B(n1311), .Z(n3891) );
  NANDN U4507 ( .A(n1311), .B(A[410]), .Z(n3889) );
  AND U4508 ( .A(n3892), .B(n3893), .Z(n1311) );
  NANDN U4509 ( .A(B[409]), .B(n3894), .Z(n3893) );
  NANDN U4510 ( .A(A[409]), .B(n1315), .Z(n3894) );
  NANDN U4511 ( .A(n1315), .B(A[409]), .Z(n3892) );
  AND U4512 ( .A(n3895), .B(n3896), .Z(n1315) );
  NANDN U4513 ( .A(B[408]), .B(n3897), .Z(n3896) );
  NANDN U4514 ( .A(A[408]), .B(n1317), .Z(n3897) );
  NANDN U4515 ( .A(n1317), .B(A[408]), .Z(n3895) );
  AND U4516 ( .A(n3898), .B(n3899), .Z(n1317) );
  NANDN U4517 ( .A(B[407]), .B(n3900), .Z(n3899) );
  NANDN U4518 ( .A(A[407]), .B(n1319), .Z(n3900) );
  NANDN U4519 ( .A(n1319), .B(A[407]), .Z(n3898) );
  AND U4520 ( .A(n3901), .B(n3902), .Z(n1319) );
  NANDN U4521 ( .A(B[406]), .B(n3903), .Z(n3902) );
  NANDN U4522 ( .A(A[406]), .B(n1321), .Z(n3903) );
  NANDN U4523 ( .A(n1321), .B(A[406]), .Z(n3901) );
  AND U4524 ( .A(n3904), .B(n3905), .Z(n1321) );
  NANDN U4525 ( .A(B[405]), .B(n3906), .Z(n3905) );
  NANDN U4526 ( .A(A[405]), .B(n1323), .Z(n3906) );
  NANDN U4527 ( .A(n1323), .B(A[405]), .Z(n3904) );
  AND U4528 ( .A(n3907), .B(n3908), .Z(n1323) );
  NANDN U4529 ( .A(B[404]), .B(n3909), .Z(n3908) );
  NANDN U4530 ( .A(A[404]), .B(n1325), .Z(n3909) );
  NANDN U4531 ( .A(n1325), .B(A[404]), .Z(n3907) );
  AND U4532 ( .A(n3910), .B(n3911), .Z(n1325) );
  NANDN U4533 ( .A(B[403]), .B(n3912), .Z(n3911) );
  NANDN U4534 ( .A(A[403]), .B(n1327), .Z(n3912) );
  NANDN U4535 ( .A(n1327), .B(A[403]), .Z(n3910) );
  AND U4536 ( .A(n3913), .B(n3914), .Z(n1327) );
  NANDN U4537 ( .A(B[402]), .B(n3915), .Z(n3914) );
  NANDN U4538 ( .A(A[402]), .B(n1329), .Z(n3915) );
  NANDN U4539 ( .A(n1329), .B(A[402]), .Z(n3913) );
  AND U4540 ( .A(n3916), .B(n3917), .Z(n1329) );
  NANDN U4541 ( .A(B[401]), .B(n3918), .Z(n3917) );
  NANDN U4542 ( .A(A[401]), .B(n1331), .Z(n3918) );
  NANDN U4543 ( .A(n1331), .B(A[401]), .Z(n3916) );
  AND U4544 ( .A(n3919), .B(n3920), .Z(n1331) );
  NANDN U4545 ( .A(B[400]), .B(n3921), .Z(n3920) );
  NANDN U4546 ( .A(A[400]), .B(n1333), .Z(n3921) );
  NANDN U4547 ( .A(n1333), .B(A[400]), .Z(n3919) );
  AND U4548 ( .A(n3922), .B(n3923), .Z(n1333) );
  NANDN U4549 ( .A(B[399]), .B(n3924), .Z(n3923) );
  NANDN U4550 ( .A(A[399]), .B(n1339), .Z(n3924) );
  NANDN U4551 ( .A(n1339), .B(A[399]), .Z(n3922) );
  AND U4552 ( .A(n3925), .B(n3926), .Z(n1339) );
  NANDN U4553 ( .A(B[398]), .B(n3927), .Z(n3926) );
  NANDN U4554 ( .A(A[398]), .B(n1341), .Z(n3927) );
  NANDN U4555 ( .A(n1341), .B(A[398]), .Z(n3925) );
  AND U4556 ( .A(n3928), .B(n3929), .Z(n1341) );
  NANDN U4557 ( .A(B[397]), .B(n3930), .Z(n3929) );
  NANDN U4558 ( .A(A[397]), .B(n1343), .Z(n3930) );
  NANDN U4559 ( .A(n1343), .B(A[397]), .Z(n3928) );
  AND U4560 ( .A(n3931), .B(n3932), .Z(n1343) );
  NANDN U4561 ( .A(B[396]), .B(n3933), .Z(n3932) );
  NANDN U4562 ( .A(A[396]), .B(n1345), .Z(n3933) );
  NANDN U4563 ( .A(n1345), .B(A[396]), .Z(n3931) );
  AND U4564 ( .A(n3934), .B(n3935), .Z(n1345) );
  NANDN U4565 ( .A(B[395]), .B(n3936), .Z(n3935) );
  NANDN U4566 ( .A(A[395]), .B(n1347), .Z(n3936) );
  NANDN U4567 ( .A(n1347), .B(A[395]), .Z(n3934) );
  AND U4568 ( .A(n3937), .B(n3938), .Z(n1347) );
  NANDN U4569 ( .A(B[394]), .B(n3939), .Z(n3938) );
  NANDN U4570 ( .A(A[394]), .B(n1349), .Z(n3939) );
  NANDN U4571 ( .A(n1349), .B(A[394]), .Z(n3937) );
  AND U4572 ( .A(n3940), .B(n3941), .Z(n1349) );
  NANDN U4573 ( .A(B[393]), .B(n3942), .Z(n3941) );
  NANDN U4574 ( .A(A[393]), .B(n1351), .Z(n3942) );
  NANDN U4575 ( .A(n1351), .B(A[393]), .Z(n3940) );
  AND U4576 ( .A(n3943), .B(n3944), .Z(n1351) );
  NANDN U4577 ( .A(B[392]), .B(n3945), .Z(n3944) );
  NANDN U4578 ( .A(A[392]), .B(n1353), .Z(n3945) );
  NANDN U4579 ( .A(n1353), .B(A[392]), .Z(n3943) );
  AND U4580 ( .A(n3946), .B(n3947), .Z(n1353) );
  NANDN U4581 ( .A(B[391]), .B(n3948), .Z(n3947) );
  NANDN U4582 ( .A(A[391]), .B(n1355), .Z(n3948) );
  NANDN U4583 ( .A(n1355), .B(A[391]), .Z(n3946) );
  AND U4584 ( .A(n3949), .B(n3950), .Z(n1355) );
  NANDN U4585 ( .A(B[390]), .B(n3951), .Z(n3950) );
  NANDN U4586 ( .A(A[390]), .B(n1357), .Z(n3951) );
  NANDN U4587 ( .A(n1357), .B(A[390]), .Z(n3949) );
  AND U4588 ( .A(n3952), .B(n3953), .Z(n1357) );
  NANDN U4589 ( .A(B[389]), .B(n3954), .Z(n3953) );
  NANDN U4590 ( .A(A[389]), .B(n1361), .Z(n3954) );
  NANDN U4591 ( .A(n1361), .B(A[389]), .Z(n3952) );
  AND U4592 ( .A(n3955), .B(n3956), .Z(n1361) );
  NANDN U4593 ( .A(B[388]), .B(n3957), .Z(n3956) );
  NANDN U4594 ( .A(A[388]), .B(n1363), .Z(n3957) );
  NANDN U4595 ( .A(n1363), .B(A[388]), .Z(n3955) );
  AND U4596 ( .A(n3958), .B(n3959), .Z(n1363) );
  NANDN U4597 ( .A(B[387]), .B(n3960), .Z(n3959) );
  NANDN U4598 ( .A(A[387]), .B(n1365), .Z(n3960) );
  NANDN U4599 ( .A(n1365), .B(A[387]), .Z(n3958) );
  AND U4600 ( .A(n3961), .B(n3962), .Z(n1365) );
  NANDN U4601 ( .A(B[386]), .B(n3963), .Z(n3962) );
  NANDN U4602 ( .A(A[386]), .B(n1367), .Z(n3963) );
  NANDN U4603 ( .A(n1367), .B(A[386]), .Z(n3961) );
  AND U4604 ( .A(n3964), .B(n3965), .Z(n1367) );
  NANDN U4605 ( .A(B[385]), .B(n3966), .Z(n3965) );
  NANDN U4606 ( .A(A[385]), .B(n1369), .Z(n3966) );
  NANDN U4607 ( .A(n1369), .B(A[385]), .Z(n3964) );
  AND U4608 ( .A(n3967), .B(n3968), .Z(n1369) );
  NANDN U4609 ( .A(B[384]), .B(n3969), .Z(n3968) );
  NANDN U4610 ( .A(A[384]), .B(n1371), .Z(n3969) );
  NANDN U4611 ( .A(n1371), .B(A[384]), .Z(n3967) );
  AND U4612 ( .A(n3970), .B(n3971), .Z(n1371) );
  NANDN U4613 ( .A(B[383]), .B(n3972), .Z(n3971) );
  NANDN U4614 ( .A(A[383]), .B(n1373), .Z(n3972) );
  NANDN U4615 ( .A(n1373), .B(A[383]), .Z(n3970) );
  AND U4616 ( .A(n3973), .B(n3974), .Z(n1373) );
  NANDN U4617 ( .A(B[382]), .B(n3975), .Z(n3974) );
  NANDN U4618 ( .A(A[382]), .B(n1375), .Z(n3975) );
  NANDN U4619 ( .A(n1375), .B(A[382]), .Z(n3973) );
  AND U4620 ( .A(n3976), .B(n3977), .Z(n1375) );
  NANDN U4621 ( .A(B[381]), .B(n3978), .Z(n3977) );
  NANDN U4622 ( .A(A[381]), .B(n1377), .Z(n3978) );
  NANDN U4623 ( .A(n1377), .B(A[381]), .Z(n3976) );
  AND U4624 ( .A(n3979), .B(n3980), .Z(n1377) );
  NANDN U4625 ( .A(B[380]), .B(n3981), .Z(n3980) );
  NANDN U4626 ( .A(A[380]), .B(n1379), .Z(n3981) );
  NANDN U4627 ( .A(n1379), .B(A[380]), .Z(n3979) );
  AND U4628 ( .A(n3982), .B(n3983), .Z(n1379) );
  NANDN U4629 ( .A(B[379]), .B(n3984), .Z(n3983) );
  NANDN U4630 ( .A(A[379]), .B(n1383), .Z(n3984) );
  NANDN U4631 ( .A(n1383), .B(A[379]), .Z(n3982) );
  AND U4632 ( .A(n3985), .B(n3986), .Z(n1383) );
  NANDN U4633 ( .A(B[378]), .B(n3987), .Z(n3986) );
  NANDN U4634 ( .A(A[378]), .B(n1385), .Z(n3987) );
  NANDN U4635 ( .A(n1385), .B(A[378]), .Z(n3985) );
  AND U4636 ( .A(n3988), .B(n3989), .Z(n1385) );
  NANDN U4637 ( .A(B[377]), .B(n3990), .Z(n3989) );
  NANDN U4638 ( .A(A[377]), .B(n1387), .Z(n3990) );
  NANDN U4639 ( .A(n1387), .B(A[377]), .Z(n3988) );
  AND U4640 ( .A(n3991), .B(n3992), .Z(n1387) );
  NANDN U4641 ( .A(B[376]), .B(n3993), .Z(n3992) );
  NANDN U4642 ( .A(A[376]), .B(n1389), .Z(n3993) );
  NANDN U4643 ( .A(n1389), .B(A[376]), .Z(n3991) );
  AND U4644 ( .A(n3994), .B(n3995), .Z(n1389) );
  NANDN U4645 ( .A(B[375]), .B(n3996), .Z(n3995) );
  NANDN U4646 ( .A(A[375]), .B(n1391), .Z(n3996) );
  NANDN U4647 ( .A(n1391), .B(A[375]), .Z(n3994) );
  AND U4648 ( .A(n3997), .B(n3998), .Z(n1391) );
  NANDN U4649 ( .A(B[374]), .B(n3999), .Z(n3998) );
  NANDN U4650 ( .A(A[374]), .B(n1393), .Z(n3999) );
  NANDN U4651 ( .A(n1393), .B(A[374]), .Z(n3997) );
  AND U4652 ( .A(n4000), .B(n4001), .Z(n1393) );
  NANDN U4653 ( .A(B[373]), .B(n4002), .Z(n4001) );
  NANDN U4654 ( .A(A[373]), .B(n1395), .Z(n4002) );
  NANDN U4655 ( .A(n1395), .B(A[373]), .Z(n4000) );
  AND U4656 ( .A(n4003), .B(n4004), .Z(n1395) );
  NANDN U4657 ( .A(B[372]), .B(n4005), .Z(n4004) );
  NANDN U4658 ( .A(A[372]), .B(n1397), .Z(n4005) );
  NANDN U4659 ( .A(n1397), .B(A[372]), .Z(n4003) );
  AND U4660 ( .A(n4006), .B(n4007), .Z(n1397) );
  NANDN U4661 ( .A(B[371]), .B(n4008), .Z(n4007) );
  NANDN U4662 ( .A(A[371]), .B(n1399), .Z(n4008) );
  NANDN U4663 ( .A(n1399), .B(A[371]), .Z(n4006) );
  AND U4664 ( .A(n4009), .B(n4010), .Z(n1399) );
  NANDN U4665 ( .A(B[370]), .B(n4011), .Z(n4010) );
  NANDN U4666 ( .A(A[370]), .B(n1401), .Z(n4011) );
  NANDN U4667 ( .A(n1401), .B(A[370]), .Z(n4009) );
  AND U4668 ( .A(n4012), .B(n4013), .Z(n1401) );
  NANDN U4669 ( .A(B[369]), .B(n4014), .Z(n4013) );
  NANDN U4670 ( .A(A[369]), .B(n1405), .Z(n4014) );
  NANDN U4671 ( .A(n1405), .B(A[369]), .Z(n4012) );
  AND U4672 ( .A(n4015), .B(n4016), .Z(n1405) );
  NANDN U4673 ( .A(B[368]), .B(n4017), .Z(n4016) );
  NANDN U4674 ( .A(A[368]), .B(n1407), .Z(n4017) );
  NANDN U4675 ( .A(n1407), .B(A[368]), .Z(n4015) );
  AND U4676 ( .A(n4018), .B(n4019), .Z(n1407) );
  NANDN U4677 ( .A(B[367]), .B(n4020), .Z(n4019) );
  NANDN U4678 ( .A(A[367]), .B(n1409), .Z(n4020) );
  NANDN U4679 ( .A(n1409), .B(A[367]), .Z(n4018) );
  AND U4680 ( .A(n4021), .B(n4022), .Z(n1409) );
  NANDN U4681 ( .A(B[366]), .B(n4023), .Z(n4022) );
  NANDN U4682 ( .A(A[366]), .B(n1411), .Z(n4023) );
  NANDN U4683 ( .A(n1411), .B(A[366]), .Z(n4021) );
  AND U4684 ( .A(n4024), .B(n4025), .Z(n1411) );
  NANDN U4685 ( .A(B[365]), .B(n4026), .Z(n4025) );
  NANDN U4686 ( .A(A[365]), .B(n1413), .Z(n4026) );
  NANDN U4687 ( .A(n1413), .B(A[365]), .Z(n4024) );
  AND U4688 ( .A(n4027), .B(n4028), .Z(n1413) );
  NANDN U4689 ( .A(B[364]), .B(n4029), .Z(n4028) );
  NANDN U4690 ( .A(A[364]), .B(n1415), .Z(n4029) );
  NANDN U4691 ( .A(n1415), .B(A[364]), .Z(n4027) );
  AND U4692 ( .A(n4030), .B(n4031), .Z(n1415) );
  NANDN U4693 ( .A(B[363]), .B(n4032), .Z(n4031) );
  NANDN U4694 ( .A(A[363]), .B(n1417), .Z(n4032) );
  NANDN U4695 ( .A(n1417), .B(A[363]), .Z(n4030) );
  AND U4696 ( .A(n4033), .B(n4034), .Z(n1417) );
  NANDN U4697 ( .A(B[362]), .B(n4035), .Z(n4034) );
  NANDN U4698 ( .A(A[362]), .B(n1419), .Z(n4035) );
  NANDN U4699 ( .A(n1419), .B(A[362]), .Z(n4033) );
  AND U4700 ( .A(n4036), .B(n4037), .Z(n1419) );
  NANDN U4701 ( .A(B[361]), .B(n4038), .Z(n4037) );
  NANDN U4702 ( .A(A[361]), .B(n1421), .Z(n4038) );
  NANDN U4703 ( .A(n1421), .B(A[361]), .Z(n4036) );
  AND U4704 ( .A(n4039), .B(n4040), .Z(n1421) );
  NANDN U4705 ( .A(B[360]), .B(n4041), .Z(n4040) );
  NANDN U4706 ( .A(A[360]), .B(n1423), .Z(n4041) );
  NANDN U4707 ( .A(n1423), .B(A[360]), .Z(n4039) );
  AND U4708 ( .A(n4042), .B(n4043), .Z(n1423) );
  NANDN U4709 ( .A(B[359]), .B(n4044), .Z(n4043) );
  NANDN U4710 ( .A(A[359]), .B(n1427), .Z(n4044) );
  NANDN U4711 ( .A(n1427), .B(A[359]), .Z(n4042) );
  AND U4712 ( .A(n4045), .B(n4046), .Z(n1427) );
  NANDN U4713 ( .A(B[358]), .B(n4047), .Z(n4046) );
  NANDN U4714 ( .A(A[358]), .B(n1429), .Z(n4047) );
  NANDN U4715 ( .A(n1429), .B(A[358]), .Z(n4045) );
  AND U4716 ( .A(n4048), .B(n4049), .Z(n1429) );
  NANDN U4717 ( .A(B[357]), .B(n4050), .Z(n4049) );
  NANDN U4718 ( .A(A[357]), .B(n1431), .Z(n4050) );
  NANDN U4719 ( .A(n1431), .B(A[357]), .Z(n4048) );
  AND U4720 ( .A(n4051), .B(n4052), .Z(n1431) );
  NANDN U4721 ( .A(B[356]), .B(n4053), .Z(n4052) );
  NANDN U4722 ( .A(A[356]), .B(n1433), .Z(n4053) );
  NANDN U4723 ( .A(n1433), .B(A[356]), .Z(n4051) );
  AND U4724 ( .A(n4054), .B(n4055), .Z(n1433) );
  NANDN U4725 ( .A(B[355]), .B(n4056), .Z(n4055) );
  NANDN U4726 ( .A(A[355]), .B(n1435), .Z(n4056) );
  NANDN U4727 ( .A(n1435), .B(A[355]), .Z(n4054) );
  AND U4728 ( .A(n4057), .B(n4058), .Z(n1435) );
  NANDN U4729 ( .A(B[354]), .B(n4059), .Z(n4058) );
  NANDN U4730 ( .A(A[354]), .B(n1437), .Z(n4059) );
  NANDN U4731 ( .A(n1437), .B(A[354]), .Z(n4057) );
  AND U4732 ( .A(n4060), .B(n4061), .Z(n1437) );
  NANDN U4733 ( .A(B[353]), .B(n4062), .Z(n4061) );
  NANDN U4734 ( .A(A[353]), .B(n1439), .Z(n4062) );
  NANDN U4735 ( .A(n1439), .B(A[353]), .Z(n4060) );
  AND U4736 ( .A(n4063), .B(n4064), .Z(n1439) );
  NANDN U4737 ( .A(B[352]), .B(n4065), .Z(n4064) );
  NANDN U4738 ( .A(A[352]), .B(n1441), .Z(n4065) );
  NANDN U4739 ( .A(n1441), .B(A[352]), .Z(n4063) );
  AND U4740 ( .A(n4066), .B(n4067), .Z(n1441) );
  NANDN U4741 ( .A(B[351]), .B(n4068), .Z(n4067) );
  NANDN U4742 ( .A(A[351]), .B(n1443), .Z(n4068) );
  NANDN U4743 ( .A(n1443), .B(A[351]), .Z(n4066) );
  AND U4744 ( .A(n4069), .B(n4070), .Z(n1443) );
  NANDN U4745 ( .A(B[350]), .B(n4071), .Z(n4070) );
  NANDN U4746 ( .A(A[350]), .B(n1445), .Z(n4071) );
  NANDN U4747 ( .A(n1445), .B(A[350]), .Z(n4069) );
  AND U4748 ( .A(n4072), .B(n4073), .Z(n1445) );
  NANDN U4749 ( .A(B[349]), .B(n4074), .Z(n4073) );
  NANDN U4750 ( .A(A[349]), .B(n1449), .Z(n4074) );
  NANDN U4751 ( .A(n1449), .B(A[349]), .Z(n4072) );
  AND U4752 ( .A(n4075), .B(n4076), .Z(n1449) );
  NANDN U4753 ( .A(B[348]), .B(n4077), .Z(n4076) );
  NANDN U4754 ( .A(A[348]), .B(n1451), .Z(n4077) );
  NANDN U4755 ( .A(n1451), .B(A[348]), .Z(n4075) );
  AND U4756 ( .A(n4078), .B(n4079), .Z(n1451) );
  NANDN U4757 ( .A(B[347]), .B(n4080), .Z(n4079) );
  NANDN U4758 ( .A(A[347]), .B(n1453), .Z(n4080) );
  NANDN U4759 ( .A(n1453), .B(A[347]), .Z(n4078) );
  AND U4760 ( .A(n4081), .B(n4082), .Z(n1453) );
  NANDN U4761 ( .A(B[346]), .B(n4083), .Z(n4082) );
  NANDN U4762 ( .A(A[346]), .B(n1455), .Z(n4083) );
  NANDN U4763 ( .A(n1455), .B(A[346]), .Z(n4081) );
  AND U4764 ( .A(n4084), .B(n4085), .Z(n1455) );
  NANDN U4765 ( .A(B[345]), .B(n4086), .Z(n4085) );
  NANDN U4766 ( .A(A[345]), .B(n1457), .Z(n4086) );
  NANDN U4767 ( .A(n1457), .B(A[345]), .Z(n4084) );
  AND U4768 ( .A(n4087), .B(n4088), .Z(n1457) );
  NANDN U4769 ( .A(B[344]), .B(n4089), .Z(n4088) );
  NANDN U4770 ( .A(A[344]), .B(n1459), .Z(n4089) );
  NANDN U4771 ( .A(n1459), .B(A[344]), .Z(n4087) );
  AND U4772 ( .A(n4090), .B(n4091), .Z(n1459) );
  NANDN U4773 ( .A(B[343]), .B(n4092), .Z(n4091) );
  NANDN U4774 ( .A(A[343]), .B(n1461), .Z(n4092) );
  NANDN U4775 ( .A(n1461), .B(A[343]), .Z(n4090) );
  AND U4776 ( .A(n4093), .B(n4094), .Z(n1461) );
  NANDN U4777 ( .A(B[342]), .B(n4095), .Z(n4094) );
  NANDN U4778 ( .A(A[342]), .B(n1463), .Z(n4095) );
  NANDN U4779 ( .A(n1463), .B(A[342]), .Z(n4093) );
  AND U4780 ( .A(n4096), .B(n4097), .Z(n1463) );
  NANDN U4781 ( .A(B[341]), .B(n4098), .Z(n4097) );
  NANDN U4782 ( .A(A[341]), .B(n1465), .Z(n4098) );
  NANDN U4783 ( .A(n1465), .B(A[341]), .Z(n4096) );
  AND U4784 ( .A(n4099), .B(n4100), .Z(n1465) );
  NANDN U4785 ( .A(B[340]), .B(n4101), .Z(n4100) );
  NANDN U4786 ( .A(A[340]), .B(n1467), .Z(n4101) );
  NANDN U4787 ( .A(n1467), .B(A[340]), .Z(n4099) );
  AND U4788 ( .A(n4102), .B(n4103), .Z(n1467) );
  NANDN U4789 ( .A(B[339]), .B(n4104), .Z(n4103) );
  NANDN U4790 ( .A(A[339]), .B(n1471), .Z(n4104) );
  NANDN U4791 ( .A(n1471), .B(A[339]), .Z(n4102) );
  AND U4792 ( .A(n4105), .B(n4106), .Z(n1471) );
  NANDN U4793 ( .A(B[338]), .B(n4107), .Z(n4106) );
  NANDN U4794 ( .A(A[338]), .B(n1473), .Z(n4107) );
  NANDN U4795 ( .A(n1473), .B(A[338]), .Z(n4105) );
  AND U4796 ( .A(n4108), .B(n4109), .Z(n1473) );
  NANDN U4797 ( .A(B[337]), .B(n4110), .Z(n4109) );
  NANDN U4798 ( .A(A[337]), .B(n1475), .Z(n4110) );
  NANDN U4799 ( .A(n1475), .B(A[337]), .Z(n4108) );
  AND U4800 ( .A(n4111), .B(n4112), .Z(n1475) );
  NANDN U4801 ( .A(B[336]), .B(n4113), .Z(n4112) );
  NANDN U4802 ( .A(A[336]), .B(n1477), .Z(n4113) );
  NANDN U4803 ( .A(n1477), .B(A[336]), .Z(n4111) );
  AND U4804 ( .A(n4114), .B(n4115), .Z(n1477) );
  NANDN U4805 ( .A(B[335]), .B(n4116), .Z(n4115) );
  NANDN U4806 ( .A(A[335]), .B(n1479), .Z(n4116) );
  NANDN U4807 ( .A(n1479), .B(A[335]), .Z(n4114) );
  AND U4808 ( .A(n4117), .B(n4118), .Z(n1479) );
  NANDN U4809 ( .A(B[334]), .B(n4119), .Z(n4118) );
  NANDN U4810 ( .A(A[334]), .B(n1481), .Z(n4119) );
  NANDN U4811 ( .A(n1481), .B(A[334]), .Z(n4117) );
  AND U4812 ( .A(n4120), .B(n4121), .Z(n1481) );
  NANDN U4813 ( .A(B[333]), .B(n4122), .Z(n4121) );
  NANDN U4814 ( .A(A[333]), .B(n1483), .Z(n4122) );
  NANDN U4815 ( .A(n1483), .B(A[333]), .Z(n4120) );
  AND U4816 ( .A(n4123), .B(n4124), .Z(n1483) );
  NANDN U4817 ( .A(B[332]), .B(n4125), .Z(n4124) );
  NANDN U4818 ( .A(A[332]), .B(n1485), .Z(n4125) );
  NANDN U4819 ( .A(n1485), .B(A[332]), .Z(n4123) );
  AND U4820 ( .A(n4126), .B(n4127), .Z(n1485) );
  NANDN U4821 ( .A(B[331]), .B(n4128), .Z(n4127) );
  NANDN U4822 ( .A(A[331]), .B(n1487), .Z(n4128) );
  NANDN U4823 ( .A(n1487), .B(A[331]), .Z(n4126) );
  AND U4824 ( .A(n4129), .B(n4130), .Z(n1487) );
  NANDN U4825 ( .A(B[330]), .B(n4131), .Z(n4130) );
  NANDN U4826 ( .A(A[330]), .B(n1489), .Z(n4131) );
  NANDN U4827 ( .A(n1489), .B(A[330]), .Z(n4129) );
  AND U4828 ( .A(n4132), .B(n4133), .Z(n1489) );
  NANDN U4829 ( .A(B[329]), .B(n4134), .Z(n4133) );
  NANDN U4830 ( .A(A[329]), .B(n1493), .Z(n4134) );
  NANDN U4831 ( .A(n1493), .B(A[329]), .Z(n4132) );
  AND U4832 ( .A(n4135), .B(n4136), .Z(n1493) );
  NANDN U4833 ( .A(B[328]), .B(n4137), .Z(n4136) );
  NANDN U4834 ( .A(A[328]), .B(n1495), .Z(n4137) );
  NANDN U4835 ( .A(n1495), .B(A[328]), .Z(n4135) );
  AND U4836 ( .A(n4138), .B(n4139), .Z(n1495) );
  NANDN U4837 ( .A(B[327]), .B(n4140), .Z(n4139) );
  NANDN U4838 ( .A(A[327]), .B(n1497), .Z(n4140) );
  NANDN U4839 ( .A(n1497), .B(A[327]), .Z(n4138) );
  AND U4840 ( .A(n4141), .B(n4142), .Z(n1497) );
  NANDN U4841 ( .A(B[326]), .B(n4143), .Z(n4142) );
  NANDN U4842 ( .A(A[326]), .B(n1499), .Z(n4143) );
  NANDN U4843 ( .A(n1499), .B(A[326]), .Z(n4141) );
  AND U4844 ( .A(n4144), .B(n4145), .Z(n1499) );
  NANDN U4845 ( .A(B[325]), .B(n4146), .Z(n4145) );
  NANDN U4846 ( .A(A[325]), .B(n1501), .Z(n4146) );
  NANDN U4847 ( .A(n1501), .B(A[325]), .Z(n4144) );
  AND U4848 ( .A(n4147), .B(n4148), .Z(n1501) );
  NANDN U4849 ( .A(B[324]), .B(n4149), .Z(n4148) );
  NANDN U4850 ( .A(A[324]), .B(n1503), .Z(n4149) );
  NANDN U4851 ( .A(n1503), .B(A[324]), .Z(n4147) );
  AND U4852 ( .A(n4150), .B(n4151), .Z(n1503) );
  NANDN U4853 ( .A(B[323]), .B(n4152), .Z(n4151) );
  NANDN U4854 ( .A(A[323]), .B(n1505), .Z(n4152) );
  NANDN U4855 ( .A(n1505), .B(A[323]), .Z(n4150) );
  AND U4856 ( .A(n4153), .B(n4154), .Z(n1505) );
  NANDN U4857 ( .A(B[322]), .B(n4155), .Z(n4154) );
  NANDN U4858 ( .A(A[322]), .B(n1507), .Z(n4155) );
  NANDN U4859 ( .A(n1507), .B(A[322]), .Z(n4153) );
  AND U4860 ( .A(n4156), .B(n4157), .Z(n1507) );
  NANDN U4861 ( .A(B[321]), .B(n4158), .Z(n4157) );
  NANDN U4862 ( .A(A[321]), .B(n1509), .Z(n4158) );
  NANDN U4863 ( .A(n1509), .B(A[321]), .Z(n4156) );
  AND U4864 ( .A(n4159), .B(n4160), .Z(n1509) );
  NANDN U4865 ( .A(B[320]), .B(n4161), .Z(n4160) );
  NANDN U4866 ( .A(A[320]), .B(n1511), .Z(n4161) );
  NANDN U4867 ( .A(n1511), .B(A[320]), .Z(n4159) );
  AND U4868 ( .A(n4162), .B(n4163), .Z(n1511) );
  NANDN U4869 ( .A(B[319]), .B(n4164), .Z(n4163) );
  NANDN U4870 ( .A(A[319]), .B(n1515), .Z(n4164) );
  NANDN U4871 ( .A(n1515), .B(A[319]), .Z(n4162) );
  AND U4872 ( .A(n4165), .B(n4166), .Z(n1515) );
  NANDN U4873 ( .A(B[318]), .B(n4167), .Z(n4166) );
  NANDN U4874 ( .A(A[318]), .B(n1517), .Z(n4167) );
  NANDN U4875 ( .A(n1517), .B(A[318]), .Z(n4165) );
  AND U4876 ( .A(n4168), .B(n4169), .Z(n1517) );
  NANDN U4877 ( .A(B[317]), .B(n4170), .Z(n4169) );
  NANDN U4878 ( .A(A[317]), .B(n1519), .Z(n4170) );
  NANDN U4879 ( .A(n1519), .B(A[317]), .Z(n4168) );
  AND U4880 ( .A(n4171), .B(n4172), .Z(n1519) );
  NANDN U4881 ( .A(B[316]), .B(n4173), .Z(n4172) );
  NANDN U4882 ( .A(A[316]), .B(n1521), .Z(n4173) );
  NANDN U4883 ( .A(n1521), .B(A[316]), .Z(n4171) );
  AND U4884 ( .A(n4174), .B(n4175), .Z(n1521) );
  NANDN U4885 ( .A(B[315]), .B(n4176), .Z(n4175) );
  NANDN U4886 ( .A(A[315]), .B(n1523), .Z(n4176) );
  NANDN U4887 ( .A(n1523), .B(A[315]), .Z(n4174) );
  AND U4888 ( .A(n4177), .B(n4178), .Z(n1523) );
  NANDN U4889 ( .A(B[314]), .B(n4179), .Z(n4178) );
  NANDN U4890 ( .A(A[314]), .B(n1525), .Z(n4179) );
  NANDN U4891 ( .A(n1525), .B(A[314]), .Z(n4177) );
  AND U4892 ( .A(n4180), .B(n4181), .Z(n1525) );
  NANDN U4893 ( .A(B[313]), .B(n4182), .Z(n4181) );
  NANDN U4894 ( .A(A[313]), .B(n1527), .Z(n4182) );
  NANDN U4895 ( .A(n1527), .B(A[313]), .Z(n4180) );
  AND U4896 ( .A(n4183), .B(n4184), .Z(n1527) );
  NANDN U4897 ( .A(B[312]), .B(n4185), .Z(n4184) );
  NANDN U4898 ( .A(A[312]), .B(n1529), .Z(n4185) );
  NANDN U4899 ( .A(n1529), .B(A[312]), .Z(n4183) );
  AND U4900 ( .A(n4186), .B(n4187), .Z(n1529) );
  NANDN U4901 ( .A(B[311]), .B(n4188), .Z(n4187) );
  NANDN U4902 ( .A(A[311]), .B(n1531), .Z(n4188) );
  NANDN U4903 ( .A(n1531), .B(A[311]), .Z(n4186) );
  AND U4904 ( .A(n4189), .B(n4190), .Z(n1531) );
  NANDN U4905 ( .A(B[310]), .B(n4191), .Z(n4190) );
  NANDN U4906 ( .A(A[310]), .B(n1533), .Z(n4191) );
  NANDN U4907 ( .A(n1533), .B(A[310]), .Z(n4189) );
  AND U4908 ( .A(n4192), .B(n4193), .Z(n1533) );
  NANDN U4909 ( .A(B[309]), .B(n4194), .Z(n4193) );
  NANDN U4910 ( .A(A[309]), .B(n1537), .Z(n4194) );
  NANDN U4911 ( .A(n1537), .B(A[309]), .Z(n4192) );
  AND U4912 ( .A(n4195), .B(n4196), .Z(n1537) );
  NANDN U4913 ( .A(B[308]), .B(n4197), .Z(n4196) );
  NANDN U4914 ( .A(A[308]), .B(n1539), .Z(n4197) );
  NANDN U4915 ( .A(n1539), .B(A[308]), .Z(n4195) );
  AND U4916 ( .A(n4198), .B(n4199), .Z(n1539) );
  NANDN U4917 ( .A(B[307]), .B(n4200), .Z(n4199) );
  NANDN U4918 ( .A(A[307]), .B(n1541), .Z(n4200) );
  NANDN U4919 ( .A(n1541), .B(A[307]), .Z(n4198) );
  AND U4920 ( .A(n4201), .B(n4202), .Z(n1541) );
  NANDN U4921 ( .A(B[306]), .B(n4203), .Z(n4202) );
  NANDN U4922 ( .A(A[306]), .B(n1543), .Z(n4203) );
  NANDN U4923 ( .A(n1543), .B(A[306]), .Z(n4201) );
  AND U4924 ( .A(n4204), .B(n4205), .Z(n1543) );
  NANDN U4925 ( .A(B[305]), .B(n4206), .Z(n4205) );
  NANDN U4926 ( .A(A[305]), .B(n1545), .Z(n4206) );
  NANDN U4927 ( .A(n1545), .B(A[305]), .Z(n4204) );
  AND U4928 ( .A(n4207), .B(n4208), .Z(n1545) );
  NANDN U4929 ( .A(B[304]), .B(n4209), .Z(n4208) );
  NANDN U4930 ( .A(A[304]), .B(n1547), .Z(n4209) );
  NANDN U4931 ( .A(n1547), .B(A[304]), .Z(n4207) );
  AND U4932 ( .A(n4210), .B(n4211), .Z(n1547) );
  NANDN U4933 ( .A(B[303]), .B(n4212), .Z(n4211) );
  NANDN U4934 ( .A(A[303]), .B(n1549), .Z(n4212) );
  NANDN U4935 ( .A(n1549), .B(A[303]), .Z(n4210) );
  AND U4936 ( .A(n4213), .B(n4214), .Z(n1549) );
  NANDN U4937 ( .A(B[302]), .B(n4215), .Z(n4214) );
  NANDN U4938 ( .A(A[302]), .B(n1551), .Z(n4215) );
  NANDN U4939 ( .A(n1551), .B(A[302]), .Z(n4213) );
  AND U4940 ( .A(n4216), .B(n4217), .Z(n1551) );
  NANDN U4941 ( .A(B[301]), .B(n4218), .Z(n4217) );
  NANDN U4942 ( .A(A[301]), .B(n1553), .Z(n4218) );
  NANDN U4943 ( .A(n1553), .B(A[301]), .Z(n4216) );
  AND U4944 ( .A(n4219), .B(n4220), .Z(n1553) );
  NANDN U4945 ( .A(B[300]), .B(n4221), .Z(n4220) );
  NANDN U4946 ( .A(A[300]), .B(n1555), .Z(n4221) );
  NANDN U4947 ( .A(n1555), .B(A[300]), .Z(n4219) );
  AND U4948 ( .A(n4222), .B(n4223), .Z(n1555) );
  NANDN U4949 ( .A(B[299]), .B(n4224), .Z(n4223) );
  NANDN U4950 ( .A(A[299]), .B(n1561), .Z(n4224) );
  NANDN U4951 ( .A(n1561), .B(A[299]), .Z(n4222) );
  AND U4952 ( .A(n4225), .B(n4226), .Z(n1561) );
  NANDN U4953 ( .A(B[298]), .B(n4227), .Z(n4226) );
  NANDN U4954 ( .A(A[298]), .B(n1563), .Z(n4227) );
  NANDN U4955 ( .A(n1563), .B(A[298]), .Z(n4225) );
  AND U4956 ( .A(n4228), .B(n4229), .Z(n1563) );
  NANDN U4957 ( .A(B[297]), .B(n4230), .Z(n4229) );
  NANDN U4958 ( .A(A[297]), .B(n1565), .Z(n4230) );
  NANDN U4959 ( .A(n1565), .B(A[297]), .Z(n4228) );
  AND U4960 ( .A(n4231), .B(n4232), .Z(n1565) );
  NANDN U4961 ( .A(B[296]), .B(n4233), .Z(n4232) );
  NANDN U4962 ( .A(A[296]), .B(n1567), .Z(n4233) );
  NANDN U4963 ( .A(n1567), .B(A[296]), .Z(n4231) );
  AND U4964 ( .A(n4234), .B(n4235), .Z(n1567) );
  NANDN U4965 ( .A(B[295]), .B(n4236), .Z(n4235) );
  NANDN U4966 ( .A(A[295]), .B(n1569), .Z(n4236) );
  NANDN U4967 ( .A(n1569), .B(A[295]), .Z(n4234) );
  AND U4968 ( .A(n4237), .B(n4238), .Z(n1569) );
  NANDN U4969 ( .A(B[294]), .B(n4239), .Z(n4238) );
  NANDN U4970 ( .A(A[294]), .B(n1571), .Z(n4239) );
  NANDN U4971 ( .A(n1571), .B(A[294]), .Z(n4237) );
  AND U4972 ( .A(n4240), .B(n4241), .Z(n1571) );
  NANDN U4973 ( .A(B[293]), .B(n4242), .Z(n4241) );
  NANDN U4974 ( .A(A[293]), .B(n1573), .Z(n4242) );
  NANDN U4975 ( .A(n1573), .B(A[293]), .Z(n4240) );
  AND U4976 ( .A(n4243), .B(n4244), .Z(n1573) );
  NANDN U4977 ( .A(B[292]), .B(n4245), .Z(n4244) );
  NANDN U4978 ( .A(A[292]), .B(n1575), .Z(n4245) );
  NANDN U4979 ( .A(n1575), .B(A[292]), .Z(n4243) );
  AND U4980 ( .A(n4246), .B(n4247), .Z(n1575) );
  NANDN U4981 ( .A(B[291]), .B(n4248), .Z(n4247) );
  NANDN U4982 ( .A(A[291]), .B(n1577), .Z(n4248) );
  NANDN U4983 ( .A(n1577), .B(A[291]), .Z(n4246) );
  AND U4984 ( .A(n4249), .B(n4250), .Z(n1577) );
  NANDN U4985 ( .A(B[290]), .B(n4251), .Z(n4250) );
  NANDN U4986 ( .A(A[290]), .B(n1579), .Z(n4251) );
  NANDN U4987 ( .A(n1579), .B(A[290]), .Z(n4249) );
  AND U4988 ( .A(n4252), .B(n4253), .Z(n1579) );
  NANDN U4989 ( .A(B[289]), .B(n4254), .Z(n4253) );
  NANDN U4990 ( .A(A[289]), .B(n1583), .Z(n4254) );
  NANDN U4991 ( .A(n1583), .B(A[289]), .Z(n4252) );
  AND U4992 ( .A(n4255), .B(n4256), .Z(n1583) );
  NANDN U4993 ( .A(B[288]), .B(n4257), .Z(n4256) );
  NANDN U4994 ( .A(A[288]), .B(n1585), .Z(n4257) );
  NANDN U4995 ( .A(n1585), .B(A[288]), .Z(n4255) );
  AND U4996 ( .A(n4258), .B(n4259), .Z(n1585) );
  NANDN U4997 ( .A(B[287]), .B(n4260), .Z(n4259) );
  NANDN U4998 ( .A(A[287]), .B(n1587), .Z(n4260) );
  NANDN U4999 ( .A(n1587), .B(A[287]), .Z(n4258) );
  AND U5000 ( .A(n4261), .B(n4262), .Z(n1587) );
  NANDN U5001 ( .A(B[286]), .B(n4263), .Z(n4262) );
  NANDN U5002 ( .A(A[286]), .B(n1589), .Z(n4263) );
  NANDN U5003 ( .A(n1589), .B(A[286]), .Z(n4261) );
  AND U5004 ( .A(n4264), .B(n4265), .Z(n1589) );
  NANDN U5005 ( .A(B[285]), .B(n4266), .Z(n4265) );
  NANDN U5006 ( .A(A[285]), .B(n1591), .Z(n4266) );
  NANDN U5007 ( .A(n1591), .B(A[285]), .Z(n4264) );
  AND U5008 ( .A(n4267), .B(n4268), .Z(n1591) );
  NANDN U5009 ( .A(B[284]), .B(n4269), .Z(n4268) );
  NANDN U5010 ( .A(A[284]), .B(n1593), .Z(n4269) );
  NANDN U5011 ( .A(n1593), .B(A[284]), .Z(n4267) );
  AND U5012 ( .A(n4270), .B(n4271), .Z(n1593) );
  NANDN U5013 ( .A(B[283]), .B(n4272), .Z(n4271) );
  NANDN U5014 ( .A(A[283]), .B(n1595), .Z(n4272) );
  NANDN U5015 ( .A(n1595), .B(A[283]), .Z(n4270) );
  AND U5016 ( .A(n4273), .B(n4274), .Z(n1595) );
  NANDN U5017 ( .A(B[282]), .B(n4275), .Z(n4274) );
  NANDN U5018 ( .A(A[282]), .B(n1597), .Z(n4275) );
  NANDN U5019 ( .A(n1597), .B(A[282]), .Z(n4273) );
  AND U5020 ( .A(n4276), .B(n4277), .Z(n1597) );
  NANDN U5021 ( .A(B[281]), .B(n4278), .Z(n4277) );
  NANDN U5022 ( .A(A[281]), .B(n1599), .Z(n4278) );
  NANDN U5023 ( .A(n1599), .B(A[281]), .Z(n4276) );
  AND U5024 ( .A(n4279), .B(n4280), .Z(n1599) );
  NANDN U5025 ( .A(B[280]), .B(n4281), .Z(n4280) );
  NANDN U5026 ( .A(A[280]), .B(n1601), .Z(n4281) );
  NANDN U5027 ( .A(n1601), .B(A[280]), .Z(n4279) );
  AND U5028 ( .A(n4282), .B(n4283), .Z(n1601) );
  NANDN U5029 ( .A(B[279]), .B(n4284), .Z(n4283) );
  NANDN U5030 ( .A(A[279]), .B(n1605), .Z(n4284) );
  NANDN U5031 ( .A(n1605), .B(A[279]), .Z(n4282) );
  AND U5032 ( .A(n4285), .B(n4286), .Z(n1605) );
  NANDN U5033 ( .A(B[278]), .B(n4287), .Z(n4286) );
  NANDN U5034 ( .A(A[278]), .B(n1607), .Z(n4287) );
  NANDN U5035 ( .A(n1607), .B(A[278]), .Z(n4285) );
  AND U5036 ( .A(n4288), .B(n4289), .Z(n1607) );
  NANDN U5037 ( .A(B[277]), .B(n4290), .Z(n4289) );
  NANDN U5038 ( .A(A[277]), .B(n1609), .Z(n4290) );
  NANDN U5039 ( .A(n1609), .B(A[277]), .Z(n4288) );
  AND U5040 ( .A(n4291), .B(n4292), .Z(n1609) );
  NANDN U5041 ( .A(B[276]), .B(n4293), .Z(n4292) );
  NANDN U5042 ( .A(A[276]), .B(n1611), .Z(n4293) );
  NANDN U5043 ( .A(n1611), .B(A[276]), .Z(n4291) );
  AND U5044 ( .A(n4294), .B(n4295), .Z(n1611) );
  NANDN U5045 ( .A(B[275]), .B(n4296), .Z(n4295) );
  NANDN U5046 ( .A(A[275]), .B(n1613), .Z(n4296) );
  NANDN U5047 ( .A(n1613), .B(A[275]), .Z(n4294) );
  AND U5048 ( .A(n4297), .B(n4298), .Z(n1613) );
  NANDN U5049 ( .A(B[274]), .B(n4299), .Z(n4298) );
  NANDN U5050 ( .A(A[274]), .B(n1615), .Z(n4299) );
  NANDN U5051 ( .A(n1615), .B(A[274]), .Z(n4297) );
  AND U5052 ( .A(n4300), .B(n4301), .Z(n1615) );
  NANDN U5053 ( .A(B[273]), .B(n4302), .Z(n4301) );
  NANDN U5054 ( .A(A[273]), .B(n1617), .Z(n4302) );
  NANDN U5055 ( .A(n1617), .B(A[273]), .Z(n4300) );
  AND U5056 ( .A(n4303), .B(n4304), .Z(n1617) );
  NANDN U5057 ( .A(B[272]), .B(n4305), .Z(n4304) );
  NANDN U5058 ( .A(A[272]), .B(n1619), .Z(n4305) );
  NANDN U5059 ( .A(n1619), .B(A[272]), .Z(n4303) );
  AND U5060 ( .A(n4306), .B(n4307), .Z(n1619) );
  NANDN U5061 ( .A(B[271]), .B(n4308), .Z(n4307) );
  NANDN U5062 ( .A(A[271]), .B(n1621), .Z(n4308) );
  NANDN U5063 ( .A(n1621), .B(A[271]), .Z(n4306) );
  AND U5064 ( .A(n4309), .B(n4310), .Z(n1621) );
  NANDN U5065 ( .A(B[270]), .B(n4311), .Z(n4310) );
  NANDN U5066 ( .A(A[270]), .B(n1623), .Z(n4311) );
  NANDN U5067 ( .A(n1623), .B(A[270]), .Z(n4309) );
  AND U5068 ( .A(n4312), .B(n4313), .Z(n1623) );
  NANDN U5069 ( .A(B[269]), .B(n4314), .Z(n4313) );
  NANDN U5070 ( .A(A[269]), .B(n1627), .Z(n4314) );
  NANDN U5071 ( .A(n1627), .B(A[269]), .Z(n4312) );
  AND U5072 ( .A(n4315), .B(n4316), .Z(n1627) );
  NANDN U5073 ( .A(B[268]), .B(n4317), .Z(n4316) );
  NANDN U5074 ( .A(A[268]), .B(n1629), .Z(n4317) );
  NANDN U5075 ( .A(n1629), .B(A[268]), .Z(n4315) );
  AND U5076 ( .A(n4318), .B(n4319), .Z(n1629) );
  NANDN U5077 ( .A(B[267]), .B(n4320), .Z(n4319) );
  NANDN U5078 ( .A(A[267]), .B(n1631), .Z(n4320) );
  NANDN U5079 ( .A(n1631), .B(A[267]), .Z(n4318) );
  AND U5080 ( .A(n4321), .B(n4322), .Z(n1631) );
  NANDN U5081 ( .A(B[266]), .B(n4323), .Z(n4322) );
  NANDN U5082 ( .A(A[266]), .B(n1633), .Z(n4323) );
  NANDN U5083 ( .A(n1633), .B(A[266]), .Z(n4321) );
  AND U5084 ( .A(n4324), .B(n4325), .Z(n1633) );
  NANDN U5085 ( .A(B[265]), .B(n4326), .Z(n4325) );
  NANDN U5086 ( .A(A[265]), .B(n1635), .Z(n4326) );
  NANDN U5087 ( .A(n1635), .B(A[265]), .Z(n4324) );
  AND U5088 ( .A(n4327), .B(n4328), .Z(n1635) );
  NANDN U5089 ( .A(B[264]), .B(n4329), .Z(n4328) );
  NANDN U5090 ( .A(A[264]), .B(n1637), .Z(n4329) );
  NANDN U5091 ( .A(n1637), .B(A[264]), .Z(n4327) );
  AND U5092 ( .A(n4330), .B(n4331), .Z(n1637) );
  NANDN U5093 ( .A(B[263]), .B(n4332), .Z(n4331) );
  NANDN U5094 ( .A(A[263]), .B(n1639), .Z(n4332) );
  NANDN U5095 ( .A(n1639), .B(A[263]), .Z(n4330) );
  AND U5096 ( .A(n4333), .B(n4334), .Z(n1639) );
  NANDN U5097 ( .A(B[262]), .B(n4335), .Z(n4334) );
  NANDN U5098 ( .A(A[262]), .B(n1641), .Z(n4335) );
  NANDN U5099 ( .A(n1641), .B(A[262]), .Z(n4333) );
  AND U5100 ( .A(n4336), .B(n4337), .Z(n1641) );
  NANDN U5101 ( .A(B[261]), .B(n4338), .Z(n4337) );
  NANDN U5102 ( .A(A[261]), .B(n1643), .Z(n4338) );
  NANDN U5103 ( .A(n1643), .B(A[261]), .Z(n4336) );
  AND U5104 ( .A(n4339), .B(n4340), .Z(n1643) );
  NANDN U5105 ( .A(B[260]), .B(n4341), .Z(n4340) );
  NANDN U5106 ( .A(A[260]), .B(n1645), .Z(n4341) );
  NANDN U5107 ( .A(n1645), .B(A[260]), .Z(n4339) );
  AND U5108 ( .A(n4342), .B(n4343), .Z(n1645) );
  NANDN U5109 ( .A(B[259]), .B(n4344), .Z(n4343) );
  NANDN U5110 ( .A(A[259]), .B(n1649), .Z(n4344) );
  NANDN U5111 ( .A(n1649), .B(A[259]), .Z(n4342) );
  AND U5112 ( .A(n4345), .B(n4346), .Z(n1649) );
  NANDN U5113 ( .A(B[258]), .B(n4347), .Z(n4346) );
  NANDN U5114 ( .A(A[258]), .B(n1651), .Z(n4347) );
  NANDN U5115 ( .A(n1651), .B(A[258]), .Z(n4345) );
  AND U5116 ( .A(n4348), .B(n4349), .Z(n1651) );
  NANDN U5117 ( .A(B[257]), .B(n4350), .Z(n4349) );
  NANDN U5118 ( .A(A[257]), .B(n1653), .Z(n4350) );
  NANDN U5119 ( .A(n1653), .B(A[257]), .Z(n4348) );
  AND U5120 ( .A(n4351), .B(n4352), .Z(n1653) );
  NANDN U5121 ( .A(B[256]), .B(n4353), .Z(n4352) );
  NANDN U5122 ( .A(A[256]), .B(n1655), .Z(n4353) );
  NANDN U5123 ( .A(n1655), .B(A[256]), .Z(n4351) );
  AND U5124 ( .A(n4354), .B(n4355), .Z(n1655) );
  NANDN U5125 ( .A(B[255]), .B(n4356), .Z(n4355) );
  NANDN U5126 ( .A(A[255]), .B(n1657), .Z(n4356) );
  NANDN U5127 ( .A(n1657), .B(A[255]), .Z(n4354) );
  AND U5128 ( .A(n4357), .B(n4358), .Z(n1657) );
  NANDN U5129 ( .A(B[254]), .B(n4359), .Z(n4358) );
  NANDN U5130 ( .A(A[254]), .B(n1659), .Z(n4359) );
  NANDN U5131 ( .A(n1659), .B(A[254]), .Z(n4357) );
  AND U5132 ( .A(n4360), .B(n4361), .Z(n1659) );
  NANDN U5133 ( .A(B[253]), .B(n4362), .Z(n4361) );
  NANDN U5134 ( .A(A[253]), .B(n1661), .Z(n4362) );
  NANDN U5135 ( .A(n1661), .B(A[253]), .Z(n4360) );
  AND U5136 ( .A(n4363), .B(n4364), .Z(n1661) );
  NANDN U5137 ( .A(B[252]), .B(n4365), .Z(n4364) );
  NANDN U5138 ( .A(A[252]), .B(n1663), .Z(n4365) );
  NANDN U5139 ( .A(n1663), .B(A[252]), .Z(n4363) );
  AND U5140 ( .A(n4366), .B(n4367), .Z(n1663) );
  NANDN U5141 ( .A(B[251]), .B(n4368), .Z(n4367) );
  NANDN U5142 ( .A(A[251]), .B(n1665), .Z(n4368) );
  NANDN U5143 ( .A(n1665), .B(A[251]), .Z(n4366) );
  AND U5144 ( .A(n4369), .B(n4370), .Z(n1665) );
  NANDN U5145 ( .A(B[250]), .B(n4371), .Z(n4370) );
  NANDN U5146 ( .A(A[250]), .B(n1667), .Z(n4371) );
  NANDN U5147 ( .A(n1667), .B(A[250]), .Z(n4369) );
  AND U5148 ( .A(n4372), .B(n4373), .Z(n1667) );
  NANDN U5149 ( .A(B[249]), .B(n4374), .Z(n4373) );
  NANDN U5150 ( .A(A[249]), .B(n1671), .Z(n4374) );
  NANDN U5151 ( .A(n1671), .B(A[249]), .Z(n4372) );
  AND U5152 ( .A(n4375), .B(n4376), .Z(n1671) );
  NANDN U5153 ( .A(B[248]), .B(n4377), .Z(n4376) );
  NANDN U5154 ( .A(A[248]), .B(n1673), .Z(n4377) );
  NANDN U5155 ( .A(n1673), .B(A[248]), .Z(n4375) );
  AND U5156 ( .A(n4378), .B(n4379), .Z(n1673) );
  NANDN U5157 ( .A(B[247]), .B(n4380), .Z(n4379) );
  NANDN U5158 ( .A(A[247]), .B(n1675), .Z(n4380) );
  NANDN U5159 ( .A(n1675), .B(A[247]), .Z(n4378) );
  AND U5160 ( .A(n4381), .B(n4382), .Z(n1675) );
  NANDN U5161 ( .A(B[246]), .B(n4383), .Z(n4382) );
  NANDN U5162 ( .A(A[246]), .B(n1677), .Z(n4383) );
  NANDN U5163 ( .A(n1677), .B(A[246]), .Z(n4381) );
  AND U5164 ( .A(n4384), .B(n4385), .Z(n1677) );
  NANDN U5165 ( .A(B[245]), .B(n4386), .Z(n4385) );
  NANDN U5166 ( .A(A[245]), .B(n1679), .Z(n4386) );
  NANDN U5167 ( .A(n1679), .B(A[245]), .Z(n4384) );
  AND U5168 ( .A(n4387), .B(n4388), .Z(n1679) );
  NANDN U5169 ( .A(B[244]), .B(n4389), .Z(n4388) );
  NANDN U5170 ( .A(A[244]), .B(n1681), .Z(n4389) );
  NANDN U5171 ( .A(n1681), .B(A[244]), .Z(n4387) );
  AND U5172 ( .A(n4390), .B(n4391), .Z(n1681) );
  NANDN U5173 ( .A(B[243]), .B(n4392), .Z(n4391) );
  NANDN U5174 ( .A(A[243]), .B(n1683), .Z(n4392) );
  NANDN U5175 ( .A(n1683), .B(A[243]), .Z(n4390) );
  AND U5176 ( .A(n4393), .B(n4394), .Z(n1683) );
  NANDN U5177 ( .A(B[242]), .B(n4395), .Z(n4394) );
  NANDN U5178 ( .A(A[242]), .B(n1685), .Z(n4395) );
  NANDN U5179 ( .A(n1685), .B(A[242]), .Z(n4393) );
  AND U5180 ( .A(n4396), .B(n4397), .Z(n1685) );
  NANDN U5181 ( .A(B[241]), .B(n4398), .Z(n4397) );
  NANDN U5182 ( .A(A[241]), .B(n1687), .Z(n4398) );
  NANDN U5183 ( .A(n1687), .B(A[241]), .Z(n4396) );
  AND U5184 ( .A(n4399), .B(n4400), .Z(n1687) );
  NANDN U5185 ( .A(B[240]), .B(n4401), .Z(n4400) );
  NANDN U5186 ( .A(A[240]), .B(n1689), .Z(n4401) );
  NANDN U5187 ( .A(n1689), .B(A[240]), .Z(n4399) );
  AND U5188 ( .A(n4402), .B(n4403), .Z(n1689) );
  NANDN U5189 ( .A(B[239]), .B(n4404), .Z(n4403) );
  NANDN U5190 ( .A(A[239]), .B(n1693), .Z(n4404) );
  NANDN U5191 ( .A(n1693), .B(A[239]), .Z(n4402) );
  AND U5192 ( .A(n4405), .B(n4406), .Z(n1693) );
  NANDN U5193 ( .A(B[238]), .B(n4407), .Z(n4406) );
  NANDN U5194 ( .A(A[238]), .B(n1695), .Z(n4407) );
  NANDN U5195 ( .A(n1695), .B(A[238]), .Z(n4405) );
  AND U5196 ( .A(n4408), .B(n4409), .Z(n1695) );
  NANDN U5197 ( .A(B[237]), .B(n4410), .Z(n4409) );
  NANDN U5198 ( .A(A[237]), .B(n1697), .Z(n4410) );
  NANDN U5199 ( .A(n1697), .B(A[237]), .Z(n4408) );
  AND U5200 ( .A(n4411), .B(n4412), .Z(n1697) );
  NANDN U5201 ( .A(B[236]), .B(n4413), .Z(n4412) );
  NANDN U5202 ( .A(A[236]), .B(n1699), .Z(n4413) );
  NANDN U5203 ( .A(n1699), .B(A[236]), .Z(n4411) );
  AND U5204 ( .A(n4414), .B(n4415), .Z(n1699) );
  NANDN U5205 ( .A(B[235]), .B(n4416), .Z(n4415) );
  NANDN U5206 ( .A(A[235]), .B(n1701), .Z(n4416) );
  NANDN U5207 ( .A(n1701), .B(A[235]), .Z(n4414) );
  AND U5208 ( .A(n4417), .B(n4418), .Z(n1701) );
  NANDN U5209 ( .A(B[234]), .B(n4419), .Z(n4418) );
  NANDN U5210 ( .A(A[234]), .B(n1703), .Z(n4419) );
  NANDN U5211 ( .A(n1703), .B(A[234]), .Z(n4417) );
  AND U5212 ( .A(n4420), .B(n4421), .Z(n1703) );
  NANDN U5213 ( .A(B[233]), .B(n4422), .Z(n4421) );
  NANDN U5214 ( .A(A[233]), .B(n1705), .Z(n4422) );
  NANDN U5215 ( .A(n1705), .B(A[233]), .Z(n4420) );
  AND U5216 ( .A(n4423), .B(n4424), .Z(n1705) );
  NANDN U5217 ( .A(B[232]), .B(n4425), .Z(n4424) );
  NANDN U5218 ( .A(A[232]), .B(n1707), .Z(n4425) );
  NANDN U5219 ( .A(n1707), .B(A[232]), .Z(n4423) );
  AND U5220 ( .A(n4426), .B(n4427), .Z(n1707) );
  NANDN U5221 ( .A(B[231]), .B(n4428), .Z(n4427) );
  NANDN U5222 ( .A(A[231]), .B(n1709), .Z(n4428) );
  NANDN U5223 ( .A(n1709), .B(A[231]), .Z(n4426) );
  AND U5224 ( .A(n4429), .B(n4430), .Z(n1709) );
  NANDN U5225 ( .A(B[230]), .B(n4431), .Z(n4430) );
  NANDN U5226 ( .A(A[230]), .B(n1711), .Z(n4431) );
  NANDN U5227 ( .A(n1711), .B(A[230]), .Z(n4429) );
  AND U5228 ( .A(n4432), .B(n4433), .Z(n1711) );
  NANDN U5229 ( .A(B[229]), .B(n4434), .Z(n4433) );
  NANDN U5230 ( .A(A[229]), .B(n1715), .Z(n4434) );
  NANDN U5231 ( .A(n1715), .B(A[229]), .Z(n4432) );
  AND U5232 ( .A(n4435), .B(n4436), .Z(n1715) );
  NANDN U5233 ( .A(B[228]), .B(n4437), .Z(n4436) );
  NANDN U5234 ( .A(A[228]), .B(n1717), .Z(n4437) );
  NANDN U5235 ( .A(n1717), .B(A[228]), .Z(n4435) );
  AND U5236 ( .A(n4438), .B(n4439), .Z(n1717) );
  NANDN U5237 ( .A(B[227]), .B(n4440), .Z(n4439) );
  NANDN U5238 ( .A(A[227]), .B(n1719), .Z(n4440) );
  NANDN U5239 ( .A(n1719), .B(A[227]), .Z(n4438) );
  AND U5240 ( .A(n4441), .B(n4442), .Z(n1719) );
  NANDN U5241 ( .A(B[226]), .B(n4443), .Z(n4442) );
  NANDN U5242 ( .A(A[226]), .B(n1721), .Z(n4443) );
  NANDN U5243 ( .A(n1721), .B(A[226]), .Z(n4441) );
  AND U5244 ( .A(n4444), .B(n4445), .Z(n1721) );
  NANDN U5245 ( .A(B[225]), .B(n4446), .Z(n4445) );
  NANDN U5246 ( .A(A[225]), .B(n1723), .Z(n4446) );
  NANDN U5247 ( .A(n1723), .B(A[225]), .Z(n4444) );
  AND U5248 ( .A(n4447), .B(n4448), .Z(n1723) );
  NANDN U5249 ( .A(B[224]), .B(n4449), .Z(n4448) );
  NANDN U5250 ( .A(A[224]), .B(n1725), .Z(n4449) );
  NANDN U5251 ( .A(n1725), .B(A[224]), .Z(n4447) );
  AND U5252 ( .A(n4450), .B(n4451), .Z(n1725) );
  NANDN U5253 ( .A(B[223]), .B(n4452), .Z(n4451) );
  NANDN U5254 ( .A(A[223]), .B(n1727), .Z(n4452) );
  NANDN U5255 ( .A(n1727), .B(A[223]), .Z(n4450) );
  AND U5256 ( .A(n4453), .B(n4454), .Z(n1727) );
  NANDN U5257 ( .A(B[222]), .B(n4455), .Z(n4454) );
  NANDN U5258 ( .A(A[222]), .B(n1729), .Z(n4455) );
  NANDN U5259 ( .A(n1729), .B(A[222]), .Z(n4453) );
  AND U5260 ( .A(n4456), .B(n4457), .Z(n1729) );
  NANDN U5261 ( .A(B[221]), .B(n4458), .Z(n4457) );
  NANDN U5262 ( .A(A[221]), .B(n1731), .Z(n4458) );
  NANDN U5263 ( .A(n1731), .B(A[221]), .Z(n4456) );
  AND U5264 ( .A(n4459), .B(n4460), .Z(n1731) );
  NANDN U5265 ( .A(B[220]), .B(n4461), .Z(n4460) );
  NANDN U5266 ( .A(A[220]), .B(n1733), .Z(n4461) );
  NANDN U5267 ( .A(n1733), .B(A[220]), .Z(n4459) );
  AND U5268 ( .A(n4462), .B(n4463), .Z(n1733) );
  NANDN U5269 ( .A(B[219]), .B(n4464), .Z(n4463) );
  NANDN U5270 ( .A(A[219]), .B(n1737), .Z(n4464) );
  NANDN U5271 ( .A(n1737), .B(A[219]), .Z(n4462) );
  AND U5272 ( .A(n4465), .B(n4466), .Z(n1737) );
  NANDN U5273 ( .A(B[218]), .B(n4467), .Z(n4466) );
  NANDN U5274 ( .A(A[218]), .B(n1739), .Z(n4467) );
  NANDN U5275 ( .A(n1739), .B(A[218]), .Z(n4465) );
  AND U5276 ( .A(n4468), .B(n4469), .Z(n1739) );
  NANDN U5277 ( .A(B[217]), .B(n4470), .Z(n4469) );
  NANDN U5278 ( .A(A[217]), .B(n1741), .Z(n4470) );
  NANDN U5279 ( .A(n1741), .B(A[217]), .Z(n4468) );
  AND U5280 ( .A(n4471), .B(n4472), .Z(n1741) );
  NANDN U5281 ( .A(B[216]), .B(n4473), .Z(n4472) );
  NANDN U5282 ( .A(A[216]), .B(n1743), .Z(n4473) );
  NANDN U5283 ( .A(n1743), .B(A[216]), .Z(n4471) );
  AND U5284 ( .A(n4474), .B(n4475), .Z(n1743) );
  NANDN U5285 ( .A(B[215]), .B(n4476), .Z(n4475) );
  NANDN U5286 ( .A(A[215]), .B(n1745), .Z(n4476) );
  NANDN U5287 ( .A(n1745), .B(A[215]), .Z(n4474) );
  AND U5288 ( .A(n4477), .B(n4478), .Z(n1745) );
  NANDN U5289 ( .A(B[214]), .B(n4479), .Z(n4478) );
  NANDN U5290 ( .A(A[214]), .B(n1747), .Z(n4479) );
  NANDN U5291 ( .A(n1747), .B(A[214]), .Z(n4477) );
  AND U5292 ( .A(n4480), .B(n4481), .Z(n1747) );
  NANDN U5293 ( .A(B[213]), .B(n4482), .Z(n4481) );
  NANDN U5294 ( .A(A[213]), .B(n1749), .Z(n4482) );
  NANDN U5295 ( .A(n1749), .B(A[213]), .Z(n4480) );
  AND U5296 ( .A(n4483), .B(n4484), .Z(n1749) );
  NANDN U5297 ( .A(B[212]), .B(n4485), .Z(n4484) );
  NANDN U5298 ( .A(A[212]), .B(n1751), .Z(n4485) );
  NANDN U5299 ( .A(n1751), .B(A[212]), .Z(n4483) );
  AND U5300 ( .A(n4486), .B(n4487), .Z(n1751) );
  NANDN U5301 ( .A(B[211]), .B(n4488), .Z(n4487) );
  NANDN U5302 ( .A(A[211]), .B(n1753), .Z(n4488) );
  NANDN U5303 ( .A(n1753), .B(A[211]), .Z(n4486) );
  AND U5304 ( .A(n4489), .B(n4490), .Z(n1753) );
  NANDN U5305 ( .A(B[210]), .B(n4491), .Z(n4490) );
  NANDN U5306 ( .A(A[210]), .B(n1755), .Z(n4491) );
  NANDN U5307 ( .A(n1755), .B(A[210]), .Z(n4489) );
  AND U5308 ( .A(n4492), .B(n4493), .Z(n1755) );
  NANDN U5309 ( .A(B[209]), .B(n4494), .Z(n4493) );
  NANDN U5310 ( .A(A[209]), .B(n1759), .Z(n4494) );
  NANDN U5311 ( .A(n1759), .B(A[209]), .Z(n4492) );
  AND U5312 ( .A(n4495), .B(n4496), .Z(n1759) );
  NANDN U5313 ( .A(B[208]), .B(n4497), .Z(n4496) );
  NANDN U5314 ( .A(A[208]), .B(n1761), .Z(n4497) );
  NANDN U5315 ( .A(n1761), .B(A[208]), .Z(n4495) );
  AND U5316 ( .A(n4498), .B(n4499), .Z(n1761) );
  NANDN U5317 ( .A(B[207]), .B(n4500), .Z(n4499) );
  NANDN U5318 ( .A(A[207]), .B(n1763), .Z(n4500) );
  NANDN U5319 ( .A(n1763), .B(A[207]), .Z(n4498) );
  AND U5320 ( .A(n4501), .B(n4502), .Z(n1763) );
  NANDN U5321 ( .A(B[206]), .B(n4503), .Z(n4502) );
  NANDN U5322 ( .A(A[206]), .B(n1765), .Z(n4503) );
  NANDN U5323 ( .A(n1765), .B(A[206]), .Z(n4501) );
  AND U5324 ( .A(n4504), .B(n4505), .Z(n1765) );
  NANDN U5325 ( .A(B[205]), .B(n4506), .Z(n4505) );
  NANDN U5326 ( .A(A[205]), .B(n1767), .Z(n4506) );
  NANDN U5327 ( .A(n1767), .B(A[205]), .Z(n4504) );
  AND U5328 ( .A(n4507), .B(n4508), .Z(n1767) );
  NANDN U5329 ( .A(B[204]), .B(n4509), .Z(n4508) );
  NANDN U5330 ( .A(A[204]), .B(n1769), .Z(n4509) );
  NANDN U5331 ( .A(n1769), .B(A[204]), .Z(n4507) );
  AND U5332 ( .A(n4510), .B(n4511), .Z(n1769) );
  NANDN U5333 ( .A(B[203]), .B(n4512), .Z(n4511) );
  NANDN U5334 ( .A(A[203]), .B(n1771), .Z(n4512) );
  NANDN U5335 ( .A(n1771), .B(A[203]), .Z(n4510) );
  AND U5336 ( .A(n4513), .B(n4514), .Z(n1771) );
  NANDN U5337 ( .A(B[202]), .B(n4515), .Z(n4514) );
  NANDN U5338 ( .A(A[202]), .B(n1773), .Z(n4515) );
  NANDN U5339 ( .A(n1773), .B(A[202]), .Z(n4513) );
  AND U5340 ( .A(n4516), .B(n4517), .Z(n1773) );
  NANDN U5341 ( .A(B[201]), .B(n4518), .Z(n4517) );
  NANDN U5342 ( .A(A[201]), .B(n1775), .Z(n4518) );
  NANDN U5343 ( .A(n1775), .B(A[201]), .Z(n4516) );
  AND U5344 ( .A(n4519), .B(n4520), .Z(n1775) );
  NANDN U5345 ( .A(B[200]), .B(n4521), .Z(n4520) );
  NANDN U5346 ( .A(A[200]), .B(n1777), .Z(n4521) );
  NANDN U5347 ( .A(n1777), .B(A[200]), .Z(n4519) );
  AND U5348 ( .A(n4522), .B(n4523), .Z(n1777) );
  NANDN U5349 ( .A(B[199]), .B(n4524), .Z(n4523) );
  NANDN U5350 ( .A(A[199]), .B(n1782), .Z(n4524) );
  NANDN U5351 ( .A(n1782), .B(A[199]), .Z(n4522) );
  AND U5352 ( .A(n4525), .B(n4526), .Z(n1782) );
  NANDN U5353 ( .A(B[198]), .B(n4527), .Z(n4526) );
  NANDN U5354 ( .A(A[198]), .B(n1784), .Z(n4527) );
  NANDN U5355 ( .A(n1784), .B(A[198]), .Z(n4525) );
  AND U5356 ( .A(n4528), .B(n4529), .Z(n1784) );
  NANDN U5357 ( .A(B[197]), .B(n4530), .Z(n4529) );
  NANDN U5358 ( .A(A[197]), .B(n1786), .Z(n4530) );
  NANDN U5359 ( .A(n1786), .B(A[197]), .Z(n4528) );
  AND U5360 ( .A(n4531), .B(n4532), .Z(n1786) );
  NANDN U5361 ( .A(B[196]), .B(n4533), .Z(n4532) );
  NANDN U5362 ( .A(A[196]), .B(n1788), .Z(n4533) );
  NANDN U5363 ( .A(n1788), .B(A[196]), .Z(n4531) );
  AND U5364 ( .A(n4534), .B(n4535), .Z(n1788) );
  NANDN U5365 ( .A(B[195]), .B(n4536), .Z(n4535) );
  NANDN U5366 ( .A(A[195]), .B(n1790), .Z(n4536) );
  NANDN U5367 ( .A(n1790), .B(A[195]), .Z(n4534) );
  AND U5368 ( .A(n4537), .B(n4538), .Z(n1790) );
  NANDN U5369 ( .A(B[194]), .B(n4539), .Z(n4538) );
  NANDN U5370 ( .A(A[194]), .B(n1792), .Z(n4539) );
  NANDN U5371 ( .A(n1792), .B(A[194]), .Z(n4537) );
  AND U5372 ( .A(n4540), .B(n4541), .Z(n1792) );
  NANDN U5373 ( .A(B[193]), .B(n4542), .Z(n4541) );
  NANDN U5374 ( .A(A[193]), .B(n1794), .Z(n4542) );
  NANDN U5375 ( .A(n1794), .B(A[193]), .Z(n4540) );
  AND U5376 ( .A(n4543), .B(n4544), .Z(n1794) );
  NANDN U5377 ( .A(B[192]), .B(n4545), .Z(n4544) );
  NANDN U5378 ( .A(A[192]), .B(n1796), .Z(n4545) );
  NANDN U5379 ( .A(n1796), .B(A[192]), .Z(n4543) );
  AND U5380 ( .A(n4546), .B(n4547), .Z(n1796) );
  NANDN U5381 ( .A(B[191]), .B(n4548), .Z(n4547) );
  NANDN U5382 ( .A(A[191]), .B(n1798), .Z(n4548) );
  NANDN U5383 ( .A(n1798), .B(A[191]), .Z(n4546) );
  AND U5384 ( .A(n4549), .B(n4550), .Z(n1798) );
  NANDN U5385 ( .A(B[190]), .B(n4551), .Z(n4550) );
  NANDN U5386 ( .A(A[190]), .B(n1800), .Z(n4551) );
  NANDN U5387 ( .A(n1800), .B(A[190]), .Z(n4549) );
  AND U5388 ( .A(n4552), .B(n4553), .Z(n1800) );
  NANDN U5389 ( .A(B[189]), .B(n4554), .Z(n4553) );
  NANDN U5390 ( .A(A[189]), .B(n1804), .Z(n4554) );
  NANDN U5391 ( .A(n1804), .B(A[189]), .Z(n4552) );
  AND U5392 ( .A(n4555), .B(n4556), .Z(n1804) );
  NANDN U5393 ( .A(B[188]), .B(n4557), .Z(n4556) );
  NANDN U5394 ( .A(A[188]), .B(n1806), .Z(n4557) );
  NANDN U5395 ( .A(n1806), .B(A[188]), .Z(n4555) );
  AND U5396 ( .A(n4558), .B(n4559), .Z(n1806) );
  NANDN U5397 ( .A(B[187]), .B(n4560), .Z(n4559) );
  NANDN U5398 ( .A(A[187]), .B(n1808), .Z(n4560) );
  NANDN U5399 ( .A(n1808), .B(A[187]), .Z(n4558) );
  AND U5400 ( .A(n4561), .B(n4562), .Z(n1808) );
  NANDN U5401 ( .A(B[186]), .B(n4563), .Z(n4562) );
  NANDN U5402 ( .A(A[186]), .B(n1810), .Z(n4563) );
  NANDN U5403 ( .A(n1810), .B(A[186]), .Z(n4561) );
  AND U5404 ( .A(n4564), .B(n4565), .Z(n1810) );
  NANDN U5405 ( .A(B[185]), .B(n4566), .Z(n4565) );
  NANDN U5406 ( .A(A[185]), .B(n1812), .Z(n4566) );
  NANDN U5407 ( .A(n1812), .B(A[185]), .Z(n4564) );
  AND U5408 ( .A(n4567), .B(n4568), .Z(n1812) );
  NANDN U5409 ( .A(B[184]), .B(n4569), .Z(n4568) );
  NANDN U5410 ( .A(A[184]), .B(n1814), .Z(n4569) );
  NANDN U5411 ( .A(n1814), .B(A[184]), .Z(n4567) );
  AND U5412 ( .A(n4570), .B(n4571), .Z(n1814) );
  NANDN U5413 ( .A(B[183]), .B(n4572), .Z(n4571) );
  NANDN U5414 ( .A(A[183]), .B(n1816), .Z(n4572) );
  NANDN U5415 ( .A(n1816), .B(A[183]), .Z(n4570) );
  AND U5416 ( .A(n4573), .B(n4574), .Z(n1816) );
  NANDN U5417 ( .A(B[182]), .B(n4575), .Z(n4574) );
  NANDN U5418 ( .A(A[182]), .B(n1818), .Z(n4575) );
  NANDN U5419 ( .A(n1818), .B(A[182]), .Z(n4573) );
  AND U5420 ( .A(n4576), .B(n4577), .Z(n1818) );
  NANDN U5421 ( .A(B[181]), .B(n4578), .Z(n4577) );
  NANDN U5422 ( .A(A[181]), .B(n1820), .Z(n4578) );
  NANDN U5423 ( .A(n1820), .B(A[181]), .Z(n4576) );
  AND U5424 ( .A(n4579), .B(n4580), .Z(n1820) );
  NANDN U5425 ( .A(B[180]), .B(n4581), .Z(n4580) );
  NANDN U5426 ( .A(A[180]), .B(n1822), .Z(n4581) );
  NANDN U5427 ( .A(n1822), .B(A[180]), .Z(n4579) );
  AND U5428 ( .A(n4582), .B(n4583), .Z(n1822) );
  NANDN U5429 ( .A(B[179]), .B(n4584), .Z(n4583) );
  NANDN U5430 ( .A(A[179]), .B(n1826), .Z(n4584) );
  NANDN U5431 ( .A(n1826), .B(A[179]), .Z(n4582) );
  AND U5432 ( .A(n4585), .B(n4586), .Z(n1826) );
  NANDN U5433 ( .A(B[178]), .B(n4587), .Z(n4586) );
  NANDN U5434 ( .A(A[178]), .B(n1828), .Z(n4587) );
  NANDN U5435 ( .A(n1828), .B(A[178]), .Z(n4585) );
  AND U5436 ( .A(n4588), .B(n4589), .Z(n1828) );
  NANDN U5437 ( .A(B[177]), .B(n4590), .Z(n4589) );
  NANDN U5438 ( .A(A[177]), .B(n1830), .Z(n4590) );
  NANDN U5439 ( .A(n1830), .B(A[177]), .Z(n4588) );
  AND U5440 ( .A(n4591), .B(n4592), .Z(n1830) );
  NANDN U5441 ( .A(B[176]), .B(n4593), .Z(n4592) );
  NANDN U5442 ( .A(A[176]), .B(n1832), .Z(n4593) );
  NANDN U5443 ( .A(n1832), .B(A[176]), .Z(n4591) );
  AND U5444 ( .A(n4594), .B(n4595), .Z(n1832) );
  NANDN U5445 ( .A(B[175]), .B(n4596), .Z(n4595) );
  NANDN U5446 ( .A(A[175]), .B(n1834), .Z(n4596) );
  NANDN U5447 ( .A(n1834), .B(A[175]), .Z(n4594) );
  AND U5448 ( .A(n4597), .B(n4598), .Z(n1834) );
  NANDN U5449 ( .A(B[174]), .B(n4599), .Z(n4598) );
  NANDN U5450 ( .A(A[174]), .B(n1836), .Z(n4599) );
  NANDN U5451 ( .A(n1836), .B(A[174]), .Z(n4597) );
  AND U5452 ( .A(n4600), .B(n4601), .Z(n1836) );
  NANDN U5453 ( .A(B[173]), .B(n4602), .Z(n4601) );
  NANDN U5454 ( .A(A[173]), .B(n1838), .Z(n4602) );
  NANDN U5455 ( .A(n1838), .B(A[173]), .Z(n4600) );
  AND U5456 ( .A(n4603), .B(n4604), .Z(n1838) );
  NANDN U5457 ( .A(B[172]), .B(n4605), .Z(n4604) );
  NANDN U5458 ( .A(A[172]), .B(n1840), .Z(n4605) );
  NANDN U5459 ( .A(n1840), .B(A[172]), .Z(n4603) );
  AND U5460 ( .A(n4606), .B(n4607), .Z(n1840) );
  NANDN U5461 ( .A(B[171]), .B(n4608), .Z(n4607) );
  NANDN U5462 ( .A(A[171]), .B(n1842), .Z(n4608) );
  NANDN U5463 ( .A(n1842), .B(A[171]), .Z(n4606) );
  AND U5464 ( .A(n4609), .B(n4610), .Z(n1842) );
  NANDN U5465 ( .A(B[170]), .B(n4611), .Z(n4610) );
  NANDN U5466 ( .A(A[170]), .B(n1844), .Z(n4611) );
  NANDN U5467 ( .A(n1844), .B(A[170]), .Z(n4609) );
  AND U5468 ( .A(n4612), .B(n4613), .Z(n1844) );
  NANDN U5469 ( .A(B[169]), .B(n4614), .Z(n4613) );
  NANDN U5470 ( .A(A[169]), .B(n1848), .Z(n4614) );
  NANDN U5471 ( .A(n1848), .B(A[169]), .Z(n4612) );
  AND U5472 ( .A(n4615), .B(n4616), .Z(n1848) );
  NANDN U5473 ( .A(B[168]), .B(n4617), .Z(n4616) );
  NANDN U5474 ( .A(A[168]), .B(n1850), .Z(n4617) );
  NANDN U5475 ( .A(n1850), .B(A[168]), .Z(n4615) );
  AND U5476 ( .A(n4618), .B(n4619), .Z(n1850) );
  NANDN U5477 ( .A(B[167]), .B(n4620), .Z(n4619) );
  NANDN U5478 ( .A(A[167]), .B(n1852), .Z(n4620) );
  NANDN U5479 ( .A(n1852), .B(A[167]), .Z(n4618) );
  AND U5480 ( .A(n4621), .B(n4622), .Z(n1852) );
  NANDN U5481 ( .A(B[166]), .B(n4623), .Z(n4622) );
  NANDN U5482 ( .A(A[166]), .B(n1854), .Z(n4623) );
  NANDN U5483 ( .A(n1854), .B(A[166]), .Z(n4621) );
  AND U5484 ( .A(n4624), .B(n4625), .Z(n1854) );
  NANDN U5485 ( .A(B[165]), .B(n4626), .Z(n4625) );
  NANDN U5486 ( .A(A[165]), .B(n1856), .Z(n4626) );
  NANDN U5487 ( .A(n1856), .B(A[165]), .Z(n4624) );
  AND U5488 ( .A(n4627), .B(n4628), .Z(n1856) );
  NANDN U5489 ( .A(B[164]), .B(n4629), .Z(n4628) );
  NANDN U5490 ( .A(A[164]), .B(n1858), .Z(n4629) );
  NANDN U5491 ( .A(n1858), .B(A[164]), .Z(n4627) );
  AND U5492 ( .A(n4630), .B(n4631), .Z(n1858) );
  NANDN U5493 ( .A(B[163]), .B(n4632), .Z(n4631) );
  NANDN U5494 ( .A(A[163]), .B(n1860), .Z(n4632) );
  NANDN U5495 ( .A(n1860), .B(A[163]), .Z(n4630) );
  AND U5496 ( .A(n4633), .B(n4634), .Z(n1860) );
  NANDN U5497 ( .A(B[162]), .B(n4635), .Z(n4634) );
  NANDN U5498 ( .A(A[162]), .B(n1862), .Z(n4635) );
  NANDN U5499 ( .A(n1862), .B(A[162]), .Z(n4633) );
  AND U5500 ( .A(n4636), .B(n4637), .Z(n1862) );
  NANDN U5501 ( .A(B[161]), .B(n4638), .Z(n4637) );
  NANDN U5502 ( .A(A[161]), .B(n1864), .Z(n4638) );
  NANDN U5503 ( .A(n1864), .B(A[161]), .Z(n4636) );
  AND U5504 ( .A(n4639), .B(n4640), .Z(n1864) );
  NANDN U5505 ( .A(B[160]), .B(n4641), .Z(n4640) );
  NANDN U5506 ( .A(A[160]), .B(n1866), .Z(n4641) );
  NANDN U5507 ( .A(n1866), .B(A[160]), .Z(n4639) );
  AND U5508 ( .A(n4642), .B(n4643), .Z(n1866) );
  NANDN U5509 ( .A(B[159]), .B(n4644), .Z(n4643) );
  NANDN U5510 ( .A(A[159]), .B(n1870), .Z(n4644) );
  NANDN U5511 ( .A(n1870), .B(A[159]), .Z(n4642) );
  AND U5512 ( .A(n4645), .B(n4646), .Z(n1870) );
  NANDN U5513 ( .A(B[158]), .B(n4647), .Z(n4646) );
  NANDN U5514 ( .A(A[158]), .B(n1872), .Z(n4647) );
  NANDN U5515 ( .A(n1872), .B(A[158]), .Z(n4645) );
  AND U5516 ( .A(n4648), .B(n4649), .Z(n1872) );
  NANDN U5517 ( .A(B[157]), .B(n4650), .Z(n4649) );
  NANDN U5518 ( .A(A[157]), .B(n1874), .Z(n4650) );
  NANDN U5519 ( .A(n1874), .B(A[157]), .Z(n4648) );
  AND U5520 ( .A(n4651), .B(n4652), .Z(n1874) );
  NANDN U5521 ( .A(B[156]), .B(n4653), .Z(n4652) );
  NANDN U5522 ( .A(A[156]), .B(n1876), .Z(n4653) );
  NANDN U5523 ( .A(n1876), .B(A[156]), .Z(n4651) );
  AND U5524 ( .A(n4654), .B(n4655), .Z(n1876) );
  NANDN U5525 ( .A(B[155]), .B(n4656), .Z(n4655) );
  NANDN U5526 ( .A(A[155]), .B(n1878), .Z(n4656) );
  NANDN U5527 ( .A(n1878), .B(A[155]), .Z(n4654) );
  AND U5528 ( .A(n4657), .B(n4658), .Z(n1878) );
  NANDN U5529 ( .A(B[154]), .B(n4659), .Z(n4658) );
  NANDN U5530 ( .A(A[154]), .B(n1880), .Z(n4659) );
  NANDN U5531 ( .A(n1880), .B(A[154]), .Z(n4657) );
  AND U5532 ( .A(n4660), .B(n4661), .Z(n1880) );
  NANDN U5533 ( .A(B[153]), .B(n4662), .Z(n4661) );
  NANDN U5534 ( .A(A[153]), .B(n1882), .Z(n4662) );
  NANDN U5535 ( .A(n1882), .B(A[153]), .Z(n4660) );
  AND U5536 ( .A(n4663), .B(n4664), .Z(n1882) );
  NANDN U5537 ( .A(B[152]), .B(n4665), .Z(n4664) );
  NANDN U5538 ( .A(A[152]), .B(n1884), .Z(n4665) );
  NANDN U5539 ( .A(n1884), .B(A[152]), .Z(n4663) );
  AND U5540 ( .A(n4666), .B(n4667), .Z(n1884) );
  NANDN U5541 ( .A(B[151]), .B(n4668), .Z(n4667) );
  NANDN U5542 ( .A(A[151]), .B(n1886), .Z(n4668) );
  NANDN U5543 ( .A(n1886), .B(A[151]), .Z(n4666) );
  AND U5544 ( .A(n4669), .B(n4670), .Z(n1886) );
  NANDN U5545 ( .A(B[150]), .B(n4671), .Z(n4670) );
  NANDN U5546 ( .A(A[150]), .B(n1888), .Z(n4671) );
  NANDN U5547 ( .A(n1888), .B(A[150]), .Z(n4669) );
  AND U5548 ( .A(n4672), .B(n4673), .Z(n1888) );
  NANDN U5549 ( .A(B[149]), .B(n4674), .Z(n4673) );
  NANDN U5550 ( .A(A[149]), .B(n1892), .Z(n4674) );
  NANDN U5551 ( .A(n1892), .B(A[149]), .Z(n4672) );
  AND U5552 ( .A(n4675), .B(n4676), .Z(n1892) );
  NANDN U5553 ( .A(B[148]), .B(n4677), .Z(n4676) );
  NANDN U5554 ( .A(A[148]), .B(n1894), .Z(n4677) );
  NANDN U5555 ( .A(n1894), .B(A[148]), .Z(n4675) );
  AND U5556 ( .A(n4678), .B(n4679), .Z(n1894) );
  NANDN U5557 ( .A(B[147]), .B(n4680), .Z(n4679) );
  NANDN U5558 ( .A(A[147]), .B(n1896), .Z(n4680) );
  NANDN U5559 ( .A(n1896), .B(A[147]), .Z(n4678) );
  AND U5560 ( .A(n4681), .B(n4682), .Z(n1896) );
  NANDN U5561 ( .A(B[146]), .B(n4683), .Z(n4682) );
  NANDN U5562 ( .A(A[146]), .B(n1898), .Z(n4683) );
  NANDN U5563 ( .A(n1898), .B(A[146]), .Z(n4681) );
  AND U5564 ( .A(n4684), .B(n4685), .Z(n1898) );
  NANDN U5565 ( .A(B[145]), .B(n4686), .Z(n4685) );
  NANDN U5566 ( .A(A[145]), .B(n1900), .Z(n4686) );
  NANDN U5567 ( .A(n1900), .B(A[145]), .Z(n4684) );
  AND U5568 ( .A(n4687), .B(n4688), .Z(n1900) );
  NANDN U5569 ( .A(B[144]), .B(n4689), .Z(n4688) );
  NANDN U5570 ( .A(A[144]), .B(n1902), .Z(n4689) );
  NANDN U5571 ( .A(n1902), .B(A[144]), .Z(n4687) );
  AND U5572 ( .A(n4690), .B(n4691), .Z(n1902) );
  NANDN U5573 ( .A(B[143]), .B(n4692), .Z(n4691) );
  NANDN U5574 ( .A(A[143]), .B(n1904), .Z(n4692) );
  NANDN U5575 ( .A(n1904), .B(A[143]), .Z(n4690) );
  AND U5576 ( .A(n4693), .B(n4694), .Z(n1904) );
  NANDN U5577 ( .A(B[142]), .B(n4695), .Z(n4694) );
  NANDN U5578 ( .A(A[142]), .B(n1906), .Z(n4695) );
  NANDN U5579 ( .A(n1906), .B(A[142]), .Z(n4693) );
  AND U5580 ( .A(n4696), .B(n4697), .Z(n1906) );
  NANDN U5581 ( .A(B[141]), .B(n4698), .Z(n4697) );
  NANDN U5582 ( .A(A[141]), .B(n1908), .Z(n4698) );
  NANDN U5583 ( .A(n1908), .B(A[141]), .Z(n4696) );
  AND U5584 ( .A(n4699), .B(n4700), .Z(n1908) );
  NANDN U5585 ( .A(B[140]), .B(n4701), .Z(n4700) );
  NANDN U5586 ( .A(A[140]), .B(n1910), .Z(n4701) );
  NANDN U5587 ( .A(n1910), .B(A[140]), .Z(n4699) );
  AND U5588 ( .A(n4702), .B(n4703), .Z(n1910) );
  NANDN U5589 ( .A(B[139]), .B(n4704), .Z(n4703) );
  NANDN U5590 ( .A(A[139]), .B(n1914), .Z(n4704) );
  NANDN U5591 ( .A(n1914), .B(A[139]), .Z(n4702) );
  AND U5592 ( .A(n4705), .B(n4706), .Z(n1914) );
  NANDN U5593 ( .A(B[138]), .B(n4707), .Z(n4706) );
  NANDN U5594 ( .A(A[138]), .B(n1916), .Z(n4707) );
  NANDN U5595 ( .A(n1916), .B(A[138]), .Z(n4705) );
  AND U5596 ( .A(n4708), .B(n4709), .Z(n1916) );
  NANDN U5597 ( .A(B[137]), .B(n4710), .Z(n4709) );
  NANDN U5598 ( .A(A[137]), .B(n1918), .Z(n4710) );
  NANDN U5599 ( .A(n1918), .B(A[137]), .Z(n4708) );
  AND U5600 ( .A(n4711), .B(n4712), .Z(n1918) );
  NANDN U5601 ( .A(B[136]), .B(n4713), .Z(n4712) );
  NANDN U5602 ( .A(A[136]), .B(n1920), .Z(n4713) );
  NANDN U5603 ( .A(n1920), .B(A[136]), .Z(n4711) );
  AND U5604 ( .A(n4714), .B(n4715), .Z(n1920) );
  NANDN U5605 ( .A(B[135]), .B(n4716), .Z(n4715) );
  NANDN U5606 ( .A(A[135]), .B(n1922), .Z(n4716) );
  NANDN U5607 ( .A(n1922), .B(A[135]), .Z(n4714) );
  AND U5608 ( .A(n4717), .B(n4718), .Z(n1922) );
  NANDN U5609 ( .A(B[134]), .B(n4719), .Z(n4718) );
  NANDN U5610 ( .A(A[134]), .B(n1924), .Z(n4719) );
  NANDN U5611 ( .A(n1924), .B(A[134]), .Z(n4717) );
  AND U5612 ( .A(n4720), .B(n4721), .Z(n1924) );
  NANDN U5613 ( .A(B[133]), .B(n4722), .Z(n4721) );
  NANDN U5614 ( .A(A[133]), .B(n1926), .Z(n4722) );
  NANDN U5615 ( .A(n1926), .B(A[133]), .Z(n4720) );
  AND U5616 ( .A(n4723), .B(n4724), .Z(n1926) );
  NANDN U5617 ( .A(B[132]), .B(n4725), .Z(n4724) );
  NANDN U5618 ( .A(A[132]), .B(n1928), .Z(n4725) );
  NANDN U5619 ( .A(n1928), .B(A[132]), .Z(n4723) );
  AND U5620 ( .A(n4726), .B(n4727), .Z(n1928) );
  NANDN U5621 ( .A(B[131]), .B(n4728), .Z(n4727) );
  NANDN U5622 ( .A(A[131]), .B(n1930), .Z(n4728) );
  NANDN U5623 ( .A(n1930), .B(A[131]), .Z(n4726) );
  AND U5624 ( .A(n4729), .B(n4730), .Z(n1930) );
  NANDN U5625 ( .A(B[130]), .B(n4731), .Z(n4730) );
  NANDN U5626 ( .A(A[130]), .B(n1932), .Z(n4731) );
  NANDN U5627 ( .A(n1932), .B(A[130]), .Z(n4729) );
  AND U5628 ( .A(n4732), .B(n4733), .Z(n1932) );
  NANDN U5629 ( .A(B[129]), .B(n4734), .Z(n4733) );
  NANDN U5630 ( .A(A[129]), .B(n1936), .Z(n4734) );
  NANDN U5631 ( .A(n1936), .B(A[129]), .Z(n4732) );
  AND U5632 ( .A(n4735), .B(n4736), .Z(n1936) );
  NANDN U5633 ( .A(B[128]), .B(n4737), .Z(n4736) );
  NANDN U5634 ( .A(A[128]), .B(n1938), .Z(n4737) );
  NANDN U5635 ( .A(n1938), .B(A[128]), .Z(n4735) );
  AND U5636 ( .A(n4738), .B(n4739), .Z(n1938) );
  NANDN U5637 ( .A(B[127]), .B(n4740), .Z(n4739) );
  NANDN U5638 ( .A(A[127]), .B(n1940), .Z(n4740) );
  NANDN U5639 ( .A(n1940), .B(A[127]), .Z(n4738) );
  AND U5640 ( .A(n4741), .B(n4742), .Z(n1940) );
  NANDN U5641 ( .A(B[126]), .B(n4743), .Z(n4742) );
  NANDN U5642 ( .A(A[126]), .B(n1942), .Z(n4743) );
  NANDN U5643 ( .A(n1942), .B(A[126]), .Z(n4741) );
  AND U5644 ( .A(n4744), .B(n4745), .Z(n1942) );
  NANDN U5645 ( .A(B[125]), .B(n4746), .Z(n4745) );
  NANDN U5646 ( .A(A[125]), .B(n1944), .Z(n4746) );
  NANDN U5647 ( .A(n1944), .B(A[125]), .Z(n4744) );
  AND U5648 ( .A(n4747), .B(n4748), .Z(n1944) );
  NANDN U5649 ( .A(B[124]), .B(n4749), .Z(n4748) );
  NANDN U5650 ( .A(A[124]), .B(n1946), .Z(n4749) );
  NANDN U5651 ( .A(n1946), .B(A[124]), .Z(n4747) );
  AND U5652 ( .A(n4750), .B(n4751), .Z(n1946) );
  NANDN U5653 ( .A(B[123]), .B(n4752), .Z(n4751) );
  NANDN U5654 ( .A(A[123]), .B(n1948), .Z(n4752) );
  NANDN U5655 ( .A(n1948), .B(A[123]), .Z(n4750) );
  AND U5656 ( .A(n4753), .B(n4754), .Z(n1948) );
  NANDN U5657 ( .A(B[122]), .B(n4755), .Z(n4754) );
  NANDN U5658 ( .A(A[122]), .B(n1950), .Z(n4755) );
  NANDN U5659 ( .A(n1950), .B(A[122]), .Z(n4753) );
  AND U5660 ( .A(n4756), .B(n4757), .Z(n1950) );
  NANDN U5661 ( .A(B[121]), .B(n4758), .Z(n4757) );
  NANDN U5662 ( .A(A[121]), .B(n1952), .Z(n4758) );
  NANDN U5663 ( .A(n1952), .B(A[121]), .Z(n4756) );
  AND U5664 ( .A(n4759), .B(n4760), .Z(n1952) );
  NANDN U5665 ( .A(B[120]), .B(n4761), .Z(n4760) );
  NANDN U5666 ( .A(A[120]), .B(n1954), .Z(n4761) );
  NANDN U5667 ( .A(n1954), .B(A[120]), .Z(n4759) );
  AND U5668 ( .A(n4762), .B(n4763), .Z(n1954) );
  NANDN U5669 ( .A(B[119]), .B(n4764), .Z(n4763) );
  NANDN U5670 ( .A(A[119]), .B(n1958), .Z(n4764) );
  NANDN U5671 ( .A(n1958), .B(A[119]), .Z(n4762) );
  AND U5672 ( .A(n4765), .B(n4766), .Z(n1958) );
  NANDN U5673 ( .A(B[118]), .B(n4767), .Z(n4766) );
  NANDN U5674 ( .A(A[118]), .B(n1960), .Z(n4767) );
  NANDN U5675 ( .A(n1960), .B(A[118]), .Z(n4765) );
  AND U5676 ( .A(n4768), .B(n4769), .Z(n1960) );
  NANDN U5677 ( .A(B[117]), .B(n4770), .Z(n4769) );
  NANDN U5678 ( .A(A[117]), .B(n1962), .Z(n4770) );
  NANDN U5679 ( .A(n1962), .B(A[117]), .Z(n4768) );
  AND U5680 ( .A(n4771), .B(n4772), .Z(n1962) );
  NANDN U5681 ( .A(B[116]), .B(n4773), .Z(n4772) );
  NANDN U5682 ( .A(A[116]), .B(n1964), .Z(n4773) );
  NANDN U5683 ( .A(n1964), .B(A[116]), .Z(n4771) );
  AND U5684 ( .A(n4774), .B(n4775), .Z(n1964) );
  NANDN U5685 ( .A(B[115]), .B(n4776), .Z(n4775) );
  NANDN U5686 ( .A(A[115]), .B(n1966), .Z(n4776) );
  NANDN U5687 ( .A(n1966), .B(A[115]), .Z(n4774) );
  AND U5688 ( .A(n4777), .B(n4778), .Z(n1966) );
  NANDN U5689 ( .A(B[114]), .B(n4779), .Z(n4778) );
  NANDN U5690 ( .A(A[114]), .B(n1968), .Z(n4779) );
  NANDN U5691 ( .A(n1968), .B(A[114]), .Z(n4777) );
  AND U5692 ( .A(n4780), .B(n4781), .Z(n1968) );
  NANDN U5693 ( .A(B[113]), .B(n4782), .Z(n4781) );
  NANDN U5694 ( .A(A[113]), .B(n1970), .Z(n4782) );
  NANDN U5695 ( .A(n1970), .B(A[113]), .Z(n4780) );
  AND U5696 ( .A(n4783), .B(n4784), .Z(n1970) );
  NANDN U5697 ( .A(B[112]), .B(n4785), .Z(n4784) );
  NANDN U5698 ( .A(A[112]), .B(n1972), .Z(n4785) );
  NANDN U5699 ( .A(n1972), .B(A[112]), .Z(n4783) );
  AND U5700 ( .A(n4786), .B(n4787), .Z(n1972) );
  NANDN U5701 ( .A(B[111]), .B(n4788), .Z(n4787) );
  NANDN U5702 ( .A(A[111]), .B(n1974), .Z(n4788) );
  NANDN U5703 ( .A(n1974), .B(A[111]), .Z(n4786) );
  AND U5704 ( .A(n4789), .B(n4790), .Z(n1974) );
  NANDN U5705 ( .A(B[110]), .B(n4791), .Z(n4790) );
  NANDN U5706 ( .A(A[110]), .B(n1976), .Z(n4791) );
  NANDN U5707 ( .A(n1976), .B(A[110]), .Z(n4789) );
  AND U5708 ( .A(n4792), .B(n4793), .Z(n1976) );
  NANDN U5709 ( .A(B[109]), .B(n4794), .Z(n4793) );
  NANDN U5710 ( .A(A[109]), .B(n1980), .Z(n4794) );
  NANDN U5711 ( .A(n1980), .B(A[109]), .Z(n4792) );
  AND U5712 ( .A(n4795), .B(n4796), .Z(n1980) );
  NANDN U5713 ( .A(B[108]), .B(n4797), .Z(n4796) );
  NANDN U5714 ( .A(A[108]), .B(n1982), .Z(n4797) );
  NANDN U5715 ( .A(n1982), .B(A[108]), .Z(n4795) );
  AND U5716 ( .A(n4798), .B(n4799), .Z(n1982) );
  NANDN U5717 ( .A(B[107]), .B(n4800), .Z(n4799) );
  NANDN U5718 ( .A(A[107]), .B(n1984), .Z(n4800) );
  NANDN U5719 ( .A(n1984), .B(A[107]), .Z(n4798) );
  AND U5720 ( .A(n4801), .B(n4802), .Z(n1984) );
  NANDN U5721 ( .A(B[106]), .B(n4803), .Z(n4802) );
  NANDN U5722 ( .A(A[106]), .B(n1986), .Z(n4803) );
  NANDN U5723 ( .A(n1986), .B(A[106]), .Z(n4801) );
  AND U5724 ( .A(n4804), .B(n4805), .Z(n1986) );
  NANDN U5725 ( .A(B[105]), .B(n4806), .Z(n4805) );
  NANDN U5726 ( .A(A[105]), .B(n1988), .Z(n4806) );
  NANDN U5727 ( .A(n1988), .B(A[105]), .Z(n4804) );
  AND U5728 ( .A(n4807), .B(n4808), .Z(n1988) );
  NANDN U5729 ( .A(B[104]), .B(n4809), .Z(n4808) );
  NANDN U5730 ( .A(A[104]), .B(n1990), .Z(n4809) );
  NANDN U5731 ( .A(n1990), .B(A[104]), .Z(n4807) );
  AND U5732 ( .A(n4810), .B(n4811), .Z(n1990) );
  NANDN U5733 ( .A(B[103]), .B(n4812), .Z(n4811) );
  NANDN U5734 ( .A(A[103]), .B(n1992), .Z(n4812) );
  NANDN U5735 ( .A(n1992), .B(A[103]), .Z(n4810) );
  AND U5736 ( .A(n4813), .B(n4814), .Z(n1992) );
  NANDN U5737 ( .A(B[102]), .B(n4815), .Z(n4814) );
  NANDN U5738 ( .A(A[102]), .B(n1994), .Z(n4815) );
  NANDN U5739 ( .A(n1994), .B(A[102]), .Z(n4813) );
  AND U5740 ( .A(n4816), .B(n4817), .Z(n1994) );
  NANDN U5741 ( .A(B[101]), .B(n4818), .Z(n4817) );
  NANDN U5742 ( .A(A[101]), .B(n2022), .Z(n4818) );
  NANDN U5743 ( .A(n2022), .B(A[101]), .Z(n4816) );
  AND U5744 ( .A(n4819), .B(n4820), .Z(n2022) );
  NANDN U5745 ( .A(B[100]), .B(n4821), .Z(n4820) );
  NANDN U5746 ( .A(A[100]), .B(n2074), .Z(n4821) );
  NANDN U5747 ( .A(n2074), .B(A[100]), .Z(n4819) );
  AND U5748 ( .A(n4822), .B(n4823), .Z(n2074) );
  NANDN U5749 ( .A(B[99]), .B(n4824), .Z(n4823) );
  OR U5750 ( .A(n5), .B(A[99]), .Z(n4824) );
  NAND U5751 ( .A(A[99]), .B(n5), .Z(n4822) );
  NAND U5752 ( .A(n4825), .B(n4826), .Z(n5) );
  NANDN U5753 ( .A(B[98]), .B(n4827), .Z(n4826) );
  NANDN U5754 ( .A(A[98]), .B(n27), .Z(n4827) );
  NANDN U5755 ( .A(n27), .B(A[98]), .Z(n4825) );
  AND U5756 ( .A(n4828), .B(n4829), .Z(n27) );
  NANDN U5757 ( .A(B[97]), .B(n4830), .Z(n4829) );
  NANDN U5758 ( .A(A[97]), .B(n49), .Z(n4830) );
  NANDN U5759 ( .A(n49), .B(A[97]), .Z(n4828) );
  AND U5760 ( .A(n4831), .B(n4832), .Z(n49) );
  NANDN U5761 ( .A(B[96]), .B(n4833), .Z(n4832) );
  NANDN U5762 ( .A(A[96]), .B(n71), .Z(n4833) );
  NANDN U5763 ( .A(n71), .B(A[96]), .Z(n4831) );
  AND U5764 ( .A(n4834), .B(n4835), .Z(n71) );
  NANDN U5765 ( .A(B[95]), .B(n4836), .Z(n4835) );
  NANDN U5766 ( .A(A[95]), .B(n93), .Z(n4836) );
  NANDN U5767 ( .A(n93), .B(A[95]), .Z(n4834) );
  AND U5768 ( .A(n4837), .B(n4838), .Z(n93) );
  NANDN U5769 ( .A(B[94]), .B(n4839), .Z(n4838) );
  NANDN U5770 ( .A(A[94]), .B(n115), .Z(n4839) );
  NANDN U5771 ( .A(n115), .B(A[94]), .Z(n4837) );
  AND U5772 ( .A(n4840), .B(n4841), .Z(n115) );
  NANDN U5773 ( .A(B[93]), .B(n4842), .Z(n4841) );
  NANDN U5774 ( .A(A[93]), .B(n137), .Z(n4842) );
  NANDN U5775 ( .A(n137), .B(A[93]), .Z(n4840) );
  AND U5776 ( .A(n4843), .B(n4844), .Z(n137) );
  NANDN U5777 ( .A(B[92]), .B(n4845), .Z(n4844) );
  NANDN U5778 ( .A(A[92]), .B(n159), .Z(n4845) );
  NANDN U5779 ( .A(n159), .B(A[92]), .Z(n4843) );
  AND U5780 ( .A(n4846), .B(n4847), .Z(n159) );
  NANDN U5781 ( .A(B[91]), .B(n4848), .Z(n4847) );
  NANDN U5782 ( .A(A[91]), .B(n181), .Z(n4848) );
  NANDN U5783 ( .A(n181), .B(A[91]), .Z(n4846) );
  AND U5784 ( .A(n4849), .B(n4850), .Z(n181) );
  NANDN U5785 ( .A(B[90]), .B(n4851), .Z(n4850) );
  NANDN U5786 ( .A(A[90]), .B(n203), .Z(n4851) );
  NANDN U5787 ( .A(n203), .B(A[90]), .Z(n4849) );
  AND U5788 ( .A(n4852), .B(n4853), .Z(n203) );
  NANDN U5789 ( .A(B[89]), .B(n4854), .Z(n4853) );
  NANDN U5790 ( .A(A[89]), .B(n227), .Z(n4854) );
  NANDN U5791 ( .A(n227), .B(A[89]), .Z(n4852) );
  AND U5792 ( .A(n4855), .B(n4856), .Z(n227) );
  NANDN U5793 ( .A(B[88]), .B(n4857), .Z(n4856) );
  NANDN U5794 ( .A(A[88]), .B(n249), .Z(n4857) );
  NANDN U5795 ( .A(n249), .B(A[88]), .Z(n4855) );
  AND U5796 ( .A(n4858), .B(n4859), .Z(n249) );
  NANDN U5797 ( .A(B[87]), .B(n4860), .Z(n4859) );
  NANDN U5798 ( .A(A[87]), .B(n271), .Z(n4860) );
  NANDN U5799 ( .A(n271), .B(A[87]), .Z(n4858) );
  AND U5800 ( .A(n4861), .B(n4862), .Z(n271) );
  NANDN U5801 ( .A(B[86]), .B(n4863), .Z(n4862) );
  NANDN U5802 ( .A(A[86]), .B(n293), .Z(n4863) );
  NANDN U5803 ( .A(n293), .B(A[86]), .Z(n4861) );
  AND U5804 ( .A(n4864), .B(n4865), .Z(n293) );
  NANDN U5805 ( .A(B[85]), .B(n4866), .Z(n4865) );
  NANDN U5806 ( .A(A[85]), .B(n315), .Z(n4866) );
  NANDN U5807 ( .A(n315), .B(A[85]), .Z(n4864) );
  AND U5808 ( .A(n4867), .B(n4868), .Z(n315) );
  NANDN U5809 ( .A(B[84]), .B(n4869), .Z(n4868) );
  NANDN U5810 ( .A(A[84]), .B(n337), .Z(n4869) );
  NANDN U5811 ( .A(n337), .B(A[84]), .Z(n4867) );
  AND U5812 ( .A(n4870), .B(n4871), .Z(n337) );
  NANDN U5813 ( .A(B[83]), .B(n4872), .Z(n4871) );
  NANDN U5814 ( .A(A[83]), .B(n359), .Z(n4872) );
  NANDN U5815 ( .A(n359), .B(A[83]), .Z(n4870) );
  AND U5816 ( .A(n4873), .B(n4874), .Z(n359) );
  NANDN U5817 ( .A(B[82]), .B(n4875), .Z(n4874) );
  NANDN U5818 ( .A(A[82]), .B(n381), .Z(n4875) );
  NANDN U5819 ( .A(n381), .B(A[82]), .Z(n4873) );
  AND U5820 ( .A(n4876), .B(n4877), .Z(n381) );
  NANDN U5821 ( .A(B[81]), .B(n4878), .Z(n4877) );
  NANDN U5822 ( .A(A[81]), .B(n403), .Z(n4878) );
  NANDN U5823 ( .A(n403), .B(A[81]), .Z(n4876) );
  AND U5824 ( .A(n4879), .B(n4880), .Z(n403) );
  NANDN U5825 ( .A(B[80]), .B(n4881), .Z(n4880) );
  NANDN U5826 ( .A(A[80]), .B(n425), .Z(n4881) );
  NANDN U5827 ( .A(n425), .B(A[80]), .Z(n4879) );
  AND U5828 ( .A(n4882), .B(n4883), .Z(n425) );
  NANDN U5829 ( .A(B[79]), .B(n4884), .Z(n4883) );
  NANDN U5830 ( .A(A[79]), .B(n449), .Z(n4884) );
  NANDN U5831 ( .A(n449), .B(A[79]), .Z(n4882) );
  AND U5832 ( .A(n4885), .B(n4886), .Z(n449) );
  NANDN U5833 ( .A(B[78]), .B(n4887), .Z(n4886) );
  NANDN U5834 ( .A(A[78]), .B(n471), .Z(n4887) );
  NANDN U5835 ( .A(n471), .B(A[78]), .Z(n4885) );
  AND U5836 ( .A(n4888), .B(n4889), .Z(n471) );
  NANDN U5837 ( .A(B[77]), .B(n4890), .Z(n4889) );
  NANDN U5838 ( .A(A[77]), .B(n493), .Z(n4890) );
  NANDN U5839 ( .A(n493), .B(A[77]), .Z(n4888) );
  AND U5840 ( .A(n4891), .B(n4892), .Z(n493) );
  NANDN U5841 ( .A(B[76]), .B(n4893), .Z(n4892) );
  NANDN U5842 ( .A(A[76]), .B(n515), .Z(n4893) );
  NANDN U5843 ( .A(n515), .B(A[76]), .Z(n4891) );
  AND U5844 ( .A(n4894), .B(n4895), .Z(n515) );
  NANDN U5845 ( .A(B[75]), .B(n4896), .Z(n4895) );
  NANDN U5846 ( .A(A[75]), .B(n537), .Z(n4896) );
  NANDN U5847 ( .A(n537), .B(A[75]), .Z(n4894) );
  AND U5848 ( .A(n4897), .B(n4898), .Z(n537) );
  NANDN U5849 ( .A(B[74]), .B(n4899), .Z(n4898) );
  NANDN U5850 ( .A(A[74]), .B(n559), .Z(n4899) );
  NANDN U5851 ( .A(n559), .B(A[74]), .Z(n4897) );
  AND U5852 ( .A(n4900), .B(n4901), .Z(n559) );
  NANDN U5853 ( .A(B[73]), .B(n4902), .Z(n4901) );
  NANDN U5854 ( .A(A[73]), .B(n581), .Z(n4902) );
  NANDN U5855 ( .A(n581), .B(A[73]), .Z(n4900) );
  AND U5856 ( .A(n4903), .B(n4904), .Z(n581) );
  NANDN U5857 ( .A(B[72]), .B(n4905), .Z(n4904) );
  NANDN U5858 ( .A(A[72]), .B(n603), .Z(n4905) );
  NANDN U5859 ( .A(n603), .B(A[72]), .Z(n4903) );
  AND U5860 ( .A(n4906), .B(n4907), .Z(n603) );
  NANDN U5861 ( .A(B[71]), .B(n4908), .Z(n4907) );
  NANDN U5862 ( .A(A[71]), .B(n625), .Z(n4908) );
  NANDN U5863 ( .A(n625), .B(A[71]), .Z(n4906) );
  AND U5864 ( .A(n4909), .B(n4910), .Z(n625) );
  NANDN U5865 ( .A(B[70]), .B(n4911), .Z(n4910) );
  NANDN U5866 ( .A(A[70]), .B(n647), .Z(n4911) );
  NANDN U5867 ( .A(n647), .B(A[70]), .Z(n4909) );
  AND U5868 ( .A(n4912), .B(n4913), .Z(n647) );
  NANDN U5869 ( .A(B[69]), .B(n4914), .Z(n4913) );
  NANDN U5870 ( .A(A[69]), .B(n671), .Z(n4914) );
  NANDN U5871 ( .A(n671), .B(A[69]), .Z(n4912) );
  AND U5872 ( .A(n4915), .B(n4916), .Z(n671) );
  NANDN U5873 ( .A(B[68]), .B(n4917), .Z(n4916) );
  NANDN U5874 ( .A(A[68]), .B(n693), .Z(n4917) );
  NANDN U5875 ( .A(n693), .B(A[68]), .Z(n4915) );
  AND U5876 ( .A(n4918), .B(n4919), .Z(n693) );
  NANDN U5877 ( .A(B[67]), .B(n4920), .Z(n4919) );
  NANDN U5878 ( .A(A[67]), .B(n715), .Z(n4920) );
  NANDN U5879 ( .A(n715), .B(A[67]), .Z(n4918) );
  AND U5880 ( .A(n4921), .B(n4922), .Z(n715) );
  NANDN U5881 ( .A(B[66]), .B(n4923), .Z(n4922) );
  NANDN U5882 ( .A(A[66]), .B(n737), .Z(n4923) );
  NANDN U5883 ( .A(n737), .B(A[66]), .Z(n4921) );
  AND U5884 ( .A(n4924), .B(n4925), .Z(n737) );
  NANDN U5885 ( .A(B[65]), .B(n4926), .Z(n4925) );
  NANDN U5886 ( .A(A[65]), .B(n759), .Z(n4926) );
  NANDN U5887 ( .A(n759), .B(A[65]), .Z(n4924) );
  AND U5888 ( .A(n4927), .B(n4928), .Z(n759) );
  NANDN U5889 ( .A(B[64]), .B(n4929), .Z(n4928) );
  NANDN U5890 ( .A(A[64]), .B(n781), .Z(n4929) );
  NANDN U5891 ( .A(n781), .B(A[64]), .Z(n4927) );
  AND U5892 ( .A(n4930), .B(n4931), .Z(n781) );
  NANDN U5893 ( .A(B[63]), .B(n4932), .Z(n4931) );
  NANDN U5894 ( .A(A[63]), .B(n803), .Z(n4932) );
  NANDN U5895 ( .A(n803), .B(A[63]), .Z(n4930) );
  AND U5896 ( .A(n4933), .B(n4934), .Z(n803) );
  NANDN U5897 ( .A(B[62]), .B(n4935), .Z(n4934) );
  NANDN U5898 ( .A(A[62]), .B(n825), .Z(n4935) );
  NANDN U5899 ( .A(n825), .B(A[62]), .Z(n4933) );
  AND U5900 ( .A(n4936), .B(n4937), .Z(n825) );
  NANDN U5901 ( .A(B[61]), .B(n4938), .Z(n4937) );
  NANDN U5902 ( .A(A[61]), .B(n847), .Z(n4938) );
  NANDN U5903 ( .A(n847), .B(A[61]), .Z(n4936) );
  AND U5904 ( .A(n4939), .B(n4940), .Z(n847) );
  NANDN U5905 ( .A(B[60]), .B(n4941), .Z(n4940) );
  NANDN U5906 ( .A(A[60]), .B(n869), .Z(n4941) );
  NANDN U5907 ( .A(n869), .B(A[60]), .Z(n4939) );
  AND U5908 ( .A(n4942), .B(n4943), .Z(n869) );
  NANDN U5909 ( .A(B[59]), .B(n4944), .Z(n4943) );
  NANDN U5910 ( .A(A[59]), .B(n893), .Z(n4944) );
  NANDN U5911 ( .A(n893), .B(A[59]), .Z(n4942) );
  AND U5912 ( .A(n4945), .B(n4946), .Z(n893) );
  NANDN U5913 ( .A(B[58]), .B(n4947), .Z(n4946) );
  NANDN U5914 ( .A(A[58]), .B(n915), .Z(n4947) );
  NANDN U5915 ( .A(n915), .B(A[58]), .Z(n4945) );
  AND U5916 ( .A(n4948), .B(n4949), .Z(n915) );
  NANDN U5917 ( .A(B[57]), .B(n4950), .Z(n4949) );
  NANDN U5918 ( .A(A[57]), .B(n937), .Z(n4950) );
  NANDN U5919 ( .A(n937), .B(A[57]), .Z(n4948) );
  AND U5920 ( .A(n4951), .B(n4952), .Z(n937) );
  NANDN U5921 ( .A(B[56]), .B(n4953), .Z(n4952) );
  NANDN U5922 ( .A(A[56]), .B(n959), .Z(n4953) );
  NANDN U5923 ( .A(n959), .B(A[56]), .Z(n4951) );
  AND U5924 ( .A(n4954), .B(n4955), .Z(n959) );
  NANDN U5925 ( .A(B[55]), .B(n4956), .Z(n4955) );
  NANDN U5926 ( .A(A[55]), .B(n981), .Z(n4956) );
  NANDN U5927 ( .A(n981), .B(A[55]), .Z(n4954) );
  AND U5928 ( .A(n4957), .B(n4958), .Z(n981) );
  NANDN U5929 ( .A(B[54]), .B(n4959), .Z(n4958) );
  NANDN U5930 ( .A(A[54]), .B(n1003), .Z(n4959) );
  NANDN U5931 ( .A(n1003), .B(A[54]), .Z(n4957) );
  AND U5932 ( .A(n4960), .B(n4961), .Z(n1003) );
  NANDN U5933 ( .A(B[53]), .B(n4962), .Z(n4961) );
  NANDN U5934 ( .A(A[53]), .B(n1025), .Z(n4962) );
  NANDN U5935 ( .A(n1025), .B(A[53]), .Z(n4960) );
  AND U5936 ( .A(n4963), .B(n4964), .Z(n1025) );
  NANDN U5937 ( .A(B[52]), .B(n4965), .Z(n4964) );
  NANDN U5938 ( .A(A[52]), .B(n1047), .Z(n4965) );
  NANDN U5939 ( .A(n1047), .B(A[52]), .Z(n4963) );
  AND U5940 ( .A(n4966), .B(n4967), .Z(n1047) );
  NANDN U5941 ( .A(B[51]), .B(n4968), .Z(n4967) );
  NANDN U5942 ( .A(A[51]), .B(n1069), .Z(n4968) );
  NANDN U5943 ( .A(n1069), .B(A[51]), .Z(n4966) );
  AND U5944 ( .A(n4969), .B(n4970), .Z(n1069) );
  NANDN U5945 ( .A(B[50]), .B(n4971), .Z(n4970) );
  NANDN U5946 ( .A(A[50]), .B(n1091), .Z(n4971) );
  NANDN U5947 ( .A(n1091), .B(A[50]), .Z(n4969) );
  AND U5948 ( .A(n4972), .B(n4973), .Z(n1091) );
  NANDN U5949 ( .A(B[49]), .B(n4974), .Z(n4973) );
  NANDN U5950 ( .A(A[49]), .B(n1115), .Z(n4974) );
  NANDN U5951 ( .A(n1115), .B(A[49]), .Z(n4972) );
  AND U5952 ( .A(n4975), .B(n4976), .Z(n1115) );
  NANDN U5953 ( .A(B[48]), .B(n4977), .Z(n4976) );
  NANDN U5954 ( .A(A[48]), .B(n1137), .Z(n4977) );
  NANDN U5955 ( .A(n1137), .B(A[48]), .Z(n4975) );
  AND U5956 ( .A(n4978), .B(n4979), .Z(n1137) );
  NANDN U5957 ( .A(B[47]), .B(n4980), .Z(n4979) );
  NANDN U5958 ( .A(A[47]), .B(n1159), .Z(n4980) );
  NANDN U5959 ( .A(n1159), .B(A[47]), .Z(n4978) );
  AND U5960 ( .A(n4981), .B(n4982), .Z(n1159) );
  NANDN U5961 ( .A(B[46]), .B(n4983), .Z(n4982) );
  NANDN U5962 ( .A(A[46]), .B(n1181), .Z(n4983) );
  NANDN U5963 ( .A(n1181), .B(A[46]), .Z(n4981) );
  AND U5964 ( .A(n4984), .B(n4985), .Z(n1181) );
  NANDN U5965 ( .A(B[45]), .B(n4986), .Z(n4985) );
  NANDN U5966 ( .A(A[45]), .B(n1203), .Z(n4986) );
  NANDN U5967 ( .A(n1203), .B(A[45]), .Z(n4984) );
  AND U5968 ( .A(n4987), .B(n4988), .Z(n1203) );
  NANDN U5969 ( .A(B[44]), .B(n4989), .Z(n4988) );
  NANDN U5970 ( .A(A[44]), .B(n1225), .Z(n4989) );
  NANDN U5971 ( .A(n1225), .B(A[44]), .Z(n4987) );
  AND U5972 ( .A(n4990), .B(n4991), .Z(n1225) );
  NANDN U5973 ( .A(B[43]), .B(n4992), .Z(n4991) );
  NANDN U5974 ( .A(A[43]), .B(n1247), .Z(n4992) );
  NANDN U5975 ( .A(n1247), .B(A[43]), .Z(n4990) );
  AND U5976 ( .A(n4993), .B(n4994), .Z(n1247) );
  NANDN U5977 ( .A(B[42]), .B(n4995), .Z(n4994) );
  NANDN U5978 ( .A(A[42]), .B(n1269), .Z(n4995) );
  NANDN U5979 ( .A(n1269), .B(A[42]), .Z(n4993) );
  AND U5980 ( .A(n4996), .B(n4997), .Z(n1269) );
  NANDN U5981 ( .A(B[41]), .B(n4998), .Z(n4997) );
  NANDN U5982 ( .A(A[41]), .B(n1291), .Z(n4998) );
  NANDN U5983 ( .A(n1291), .B(A[41]), .Z(n4996) );
  AND U5984 ( .A(n4999), .B(n5000), .Z(n1291) );
  NANDN U5985 ( .A(B[40]), .B(n5001), .Z(n5000) );
  NANDN U5986 ( .A(A[40]), .B(n1313), .Z(n5001) );
  NANDN U5987 ( .A(n1313), .B(A[40]), .Z(n4999) );
  AND U5988 ( .A(n5002), .B(n5003), .Z(n1313) );
  NANDN U5989 ( .A(B[39]), .B(n5004), .Z(n5003) );
  NANDN U5990 ( .A(A[39]), .B(n1337), .Z(n5004) );
  NANDN U5991 ( .A(n1337), .B(A[39]), .Z(n5002) );
  AND U5992 ( .A(n5005), .B(n5006), .Z(n1337) );
  NANDN U5993 ( .A(B[38]), .B(n5007), .Z(n5006) );
  NANDN U5994 ( .A(A[38]), .B(n1359), .Z(n5007) );
  NANDN U5995 ( .A(n1359), .B(A[38]), .Z(n5005) );
  AND U5996 ( .A(n5008), .B(n5009), .Z(n1359) );
  NANDN U5997 ( .A(B[37]), .B(n5010), .Z(n5009) );
  NANDN U5998 ( .A(A[37]), .B(n1381), .Z(n5010) );
  NANDN U5999 ( .A(n1381), .B(A[37]), .Z(n5008) );
  AND U6000 ( .A(n5011), .B(n5012), .Z(n1381) );
  NANDN U6001 ( .A(B[36]), .B(n5013), .Z(n5012) );
  NANDN U6002 ( .A(A[36]), .B(n1403), .Z(n5013) );
  NANDN U6003 ( .A(n1403), .B(A[36]), .Z(n5011) );
  AND U6004 ( .A(n5014), .B(n5015), .Z(n1403) );
  NANDN U6005 ( .A(B[35]), .B(n5016), .Z(n5015) );
  NANDN U6006 ( .A(A[35]), .B(n1425), .Z(n5016) );
  NANDN U6007 ( .A(n1425), .B(A[35]), .Z(n5014) );
  AND U6008 ( .A(n5017), .B(n5018), .Z(n1425) );
  NANDN U6009 ( .A(B[34]), .B(n5019), .Z(n5018) );
  NANDN U6010 ( .A(A[34]), .B(n1447), .Z(n5019) );
  NANDN U6011 ( .A(n1447), .B(A[34]), .Z(n5017) );
  AND U6012 ( .A(n5020), .B(n5021), .Z(n1447) );
  NANDN U6013 ( .A(B[33]), .B(n5022), .Z(n5021) );
  NANDN U6014 ( .A(A[33]), .B(n1469), .Z(n5022) );
  NANDN U6015 ( .A(n1469), .B(A[33]), .Z(n5020) );
  AND U6016 ( .A(n5023), .B(n5024), .Z(n1469) );
  NANDN U6017 ( .A(B[32]), .B(n5025), .Z(n5024) );
  NANDN U6018 ( .A(A[32]), .B(n1491), .Z(n5025) );
  NANDN U6019 ( .A(n1491), .B(A[32]), .Z(n5023) );
  AND U6020 ( .A(n5026), .B(n5027), .Z(n1491) );
  NANDN U6021 ( .A(B[31]), .B(n5028), .Z(n5027) );
  NANDN U6022 ( .A(A[31]), .B(n1513), .Z(n5028) );
  NANDN U6023 ( .A(n1513), .B(A[31]), .Z(n5026) );
  AND U6024 ( .A(n5029), .B(n5030), .Z(n1513) );
  NANDN U6025 ( .A(B[30]), .B(n5031), .Z(n5030) );
  NANDN U6026 ( .A(A[30]), .B(n1535), .Z(n5031) );
  NANDN U6027 ( .A(n1535), .B(A[30]), .Z(n5029) );
  AND U6028 ( .A(n5032), .B(n5033), .Z(n1535) );
  NANDN U6029 ( .A(B[29]), .B(n5034), .Z(n5033) );
  NANDN U6030 ( .A(A[29]), .B(n1559), .Z(n5034) );
  NANDN U6031 ( .A(n1559), .B(A[29]), .Z(n5032) );
  AND U6032 ( .A(n5035), .B(n5036), .Z(n1559) );
  NANDN U6033 ( .A(B[28]), .B(n5037), .Z(n5036) );
  NANDN U6034 ( .A(A[28]), .B(n1581), .Z(n5037) );
  NANDN U6035 ( .A(n1581), .B(A[28]), .Z(n5035) );
  AND U6036 ( .A(n5038), .B(n5039), .Z(n1581) );
  NANDN U6037 ( .A(B[27]), .B(n5040), .Z(n5039) );
  NANDN U6038 ( .A(A[27]), .B(n1603), .Z(n5040) );
  NANDN U6039 ( .A(n1603), .B(A[27]), .Z(n5038) );
  AND U6040 ( .A(n5041), .B(n5042), .Z(n1603) );
  NANDN U6041 ( .A(B[26]), .B(n5043), .Z(n5042) );
  NANDN U6042 ( .A(A[26]), .B(n1625), .Z(n5043) );
  NANDN U6043 ( .A(n1625), .B(A[26]), .Z(n5041) );
  AND U6044 ( .A(n5044), .B(n5045), .Z(n1625) );
  NANDN U6045 ( .A(B[25]), .B(n5046), .Z(n5045) );
  NANDN U6046 ( .A(A[25]), .B(n1647), .Z(n5046) );
  NANDN U6047 ( .A(n1647), .B(A[25]), .Z(n5044) );
  AND U6048 ( .A(n5047), .B(n5048), .Z(n1647) );
  NANDN U6049 ( .A(B[24]), .B(n5049), .Z(n5048) );
  NANDN U6050 ( .A(A[24]), .B(n1669), .Z(n5049) );
  NANDN U6051 ( .A(n1669), .B(A[24]), .Z(n5047) );
  AND U6052 ( .A(n5050), .B(n5051), .Z(n1669) );
  NANDN U6053 ( .A(B[23]), .B(n5052), .Z(n5051) );
  NANDN U6054 ( .A(A[23]), .B(n1691), .Z(n5052) );
  NANDN U6055 ( .A(n1691), .B(A[23]), .Z(n5050) );
  AND U6056 ( .A(n5053), .B(n5054), .Z(n1691) );
  NANDN U6057 ( .A(B[22]), .B(n5055), .Z(n5054) );
  NANDN U6058 ( .A(A[22]), .B(n1713), .Z(n5055) );
  NANDN U6059 ( .A(n1713), .B(A[22]), .Z(n5053) );
  AND U6060 ( .A(n5056), .B(n5057), .Z(n1713) );
  NANDN U6061 ( .A(B[21]), .B(n5058), .Z(n5057) );
  NANDN U6062 ( .A(A[21]), .B(n1735), .Z(n5058) );
  NANDN U6063 ( .A(n1735), .B(A[21]), .Z(n5056) );
  AND U6064 ( .A(n5059), .B(n5060), .Z(n1735) );
  NANDN U6065 ( .A(B[20]), .B(n5061), .Z(n5060) );
  NANDN U6066 ( .A(A[20]), .B(n1757), .Z(n5061) );
  NANDN U6067 ( .A(n1757), .B(A[20]), .Z(n5059) );
  AND U6068 ( .A(n5062), .B(n5063), .Z(n1757) );
  NANDN U6069 ( .A(B[19]), .B(n5064), .Z(n5063) );
  NANDN U6070 ( .A(A[19]), .B(n1780), .Z(n5064) );
  NANDN U6071 ( .A(n1780), .B(A[19]), .Z(n5062) );
  AND U6072 ( .A(n5065), .B(n5066), .Z(n1780) );
  NANDN U6073 ( .A(B[18]), .B(n5067), .Z(n5066) );
  NANDN U6074 ( .A(A[18]), .B(n1802), .Z(n5067) );
  NANDN U6075 ( .A(n1802), .B(A[18]), .Z(n5065) );
  AND U6076 ( .A(n5068), .B(n5069), .Z(n1802) );
  NANDN U6077 ( .A(B[17]), .B(n5070), .Z(n5069) );
  NANDN U6078 ( .A(A[17]), .B(n1824), .Z(n5070) );
  NANDN U6079 ( .A(n1824), .B(A[17]), .Z(n5068) );
  AND U6080 ( .A(n5071), .B(n5072), .Z(n1824) );
  NANDN U6081 ( .A(B[16]), .B(n5073), .Z(n5072) );
  NANDN U6082 ( .A(A[16]), .B(n1846), .Z(n5073) );
  NANDN U6083 ( .A(n1846), .B(A[16]), .Z(n5071) );
  AND U6084 ( .A(n5074), .B(n5075), .Z(n1846) );
  NANDN U6085 ( .A(B[15]), .B(n5076), .Z(n5075) );
  NANDN U6086 ( .A(A[15]), .B(n1868), .Z(n5076) );
  NANDN U6087 ( .A(n1868), .B(A[15]), .Z(n5074) );
  AND U6088 ( .A(n5077), .B(n5078), .Z(n1868) );
  NANDN U6089 ( .A(B[14]), .B(n5079), .Z(n5078) );
  NANDN U6090 ( .A(A[14]), .B(n1890), .Z(n5079) );
  NANDN U6091 ( .A(n1890), .B(A[14]), .Z(n5077) );
  AND U6092 ( .A(n5080), .B(n5081), .Z(n1890) );
  NANDN U6093 ( .A(B[13]), .B(n5082), .Z(n5081) );
  NANDN U6094 ( .A(A[13]), .B(n1912), .Z(n5082) );
  NANDN U6095 ( .A(n1912), .B(A[13]), .Z(n5080) );
  AND U6096 ( .A(n5083), .B(n5084), .Z(n1912) );
  NANDN U6097 ( .A(B[12]), .B(n5085), .Z(n5084) );
  NANDN U6098 ( .A(A[12]), .B(n1934), .Z(n5085) );
  NANDN U6099 ( .A(n1934), .B(A[12]), .Z(n5083) );
  AND U6100 ( .A(n5086), .B(n5087), .Z(n1934) );
  NANDN U6101 ( .A(B[11]), .B(n5088), .Z(n5087) );
  NANDN U6102 ( .A(A[11]), .B(n1956), .Z(n5088) );
  NANDN U6103 ( .A(n1956), .B(A[11]), .Z(n5086) );
  AND U6104 ( .A(n5089), .B(n5090), .Z(n1956) );
  NANDN U6105 ( .A(B[10]), .B(n5091), .Z(n5090) );
  NANDN U6106 ( .A(A[10]), .B(n1978), .Z(n5091) );
  NANDN U6107 ( .A(n1978), .B(A[10]), .Z(n5089) );
  AND U6108 ( .A(n5092), .B(n5093), .Z(n1978) );
  NANDN U6109 ( .A(B[9]), .B(n5094), .Z(n5093) );
  OR U6110 ( .A(n3), .B(A[9]), .Z(n5094) );
  NAND U6111 ( .A(A[9]), .B(n3), .Z(n5092) );
  NAND U6112 ( .A(n5095), .B(n5096), .Z(n3) );
  NANDN U6113 ( .A(B[8]), .B(n5097), .Z(n5096) );
  NANDN U6114 ( .A(A[8]), .B(n225), .Z(n5097) );
  NANDN U6115 ( .A(n225), .B(A[8]), .Z(n5095) );
  AND U6116 ( .A(n5098), .B(n5099), .Z(n225) );
  NANDN U6117 ( .A(B[7]), .B(n5100), .Z(n5099) );
  NANDN U6118 ( .A(A[7]), .B(n447), .Z(n5100) );
  NANDN U6119 ( .A(n447), .B(A[7]), .Z(n5098) );
  AND U6120 ( .A(n5101), .B(n5102), .Z(n447) );
  NANDN U6121 ( .A(B[6]), .B(n5103), .Z(n5102) );
  NANDN U6122 ( .A(A[6]), .B(n669), .Z(n5103) );
  NANDN U6123 ( .A(n669), .B(A[6]), .Z(n5101) );
  AND U6124 ( .A(n5104), .B(n5105), .Z(n669) );
  NANDN U6125 ( .A(B[5]), .B(n5106), .Z(n5105) );
  NANDN U6126 ( .A(A[5]), .B(n891), .Z(n5106) );
  NANDN U6127 ( .A(n891), .B(A[5]), .Z(n5104) );
  AND U6128 ( .A(n5107), .B(n5108), .Z(n891) );
  NANDN U6129 ( .A(B[4]), .B(n5109), .Z(n5108) );
  NANDN U6130 ( .A(A[4]), .B(n1113), .Z(n5109) );
  NANDN U6131 ( .A(n1113), .B(A[4]), .Z(n5107) );
  AND U6132 ( .A(n5110), .B(n5111), .Z(n1113) );
  NANDN U6133 ( .A(B[3]), .B(n5112), .Z(n5111) );
  NANDN U6134 ( .A(A[3]), .B(n1335), .Z(n5112) );
  NANDN U6135 ( .A(n1335), .B(A[3]), .Z(n5110) );
  AND U6136 ( .A(n5113), .B(n5114), .Z(n1335) );
  NANDN U6137 ( .A(B[2]), .B(n5115), .Z(n5114) );
  NANDN U6138 ( .A(A[2]), .B(n1557), .Z(n5115) );
  NANDN U6139 ( .A(n1557), .B(A[2]), .Z(n5113) );
  AND U6140 ( .A(n5116), .B(n5117), .Z(n1557) );
  NANDN U6141 ( .A(B[1]), .B(n5118), .Z(n5117) );
  NAND U6142 ( .A(n2), .B(n1), .Z(n5118) );
  NAND U6143 ( .A(A[1]), .B(n5119), .Z(n5116) );
  NAND U6144 ( .A(n5119), .B(n5120), .Z(DIFF[0]) );
  NANDN U6145 ( .A(B[0]), .B(A[0]), .Z(n5120) );
  NANDN U6146 ( .A(A[0]), .B(B[0]), .Z(n5119) );
endmodule


module modmult_step_N1024_DW01_cmp2_1 ( A, B, LEQ, TC, LT_LE, GE_GT );
  input [1025:0] A;
  input [1025:0] B;
  input LEQ, TC;
  output LT_LE, GE_GT;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094;

  NAND U1 ( .A(n1), .B(n2), .Z(LT_LE) );
  NOR U2 ( .A(B[1025]), .B(B[1024]), .Z(n2) );
  AND U3 ( .A(n3), .B(n4), .Z(n1) );
  NAND U4 ( .A(n5), .B(n6), .Z(n4) );
  NANDN U5 ( .A(B[1023]), .B(A[1023]), .Z(n6) );
  NAND U6 ( .A(n7), .B(n8), .Z(n5) );
  NANDN U7 ( .A(A[1022]), .B(B[1022]), .Z(n8) );
  NAND U8 ( .A(n9), .B(n10), .Z(n7) );
  NANDN U9 ( .A(B[1022]), .B(A[1022]), .Z(n10) );
  AND U10 ( .A(n11), .B(n12), .Z(n9) );
  NAND U11 ( .A(n13), .B(n14), .Z(n12) );
  NANDN U12 ( .A(A[1021]), .B(B[1021]), .Z(n14) );
  AND U13 ( .A(n15), .B(n16), .Z(n13) );
  NANDN U14 ( .A(A[1020]), .B(B[1020]), .Z(n16) );
  NAND U15 ( .A(n17), .B(n18), .Z(n15) );
  NANDN U16 ( .A(B[1020]), .B(A[1020]), .Z(n18) );
  AND U17 ( .A(n19), .B(n20), .Z(n17) );
  NAND U18 ( .A(n21), .B(n22), .Z(n20) );
  NANDN U19 ( .A(A[1019]), .B(B[1019]), .Z(n22) );
  AND U20 ( .A(n23), .B(n24), .Z(n21) );
  NANDN U21 ( .A(A[1018]), .B(B[1018]), .Z(n24) );
  NAND U22 ( .A(n25), .B(n26), .Z(n23) );
  NANDN U23 ( .A(B[1018]), .B(A[1018]), .Z(n26) );
  AND U24 ( .A(n27), .B(n28), .Z(n25) );
  NAND U25 ( .A(n29), .B(n30), .Z(n28) );
  NANDN U26 ( .A(A[1017]), .B(B[1017]), .Z(n30) );
  AND U27 ( .A(n31), .B(n32), .Z(n29) );
  NANDN U28 ( .A(A[1016]), .B(B[1016]), .Z(n32) );
  NAND U29 ( .A(n33), .B(n34), .Z(n31) );
  NANDN U30 ( .A(B[1016]), .B(A[1016]), .Z(n34) );
  AND U31 ( .A(n35), .B(n36), .Z(n33) );
  NAND U32 ( .A(n37), .B(n38), .Z(n36) );
  NANDN U33 ( .A(A[1015]), .B(B[1015]), .Z(n38) );
  AND U34 ( .A(n39), .B(n40), .Z(n37) );
  NANDN U35 ( .A(A[1014]), .B(B[1014]), .Z(n40) );
  NAND U36 ( .A(n41), .B(n42), .Z(n39) );
  NANDN U37 ( .A(B[1014]), .B(A[1014]), .Z(n42) );
  AND U38 ( .A(n43), .B(n44), .Z(n41) );
  NAND U39 ( .A(n45), .B(n46), .Z(n44) );
  NANDN U40 ( .A(A[1013]), .B(B[1013]), .Z(n46) );
  AND U41 ( .A(n47), .B(n48), .Z(n45) );
  NANDN U42 ( .A(A[1012]), .B(B[1012]), .Z(n48) );
  NAND U43 ( .A(n49), .B(n50), .Z(n47) );
  NANDN U44 ( .A(B[1012]), .B(A[1012]), .Z(n50) );
  AND U45 ( .A(n51), .B(n52), .Z(n49) );
  NAND U46 ( .A(n53), .B(n54), .Z(n52) );
  NANDN U47 ( .A(A[1011]), .B(B[1011]), .Z(n54) );
  AND U48 ( .A(n55), .B(n56), .Z(n53) );
  NANDN U49 ( .A(A[1010]), .B(B[1010]), .Z(n56) );
  NAND U50 ( .A(n57), .B(n58), .Z(n55) );
  NANDN U51 ( .A(B[1010]), .B(A[1010]), .Z(n58) );
  AND U52 ( .A(n59), .B(n60), .Z(n57) );
  NAND U53 ( .A(n61), .B(n62), .Z(n60) );
  NANDN U54 ( .A(A[1009]), .B(B[1009]), .Z(n62) );
  AND U55 ( .A(n63), .B(n64), .Z(n61) );
  NANDN U56 ( .A(A[1008]), .B(B[1008]), .Z(n64) );
  NAND U57 ( .A(n65), .B(n66), .Z(n63) );
  NANDN U58 ( .A(B[1008]), .B(A[1008]), .Z(n66) );
  AND U59 ( .A(n67), .B(n68), .Z(n65) );
  NAND U60 ( .A(n69), .B(n70), .Z(n68) );
  NANDN U61 ( .A(A[1007]), .B(B[1007]), .Z(n70) );
  AND U62 ( .A(n71), .B(n72), .Z(n69) );
  NANDN U63 ( .A(A[1006]), .B(B[1006]), .Z(n72) );
  NAND U64 ( .A(n73), .B(n74), .Z(n71) );
  NANDN U65 ( .A(B[1006]), .B(A[1006]), .Z(n74) );
  AND U66 ( .A(n75), .B(n76), .Z(n73) );
  NAND U67 ( .A(n77), .B(n78), .Z(n76) );
  NANDN U68 ( .A(A[1005]), .B(B[1005]), .Z(n78) );
  AND U69 ( .A(n79), .B(n80), .Z(n77) );
  NANDN U70 ( .A(A[1004]), .B(B[1004]), .Z(n80) );
  NAND U71 ( .A(n81), .B(n82), .Z(n79) );
  NANDN U72 ( .A(B[1004]), .B(A[1004]), .Z(n82) );
  AND U73 ( .A(n83), .B(n84), .Z(n81) );
  NAND U74 ( .A(n85), .B(n86), .Z(n84) );
  NANDN U75 ( .A(A[1003]), .B(B[1003]), .Z(n86) );
  AND U76 ( .A(n87), .B(n88), .Z(n85) );
  NANDN U77 ( .A(A[1002]), .B(B[1002]), .Z(n88) );
  NAND U78 ( .A(n89), .B(n90), .Z(n87) );
  NANDN U79 ( .A(B[1002]), .B(A[1002]), .Z(n90) );
  AND U80 ( .A(n91), .B(n92), .Z(n89) );
  NAND U81 ( .A(n93), .B(n94), .Z(n92) );
  NANDN U82 ( .A(A[1001]), .B(B[1001]), .Z(n94) );
  AND U83 ( .A(n95), .B(n96), .Z(n93) );
  NANDN U84 ( .A(A[1000]), .B(B[1000]), .Z(n96) );
  NAND U85 ( .A(n97), .B(n98), .Z(n95) );
  NANDN U86 ( .A(B[999]), .B(A[999]), .Z(n98) );
  AND U87 ( .A(n99), .B(n100), .Z(n97) );
  NAND U88 ( .A(n101), .B(n102), .Z(n100) );
  NANDN U89 ( .A(A[999]), .B(B[999]), .Z(n102) );
  AND U90 ( .A(n103), .B(n104), .Z(n101) );
  NANDN U91 ( .A(A[998]), .B(B[998]), .Z(n104) );
  NAND U92 ( .A(n105), .B(n106), .Z(n103) );
  NANDN U93 ( .A(B[998]), .B(A[998]), .Z(n106) );
  AND U94 ( .A(n107), .B(n108), .Z(n105) );
  NAND U95 ( .A(n109), .B(n110), .Z(n108) );
  NANDN U96 ( .A(A[997]), .B(B[997]), .Z(n110) );
  AND U97 ( .A(n111), .B(n112), .Z(n109) );
  NANDN U98 ( .A(A[996]), .B(B[996]), .Z(n112) );
  NAND U99 ( .A(n113), .B(n114), .Z(n111) );
  NANDN U100 ( .A(B[996]), .B(A[996]), .Z(n114) );
  AND U101 ( .A(n115), .B(n116), .Z(n113) );
  NAND U102 ( .A(n117), .B(n118), .Z(n116) );
  NANDN U103 ( .A(A[995]), .B(B[995]), .Z(n118) );
  AND U104 ( .A(n119), .B(n120), .Z(n117) );
  NANDN U105 ( .A(A[994]), .B(B[994]), .Z(n120) );
  NAND U106 ( .A(n121), .B(n122), .Z(n119) );
  NANDN U107 ( .A(B[994]), .B(A[994]), .Z(n122) );
  AND U108 ( .A(n123), .B(n124), .Z(n121) );
  NAND U109 ( .A(n125), .B(n126), .Z(n124) );
  NANDN U110 ( .A(A[993]), .B(B[993]), .Z(n126) );
  AND U111 ( .A(n127), .B(n128), .Z(n125) );
  NANDN U112 ( .A(A[992]), .B(B[992]), .Z(n128) );
  NAND U113 ( .A(n129), .B(n130), .Z(n127) );
  NANDN U114 ( .A(B[992]), .B(A[992]), .Z(n130) );
  AND U115 ( .A(n131), .B(n132), .Z(n129) );
  NAND U116 ( .A(n133), .B(n134), .Z(n132) );
  NANDN U117 ( .A(A[991]), .B(B[991]), .Z(n134) );
  AND U118 ( .A(n135), .B(n136), .Z(n133) );
  NANDN U119 ( .A(A[990]), .B(B[990]), .Z(n136) );
  NAND U120 ( .A(n137), .B(n138), .Z(n135) );
  NANDN U121 ( .A(B[990]), .B(A[990]), .Z(n138) );
  AND U122 ( .A(n139), .B(n140), .Z(n137) );
  NAND U123 ( .A(n141), .B(n142), .Z(n140) );
  NANDN U124 ( .A(A[989]), .B(B[989]), .Z(n142) );
  AND U125 ( .A(n143), .B(n144), .Z(n141) );
  NANDN U126 ( .A(A[988]), .B(B[988]), .Z(n144) );
  NAND U127 ( .A(n145), .B(n146), .Z(n143) );
  NANDN U128 ( .A(B[988]), .B(A[988]), .Z(n146) );
  AND U129 ( .A(n147), .B(n148), .Z(n145) );
  NAND U130 ( .A(n149), .B(n150), .Z(n148) );
  NANDN U131 ( .A(A[987]), .B(B[987]), .Z(n150) );
  AND U132 ( .A(n151), .B(n152), .Z(n149) );
  NANDN U133 ( .A(A[986]), .B(B[986]), .Z(n152) );
  NAND U134 ( .A(n153), .B(n154), .Z(n151) );
  NANDN U135 ( .A(B[986]), .B(A[986]), .Z(n154) );
  AND U136 ( .A(n155), .B(n156), .Z(n153) );
  NAND U137 ( .A(n157), .B(n158), .Z(n156) );
  NANDN U138 ( .A(A[985]), .B(B[985]), .Z(n158) );
  AND U139 ( .A(n159), .B(n160), .Z(n157) );
  NANDN U140 ( .A(A[984]), .B(B[984]), .Z(n160) );
  NAND U141 ( .A(n161), .B(n162), .Z(n159) );
  NANDN U142 ( .A(B[984]), .B(A[984]), .Z(n162) );
  AND U143 ( .A(n163), .B(n164), .Z(n161) );
  NAND U144 ( .A(n165), .B(n166), .Z(n164) );
  NANDN U145 ( .A(A[983]), .B(B[983]), .Z(n166) );
  AND U146 ( .A(n167), .B(n168), .Z(n165) );
  NANDN U147 ( .A(A[982]), .B(B[982]), .Z(n168) );
  NAND U148 ( .A(n169), .B(n170), .Z(n167) );
  NANDN U149 ( .A(B[982]), .B(A[982]), .Z(n170) );
  AND U150 ( .A(n171), .B(n172), .Z(n169) );
  NAND U151 ( .A(n173), .B(n174), .Z(n172) );
  NANDN U152 ( .A(A[981]), .B(B[981]), .Z(n174) );
  AND U153 ( .A(n175), .B(n176), .Z(n173) );
  NANDN U154 ( .A(A[980]), .B(B[980]), .Z(n176) );
  NAND U155 ( .A(n177), .B(n178), .Z(n175) );
  NANDN U156 ( .A(B[980]), .B(A[980]), .Z(n178) );
  AND U157 ( .A(n179), .B(n180), .Z(n177) );
  NAND U158 ( .A(n181), .B(n182), .Z(n180) );
  NANDN U159 ( .A(A[979]), .B(B[979]), .Z(n182) );
  AND U160 ( .A(n183), .B(n184), .Z(n181) );
  NANDN U161 ( .A(A[978]), .B(B[978]), .Z(n184) );
  NAND U162 ( .A(n185), .B(n186), .Z(n183) );
  NANDN U163 ( .A(B[978]), .B(A[978]), .Z(n186) );
  AND U164 ( .A(n187), .B(n188), .Z(n185) );
  NAND U165 ( .A(n189), .B(n190), .Z(n188) );
  NANDN U166 ( .A(A[977]), .B(B[977]), .Z(n190) );
  AND U167 ( .A(n191), .B(n192), .Z(n189) );
  NANDN U168 ( .A(A[976]), .B(B[976]), .Z(n192) );
  NAND U169 ( .A(n193), .B(n194), .Z(n191) );
  NANDN U170 ( .A(B[976]), .B(A[976]), .Z(n194) );
  AND U171 ( .A(n195), .B(n196), .Z(n193) );
  NAND U172 ( .A(n197), .B(n198), .Z(n196) );
  NANDN U173 ( .A(A[975]), .B(B[975]), .Z(n198) );
  AND U174 ( .A(n199), .B(n200), .Z(n197) );
  NANDN U175 ( .A(A[974]), .B(B[974]), .Z(n200) );
  NAND U176 ( .A(n201), .B(n202), .Z(n199) );
  NANDN U177 ( .A(B[974]), .B(A[974]), .Z(n202) );
  AND U178 ( .A(n203), .B(n204), .Z(n201) );
  NAND U179 ( .A(n205), .B(n206), .Z(n204) );
  NANDN U180 ( .A(A[973]), .B(B[973]), .Z(n206) );
  AND U181 ( .A(n207), .B(n208), .Z(n205) );
  NANDN U182 ( .A(A[972]), .B(B[972]), .Z(n208) );
  NAND U183 ( .A(n209), .B(n210), .Z(n207) );
  NANDN U184 ( .A(B[972]), .B(A[972]), .Z(n210) );
  AND U185 ( .A(n211), .B(n212), .Z(n209) );
  NAND U186 ( .A(n213), .B(n214), .Z(n212) );
  NANDN U187 ( .A(A[971]), .B(B[971]), .Z(n214) );
  AND U188 ( .A(n215), .B(n216), .Z(n213) );
  NANDN U189 ( .A(A[970]), .B(B[970]), .Z(n216) );
  NAND U190 ( .A(n217), .B(n218), .Z(n215) );
  NANDN U191 ( .A(B[970]), .B(A[970]), .Z(n218) );
  AND U192 ( .A(n219), .B(n220), .Z(n217) );
  NAND U193 ( .A(n221), .B(n222), .Z(n220) );
  NANDN U194 ( .A(A[969]), .B(B[969]), .Z(n222) );
  AND U195 ( .A(n223), .B(n224), .Z(n221) );
  NANDN U196 ( .A(A[968]), .B(B[968]), .Z(n224) );
  NAND U197 ( .A(n225), .B(n226), .Z(n223) );
  NANDN U198 ( .A(B[968]), .B(A[968]), .Z(n226) );
  AND U199 ( .A(n227), .B(n228), .Z(n225) );
  NAND U200 ( .A(n229), .B(n230), .Z(n228) );
  NANDN U201 ( .A(A[967]), .B(B[967]), .Z(n230) );
  AND U202 ( .A(n231), .B(n232), .Z(n229) );
  NANDN U203 ( .A(A[966]), .B(B[966]), .Z(n232) );
  NAND U204 ( .A(n233), .B(n234), .Z(n231) );
  NANDN U205 ( .A(B[966]), .B(A[966]), .Z(n234) );
  AND U206 ( .A(n235), .B(n236), .Z(n233) );
  NAND U207 ( .A(n237), .B(n238), .Z(n236) );
  NANDN U208 ( .A(A[965]), .B(B[965]), .Z(n238) );
  AND U209 ( .A(n239), .B(n240), .Z(n237) );
  NANDN U210 ( .A(A[964]), .B(B[964]), .Z(n240) );
  NAND U211 ( .A(n241), .B(n242), .Z(n239) );
  NANDN U212 ( .A(B[964]), .B(A[964]), .Z(n242) );
  AND U213 ( .A(n243), .B(n244), .Z(n241) );
  NAND U214 ( .A(n245), .B(n246), .Z(n244) );
  NANDN U215 ( .A(A[963]), .B(B[963]), .Z(n246) );
  AND U216 ( .A(n247), .B(n248), .Z(n245) );
  NANDN U217 ( .A(A[962]), .B(B[962]), .Z(n248) );
  NAND U218 ( .A(n249), .B(n250), .Z(n247) );
  NANDN U219 ( .A(B[962]), .B(A[962]), .Z(n250) );
  AND U220 ( .A(n251), .B(n252), .Z(n249) );
  NAND U221 ( .A(n253), .B(n254), .Z(n252) );
  NANDN U222 ( .A(A[961]), .B(B[961]), .Z(n254) );
  AND U223 ( .A(n255), .B(n256), .Z(n253) );
  NANDN U224 ( .A(A[960]), .B(B[960]), .Z(n256) );
  NAND U225 ( .A(n257), .B(n258), .Z(n255) );
  NANDN U226 ( .A(B[960]), .B(A[960]), .Z(n258) );
  AND U227 ( .A(n259), .B(n260), .Z(n257) );
  NAND U228 ( .A(n261), .B(n262), .Z(n260) );
  NANDN U229 ( .A(A[959]), .B(B[959]), .Z(n262) );
  AND U230 ( .A(n263), .B(n264), .Z(n261) );
  NANDN U231 ( .A(A[958]), .B(B[958]), .Z(n264) );
  NAND U232 ( .A(n265), .B(n266), .Z(n263) );
  NANDN U233 ( .A(B[958]), .B(A[958]), .Z(n266) );
  AND U234 ( .A(n267), .B(n268), .Z(n265) );
  NAND U235 ( .A(n269), .B(n270), .Z(n268) );
  NANDN U236 ( .A(A[957]), .B(B[957]), .Z(n270) );
  AND U237 ( .A(n271), .B(n272), .Z(n269) );
  NANDN U238 ( .A(A[956]), .B(B[956]), .Z(n272) );
  NAND U239 ( .A(n273), .B(n274), .Z(n271) );
  NANDN U240 ( .A(B[956]), .B(A[956]), .Z(n274) );
  AND U241 ( .A(n275), .B(n276), .Z(n273) );
  NAND U242 ( .A(n277), .B(n278), .Z(n276) );
  NANDN U243 ( .A(A[955]), .B(B[955]), .Z(n278) );
  AND U244 ( .A(n279), .B(n280), .Z(n277) );
  NANDN U245 ( .A(A[954]), .B(B[954]), .Z(n280) );
  NAND U246 ( .A(n281), .B(n282), .Z(n279) );
  NANDN U247 ( .A(B[954]), .B(A[954]), .Z(n282) );
  AND U248 ( .A(n283), .B(n284), .Z(n281) );
  NAND U249 ( .A(n285), .B(n286), .Z(n284) );
  NANDN U250 ( .A(A[953]), .B(B[953]), .Z(n286) );
  AND U251 ( .A(n287), .B(n288), .Z(n285) );
  NANDN U252 ( .A(A[952]), .B(B[952]), .Z(n288) );
  NAND U253 ( .A(n289), .B(n290), .Z(n287) );
  NANDN U254 ( .A(B[952]), .B(A[952]), .Z(n290) );
  AND U255 ( .A(n291), .B(n292), .Z(n289) );
  NAND U256 ( .A(n293), .B(n294), .Z(n292) );
  NANDN U257 ( .A(A[951]), .B(B[951]), .Z(n294) );
  AND U258 ( .A(n295), .B(n296), .Z(n293) );
  NANDN U259 ( .A(A[950]), .B(B[950]), .Z(n296) );
  NAND U260 ( .A(n297), .B(n298), .Z(n295) );
  NANDN U261 ( .A(B[950]), .B(A[950]), .Z(n298) );
  AND U262 ( .A(n299), .B(n300), .Z(n297) );
  NAND U263 ( .A(n301), .B(n302), .Z(n300) );
  NANDN U264 ( .A(A[949]), .B(B[949]), .Z(n302) );
  AND U265 ( .A(n303), .B(n304), .Z(n301) );
  NANDN U266 ( .A(A[948]), .B(B[948]), .Z(n304) );
  NAND U267 ( .A(n305), .B(n306), .Z(n303) );
  NANDN U268 ( .A(B[948]), .B(A[948]), .Z(n306) );
  AND U269 ( .A(n307), .B(n308), .Z(n305) );
  NAND U270 ( .A(n309), .B(n310), .Z(n308) );
  NANDN U271 ( .A(A[947]), .B(B[947]), .Z(n310) );
  AND U272 ( .A(n311), .B(n312), .Z(n309) );
  NANDN U273 ( .A(A[946]), .B(B[946]), .Z(n312) );
  NAND U274 ( .A(n313), .B(n314), .Z(n311) );
  NANDN U275 ( .A(B[946]), .B(A[946]), .Z(n314) );
  AND U276 ( .A(n315), .B(n316), .Z(n313) );
  NAND U277 ( .A(n317), .B(n318), .Z(n316) );
  NANDN U278 ( .A(A[945]), .B(B[945]), .Z(n318) );
  AND U279 ( .A(n319), .B(n320), .Z(n317) );
  NANDN U280 ( .A(A[944]), .B(B[944]), .Z(n320) );
  NAND U281 ( .A(n321), .B(n322), .Z(n319) );
  NANDN U282 ( .A(B[944]), .B(A[944]), .Z(n322) );
  AND U283 ( .A(n323), .B(n324), .Z(n321) );
  NAND U284 ( .A(n325), .B(n326), .Z(n324) );
  NANDN U285 ( .A(A[943]), .B(B[943]), .Z(n326) );
  AND U286 ( .A(n327), .B(n328), .Z(n325) );
  NANDN U287 ( .A(A[942]), .B(B[942]), .Z(n328) );
  NAND U288 ( .A(n329), .B(n330), .Z(n327) );
  NANDN U289 ( .A(B[942]), .B(A[942]), .Z(n330) );
  AND U290 ( .A(n331), .B(n332), .Z(n329) );
  NAND U291 ( .A(n333), .B(n334), .Z(n332) );
  NANDN U292 ( .A(A[941]), .B(B[941]), .Z(n334) );
  AND U293 ( .A(n335), .B(n336), .Z(n333) );
  NANDN U294 ( .A(A[940]), .B(B[940]), .Z(n336) );
  NAND U295 ( .A(n337), .B(n338), .Z(n335) );
  NANDN U296 ( .A(B[940]), .B(A[940]), .Z(n338) );
  AND U297 ( .A(n339), .B(n340), .Z(n337) );
  NAND U298 ( .A(n341), .B(n342), .Z(n340) );
  NANDN U299 ( .A(A[939]), .B(B[939]), .Z(n342) );
  AND U300 ( .A(n343), .B(n344), .Z(n341) );
  NANDN U301 ( .A(A[938]), .B(B[938]), .Z(n344) );
  NAND U302 ( .A(n345), .B(n346), .Z(n343) );
  NANDN U303 ( .A(B[938]), .B(A[938]), .Z(n346) );
  AND U304 ( .A(n347), .B(n348), .Z(n345) );
  NAND U305 ( .A(n349), .B(n350), .Z(n348) );
  NANDN U306 ( .A(A[937]), .B(B[937]), .Z(n350) );
  AND U307 ( .A(n351), .B(n352), .Z(n349) );
  NANDN U308 ( .A(A[936]), .B(B[936]), .Z(n352) );
  NAND U309 ( .A(n353), .B(n354), .Z(n351) );
  NANDN U310 ( .A(B[936]), .B(A[936]), .Z(n354) );
  AND U311 ( .A(n355), .B(n356), .Z(n353) );
  NAND U312 ( .A(n357), .B(n358), .Z(n356) );
  NANDN U313 ( .A(A[935]), .B(B[935]), .Z(n358) );
  AND U314 ( .A(n359), .B(n360), .Z(n357) );
  NANDN U315 ( .A(A[934]), .B(B[934]), .Z(n360) );
  NAND U316 ( .A(n361), .B(n362), .Z(n359) );
  NANDN U317 ( .A(B[934]), .B(A[934]), .Z(n362) );
  AND U318 ( .A(n363), .B(n364), .Z(n361) );
  NAND U319 ( .A(n365), .B(n366), .Z(n364) );
  NANDN U320 ( .A(A[933]), .B(B[933]), .Z(n366) );
  AND U321 ( .A(n367), .B(n368), .Z(n365) );
  NANDN U322 ( .A(A[932]), .B(B[932]), .Z(n368) );
  NAND U323 ( .A(n369), .B(n370), .Z(n367) );
  NANDN U324 ( .A(B[932]), .B(A[932]), .Z(n370) );
  AND U325 ( .A(n371), .B(n372), .Z(n369) );
  NAND U326 ( .A(n373), .B(n374), .Z(n372) );
  NANDN U327 ( .A(A[931]), .B(B[931]), .Z(n374) );
  AND U328 ( .A(n375), .B(n376), .Z(n373) );
  NANDN U329 ( .A(A[930]), .B(B[930]), .Z(n376) );
  NAND U330 ( .A(n377), .B(n378), .Z(n375) );
  NANDN U331 ( .A(B[930]), .B(A[930]), .Z(n378) );
  AND U332 ( .A(n379), .B(n380), .Z(n377) );
  NAND U333 ( .A(n381), .B(n382), .Z(n380) );
  NANDN U334 ( .A(A[929]), .B(B[929]), .Z(n382) );
  AND U335 ( .A(n383), .B(n384), .Z(n381) );
  NANDN U336 ( .A(A[928]), .B(B[928]), .Z(n384) );
  NAND U337 ( .A(n385), .B(n386), .Z(n383) );
  NANDN U338 ( .A(B[928]), .B(A[928]), .Z(n386) );
  AND U339 ( .A(n387), .B(n388), .Z(n385) );
  NAND U340 ( .A(n389), .B(n390), .Z(n388) );
  NANDN U341 ( .A(A[927]), .B(B[927]), .Z(n390) );
  AND U342 ( .A(n391), .B(n392), .Z(n389) );
  NANDN U343 ( .A(A[926]), .B(B[926]), .Z(n392) );
  NAND U344 ( .A(n393), .B(n394), .Z(n391) );
  NANDN U345 ( .A(B[926]), .B(A[926]), .Z(n394) );
  AND U346 ( .A(n395), .B(n396), .Z(n393) );
  NAND U347 ( .A(n397), .B(n398), .Z(n396) );
  NANDN U348 ( .A(A[925]), .B(B[925]), .Z(n398) );
  AND U349 ( .A(n399), .B(n400), .Z(n397) );
  NANDN U350 ( .A(A[924]), .B(B[924]), .Z(n400) );
  NAND U351 ( .A(n401), .B(n402), .Z(n399) );
  NANDN U352 ( .A(B[924]), .B(A[924]), .Z(n402) );
  AND U353 ( .A(n403), .B(n404), .Z(n401) );
  NAND U354 ( .A(n405), .B(n406), .Z(n404) );
  NANDN U355 ( .A(A[923]), .B(B[923]), .Z(n406) );
  AND U356 ( .A(n407), .B(n408), .Z(n405) );
  NANDN U357 ( .A(A[922]), .B(B[922]), .Z(n408) );
  NAND U358 ( .A(n409), .B(n410), .Z(n407) );
  NANDN U359 ( .A(B[922]), .B(A[922]), .Z(n410) );
  AND U360 ( .A(n411), .B(n412), .Z(n409) );
  NAND U361 ( .A(n413), .B(n414), .Z(n412) );
  NANDN U362 ( .A(A[921]), .B(B[921]), .Z(n414) );
  AND U363 ( .A(n415), .B(n416), .Z(n413) );
  NANDN U364 ( .A(A[920]), .B(B[920]), .Z(n416) );
  NAND U365 ( .A(n417), .B(n418), .Z(n415) );
  NANDN U366 ( .A(B[920]), .B(A[920]), .Z(n418) );
  AND U367 ( .A(n419), .B(n420), .Z(n417) );
  NAND U368 ( .A(n421), .B(n422), .Z(n420) );
  NANDN U369 ( .A(A[919]), .B(B[919]), .Z(n422) );
  AND U370 ( .A(n423), .B(n424), .Z(n421) );
  NANDN U371 ( .A(A[918]), .B(B[918]), .Z(n424) );
  NAND U372 ( .A(n425), .B(n426), .Z(n423) );
  NANDN U373 ( .A(B[918]), .B(A[918]), .Z(n426) );
  AND U374 ( .A(n427), .B(n428), .Z(n425) );
  NAND U375 ( .A(n429), .B(n430), .Z(n428) );
  NANDN U376 ( .A(A[917]), .B(B[917]), .Z(n430) );
  AND U377 ( .A(n431), .B(n432), .Z(n429) );
  NANDN U378 ( .A(A[916]), .B(B[916]), .Z(n432) );
  NAND U379 ( .A(n433), .B(n434), .Z(n431) );
  NANDN U380 ( .A(B[916]), .B(A[916]), .Z(n434) );
  AND U381 ( .A(n435), .B(n436), .Z(n433) );
  NAND U382 ( .A(n437), .B(n438), .Z(n436) );
  NANDN U383 ( .A(A[915]), .B(B[915]), .Z(n438) );
  AND U384 ( .A(n439), .B(n440), .Z(n437) );
  NANDN U385 ( .A(A[914]), .B(B[914]), .Z(n440) );
  NAND U386 ( .A(n441), .B(n442), .Z(n439) );
  NANDN U387 ( .A(B[914]), .B(A[914]), .Z(n442) );
  AND U388 ( .A(n443), .B(n444), .Z(n441) );
  NAND U389 ( .A(n445), .B(n446), .Z(n444) );
  NANDN U390 ( .A(A[913]), .B(B[913]), .Z(n446) );
  AND U391 ( .A(n447), .B(n448), .Z(n445) );
  NANDN U392 ( .A(A[912]), .B(B[912]), .Z(n448) );
  NAND U393 ( .A(n449), .B(n450), .Z(n447) );
  NANDN U394 ( .A(B[912]), .B(A[912]), .Z(n450) );
  AND U395 ( .A(n451), .B(n452), .Z(n449) );
  NAND U396 ( .A(n453), .B(n454), .Z(n452) );
  NANDN U397 ( .A(A[911]), .B(B[911]), .Z(n454) );
  AND U398 ( .A(n455), .B(n456), .Z(n453) );
  NANDN U399 ( .A(A[910]), .B(B[910]), .Z(n456) );
  NAND U400 ( .A(n457), .B(n458), .Z(n455) );
  NANDN U401 ( .A(B[910]), .B(A[910]), .Z(n458) );
  AND U402 ( .A(n459), .B(n460), .Z(n457) );
  NAND U403 ( .A(n461), .B(n462), .Z(n460) );
  NANDN U404 ( .A(A[909]), .B(B[909]), .Z(n462) );
  AND U405 ( .A(n463), .B(n464), .Z(n461) );
  NANDN U406 ( .A(A[908]), .B(B[908]), .Z(n464) );
  NAND U407 ( .A(n465), .B(n466), .Z(n463) );
  NANDN U408 ( .A(B[908]), .B(A[908]), .Z(n466) );
  AND U409 ( .A(n467), .B(n468), .Z(n465) );
  NAND U410 ( .A(n469), .B(n470), .Z(n468) );
  NANDN U411 ( .A(A[907]), .B(B[907]), .Z(n470) );
  AND U412 ( .A(n471), .B(n472), .Z(n469) );
  NANDN U413 ( .A(A[906]), .B(B[906]), .Z(n472) );
  NAND U414 ( .A(n473), .B(n474), .Z(n471) );
  NANDN U415 ( .A(B[906]), .B(A[906]), .Z(n474) );
  AND U416 ( .A(n475), .B(n476), .Z(n473) );
  NAND U417 ( .A(n477), .B(n478), .Z(n476) );
  NANDN U418 ( .A(A[905]), .B(B[905]), .Z(n478) );
  AND U419 ( .A(n479), .B(n480), .Z(n477) );
  NANDN U420 ( .A(A[904]), .B(B[904]), .Z(n480) );
  NAND U421 ( .A(n481), .B(n482), .Z(n479) );
  NANDN U422 ( .A(B[904]), .B(A[904]), .Z(n482) );
  AND U423 ( .A(n483), .B(n484), .Z(n481) );
  NAND U424 ( .A(n485), .B(n486), .Z(n484) );
  NANDN U425 ( .A(A[903]), .B(B[903]), .Z(n486) );
  AND U426 ( .A(n487), .B(n488), .Z(n485) );
  NANDN U427 ( .A(A[902]), .B(B[902]), .Z(n488) );
  NAND U428 ( .A(n489), .B(n490), .Z(n487) );
  NANDN U429 ( .A(B[902]), .B(A[902]), .Z(n490) );
  AND U430 ( .A(n491), .B(n492), .Z(n489) );
  NAND U431 ( .A(n493), .B(n494), .Z(n492) );
  NANDN U432 ( .A(A[901]), .B(B[901]), .Z(n494) );
  AND U433 ( .A(n495), .B(n496), .Z(n493) );
  NANDN U434 ( .A(A[900]), .B(B[900]), .Z(n496) );
  NAND U435 ( .A(n497), .B(n498), .Z(n495) );
  NANDN U436 ( .A(B[900]), .B(A[900]), .Z(n498) );
  AND U437 ( .A(n499), .B(n500), .Z(n497) );
  NAND U438 ( .A(n501), .B(n502), .Z(n500) );
  NANDN U439 ( .A(A[899]), .B(B[899]), .Z(n502) );
  AND U440 ( .A(n503), .B(n504), .Z(n501) );
  NANDN U441 ( .A(A[898]), .B(B[898]), .Z(n504) );
  NAND U442 ( .A(n505), .B(n506), .Z(n503) );
  NANDN U443 ( .A(B[898]), .B(A[898]), .Z(n506) );
  AND U444 ( .A(n507), .B(n508), .Z(n505) );
  NAND U445 ( .A(n509), .B(n510), .Z(n508) );
  NANDN U446 ( .A(A[897]), .B(B[897]), .Z(n510) );
  AND U447 ( .A(n511), .B(n512), .Z(n509) );
  NANDN U448 ( .A(A[896]), .B(B[896]), .Z(n512) );
  NAND U449 ( .A(n513), .B(n514), .Z(n511) );
  NANDN U450 ( .A(B[896]), .B(A[896]), .Z(n514) );
  AND U451 ( .A(n515), .B(n516), .Z(n513) );
  NAND U452 ( .A(n517), .B(n518), .Z(n516) );
  NANDN U453 ( .A(A[895]), .B(B[895]), .Z(n518) );
  AND U454 ( .A(n519), .B(n520), .Z(n517) );
  NANDN U455 ( .A(A[894]), .B(B[894]), .Z(n520) );
  NAND U456 ( .A(n521), .B(n522), .Z(n519) );
  NANDN U457 ( .A(B[894]), .B(A[894]), .Z(n522) );
  AND U458 ( .A(n523), .B(n524), .Z(n521) );
  NAND U459 ( .A(n525), .B(n526), .Z(n524) );
  NANDN U460 ( .A(A[893]), .B(B[893]), .Z(n526) );
  AND U461 ( .A(n527), .B(n528), .Z(n525) );
  NANDN U462 ( .A(A[892]), .B(B[892]), .Z(n528) );
  NAND U463 ( .A(n529), .B(n530), .Z(n527) );
  NANDN U464 ( .A(B[892]), .B(A[892]), .Z(n530) );
  AND U465 ( .A(n531), .B(n532), .Z(n529) );
  NAND U466 ( .A(n533), .B(n534), .Z(n532) );
  NANDN U467 ( .A(A[891]), .B(B[891]), .Z(n534) );
  AND U468 ( .A(n535), .B(n536), .Z(n533) );
  NANDN U469 ( .A(A[890]), .B(B[890]), .Z(n536) );
  NAND U470 ( .A(n537), .B(n538), .Z(n535) );
  NANDN U471 ( .A(B[890]), .B(A[890]), .Z(n538) );
  AND U472 ( .A(n539), .B(n540), .Z(n537) );
  NAND U473 ( .A(n541), .B(n542), .Z(n540) );
  NANDN U474 ( .A(A[889]), .B(B[889]), .Z(n542) );
  AND U475 ( .A(n543), .B(n544), .Z(n541) );
  NANDN U476 ( .A(A[888]), .B(B[888]), .Z(n544) );
  NAND U477 ( .A(n545), .B(n546), .Z(n543) );
  NANDN U478 ( .A(B[888]), .B(A[888]), .Z(n546) );
  AND U479 ( .A(n547), .B(n548), .Z(n545) );
  NAND U480 ( .A(n549), .B(n550), .Z(n548) );
  NANDN U481 ( .A(A[887]), .B(B[887]), .Z(n550) );
  AND U482 ( .A(n551), .B(n552), .Z(n549) );
  NANDN U483 ( .A(A[886]), .B(B[886]), .Z(n552) );
  NAND U484 ( .A(n553), .B(n554), .Z(n551) );
  NANDN U485 ( .A(B[886]), .B(A[886]), .Z(n554) );
  AND U486 ( .A(n555), .B(n556), .Z(n553) );
  NAND U487 ( .A(n557), .B(n558), .Z(n556) );
  NANDN U488 ( .A(A[885]), .B(B[885]), .Z(n558) );
  AND U489 ( .A(n559), .B(n560), .Z(n557) );
  NANDN U490 ( .A(A[884]), .B(B[884]), .Z(n560) );
  NAND U491 ( .A(n561), .B(n562), .Z(n559) );
  NANDN U492 ( .A(B[884]), .B(A[884]), .Z(n562) );
  AND U493 ( .A(n563), .B(n564), .Z(n561) );
  NAND U494 ( .A(n565), .B(n566), .Z(n564) );
  NANDN U495 ( .A(A[883]), .B(B[883]), .Z(n566) );
  AND U496 ( .A(n567), .B(n568), .Z(n565) );
  NANDN U497 ( .A(A[882]), .B(B[882]), .Z(n568) );
  NAND U498 ( .A(n569), .B(n570), .Z(n567) );
  NANDN U499 ( .A(B[882]), .B(A[882]), .Z(n570) );
  AND U500 ( .A(n571), .B(n572), .Z(n569) );
  NAND U501 ( .A(n573), .B(n574), .Z(n572) );
  NANDN U502 ( .A(A[881]), .B(B[881]), .Z(n574) );
  AND U503 ( .A(n575), .B(n576), .Z(n573) );
  NANDN U504 ( .A(A[880]), .B(B[880]), .Z(n576) );
  NAND U505 ( .A(n577), .B(n578), .Z(n575) );
  NANDN U506 ( .A(B[880]), .B(A[880]), .Z(n578) );
  AND U507 ( .A(n579), .B(n580), .Z(n577) );
  NAND U508 ( .A(n581), .B(n582), .Z(n580) );
  NANDN U509 ( .A(A[879]), .B(B[879]), .Z(n582) );
  AND U510 ( .A(n583), .B(n584), .Z(n581) );
  NANDN U511 ( .A(A[878]), .B(B[878]), .Z(n584) );
  NAND U512 ( .A(n585), .B(n586), .Z(n583) );
  NANDN U513 ( .A(B[878]), .B(A[878]), .Z(n586) );
  AND U514 ( .A(n587), .B(n588), .Z(n585) );
  NAND U515 ( .A(n589), .B(n590), .Z(n588) );
  NANDN U516 ( .A(A[877]), .B(B[877]), .Z(n590) );
  AND U517 ( .A(n591), .B(n592), .Z(n589) );
  NANDN U518 ( .A(A[876]), .B(B[876]), .Z(n592) );
  NAND U519 ( .A(n593), .B(n594), .Z(n591) );
  NANDN U520 ( .A(B[876]), .B(A[876]), .Z(n594) );
  AND U521 ( .A(n595), .B(n596), .Z(n593) );
  NAND U522 ( .A(n597), .B(n598), .Z(n596) );
  NANDN U523 ( .A(A[875]), .B(B[875]), .Z(n598) );
  AND U524 ( .A(n599), .B(n600), .Z(n597) );
  NANDN U525 ( .A(A[874]), .B(B[874]), .Z(n600) );
  NAND U526 ( .A(n601), .B(n602), .Z(n599) );
  NANDN U527 ( .A(B[874]), .B(A[874]), .Z(n602) );
  AND U528 ( .A(n603), .B(n604), .Z(n601) );
  NAND U529 ( .A(n605), .B(n606), .Z(n604) );
  NANDN U530 ( .A(A[873]), .B(B[873]), .Z(n606) );
  AND U531 ( .A(n607), .B(n608), .Z(n605) );
  NANDN U532 ( .A(A[872]), .B(B[872]), .Z(n608) );
  NAND U533 ( .A(n609), .B(n610), .Z(n607) );
  NANDN U534 ( .A(B[872]), .B(A[872]), .Z(n610) );
  AND U535 ( .A(n611), .B(n612), .Z(n609) );
  NAND U536 ( .A(n613), .B(n614), .Z(n612) );
  NANDN U537 ( .A(A[871]), .B(B[871]), .Z(n614) );
  AND U538 ( .A(n615), .B(n616), .Z(n613) );
  NANDN U539 ( .A(A[870]), .B(B[870]), .Z(n616) );
  NAND U540 ( .A(n617), .B(n618), .Z(n615) );
  NANDN U541 ( .A(B[870]), .B(A[870]), .Z(n618) );
  AND U542 ( .A(n619), .B(n620), .Z(n617) );
  NAND U543 ( .A(n621), .B(n622), .Z(n620) );
  NANDN U544 ( .A(A[869]), .B(B[869]), .Z(n622) );
  AND U545 ( .A(n623), .B(n624), .Z(n621) );
  NANDN U546 ( .A(A[868]), .B(B[868]), .Z(n624) );
  NAND U547 ( .A(n625), .B(n626), .Z(n623) );
  NANDN U548 ( .A(B[868]), .B(A[868]), .Z(n626) );
  AND U549 ( .A(n627), .B(n628), .Z(n625) );
  NAND U550 ( .A(n629), .B(n630), .Z(n628) );
  NANDN U551 ( .A(A[867]), .B(B[867]), .Z(n630) );
  AND U552 ( .A(n631), .B(n632), .Z(n629) );
  NANDN U553 ( .A(A[866]), .B(B[866]), .Z(n632) );
  NAND U554 ( .A(n633), .B(n634), .Z(n631) );
  NANDN U555 ( .A(B[866]), .B(A[866]), .Z(n634) );
  AND U556 ( .A(n635), .B(n636), .Z(n633) );
  NAND U557 ( .A(n637), .B(n638), .Z(n636) );
  NANDN U558 ( .A(A[865]), .B(B[865]), .Z(n638) );
  AND U559 ( .A(n639), .B(n640), .Z(n637) );
  NANDN U560 ( .A(A[864]), .B(B[864]), .Z(n640) );
  NAND U561 ( .A(n641), .B(n642), .Z(n639) );
  NANDN U562 ( .A(B[864]), .B(A[864]), .Z(n642) );
  AND U563 ( .A(n643), .B(n644), .Z(n641) );
  NAND U564 ( .A(n645), .B(n646), .Z(n644) );
  NANDN U565 ( .A(A[863]), .B(B[863]), .Z(n646) );
  AND U566 ( .A(n647), .B(n648), .Z(n645) );
  NANDN U567 ( .A(A[862]), .B(B[862]), .Z(n648) );
  NAND U568 ( .A(n649), .B(n650), .Z(n647) );
  NANDN U569 ( .A(B[862]), .B(A[862]), .Z(n650) );
  AND U570 ( .A(n651), .B(n652), .Z(n649) );
  NAND U571 ( .A(n653), .B(n654), .Z(n652) );
  NANDN U572 ( .A(A[861]), .B(B[861]), .Z(n654) );
  AND U573 ( .A(n655), .B(n656), .Z(n653) );
  NANDN U574 ( .A(A[860]), .B(B[860]), .Z(n656) );
  NAND U575 ( .A(n657), .B(n658), .Z(n655) );
  NANDN U576 ( .A(B[860]), .B(A[860]), .Z(n658) );
  AND U577 ( .A(n659), .B(n660), .Z(n657) );
  NAND U578 ( .A(n661), .B(n662), .Z(n660) );
  NANDN U579 ( .A(A[859]), .B(B[859]), .Z(n662) );
  AND U580 ( .A(n663), .B(n664), .Z(n661) );
  NANDN U581 ( .A(A[858]), .B(B[858]), .Z(n664) );
  NAND U582 ( .A(n665), .B(n666), .Z(n663) );
  NANDN U583 ( .A(B[858]), .B(A[858]), .Z(n666) );
  AND U584 ( .A(n667), .B(n668), .Z(n665) );
  NAND U585 ( .A(n669), .B(n670), .Z(n668) );
  NANDN U586 ( .A(A[857]), .B(B[857]), .Z(n670) );
  AND U587 ( .A(n671), .B(n672), .Z(n669) );
  NANDN U588 ( .A(A[856]), .B(B[856]), .Z(n672) );
  NAND U589 ( .A(n673), .B(n674), .Z(n671) );
  NANDN U590 ( .A(B[856]), .B(A[856]), .Z(n674) );
  AND U591 ( .A(n675), .B(n676), .Z(n673) );
  NAND U592 ( .A(n677), .B(n678), .Z(n676) );
  NANDN U593 ( .A(A[855]), .B(B[855]), .Z(n678) );
  AND U594 ( .A(n679), .B(n680), .Z(n677) );
  NANDN U595 ( .A(A[854]), .B(B[854]), .Z(n680) );
  NAND U596 ( .A(n681), .B(n682), .Z(n679) );
  NANDN U597 ( .A(B[854]), .B(A[854]), .Z(n682) );
  AND U598 ( .A(n683), .B(n684), .Z(n681) );
  NAND U599 ( .A(n685), .B(n686), .Z(n684) );
  NANDN U600 ( .A(A[853]), .B(B[853]), .Z(n686) );
  AND U601 ( .A(n687), .B(n688), .Z(n685) );
  NANDN U602 ( .A(A[852]), .B(B[852]), .Z(n688) );
  NAND U603 ( .A(n689), .B(n690), .Z(n687) );
  NANDN U604 ( .A(B[852]), .B(A[852]), .Z(n690) );
  AND U605 ( .A(n691), .B(n692), .Z(n689) );
  NAND U606 ( .A(n693), .B(n694), .Z(n692) );
  NANDN U607 ( .A(A[851]), .B(B[851]), .Z(n694) );
  AND U608 ( .A(n695), .B(n696), .Z(n693) );
  NANDN U609 ( .A(A[850]), .B(B[850]), .Z(n696) );
  NAND U610 ( .A(n697), .B(n698), .Z(n695) );
  NANDN U611 ( .A(B[850]), .B(A[850]), .Z(n698) );
  AND U612 ( .A(n699), .B(n700), .Z(n697) );
  NAND U613 ( .A(n701), .B(n702), .Z(n700) );
  NANDN U614 ( .A(A[849]), .B(B[849]), .Z(n702) );
  AND U615 ( .A(n703), .B(n704), .Z(n701) );
  NANDN U616 ( .A(A[848]), .B(B[848]), .Z(n704) );
  NAND U617 ( .A(n705), .B(n706), .Z(n703) );
  NANDN U618 ( .A(B[848]), .B(A[848]), .Z(n706) );
  AND U619 ( .A(n707), .B(n708), .Z(n705) );
  NAND U620 ( .A(n709), .B(n710), .Z(n708) );
  NANDN U621 ( .A(A[847]), .B(B[847]), .Z(n710) );
  AND U622 ( .A(n711), .B(n712), .Z(n709) );
  NANDN U623 ( .A(A[846]), .B(B[846]), .Z(n712) );
  NAND U624 ( .A(n713), .B(n714), .Z(n711) );
  NANDN U625 ( .A(B[846]), .B(A[846]), .Z(n714) );
  AND U626 ( .A(n715), .B(n716), .Z(n713) );
  NAND U627 ( .A(n717), .B(n718), .Z(n716) );
  NANDN U628 ( .A(A[845]), .B(B[845]), .Z(n718) );
  AND U629 ( .A(n719), .B(n720), .Z(n717) );
  NANDN U630 ( .A(A[844]), .B(B[844]), .Z(n720) );
  NAND U631 ( .A(n721), .B(n722), .Z(n719) );
  NANDN U632 ( .A(B[844]), .B(A[844]), .Z(n722) );
  AND U633 ( .A(n723), .B(n724), .Z(n721) );
  NAND U634 ( .A(n725), .B(n726), .Z(n724) );
  NANDN U635 ( .A(A[843]), .B(B[843]), .Z(n726) );
  AND U636 ( .A(n727), .B(n728), .Z(n725) );
  NANDN U637 ( .A(A[842]), .B(B[842]), .Z(n728) );
  NAND U638 ( .A(n729), .B(n730), .Z(n727) );
  NANDN U639 ( .A(B[842]), .B(A[842]), .Z(n730) );
  AND U640 ( .A(n731), .B(n732), .Z(n729) );
  NAND U641 ( .A(n733), .B(n734), .Z(n732) );
  NANDN U642 ( .A(A[841]), .B(B[841]), .Z(n734) );
  AND U643 ( .A(n735), .B(n736), .Z(n733) );
  NANDN U644 ( .A(A[840]), .B(B[840]), .Z(n736) );
  NAND U645 ( .A(n737), .B(n738), .Z(n735) );
  NANDN U646 ( .A(B[840]), .B(A[840]), .Z(n738) );
  AND U647 ( .A(n739), .B(n740), .Z(n737) );
  NAND U648 ( .A(n741), .B(n742), .Z(n740) );
  NANDN U649 ( .A(A[839]), .B(B[839]), .Z(n742) );
  AND U650 ( .A(n743), .B(n744), .Z(n741) );
  NANDN U651 ( .A(A[838]), .B(B[838]), .Z(n744) );
  NAND U652 ( .A(n745), .B(n746), .Z(n743) );
  NANDN U653 ( .A(B[838]), .B(A[838]), .Z(n746) );
  AND U654 ( .A(n747), .B(n748), .Z(n745) );
  NAND U655 ( .A(n749), .B(n750), .Z(n748) );
  NANDN U656 ( .A(A[837]), .B(B[837]), .Z(n750) );
  AND U657 ( .A(n751), .B(n752), .Z(n749) );
  NANDN U658 ( .A(A[836]), .B(B[836]), .Z(n752) );
  NAND U659 ( .A(n753), .B(n754), .Z(n751) );
  NANDN U660 ( .A(B[836]), .B(A[836]), .Z(n754) );
  AND U661 ( .A(n755), .B(n756), .Z(n753) );
  NAND U662 ( .A(n757), .B(n758), .Z(n756) );
  NANDN U663 ( .A(A[835]), .B(B[835]), .Z(n758) );
  AND U664 ( .A(n759), .B(n760), .Z(n757) );
  NANDN U665 ( .A(A[834]), .B(B[834]), .Z(n760) );
  NAND U666 ( .A(n761), .B(n762), .Z(n759) );
  NANDN U667 ( .A(B[834]), .B(A[834]), .Z(n762) );
  AND U668 ( .A(n763), .B(n764), .Z(n761) );
  NAND U669 ( .A(n765), .B(n766), .Z(n764) );
  NANDN U670 ( .A(A[833]), .B(B[833]), .Z(n766) );
  AND U671 ( .A(n767), .B(n768), .Z(n765) );
  NANDN U672 ( .A(A[832]), .B(B[832]), .Z(n768) );
  NAND U673 ( .A(n769), .B(n770), .Z(n767) );
  NANDN U674 ( .A(B[832]), .B(A[832]), .Z(n770) );
  AND U675 ( .A(n771), .B(n772), .Z(n769) );
  NAND U676 ( .A(n773), .B(n774), .Z(n772) );
  NANDN U677 ( .A(A[831]), .B(B[831]), .Z(n774) );
  AND U678 ( .A(n775), .B(n776), .Z(n773) );
  NANDN U679 ( .A(A[830]), .B(B[830]), .Z(n776) );
  NAND U680 ( .A(n777), .B(n778), .Z(n775) );
  NANDN U681 ( .A(B[830]), .B(A[830]), .Z(n778) );
  AND U682 ( .A(n779), .B(n780), .Z(n777) );
  NAND U683 ( .A(n781), .B(n782), .Z(n780) );
  NANDN U684 ( .A(A[829]), .B(B[829]), .Z(n782) );
  AND U685 ( .A(n783), .B(n784), .Z(n781) );
  NANDN U686 ( .A(A[828]), .B(B[828]), .Z(n784) );
  NAND U687 ( .A(n785), .B(n786), .Z(n783) );
  NANDN U688 ( .A(B[828]), .B(A[828]), .Z(n786) );
  AND U689 ( .A(n787), .B(n788), .Z(n785) );
  NAND U690 ( .A(n789), .B(n790), .Z(n788) );
  NANDN U691 ( .A(A[827]), .B(B[827]), .Z(n790) );
  AND U692 ( .A(n791), .B(n792), .Z(n789) );
  NANDN U693 ( .A(A[826]), .B(B[826]), .Z(n792) );
  NAND U694 ( .A(n793), .B(n794), .Z(n791) );
  NANDN U695 ( .A(B[826]), .B(A[826]), .Z(n794) );
  AND U696 ( .A(n795), .B(n796), .Z(n793) );
  NAND U697 ( .A(n797), .B(n798), .Z(n796) );
  NANDN U698 ( .A(A[825]), .B(B[825]), .Z(n798) );
  AND U699 ( .A(n799), .B(n800), .Z(n797) );
  NANDN U700 ( .A(A[824]), .B(B[824]), .Z(n800) );
  NAND U701 ( .A(n801), .B(n802), .Z(n799) );
  NANDN U702 ( .A(B[824]), .B(A[824]), .Z(n802) );
  AND U703 ( .A(n803), .B(n804), .Z(n801) );
  NAND U704 ( .A(n805), .B(n806), .Z(n804) );
  NANDN U705 ( .A(A[823]), .B(B[823]), .Z(n806) );
  AND U706 ( .A(n807), .B(n808), .Z(n805) );
  NANDN U707 ( .A(A[822]), .B(B[822]), .Z(n808) );
  NAND U708 ( .A(n809), .B(n810), .Z(n807) );
  NANDN U709 ( .A(B[822]), .B(A[822]), .Z(n810) );
  AND U710 ( .A(n811), .B(n812), .Z(n809) );
  NAND U711 ( .A(n813), .B(n814), .Z(n812) );
  NANDN U712 ( .A(A[821]), .B(B[821]), .Z(n814) );
  AND U713 ( .A(n815), .B(n816), .Z(n813) );
  NANDN U714 ( .A(A[820]), .B(B[820]), .Z(n816) );
  NAND U715 ( .A(n817), .B(n818), .Z(n815) );
  NANDN U716 ( .A(B[820]), .B(A[820]), .Z(n818) );
  AND U717 ( .A(n819), .B(n820), .Z(n817) );
  NAND U718 ( .A(n821), .B(n822), .Z(n820) );
  NANDN U719 ( .A(A[819]), .B(B[819]), .Z(n822) );
  AND U720 ( .A(n823), .B(n824), .Z(n821) );
  NANDN U721 ( .A(A[818]), .B(B[818]), .Z(n824) );
  NAND U722 ( .A(n825), .B(n826), .Z(n823) );
  NANDN U723 ( .A(B[818]), .B(A[818]), .Z(n826) );
  AND U724 ( .A(n827), .B(n828), .Z(n825) );
  NAND U725 ( .A(n829), .B(n830), .Z(n828) );
  NANDN U726 ( .A(A[817]), .B(B[817]), .Z(n830) );
  AND U727 ( .A(n831), .B(n832), .Z(n829) );
  NANDN U728 ( .A(A[816]), .B(B[816]), .Z(n832) );
  NAND U729 ( .A(n833), .B(n834), .Z(n831) );
  NANDN U730 ( .A(B[816]), .B(A[816]), .Z(n834) );
  AND U731 ( .A(n835), .B(n836), .Z(n833) );
  NAND U732 ( .A(n837), .B(n838), .Z(n836) );
  NANDN U733 ( .A(A[815]), .B(B[815]), .Z(n838) );
  AND U734 ( .A(n839), .B(n840), .Z(n837) );
  NANDN U735 ( .A(A[814]), .B(B[814]), .Z(n840) );
  NAND U736 ( .A(n841), .B(n842), .Z(n839) );
  NANDN U737 ( .A(B[814]), .B(A[814]), .Z(n842) );
  AND U738 ( .A(n843), .B(n844), .Z(n841) );
  NAND U739 ( .A(n845), .B(n846), .Z(n844) );
  NANDN U740 ( .A(A[813]), .B(B[813]), .Z(n846) );
  AND U741 ( .A(n847), .B(n848), .Z(n845) );
  NANDN U742 ( .A(A[812]), .B(B[812]), .Z(n848) );
  NAND U743 ( .A(n849), .B(n850), .Z(n847) );
  NANDN U744 ( .A(B[812]), .B(A[812]), .Z(n850) );
  AND U745 ( .A(n851), .B(n852), .Z(n849) );
  NAND U746 ( .A(n853), .B(n854), .Z(n852) );
  NANDN U747 ( .A(A[811]), .B(B[811]), .Z(n854) );
  AND U748 ( .A(n855), .B(n856), .Z(n853) );
  NANDN U749 ( .A(A[810]), .B(B[810]), .Z(n856) );
  NAND U750 ( .A(n857), .B(n858), .Z(n855) );
  NANDN U751 ( .A(B[810]), .B(A[810]), .Z(n858) );
  AND U752 ( .A(n859), .B(n860), .Z(n857) );
  NAND U753 ( .A(n861), .B(n862), .Z(n860) );
  NANDN U754 ( .A(A[809]), .B(B[809]), .Z(n862) );
  AND U755 ( .A(n863), .B(n864), .Z(n861) );
  NANDN U756 ( .A(A[808]), .B(B[808]), .Z(n864) );
  NAND U757 ( .A(n865), .B(n866), .Z(n863) );
  NANDN U758 ( .A(B[808]), .B(A[808]), .Z(n866) );
  AND U759 ( .A(n867), .B(n868), .Z(n865) );
  NAND U760 ( .A(n869), .B(n870), .Z(n868) );
  NANDN U761 ( .A(A[807]), .B(B[807]), .Z(n870) );
  AND U762 ( .A(n871), .B(n872), .Z(n869) );
  NANDN U763 ( .A(A[806]), .B(B[806]), .Z(n872) );
  NAND U764 ( .A(n873), .B(n874), .Z(n871) );
  NANDN U765 ( .A(B[806]), .B(A[806]), .Z(n874) );
  AND U766 ( .A(n875), .B(n876), .Z(n873) );
  NAND U767 ( .A(n877), .B(n878), .Z(n876) );
  NANDN U768 ( .A(A[805]), .B(B[805]), .Z(n878) );
  AND U769 ( .A(n879), .B(n880), .Z(n877) );
  NANDN U770 ( .A(A[804]), .B(B[804]), .Z(n880) );
  NAND U771 ( .A(n881), .B(n882), .Z(n879) );
  NANDN U772 ( .A(B[804]), .B(A[804]), .Z(n882) );
  AND U773 ( .A(n883), .B(n884), .Z(n881) );
  NAND U774 ( .A(n885), .B(n886), .Z(n884) );
  NANDN U775 ( .A(A[803]), .B(B[803]), .Z(n886) );
  AND U776 ( .A(n887), .B(n888), .Z(n885) );
  NANDN U777 ( .A(A[802]), .B(B[802]), .Z(n888) );
  NAND U778 ( .A(n889), .B(n890), .Z(n887) );
  NANDN U779 ( .A(B[802]), .B(A[802]), .Z(n890) );
  AND U780 ( .A(n891), .B(n892), .Z(n889) );
  NAND U781 ( .A(n893), .B(n894), .Z(n892) );
  NANDN U782 ( .A(A[801]), .B(B[801]), .Z(n894) );
  AND U783 ( .A(n895), .B(n896), .Z(n893) );
  NANDN U784 ( .A(A[800]), .B(B[800]), .Z(n896) );
  NAND U785 ( .A(n897), .B(n898), .Z(n895) );
  NANDN U786 ( .A(B[800]), .B(A[800]), .Z(n898) );
  AND U787 ( .A(n899), .B(n900), .Z(n897) );
  NAND U788 ( .A(n901), .B(n902), .Z(n900) );
  NANDN U789 ( .A(A[799]), .B(B[799]), .Z(n902) );
  AND U790 ( .A(n903), .B(n904), .Z(n901) );
  NANDN U791 ( .A(A[798]), .B(B[798]), .Z(n904) );
  NAND U792 ( .A(n905), .B(n906), .Z(n903) );
  NANDN U793 ( .A(B[798]), .B(A[798]), .Z(n906) );
  AND U794 ( .A(n907), .B(n908), .Z(n905) );
  NAND U795 ( .A(n909), .B(n910), .Z(n908) );
  NANDN U796 ( .A(A[797]), .B(B[797]), .Z(n910) );
  AND U797 ( .A(n911), .B(n912), .Z(n909) );
  NANDN U798 ( .A(A[796]), .B(B[796]), .Z(n912) );
  NAND U799 ( .A(n913), .B(n914), .Z(n911) );
  NANDN U800 ( .A(B[796]), .B(A[796]), .Z(n914) );
  AND U801 ( .A(n915), .B(n916), .Z(n913) );
  NAND U802 ( .A(n917), .B(n918), .Z(n916) );
  NANDN U803 ( .A(A[795]), .B(B[795]), .Z(n918) );
  AND U804 ( .A(n919), .B(n920), .Z(n917) );
  NANDN U805 ( .A(A[794]), .B(B[794]), .Z(n920) );
  NAND U806 ( .A(n921), .B(n922), .Z(n919) );
  NANDN U807 ( .A(B[794]), .B(A[794]), .Z(n922) );
  AND U808 ( .A(n923), .B(n924), .Z(n921) );
  NAND U809 ( .A(n925), .B(n926), .Z(n924) );
  NANDN U810 ( .A(A[793]), .B(B[793]), .Z(n926) );
  AND U811 ( .A(n927), .B(n928), .Z(n925) );
  NANDN U812 ( .A(A[792]), .B(B[792]), .Z(n928) );
  NAND U813 ( .A(n929), .B(n930), .Z(n927) );
  NANDN U814 ( .A(B[792]), .B(A[792]), .Z(n930) );
  AND U815 ( .A(n931), .B(n932), .Z(n929) );
  NAND U816 ( .A(n933), .B(n934), .Z(n932) );
  NANDN U817 ( .A(A[791]), .B(B[791]), .Z(n934) );
  AND U818 ( .A(n935), .B(n936), .Z(n933) );
  NANDN U819 ( .A(A[790]), .B(B[790]), .Z(n936) );
  NAND U820 ( .A(n937), .B(n938), .Z(n935) );
  NANDN U821 ( .A(B[790]), .B(A[790]), .Z(n938) );
  AND U822 ( .A(n939), .B(n940), .Z(n937) );
  NAND U823 ( .A(n941), .B(n942), .Z(n940) );
  NANDN U824 ( .A(A[789]), .B(B[789]), .Z(n942) );
  AND U825 ( .A(n943), .B(n944), .Z(n941) );
  NANDN U826 ( .A(A[788]), .B(B[788]), .Z(n944) );
  NAND U827 ( .A(n945), .B(n946), .Z(n943) );
  NANDN U828 ( .A(B[788]), .B(A[788]), .Z(n946) );
  AND U829 ( .A(n947), .B(n948), .Z(n945) );
  NAND U830 ( .A(n949), .B(n950), .Z(n948) );
  NANDN U831 ( .A(A[787]), .B(B[787]), .Z(n950) );
  AND U832 ( .A(n951), .B(n952), .Z(n949) );
  NANDN U833 ( .A(A[786]), .B(B[786]), .Z(n952) );
  NAND U834 ( .A(n953), .B(n954), .Z(n951) );
  NANDN U835 ( .A(B[786]), .B(A[786]), .Z(n954) );
  AND U836 ( .A(n955), .B(n956), .Z(n953) );
  NAND U837 ( .A(n957), .B(n958), .Z(n956) );
  NANDN U838 ( .A(A[785]), .B(B[785]), .Z(n958) );
  AND U839 ( .A(n959), .B(n960), .Z(n957) );
  NANDN U840 ( .A(A[784]), .B(B[784]), .Z(n960) );
  NAND U841 ( .A(n961), .B(n962), .Z(n959) );
  NANDN U842 ( .A(B[784]), .B(A[784]), .Z(n962) );
  AND U843 ( .A(n963), .B(n964), .Z(n961) );
  NAND U844 ( .A(n965), .B(n966), .Z(n964) );
  NANDN U845 ( .A(A[783]), .B(B[783]), .Z(n966) );
  AND U846 ( .A(n967), .B(n968), .Z(n965) );
  NANDN U847 ( .A(A[782]), .B(B[782]), .Z(n968) );
  NAND U848 ( .A(n969), .B(n970), .Z(n967) );
  NANDN U849 ( .A(B[782]), .B(A[782]), .Z(n970) );
  AND U850 ( .A(n971), .B(n972), .Z(n969) );
  NAND U851 ( .A(n973), .B(n974), .Z(n972) );
  NANDN U852 ( .A(A[781]), .B(B[781]), .Z(n974) );
  AND U853 ( .A(n975), .B(n976), .Z(n973) );
  NANDN U854 ( .A(A[780]), .B(B[780]), .Z(n976) );
  NAND U855 ( .A(n977), .B(n978), .Z(n975) );
  NANDN U856 ( .A(B[780]), .B(A[780]), .Z(n978) );
  AND U857 ( .A(n979), .B(n980), .Z(n977) );
  NAND U858 ( .A(n981), .B(n982), .Z(n980) );
  NANDN U859 ( .A(A[779]), .B(B[779]), .Z(n982) );
  AND U860 ( .A(n983), .B(n984), .Z(n981) );
  NANDN U861 ( .A(A[778]), .B(B[778]), .Z(n984) );
  NAND U862 ( .A(n985), .B(n986), .Z(n983) );
  NANDN U863 ( .A(B[778]), .B(A[778]), .Z(n986) );
  AND U864 ( .A(n987), .B(n988), .Z(n985) );
  NAND U865 ( .A(n989), .B(n990), .Z(n988) );
  NANDN U866 ( .A(A[777]), .B(B[777]), .Z(n990) );
  AND U867 ( .A(n991), .B(n992), .Z(n989) );
  NANDN U868 ( .A(A[776]), .B(B[776]), .Z(n992) );
  NAND U869 ( .A(n993), .B(n994), .Z(n991) );
  NANDN U870 ( .A(B[776]), .B(A[776]), .Z(n994) );
  AND U871 ( .A(n995), .B(n996), .Z(n993) );
  NAND U872 ( .A(n997), .B(n998), .Z(n996) );
  NANDN U873 ( .A(A[775]), .B(B[775]), .Z(n998) );
  AND U874 ( .A(n999), .B(n1000), .Z(n997) );
  NANDN U875 ( .A(A[774]), .B(B[774]), .Z(n1000) );
  NAND U876 ( .A(n1001), .B(n1002), .Z(n999) );
  NANDN U877 ( .A(B[774]), .B(A[774]), .Z(n1002) );
  AND U878 ( .A(n1003), .B(n1004), .Z(n1001) );
  NAND U879 ( .A(n1005), .B(n1006), .Z(n1004) );
  NANDN U880 ( .A(A[773]), .B(B[773]), .Z(n1006) );
  AND U881 ( .A(n1007), .B(n1008), .Z(n1005) );
  NANDN U882 ( .A(A[772]), .B(B[772]), .Z(n1008) );
  NAND U883 ( .A(n1009), .B(n1010), .Z(n1007) );
  NANDN U884 ( .A(B[772]), .B(A[772]), .Z(n1010) );
  AND U885 ( .A(n1011), .B(n1012), .Z(n1009) );
  NAND U886 ( .A(n1013), .B(n1014), .Z(n1012) );
  NANDN U887 ( .A(A[771]), .B(B[771]), .Z(n1014) );
  AND U888 ( .A(n1015), .B(n1016), .Z(n1013) );
  NANDN U889 ( .A(A[770]), .B(B[770]), .Z(n1016) );
  NAND U890 ( .A(n1017), .B(n1018), .Z(n1015) );
  NANDN U891 ( .A(B[770]), .B(A[770]), .Z(n1018) );
  AND U892 ( .A(n1019), .B(n1020), .Z(n1017) );
  NAND U893 ( .A(n1021), .B(n1022), .Z(n1020) );
  NANDN U894 ( .A(A[769]), .B(B[769]), .Z(n1022) );
  AND U895 ( .A(n1023), .B(n1024), .Z(n1021) );
  NANDN U896 ( .A(A[768]), .B(B[768]), .Z(n1024) );
  NAND U897 ( .A(n1025), .B(n1026), .Z(n1023) );
  NANDN U898 ( .A(B[768]), .B(A[768]), .Z(n1026) );
  AND U899 ( .A(n1027), .B(n1028), .Z(n1025) );
  NAND U900 ( .A(n1029), .B(n1030), .Z(n1028) );
  NANDN U901 ( .A(A[767]), .B(B[767]), .Z(n1030) );
  AND U902 ( .A(n1031), .B(n1032), .Z(n1029) );
  NANDN U903 ( .A(A[766]), .B(B[766]), .Z(n1032) );
  NAND U904 ( .A(n1033), .B(n1034), .Z(n1031) );
  NANDN U905 ( .A(B[766]), .B(A[766]), .Z(n1034) );
  AND U906 ( .A(n1035), .B(n1036), .Z(n1033) );
  NAND U907 ( .A(n1037), .B(n1038), .Z(n1036) );
  NANDN U908 ( .A(A[765]), .B(B[765]), .Z(n1038) );
  AND U909 ( .A(n1039), .B(n1040), .Z(n1037) );
  NANDN U910 ( .A(A[764]), .B(B[764]), .Z(n1040) );
  NAND U911 ( .A(n1041), .B(n1042), .Z(n1039) );
  NANDN U912 ( .A(B[764]), .B(A[764]), .Z(n1042) );
  AND U913 ( .A(n1043), .B(n1044), .Z(n1041) );
  NAND U914 ( .A(n1045), .B(n1046), .Z(n1044) );
  NANDN U915 ( .A(A[763]), .B(B[763]), .Z(n1046) );
  AND U916 ( .A(n1047), .B(n1048), .Z(n1045) );
  NANDN U917 ( .A(A[762]), .B(B[762]), .Z(n1048) );
  NAND U918 ( .A(n1049), .B(n1050), .Z(n1047) );
  NANDN U919 ( .A(B[762]), .B(A[762]), .Z(n1050) );
  AND U920 ( .A(n1051), .B(n1052), .Z(n1049) );
  NAND U921 ( .A(n1053), .B(n1054), .Z(n1052) );
  NANDN U922 ( .A(A[761]), .B(B[761]), .Z(n1054) );
  AND U923 ( .A(n1055), .B(n1056), .Z(n1053) );
  NANDN U924 ( .A(A[760]), .B(B[760]), .Z(n1056) );
  NAND U925 ( .A(n1057), .B(n1058), .Z(n1055) );
  NANDN U926 ( .A(B[760]), .B(A[760]), .Z(n1058) );
  AND U927 ( .A(n1059), .B(n1060), .Z(n1057) );
  NAND U928 ( .A(n1061), .B(n1062), .Z(n1060) );
  NANDN U929 ( .A(A[759]), .B(B[759]), .Z(n1062) );
  AND U930 ( .A(n1063), .B(n1064), .Z(n1061) );
  NANDN U931 ( .A(A[758]), .B(B[758]), .Z(n1064) );
  NAND U932 ( .A(n1065), .B(n1066), .Z(n1063) );
  NANDN U933 ( .A(B[758]), .B(A[758]), .Z(n1066) );
  AND U934 ( .A(n1067), .B(n1068), .Z(n1065) );
  NAND U935 ( .A(n1069), .B(n1070), .Z(n1068) );
  NANDN U936 ( .A(A[757]), .B(B[757]), .Z(n1070) );
  AND U937 ( .A(n1071), .B(n1072), .Z(n1069) );
  NANDN U938 ( .A(A[756]), .B(B[756]), .Z(n1072) );
  NAND U939 ( .A(n1073), .B(n1074), .Z(n1071) );
  NANDN U940 ( .A(B[756]), .B(A[756]), .Z(n1074) );
  AND U941 ( .A(n1075), .B(n1076), .Z(n1073) );
  NAND U942 ( .A(n1077), .B(n1078), .Z(n1076) );
  NANDN U943 ( .A(A[755]), .B(B[755]), .Z(n1078) );
  AND U944 ( .A(n1079), .B(n1080), .Z(n1077) );
  NANDN U945 ( .A(A[754]), .B(B[754]), .Z(n1080) );
  NAND U946 ( .A(n1081), .B(n1082), .Z(n1079) );
  NANDN U947 ( .A(B[754]), .B(A[754]), .Z(n1082) );
  AND U948 ( .A(n1083), .B(n1084), .Z(n1081) );
  NAND U949 ( .A(n1085), .B(n1086), .Z(n1084) );
  NANDN U950 ( .A(A[753]), .B(B[753]), .Z(n1086) );
  AND U951 ( .A(n1087), .B(n1088), .Z(n1085) );
  NANDN U952 ( .A(A[752]), .B(B[752]), .Z(n1088) );
  NAND U953 ( .A(n1089), .B(n1090), .Z(n1087) );
  NANDN U954 ( .A(B[752]), .B(A[752]), .Z(n1090) );
  AND U955 ( .A(n1091), .B(n1092), .Z(n1089) );
  NAND U956 ( .A(n1093), .B(n1094), .Z(n1092) );
  NANDN U957 ( .A(A[751]), .B(B[751]), .Z(n1094) );
  AND U958 ( .A(n1095), .B(n1096), .Z(n1093) );
  NANDN U959 ( .A(A[750]), .B(B[750]), .Z(n1096) );
  NAND U960 ( .A(n1097), .B(n1098), .Z(n1095) );
  NANDN U961 ( .A(B[750]), .B(A[750]), .Z(n1098) );
  AND U962 ( .A(n1099), .B(n1100), .Z(n1097) );
  NAND U963 ( .A(n1101), .B(n1102), .Z(n1100) );
  NANDN U964 ( .A(A[749]), .B(B[749]), .Z(n1102) );
  AND U965 ( .A(n1103), .B(n1104), .Z(n1101) );
  NANDN U966 ( .A(A[748]), .B(B[748]), .Z(n1104) );
  NAND U967 ( .A(n1105), .B(n1106), .Z(n1103) );
  NANDN U968 ( .A(B[748]), .B(A[748]), .Z(n1106) );
  AND U969 ( .A(n1107), .B(n1108), .Z(n1105) );
  NAND U970 ( .A(n1109), .B(n1110), .Z(n1108) );
  NANDN U971 ( .A(A[747]), .B(B[747]), .Z(n1110) );
  AND U972 ( .A(n1111), .B(n1112), .Z(n1109) );
  NANDN U973 ( .A(A[746]), .B(B[746]), .Z(n1112) );
  NAND U974 ( .A(n1113), .B(n1114), .Z(n1111) );
  NANDN U975 ( .A(B[746]), .B(A[746]), .Z(n1114) );
  AND U976 ( .A(n1115), .B(n1116), .Z(n1113) );
  NAND U977 ( .A(n1117), .B(n1118), .Z(n1116) );
  NANDN U978 ( .A(A[745]), .B(B[745]), .Z(n1118) );
  AND U979 ( .A(n1119), .B(n1120), .Z(n1117) );
  NANDN U980 ( .A(A[744]), .B(B[744]), .Z(n1120) );
  NAND U981 ( .A(n1121), .B(n1122), .Z(n1119) );
  NANDN U982 ( .A(B[744]), .B(A[744]), .Z(n1122) );
  AND U983 ( .A(n1123), .B(n1124), .Z(n1121) );
  NAND U984 ( .A(n1125), .B(n1126), .Z(n1124) );
  NANDN U985 ( .A(A[743]), .B(B[743]), .Z(n1126) );
  AND U986 ( .A(n1127), .B(n1128), .Z(n1125) );
  NANDN U987 ( .A(A[742]), .B(B[742]), .Z(n1128) );
  NAND U988 ( .A(n1129), .B(n1130), .Z(n1127) );
  NANDN U989 ( .A(B[742]), .B(A[742]), .Z(n1130) );
  AND U990 ( .A(n1131), .B(n1132), .Z(n1129) );
  NAND U991 ( .A(n1133), .B(n1134), .Z(n1132) );
  NANDN U992 ( .A(A[741]), .B(B[741]), .Z(n1134) );
  AND U993 ( .A(n1135), .B(n1136), .Z(n1133) );
  NANDN U994 ( .A(A[740]), .B(B[740]), .Z(n1136) );
  NAND U995 ( .A(n1137), .B(n1138), .Z(n1135) );
  NANDN U996 ( .A(B[740]), .B(A[740]), .Z(n1138) );
  AND U997 ( .A(n1139), .B(n1140), .Z(n1137) );
  NAND U998 ( .A(n1141), .B(n1142), .Z(n1140) );
  NANDN U999 ( .A(A[739]), .B(B[739]), .Z(n1142) );
  AND U1000 ( .A(n1143), .B(n1144), .Z(n1141) );
  NANDN U1001 ( .A(A[738]), .B(B[738]), .Z(n1144) );
  NAND U1002 ( .A(n1145), .B(n1146), .Z(n1143) );
  NANDN U1003 ( .A(B[738]), .B(A[738]), .Z(n1146) );
  AND U1004 ( .A(n1147), .B(n1148), .Z(n1145) );
  NAND U1005 ( .A(n1149), .B(n1150), .Z(n1148) );
  NANDN U1006 ( .A(A[737]), .B(B[737]), .Z(n1150) );
  AND U1007 ( .A(n1151), .B(n1152), .Z(n1149) );
  NANDN U1008 ( .A(A[736]), .B(B[736]), .Z(n1152) );
  NAND U1009 ( .A(n1153), .B(n1154), .Z(n1151) );
  NANDN U1010 ( .A(B[736]), .B(A[736]), .Z(n1154) );
  AND U1011 ( .A(n1155), .B(n1156), .Z(n1153) );
  NAND U1012 ( .A(n1157), .B(n1158), .Z(n1156) );
  NANDN U1013 ( .A(A[735]), .B(B[735]), .Z(n1158) );
  AND U1014 ( .A(n1159), .B(n1160), .Z(n1157) );
  NANDN U1015 ( .A(A[734]), .B(B[734]), .Z(n1160) );
  NAND U1016 ( .A(n1161), .B(n1162), .Z(n1159) );
  NANDN U1017 ( .A(B[734]), .B(A[734]), .Z(n1162) );
  AND U1018 ( .A(n1163), .B(n1164), .Z(n1161) );
  NAND U1019 ( .A(n1165), .B(n1166), .Z(n1164) );
  NANDN U1020 ( .A(A[733]), .B(B[733]), .Z(n1166) );
  AND U1021 ( .A(n1167), .B(n1168), .Z(n1165) );
  NANDN U1022 ( .A(A[732]), .B(B[732]), .Z(n1168) );
  NAND U1023 ( .A(n1169), .B(n1170), .Z(n1167) );
  NANDN U1024 ( .A(B[732]), .B(A[732]), .Z(n1170) );
  AND U1025 ( .A(n1171), .B(n1172), .Z(n1169) );
  NAND U1026 ( .A(n1173), .B(n1174), .Z(n1172) );
  NANDN U1027 ( .A(A[731]), .B(B[731]), .Z(n1174) );
  AND U1028 ( .A(n1175), .B(n1176), .Z(n1173) );
  NANDN U1029 ( .A(A[730]), .B(B[730]), .Z(n1176) );
  NAND U1030 ( .A(n1177), .B(n1178), .Z(n1175) );
  NANDN U1031 ( .A(B[730]), .B(A[730]), .Z(n1178) );
  AND U1032 ( .A(n1179), .B(n1180), .Z(n1177) );
  NAND U1033 ( .A(n1181), .B(n1182), .Z(n1180) );
  NANDN U1034 ( .A(A[729]), .B(B[729]), .Z(n1182) );
  AND U1035 ( .A(n1183), .B(n1184), .Z(n1181) );
  NANDN U1036 ( .A(A[728]), .B(B[728]), .Z(n1184) );
  NAND U1037 ( .A(n1185), .B(n1186), .Z(n1183) );
  NANDN U1038 ( .A(B[728]), .B(A[728]), .Z(n1186) );
  AND U1039 ( .A(n1187), .B(n1188), .Z(n1185) );
  NAND U1040 ( .A(n1189), .B(n1190), .Z(n1188) );
  NANDN U1041 ( .A(A[727]), .B(B[727]), .Z(n1190) );
  AND U1042 ( .A(n1191), .B(n1192), .Z(n1189) );
  NANDN U1043 ( .A(A[726]), .B(B[726]), .Z(n1192) );
  NAND U1044 ( .A(n1193), .B(n1194), .Z(n1191) );
  NANDN U1045 ( .A(B[726]), .B(A[726]), .Z(n1194) );
  AND U1046 ( .A(n1195), .B(n1196), .Z(n1193) );
  NAND U1047 ( .A(n1197), .B(n1198), .Z(n1196) );
  NANDN U1048 ( .A(A[725]), .B(B[725]), .Z(n1198) );
  AND U1049 ( .A(n1199), .B(n1200), .Z(n1197) );
  NANDN U1050 ( .A(A[724]), .B(B[724]), .Z(n1200) );
  NAND U1051 ( .A(n1201), .B(n1202), .Z(n1199) );
  NANDN U1052 ( .A(B[724]), .B(A[724]), .Z(n1202) );
  AND U1053 ( .A(n1203), .B(n1204), .Z(n1201) );
  NAND U1054 ( .A(n1205), .B(n1206), .Z(n1204) );
  NANDN U1055 ( .A(A[723]), .B(B[723]), .Z(n1206) );
  AND U1056 ( .A(n1207), .B(n1208), .Z(n1205) );
  NANDN U1057 ( .A(A[722]), .B(B[722]), .Z(n1208) );
  NAND U1058 ( .A(n1209), .B(n1210), .Z(n1207) );
  NANDN U1059 ( .A(B[722]), .B(A[722]), .Z(n1210) );
  AND U1060 ( .A(n1211), .B(n1212), .Z(n1209) );
  NAND U1061 ( .A(n1213), .B(n1214), .Z(n1212) );
  NANDN U1062 ( .A(A[721]), .B(B[721]), .Z(n1214) );
  AND U1063 ( .A(n1215), .B(n1216), .Z(n1213) );
  NANDN U1064 ( .A(A[720]), .B(B[720]), .Z(n1216) );
  NAND U1065 ( .A(n1217), .B(n1218), .Z(n1215) );
  NANDN U1066 ( .A(B[720]), .B(A[720]), .Z(n1218) );
  AND U1067 ( .A(n1219), .B(n1220), .Z(n1217) );
  NAND U1068 ( .A(n1221), .B(n1222), .Z(n1220) );
  NANDN U1069 ( .A(A[719]), .B(B[719]), .Z(n1222) );
  AND U1070 ( .A(n1223), .B(n1224), .Z(n1221) );
  NANDN U1071 ( .A(A[718]), .B(B[718]), .Z(n1224) );
  NAND U1072 ( .A(n1225), .B(n1226), .Z(n1223) );
  NANDN U1073 ( .A(B[718]), .B(A[718]), .Z(n1226) );
  AND U1074 ( .A(n1227), .B(n1228), .Z(n1225) );
  NAND U1075 ( .A(n1229), .B(n1230), .Z(n1228) );
  NANDN U1076 ( .A(A[717]), .B(B[717]), .Z(n1230) );
  AND U1077 ( .A(n1231), .B(n1232), .Z(n1229) );
  NANDN U1078 ( .A(A[716]), .B(B[716]), .Z(n1232) );
  NAND U1079 ( .A(n1233), .B(n1234), .Z(n1231) );
  NANDN U1080 ( .A(B[716]), .B(A[716]), .Z(n1234) );
  AND U1081 ( .A(n1235), .B(n1236), .Z(n1233) );
  NAND U1082 ( .A(n1237), .B(n1238), .Z(n1236) );
  NANDN U1083 ( .A(A[715]), .B(B[715]), .Z(n1238) );
  AND U1084 ( .A(n1239), .B(n1240), .Z(n1237) );
  NANDN U1085 ( .A(A[714]), .B(B[714]), .Z(n1240) );
  NAND U1086 ( .A(n1241), .B(n1242), .Z(n1239) );
  NANDN U1087 ( .A(B[714]), .B(A[714]), .Z(n1242) );
  AND U1088 ( .A(n1243), .B(n1244), .Z(n1241) );
  NAND U1089 ( .A(n1245), .B(n1246), .Z(n1244) );
  NANDN U1090 ( .A(A[713]), .B(B[713]), .Z(n1246) );
  AND U1091 ( .A(n1247), .B(n1248), .Z(n1245) );
  NANDN U1092 ( .A(A[712]), .B(B[712]), .Z(n1248) );
  NAND U1093 ( .A(n1249), .B(n1250), .Z(n1247) );
  NANDN U1094 ( .A(B[712]), .B(A[712]), .Z(n1250) );
  AND U1095 ( .A(n1251), .B(n1252), .Z(n1249) );
  NAND U1096 ( .A(n1253), .B(n1254), .Z(n1252) );
  NANDN U1097 ( .A(A[711]), .B(B[711]), .Z(n1254) );
  AND U1098 ( .A(n1255), .B(n1256), .Z(n1253) );
  NANDN U1099 ( .A(A[710]), .B(B[710]), .Z(n1256) );
  NAND U1100 ( .A(n1257), .B(n1258), .Z(n1255) );
  NANDN U1101 ( .A(B[710]), .B(A[710]), .Z(n1258) );
  AND U1102 ( .A(n1259), .B(n1260), .Z(n1257) );
  NAND U1103 ( .A(n1261), .B(n1262), .Z(n1260) );
  NANDN U1104 ( .A(A[709]), .B(B[709]), .Z(n1262) );
  AND U1105 ( .A(n1263), .B(n1264), .Z(n1261) );
  NANDN U1106 ( .A(A[708]), .B(B[708]), .Z(n1264) );
  NAND U1107 ( .A(n1265), .B(n1266), .Z(n1263) );
  NANDN U1108 ( .A(B[708]), .B(A[708]), .Z(n1266) );
  AND U1109 ( .A(n1267), .B(n1268), .Z(n1265) );
  NAND U1110 ( .A(n1269), .B(n1270), .Z(n1268) );
  NANDN U1111 ( .A(A[707]), .B(B[707]), .Z(n1270) );
  AND U1112 ( .A(n1271), .B(n1272), .Z(n1269) );
  NANDN U1113 ( .A(A[706]), .B(B[706]), .Z(n1272) );
  NAND U1114 ( .A(n1273), .B(n1274), .Z(n1271) );
  NANDN U1115 ( .A(B[706]), .B(A[706]), .Z(n1274) );
  AND U1116 ( .A(n1275), .B(n1276), .Z(n1273) );
  NAND U1117 ( .A(n1277), .B(n1278), .Z(n1276) );
  NANDN U1118 ( .A(A[705]), .B(B[705]), .Z(n1278) );
  AND U1119 ( .A(n1279), .B(n1280), .Z(n1277) );
  NANDN U1120 ( .A(A[704]), .B(B[704]), .Z(n1280) );
  NAND U1121 ( .A(n1281), .B(n1282), .Z(n1279) );
  NANDN U1122 ( .A(B[704]), .B(A[704]), .Z(n1282) );
  AND U1123 ( .A(n1283), .B(n1284), .Z(n1281) );
  NAND U1124 ( .A(n1285), .B(n1286), .Z(n1284) );
  NANDN U1125 ( .A(A[703]), .B(B[703]), .Z(n1286) );
  AND U1126 ( .A(n1287), .B(n1288), .Z(n1285) );
  NANDN U1127 ( .A(A[702]), .B(B[702]), .Z(n1288) );
  NAND U1128 ( .A(n1289), .B(n1290), .Z(n1287) );
  NANDN U1129 ( .A(B[702]), .B(A[702]), .Z(n1290) );
  AND U1130 ( .A(n1291), .B(n1292), .Z(n1289) );
  NAND U1131 ( .A(n1293), .B(n1294), .Z(n1292) );
  NANDN U1132 ( .A(A[701]), .B(B[701]), .Z(n1294) );
  AND U1133 ( .A(n1295), .B(n1296), .Z(n1293) );
  NANDN U1134 ( .A(A[700]), .B(B[700]), .Z(n1296) );
  NAND U1135 ( .A(n1297), .B(n1298), .Z(n1295) );
  NANDN U1136 ( .A(B[700]), .B(A[700]), .Z(n1298) );
  AND U1137 ( .A(n1299), .B(n1300), .Z(n1297) );
  NAND U1138 ( .A(n1301), .B(n1302), .Z(n1300) );
  NANDN U1139 ( .A(A[699]), .B(B[699]), .Z(n1302) );
  AND U1140 ( .A(n1303), .B(n1304), .Z(n1301) );
  NANDN U1141 ( .A(A[698]), .B(B[698]), .Z(n1304) );
  NAND U1142 ( .A(n1305), .B(n1306), .Z(n1303) );
  NANDN U1143 ( .A(B[698]), .B(A[698]), .Z(n1306) );
  AND U1144 ( .A(n1307), .B(n1308), .Z(n1305) );
  NAND U1145 ( .A(n1309), .B(n1310), .Z(n1308) );
  NANDN U1146 ( .A(A[697]), .B(B[697]), .Z(n1310) );
  AND U1147 ( .A(n1311), .B(n1312), .Z(n1309) );
  NANDN U1148 ( .A(A[696]), .B(B[696]), .Z(n1312) );
  NAND U1149 ( .A(n1313), .B(n1314), .Z(n1311) );
  NANDN U1150 ( .A(B[696]), .B(A[696]), .Z(n1314) );
  AND U1151 ( .A(n1315), .B(n1316), .Z(n1313) );
  NAND U1152 ( .A(n1317), .B(n1318), .Z(n1316) );
  NANDN U1153 ( .A(A[695]), .B(B[695]), .Z(n1318) );
  AND U1154 ( .A(n1319), .B(n1320), .Z(n1317) );
  NANDN U1155 ( .A(A[694]), .B(B[694]), .Z(n1320) );
  NAND U1156 ( .A(n1321), .B(n1322), .Z(n1319) );
  NANDN U1157 ( .A(B[694]), .B(A[694]), .Z(n1322) );
  AND U1158 ( .A(n1323), .B(n1324), .Z(n1321) );
  NAND U1159 ( .A(n1325), .B(n1326), .Z(n1324) );
  NANDN U1160 ( .A(A[693]), .B(B[693]), .Z(n1326) );
  AND U1161 ( .A(n1327), .B(n1328), .Z(n1325) );
  NANDN U1162 ( .A(A[692]), .B(B[692]), .Z(n1328) );
  NAND U1163 ( .A(n1329), .B(n1330), .Z(n1327) );
  NANDN U1164 ( .A(B[692]), .B(A[692]), .Z(n1330) );
  AND U1165 ( .A(n1331), .B(n1332), .Z(n1329) );
  NAND U1166 ( .A(n1333), .B(n1334), .Z(n1332) );
  NANDN U1167 ( .A(A[691]), .B(B[691]), .Z(n1334) );
  AND U1168 ( .A(n1335), .B(n1336), .Z(n1333) );
  NANDN U1169 ( .A(A[690]), .B(B[690]), .Z(n1336) );
  NAND U1170 ( .A(n1337), .B(n1338), .Z(n1335) );
  NANDN U1171 ( .A(B[690]), .B(A[690]), .Z(n1338) );
  AND U1172 ( .A(n1339), .B(n1340), .Z(n1337) );
  NAND U1173 ( .A(n1341), .B(n1342), .Z(n1340) );
  NANDN U1174 ( .A(A[689]), .B(B[689]), .Z(n1342) );
  AND U1175 ( .A(n1343), .B(n1344), .Z(n1341) );
  NANDN U1176 ( .A(A[688]), .B(B[688]), .Z(n1344) );
  NAND U1177 ( .A(n1345), .B(n1346), .Z(n1343) );
  NANDN U1178 ( .A(B[688]), .B(A[688]), .Z(n1346) );
  AND U1179 ( .A(n1347), .B(n1348), .Z(n1345) );
  NAND U1180 ( .A(n1349), .B(n1350), .Z(n1348) );
  NANDN U1181 ( .A(A[687]), .B(B[687]), .Z(n1350) );
  AND U1182 ( .A(n1351), .B(n1352), .Z(n1349) );
  NANDN U1183 ( .A(A[686]), .B(B[686]), .Z(n1352) );
  NAND U1184 ( .A(n1353), .B(n1354), .Z(n1351) );
  NANDN U1185 ( .A(B[686]), .B(A[686]), .Z(n1354) );
  AND U1186 ( .A(n1355), .B(n1356), .Z(n1353) );
  NAND U1187 ( .A(n1357), .B(n1358), .Z(n1356) );
  NANDN U1188 ( .A(A[685]), .B(B[685]), .Z(n1358) );
  AND U1189 ( .A(n1359), .B(n1360), .Z(n1357) );
  NANDN U1190 ( .A(A[684]), .B(B[684]), .Z(n1360) );
  NAND U1191 ( .A(n1361), .B(n1362), .Z(n1359) );
  NANDN U1192 ( .A(B[684]), .B(A[684]), .Z(n1362) );
  AND U1193 ( .A(n1363), .B(n1364), .Z(n1361) );
  NAND U1194 ( .A(n1365), .B(n1366), .Z(n1364) );
  NANDN U1195 ( .A(A[683]), .B(B[683]), .Z(n1366) );
  AND U1196 ( .A(n1367), .B(n1368), .Z(n1365) );
  NANDN U1197 ( .A(A[682]), .B(B[682]), .Z(n1368) );
  NAND U1198 ( .A(n1369), .B(n1370), .Z(n1367) );
  NANDN U1199 ( .A(B[682]), .B(A[682]), .Z(n1370) );
  AND U1200 ( .A(n1371), .B(n1372), .Z(n1369) );
  NAND U1201 ( .A(n1373), .B(n1374), .Z(n1372) );
  NANDN U1202 ( .A(A[681]), .B(B[681]), .Z(n1374) );
  AND U1203 ( .A(n1375), .B(n1376), .Z(n1373) );
  NANDN U1204 ( .A(A[680]), .B(B[680]), .Z(n1376) );
  NAND U1205 ( .A(n1377), .B(n1378), .Z(n1375) );
  NANDN U1206 ( .A(B[680]), .B(A[680]), .Z(n1378) );
  AND U1207 ( .A(n1379), .B(n1380), .Z(n1377) );
  NAND U1208 ( .A(n1381), .B(n1382), .Z(n1380) );
  NANDN U1209 ( .A(A[679]), .B(B[679]), .Z(n1382) );
  AND U1210 ( .A(n1383), .B(n1384), .Z(n1381) );
  NANDN U1211 ( .A(A[678]), .B(B[678]), .Z(n1384) );
  NAND U1212 ( .A(n1385), .B(n1386), .Z(n1383) );
  NANDN U1213 ( .A(B[678]), .B(A[678]), .Z(n1386) );
  AND U1214 ( .A(n1387), .B(n1388), .Z(n1385) );
  NAND U1215 ( .A(n1389), .B(n1390), .Z(n1388) );
  NANDN U1216 ( .A(A[677]), .B(B[677]), .Z(n1390) );
  AND U1217 ( .A(n1391), .B(n1392), .Z(n1389) );
  NANDN U1218 ( .A(A[676]), .B(B[676]), .Z(n1392) );
  NAND U1219 ( .A(n1393), .B(n1394), .Z(n1391) );
  NANDN U1220 ( .A(B[676]), .B(A[676]), .Z(n1394) );
  AND U1221 ( .A(n1395), .B(n1396), .Z(n1393) );
  NAND U1222 ( .A(n1397), .B(n1398), .Z(n1396) );
  NANDN U1223 ( .A(A[675]), .B(B[675]), .Z(n1398) );
  AND U1224 ( .A(n1399), .B(n1400), .Z(n1397) );
  NANDN U1225 ( .A(A[674]), .B(B[674]), .Z(n1400) );
  NAND U1226 ( .A(n1401), .B(n1402), .Z(n1399) );
  NANDN U1227 ( .A(B[674]), .B(A[674]), .Z(n1402) );
  AND U1228 ( .A(n1403), .B(n1404), .Z(n1401) );
  NAND U1229 ( .A(n1405), .B(n1406), .Z(n1404) );
  NANDN U1230 ( .A(A[673]), .B(B[673]), .Z(n1406) );
  AND U1231 ( .A(n1407), .B(n1408), .Z(n1405) );
  NANDN U1232 ( .A(A[672]), .B(B[672]), .Z(n1408) );
  NAND U1233 ( .A(n1409), .B(n1410), .Z(n1407) );
  NANDN U1234 ( .A(B[672]), .B(A[672]), .Z(n1410) );
  AND U1235 ( .A(n1411), .B(n1412), .Z(n1409) );
  NAND U1236 ( .A(n1413), .B(n1414), .Z(n1412) );
  NANDN U1237 ( .A(A[671]), .B(B[671]), .Z(n1414) );
  AND U1238 ( .A(n1415), .B(n1416), .Z(n1413) );
  NANDN U1239 ( .A(A[670]), .B(B[670]), .Z(n1416) );
  NAND U1240 ( .A(n1417), .B(n1418), .Z(n1415) );
  NANDN U1241 ( .A(B[670]), .B(A[670]), .Z(n1418) );
  AND U1242 ( .A(n1419), .B(n1420), .Z(n1417) );
  NAND U1243 ( .A(n1421), .B(n1422), .Z(n1420) );
  NANDN U1244 ( .A(A[669]), .B(B[669]), .Z(n1422) );
  AND U1245 ( .A(n1423), .B(n1424), .Z(n1421) );
  NANDN U1246 ( .A(A[668]), .B(B[668]), .Z(n1424) );
  NAND U1247 ( .A(n1425), .B(n1426), .Z(n1423) );
  NANDN U1248 ( .A(B[668]), .B(A[668]), .Z(n1426) );
  AND U1249 ( .A(n1427), .B(n1428), .Z(n1425) );
  NAND U1250 ( .A(n1429), .B(n1430), .Z(n1428) );
  NANDN U1251 ( .A(A[667]), .B(B[667]), .Z(n1430) );
  AND U1252 ( .A(n1431), .B(n1432), .Z(n1429) );
  NANDN U1253 ( .A(A[666]), .B(B[666]), .Z(n1432) );
  NAND U1254 ( .A(n1433), .B(n1434), .Z(n1431) );
  NANDN U1255 ( .A(B[666]), .B(A[666]), .Z(n1434) );
  AND U1256 ( .A(n1435), .B(n1436), .Z(n1433) );
  NAND U1257 ( .A(n1437), .B(n1438), .Z(n1436) );
  NANDN U1258 ( .A(A[665]), .B(B[665]), .Z(n1438) );
  AND U1259 ( .A(n1439), .B(n1440), .Z(n1437) );
  NANDN U1260 ( .A(A[664]), .B(B[664]), .Z(n1440) );
  NAND U1261 ( .A(n1441), .B(n1442), .Z(n1439) );
  NANDN U1262 ( .A(B[664]), .B(A[664]), .Z(n1442) );
  AND U1263 ( .A(n1443), .B(n1444), .Z(n1441) );
  NAND U1264 ( .A(n1445), .B(n1446), .Z(n1444) );
  NANDN U1265 ( .A(A[663]), .B(B[663]), .Z(n1446) );
  AND U1266 ( .A(n1447), .B(n1448), .Z(n1445) );
  NANDN U1267 ( .A(A[662]), .B(B[662]), .Z(n1448) );
  NAND U1268 ( .A(n1449), .B(n1450), .Z(n1447) );
  NANDN U1269 ( .A(B[662]), .B(A[662]), .Z(n1450) );
  AND U1270 ( .A(n1451), .B(n1452), .Z(n1449) );
  NAND U1271 ( .A(n1453), .B(n1454), .Z(n1452) );
  NANDN U1272 ( .A(A[661]), .B(B[661]), .Z(n1454) );
  AND U1273 ( .A(n1455), .B(n1456), .Z(n1453) );
  NANDN U1274 ( .A(A[660]), .B(B[660]), .Z(n1456) );
  NAND U1275 ( .A(n1457), .B(n1458), .Z(n1455) );
  NANDN U1276 ( .A(B[660]), .B(A[660]), .Z(n1458) );
  AND U1277 ( .A(n1459), .B(n1460), .Z(n1457) );
  NAND U1278 ( .A(n1461), .B(n1462), .Z(n1460) );
  NANDN U1279 ( .A(A[659]), .B(B[659]), .Z(n1462) );
  AND U1280 ( .A(n1463), .B(n1464), .Z(n1461) );
  NANDN U1281 ( .A(A[658]), .B(B[658]), .Z(n1464) );
  NAND U1282 ( .A(n1465), .B(n1466), .Z(n1463) );
  NANDN U1283 ( .A(B[658]), .B(A[658]), .Z(n1466) );
  AND U1284 ( .A(n1467), .B(n1468), .Z(n1465) );
  NAND U1285 ( .A(n1469), .B(n1470), .Z(n1468) );
  NANDN U1286 ( .A(A[657]), .B(B[657]), .Z(n1470) );
  AND U1287 ( .A(n1471), .B(n1472), .Z(n1469) );
  NANDN U1288 ( .A(A[656]), .B(B[656]), .Z(n1472) );
  NAND U1289 ( .A(n1473), .B(n1474), .Z(n1471) );
  NANDN U1290 ( .A(B[656]), .B(A[656]), .Z(n1474) );
  AND U1291 ( .A(n1475), .B(n1476), .Z(n1473) );
  NAND U1292 ( .A(n1477), .B(n1478), .Z(n1476) );
  NANDN U1293 ( .A(A[655]), .B(B[655]), .Z(n1478) );
  AND U1294 ( .A(n1479), .B(n1480), .Z(n1477) );
  NANDN U1295 ( .A(A[654]), .B(B[654]), .Z(n1480) );
  NAND U1296 ( .A(n1481), .B(n1482), .Z(n1479) );
  NANDN U1297 ( .A(B[654]), .B(A[654]), .Z(n1482) );
  AND U1298 ( .A(n1483), .B(n1484), .Z(n1481) );
  NAND U1299 ( .A(n1485), .B(n1486), .Z(n1484) );
  NANDN U1300 ( .A(A[653]), .B(B[653]), .Z(n1486) );
  AND U1301 ( .A(n1487), .B(n1488), .Z(n1485) );
  NANDN U1302 ( .A(A[652]), .B(B[652]), .Z(n1488) );
  NAND U1303 ( .A(n1489), .B(n1490), .Z(n1487) );
  NANDN U1304 ( .A(B[652]), .B(A[652]), .Z(n1490) );
  AND U1305 ( .A(n1491), .B(n1492), .Z(n1489) );
  NAND U1306 ( .A(n1493), .B(n1494), .Z(n1492) );
  NANDN U1307 ( .A(A[651]), .B(B[651]), .Z(n1494) );
  AND U1308 ( .A(n1495), .B(n1496), .Z(n1493) );
  NANDN U1309 ( .A(A[650]), .B(B[650]), .Z(n1496) );
  NAND U1310 ( .A(n1497), .B(n1498), .Z(n1495) );
  NANDN U1311 ( .A(B[650]), .B(A[650]), .Z(n1498) );
  AND U1312 ( .A(n1499), .B(n1500), .Z(n1497) );
  NAND U1313 ( .A(n1501), .B(n1502), .Z(n1500) );
  NANDN U1314 ( .A(A[649]), .B(B[649]), .Z(n1502) );
  AND U1315 ( .A(n1503), .B(n1504), .Z(n1501) );
  NANDN U1316 ( .A(A[648]), .B(B[648]), .Z(n1504) );
  NAND U1317 ( .A(n1505), .B(n1506), .Z(n1503) );
  NANDN U1318 ( .A(B[648]), .B(A[648]), .Z(n1506) );
  AND U1319 ( .A(n1507), .B(n1508), .Z(n1505) );
  NAND U1320 ( .A(n1509), .B(n1510), .Z(n1508) );
  NANDN U1321 ( .A(A[647]), .B(B[647]), .Z(n1510) );
  AND U1322 ( .A(n1511), .B(n1512), .Z(n1509) );
  NANDN U1323 ( .A(A[646]), .B(B[646]), .Z(n1512) );
  NAND U1324 ( .A(n1513), .B(n1514), .Z(n1511) );
  NANDN U1325 ( .A(B[646]), .B(A[646]), .Z(n1514) );
  AND U1326 ( .A(n1515), .B(n1516), .Z(n1513) );
  NAND U1327 ( .A(n1517), .B(n1518), .Z(n1516) );
  NANDN U1328 ( .A(A[645]), .B(B[645]), .Z(n1518) );
  AND U1329 ( .A(n1519), .B(n1520), .Z(n1517) );
  NANDN U1330 ( .A(A[644]), .B(B[644]), .Z(n1520) );
  NAND U1331 ( .A(n1521), .B(n1522), .Z(n1519) );
  NANDN U1332 ( .A(B[644]), .B(A[644]), .Z(n1522) );
  AND U1333 ( .A(n1523), .B(n1524), .Z(n1521) );
  NAND U1334 ( .A(n1525), .B(n1526), .Z(n1524) );
  NANDN U1335 ( .A(A[643]), .B(B[643]), .Z(n1526) );
  AND U1336 ( .A(n1527), .B(n1528), .Z(n1525) );
  NANDN U1337 ( .A(A[642]), .B(B[642]), .Z(n1528) );
  NAND U1338 ( .A(n1529), .B(n1530), .Z(n1527) );
  NANDN U1339 ( .A(B[642]), .B(A[642]), .Z(n1530) );
  AND U1340 ( .A(n1531), .B(n1532), .Z(n1529) );
  NAND U1341 ( .A(n1533), .B(n1534), .Z(n1532) );
  NANDN U1342 ( .A(A[641]), .B(B[641]), .Z(n1534) );
  AND U1343 ( .A(n1535), .B(n1536), .Z(n1533) );
  NANDN U1344 ( .A(A[640]), .B(B[640]), .Z(n1536) );
  NAND U1345 ( .A(n1537), .B(n1538), .Z(n1535) );
  NANDN U1346 ( .A(B[640]), .B(A[640]), .Z(n1538) );
  AND U1347 ( .A(n1539), .B(n1540), .Z(n1537) );
  NAND U1348 ( .A(n1541), .B(n1542), .Z(n1540) );
  NANDN U1349 ( .A(A[639]), .B(B[639]), .Z(n1542) );
  AND U1350 ( .A(n1543), .B(n1544), .Z(n1541) );
  NANDN U1351 ( .A(A[638]), .B(B[638]), .Z(n1544) );
  NAND U1352 ( .A(n1545), .B(n1546), .Z(n1543) );
  NANDN U1353 ( .A(B[638]), .B(A[638]), .Z(n1546) );
  AND U1354 ( .A(n1547), .B(n1548), .Z(n1545) );
  NAND U1355 ( .A(n1549), .B(n1550), .Z(n1548) );
  NANDN U1356 ( .A(A[637]), .B(B[637]), .Z(n1550) );
  AND U1357 ( .A(n1551), .B(n1552), .Z(n1549) );
  NANDN U1358 ( .A(A[636]), .B(B[636]), .Z(n1552) );
  NAND U1359 ( .A(n1553), .B(n1554), .Z(n1551) );
  NANDN U1360 ( .A(B[636]), .B(A[636]), .Z(n1554) );
  AND U1361 ( .A(n1555), .B(n1556), .Z(n1553) );
  NAND U1362 ( .A(n1557), .B(n1558), .Z(n1556) );
  NANDN U1363 ( .A(A[635]), .B(B[635]), .Z(n1558) );
  AND U1364 ( .A(n1559), .B(n1560), .Z(n1557) );
  NANDN U1365 ( .A(A[634]), .B(B[634]), .Z(n1560) );
  NAND U1366 ( .A(n1561), .B(n1562), .Z(n1559) );
  NANDN U1367 ( .A(B[634]), .B(A[634]), .Z(n1562) );
  AND U1368 ( .A(n1563), .B(n1564), .Z(n1561) );
  NAND U1369 ( .A(n1565), .B(n1566), .Z(n1564) );
  NANDN U1370 ( .A(A[633]), .B(B[633]), .Z(n1566) );
  AND U1371 ( .A(n1567), .B(n1568), .Z(n1565) );
  NANDN U1372 ( .A(A[632]), .B(B[632]), .Z(n1568) );
  NAND U1373 ( .A(n1569), .B(n1570), .Z(n1567) );
  NANDN U1374 ( .A(B[632]), .B(A[632]), .Z(n1570) );
  AND U1375 ( .A(n1571), .B(n1572), .Z(n1569) );
  NAND U1376 ( .A(n1573), .B(n1574), .Z(n1572) );
  NANDN U1377 ( .A(A[631]), .B(B[631]), .Z(n1574) );
  AND U1378 ( .A(n1575), .B(n1576), .Z(n1573) );
  NANDN U1379 ( .A(A[630]), .B(B[630]), .Z(n1576) );
  NAND U1380 ( .A(n1577), .B(n1578), .Z(n1575) );
  NANDN U1381 ( .A(B[630]), .B(A[630]), .Z(n1578) );
  AND U1382 ( .A(n1579), .B(n1580), .Z(n1577) );
  NAND U1383 ( .A(n1581), .B(n1582), .Z(n1580) );
  NANDN U1384 ( .A(A[629]), .B(B[629]), .Z(n1582) );
  AND U1385 ( .A(n1583), .B(n1584), .Z(n1581) );
  NANDN U1386 ( .A(A[628]), .B(B[628]), .Z(n1584) );
  NAND U1387 ( .A(n1585), .B(n1586), .Z(n1583) );
  NANDN U1388 ( .A(B[628]), .B(A[628]), .Z(n1586) );
  AND U1389 ( .A(n1587), .B(n1588), .Z(n1585) );
  NAND U1390 ( .A(n1589), .B(n1590), .Z(n1588) );
  NANDN U1391 ( .A(A[627]), .B(B[627]), .Z(n1590) );
  AND U1392 ( .A(n1591), .B(n1592), .Z(n1589) );
  NANDN U1393 ( .A(A[626]), .B(B[626]), .Z(n1592) );
  NAND U1394 ( .A(n1593), .B(n1594), .Z(n1591) );
  NANDN U1395 ( .A(B[626]), .B(A[626]), .Z(n1594) );
  AND U1396 ( .A(n1595), .B(n1596), .Z(n1593) );
  NAND U1397 ( .A(n1597), .B(n1598), .Z(n1596) );
  NANDN U1398 ( .A(A[625]), .B(B[625]), .Z(n1598) );
  AND U1399 ( .A(n1599), .B(n1600), .Z(n1597) );
  NANDN U1400 ( .A(A[624]), .B(B[624]), .Z(n1600) );
  NAND U1401 ( .A(n1601), .B(n1602), .Z(n1599) );
  NANDN U1402 ( .A(B[624]), .B(A[624]), .Z(n1602) );
  AND U1403 ( .A(n1603), .B(n1604), .Z(n1601) );
  NAND U1404 ( .A(n1605), .B(n1606), .Z(n1604) );
  NANDN U1405 ( .A(A[623]), .B(B[623]), .Z(n1606) );
  AND U1406 ( .A(n1607), .B(n1608), .Z(n1605) );
  NANDN U1407 ( .A(A[622]), .B(B[622]), .Z(n1608) );
  NAND U1408 ( .A(n1609), .B(n1610), .Z(n1607) );
  NANDN U1409 ( .A(B[622]), .B(A[622]), .Z(n1610) );
  AND U1410 ( .A(n1611), .B(n1612), .Z(n1609) );
  NAND U1411 ( .A(n1613), .B(n1614), .Z(n1612) );
  NANDN U1412 ( .A(A[621]), .B(B[621]), .Z(n1614) );
  AND U1413 ( .A(n1615), .B(n1616), .Z(n1613) );
  NANDN U1414 ( .A(A[620]), .B(B[620]), .Z(n1616) );
  NAND U1415 ( .A(n1617), .B(n1618), .Z(n1615) );
  NANDN U1416 ( .A(B[620]), .B(A[620]), .Z(n1618) );
  AND U1417 ( .A(n1619), .B(n1620), .Z(n1617) );
  NAND U1418 ( .A(n1621), .B(n1622), .Z(n1620) );
  NANDN U1419 ( .A(A[619]), .B(B[619]), .Z(n1622) );
  AND U1420 ( .A(n1623), .B(n1624), .Z(n1621) );
  NANDN U1421 ( .A(A[618]), .B(B[618]), .Z(n1624) );
  NAND U1422 ( .A(n1625), .B(n1626), .Z(n1623) );
  NANDN U1423 ( .A(B[618]), .B(A[618]), .Z(n1626) );
  AND U1424 ( .A(n1627), .B(n1628), .Z(n1625) );
  NAND U1425 ( .A(n1629), .B(n1630), .Z(n1628) );
  NANDN U1426 ( .A(A[617]), .B(B[617]), .Z(n1630) );
  AND U1427 ( .A(n1631), .B(n1632), .Z(n1629) );
  NANDN U1428 ( .A(A[616]), .B(B[616]), .Z(n1632) );
  NAND U1429 ( .A(n1633), .B(n1634), .Z(n1631) );
  NANDN U1430 ( .A(B[616]), .B(A[616]), .Z(n1634) );
  AND U1431 ( .A(n1635), .B(n1636), .Z(n1633) );
  NAND U1432 ( .A(n1637), .B(n1638), .Z(n1636) );
  NANDN U1433 ( .A(A[615]), .B(B[615]), .Z(n1638) );
  AND U1434 ( .A(n1639), .B(n1640), .Z(n1637) );
  NANDN U1435 ( .A(A[614]), .B(B[614]), .Z(n1640) );
  NAND U1436 ( .A(n1641), .B(n1642), .Z(n1639) );
  NANDN U1437 ( .A(B[614]), .B(A[614]), .Z(n1642) );
  AND U1438 ( .A(n1643), .B(n1644), .Z(n1641) );
  NAND U1439 ( .A(n1645), .B(n1646), .Z(n1644) );
  NANDN U1440 ( .A(A[613]), .B(B[613]), .Z(n1646) );
  AND U1441 ( .A(n1647), .B(n1648), .Z(n1645) );
  NANDN U1442 ( .A(A[612]), .B(B[612]), .Z(n1648) );
  NAND U1443 ( .A(n1649), .B(n1650), .Z(n1647) );
  NANDN U1444 ( .A(B[612]), .B(A[612]), .Z(n1650) );
  AND U1445 ( .A(n1651), .B(n1652), .Z(n1649) );
  NAND U1446 ( .A(n1653), .B(n1654), .Z(n1652) );
  NANDN U1447 ( .A(A[611]), .B(B[611]), .Z(n1654) );
  AND U1448 ( .A(n1655), .B(n1656), .Z(n1653) );
  NANDN U1449 ( .A(A[610]), .B(B[610]), .Z(n1656) );
  NAND U1450 ( .A(n1657), .B(n1658), .Z(n1655) );
  NANDN U1451 ( .A(B[610]), .B(A[610]), .Z(n1658) );
  AND U1452 ( .A(n1659), .B(n1660), .Z(n1657) );
  NAND U1453 ( .A(n1661), .B(n1662), .Z(n1660) );
  NANDN U1454 ( .A(A[609]), .B(B[609]), .Z(n1662) );
  AND U1455 ( .A(n1663), .B(n1664), .Z(n1661) );
  NANDN U1456 ( .A(A[608]), .B(B[608]), .Z(n1664) );
  NAND U1457 ( .A(n1665), .B(n1666), .Z(n1663) );
  NANDN U1458 ( .A(B[608]), .B(A[608]), .Z(n1666) );
  AND U1459 ( .A(n1667), .B(n1668), .Z(n1665) );
  NAND U1460 ( .A(n1669), .B(n1670), .Z(n1668) );
  NANDN U1461 ( .A(A[607]), .B(B[607]), .Z(n1670) );
  AND U1462 ( .A(n1671), .B(n1672), .Z(n1669) );
  NANDN U1463 ( .A(A[606]), .B(B[606]), .Z(n1672) );
  NAND U1464 ( .A(n1673), .B(n1674), .Z(n1671) );
  NANDN U1465 ( .A(B[606]), .B(A[606]), .Z(n1674) );
  AND U1466 ( .A(n1675), .B(n1676), .Z(n1673) );
  NAND U1467 ( .A(n1677), .B(n1678), .Z(n1676) );
  NANDN U1468 ( .A(A[605]), .B(B[605]), .Z(n1678) );
  AND U1469 ( .A(n1679), .B(n1680), .Z(n1677) );
  NANDN U1470 ( .A(A[604]), .B(B[604]), .Z(n1680) );
  NAND U1471 ( .A(n1681), .B(n1682), .Z(n1679) );
  NANDN U1472 ( .A(B[604]), .B(A[604]), .Z(n1682) );
  AND U1473 ( .A(n1683), .B(n1684), .Z(n1681) );
  NAND U1474 ( .A(n1685), .B(n1686), .Z(n1684) );
  NANDN U1475 ( .A(A[603]), .B(B[603]), .Z(n1686) );
  AND U1476 ( .A(n1687), .B(n1688), .Z(n1685) );
  NANDN U1477 ( .A(A[602]), .B(B[602]), .Z(n1688) );
  NAND U1478 ( .A(n1689), .B(n1690), .Z(n1687) );
  NANDN U1479 ( .A(B[602]), .B(A[602]), .Z(n1690) );
  AND U1480 ( .A(n1691), .B(n1692), .Z(n1689) );
  NAND U1481 ( .A(n1693), .B(n1694), .Z(n1692) );
  NANDN U1482 ( .A(A[601]), .B(B[601]), .Z(n1694) );
  AND U1483 ( .A(n1695), .B(n1696), .Z(n1693) );
  NANDN U1484 ( .A(A[600]), .B(B[600]), .Z(n1696) );
  NAND U1485 ( .A(n1697), .B(n1698), .Z(n1695) );
  NANDN U1486 ( .A(B[600]), .B(A[600]), .Z(n1698) );
  AND U1487 ( .A(n1699), .B(n1700), .Z(n1697) );
  NAND U1488 ( .A(n1701), .B(n1702), .Z(n1700) );
  NANDN U1489 ( .A(A[599]), .B(B[599]), .Z(n1702) );
  AND U1490 ( .A(n1703), .B(n1704), .Z(n1701) );
  NANDN U1491 ( .A(A[598]), .B(B[598]), .Z(n1704) );
  NAND U1492 ( .A(n1705), .B(n1706), .Z(n1703) );
  NANDN U1493 ( .A(B[598]), .B(A[598]), .Z(n1706) );
  AND U1494 ( .A(n1707), .B(n1708), .Z(n1705) );
  NAND U1495 ( .A(n1709), .B(n1710), .Z(n1708) );
  NANDN U1496 ( .A(A[597]), .B(B[597]), .Z(n1710) );
  AND U1497 ( .A(n1711), .B(n1712), .Z(n1709) );
  NANDN U1498 ( .A(A[596]), .B(B[596]), .Z(n1712) );
  NAND U1499 ( .A(n1713), .B(n1714), .Z(n1711) );
  NANDN U1500 ( .A(B[596]), .B(A[596]), .Z(n1714) );
  AND U1501 ( .A(n1715), .B(n1716), .Z(n1713) );
  NAND U1502 ( .A(n1717), .B(n1718), .Z(n1716) );
  NANDN U1503 ( .A(A[595]), .B(B[595]), .Z(n1718) );
  AND U1504 ( .A(n1719), .B(n1720), .Z(n1717) );
  NANDN U1505 ( .A(A[594]), .B(B[594]), .Z(n1720) );
  NAND U1506 ( .A(n1721), .B(n1722), .Z(n1719) );
  NANDN U1507 ( .A(B[594]), .B(A[594]), .Z(n1722) );
  AND U1508 ( .A(n1723), .B(n1724), .Z(n1721) );
  NAND U1509 ( .A(n1725), .B(n1726), .Z(n1724) );
  NANDN U1510 ( .A(A[593]), .B(B[593]), .Z(n1726) );
  AND U1511 ( .A(n1727), .B(n1728), .Z(n1725) );
  NANDN U1512 ( .A(A[592]), .B(B[592]), .Z(n1728) );
  NAND U1513 ( .A(n1729), .B(n1730), .Z(n1727) );
  NANDN U1514 ( .A(B[592]), .B(A[592]), .Z(n1730) );
  AND U1515 ( .A(n1731), .B(n1732), .Z(n1729) );
  NAND U1516 ( .A(n1733), .B(n1734), .Z(n1732) );
  NANDN U1517 ( .A(A[591]), .B(B[591]), .Z(n1734) );
  AND U1518 ( .A(n1735), .B(n1736), .Z(n1733) );
  NANDN U1519 ( .A(A[590]), .B(B[590]), .Z(n1736) );
  NAND U1520 ( .A(n1737), .B(n1738), .Z(n1735) );
  NANDN U1521 ( .A(B[590]), .B(A[590]), .Z(n1738) );
  AND U1522 ( .A(n1739), .B(n1740), .Z(n1737) );
  NAND U1523 ( .A(n1741), .B(n1742), .Z(n1740) );
  NANDN U1524 ( .A(A[589]), .B(B[589]), .Z(n1742) );
  AND U1525 ( .A(n1743), .B(n1744), .Z(n1741) );
  NANDN U1526 ( .A(A[588]), .B(B[588]), .Z(n1744) );
  NAND U1527 ( .A(n1745), .B(n1746), .Z(n1743) );
  NANDN U1528 ( .A(B[588]), .B(A[588]), .Z(n1746) );
  AND U1529 ( .A(n1747), .B(n1748), .Z(n1745) );
  NAND U1530 ( .A(n1749), .B(n1750), .Z(n1748) );
  NANDN U1531 ( .A(A[587]), .B(B[587]), .Z(n1750) );
  AND U1532 ( .A(n1751), .B(n1752), .Z(n1749) );
  NANDN U1533 ( .A(A[586]), .B(B[586]), .Z(n1752) );
  NAND U1534 ( .A(n1753), .B(n1754), .Z(n1751) );
  NANDN U1535 ( .A(B[586]), .B(A[586]), .Z(n1754) );
  AND U1536 ( .A(n1755), .B(n1756), .Z(n1753) );
  NAND U1537 ( .A(n1757), .B(n1758), .Z(n1756) );
  NANDN U1538 ( .A(A[585]), .B(B[585]), .Z(n1758) );
  AND U1539 ( .A(n1759), .B(n1760), .Z(n1757) );
  NANDN U1540 ( .A(A[584]), .B(B[584]), .Z(n1760) );
  NAND U1541 ( .A(n1761), .B(n1762), .Z(n1759) );
  NANDN U1542 ( .A(B[584]), .B(A[584]), .Z(n1762) );
  AND U1543 ( .A(n1763), .B(n1764), .Z(n1761) );
  NAND U1544 ( .A(n1765), .B(n1766), .Z(n1764) );
  NANDN U1545 ( .A(A[583]), .B(B[583]), .Z(n1766) );
  AND U1546 ( .A(n1767), .B(n1768), .Z(n1765) );
  NANDN U1547 ( .A(A[582]), .B(B[582]), .Z(n1768) );
  NAND U1548 ( .A(n1769), .B(n1770), .Z(n1767) );
  NANDN U1549 ( .A(B[582]), .B(A[582]), .Z(n1770) );
  AND U1550 ( .A(n1771), .B(n1772), .Z(n1769) );
  NAND U1551 ( .A(n1773), .B(n1774), .Z(n1772) );
  NANDN U1552 ( .A(A[581]), .B(B[581]), .Z(n1774) );
  AND U1553 ( .A(n1775), .B(n1776), .Z(n1773) );
  NANDN U1554 ( .A(A[580]), .B(B[580]), .Z(n1776) );
  NAND U1555 ( .A(n1777), .B(n1778), .Z(n1775) );
  NANDN U1556 ( .A(B[580]), .B(A[580]), .Z(n1778) );
  AND U1557 ( .A(n1779), .B(n1780), .Z(n1777) );
  NAND U1558 ( .A(n1781), .B(n1782), .Z(n1780) );
  NANDN U1559 ( .A(A[579]), .B(B[579]), .Z(n1782) );
  AND U1560 ( .A(n1783), .B(n1784), .Z(n1781) );
  NANDN U1561 ( .A(A[578]), .B(B[578]), .Z(n1784) );
  NAND U1562 ( .A(n1785), .B(n1786), .Z(n1783) );
  NANDN U1563 ( .A(B[578]), .B(A[578]), .Z(n1786) );
  AND U1564 ( .A(n1787), .B(n1788), .Z(n1785) );
  NAND U1565 ( .A(n1789), .B(n1790), .Z(n1788) );
  NANDN U1566 ( .A(A[577]), .B(B[577]), .Z(n1790) );
  AND U1567 ( .A(n1791), .B(n1792), .Z(n1789) );
  NANDN U1568 ( .A(A[576]), .B(B[576]), .Z(n1792) );
  NAND U1569 ( .A(n1793), .B(n1794), .Z(n1791) );
  NANDN U1570 ( .A(B[576]), .B(A[576]), .Z(n1794) );
  AND U1571 ( .A(n1795), .B(n1796), .Z(n1793) );
  NAND U1572 ( .A(n1797), .B(n1798), .Z(n1796) );
  NANDN U1573 ( .A(A[575]), .B(B[575]), .Z(n1798) );
  AND U1574 ( .A(n1799), .B(n1800), .Z(n1797) );
  NANDN U1575 ( .A(A[574]), .B(B[574]), .Z(n1800) );
  NAND U1576 ( .A(n1801), .B(n1802), .Z(n1799) );
  NANDN U1577 ( .A(B[574]), .B(A[574]), .Z(n1802) );
  AND U1578 ( .A(n1803), .B(n1804), .Z(n1801) );
  NAND U1579 ( .A(n1805), .B(n1806), .Z(n1804) );
  NANDN U1580 ( .A(A[573]), .B(B[573]), .Z(n1806) );
  AND U1581 ( .A(n1807), .B(n1808), .Z(n1805) );
  NANDN U1582 ( .A(A[572]), .B(B[572]), .Z(n1808) );
  NAND U1583 ( .A(n1809), .B(n1810), .Z(n1807) );
  NANDN U1584 ( .A(B[572]), .B(A[572]), .Z(n1810) );
  AND U1585 ( .A(n1811), .B(n1812), .Z(n1809) );
  NAND U1586 ( .A(n1813), .B(n1814), .Z(n1812) );
  NANDN U1587 ( .A(A[571]), .B(B[571]), .Z(n1814) );
  AND U1588 ( .A(n1815), .B(n1816), .Z(n1813) );
  NANDN U1589 ( .A(A[570]), .B(B[570]), .Z(n1816) );
  NAND U1590 ( .A(n1817), .B(n1818), .Z(n1815) );
  NANDN U1591 ( .A(B[570]), .B(A[570]), .Z(n1818) );
  AND U1592 ( .A(n1819), .B(n1820), .Z(n1817) );
  NAND U1593 ( .A(n1821), .B(n1822), .Z(n1820) );
  NANDN U1594 ( .A(A[569]), .B(B[569]), .Z(n1822) );
  AND U1595 ( .A(n1823), .B(n1824), .Z(n1821) );
  NANDN U1596 ( .A(A[568]), .B(B[568]), .Z(n1824) );
  NAND U1597 ( .A(n1825), .B(n1826), .Z(n1823) );
  NANDN U1598 ( .A(B[568]), .B(A[568]), .Z(n1826) );
  AND U1599 ( .A(n1827), .B(n1828), .Z(n1825) );
  NAND U1600 ( .A(n1829), .B(n1830), .Z(n1828) );
  NANDN U1601 ( .A(A[567]), .B(B[567]), .Z(n1830) );
  AND U1602 ( .A(n1831), .B(n1832), .Z(n1829) );
  NANDN U1603 ( .A(A[566]), .B(B[566]), .Z(n1832) );
  NAND U1604 ( .A(n1833), .B(n1834), .Z(n1831) );
  NANDN U1605 ( .A(B[566]), .B(A[566]), .Z(n1834) );
  AND U1606 ( .A(n1835), .B(n1836), .Z(n1833) );
  NAND U1607 ( .A(n1837), .B(n1838), .Z(n1836) );
  NANDN U1608 ( .A(A[565]), .B(B[565]), .Z(n1838) );
  AND U1609 ( .A(n1839), .B(n1840), .Z(n1837) );
  NANDN U1610 ( .A(A[564]), .B(B[564]), .Z(n1840) );
  NAND U1611 ( .A(n1841), .B(n1842), .Z(n1839) );
  NANDN U1612 ( .A(B[564]), .B(A[564]), .Z(n1842) );
  AND U1613 ( .A(n1843), .B(n1844), .Z(n1841) );
  NAND U1614 ( .A(n1845), .B(n1846), .Z(n1844) );
  NANDN U1615 ( .A(A[563]), .B(B[563]), .Z(n1846) );
  AND U1616 ( .A(n1847), .B(n1848), .Z(n1845) );
  NANDN U1617 ( .A(A[562]), .B(B[562]), .Z(n1848) );
  NAND U1618 ( .A(n1849), .B(n1850), .Z(n1847) );
  NANDN U1619 ( .A(B[562]), .B(A[562]), .Z(n1850) );
  AND U1620 ( .A(n1851), .B(n1852), .Z(n1849) );
  NAND U1621 ( .A(n1853), .B(n1854), .Z(n1852) );
  NANDN U1622 ( .A(A[561]), .B(B[561]), .Z(n1854) );
  AND U1623 ( .A(n1855), .B(n1856), .Z(n1853) );
  NANDN U1624 ( .A(A[560]), .B(B[560]), .Z(n1856) );
  NAND U1625 ( .A(n1857), .B(n1858), .Z(n1855) );
  NANDN U1626 ( .A(B[560]), .B(A[560]), .Z(n1858) );
  AND U1627 ( .A(n1859), .B(n1860), .Z(n1857) );
  NAND U1628 ( .A(n1861), .B(n1862), .Z(n1860) );
  NANDN U1629 ( .A(A[559]), .B(B[559]), .Z(n1862) );
  AND U1630 ( .A(n1863), .B(n1864), .Z(n1861) );
  NANDN U1631 ( .A(A[558]), .B(B[558]), .Z(n1864) );
  NAND U1632 ( .A(n1865), .B(n1866), .Z(n1863) );
  NANDN U1633 ( .A(B[558]), .B(A[558]), .Z(n1866) );
  AND U1634 ( .A(n1867), .B(n1868), .Z(n1865) );
  NAND U1635 ( .A(n1869), .B(n1870), .Z(n1868) );
  NANDN U1636 ( .A(A[557]), .B(B[557]), .Z(n1870) );
  AND U1637 ( .A(n1871), .B(n1872), .Z(n1869) );
  NANDN U1638 ( .A(A[556]), .B(B[556]), .Z(n1872) );
  NAND U1639 ( .A(n1873), .B(n1874), .Z(n1871) );
  NANDN U1640 ( .A(B[556]), .B(A[556]), .Z(n1874) );
  AND U1641 ( .A(n1875), .B(n1876), .Z(n1873) );
  NAND U1642 ( .A(n1877), .B(n1878), .Z(n1876) );
  NANDN U1643 ( .A(A[555]), .B(B[555]), .Z(n1878) );
  AND U1644 ( .A(n1879), .B(n1880), .Z(n1877) );
  NANDN U1645 ( .A(A[554]), .B(B[554]), .Z(n1880) );
  NAND U1646 ( .A(n1881), .B(n1882), .Z(n1879) );
  NANDN U1647 ( .A(B[554]), .B(A[554]), .Z(n1882) );
  AND U1648 ( .A(n1883), .B(n1884), .Z(n1881) );
  NAND U1649 ( .A(n1885), .B(n1886), .Z(n1884) );
  NANDN U1650 ( .A(A[553]), .B(B[553]), .Z(n1886) );
  AND U1651 ( .A(n1887), .B(n1888), .Z(n1885) );
  NANDN U1652 ( .A(A[552]), .B(B[552]), .Z(n1888) );
  NAND U1653 ( .A(n1889), .B(n1890), .Z(n1887) );
  NANDN U1654 ( .A(B[552]), .B(A[552]), .Z(n1890) );
  AND U1655 ( .A(n1891), .B(n1892), .Z(n1889) );
  NAND U1656 ( .A(n1893), .B(n1894), .Z(n1892) );
  NANDN U1657 ( .A(A[551]), .B(B[551]), .Z(n1894) );
  AND U1658 ( .A(n1895), .B(n1896), .Z(n1893) );
  NANDN U1659 ( .A(A[550]), .B(B[550]), .Z(n1896) );
  NAND U1660 ( .A(n1897), .B(n1898), .Z(n1895) );
  NANDN U1661 ( .A(B[550]), .B(A[550]), .Z(n1898) );
  AND U1662 ( .A(n1899), .B(n1900), .Z(n1897) );
  NAND U1663 ( .A(n1901), .B(n1902), .Z(n1900) );
  NANDN U1664 ( .A(A[549]), .B(B[549]), .Z(n1902) );
  AND U1665 ( .A(n1903), .B(n1904), .Z(n1901) );
  NANDN U1666 ( .A(A[548]), .B(B[548]), .Z(n1904) );
  NAND U1667 ( .A(n1905), .B(n1906), .Z(n1903) );
  NANDN U1668 ( .A(B[548]), .B(A[548]), .Z(n1906) );
  AND U1669 ( .A(n1907), .B(n1908), .Z(n1905) );
  NAND U1670 ( .A(n1909), .B(n1910), .Z(n1908) );
  NANDN U1671 ( .A(A[547]), .B(B[547]), .Z(n1910) );
  AND U1672 ( .A(n1911), .B(n1912), .Z(n1909) );
  NANDN U1673 ( .A(A[546]), .B(B[546]), .Z(n1912) );
  NAND U1674 ( .A(n1913), .B(n1914), .Z(n1911) );
  NANDN U1675 ( .A(B[546]), .B(A[546]), .Z(n1914) );
  AND U1676 ( .A(n1915), .B(n1916), .Z(n1913) );
  NAND U1677 ( .A(n1917), .B(n1918), .Z(n1916) );
  NANDN U1678 ( .A(A[545]), .B(B[545]), .Z(n1918) );
  AND U1679 ( .A(n1919), .B(n1920), .Z(n1917) );
  NANDN U1680 ( .A(A[544]), .B(B[544]), .Z(n1920) );
  NAND U1681 ( .A(n1921), .B(n1922), .Z(n1919) );
  NANDN U1682 ( .A(B[544]), .B(A[544]), .Z(n1922) );
  AND U1683 ( .A(n1923), .B(n1924), .Z(n1921) );
  NAND U1684 ( .A(n1925), .B(n1926), .Z(n1924) );
  NANDN U1685 ( .A(A[543]), .B(B[543]), .Z(n1926) );
  AND U1686 ( .A(n1927), .B(n1928), .Z(n1925) );
  NANDN U1687 ( .A(A[542]), .B(B[542]), .Z(n1928) );
  NAND U1688 ( .A(n1929), .B(n1930), .Z(n1927) );
  NANDN U1689 ( .A(B[542]), .B(A[542]), .Z(n1930) );
  AND U1690 ( .A(n1931), .B(n1932), .Z(n1929) );
  NAND U1691 ( .A(n1933), .B(n1934), .Z(n1932) );
  NANDN U1692 ( .A(A[541]), .B(B[541]), .Z(n1934) );
  AND U1693 ( .A(n1935), .B(n1936), .Z(n1933) );
  NANDN U1694 ( .A(A[540]), .B(B[540]), .Z(n1936) );
  NAND U1695 ( .A(n1937), .B(n1938), .Z(n1935) );
  NANDN U1696 ( .A(B[540]), .B(A[540]), .Z(n1938) );
  AND U1697 ( .A(n1939), .B(n1940), .Z(n1937) );
  NAND U1698 ( .A(n1941), .B(n1942), .Z(n1940) );
  NANDN U1699 ( .A(A[539]), .B(B[539]), .Z(n1942) );
  AND U1700 ( .A(n1943), .B(n1944), .Z(n1941) );
  NANDN U1701 ( .A(A[538]), .B(B[538]), .Z(n1944) );
  NAND U1702 ( .A(n1945), .B(n1946), .Z(n1943) );
  NANDN U1703 ( .A(B[538]), .B(A[538]), .Z(n1946) );
  AND U1704 ( .A(n1947), .B(n1948), .Z(n1945) );
  NAND U1705 ( .A(n1949), .B(n1950), .Z(n1948) );
  NANDN U1706 ( .A(A[537]), .B(B[537]), .Z(n1950) );
  AND U1707 ( .A(n1951), .B(n1952), .Z(n1949) );
  NANDN U1708 ( .A(A[536]), .B(B[536]), .Z(n1952) );
  NAND U1709 ( .A(n1953), .B(n1954), .Z(n1951) );
  NANDN U1710 ( .A(B[536]), .B(A[536]), .Z(n1954) );
  AND U1711 ( .A(n1955), .B(n1956), .Z(n1953) );
  NAND U1712 ( .A(n1957), .B(n1958), .Z(n1956) );
  NANDN U1713 ( .A(A[535]), .B(B[535]), .Z(n1958) );
  AND U1714 ( .A(n1959), .B(n1960), .Z(n1957) );
  NANDN U1715 ( .A(A[534]), .B(B[534]), .Z(n1960) );
  NAND U1716 ( .A(n1961), .B(n1962), .Z(n1959) );
  NANDN U1717 ( .A(B[534]), .B(A[534]), .Z(n1962) );
  AND U1718 ( .A(n1963), .B(n1964), .Z(n1961) );
  NAND U1719 ( .A(n1965), .B(n1966), .Z(n1964) );
  NANDN U1720 ( .A(A[533]), .B(B[533]), .Z(n1966) );
  AND U1721 ( .A(n1967), .B(n1968), .Z(n1965) );
  NANDN U1722 ( .A(A[532]), .B(B[532]), .Z(n1968) );
  NAND U1723 ( .A(n1969), .B(n1970), .Z(n1967) );
  NANDN U1724 ( .A(B[532]), .B(A[532]), .Z(n1970) );
  AND U1725 ( .A(n1971), .B(n1972), .Z(n1969) );
  NAND U1726 ( .A(n1973), .B(n1974), .Z(n1972) );
  NANDN U1727 ( .A(A[531]), .B(B[531]), .Z(n1974) );
  AND U1728 ( .A(n1975), .B(n1976), .Z(n1973) );
  NANDN U1729 ( .A(A[530]), .B(B[530]), .Z(n1976) );
  NAND U1730 ( .A(n1977), .B(n1978), .Z(n1975) );
  NANDN U1731 ( .A(B[530]), .B(A[530]), .Z(n1978) );
  AND U1732 ( .A(n1979), .B(n1980), .Z(n1977) );
  NAND U1733 ( .A(n1981), .B(n1982), .Z(n1980) );
  NANDN U1734 ( .A(A[529]), .B(B[529]), .Z(n1982) );
  AND U1735 ( .A(n1983), .B(n1984), .Z(n1981) );
  NANDN U1736 ( .A(A[528]), .B(B[528]), .Z(n1984) );
  NAND U1737 ( .A(n1985), .B(n1986), .Z(n1983) );
  NANDN U1738 ( .A(B[528]), .B(A[528]), .Z(n1986) );
  AND U1739 ( .A(n1987), .B(n1988), .Z(n1985) );
  NAND U1740 ( .A(n1989), .B(n1990), .Z(n1988) );
  NANDN U1741 ( .A(A[527]), .B(B[527]), .Z(n1990) );
  AND U1742 ( .A(n1991), .B(n1992), .Z(n1989) );
  NANDN U1743 ( .A(A[526]), .B(B[526]), .Z(n1992) );
  NAND U1744 ( .A(n1993), .B(n1994), .Z(n1991) );
  NANDN U1745 ( .A(B[526]), .B(A[526]), .Z(n1994) );
  AND U1746 ( .A(n1995), .B(n1996), .Z(n1993) );
  NAND U1747 ( .A(n1997), .B(n1998), .Z(n1996) );
  NANDN U1748 ( .A(A[525]), .B(B[525]), .Z(n1998) );
  AND U1749 ( .A(n1999), .B(n2000), .Z(n1997) );
  NANDN U1750 ( .A(A[524]), .B(B[524]), .Z(n2000) );
  NAND U1751 ( .A(n2001), .B(n2002), .Z(n1999) );
  NANDN U1752 ( .A(B[524]), .B(A[524]), .Z(n2002) );
  AND U1753 ( .A(n2003), .B(n2004), .Z(n2001) );
  NAND U1754 ( .A(n2005), .B(n2006), .Z(n2004) );
  NANDN U1755 ( .A(A[523]), .B(B[523]), .Z(n2006) );
  AND U1756 ( .A(n2007), .B(n2008), .Z(n2005) );
  NANDN U1757 ( .A(A[522]), .B(B[522]), .Z(n2008) );
  NAND U1758 ( .A(n2009), .B(n2010), .Z(n2007) );
  NANDN U1759 ( .A(B[522]), .B(A[522]), .Z(n2010) );
  AND U1760 ( .A(n2011), .B(n2012), .Z(n2009) );
  NAND U1761 ( .A(n2013), .B(n2014), .Z(n2012) );
  NANDN U1762 ( .A(A[521]), .B(B[521]), .Z(n2014) );
  AND U1763 ( .A(n2015), .B(n2016), .Z(n2013) );
  NANDN U1764 ( .A(A[520]), .B(B[520]), .Z(n2016) );
  NAND U1765 ( .A(n2017), .B(n2018), .Z(n2015) );
  NANDN U1766 ( .A(B[520]), .B(A[520]), .Z(n2018) );
  AND U1767 ( .A(n2019), .B(n2020), .Z(n2017) );
  NAND U1768 ( .A(n2021), .B(n2022), .Z(n2020) );
  NANDN U1769 ( .A(A[519]), .B(B[519]), .Z(n2022) );
  AND U1770 ( .A(n2023), .B(n2024), .Z(n2021) );
  NANDN U1771 ( .A(A[518]), .B(B[518]), .Z(n2024) );
  NAND U1772 ( .A(n2025), .B(n2026), .Z(n2023) );
  NANDN U1773 ( .A(B[518]), .B(A[518]), .Z(n2026) );
  AND U1774 ( .A(n2027), .B(n2028), .Z(n2025) );
  NAND U1775 ( .A(n2029), .B(n2030), .Z(n2028) );
  NANDN U1776 ( .A(A[517]), .B(B[517]), .Z(n2030) );
  AND U1777 ( .A(n2031), .B(n2032), .Z(n2029) );
  NANDN U1778 ( .A(A[516]), .B(B[516]), .Z(n2032) );
  NAND U1779 ( .A(n2033), .B(n2034), .Z(n2031) );
  NANDN U1780 ( .A(B[516]), .B(A[516]), .Z(n2034) );
  AND U1781 ( .A(n2035), .B(n2036), .Z(n2033) );
  NAND U1782 ( .A(n2037), .B(n2038), .Z(n2036) );
  NANDN U1783 ( .A(A[515]), .B(B[515]), .Z(n2038) );
  AND U1784 ( .A(n2039), .B(n2040), .Z(n2037) );
  NANDN U1785 ( .A(A[514]), .B(B[514]), .Z(n2040) );
  NAND U1786 ( .A(n2041), .B(n2042), .Z(n2039) );
  NANDN U1787 ( .A(B[514]), .B(A[514]), .Z(n2042) );
  AND U1788 ( .A(n2043), .B(n2044), .Z(n2041) );
  NAND U1789 ( .A(n2045), .B(n2046), .Z(n2044) );
  NANDN U1790 ( .A(A[513]), .B(B[513]), .Z(n2046) );
  AND U1791 ( .A(n2047), .B(n2048), .Z(n2045) );
  NANDN U1792 ( .A(A[512]), .B(B[512]), .Z(n2048) );
  NAND U1793 ( .A(n2049), .B(n2050), .Z(n2047) );
  NANDN U1794 ( .A(B[512]), .B(A[512]), .Z(n2050) );
  AND U1795 ( .A(n2051), .B(n2052), .Z(n2049) );
  NAND U1796 ( .A(n2053), .B(n2054), .Z(n2052) );
  NANDN U1797 ( .A(A[511]), .B(B[511]), .Z(n2054) );
  AND U1798 ( .A(n2055), .B(n2056), .Z(n2053) );
  NANDN U1799 ( .A(A[510]), .B(B[510]), .Z(n2056) );
  NAND U1800 ( .A(n2057), .B(n2058), .Z(n2055) );
  NANDN U1801 ( .A(B[510]), .B(A[510]), .Z(n2058) );
  AND U1802 ( .A(n2059), .B(n2060), .Z(n2057) );
  NAND U1803 ( .A(n2061), .B(n2062), .Z(n2060) );
  NANDN U1804 ( .A(A[509]), .B(B[509]), .Z(n2062) );
  AND U1805 ( .A(n2063), .B(n2064), .Z(n2061) );
  NANDN U1806 ( .A(A[508]), .B(B[508]), .Z(n2064) );
  NAND U1807 ( .A(n2065), .B(n2066), .Z(n2063) );
  NANDN U1808 ( .A(B[508]), .B(A[508]), .Z(n2066) );
  AND U1809 ( .A(n2067), .B(n2068), .Z(n2065) );
  NAND U1810 ( .A(n2069), .B(n2070), .Z(n2068) );
  NANDN U1811 ( .A(A[507]), .B(B[507]), .Z(n2070) );
  AND U1812 ( .A(n2071), .B(n2072), .Z(n2069) );
  NANDN U1813 ( .A(A[506]), .B(B[506]), .Z(n2072) );
  NAND U1814 ( .A(n2073), .B(n2074), .Z(n2071) );
  NANDN U1815 ( .A(B[506]), .B(A[506]), .Z(n2074) );
  AND U1816 ( .A(n2075), .B(n2076), .Z(n2073) );
  NAND U1817 ( .A(n2077), .B(n2078), .Z(n2076) );
  NANDN U1818 ( .A(A[505]), .B(B[505]), .Z(n2078) );
  AND U1819 ( .A(n2079), .B(n2080), .Z(n2077) );
  NANDN U1820 ( .A(A[504]), .B(B[504]), .Z(n2080) );
  NAND U1821 ( .A(n2081), .B(n2082), .Z(n2079) );
  NANDN U1822 ( .A(B[504]), .B(A[504]), .Z(n2082) );
  AND U1823 ( .A(n2083), .B(n2084), .Z(n2081) );
  NAND U1824 ( .A(n2085), .B(n2086), .Z(n2084) );
  NANDN U1825 ( .A(A[503]), .B(B[503]), .Z(n2086) );
  AND U1826 ( .A(n2087), .B(n2088), .Z(n2085) );
  NANDN U1827 ( .A(A[502]), .B(B[502]), .Z(n2088) );
  NAND U1828 ( .A(n2089), .B(n2090), .Z(n2087) );
  NANDN U1829 ( .A(B[502]), .B(A[502]), .Z(n2090) );
  AND U1830 ( .A(n2091), .B(n2092), .Z(n2089) );
  NAND U1831 ( .A(n2093), .B(n2094), .Z(n2092) );
  NANDN U1832 ( .A(A[501]), .B(B[501]), .Z(n2094) );
  AND U1833 ( .A(n2095), .B(n2096), .Z(n2093) );
  NANDN U1834 ( .A(A[500]), .B(B[500]), .Z(n2096) );
  NAND U1835 ( .A(n2097), .B(n2098), .Z(n2095) );
  NANDN U1836 ( .A(B[500]), .B(A[500]), .Z(n2098) );
  AND U1837 ( .A(n2099), .B(n2100), .Z(n2097) );
  NAND U1838 ( .A(n2101), .B(n2102), .Z(n2100) );
  NANDN U1839 ( .A(A[499]), .B(B[499]), .Z(n2102) );
  AND U1840 ( .A(n2103), .B(n2104), .Z(n2101) );
  NANDN U1841 ( .A(A[498]), .B(B[498]), .Z(n2104) );
  NAND U1842 ( .A(n2105), .B(n2106), .Z(n2103) );
  NANDN U1843 ( .A(B[498]), .B(A[498]), .Z(n2106) );
  AND U1844 ( .A(n2107), .B(n2108), .Z(n2105) );
  NAND U1845 ( .A(n2109), .B(n2110), .Z(n2108) );
  NANDN U1846 ( .A(A[497]), .B(B[497]), .Z(n2110) );
  AND U1847 ( .A(n2111), .B(n2112), .Z(n2109) );
  NANDN U1848 ( .A(A[496]), .B(B[496]), .Z(n2112) );
  NAND U1849 ( .A(n2113), .B(n2114), .Z(n2111) );
  NANDN U1850 ( .A(B[496]), .B(A[496]), .Z(n2114) );
  AND U1851 ( .A(n2115), .B(n2116), .Z(n2113) );
  NAND U1852 ( .A(n2117), .B(n2118), .Z(n2116) );
  NANDN U1853 ( .A(A[495]), .B(B[495]), .Z(n2118) );
  AND U1854 ( .A(n2119), .B(n2120), .Z(n2117) );
  NANDN U1855 ( .A(A[494]), .B(B[494]), .Z(n2120) );
  NAND U1856 ( .A(n2121), .B(n2122), .Z(n2119) );
  NANDN U1857 ( .A(B[494]), .B(A[494]), .Z(n2122) );
  AND U1858 ( .A(n2123), .B(n2124), .Z(n2121) );
  NAND U1859 ( .A(n2125), .B(n2126), .Z(n2124) );
  NANDN U1860 ( .A(A[493]), .B(B[493]), .Z(n2126) );
  AND U1861 ( .A(n2127), .B(n2128), .Z(n2125) );
  NANDN U1862 ( .A(A[492]), .B(B[492]), .Z(n2128) );
  NAND U1863 ( .A(n2129), .B(n2130), .Z(n2127) );
  NANDN U1864 ( .A(B[492]), .B(A[492]), .Z(n2130) );
  AND U1865 ( .A(n2131), .B(n2132), .Z(n2129) );
  NAND U1866 ( .A(n2133), .B(n2134), .Z(n2132) );
  NANDN U1867 ( .A(A[491]), .B(B[491]), .Z(n2134) );
  AND U1868 ( .A(n2135), .B(n2136), .Z(n2133) );
  NANDN U1869 ( .A(A[490]), .B(B[490]), .Z(n2136) );
  NAND U1870 ( .A(n2137), .B(n2138), .Z(n2135) );
  NANDN U1871 ( .A(B[490]), .B(A[490]), .Z(n2138) );
  AND U1872 ( .A(n2139), .B(n2140), .Z(n2137) );
  NAND U1873 ( .A(n2141), .B(n2142), .Z(n2140) );
  NANDN U1874 ( .A(A[489]), .B(B[489]), .Z(n2142) );
  AND U1875 ( .A(n2143), .B(n2144), .Z(n2141) );
  NANDN U1876 ( .A(A[488]), .B(B[488]), .Z(n2144) );
  NAND U1877 ( .A(n2145), .B(n2146), .Z(n2143) );
  NANDN U1878 ( .A(B[488]), .B(A[488]), .Z(n2146) );
  AND U1879 ( .A(n2147), .B(n2148), .Z(n2145) );
  NAND U1880 ( .A(n2149), .B(n2150), .Z(n2148) );
  NANDN U1881 ( .A(A[487]), .B(B[487]), .Z(n2150) );
  AND U1882 ( .A(n2151), .B(n2152), .Z(n2149) );
  NANDN U1883 ( .A(A[486]), .B(B[486]), .Z(n2152) );
  NAND U1884 ( .A(n2153), .B(n2154), .Z(n2151) );
  NANDN U1885 ( .A(B[486]), .B(A[486]), .Z(n2154) );
  AND U1886 ( .A(n2155), .B(n2156), .Z(n2153) );
  NAND U1887 ( .A(n2157), .B(n2158), .Z(n2156) );
  NANDN U1888 ( .A(A[485]), .B(B[485]), .Z(n2158) );
  AND U1889 ( .A(n2159), .B(n2160), .Z(n2157) );
  NANDN U1890 ( .A(A[484]), .B(B[484]), .Z(n2160) );
  NAND U1891 ( .A(n2161), .B(n2162), .Z(n2159) );
  NANDN U1892 ( .A(B[484]), .B(A[484]), .Z(n2162) );
  AND U1893 ( .A(n2163), .B(n2164), .Z(n2161) );
  NAND U1894 ( .A(n2165), .B(n2166), .Z(n2164) );
  NANDN U1895 ( .A(A[483]), .B(B[483]), .Z(n2166) );
  AND U1896 ( .A(n2167), .B(n2168), .Z(n2165) );
  NANDN U1897 ( .A(A[482]), .B(B[482]), .Z(n2168) );
  NAND U1898 ( .A(n2169), .B(n2170), .Z(n2167) );
  NANDN U1899 ( .A(B[482]), .B(A[482]), .Z(n2170) );
  AND U1900 ( .A(n2171), .B(n2172), .Z(n2169) );
  NAND U1901 ( .A(n2173), .B(n2174), .Z(n2172) );
  NANDN U1902 ( .A(A[481]), .B(B[481]), .Z(n2174) );
  AND U1903 ( .A(n2175), .B(n2176), .Z(n2173) );
  NANDN U1904 ( .A(A[480]), .B(B[480]), .Z(n2176) );
  NAND U1905 ( .A(n2177), .B(n2178), .Z(n2175) );
  NANDN U1906 ( .A(B[480]), .B(A[480]), .Z(n2178) );
  AND U1907 ( .A(n2179), .B(n2180), .Z(n2177) );
  NAND U1908 ( .A(n2181), .B(n2182), .Z(n2180) );
  NANDN U1909 ( .A(A[479]), .B(B[479]), .Z(n2182) );
  AND U1910 ( .A(n2183), .B(n2184), .Z(n2181) );
  NANDN U1911 ( .A(A[478]), .B(B[478]), .Z(n2184) );
  NAND U1912 ( .A(n2185), .B(n2186), .Z(n2183) );
  NANDN U1913 ( .A(B[478]), .B(A[478]), .Z(n2186) );
  AND U1914 ( .A(n2187), .B(n2188), .Z(n2185) );
  NAND U1915 ( .A(n2189), .B(n2190), .Z(n2188) );
  NANDN U1916 ( .A(A[477]), .B(B[477]), .Z(n2190) );
  AND U1917 ( .A(n2191), .B(n2192), .Z(n2189) );
  NANDN U1918 ( .A(A[476]), .B(B[476]), .Z(n2192) );
  NAND U1919 ( .A(n2193), .B(n2194), .Z(n2191) );
  NANDN U1920 ( .A(B[476]), .B(A[476]), .Z(n2194) );
  AND U1921 ( .A(n2195), .B(n2196), .Z(n2193) );
  NAND U1922 ( .A(n2197), .B(n2198), .Z(n2196) );
  NANDN U1923 ( .A(A[475]), .B(B[475]), .Z(n2198) );
  AND U1924 ( .A(n2199), .B(n2200), .Z(n2197) );
  NANDN U1925 ( .A(A[474]), .B(B[474]), .Z(n2200) );
  NAND U1926 ( .A(n2201), .B(n2202), .Z(n2199) );
  NANDN U1927 ( .A(B[474]), .B(A[474]), .Z(n2202) );
  AND U1928 ( .A(n2203), .B(n2204), .Z(n2201) );
  NAND U1929 ( .A(n2205), .B(n2206), .Z(n2204) );
  NANDN U1930 ( .A(A[473]), .B(B[473]), .Z(n2206) );
  AND U1931 ( .A(n2207), .B(n2208), .Z(n2205) );
  NANDN U1932 ( .A(A[472]), .B(B[472]), .Z(n2208) );
  NAND U1933 ( .A(n2209), .B(n2210), .Z(n2207) );
  NANDN U1934 ( .A(B[472]), .B(A[472]), .Z(n2210) );
  AND U1935 ( .A(n2211), .B(n2212), .Z(n2209) );
  NAND U1936 ( .A(n2213), .B(n2214), .Z(n2212) );
  NANDN U1937 ( .A(A[471]), .B(B[471]), .Z(n2214) );
  AND U1938 ( .A(n2215), .B(n2216), .Z(n2213) );
  NANDN U1939 ( .A(A[470]), .B(B[470]), .Z(n2216) );
  NAND U1940 ( .A(n2217), .B(n2218), .Z(n2215) );
  NANDN U1941 ( .A(B[470]), .B(A[470]), .Z(n2218) );
  AND U1942 ( .A(n2219), .B(n2220), .Z(n2217) );
  NAND U1943 ( .A(n2221), .B(n2222), .Z(n2220) );
  NANDN U1944 ( .A(A[469]), .B(B[469]), .Z(n2222) );
  AND U1945 ( .A(n2223), .B(n2224), .Z(n2221) );
  NANDN U1946 ( .A(A[468]), .B(B[468]), .Z(n2224) );
  NAND U1947 ( .A(n2225), .B(n2226), .Z(n2223) );
  NANDN U1948 ( .A(B[468]), .B(A[468]), .Z(n2226) );
  AND U1949 ( .A(n2227), .B(n2228), .Z(n2225) );
  NAND U1950 ( .A(n2229), .B(n2230), .Z(n2228) );
  NANDN U1951 ( .A(A[467]), .B(B[467]), .Z(n2230) );
  AND U1952 ( .A(n2231), .B(n2232), .Z(n2229) );
  NANDN U1953 ( .A(A[466]), .B(B[466]), .Z(n2232) );
  NAND U1954 ( .A(n2233), .B(n2234), .Z(n2231) );
  NANDN U1955 ( .A(B[466]), .B(A[466]), .Z(n2234) );
  AND U1956 ( .A(n2235), .B(n2236), .Z(n2233) );
  NAND U1957 ( .A(n2237), .B(n2238), .Z(n2236) );
  NANDN U1958 ( .A(A[465]), .B(B[465]), .Z(n2238) );
  AND U1959 ( .A(n2239), .B(n2240), .Z(n2237) );
  NANDN U1960 ( .A(A[464]), .B(B[464]), .Z(n2240) );
  NAND U1961 ( .A(n2241), .B(n2242), .Z(n2239) );
  NANDN U1962 ( .A(B[464]), .B(A[464]), .Z(n2242) );
  AND U1963 ( .A(n2243), .B(n2244), .Z(n2241) );
  NAND U1964 ( .A(n2245), .B(n2246), .Z(n2244) );
  NANDN U1965 ( .A(A[463]), .B(B[463]), .Z(n2246) );
  AND U1966 ( .A(n2247), .B(n2248), .Z(n2245) );
  NANDN U1967 ( .A(A[462]), .B(B[462]), .Z(n2248) );
  NAND U1968 ( .A(n2249), .B(n2250), .Z(n2247) );
  NANDN U1969 ( .A(B[462]), .B(A[462]), .Z(n2250) );
  AND U1970 ( .A(n2251), .B(n2252), .Z(n2249) );
  NAND U1971 ( .A(n2253), .B(n2254), .Z(n2252) );
  NANDN U1972 ( .A(A[461]), .B(B[461]), .Z(n2254) );
  AND U1973 ( .A(n2255), .B(n2256), .Z(n2253) );
  NANDN U1974 ( .A(A[460]), .B(B[460]), .Z(n2256) );
  NAND U1975 ( .A(n2257), .B(n2258), .Z(n2255) );
  NANDN U1976 ( .A(B[460]), .B(A[460]), .Z(n2258) );
  AND U1977 ( .A(n2259), .B(n2260), .Z(n2257) );
  NAND U1978 ( .A(n2261), .B(n2262), .Z(n2260) );
  NANDN U1979 ( .A(A[459]), .B(B[459]), .Z(n2262) );
  AND U1980 ( .A(n2263), .B(n2264), .Z(n2261) );
  NANDN U1981 ( .A(A[458]), .B(B[458]), .Z(n2264) );
  NAND U1982 ( .A(n2265), .B(n2266), .Z(n2263) );
  NANDN U1983 ( .A(B[458]), .B(A[458]), .Z(n2266) );
  AND U1984 ( .A(n2267), .B(n2268), .Z(n2265) );
  NAND U1985 ( .A(n2269), .B(n2270), .Z(n2268) );
  NANDN U1986 ( .A(A[457]), .B(B[457]), .Z(n2270) );
  AND U1987 ( .A(n2271), .B(n2272), .Z(n2269) );
  NANDN U1988 ( .A(A[456]), .B(B[456]), .Z(n2272) );
  NAND U1989 ( .A(n2273), .B(n2274), .Z(n2271) );
  NANDN U1990 ( .A(B[456]), .B(A[456]), .Z(n2274) );
  AND U1991 ( .A(n2275), .B(n2276), .Z(n2273) );
  NAND U1992 ( .A(n2277), .B(n2278), .Z(n2276) );
  NANDN U1993 ( .A(A[455]), .B(B[455]), .Z(n2278) );
  AND U1994 ( .A(n2279), .B(n2280), .Z(n2277) );
  NANDN U1995 ( .A(A[454]), .B(B[454]), .Z(n2280) );
  NAND U1996 ( .A(n2281), .B(n2282), .Z(n2279) );
  NANDN U1997 ( .A(B[454]), .B(A[454]), .Z(n2282) );
  AND U1998 ( .A(n2283), .B(n2284), .Z(n2281) );
  NAND U1999 ( .A(n2285), .B(n2286), .Z(n2284) );
  NANDN U2000 ( .A(A[453]), .B(B[453]), .Z(n2286) );
  AND U2001 ( .A(n2287), .B(n2288), .Z(n2285) );
  NANDN U2002 ( .A(A[452]), .B(B[452]), .Z(n2288) );
  NAND U2003 ( .A(n2289), .B(n2290), .Z(n2287) );
  NANDN U2004 ( .A(B[452]), .B(A[452]), .Z(n2290) );
  AND U2005 ( .A(n2291), .B(n2292), .Z(n2289) );
  NAND U2006 ( .A(n2293), .B(n2294), .Z(n2292) );
  NANDN U2007 ( .A(A[451]), .B(B[451]), .Z(n2294) );
  AND U2008 ( .A(n2295), .B(n2296), .Z(n2293) );
  NANDN U2009 ( .A(A[450]), .B(B[450]), .Z(n2296) );
  NAND U2010 ( .A(n2297), .B(n2298), .Z(n2295) );
  NANDN U2011 ( .A(B[450]), .B(A[450]), .Z(n2298) );
  AND U2012 ( .A(n2299), .B(n2300), .Z(n2297) );
  NAND U2013 ( .A(n2301), .B(n2302), .Z(n2300) );
  NANDN U2014 ( .A(A[449]), .B(B[449]), .Z(n2302) );
  AND U2015 ( .A(n2303), .B(n2304), .Z(n2301) );
  NANDN U2016 ( .A(A[448]), .B(B[448]), .Z(n2304) );
  NAND U2017 ( .A(n2305), .B(n2306), .Z(n2303) );
  NANDN U2018 ( .A(B[448]), .B(A[448]), .Z(n2306) );
  AND U2019 ( .A(n2307), .B(n2308), .Z(n2305) );
  NAND U2020 ( .A(n2309), .B(n2310), .Z(n2308) );
  NANDN U2021 ( .A(A[447]), .B(B[447]), .Z(n2310) );
  AND U2022 ( .A(n2311), .B(n2312), .Z(n2309) );
  NANDN U2023 ( .A(A[446]), .B(B[446]), .Z(n2312) );
  NAND U2024 ( .A(n2313), .B(n2314), .Z(n2311) );
  NANDN U2025 ( .A(B[446]), .B(A[446]), .Z(n2314) );
  AND U2026 ( .A(n2315), .B(n2316), .Z(n2313) );
  NAND U2027 ( .A(n2317), .B(n2318), .Z(n2316) );
  NANDN U2028 ( .A(A[445]), .B(B[445]), .Z(n2318) );
  AND U2029 ( .A(n2319), .B(n2320), .Z(n2317) );
  NANDN U2030 ( .A(A[444]), .B(B[444]), .Z(n2320) );
  NAND U2031 ( .A(n2321), .B(n2322), .Z(n2319) );
  NANDN U2032 ( .A(B[444]), .B(A[444]), .Z(n2322) );
  AND U2033 ( .A(n2323), .B(n2324), .Z(n2321) );
  NAND U2034 ( .A(n2325), .B(n2326), .Z(n2324) );
  NANDN U2035 ( .A(A[443]), .B(B[443]), .Z(n2326) );
  AND U2036 ( .A(n2327), .B(n2328), .Z(n2325) );
  NANDN U2037 ( .A(A[442]), .B(B[442]), .Z(n2328) );
  NAND U2038 ( .A(n2329), .B(n2330), .Z(n2327) );
  NANDN U2039 ( .A(B[442]), .B(A[442]), .Z(n2330) );
  AND U2040 ( .A(n2331), .B(n2332), .Z(n2329) );
  NAND U2041 ( .A(n2333), .B(n2334), .Z(n2332) );
  NANDN U2042 ( .A(A[441]), .B(B[441]), .Z(n2334) );
  AND U2043 ( .A(n2335), .B(n2336), .Z(n2333) );
  NANDN U2044 ( .A(A[440]), .B(B[440]), .Z(n2336) );
  NAND U2045 ( .A(n2337), .B(n2338), .Z(n2335) );
  NANDN U2046 ( .A(B[440]), .B(A[440]), .Z(n2338) );
  AND U2047 ( .A(n2339), .B(n2340), .Z(n2337) );
  NAND U2048 ( .A(n2341), .B(n2342), .Z(n2340) );
  NANDN U2049 ( .A(A[439]), .B(B[439]), .Z(n2342) );
  AND U2050 ( .A(n2343), .B(n2344), .Z(n2341) );
  NANDN U2051 ( .A(A[438]), .B(B[438]), .Z(n2344) );
  NAND U2052 ( .A(n2345), .B(n2346), .Z(n2343) );
  NANDN U2053 ( .A(B[438]), .B(A[438]), .Z(n2346) );
  AND U2054 ( .A(n2347), .B(n2348), .Z(n2345) );
  NAND U2055 ( .A(n2349), .B(n2350), .Z(n2348) );
  NANDN U2056 ( .A(A[437]), .B(B[437]), .Z(n2350) );
  AND U2057 ( .A(n2351), .B(n2352), .Z(n2349) );
  NANDN U2058 ( .A(A[436]), .B(B[436]), .Z(n2352) );
  NAND U2059 ( .A(n2353), .B(n2354), .Z(n2351) );
  NANDN U2060 ( .A(B[436]), .B(A[436]), .Z(n2354) );
  AND U2061 ( .A(n2355), .B(n2356), .Z(n2353) );
  NAND U2062 ( .A(n2357), .B(n2358), .Z(n2356) );
  NANDN U2063 ( .A(A[435]), .B(B[435]), .Z(n2358) );
  AND U2064 ( .A(n2359), .B(n2360), .Z(n2357) );
  NANDN U2065 ( .A(A[434]), .B(B[434]), .Z(n2360) );
  NAND U2066 ( .A(n2361), .B(n2362), .Z(n2359) );
  NANDN U2067 ( .A(B[434]), .B(A[434]), .Z(n2362) );
  AND U2068 ( .A(n2363), .B(n2364), .Z(n2361) );
  NAND U2069 ( .A(n2365), .B(n2366), .Z(n2364) );
  NANDN U2070 ( .A(A[433]), .B(B[433]), .Z(n2366) );
  AND U2071 ( .A(n2367), .B(n2368), .Z(n2365) );
  NANDN U2072 ( .A(A[432]), .B(B[432]), .Z(n2368) );
  NAND U2073 ( .A(n2369), .B(n2370), .Z(n2367) );
  NANDN U2074 ( .A(B[432]), .B(A[432]), .Z(n2370) );
  AND U2075 ( .A(n2371), .B(n2372), .Z(n2369) );
  NAND U2076 ( .A(n2373), .B(n2374), .Z(n2372) );
  NANDN U2077 ( .A(A[431]), .B(B[431]), .Z(n2374) );
  AND U2078 ( .A(n2375), .B(n2376), .Z(n2373) );
  NANDN U2079 ( .A(A[430]), .B(B[430]), .Z(n2376) );
  NAND U2080 ( .A(n2377), .B(n2378), .Z(n2375) );
  NANDN U2081 ( .A(B[430]), .B(A[430]), .Z(n2378) );
  AND U2082 ( .A(n2379), .B(n2380), .Z(n2377) );
  NAND U2083 ( .A(n2381), .B(n2382), .Z(n2380) );
  NANDN U2084 ( .A(A[429]), .B(B[429]), .Z(n2382) );
  AND U2085 ( .A(n2383), .B(n2384), .Z(n2381) );
  NANDN U2086 ( .A(A[428]), .B(B[428]), .Z(n2384) );
  NAND U2087 ( .A(n2385), .B(n2386), .Z(n2383) );
  NANDN U2088 ( .A(B[428]), .B(A[428]), .Z(n2386) );
  AND U2089 ( .A(n2387), .B(n2388), .Z(n2385) );
  NAND U2090 ( .A(n2389), .B(n2390), .Z(n2388) );
  NANDN U2091 ( .A(A[427]), .B(B[427]), .Z(n2390) );
  AND U2092 ( .A(n2391), .B(n2392), .Z(n2389) );
  NANDN U2093 ( .A(A[426]), .B(B[426]), .Z(n2392) );
  NAND U2094 ( .A(n2393), .B(n2394), .Z(n2391) );
  NANDN U2095 ( .A(B[426]), .B(A[426]), .Z(n2394) );
  AND U2096 ( .A(n2395), .B(n2396), .Z(n2393) );
  NAND U2097 ( .A(n2397), .B(n2398), .Z(n2396) );
  NANDN U2098 ( .A(A[425]), .B(B[425]), .Z(n2398) );
  AND U2099 ( .A(n2399), .B(n2400), .Z(n2397) );
  NANDN U2100 ( .A(A[424]), .B(B[424]), .Z(n2400) );
  NAND U2101 ( .A(n2401), .B(n2402), .Z(n2399) );
  NANDN U2102 ( .A(B[424]), .B(A[424]), .Z(n2402) );
  AND U2103 ( .A(n2403), .B(n2404), .Z(n2401) );
  NAND U2104 ( .A(n2405), .B(n2406), .Z(n2404) );
  NANDN U2105 ( .A(A[423]), .B(B[423]), .Z(n2406) );
  AND U2106 ( .A(n2407), .B(n2408), .Z(n2405) );
  NANDN U2107 ( .A(A[422]), .B(B[422]), .Z(n2408) );
  NAND U2108 ( .A(n2409), .B(n2410), .Z(n2407) );
  NANDN U2109 ( .A(B[422]), .B(A[422]), .Z(n2410) );
  AND U2110 ( .A(n2411), .B(n2412), .Z(n2409) );
  NAND U2111 ( .A(n2413), .B(n2414), .Z(n2412) );
  NANDN U2112 ( .A(A[421]), .B(B[421]), .Z(n2414) );
  AND U2113 ( .A(n2415), .B(n2416), .Z(n2413) );
  NANDN U2114 ( .A(A[420]), .B(B[420]), .Z(n2416) );
  NAND U2115 ( .A(n2417), .B(n2418), .Z(n2415) );
  NANDN U2116 ( .A(B[420]), .B(A[420]), .Z(n2418) );
  AND U2117 ( .A(n2419), .B(n2420), .Z(n2417) );
  NAND U2118 ( .A(n2421), .B(n2422), .Z(n2420) );
  NANDN U2119 ( .A(A[419]), .B(B[419]), .Z(n2422) );
  AND U2120 ( .A(n2423), .B(n2424), .Z(n2421) );
  NANDN U2121 ( .A(A[418]), .B(B[418]), .Z(n2424) );
  NAND U2122 ( .A(n2425), .B(n2426), .Z(n2423) );
  NANDN U2123 ( .A(B[418]), .B(A[418]), .Z(n2426) );
  AND U2124 ( .A(n2427), .B(n2428), .Z(n2425) );
  NAND U2125 ( .A(n2429), .B(n2430), .Z(n2428) );
  NANDN U2126 ( .A(A[417]), .B(B[417]), .Z(n2430) );
  AND U2127 ( .A(n2431), .B(n2432), .Z(n2429) );
  NANDN U2128 ( .A(A[416]), .B(B[416]), .Z(n2432) );
  NAND U2129 ( .A(n2433), .B(n2434), .Z(n2431) );
  NANDN U2130 ( .A(B[416]), .B(A[416]), .Z(n2434) );
  AND U2131 ( .A(n2435), .B(n2436), .Z(n2433) );
  NAND U2132 ( .A(n2437), .B(n2438), .Z(n2436) );
  NANDN U2133 ( .A(A[415]), .B(B[415]), .Z(n2438) );
  AND U2134 ( .A(n2439), .B(n2440), .Z(n2437) );
  NANDN U2135 ( .A(A[414]), .B(B[414]), .Z(n2440) );
  NAND U2136 ( .A(n2441), .B(n2442), .Z(n2439) );
  NANDN U2137 ( .A(B[414]), .B(A[414]), .Z(n2442) );
  AND U2138 ( .A(n2443), .B(n2444), .Z(n2441) );
  NAND U2139 ( .A(n2445), .B(n2446), .Z(n2444) );
  NANDN U2140 ( .A(A[413]), .B(B[413]), .Z(n2446) );
  AND U2141 ( .A(n2447), .B(n2448), .Z(n2445) );
  NANDN U2142 ( .A(A[412]), .B(B[412]), .Z(n2448) );
  NAND U2143 ( .A(n2449), .B(n2450), .Z(n2447) );
  NANDN U2144 ( .A(B[412]), .B(A[412]), .Z(n2450) );
  AND U2145 ( .A(n2451), .B(n2452), .Z(n2449) );
  NAND U2146 ( .A(n2453), .B(n2454), .Z(n2452) );
  NANDN U2147 ( .A(A[411]), .B(B[411]), .Z(n2454) );
  AND U2148 ( .A(n2455), .B(n2456), .Z(n2453) );
  NANDN U2149 ( .A(A[410]), .B(B[410]), .Z(n2456) );
  NAND U2150 ( .A(n2457), .B(n2458), .Z(n2455) );
  NANDN U2151 ( .A(B[410]), .B(A[410]), .Z(n2458) );
  AND U2152 ( .A(n2459), .B(n2460), .Z(n2457) );
  NAND U2153 ( .A(n2461), .B(n2462), .Z(n2460) );
  NANDN U2154 ( .A(A[409]), .B(B[409]), .Z(n2462) );
  AND U2155 ( .A(n2463), .B(n2464), .Z(n2461) );
  NANDN U2156 ( .A(A[408]), .B(B[408]), .Z(n2464) );
  NAND U2157 ( .A(n2465), .B(n2466), .Z(n2463) );
  NANDN U2158 ( .A(B[408]), .B(A[408]), .Z(n2466) );
  AND U2159 ( .A(n2467), .B(n2468), .Z(n2465) );
  NAND U2160 ( .A(n2469), .B(n2470), .Z(n2468) );
  NANDN U2161 ( .A(A[407]), .B(B[407]), .Z(n2470) );
  AND U2162 ( .A(n2471), .B(n2472), .Z(n2469) );
  NANDN U2163 ( .A(A[406]), .B(B[406]), .Z(n2472) );
  NAND U2164 ( .A(n2473), .B(n2474), .Z(n2471) );
  NANDN U2165 ( .A(B[406]), .B(A[406]), .Z(n2474) );
  AND U2166 ( .A(n2475), .B(n2476), .Z(n2473) );
  NAND U2167 ( .A(n2477), .B(n2478), .Z(n2476) );
  NANDN U2168 ( .A(A[405]), .B(B[405]), .Z(n2478) );
  AND U2169 ( .A(n2479), .B(n2480), .Z(n2477) );
  NANDN U2170 ( .A(A[404]), .B(B[404]), .Z(n2480) );
  NAND U2171 ( .A(n2481), .B(n2482), .Z(n2479) );
  NANDN U2172 ( .A(B[404]), .B(A[404]), .Z(n2482) );
  AND U2173 ( .A(n2483), .B(n2484), .Z(n2481) );
  NAND U2174 ( .A(n2485), .B(n2486), .Z(n2484) );
  NANDN U2175 ( .A(A[403]), .B(B[403]), .Z(n2486) );
  AND U2176 ( .A(n2487), .B(n2488), .Z(n2485) );
  NANDN U2177 ( .A(A[402]), .B(B[402]), .Z(n2488) );
  NAND U2178 ( .A(n2489), .B(n2490), .Z(n2487) );
  NANDN U2179 ( .A(B[402]), .B(A[402]), .Z(n2490) );
  AND U2180 ( .A(n2491), .B(n2492), .Z(n2489) );
  NAND U2181 ( .A(n2493), .B(n2494), .Z(n2492) );
  NANDN U2182 ( .A(A[401]), .B(B[401]), .Z(n2494) );
  AND U2183 ( .A(n2495), .B(n2496), .Z(n2493) );
  NANDN U2184 ( .A(A[400]), .B(B[400]), .Z(n2496) );
  NAND U2185 ( .A(n2497), .B(n2498), .Z(n2495) );
  NANDN U2186 ( .A(B[400]), .B(A[400]), .Z(n2498) );
  AND U2187 ( .A(n2499), .B(n2500), .Z(n2497) );
  NAND U2188 ( .A(n2501), .B(n2502), .Z(n2500) );
  NANDN U2189 ( .A(A[399]), .B(B[399]), .Z(n2502) );
  AND U2190 ( .A(n2503), .B(n2504), .Z(n2501) );
  NANDN U2191 ( .A(A[398]), .B(B[398]), .Z(n2504) );
  NAND U2192 ( .A(n2505), .B(n2506), .Z(n2503) );
  NANDN U2193 ( .A(B[398]), .B(A[398]), .Z(n2506) );
  AND U2194 ( .A(n2507), .B(n2508), .Z(n2505) );
  NAND U2195 ( .A(n2509), .B(n2510), .Z(n2508) );
  NANDN U2196 ( .A(A[397]), .B(B[397]), .Z(n2510) );
  AND U2197 ( .A(n2511), .B(n2512), .Z(n2509) );
  NANDN U2198 ( .A(A[396]), .B(B[396]), .Z(n2512) );
  NAND U2199 ( .A(n2513), .B(n2514), .Z(n2511) );
  NANDN U2200 ( .A(B[396]), .B(A[396]), .Z(n2514) );
  AND U2201 ( .A(n2515), .B(n2516), .Z(n2513) );
  NAND U2202 ( .A(n2517), .B(n2518), .Z(n2516) );
  NANDN U2203 ( .A(A[395]), .B(B[395]), .Z(n2518) );
  AND U2204 ( .A(n2519), .B(n2520), .Z(n2517) );
  NANDN U2205 ( .A(A[394]), .B(B[394]), .Z(n2520) );
  NAND U2206 ( .A(n2521), .B(n2522), .Z(n2519) );
  NANDN U2207 ( .A(B[394]), .B(A[394]), .Z(n2522) );
  AND U2208 ( .A(n2523), .B(n2524), .Z(n2521) );
  NAND U2209 ( .A(n2525), .B(n2526), .Z(n2524) );
  NANDN U2210 ( .A(A[393]), .B(B[393]), .Z(n2526) );
  AND U2211 ( .A(n2527), .B(n2528), .Z(n2525) );
  NANDN U2212 ( .A(A[392]), .B(B[392]), .Z(n2528) );
  NAND U2213 ( .A(n2529), .B(n2530), .Z(n2527) );
  NANDN U2214 ( .A(B[392]), .B(A[392]), .Z(n2530) );
  AND U2215 ( .A(n2531), .B(n2532), .Z(n2529) );
  NAND U2216 ( .A(n2533), .B(n2534), .Z(n2532) );
  NANDN U2217 ( .A(A[391]), .B(B[391]), .Z(n2534) );
  AND U2218 ( .A(n2535), .B(n2536), .Z(n2533) );
  NANDN U2219 ( .A(A[390]), .B(B[390]), .Z(n2536) );
  NAND U2220 ( .A(n2537), .B(n2538), .Z(n2535) );
  NANDN U2221 ( .A(B[390]), .B(A[390]), .Z(n2538) );
  AND U2222 ( .A(n2539), .B(n2540), .Z(n2537) );
  NAND U2223 ( .A(n2541), .B(n2542), .Z(n2540) );
  NANDN U2224 ( .A(A[389]), .B(B[389]), .Z(n2542) );
  AND U2225 ( .A(n2543), .B(n2544), .Z(n2541) );
  NANDN U2226 ( .A(A[388]), .B(B[388]), .Z(n2544) );
  NAND U2227 ( .A(n2545), .B(n2546), .Z(n2543) );
  NANDN U2228 ( .A(B[388]), .B(A[388]), .Z(n2546) );
  AND U2229 ( .A(n2547), .B(n2548), .Z(n2545) );
  NAND U2230 ( .A(n2549), .B(n2550), .Z(n2548) );
  NANDN U2231 ( .A(A[387]), .B(B[387]), .Z(n2550) );
  AND U2232 ( .A(n2551), .B(n2552), .Z(n2549) );
  NANDN U2233 ( .A(A[386]), .B(B[386]), .Z(n2552) );
  NAND U2234 ( .A(n2553), .B(n2554), .Z(n2551) );
  NANDN U2235 ( .A(B[386]), .B(A[386]), .Z(n2554) );
  AND U2236 ( .A(n2555), .B(n2556), .Z(n2553) );
  NAND U2237 ( .A(n2557), .B(n2558), .Z(n2556) );
  NANDN U2238 ( .A(A[385]), .B(B[385]), .Z(n2558) );
  AND U2239 ( .A(n2559), .B(n2560), .Z(n2557) );
  NANDN U2240 ( .A(A[384]), .B(B[384]), .Z(n2560) );
  NAND U2241 ( .A(n2561), .B(n2562), .Z(n2559) );
  NANDN U2242 ( .A(B[384]), .B(A[384]), .Z(n2562) );
  AND U2243 ( .A(n2563), .B(n2564), .Z(n2561) );
  NAND U2244 ( .A(n2565), .B(n2566), .Z(n2564) );
  NANDN U2245 ( .A(A[383]), .B(B[383]), .Z(n2566) );
  AND U2246 ( .A(n2567), .B(n2568), .Z(n2565) );
  NANDN U2247 ( .A(A[382]), .B(B[382]), .Z(n2568) );
  NAND U2248 ( .A(n2569), .B(n2570), .Z(n2567) );
  NANDN U2249 ( .A(B[382]), .B(A[382]), .Z(n2570) );
  AND U2250 ( .A(n2571), .B(n2572), .Z(n2569) );
  NAND U2251 ( .A(n2573), .B(n2574), .Z(n2572) );
  NANDN U2252 ( .A(A[381]), .B(B[381]), .Z(n2574) );
  AND U2253 ( .A(n2575), .B(n2576), .Z(n2573) );
  NANDN U2254 ( .A(A[380]), .B(B[380]), .Z(n2576) );
  NAND U2255 ( .A(n2577), .B(n2578), .Z(n2575) );
  NANDN U2256 ( .A(B[380]), .B(A[380]), .Z(n2578) );
  AND U2257 ( .A(n2579), .B(n2580), .Z(n2577) );
  NAND U2258 ( .A(n2581), .B(n2582), .Z(n2580) );
  NANDN U2259 ( .A(A[379]), .B(B[379]), .Z(n2582) );
  AND U2260 ( .A(n2583), .B(n2584), .Z(n2581) );
  NANDN U2261 ( .A(A[378]), .B(B[378]), .Z(n2584) );
  NAND U2262 ( .A(n2585), .B(n2586), .Z(n2583) );
  NANDN U2263 ( .A(B[378]), .B(A[378]), .Z(n2586) );
  AND U2264 ( .A(n2587), .B(n2588), .Z(n2585) );
  NAND U2265 ( .A(n2589), .B(n2590), .Z(n2588) );
  NANDN U2266 ( .A(A[377]), .B(B[377]), .Z(n2590) );
  AND U2267 ( .A(n2591), .B(n2592), .Z(n2589) );
  NANDN U2268 ( .A(A[376]), .B(B[376]), .Z(n2592) );
  NAND U2269 ( .A(n2593), .B(n2594), .Z(n2591) );
  NANDN U2270 ( .A(B[376]), .B(A[376]), .Z(n2594) );
  AND U2271 ( .A(n2595), .B(n2596), .Z(n2593) );
  NAND U2272 ( .A(n2597), .B(n2598), .Z(n2596) );
  NANDN U2273 ( .A(A[375]), .B(B[375]), .Z(n2598) );
  AND U2274 ( .A(n2599), .B(n2600), .Z(n2597) );
  NANDN U2275 ( .A(A[374]), .B(B[374]), .Z(n2600) );
  NAND U2276 ( .A(n2601), .B(n2602), .Z(n2599) );
  NANDN U2277 ( .A(B[374]), .B(A[374]), .Z(n2602) );
  AND U2278 ( .A(n2603), .B(n2604), .Z(n2601) );
  NAND U2279 ( .A(n2605), .B(n2606), .Z(n2604) );
  NANDN U2280 ( .A(A[373]), .B(B[373]), .Z(n2606) );
  AND U2281 ( .A(n2607), .B(n2608), .Z(n2605) );
  NANDN U2282 ( .A(A[372]), .B(B[372]), .Z(n2608) );
  NAND U2283 ( .A(n2609), .B(n2610), .Z(n2607) );
  NANDN U2284 ( .A(B[372]), .B(A[372]), .Z(n2610) );
  AND U2285 ( .A(n2611), .B(n2612), .Z(n2609) );
  NAND U2286 ( .A(n2613), .B(n2614), .Z(n2612) );
  NANDN U2287 ( .A(A[371]), .B(B[371]), .Z(n2614) );
  AND U2288 ( .A(n2615), .B(n2616), .Z(n2613) );
  NANDN U2289 ( .A(A[370]), .B(B[370]), .Z(n2616) );
  NAND U2290 ( .A(n2617), .B(n2618), .Z(n2615) );
  NANDN U2291 ( .A(B[370]), .B(A[370]), .Z(n2618) );
  AND U2292 ( .A(n2619), .B(n2620), .Z(n2617) );
  NAND U2293 ( .A(n2621), .B(n2622), .Z(n2620) );
  NANDN U2294 ( .A(A[369]), .B(B[369]), .Z(n2622) );
  AND U2295 ( .A(n2623), .B(n2624), .Z(n2621) );
  NANDN U2296 ( .A(A[368]), .B(B[368]), .Z(n2624) );
  NAND U2297 ( .A(n2625), .B(n2626), .Z(n2623) );
  NANDN U2298 ( .A(B[368]), .B(A[368]), .Z(n2626) );
  AND U2299 ( .A(n2627), .B(n2628), .Z(n2625) );
  NAND U2300 ( .A(n2629), .B(n2630), .Z(n2628) );
  NANDN U2301 ( .A(A[367]), .B(B[367]), .Z(n2630) );
  AND U2302 ( .A(n2631), .B(n2632), .Z(n2629) );
  NANDN U2303 ( .A(A[366]), .B(B[366]), .Z(n2632) );
  NAND U2304 ( .A(n2633), .B(n2634), .Z(n2631) );
  NANDN U2305 ( .A(B[366]), .B(A[366]), .Z(n2634) );
  AND U2306 ( .A(n2635), .B(n2636), .Z(n2633) );
  NAND U2307 ( .A(n2637), .B(n2638), .Z(n2636) );
  NANDN U2308 ( .A(A[365]), .B(B[365]), .Z(n2638) );
  AND U2309 ( .A(n2639), .B(n2640), .Z(n2637) );
  NANDN U2310 ( .A(A[364]), .B(B[364]), .Z(n2640) );
  NAND U2311 ( .A(n2641), .B(n2642), .Z(n2639) );
  NANDN U2312 ( .A(B[364]), .B(A[364]), .Z(n2642) );
  AND U2313 ( .A(n2643), .B(n2644), .Z(n2641) );
  NAND U2314 ( .A(n2645), .B(n2646), .Z(n2644) );
  NANDN U2315 ( .A(A[363]), .B(B[363]), .Z(n2646) );
  AND U2316 ( .A(n2647), .B(n2648), .Z(n2645) );
  NANDN U2317 ( .A(A[362]), .B(B[362]), .Z(n2648) );
  NAND U2318 ( .A(n2649), .B(n2650), .Z(n2647) );
  NANDN U2319 ( .A(B[362]), .B(A[362]), .Z(n2650) );
  AND U2320 ( .A(n2651), .B(n2652), .Z(n2649) );
  NAND U2321 ( .A(n2653), .B(n2654), .Z(n2652) );
  NANDN U2322 ( .A(A[361]), .B(B[361]), .Z(n2654) );
  AND U2323 ( .A(n2655), .B(n2656), .Z(n2653) );
  NANDN U2324 ( .A(A[360]), .B(B[360]), .Z(n2656) );
  NAND U2325 ( .A(n2657), .B(n2658), .Z(n2655) );
  NANDN U2326 ( .A(B[360]), .B(A[360]), .Z(n2658) );
  AND U2327 ( .A(n2659), .B(n2660), .Z(n2657) );
  NAND U2328 ( .A(n2661), .B(n2662), .Z(n2660) );
  NANDN U2329 ( .A(A[359]), .B(B[359]), .Z(n2662) );
  AND U2330 ( .A(n2663), .B(n2664), .Z(n2661) );
  NANDN U2331 ( .A(A[358]), .B(B[358]), .Z(n2664) );
  NAND U2332 ( .A(n2665), .B(n2666), .Z(n2663) );
  NANDN U2333 ( .A(B[358]), .B(A[358]), .Z(n2666) );
  AND U2334 ( .A(n2667), .B(n2668), .Z(n2665) );
  NAND U2335 ( .A(n2669), .B(n2670), .Z(n2668) );
  NANDN U2336 ( .A(A[357]), .B(B[357]), .Z(n2670) );
  AND U2337 ( .A(n2671), .B(n2672), .Z(n2669) );
  NANDN U2338 ( .A(A[356]), .B(B[356]), .Z(n2672) );
  NAND U2339 ( .A(n2673), .B(n2674), .Z(n2671) );
  NANDN U2340 ( .A(B[356]), .B(A[356]), .Z(n2674) );
  AND U2341 ( .A(n2675), .B(n2676), .Z(n2673) );
  NAND U2342 ( .A(n2677), .B(n2678), .Z(n2676) );
  NANDN U2343 ( .A(A[355]), .B(B[355]), .Z(n2678) );
  AND U2344 ( .A(n2679), .B(n2680), .Z(n2677) );
  NANDN U2345 ( .A(A[354]), .B(B[354]), .Z(n2680) );
  NAND U2346 ( .A(n2681), .B(n2682), .Z(n2679) );
  NANDN U2347 ( .A(B[354]), .B(A[354]), .Z(n2682) );
  AND U2348 ( .A(n2683), .B(n2684), .Z(n2681) );
  NAND U2349 ( .A(n2685), .B(n2686), .Z(n2684) );
  NANDN U2350 ( .A(A[353]), .B(B[353]), .Z(n2686) );
  AND U2351 ( .A(n2687), .B(n2688), .Z(n2685) );
  NANDN U2352 ( .A(A[352]), .B(B[352]), .Z(n2688) );
  NAND U2353 ( .A(n2689), .B(n2690), .Z(n2687) );
  NANDN U2354 ( .A(B[352]), .B(A[352]), .Z(n2690) );
  AND U2355 ( .A(n2691), .B(n2692), .Z(n2689) );
  NAND U2356 ( .A(n2693), .B(n2694), .Z(n2692) );
  NANDN U2357 ( .A(A[351]), .B(B[351]), .Z(n2694) );
  AND U2358 ( .A(n2695), .B(n2696), .Z(n2693) );
  NANDN U2359 ( .A(A[350]), .B(B[350]), .Z(n2696) );
  NAND U2360 ( .A(n2697), .B(n2698), .Z(n2695) );
  NANDN U2361 ( .A(B[350]), .B(A[350]), .Z(n2698) );
  AND U2362 ( .A(n2699), .B(n2700), .Z(n2697) );
  NAND U2363 ( .A(n2701), .B(n2702), .Z(n2700) );
  NANDN U2364 ( .A(A[349]), .B(B[349]), .Z(n2702) );
  AND U2365 ( .A(n2703), .B(n2704), .Z(n2701) );
  NANDN U2366 ( .A(A[348]), .B(B[348]), .Z(n2704) );
  NAND U2367 ( .A(n2705), .B(n2706), .Z(n2703) );
  NANDN U2368 ( .A(B[348]), .B(A[348]), .Z(n2706) );
  AND U2369 ( .A(n2707), .B(n2708), .Z(n2705) );
  NAND U2370 ( .A(n2709), .B(n2710), .Z(n2708) );
  NANDN U2371 ( .A(A[347]), .B(B[347]), .Z(n2710) );
  AND U2372 ( .A(n2711), .B(n2712), .Z(n2709) );
  NANDN U2373 ( .A(A[346]), .B(B[346]), .Z(n2712) );
  NAND U2374 ( .A(n2713), .B(n2714), .Z(n2711) );
  NANDN U2375 ( .A(B[346]), .B(A[346]), .Z(n2714) );
  AND U2376 ( .A(n2715), .B(n2716), .Z(n2713) );
  NAND U2377 ( .A(n2717), .B(n2718), .Z(n2716) );
  NANDN U2378 ( .A(A[345]), .B(B[345]), .Z(n2718) );
  AND U2379 ( .A(n2719), .B(n2720), .Z(n2717) );
  NANDN U2380 ( .A(A[344]), .B(B[344]), .Z(n2720) );
  NAND U2381 ( .A(n2721), .B(n2722), .Z(n2719) );
  NANDN U2382 ( .A(B[344]), .B(A[344]), .Z(n2722) );
  AND U2383 ( .A(n2723), .B(n2724), .Z(n2721) );
  NAND U2384 ( .A(n2725), .B(n2726), .Z(n2724) );
  NANDN U2385 ( .A(A[343]), .B(B[343]), .Z(n2726) );
  AND U2386 ( .A(n2727), .B(n2728), .Z(n2725) );
  NANDN U2387 ( .A(A[342]), .B(B[342]), .Z(n2728) );
  NAND U2388 ( .A(n2729), .B(n2730), .Z(n2727) );
  NANDN U2389 ( .A(B[342]), .B(A[342]), .Z(n2730) );
  AND U2390 ( .A(n2731), .B(n2732), .Z(n2729) );
  NAND U2391 ( .A(n2733), .B(n2734), .Z(n2732) );
  NANDN U2392 ( .A(A[341]), .B(B[341]), .Z(n2734) );
  AND U2393 ( .A(n2735), .B(n2736), .Z(n2733) );
  NANDN U2394 ( .A(A[340]), .B(B[340]), .Z(n2736) );
  NAND U2395 ( .A(n2737), .B(n2738), .Z(n2735) );
  NANDN U2396 ( .A(B[340]), .B(A[340]), .Z(n2738) );
  AND U2397 ( .A(n2739), .B(n2740), .Z(n2737) );
  NAND U2398 ( .A(n2741), .B(n2742), .Z(n2740) );
  NANDN U2399 ( .A(A[339]), .B(B[339]), .Z(n2742) );
  AND U2400 ( .A(n2743), .B(n2744), .Z(n2741) );
  NANDN U2401 ( .A(A[338]), .B(B[338]), .Z(n2744) );
  NAND U2402 ( .A(n2745), .B(n2746), .Z(n2743) );
  NANDN U2403 ( .A(B[338]), .B(A[338]), .Z(n2746) );
  AND U2404 ( .A(n2747), .B(n2748), .Z(n2745) );
  NAND U2405 ( .A(n2749), .B(n2750), .Z(n2748) );
  NANDN U2406 ( .A(A[337]), .B(B[337]), .Z(n2750) );
  AND U2407 ( .A(n2751), .B(n2752), .Z(n2749) );
  NANDN U2408 ( .A(A[336]), .B(B[336]), .Z(n2752) );
  NAND U2409 ( .A(n2753), .B(n2754), .Z(n2751) );
  NANDN U2410 ( .A(B[336]), .B(A[336]), .Z(n2754) );
  AND U2411 ( .A(n2755), .B(n2756), .Z(n2753) );
  NAND U2412 ( .A(n2757), .B(n2758), .Z(n2756) );
  NANDN U2413 ( .A(A[335]), .B(B[335]), .Z(n2758) );
  AND U2414 ( .A(n2759), .B(n2760), .Z(n2757) );
  NANDN U2415 ( .A(A[334]), .B(B[334]), .Z(n2760) );
  NAND U2416 ( .A(n2761), .B(n2762), .Z(n2759) );
  NANDN U2417 ( .A(B[334]), .B(A[334]), .Z(n2762) );
  AND U2418 ( .A(n2763), .B(n2764), .Z(n2761) );
  NAND U2419 ( .A(n2765), .B(n2766), .Z(n2764) );
  NANDN U2420 ( .A(A[333]), .B(B[333]), .Z(n2766) );
  AND U2421 ( .A(n2767), .B(n2768), .Z(n2765) );
  NANDN U2422 ( .A(A[332]), .B(B[332]), .Z(n2768) );
  NAND U2423 ( .A(n2769), .B(n2770), .Z(n2767) );
  NANDN U2424 ( .A(B[332]), .B(A[332]), .Z(n2770) );
  AND U2425 ( .A(n2771), .B(n2772), .Z(n2769) );
  NAND U2426 ( .A(n2773), .B(n2774), .Z(n2772) );
  NANDN U2427 ( .A(A[331]), .B(B[331]), .Z(n2774) );
  AND U2428 ( .A(n2775), .B(n2776), .Z(n2773) );
  NANDN U2429 ( .A(A[330]), .B(B[330]), .Z(n2776) );
  NAND U2430 ( .A(n2777), .B(n2778), .Z(n2775) );
  NANDN U2431 ( .A(B[330]), .B(A[330]), .Z(n2778) );
  AND U2432 ( .A(n2779), .B(n2780), .Z(n2777) );
  NAND U2433 ( .A(n2781), .B(n2782), .Z(n2780) );
  NANDN U2434 ( .A(A[329]), .B(B[329]), .Z(n2782) );
  AND U2435 ( .A(n2783), .B(n2784), .Z(n2781) );
  NANDN U2436 ( .A(A[328]), .B(B[328]), .Z(n2784) );
  NAND U2437 ( .A(n2785), .B(n2786), .Z(n2783) );
  NANDN U2438 ( .A(B[328]), .B(A[328]), .Z(n2786) );
  AND U2439 ( .A(n2787), .B(n2788), .Z(n2785) );
  NAND U2440 ( .A(n2789), .B(n2790), .Z(n2788) );
  NANDN U2441 ( .A(A[327]), .B(B[327]), .Z(n2790) );
  AND U2442 ( .A(n2791), .B(n2792), .Z(n2789) );
  NANDN U2443 ( .A(A[326]), .B(B[326]), .Z(n2792) );
  NAND U2444 ( .A(n2793), .B(n2794), .Z(n2791) );
  NANDN U2445 ( .A(B[326]), .B(A[326]), .Z(n2794) );
  AND U2446 ( .A(n2795), .B(n2796), .Z(n2793) );
  NAND U2447 ( .A(n2797), .B(n2798), .Z(n2796) );
  NANDN U2448 ( .A(A[325]), .B(B[325]), .Z(n2798) );
  AND U2449 ( .A(n2799), .B(n2800), .Z(n2797) );
  NANDN U2450 ( .A(A[324]), .B(B[324]), .Z(n2800) );
  NAND U2451 ( .A(n2801), .B(n2802), .Z(n2799) );
  NANDN U2452 ( .A(B[324]), .B(A[324]), .Z(n2802) );
  AND U2453 ( .A(n2803), .B(n2804), .Z(n2801) );
  NAND U2454 ( .A(n2805), .B(n2806), .Z(n2804) );
  NANDN U2455 ( .A(A[323]), .B(B[323]), .Z(n2806) );
  AND U2456 ( .A(n2807), .B(n2808), .Z(n2805) );
  NANDN U2457 ( .A(A[322]), .B(B[322]), .Z(n2808) );
  NAND U2458 ( .A(n2809), .B(n2810), .Z(n2807) );
  NANDN U2459 ( .A(B[322]), .B(A[322]), .Z(n2810) );
  AND U2460 ( .A(n2811), .B(n2812), .Z(n2809) );
  NAND U2461 ( .A(n2813), .B(n2814), .Z(n2812) );
  NANDN U2462 ( .A(A[321]), .B(B[321]), .Z(n2814) );
  AND U2463 ( .A(n2815), .B(n2816), .Z(n2813) );
  NANDN U2464 ( .A(A[320]), .B(B[320]), .Z(n2816) );
  NAND U2465 ( .A(n2817), .B(n2818), .Z(n2815) );
  NANDN U2466 ( .A(B[320]), .B(A[320]), .Z(n2818) );
  AND U2467 ( .A(n2819), .B(n2820), .Z(n2817) );
  NAND U2468 ( .A(n2821), .B(n2822), .Z(n2820) );
  NANDN U2469 ( .A(A[319]), .B(B[319]), .Z(n2822) );
  AND U2470 ( .A(n2823), .B(n2824), .Z(n2821) );
  NANDN U2471 ( .A(A[318]), .B(B[318]), .Z(n2824) );
  NAND U2472 ( .A(n2825), .B(n2826), .Z(n2823) );
  NANDN U2473 ( .A(B[318]), .B(A[318]), .Z(n2826) );
  AND U2474 ( .A(n2827), .B(n2828), .Z(n2825) );
  NAND U2475 ( .A(n2829), .B(n2830), .Z(n2828) );
  NANDN U2476 ( .A(A[317]), .B(B[317]), .Z(n2830) );
  AND U2477 ( .A(n2831), .B(n2832), .Z(n2829) );
  NANDN U2478 ( .A(A[316]), .B(B[316]), .Z(n2832) );
  NAND U2479 ( .A(n2833), .B(n2834), .Z(n2831) );
  NANDN U2480 ( .A(B[316]), .B(A[316]), .Z(n2834) );
  AND U2481 ( .A(n2835), .B(n2836), .Z(n2833) );
  NAND U2482 ( .A(n2837), .B(n2838), .Z(n2836) );
  NANDN U2483 ( .A(A[315]), .B(B[315]), .Z(n2838) );
  AND U2484 ( .A(n2839), .B(n2840), .Z(n2837) );
  NANDN U2485 ( .A(A[314]), .B(B[314]), .Z(n2840) );
  NAND U2486 ( .A(n2841), .B(n2842), .Z(n2839) );
  NANDN U2487 ( .A(B[314]), .B(A[314]), .Z(n2842) );
  AND U2488 ( .A(n2843), .B(n2844), .Z(n2841) );
  NAND U2489 ( .A(n2845), .B(n2846), .Z(n2844) );
  NANDN U2490 ( .A(A[313]), .B(B[313]), .Z(n2846) );
  AND U2491 ( .A(n2847), .B(n2848), .Z(n2845) );
  NANDN U2492 ( .A(A[312]), .B(B[312]), .Z(n2848) );
  NAND U2493 ( .A(n2849), .B(n2850), .Z(n2847) );
  NANDN U2494 ( .A(B[312]), .B(A[312]), .Z(n2850) );
  AND U2495 ( .A(n2851), .B(n2852), .Z(n2849) );
  NAND U2496 ( .A(n2853), .B(n2854), .Z(n2852) );
  NANDN U2497 ( .A(A[311]), .B(B[311]), .Z(n2854) );
  AND U2498 ( .A(n2855), .B(n2856), .Z(n2853) );
  NANDN U2499 ( .A(A[310]), .B(B[310]), .Z(n2856) );
  NAND U2500 ( .A(n2857), .B(n2858), .Z(n2855) );
  NANDN U2501 ( .A(B[310]), .B(A[310]), .Z(n2858) );
  AND U2502 ( .A(n2859), .B(n2860), .Z(n2857) );
  NAND U2503 ( .A(n2861), .B(n2862), .Z(n2860) );
  NANDN U2504 ( .A(A[309]), .B(B[309]), .Z(n2862) );
  AND U2505 ( .A(n2863), .B(n2864), .Z(n2861) );
  NANDN U2506 ( .A(A[308]), .B(B[308]), .Z(n2864) );
  NAND U2507 ( .A(n2865), .B(n2866), .Z(n2863) );
  NANDN U2508 ( .A(B[308]), .B(A[308]), .Z(n2866) );
  AND U2509 ( .A(n2867), .B(n2868), .Z(n2865) );
  NAND U2510 ( .A(n2869), .B(n2870), .Z(n2868) );
  NANDN U2511 ( .A(A[307]), .B(B[307]), .Z(n2870) );
  AND U2512 ( .A(n2871), .B(n2872), .Z(n2869) );
  NANDN U2513 ( .A(A[306]), .B(B[306]), .Z(n2872) );
  NAND U2514 ( .A(n2873), .B(n2874), .Z(n2871) );
  NANDN U2515 ( .A(B[306]), .B(A[306]), .Z(n2874) );
  AND U2516 ( .A(n2875), .B(n2876), .Z(n2873) );
  NAND U2517 ( .A(n2877), .B(n2878), .Z(n2876) );
  NANDN U2518 ( .A(A[305]), .B(B[305]), .Z(n2878) );
  AND U2519 ( .A(n2879), .B(n2880), .Z(n2877) );
  NANDN U2520 ( .A(A[304]), .B(B[304]), .Z(n2880) );
  NAND U2521 ( .A(n2881), .B(n2882), .Z(n2879) );
  NANDN U2522 ( .A(B[304]), .B(A[304]), .Z(n2882) );
  AND U2523 ( .A(n2883), .B(n2884), .Z(n2881) );
  NAND U2524 ( .A(n2885), .B(n2886), .Z(n2884) );
  NANDN U2525 ( .A(A[303]), .B(B[303]), .Z(n2886) );
  AND U2526 ( .A(n2887), .B(n2888), .Z(n2885) );
  NANDN U2527 ( .A(A[302]), .B(B[302]), .Z(n2888) );
  NAND U2528 ( .A(n2889), .B(n2890), .Z(n2887) );
  NANDN U2529 ( .A(B[302]), .B(A[302]), .Z(n2890) );
  AND U2530 ( .A(n2891), .B(n2892), .Z(n2889) );
  NAND U2531 ( .A(n2893), .B(n2894), .Z(n2892) );
  NANDN U2532 ( .A(A[301]), .B(B[301]), .Z(n2894) );
  AND U2533 ( .A(n2895), .B(n2896), .Z(n2893) );
  NANDN U2534 ( .A(A[300]), .B(B[300]), .Z(n2896) );
  NAND U2535 ( .A(n2897), .B(n2898), .Z(n2895) );
  NANDN U2536 ( .A(B[300]), .B(A[300]), .Z(n2898) );
  AND U2537 ( .A(n2899), .B(n2900), .Z(n2897) );
  NAND U2538 ( .A(n2901), .B(n2902), .Z(n2900) );
  NANDN U2539 ( .A(A[299]), .B(B[299]), .Z(n2902) );
  AND U2540 ( .A(n2903), .B(n2904), .Z(n2901) );
  NANDN U2541 ( .A(A[298]), .B(B[298]), .Z(n2904) );
  NAND U2542 ( .A(n2905), .B(n2906), .Z(n2903) );
  NANDN U2543 ( .A(B[298]), .B(A[298]), .Z(n2906) );
  AND U2544 ( .A(n2907), .B(n2908), .Z(n2905) );
  NAND U2545 ( .A(n2909), .B(n2910), .Z(n2908) );
  NANDN U2546 ( .A(A[297]), .B(B[297]), .Z(n2910) );
  AND U2547 ( .A(n2911), .B(n2912), .Z(n2909) );
  NANDN U2548 ( .A(A[296]), .B(B[296]), .Z(n2912) );
  NAND U2549 ( .A(n2913), .B(n2914), .Z(n2911) );
  NANDN U2550 ( .A(B[296]), .B(A[296]), .Z(n2914) );
  AND U2551 ( .A(n2915), .B(n2916), .Z(n2913) );
  NAND U2552 ( .A(n2917), .B(n2918), .Z(n2916) );
  NANDN U2553 ( .A(A[295]), .B(B[295]), .Z(n2918) );
  AND U2554 ( .A(n2919), .B(n2920), .Z(n2917) );
  NANDN U2555 ( .A(A[294]), .B(B[294]), .Z(n2920) );
  NAND U2556 ( .A(n2921), .B(n2922), .Z(n2919) );
  NANDN U2557 ( .A(B[294]), .B(A[294]), .Z(n2922) );
  AND U2558 ( .A(n2923), .B(n2924), .Z(n2921) );
  NAND U2559 ( .A(n2925), .B(n2926), .Z(n2924) );
  NANDN U2560 ( .A(A[293]), .B(B[293]), .Z(n2926) );
  AND U2561 ( .A(n2927), .B(n2928), .Z(n2925) );
  NANDN U2562 ( .A(A[292]), .B(B[292]), .Z(n2928) );
  NAND U2563 ( .A(n2929), .B(n2930), .Z(n2927) );
  NANDN U2564 ( .A(B[292]), .B(A[292]), .Z(n2930) );
  AND U2565 ( .A(n2931), .B(n2932), .Z(n2929) );
  NAND U2566 ( .A(n2933), .B(n2934), .Z(n2932) );
  NANDN U2567 ( .A(A[291]), .B(B[291]), .Z(n2934) );
  AND U2568 ( .A(n2935), .B(n2936), .Z(n2933) );
  NANDN U2569 ( .A(A[290]), .B(B[290]), .Z(n2936) );
  NAND U2570 ( .A(n2937), .B(n2938), .Z(n2935) );
  NANDN U2571 ( .A(B[290]), .B(A[290]), .Z(n2938) );
  AND U2572 ( .A(n2939), .B(n2940), .Z(n2937) );
  NAND U2573 ( .A(n2941), .B(n2942), .Z(n2940) );
  NANDN U2574 ( .A(A[289]), .B(B[289]), .Z(n2942) );
  AND U2575 ( .A(n2943), .B(n2944), .Z(n2941) );
  NANDN U2576 ( .A(A[288]), .B(B[288]), .Z(n2944) );
  NAND U2577 ( .A(n2945), .B(n2946), .Z(n2943) );
  NANDN U2578 ( .A(B[288]), .B(A[288]), .Z(n2946) );
  AND U2579 ( .A(n2947), .B(n2948), .Z(n2945) );
  NAND U2580 ( .A(n2949), .B(n2950), .Z(n2948) );
  NANDN U2581 ( .A(A[287]), .B(B[287]), .Z(n2950) );
  AND U2582 ( .A(n2951), .B(n2952), .Z(n2949) );
  NANDN U2583 ( .A(A[286]), .B(B[286]), .Z(n2952) );
  NAND U2584 ( .A(n2953), .B(n2954), .Z(n2951) );
  NANDN U2585 ( .A(B[286]), .B(A[286]), .Z(n2954) );
  AND U2586 ( .A(n2955), .B(n2956), .Z(n2953) );
  NAND U2587 ( .A(n2957), .B(n2958), .Z(n2956) );
  NANDN U2588 ( .A(A[285]), .B(B[285]), .Z(n2958) );
  AND U2589 ( .A(n2959), .B(n2960), .Z(n2957) );
  NANDN U2590 ( .A(A[284]), .B(B[284]), .Z(n2960) );
  NAND U2591 ( .A(n2961), .B(n2962), .Z(n2959) );
  NANDN U2592 ( .A(B[284]), .B(A[284]), .Z(n2962) );
  AND U2593 ( .A(n2963), .B(n2964), .Z(n2961) );
  NAND U2594 ( .A(n2965), .B(n2966), .Z(n2964) );
  NANDN U2595 ( .A(A[283]), .B(B[283]), .Z(n2966) );
  AND U2596 ( .A(n2967), .B(n2968), .Z(n2965) );
  NANDN U2597 ( .A(A[282]), .B(B[282]), .Z(n2968) );
  NAND U2598 ( .A(n2969), .B(n2970), .Z(n2967) );
  NANDN U2599 ( .A(B[282]), .B(A[282]), .Z(n2970) );
  AND U2600 ( .A(n2971), .B(n2972), .Z(n2969) );
  NAND U2601 ( .A(n2973), .B(n2974), .Z(n2972) );
  NANDN U2602 ( .A(A[281]), .B(B[281]), .Z(n2974) );
  AND U2603 ( .A(n2975), .B(n2976), .Z(n2973) );
  NANDN U2604 ( .A(A[280]), .B(B[280]), .Z(n2976) );
  NAND U2605 ( .A(n2977), .B(n2978), .Z(n2975) );
  NANDN U2606 ( .A(B[280]), .B(A[280]), .Z(n2978) );
  AND U2607 ( .A(n2979), .B(n2980), .Z(n2977) );
  NAND U2608 ( .A(n2981), .B(n2982), .Z(n2980) );
  NANDN U2609 ( .A(A[279]), .B(B[279]), .Z(n2982) );
  AND U2610 ( .A(n2983), .B(n2984), .Z(n2981) );
  NANDN U2611 ( .A(A[278]), .B(B[278]), .Z(n2984) );
  NAND U2612 ( .A(n2985), .B(n2986), .Z(n2983) );
  NANDN U2613 ( .A(B[278]), .B(A[278]), .Z(n2986) );
  AND U2614 ( .A(n2987), .B(n2988), .Z(n2985) );
  NAND U2615 ( .A(n2989), .B(n2990), .Z(n2988) );
  NANDN U2616 ( .A(A[277]), .B(B[277]), .Z(n2990) );
  AND U2617 ( .A(n2991), .B(n2992), .Z(n2989) );
  NANDN U2618 ( .A(A[276]), .B(B[276]), .Z(n2992) );
  NAND U2619 ( .A(n2993), .B(n2994), .Z(n2991) );
  NANDN U2620 ( .A(B[276]), .B(A[276]), .Z(n2994) );
  AND U2621 ( .A(n2995), .B(n2996), .Z(n2993) );
  NAND U2622 ( .A(n2997), .B(n2998), .Z(n2996) );
  NANDN U2623 ( .A(A[275]), .B(B[275]), .Z(n2998) );
  AND U2624 ( .A(n2999), .B(n3000), .Z(n2997) );
  NANDN U2625 ( .A(A[274]), .B(B[274]), .Z(n3000) );
  NAND U2626 ( .A(n3001), .B(n3002), .Z(n2999) );
  NANDN U2627 ( .A(B[274]), .B(A[274]), .Z(n3002) );
  AND U2628 ( .A(n3003), .B(n3004), .Z(n3001) );
  NAND U2629 ( .A(n3005), .B(n3006), .Z(n3004) );
  NANDN U2630 ( .A(A[273]), .B(B[273]), .Z(n3006) );
  AND U2631 ( .A(n3007), .B(n3008), .Z(n3005) );
  NANDN U2632 ( .A(A[272]), .B(B[272]), .Z(n3008) );
  NAND U2633 ( .A(n3009), .B(n3010), .Z(n3007) );
  NANDN U2634 ( .A(B[272]), .B(A[272]), .Z(n3010) );
  AND U2635 ( .A(n3011), .B(n3012), .Z(n3009) );
  NAND U2636 ( .A(n3013), .B(n3014), .Z(n3012) );
  NANDN U2637 ( .A(A[271]), .B(B[271]), .Z(n3014) );
  AND U2638 ( .A(n3015), .B(n3016), .Z(n3013) );
  NANDN U2639 ( .A(A[270]), .B(B[270]), .Z(n3016) );
  NAND U2640 ( .A(n3017), .B(n3018), .Z(n3015) );
  NANDN U2641 ( .A(B[270]), .B(A[270]), .Z(n3018) );
  AND U2642 ( .A(n3019), .B(n3020), .Z(n3017) );
  NAND U2643 ( .A(n3021), .B(n3022), .Z(n3020) );
  NANDN U2644 ( .A(A[269]), .B(B[269]), .Z(n3022) );
  AND U2645 ( .A(n3023), .B(n3024), .Z(n3021) );
  NANDN U2646 ( .A(A[268]), .B(B[268]), .Z(n3024) );
  NAND U2647 ( .A(n3025), .B(n3026), .Z(n3023) );
  NANDN U2648 ( .A(B[268]), .B(A[268]), .Z(n3026) );
  AND U2649 ( .A(n3027), .B(n3028), .Z(n3025) );
  NAND U2650 ( .A(n3029), .B(n3030), .Z(n3028) );
  NANDN U2651 ( .A(A[267]), .B(B[267]), .Z(n3030) );
  AND U2652 ( .A(n3031), .B(n3032), .Z(n3029) );
  NANDN U2653 ( .A(A[266]), .B(B[266]), .Z(n3032) );
  NAND U2654 ( .A(n3033), .B(n3034), .Z(n3031) );
  NANDN U2655 ( .A(B[266]), .B(A[266]), .Z(n3034) );
  AND U2656 ( .A(n3035), .B(n3036), .Z(n3033) );
  NAND U2657 ( .A(n3037), .B(n3038), .Z(n3036) );
  NANDN U2658 ( .A(A[265]), .B(B[265]), .Z(n3038) );
  AND U2659 ( .A(n3039), .B(n3040), .Z(n3037) );
  NANDN U2660 ( .A(A[264]), .B(B[264]), .Z(n3040) );
  NAND U2661 ( .A(n3041), .B(n3042), .Z(n3039) );
  NANDN U2662 ( .A(B[264]), .B(A[264]), .Z(n3042) );
  AND U2663 ( .A(n3043), .B(n3044), .Z(n3041) );
  NAND U2664 ( .A(n3045), .B(n3046), .Z(n3044) );
  NANDN U2665 ( .A(A[263]), .B(B[263]), .Z(n3046) );
  AND U2666 ( .A(n3047), .B(n3048), .Z(n3045) );
  NANDN U2667 ( .A(A[262]), .B(B[262]), .Z(n3048) );
  NAND U2668 ( .A(n3049), .B(n3050), .Z(n3047) );
  NANDN U2669 ( .A(B[262]), .B(A[262]), .Z(n3050) );
  AND U2670 ( .A(n3051), .B(n3052), .Z(n3049) );
  NAND U2671 ( .A(n3053), .B(n3054), .Z(n3052) );
  NANDN U2672 ( .A(A[261]), .B(B[261]), .Z(n3054) );
  AND U2673 ( .A(n3055), .B(n3056), .Z(n3053) );
  NANDN U2674 ( .A(A[260]), .B(B[260]), .Z(n3056) );
  NAND U2675 ( .A(n3057), .B(n3058), .Z(n3055) );
  NANDN U2676 ( .A(B[260]), .B(A[260]), .Z(n3058) );
  AND U2677 ( .A(n3059), .B(n3060), .Z(n3057) );
  NAND U2678 ( .A(n3061), .B(n3062), .Z(n3060) );
  NANDN U2679 ( .A(A[259]), .B(B[259]), .Z(n3062) );
  AND U2680 ( .A(n3063), .B(n3064), .Z(n3061) );
  NANDN U2681 ( .A(A[258]), .B(B[258]), .Z(n3064) );
  NAND U2682 ( .A(n3065), .B(n3066), .Z(n3063) );
  NANDN U2683 ( .A(B[258]), .B(A[258]), .Z(n3066) );
  AND U2684 ( .A(n3067), .B(n3068), .Z(n3065) );
  NAND U2685 ( .A(n3069), .B(n3070), .Z(n3068) );
  NANDN U2686 ( .A(A[257]), .B(B[257]), .Z(n3070) );
  AND U2687 ( .A(n3071), .B(n3072), .Z(n3069) );
  NANDN U2688 ( .A(A[256]), .B(B[256]), .Z(n3072) );
  NAND U2689 ( .A(n3073), .B(n3074), .Z(n3071) );
  NANDN U2690 ( .A(B[256]), .B(A[256]), .Z(n3074) );
  AND U2691 ( .A(n3075), .B(n3076), .Z(n3073) );
  NAND U2692 ( .A(n3077), .B(n3078), .Z(n3076) );
  NANDN U2693 ( .A(A[255]), .B(B[255]), .Z(n3078) );
  AND U2694 ( .A(n3079), .B(n3080), .Z(n3077) );
  NANDN U2695 ( .A(A[254]), .B(B[254]), .Z(n3080) );
  NAND U2696 ( .A(n3081), .B(n3082), .Z(n3079) );
  NANDN U2697 ( .A(B[254]), .B(A[254]), .Z(n3082) );
  AND U2698 ( .A(n3083), .B(n3084), .Z(n3081) );
  NAND U2699 ( .A(n3085), .B(n3086), .Z(n3084) );
  NANDN U2700 ( .A(A[253]), .B(B[253]), .Z(n3086) );
  AND U2701 ( .A(n3087), .B(n3088), .Z(n3085) );
  NANDN U2702 ( .A(A[252]), .B(B[252]), .Z(n3088) );
  NAND U2703 ( .A(n3089), .B(n3090), .Z(n3087) );
  NANDN U2704 ( .A(B[252]), .B(A[252]), .Z(n3090) );
  AND U2705 ( .A(n3091), .B(n3092), .Z(n3089) );
  NAND U2706 ( .A(n3093), .B(n3094), .Z(n3092) );
  NANDN U2707 ( .A(A[251]), .B(B[251]), .Z(n3094) );
  AND U2708 ( .A(n3095), .B(n3096), .Z(n3093) );
  NANDN U2709 ( .A(A[250]), .B(B[250]), .Z(n3096) );
  NAND U2710 ( .A(n3097), .B(n3098), .Z(n3095) );
  NANDN U2711 ( .A(B[250]), .B(A[250]), .Z(n3098) );
  AND U2712 ( .A(n3099), .B(n3100), .Z(n3097) );
  NAND U2713 ( .A(n3101), .B(n3102), .Z(n3100) );
  NANDN U2714 ( .A(A[249]), .B(B[249]), .Z(n3102) );
  AND U2715 ( .A(n3103), .B(n3104), .Z(n3101) );
  NANDN U2716 ( .A(A[248]), .B(B[248]), .Z(n3104) );
  NAND U2717 ( .A(n3105), .B(n3106), .Z(n3103) );
  NANDN U2718 ( .A(B[248]), .B(A[248]), .Z(n3106) );
  AND U2719 ( .A(n3107), .B(n3108), .Z(n3105) );
  NAND U2720 ( .A(n3109), .B(n3110), .Z(n3108) );
  NANDN U2721 ( .A(A[247]), .B(B[247]), .Z(n3110) );
  AND U2722 ( .A(n3111), .B(n3112), .Z(n3109) );
  NANDN U2723 ( .A(A[246]), .B(B[246]), .Z(n3112) );
  NAND U2724 ( .A(n3113), .B(n3114), .Z(n3111) );
  NANDN U2725 ( .A(B[246]), .B(A[246]), .Z(n3114) );
  AND U2726 ( .A(n3115), .B(n3116), .Z(n3113) );
  NAND U2727 ( .A(n3117), .B(n3118), .Z(n3116) );
  NANDN U2728 ( .A(A[245]), .B(B[245]), .Z(n3118) );
  AND U2729 ( .A(n3119), .B(n3120), .Z(n3117) );
  NANDN U2730 ( .A(A[244]), .B(B[244]), .Z(n3120) );
  NAND U2731 ( .A(n3121), .B(n3122), .Z(n3119) );
  NANDN U2732 ( .A(B[244]), .B(A[244]), .Z(n3122) );
  AND U2733 ( .A(n3123), .B(n3124), .Z(n3121) );
  NAND U2734 ( .A(n3125), .B(n3126), .Z(n3124) );
  NANDN U2735 ( .A(A[243]), .B(B[243]), .Z(n3126) );
  AND U2736 ( .A(n3127), .B(n3128), .Z(n3125) );
  NANDN U2737 ( .A(A[242]), .B(B[242]), .Z(n3128) );
  NAND U2738 ( .A(n3129), .B(n3130), .Z(n3127) );
  NANDN U2739 ( .A(B[242]), .B(A[242]), .Z(n3130) );
  AND U2740 ( .A(n3131), .B(n3132), .Z(n3129) );
  NAND U2741 ( .A(n3133), .B(n3134), .Z(n3132) );
  NANDN U2742 ( .A(A[241]), .B(B[241]), .Z(n3134) );
  AND U2743 ( .A(n3135), .B(n3136), .Z(n3133) );
  NANDN U2744 ( .A(A[240]), .B(B[240]), .Z(n3136) );
  NAND U2745 ( .A(n3137), .B(n3138), .Z(n3135) );
  NANDN U2746 ( .A(B[240]), .B(A[240]), .Z(n3138) );
  AND U2747 ( .A(n3139), .B(n3140), .Z(n3137) );
  NAND U2748 ( .A(n3141), .B(n3142), .Z(n3140) );
  NANDN U2749 ( .A(A[239]), .B(B[239]), .Z(n3142) );
  AND U2750 ( .A(n3143), .B(n3144), .Z(n3141) );
  NANDN U2751 ( .A(A[238]), .B(B[238]), .Z(n3144) );
  NAND U2752 ( .A(n3145), .B(n3146), .Z(n3143) );
  NANDN U2753 ( .A(B[238]), .B(A[238]), .Z(n3146) );
  AND U2754 ( .A(n3147), .B(n3148), .Z(n3145) );
  NAND U2755 ( .A(n3149), .B(n3150), .Z(n3148) );
  NANDN U2756 ( .A(A[237]), .B(B[237]), .Z(n3150) );
  AND U2757 ( .A(n3151), .B(n3152), .Z(n3149) );
  NANDN U2758 ( .A(A[236]), .B(B[236]), .Z(n3152) );
  NAND U2759 ( .A(n3153), .B(n3154), .Z(n3151) );
  NANDN U2760 ( .A(B[236]), .B(A[236]), .Z(n3154) );
  AND U2761 ( .A(n3155), .B(n3156), .Z(n3153) );
  NAND U2762 ( .A(n3157), .B(n3158), .Z(n3156) );
  NANDN U2763 ( .A(A[235]), .B(B[235]), .Z(n3158) );
  AND U2764 ( .A(n3159), .B(n3160), .Z(n3157) );
  NANDN U2765 ( .A(A[234]), .B(B[234]), .Z(n3160) );
  NAND U2766 ( .A(n3161), .B(n3162), .Z(n3159) );
  NANDN U2767 ( .A(B[234]), .B(A[234]), .Z(n3162) );
  AND U2768 ( .A(n3163), .B(n3164), .Z(n3161) );
  NAND U2769 ( .A(n3165), .B(n3166), .Z(n3164) );
  NANDN U2770 ( .A(A[233]), .B(B[233]), .Z(n3166) );
  AND U2771 ( .A(n3167), .B(n3168), .Z(n3165) );
  NANDN U2772 ( .A(A[232]), .B(B[232]), .Z(n3168) );
  NAND U2773 ( .A(n3169), .B(n3170), .Z(n3167) );
  NANDN U2774 ( .A(B[232]), .B(A[232]), .Z(n3170) );
  AND U2775 ( .A(n3171), .B(n3172), .Z(n3169) );
  NAND U2776 ( .A(n3173), .B(n3174), .Z(n3172) );
  NANDN U2777 ( .A(A[231]), .B(B[231]), .Z(n3174) );
  AND U2778 ( .A(n3175), .B(n3176), .Z(n3173) );
  NANDN U2779 ( .A(A[230]), .B(B[230]), .Z(n3176) );
  NAND U2780 ( .A(n3177), .B(n3178), .Z(n3175) );
  NANDN U2781 ( .A(B[230]), .B(A[230]), .Z(n3178) );
  AND U2782 ( .A(n3179), .B(n3180), .Z(n3177) );
  NAND U2783 ( .A(n3181), .B(n3182), .Z(n3180) );
  NANDN U2784 ( .A(A[229]), .B(B[229]), .Z(n3182) );
  AND U2785 ( .A(n3183), .B(n3184), .Z(n3181) );
  NANDN U2786 ( .A(A[228]), .B(B[228]), .Z(n3184) );
  NAND U2787 ( .A(n3185), .B(n3186), .Z(n3183) );
  NANDN U2788 ( .A(B[228]), .B(A[228]), .Z(n3186) );
  AND U2789 ( .A(n3187), .B(n3188), .Z(n3185) );
  NAND U2790 ( .A(n3189), .B(n3190), .Z(n3188) );
  NANDN U2791 ( .A(A[227]), .B(B[227]), .Z(n3190) );
  AND U2792 ( .A(n3191), .B(n3192), .Z(n3189) );
  NANDN U2793 ( .A(A[226]), .B(B[226]), .Z(n3192) );
  NAND U2794 ( .A(n3193), .B(n3194), .Z(n3191) );
  NANDN U2795 ( .A(B[226]), .B(A[226]), .Z(n3194) );
  AND U2796 ( .A(n3195), .B(n3196), .Z(n3193) );
  NAND U2797 ( .A(n3197), .B(n3198), .Z(n3196) );
  NANDN U2798 ( .A(A[225]), .B(B[225]), .Z(n3198) );
  AND U2799 ( .A(n3199), .B(n3200), .Z(n3197) );
  NANDN U2800 ( .A(A[224]), .B(B[224]), .Z(n3200) );
  NAND U2801 ( .A(n3201), .B(n3202), .Z(n3199) );
  NANDN U2802 ( .A(B[224]), .B(A[224]), .Z(n3202) );
  AND U2803 ( .A(n3203), .B(n3204), .Z(n3201) );
  NAND U2804 ( .A(n3205), .B(n3206), .Z(n3204) );
  NANDN U2805 ( .A(A[223]), .B(B[223]), .Z(n3206) );
  AND U2806 ( .A(n3207), .B(n3208), .Z(n3205) );
  NANDN U2807 ( .A(A[222]), .B(B[222]), .Z(n3208) );
  NAND U2808 ( .A(n3209), .B(n3210), .Z(n3207) );
  NANDN U2809 ( .A(B[222]), .B(A[222]), .Z(n3210) );
  AND U2810 ( .A(n3211), .B(n3212), .Z(n3209) );
  NAND U2811 ( .A(n3213), .B(n3214), .Z(n3212) );
  NANDN U2812 ( .A(A[221]), .B(B[221]), .Z(n3214) );
  AND U2813 ( .A(n3215), .B(n3216), .Z(n3213) );
  NANDN U2814 ( .A(A[220]), .B(B[220]), .Z(n3216) );
  NAND U2815 ( .A(n3217), .B(n3218), .Z(n3215) );
  NANDN U2816 ( .A(B[220]), .B(A[220]), .Z(n3218) );
  AND U2817 ( .A(n3219), .B(n3220), .Z(n3217) );
  NAND U2818 ( .A(n3221), .B(n3222), .Z(n3220) );
  NANDN U2819 ( .A(A[219]), .B(B[219]), .Z(n3222) );
  AND U2820 ( .A(n3223), .B(n3224), .Z(n3221) );
  NANDN U2821 ( .A(A[218]), .B(B[218]), .Z(n3224) );
  NAND U2822 ( .A(n3225), .B(n3226), .Z(n3223) );
  NANDN U2823 ( .A(B[218]), .B(A[218]), .Z(n3226) );
  AND U2824 ( .A(n3227), .B(n3228), .Z(n3225) );
  NAND U2825 ( .A(n3229), .B(n3230), .Z(n3228) );
  NANDN U2826 ( .A(A[217]), .B(B[217]), .Z(n3230) );
  AND U2827 ( .A(n3231), .B(n3232), .Z(n3229) );
  NANDN U2828 ( .A(A[216]), .B(B[216]), .Z(n3232) );
  NAND U2829 ( .A(n3233), .B(n3234), .Z(n3231) );
  NANDN U2830 ( .A(B[216]), .B(A[216]), .Z(n3234) );
  AND U2831 ( .A(n3235), .B(n3236), .Z(n3233) );
  NAND U2832 ( .A(n3237), .B(n3238), .Z(n3236) );
  NANDN U2833 ( .A(A[215]), .B(B[215]), .Z(n3238) );
  AND U2834 ( .A(n3239), .B(n3240), .Z(n3237) );
  NANDN U2835 ( .A(A[214]), .B(B[214]), .Z(n3240) );
  NAND U2836 ( .A(n3241), .B(n3242), .Z(n3239) );
  NANDN U2837 ( .A(B[214]), .B(A[214]), .Z(n3242) );
  AND U2838 ( .A(n3243), .B(n3244), .Z(n3241) );
  NAND U2839 ( .A(n3245), .B(n3246), .Z(n3244) );
  NANDN U2840 ( .A(A[213]), .B(B[213]), .Z(n3246) );
  AND U2841 ( .A(n3247), .B(n3248), .Z(n3245) );
  NANDN U2842 ( .A(A[212]), .B(B[212]), .Z(n3248) );
  NAND U2843 ( .A(n3249), .B(n3250), .Z(n3247) );
  NANDN U2844 ( .A(B[212]), .B(A[212]), .Z(n3250) );
  AND U2845 ( .A(n3251), .B(n3252), .Z(n3249) );
  NAND U2846 ( .A(n3253), .B(n3254), .Z(n3252) );
  NANDN U2847 ( .A(A[211]), .B(B[211]), .Z(n3254) );
  AND U2848 ( .A(n3255), .B(n3256), .Z(n3253) );
  NANDN U2849 ( .A(A[210]), .B(B[210]), .Z(n3256) );
  NAND U2850 ( .A(n3257), .B(n3258), .Z(n3255) );
  NANDN U2851 ( .A(B[210]), .B(A[210]), .Z(n3258) );
  AND U2852 ( .A(n3259), .B(n3260), .Z(n3257) );
  NAND U2853 ( .A(n3261), .B(n3262), .Z(n3260) );
  NANDN U2854 ( .A(A[209]), .B(B[209]), .Z(n3262) );
  AND U2855 ( .A(n3263), .B(n3264), .Z(n3261) );
  NANDN U2856 ( .A(A[208]), .B(B[208]), .Z(n3264) );
  NAND U2857 ( .A(n3265), .B(n3266), .Z(n3263) );
  NANDN U2858 ( .A(B[208]), .B(A[208]), .Z(n3266) );
  AND U2859 ( .A(n3267), .B(n3268), .Z(n3265) );
  NAND U2860 ( .A(n3269), .B(n3270), .Z(n3268) );
  NANDN U2861 ( .A(A[207]), .B(B[207]), .Z(n3270) );
  AND U2862 ( .A(n3271), .B(n3272), .Z(n3269) );
  NANDN U2863 ( .A(A[206]), .B(B[206]), .Z(n3272) );
  NAND U2864 ( .A(n3273), .B(n3274), .Z(n3271) );
  NANDN U2865 ( .A(B[206]), .B(A[206]), .Z(n3274) );
  AND U2866 ( .A(n3275), .B(n3276), .Z(n3273) );
  NAND U2867 ( .A(n3277), .B(n3278), .Z(n3276) );
  NANDN U2868 ( .A(A[205]), .B(B[205]), .Z(n3278) );
  AND U2869 ( .A(n3279), .B(n3280), .Z(n3277) );
  NANDN U2870 ( .A(A[204]), .B(B[204]), .Z(n3280) );
  NAND U2871 ( .A(n3281), .B(n3282), .Z(n3279) );
  NANDN U2872 ( .A(B[204]), .B(A[204]), .Z(n3282) );
  AND U2873 ( .A(n3283), .B(n3284), .Z(n3281) );
  NAND U2874 ( .A(n3285), .B(n3286), .Z(n3284) );
  NANDN U2875 ( .A(A[203]), .B(B[203]), .Z(n3286) );
  AND U2876 ( .A(n3287), .B(n3288), .Z(n3285) );
  NANDN U2877 ( .A(A[202]), .B(B[202]), .Z(n3288) );
  NAND U2878 ( .A(n3289), .B(n3290), .Z(n3287) );
  NANDN U2879 ( .A(B[202]), .B(A[202]), .Z(n3290) );
  AND U2880 ( .A(n3291), .B(n3292), .Z(n3289) );
  NAND U2881 ( .A(n3293), .B(n3294), .Z(n3292) );
  NANDN U2882 ( .A(A[201]), .B(B[201]), .Z(n3294) );
  AND U2883 ( .A(n3295), .B(n3296), .Z(n3293) );
  NANDN U2884 ( .A(A[200]), .B(B[200]), .Z(n3296) );
  NAND U2885 ( .A(n3297), .B(n3298), .Z(n3295) );
  NANDN U2886 ( .A(B[200]), .B(A[200]), .Z(n3298) );
  AND U2887 ( .A(n3299), .B(n3300), .Z(n3297) );
  NAND U2888 ( .A(n3301), .B(n3302), .Z(n3300) );
  NANDN U2889 ( .A(A[199]), .B(B[199]), .Z(n3302) );
  AND U2890 ( .A(n3303), .B(n3304), .Z(n3301) );
  NANDN U2891 ( .A(A[198]), .B(B[198]), .Z(n3304) );
  NAND U2892 ( .A(n3305), .B(n3306), .Z(n3303) );
  NANDN U2893 ( .A(B[198]), .B(A[198]), .Z(n3306) );
  AND U2894 ( .A(n3307), .B(n3308), .Z(n3305) );
  NAND U2895 ( .A(n3309), .B(n3310), .Z(n3308) );
  NANDN U2896 ( .A(A[197]), .B(B[197]), .Z(n3310) );
  AND U2897 ( .A(n3311), .B(n3312), .Z(n3309) );
  NANDN U2898 ( .A(A[196]), .B(B[196]), .Z(n3312) );
  NAND U2899 ( .A(n3313), .B(n3314), .Z(n3311) );
  NANDN U2900 ( .A(B[196]), .B(A[196]), .Z(n3314) );
  AND U2901 ( .A(n3315), .B(n3316), .Z(n3313) );
  NAND U2902 ( .A(n3317), .B(n3318), .Z(n3316) );
  NANDN U2903 ( .A(A[195]), .B(B[195]), .Z(n3318) );
  AND U2904 ( .A(n3319), .B(n3320), .Z(n3317) );
  NANDN U2905 ( .A(A[194]), .B(B[194]), .Z(n3320) );
  NAND U2906 ( .A(n3321), .B(n3322), .Z(n3319) );
  NANDN U2907 ( .A(B[194]), .B(A[194]), .Z(n3322) );
  AND U2908 ( .A(n3323), .B(n3324), .Z(n3321) );
  NAND U2909 ( .A(n3325), .B(n3326), .Z(n3324) );
  NANDN U2910 ( .A(A[193]), .B(B[193]), .Z(n3326) );
  AND U2911 ( .A(n3327), .B(n3328), .Z(n3325) );
  NANDN U2912 ( .A(A[192]), .B(B[192]), .Z(n3328) );
  NAND U2913 ( .A(n3329), .B(n3330), .Z(n3327) );
  NANDN U2914 ( .A(B[192]), .B(A[192]), .Z(n3330) );
  AND U2915 ( .A(n3331), .B(n3332), .Z(n3329) );
  NAND U2916 ( .A(n3333), .B(n3334), .Z(n3332) );
  NANDN U2917 ( .A(A[191]), .B(B[191]), .Z(n3334) );
  AND U2918 ( .A(n3335), .B(n3336), .Z(n3333) );
  NANDN U2919 ( .A(A[190]), .B(B[190]), .Z(n3336) );
  NAND U2920 ( .A(n3337), .B(n3338), .Z(n3335) );
  NANDN U2921 ( .A(B[190]), .B(A[190]), .Z(n3338) );
  AND U2922 ( .A(n3339), .B(n3340), .Z(n3337) );
  NAND U2923 ( .A(n3341), .B(n3342), .Z(n3340) );
  NANDN U2924 ( .A(A[189]), .B(B[189]), .Z(n3342) );
  AND U2925 ( .A(n3343), .B(n3344), .Z(n3341) );
  NANDN U2926 ( .A(A[188]), .B(B[188]), .Z(n3344) );
  NAND U2927 ( .A(n3345), .B(n3346), .Z(n3343) );
  NANDN U2928 ( .A(B[188]), .B(A[188]), .Z(n3346) );
  AND U2929 ( .A(n3347), .B(n3348), .Z(n3345) );
  NAND U2930 ( .A(n3349), .B(n3350), .Z(n3348) );
  NANDN U2931 ( .A(A[187]), .B(B[187]), .Z(n3350) );
  AND U2932 ( .A(n3351), .B(n3352), .Z(n3349) );
  NANDN U2933 ( .A(A[186]), .B(B[186]), .Z(n3352) );
  NAND U2934 ( .A(n3353), .B(n3354), .Z(n3351) );
  NANDN U2935 ( .A(B[186]), .B(A[186]), .Z(n3354) );
  AND U2936 ( .A(n3355), .B(n3356), .Z(n3353) );
  NAND U2937 ( .A(n3357), .B(n3358), .Z(n3356) );
  NANDN U2938 ( .A(A[185]), .B(B[185]), .Z(n3358) );
  AND U2939 ( .A(n3359), .B(n3360), .Z(n3357) );
  NANDN U2940 ( .A(A[184]), .B(B[184]), .Z(n3360) );
  NAND U2941 ( .A(n3361), .B(n3362), .Z(n3359) );
  NANDN U2942 ( .A(B[184]), .B(A[184]), .Z(n3362) );
  AND U2943 ( .A(n3363), .B(n3364), .Z(n3361) );
  NAND U2944 ( .A(n3365), .B(n3366), .Z(n3364) );
  NANDN U2945 ( .A(A[183]), .B(B[183]), .Z(n3366) );
  AND U2946 ( .A(n3367), .B(n3368), .Z(n3365) );
  NANDN U2947 ( .A(A[182]), .B(B[182]), .Z(n3368) );
  NAND U2948 ( .A(n3369), .B(n3370), .Z(n3367) );
  NANDN U2949 ( .A(B[182]), .B(A[182]), .Z(n3370) );
  AND U2950 ( .A(n3371), .B(n3372), .Z(n3369) );
  NAND U2951 ( .A(n3373), .B(n3374), .Z(n3372) );
  NANDN U2952 ( .A(A[181]), .B(B[181]), .Z(n3374) );
  AND U2953 ( .A(n3375), .B(n3376), .Z(n3373) );
  NANDN U2954 ( .A(A[180]), .B(B[180]), .Z(n3376) );
  NAND U2955 ( .A(n3377), .B(n3378), .Z(n3375) );
  NANDN U2956 ( .A(B[180]), .B(A[180]), .Z(n3378) );
  AND U2957 ( .A(n3379), .B(n3380), .Z(n3377) );
  NAND U2958 ( .A(n3381), .B(n3382), .Z(n3380) );
  NANDN U2959 ( .A(A[179]), .B(B[179]), .Z(n3382) );
  AND U2960 ( .A(n3383), .B(n3384), .Z(n3381) );
  NANDN U2961 ( .A(A[178]), .B(B[178]), .Z(n3384) );
  NAND U2962 ( .A(n3385), .B(n3386), .Z(n3383) );
  NANDN U2963 ( .A(B[178]), .B(A[178]), .Z(n3386) );
  AND U2964 ( .A(n3387), .B(n3388), .Z(n3385) );
  NAND U2965 ( .A(n3389), .B(n3390), .Z(n3388) );
  NANDN U2966 ( .A(A[177]), .B(B[177]), .Z(n3390) );
  AND U2967 ( .A(n3391), .B(n3392), .Z(n3389) );
  NANDN U2968 ( .A(A[176]), .B(B[176]), .Z(n3392) );
  NAND U2969 ( .A(n3393), .B(n3394), .Z(n3391) );
  NANDN U2970 ( .A(B[176]), .B(A[176]), .Z(n3394) );
  AND U2971 ( .A(n3395), .B(n3396), .Z(n3393) );
  NAND U2972 ( .A(n3397), .B(n3398), .Z(n3396) );
  NANDN U2973 ( .A(A[175]), .B(B[175]), .Z(n3398) );
  AND U2974 ( .A(n3399), .B(n3400), .Z(n3397) );
  NANDN U2975 ( .A(A[174]), .B(B[174]), .Z(n3400) );
  NAND U2976 ( .A(n3401), .B(n3402), .Z(n3399) );
  NANDN U2977 ( .A(B[174]), .B(A[174]), .Z(n3402) );
  AND U2978 ( .A(n3403), .B(n3404), .Z(n3401) );
  NAND U2979 ( .A(n3405), .B(n3406), .Z(n3404) );
  NANDN U2980 ( .A(A[173]), .B(B[173]), .Z(n3406) );
  AND U2981 ( .A(n3407), .B(n3408), .Z(n3405) );
  NANDN U2982 ( .A(A[172]), .B(B[172]), .Z(n3408) );
  NAND U2983 ( .A(n3409), .B(n3410), .Z(n3407) );
  NANDN U2984 ( .A(B[172]), .B(A[172]), .Z(n3410) );
  AND U2985 ( .A(n3411), .B(n3412), .Z(n3409) );
  NAND U2986 ( .A(n3413), .B(n3414), .Z(n3412) );
  NANDN U2987 ( .A(A[171]), .B(B[171]), .Z(n3414) );
  AND U2988 ( .A(n3415), .B(n3416), .Z(n3413) );
  NANDN U2989 ( .A(A[170]), .B(B[170]), .Z(n3416) );
  NAND U2990 ( .A(n3417), .B(n3418), .Z(n3415) );
  NANDN U2991 ( .A(B[170]), .B(A[170]), .Z(n3418) );
  AND U2992 ( .A(n3419), .B(n3420), .Z(n3417) );
  NAND U2993 ( .A(n3421), .B(n3422), .Z(n3420) );
  NANDN U2994 ( .A(A[169]), .B(B[169]), .Z(n3422) );
  AND U2995 ( .A(n3423), .B(n3424), .Z(n3421) );
  NANDN U2996 ( .A(A[168]), .B(B[168]), .Z(n3424) );
  NAND U2997 ( .A(n3425), .B(n3426), .Z(n3423) );
  NANDN U2998 ( .A(B[168]), .B(A[168]), .Z(n3426) );
  AND U2999 ( .A(n3427), .B(n3428), .Z(n3425) );
  NAND U3000 ( .A(n3429), .B(n3430), .Z(n3428) );
  NANDN U3001 ( .A(A[167]), .B(B[167]), .Z(n3430) );
  AND U3002 ( .A(n3431), .B(n3432), .Z(n3429) );
  NANDN U3003 ( .A(A[166]), .B(B[166]), .Z(n3432) );
  NAND U3004 ( .A(n3433), .B(n3434), .Z(n3431) );
  NANDN U3005 ( .A(B[166]), .B(A[166]), .Z(n3434) );
  AND U3006 ( .A(n3435), .B(n3436), .Z(n3433) );
  NAND U3007 ( .A(n3437), .B(n3438), .Z(n3436) );
  NANDN U3008 ( .A(A[165]), .B(B[165]), .Z(n3438) );
  AND U3009 ( .A(n3439), .B(n3440), .Z(n3437) );
  NANDN U3010 ( .A(A[164]), .B(B[164]), .Z(n3440) );
  NAND U3011 ( .A(n3441), .B(n3442), .Z(n3439) );
  NANDN U3012 ( .A(B[164]), .B(A[164]), .Z(n3442) );
  AND U3013 ( .A(n3443), .B(n3444), .Z(n3441) );
  NAND U3014 ( .A(n3445), .B(n3446), .Z(n3444) );
  NANDN U3015 ( .A(A[163]), .B(B[163]), .Z(n3446) );
  AND U3016 ( .A(n3447), .B(n3448), .Z(n3445) );
  NANDN U3017 ( .A(A[162]), .B(B[162]), .Z(n3448) );
  NAND U3018 ( .A(n3449), .B(n3450), .Z(n3447) );
  NANDN U3019 ( .A(B[162]), .B(A[162]), .Z(n3450) );
  AND U3020 ( .A(n3451), .B(n3452), .Z(n3449) );
  NAND U3021 ( .A(n3453), .B(n3454), .Z(n3452) );
  NANDN U3022 ( .A(A[161]), .B(B[161]), .Z(n3454) );
  AND U3023 ( .A(n3455), .B(n3456), .Z(n3453) );
  NANDN U3024 ( .A(A[160]), .B(B[160]), .Z(n3456) );
  NAND U3025 ( .A(n3457), .B(n3458), .Z(n3455) );
  NANDN U3026 ( .A(B[160]), .B(A[160]), .Z(n3458) );
  AND U3027 ( .A(n3459), .B(n3460), .Z(n3457) );
  NAND U3028 ( .A(n3461), .B(n3462), .Z(n3460) );
  NANDN U3029 ( .A(A[159]), .B(B[159]), .Z(n3462) );
  AND U3030 ( .A(n3463), .B(n3464), .Z(n3461) );
  NANDN U3031 ( .A(A[158]), .B(B[158]), .Z(n3464) );
  NAND U3032 ( .A(n3465), .B(n3466), .Z(n3463) );
  NANDN U3033 ( .A(B[158]), .B(A[158]), .Z(n3466) );
  AND U3034 ( .A(n3467), .B(n3468), .Z(n3465) );
  NAND U3035 ( .A(n3469), .B(n3470), .Z(n3468) );
  NANDN U3036 ( .A(A[157]), .B(B[157]), .Z(n3470) );
  AND U3037 ( .A(n3471), .B(n3472), .Z(n3469) );
  NANDN U3038 ( .A(A[156]), .B(B[156]), .Z(n3472) );
  NAND U3039 ( .A(n3473), .B(n3474), .Z(n3471) );
  NANDN U3040 ( .A(B[156]), .B(A[156]), .Z(n3474) );
  AND U3041 ( .A(n3475), .B(n3476), .Z(n3473) );
  NAND U3042 ( .A(n3477), .B(n3478), .Z(n3476) );
  NANDN U3043 ( .A(A[155]), .B(B[155]), .Z(n3478) );
  AND U3044 ( .A(n3479), .B(n3480), .Z(n3477) );
  NANDN U3045 ( .A(A[154]), .B(B[154]), .Z(n3480) );
  NAND U3046 ( .A(n3481), .B(n3482), .Z(n3479) );
  NANDN U3047 ( .A(B[154]), .B(A[154]), .Z(n3482) );
  AND U3048 ( .A(n3483), .B(n3484), .Z(n3481) );
  NAND U3049 ( .A(n3485), .B(n3486), .Z(n3484) );
  NANDN U3050 ( .A(A[153]), .B(B[153]), .Z(n3486) );
  AND U3051 ( .A(n3487), .B(n3488), .Z(n3485) );
  NANDN U3052 ( .A(A[152]), .B(B[152]), .Z(n3488) );
  NAND U3053 ( .A(n3489), .B(n3490), .Z(n3487) );
  NANDN U3054 ( .A(B[152]), .B(A[152]), .Z(n3490) );
  AND U3055 ( .A(n3491), .B(n3492), .Z(n3489) );
  NAND U3056 ( .A(n3493), .B(n3494), .Z(n3492) );
  NANDN U3057 ( .A(A[151]), .B(B[151]), .Z(n3494) );
  AND U3058 ( .A(n3495), .B(n3496), .Z(n3493) );
  NANDN U3059 ( .A(A[150]), .B(B[150]), .Z(n3496) );
  NAND U3060 ( .A(n3497), .B(n3498), .Z(n3495) );
  NANDN U3061 ( .A(B[150]), .B(A[150]), .Z(n3498) );
  AND U3062 ( .A(n3499), .B(n3500), .Z(n3497) );
  NAND U3063 ( .A(n3501), .B(n3502), .Z(n3500) );
  NANDN U3064 ( .A(A[149]), .B(B[149]), .Z(n3502) );
  AND U3065 ( .A(n3503), .B(n3504), .Z(n3501) );
  NANDN U3066 ( .A(A[148]), .B(B[148]), .Z(n3504) );
  NAND U3067 ( .A(n3505), .B(n3506), .Z(n3503) );
  NANDN U3068 ( .A(B[148]), .B(A[148]), .Z(n3506) );
  AND U3069 ( .A(n3507), .B(n3508), .Z(n3505) );
  NAND U3070 ( .A(n3509), .B(n3510), .Z(n3508) );
  NANDN U3071 ( .A(A[147]), .B(B[147]), .Z(n3510) );
  AND U3072 ( .A(n3511), .B(n3512), .Z(n3509) );
  NANDN U3073 ( .A(A[146]), .B(B[146]), .Z(n3512) );
  NAND U3074 ( .A(n3513), .B(n3514), .Z(n3511) );
  NANDN U3075 ( .A(B[146]), .B(A[146]), .Z(n3514) );
  AND U3076 ( .A(n3515), .B(n3516), .Z(n3513) );
  NAND U3077 ( .A(n3517), .B(n3518), .Z(n3516) );
  NANDN U3078 ( .A(A[145]), .B(B[145]), .Z(n3518) );
  AND U3079 ( .A(n3519), .B(n3520), .Z(n3517) );
  NANDN U3080 ( .A(A[144]), .B(B[144]), .Z(n3520) );
  NAND U3081 ( .A(n3521), .B(n3522), .Z(n3519) );
  NANDN U3082 ( .A(B[144]), .B(A[144]), .Z(n3522) );
  AND U3083 ( .A(n3523), .B(n3524), .Z(n3521) );
  NAND U3084 ( .A(n3525), .B(n3526), .Z(n3524) );
  NANDN U3085 ( .A(A[143]), .B(B[143]), .Z(n3526) );
  AND U3086 ( .A(n3527), .B(n3528), .Z(n3525) );
  NANDN U3087 ( .A(A[142]), .B(B[142]), .Z(n3528) );
  NAND U3088 ( .A(n3529), .B(n3530), .Z(n3527) );
  NANDN U3089 ( .A(B[142]), .B(A[142]), .Z(n3530) );
  AND U3090 ( .A(n3531), .B(n3532), .Z(n3529) );
  NAND U3091 ( .A(n3533), .B(n3534), .Z(n3532) );
  NANDN U3092 ( .A(A[141]), .B(B[141]), .Z(n3534) );
  AND U3093 ( .A(n3535), .B(n3536), .Z(n3533) );
  NANDN U3094 ( .A(A[140]), .B(B[140]), .Z(n3536) );
  NAND U3095 ( .A(n3537), .B(n3538), .Z(n3535) );
  NANDN U3096 ( .A(B[140]), .B(A[140]), .Z(n3538) );
  AND U3097 ( .A(n3539), .B(n3540), .Z(n3537) );
  NAND U3098 ( .A(n3541), .B(n3542), .Z(n3540) );
  NANDN U3099 ( .A(A[139]), .B(B[139]), .Z(n3542) );
  AND U3100 ( .A(n3543), .B(n3544), .Z(n3541) );
  NANDN U3101 ( .A(A[138]), .B(B[138]), .Z(n3544) );
  NAND U3102 ( .A(n3545), .B(n3546), .Z(n3543) );
  NANDN U3103 ( .A(B[138]), .B(A[138]), .Z(n3546) );
  AND U3104 ( .A(n3547), .B(n3548), .Z(n3545) );
  NAND U3105 ( .A(n3549), .B(n3550), .Z(n3548) );
  NANDN U3106 ( .A(A[137]), .B(B[137]), .Z(n3550) );
  AND U3107 ( .A(n3551), .B(n3552), .Z(n3549) );
  NANDN U3108 ( .A(A[136]), .B(B[136]), .Z(n3552) );
  NAND U3109 ( .A(n3553), .B(n3554), .Z(n3551) );
  NANDN U3110 ( .A(B[136]), .B(A[136]), .Z(n3554) );
  AND U3111 ( .A(n3555), .B(n3556), .Z(n3553) );
  NAND U3112 ( .A(n3557), .B(n3558), .Z(n3556) );
  NANDN U3113 ( .A(A[135]), .B(B[135]), .Z(n3558) );
  AND U3114 ( .A(n3559), .B(n3560), .Z(n3557) );
  NANDN U3115 ( .A(A[134]), .B(B[134]), .Z(n3560) );
  NAND U3116 ( .A(n3561), .B(n3562), .Z(n3559) );
  NANDN U3117 ( .A(B[134]), .B(A[134]), .Z(n3562) );
  AND U3118 ( .A(n3563), .B(n3564), .Z(n3561) );
  NAND U3119 ( .A(n3565), .B(n3566), .Z(n3564) );
  NANDN U3120 ( .A(A[133]), .B(B[133]), .Z(n3566) );
  AND U3121 ( .A(n3567), .B(n3568), .Z(n3565) );
  NANDN U3122 ( .A(A[132]), .B(B[132]), .Z(n3568) );
  NAND U3123 ( .A(n3569), .B(n3570), .Z(n3567) );
  NANDN U3124 ( .A(B[132]), .B(A[132]), .Z(n3570) );
  AND U3125 ( .A(n3571), .B(n3572), .Z(n3569) );
  NAND U3126 ( .A(n3573), .B(n3574), .Z(n3572) );
  NANDN U3127 ( .A(A[131]), .B(B[131]), .Z(n3574) );
  AND U3128 ( .A(n3575), .B(n3576), .Z(n3573) );
  NANDN U3129 ( .A(A[130]), .B(B[130]), .Z(n3576) );
  NAND U3130 ( .A(n3577), .B(n3578), .Z(n3575) );
  NANDN U3131 ( .A(B[130]), .B(A[130]), .Z(n3578) );
  AND U3132 ( .A(n3579), .B(n3580), .Z(n3577) );
  NAND U3133 ( .A(n3581), .B(n3582), .Z(n3580) );
  NANDN U3134 ( .A(A[129]), .B(B[129]), .Z(n3582) );
  AND U3135 ( .A(n3583), .B(n3584), .Z(n3581) );
  NANDN U3136 ( .A(A[128]), .B(B[128]), .Z(n3584) );
  NAND U3137 ( .A(n3585), .B(n3586), .Z(n3583) );
  NANDN U3138 ( .A(B[128]), .B(A[128]), .Z(n3586) );
  AND U3139 ( .A(n3587), .B(n3588), .Z(n3585) );
  NAND U3140 ( .A(n3589), .B(n3590), .Z(n3588) );
  NANDN U3141 ( .A(A[127]), .B(B[127]), .Z(n3590) );
  AND U3142 ( .A(n3591), .B(n3592), .Z(n3589) );
  NANDN U3143 ( .A(A[126]), .B(B[126]), .Z(n3592) );
  NAND U3144 ( .A(n3593), .B(n3594), .Z(n3591) );
  NANDN U3145 ( .A(B[126]), .B(A[126]), .Z(n3594) );
  AND U3146 ( .A(n3595), .B(n3596), .Z(n3593) );
  NAND U3147 ( .A(n3597), .B(n3598), .Z(n3596) );
  NANDN U3148 ( .A(A[125]), .B(B[125]), .Z(n3598) );
  AND U3149 ( .A(n3599), .B(n3600), .Z(n3597) );
  NANDN U3150 ( .A(A[124]), .B(B[124]), .Z(n3600) );
  NAND U3151 ( .A(n3601), .B(n3602), .Z(n3599) );
  NANDN U3152 ( .A(B[124]), .B(A[124]), .Z(n3602) );
  AND U3153 ( .A(n3603), .B(n3604), .Z(n3601) );
  NAND U3154 ( .A(n3605), .B(n3606), .Z(n3604) );
  NANDN U3155 ( .A(A[123]), .B(B[123]), .Z(n3606) );
  AND U3156 ( .A(n3607), .B(n3608), .Z(n3605) );
  NANDN U3157 ( .A(A[122]), .B(B[122]), .Z(n3608) );
  NAND U3158 ( .A(n3609), .B(n3610), .Z(n3607) );
  NANDN U3159 ( .A(B[122]), .B(A[122]), .Z(n3610) );
  AND U3160 ( .A(n3611), .B(n3612), .Z(n3609) );
  NAND U3161 ( .A(n3613), .B(n3614), .Z(n3612) );
  NANDN U3162 ( .A(A[121]), .B(B[121]), .Z(n3614) );
  AND U3163 ( .A(n3615), .B(n3616), .Z(n3613) );
  NANDN U3164 ( .A(A[120]), .B(B[120]), .Z(n3616) );
  NAND U3165 ( .A(n3617), .B(n3618), .Z(n3615) );
  NANDN U3166 ( .A(B[120]), .B(A[120]), .Z(n3618) );
  AND U3167 ( .A(n3619), .B(n3620), .Z(n3617) );
  NAND U3168 ( .A(n3621), .B(n3622), .Z(n3620) );
  NANDN U3169 ( .A(A[119]), .B(B[119]), .Z(n3622) );
  AND U3170 ( .A(n3623), .B(n3624), .Z(n3621) );
  NANDN U3171 ( .A(A[118]), .B(B[118]), .Z(n3624) );
  NAND U3172 ( .A(n3625), .B(n3626), .Z(n3623) );
  NANDN U3173 ( .A(B[118]), .B(A[118]), .Z(n3626) );
  AND U3174 ( .A(n3627), .B(n3628), .Z(n3625) );
  NAND U3175 ( .A(n3629), .B(n3630), .Z(n3628) );
  NANDN U3176 ( .A(A[117]), .B(B[117]), .Z(n3630) );
  AND U3177 ( .A(n3631), .B(n3632), .Z(n3629) );
  NANDN U3178 ( .A(A[116]), .B(B[116]), .Z(n3632) );
  NAND U3179 ( .A(n3633), .B(n3634), .Z(n3631) );
  NANDN U3180 ( .A(B[116]), .B(A[116]), .Z(n3634) );
  AND U3181 ( .A(n3635), .B(n3636), .Z(n3633) );
  NAND U3182 ( .A(n3637), .B(n3638), .Z(n3636) );
  NANDN U3183 ( .A(A[115]), .B(B[115]), .Z(n3638) );
  AND U3184 ( .A(n3639), .B(n3640), .Z(n3637) );
  NANDN U3185 ( .A(A[114]), .B(B[114]), .Z(n3640) );
  NAND U3186 ( .A(n3641), .B(n3642), .Z(n3639) );
  NANDN U3187 ( .A(B[114]), .B(A[114]), .Z(n3642) );
  AND U3188 ( .A(n3643), .B(n3644), .Z(n3641) );
  NAND U3189 ( .A(n3645), .B(n3646), .Z(n3644) );
  NANDN U3190 ( .A(A[113]), .B(B[113]), .Z(n3646) );
  AND U3191 ( .A(n3647), .B(n3648), .Z(n3645) );
  NANDN U3192 ( .A(A[112]), .B(B[112]), .Z(n3648) );
  NAND U3193 ( .A(n3649), .B(n3650), .Z(n3647) );
  NANDN U3194 ( .A(B[112]), .B(A[112]), .Z(n3650) );
  AND U3195 ( .A(n3651), .B(n3652), .Z(n3649) );
  NAND U3196 ( .A(n3653), .B(n3654), .Z(n3652) );
  NANDN U3197 ( .A(A[111]), .B(B[111]), .Z(n3654) );
  AND U3198 ( .A(n3655), .B(n3656), .Z(n3653) );
  NANDN U3199 ( .A(A[110]), .B(B[110]), .Z(n3656) );
  NAND U3200 ( .A(n3657), .B(n3658), .Z(n3655) );
  NANDN U3201 ( .A(B[110]), .B(A[110]), .Z(n3658) );
  AND U3202 ( .A(n3659), .B(n3660), .Z(n3657) );
  NAND U3203 ( .A(n3661), .B(n3662), .Z(n3660) );
  NANDN U3204 ( .A(A[109]), .B(B[109]), .Z(n3662) );
  AND U3205 ( .A(n3663), .B(n3664), .Z(n3661) );
  NANDN U3206 ( .A(A[108]), .B(B[108]), .Z(n3664) );
  NAND U3207 ( .A(n3665), .B(n3666), .Z(n3663) );
  NANDN U3208 ( .A(B[108]), .B(A[108]), .Z(n3666) );
  AND U3209 ( .A(n3667), .B(n3668), .Z(n3665) );
  NAND U3210 ( .A(n3669), .B(n3670), .Z(n3668) );
  NANDN U3211 ( .A(A[107]), .B(B[107]), .Z(n3670) );
  AND U3212 ( .A(n3671), .B(n3672), .Z(n3669) );
  NANDN U3213 ( .A(A[106]), .B(B[106]), .Z(n3672) );
  NAND U3214 ( .A(n3673), .B(n3674), .Z(n3671) );
  NANDN U3215 ( .A(B[106]), .B(A[106]), .Z(n3674) );
  AND U3216 ( .A(n3675), .B(n3676), .Z(n3673) );
  NAND U3217 ( .A(n3677), .B(n3678), .Z(n3676) );
  NANDN U3218 ( .A(A[105]), .B(B[105]), .Z(n3678) );
  AND U3219 ( .A(n3679), .B(n3680), .Z(n3677) );
  NANDN U3220 ( .A(A[104]), .B(B[104]), .Z(n3680) );
  NAND U3221 ( .A(n3681), .B(n3682), .Z(n3679) );
  NANDN U3222 ( .A(B[104]), .B(A[104]), .Z(n3682) );
  AND U3223 ( .A(n3683), .B(n3684), .Z(n3681) );
  NAND U3224 ( .A(n3685), .B(n3686), .Z(n3684) );
  NANDN U3225 ( .A(A[103]), .B(B[103]), .Z(n3686) );
  AND U3226 ( .A(n3687), .B(n3688), .Z(n3685) );
  NANDN U3227 ( .A(A[102]), .B(B[102]), .Z(n3688) );
  NAND U3228 ( .A(n3689), .B(n3690), .Z(n3687) );
  NANDN U3229 ( .A(B[102]), .B(A[102]), .Z(n3690) );
  AND U3230 ( .A(n3691), .B(n3692), .Z(n3689) );
  NAND U3231 ( .A(n3693), .B(n3694), .Z(n3692) );
  NANDN U3232 ( .A(A[101]), .B(B[101]), .Z(n3694) );
  AND U3233 ( .A(n3695), .B(n3696), .Z(n3693) );
  NANDN U3234 ( .A(A[100]), .B(B[100]), .Z(n3696) );
  NAND U3235 ( .A(n3697), .B(n3698), .Z(n3695) );
  NANDN U3236 ( .A(B[99]), .B(A[99]), .Z(n3698) );
  AND U3237 ( .A(n3699), .B(n3700), .Z(n3697) );
  NAND U3238 ( .A(n3701), .B(n3702), .Z(n3700) );
  NANDN U3239 ( .A(A[99]), .B(B[99]), .Z(n3702) );
  AND U3240 ( .A(n3703), .B(n3704), .Z(n3701) );
  NANDN U3241 ( .A(A[98]), .B(B[98]), .Z(n3704) );
  NAND U3242 ( .A(n3705), .B(n3706), .Z(n3703) );
  NANDN U3243 ( .A(B[98]), .B(A[98]), .Z(n3706) );
  AND U3244 ( .A(n3707), .B(n3708), .Z(n3705) );
  NAND U3245 ( .A(n3709), .B(n3710), .Z(n3708) );
  NANDN U3246 ( .A(A[97]), .B(B[97]), .Z(n3710) );
  AND U3247 ( .A(n3711), .B(n3712), .Z(n3709) );
  NANDN U3248 ( .A(A[96]), .B(B[96]), .Z(n3712) );
  NAND U3249 ( .A(n3713), .B(n3714), .Z(n3711) );
  NANDN U3250 ( .A(B[96]), .B(A[96]), .Z(n3714) );
  AND U3251 ( .A(n3715), .B(n3716), .Z(n3713) );
  NAND U3252 ( .A(n3717), .B(n3718), .Z(n3716) );
  NANDN U3253 ( .A(A[95]), .B(B[95]), .Z(n3718) );
  AND U3254 ( .A(n3719), .B(n3720), .Z(n3717) );
  NANDN U3255 ( .A(A[94]), .B(B[94]), .Z(n3720) );
  NAND U3256 ( .A(n3721), .B(n3722), .Z(n3719) );
  NANDN U3257 ( .A(B[94]), .B(A[94]), .Z(n3722) );
  AND U3258 ( .A(n3723), .B(n3724), .Z(n3721) );
  NAND U3259 ( .A(n3725), .B(n3726), .Z(n3724) );
  NANDN U3260 ( .A(A[93]), .B(B[93]), .Z(n3726) );
  AND U3261 ( .A(n3727), .B(n3728), .Z(n3725) );
  NANDN U3262 ( .A(A[92]), .B(B[92]), .Z(n3728) );
  NAND U3263 ( .A(n3729), .B(n3730), .Z(n3727) );
  NANDN U3264 ( .A(B[92]), .B(A[92]), .Z(n3730) );
  AND U3265 ( .A(n3731), .B(n3732), .Z(n3729) );
  NAND U3266 ( .A(n3733), .B(n3734), .Z(n3732) );
  NANDN U3267 ( .A(A[91]), .B(B[91]), .Z(n3734) );
  AND U3268 ( .A(n3735), .B(n3736), .Z(n3733) );
  NANDN U3269 ( .A(A[90]), .B(B[90]), .Z(n3736) );
  NAND U3270 ( .A(n3737), .B(n3738), .Z(n3735) );
  NANDN U3271 ( .A(B[90]), .B(A[90]), .Z(n3738) );
  AND U3272 ( .A(n3739), .B(n3740), .Z(n3737) );
  NAND U3273 ( .A(n3741), .B(n3742), .Z(n3740) );
  NANDN U3274 ( .A(A[89]), .B(B[89]), .Z(n3742) );
  AND U3275 ( .A(n3743), .B(n3744), .Z(n3741) );
  NANDN U3276 ( .A(A[88]), .B(B[88]), .Z(n3744) );
  NAND U3277 ( .A(n3745), .B(n3746), .Z(n3743) );
  NANDN U3278 ( .A(B[88]), .B(A[88]), .Z(n3746) );
  AND U3279 ( .A(n3747), .B(n3748), .Z(n3745) );
  NAND U3280 ( .A(n3749), .B(n3750), .Z(n3748) );
  NANDN U3281 ( .A(A[87]), .B(B[87]), .Z(n3750) );
  AND U3282 ( .A(n3751), .B(n3752), .Z(n3749) );
  NANDN U3283 ( .A(A[86]), .B(B[86]), .Z(n3752) );
  NAND U3284 ( .A(n3753), .B(n3754), .Z(n3751) );
  NANDN U3285 ( .A(B[86]), .B(A[86]), .Z(n3754) );
  AND U3286 ( .A(n3755), .B(n3756), .Z(n3753) );
  NAND U3287 ( .A(n3757), .B(n3758), .Z(n3756) );
  NANDN U3288 ( .A(A[85]), .B(B[85]), .Z(n3758) );
  AND U3289 ( .A(n3759), .B(n3760), .Z(n3757) );
  NANDN U3290 ( .A(A[84]), .B(B[84]), .Z(n3760) );
  NAND U3291 ( .A(n3761), .B(n3762), .Z(n3759) );
  NANDN U3292 ( .A(B[84]), .B(A[84]), .Z(n3762) );
  AND U3293 ( .A(n3763), .B(n3764), .Z(n3761) );
  NAND U3294 ( .A(n3765), .B(n3766), .Z(n3764) );
  NANDN U3295 ( .A(A[83]), .B(B[83]), .Z(n3766) );
  AND U3296 ( .A(n3767), .B(n3768), .Z(n3765) );
  NANDN U3297 ( .A(A[82]), .B(B[82]), .Z(n3768) );
  NAND U3298 ( .A(n3769), .B(n3770), .Z(n3767) );
  NANDN U3299 ( .A(B[82]), .B(A[82]), .Z(n3770) );
  AND U3300 ( .A(n3771), .B(n3772), .Z(n3769) );
  NAND U3301 ( .A(n3773), .B(n3774), .Z(n3772) );
  NANDN U3302 ( .A(A[81]), .B(B[81]), .Z(n3774) );
  AND U3303 ( .A(n3775), .B(n3776), .Z(n3773) );
  NANDN U3304 ( .A(A[80]), .B(B[80]), .Z(n3776) );
  NAND U3305 ( .A(n3777), .B(n3778), .Z(n3775) );
  NANDN U3306 ( .A(B[80]), .B(A[80]), .Z(n3778) );
  AND U3307 ( .A(n3779), .B(n3780), .Z(n3777) );
  NAND U3308 ( .A(n3781), .B(n3782), .Z(n3780) );
  NANDN U3309 ( .A(A[79]), .B(B[79]), .Z(n3782) );
  AND U3310 ( .A(n3783), .B(n3784), .Z(n3781) );
  NANDN U3311 ( .A(A[78]), .B(B[78]), .Z(n3784) );
  NAND U3312 ( .A(n3785), .B(n3786), .Z(n3783) );
  NANDN U3313 ( .A(B[78]), .B(A[78]), .Z(n3786) );
  AND U3314 ( .A(n3787), .B(n3788), .Z(n3785) );
  NAND U3315 ( .A(n3789), .B(n3790), .Z(n3788) );
  NANDN U3316 ( .A(A[77]), .B(B[77]), .Z(n3790) );
  AND U3317 ( .A(n3791), .B(n3792), .Z(n3789) );
  NANDN U3318 ( .A(A[76]), .B(B[76]), .Z(n3792) );
  NAND U3319 ( .A(n3793), .B(n3794), .Z(n3791) );
  NANDN U3320 ( .A(B[76]), .B(A[76]), .Z(n3794) );
  AND U3321 ( .A(n3795), .B(n3796), .Z(n3793) );
  NAND U3322 ( .A(n3797), .B(n3798), .Z(n3796) );
  NANDN U3323 ( .A(A[75]), .B(B[75]), .Z(n3798) );
  AND U3324 ( .A(n3799), .B(n3800), .Z(n3797) );
  NANDN U3325 ( .A(A[74]), .B(B[74]), .Z(n3800) );
  NAND U3326 ( .A(n3801), .B(n3802), .Z(n3799) );
  NANDN U3327 ( .A(B[74]), .B(A[74]), .Z(n3802) );
  AND U3328 ( .A(n3803), .B(n3804), .Z(n3801) );
  NAND U3329 ( .A(n3805), .B(n3806), .Z(n3804) );
  NANDN U3330 ( .A(A[73]), .B(B[73]), .Z(n3806) );
  AND U3331 ( .A(n3807), .B(n3808), .Z(n3805) );
  NANDN U3332 ( .A(A[72]), .B(B[72]), .Z(n3808) );
  NAND U3333 ( .A(n3809), .B(n3810), .Z(n3807) );
  NANDN U3334 ( .A(B[72]), .B(A[72]), .Z(n3810) );
  AND U3335 ( .A(n3811), .B(n3812), .Z(n3809) );
  NAND U3336 ( .A(n3813), .B(n3814), .Z(n3812) );
  NANDN U3337 ( .A(A[71]), .B(B[71]), .Z(n3814) );
  AND U3338 ( .A(n3815), .B(n3816), .Z(n3813) );
  NANDN U3339 ( .A(A[70]), .B(B[70]), .Z(n3816) );
  NAND U3340 ( .A(n3817), .B(n3818), .Z(n3815) );
  NANDN U3341 ( .A(B[70]), .B(A[70]), .Z(n3818) );
  AND U3342 ( .A(n3819), .B(n3820), .Z(n3817) );
  NAND U3343 ( .A(n3821), .B(n3822), .Z(n3820) );
  NANDN U3344 ( .A(A[69]), .B(B[69]), .Z(n3822) );
  AND U3345 ( .A(n3823), .B(n3824), .Z(n3821) );
  NANDN U3346 ( .A(A[68]), .B(B[68]), .Z(n3824) );
  NAND U3347 ( .A(n3825), .B(n3826), .Z(n3823) );
  NANDN U3348 ( .A(B[68]), .B(A[68]), .Z(n3826) );
  AND U3349 ( .A(n3827), .B(n3828), .Z(n3825) );
  NAND U3350 ( .A(n3829), .B(n3830), .Z(n3828) );
  NANDN U3351 ( .A(A[67]), .B(B[67]), .Z(n3830) );
  AND U3352 ( .A(n3831), .B(n3832), .Z(n3829) );
  NANDN U3353 ( .A(A[66]), .B(B[66]), .Z(n3832) );
  NAND U3354 ( .A(n3833), .B(n3834), .Z(n3831) );
  NANDN U3355 ( .A(B[66]), .B(A[66]), .Z(n3834) );
  AND U3356 ( .A(n3835), .B(n3836), .Z(n3833) );
  NAND U3357 ( .A(n3837), .B(n3838), .Z(n3836) );
  NANDN U3358 ( .A(A[65]), .B(B[65]), .Z(n3838) );
  AND U3359 ( .A(n3839), .B(n3840), .Z(n3837) );
  NANDN U3360 ( .A(A[64]), .B(B[64]), .Z(n3840) );
  NAND U3361 ( .A(n3841), .B(n3842), .Z(n3839) );
  NANDN U3362 ( .A(B[64]), .B(A[64]), .Z(n3842) );
  AND U3363 ( .A(n3843), .B(n3844), .Z(n3841) );
  NAND U3364 ( .A(n3845), .B(n3846), .Z(n3844) );
  NANDN U3365 ( .A(A[63]), .B(B[63]), .Z(n3846) );
  AND U3366 ( .A(n3847), .B(n3848), .Z(n3845) );
  NANDN U3367 ( .A(A[62]), .B(B[62]), .Z(n3848) );
  NAND U3368 ( .A(n3849), .B(n3850), .Z(n3847) );
  NANDN U3369 ( .A(B[62]), .B(A[62]), .Z(n3850) );
  AND U3370 ( .A(n3851), .B(n3852), .Z(n3849) );
  NAND U3371 ( .A(n3853), .B(n3854), .Z(n3852) );
  NANDN U3372 ( .A(A[61]), .B(B[61]), .Z(n3854) );
  AND U3373 ( .A(n3855), .B(n3856), .Z(n3853) );
  NANDN U3374 ( .A(A[60]), .B(B[60]), .Z(n3856) );
  NAND U3375 ( .A(n3857), .B(n3858), .Z(n3855) );
  NANDN U3376 ( .A(B[60]), .B(A[60]), .Z(n3858) );
  AND U3377 ( .A(n3859), .B(n3860), .Z(n3857) );
  NAND U3378 ( .A(n3861), .B(n3862), .Z(n3860) );
  NANDN U3379 ( .A(A[59]), .B(B[59]), .Z(n3862) );
  AND U3380 ( .A(n3863), .B(n3864), .Z(n3861) );
  NANDN U3381 ( .A(A[58]), .B(B[58]), .Z(n3864) );
  NAND U3382 ( .A(n3865), .B(n3866), .Z(n3863) );
  NANDN U3383 ( .A(B[58]), .B(A[58]), .Z(n3866) );
  AND U3384 ( .A(n3867), .B(n3868), .Z(n3865) );
  NAND U3385 ( .A(n3869), .B(n3870), .Z(n3868) );
  NANDN U3386 ( .A(A[57]), .B(B[57]), .Z(n3870) );
  AND U3387 ( .A(n3871), .B(n3872), .Z(n3869) );
  NANDN U3388 ( .A(A[56]), .B(B[56]), .Z(n3872) );
  NAND U3389 ( .A(n3873), .B(n3874), .Z(n3871) );
  NANDN U3390 ( .A(B[56]), .B(A[56]), .Z(n3874) );
  AND U3391 ( .A(n3875), .B(n3876), .Z(n3873) );
  NAND U3392 ( .A(n3877), .B(n3878), .Z(n3876) );
  NANDN U3393 ( .A(A[55]), .B(B[55]), .Z(n3878) );
  AND U3394 ( .A(n3879), .B(n3880), .Z(n3877) );
  NANDN U3395 ( .A(A[54]), .B(B[54]), .Z(n3880) );
  NAND U3396 ( .A(n3881), .B(n3882), .Z(n3879) );
  NANDN U3397 ( .A(B[54]), .B(A[54]), .Z(n3882) );
  AND U3398 ( .A(n3883), .B(n3884), .Z(n3881) );
  NAND U3399 ( .A(n3885), .B(n3886), .Z(n3884) );
  NANDN U3400 ( .A(A[53]), .B(B[53]), .Z(n3886) );
  AND U3401 ( .A(n3887), .B(n3888), .Z(n3885) );
  NANDN U3402 ( .A(A[52]), .B(B[52]), .Z(n3888) );
  NAND U3403 ( .A(n3889), .B(n3890), .Z(n3887) );
  NANDN U3404 ( .A(B[52]), .B(A[52]), .Z(n3890) );
  AND U3405 ( .A(n3891), .B(n3892), .Z(n3889) );
  NAND U3406 ( .A(n3893), .B(n3894), .Z(n3892) );
  NANDN U3407 ( .A(A[51]), .B(B[51]), .Z(n3894) );
  AND U3408 ( .A(n3895), .B(n3896), .Z(n3893) );
  NANDN U3409 ( .A(A[50]), .B(B[50]), .Z(n3896) );
  NAND U3410 ( .A(n3897), .B(n3898), .Z(n3895) );
  NANDN U3411 ( .A(B[50]), .B(A[50]), .Z(n3898) );
  AND U3412 ( .A(n3899), .B(n3900), .Z(n3897) );
  NAND U3413 ( .A(n3901), .B(n3902), .Z(n3900) );
  NANDN U3414 ( .A(A[49]), .B(B[49]), .Z(n3902) );
  AND U3415 ( .A(n3903), .B(n3904), .Z(n3901) );
  NANDN U3416 ( .A(A[48]), .B(B[48]), .Z(n3904) );
  NAND U3417 ( .A(n3905), .B(n3906), .Z(n3903) );
  NANDN U3418 ( .A(B[48]), .B(A[48]), .Z(n3906) );
  AND U3419 ( .A(n3907), .B(n3908), .Z(n3905) );
  NAND U3420 ( .A(n3909), .B(n3910), .Z(n3908) );
  NANDN U3421 ( .A(A[47]), .B(B[47]), .Z(n3910) );
  AND U3422 ( .A(n3911), .B(n3912), .Z(n3909) );
  NANDN U3423 ( .A(A[46]), .B(B[46]), .Z(n3912) );
  NAND U3424 ( .A(n3913), .B(n3914), .Z(n3911) );
  NANDN U3425 ( .A(B[46]), .B(A[46]), .Z(n3914) );
  AND U3426 ( .A(n3915), .B(n3916), .Z(n3913) );
  NAND U3427 ( .A(n3917), .B(n3918), .Z(n3916) );
  NANDN U3428 ( .A(A[45]), .B(B[45]), .Z(n3918) );
  AND U3429 ( .A(n3919), .B(n3920), .Z(n3917) );
  NANDN U3430 ( .A(A[44]), .B(B[44]), .Z(n3920) );
  NAND U3431 ( .A(n3921), .B(n3922), .Z(n3919) );
  NANDN U3432 ( .A(B[44]), .B(A[44]), .Z(n3922) );
  AND U3433 ( .A(n3923), .B(n3924), .Z(n3921) );
  NAND U3434 ( .A(n3925), .B(n3926), .Z(n3924) );
  NANDN U3435 ( .A(A[43]), .B(B[43]), .Z(n3926) );
  AND U3436 ( .A(n3927), .B(n3928), .Z(n3925) );
  NANDN U3437 ( .A(A[42]), .B(B[42]), .Z(n3928) );
  NAND U3438 ( .A(n3929), .B(n3930), .Z(n3927) );
  NANDN U3439 ( .A(B[42]), .B(A[42]), .Z(n3930) );
  AND U3440 ( .A(n3931), .B(n3932), .Z(n3929) );
  NAND U3441 ( .A(n3933), .B(n3934), .Z(n3932) );
  NANDN U3442 ( .A(A[41]), .B(B[41]), .Z(n3934) );
  AND U3443 ( .A(n3935), .B(n3936), .Z(n3933) );
  NANDN U3444 ( .A(A[40]), .B(B[40]), .Z(n3936) );
  NAND U3445 ( .A(n3937), .B(n3938), .Z(n3935) );
  NANDN U3446 ( .A(B[40]), .B(A[40]), .Z(n3938) );
  AND U3447 ( .A(n3939), .B(n3940), .Z(n3937) );
  NAND U3448 ( .A(n3941), .B(n3942), .Z(n3940) );
  NANDN U3449 ( .A(A[39]), .B(B[39]), .Z(n3942) );
  AND U3450 ( .A(n3943), .B(n3944), .Z(n3941) );
  NANDN U3451 ( .A(A[38]), .B(B[38]), .Z(n3944) );
  NAND U3452 ( .A(n3945), .B(n3946), .Z(n3943) );
  NANDN U3453 ( .A(B[38]), .B(A[38]), .Z(n3946) );
  AND U3454 ( .A(n3947), .B(n3948), .Z(n3945) );
  NAND U3455 ( .A(n3949), .B(n3950), .Z(n3948) );
  NANDN U3456 ( .A(A[37]), .B(B[37]), .Z(n3950) );
  AND U3457 ( .A(n3951), .B(n3952), .Z(n3949) );
  NANDN U3458 ( .A(A[36]), .B(B[36]), .Z(n3952) );
  NAND U3459 ( .A(n3953), .B(n3954), .Z(n3951) );
  NANDN U3460 ( .A(B[36]), .B(A[36]), .Z(n3954) );
  AND U3461 ( .A(n3955), .B(n3956), .Z(n3953) );
  NAND U3462 ( .A(n3957), .B(n3958), .Z(n3956) );
  NANDN U3463 ( .A(A[35]), .B(B[35]), .Z(n3958) );
  AND U3464 ( .A(n3959), .B(n3960), .Z(n3957) );
  NANDN U3465 ( .A(A[34]), .B(B[34]), .Z(n3960) );
  NAND U3466 ( .A(n3961), .B(n3962), .Z(n3959) );
  NANDN U3467 ( .A(B[34]), .B(A[34]), .Z(n3962) );
  AND U3468 ( .A(n3963), .B(n3964), .Z(n3961) );
  NAND U3469 ( .A(n3965), .B(n3966), .Z(n3964) );
  NANDN U3470 ( .A(A[33]), .B(B[33]), .Z(n3966) );
  AND U3471 ( .A(n3967), .B(n3968), .Z(n3965) );
  NANDN U3472 ( .A(A[32]), .B(B[32]), .Z(n3968) );
  NAND U3473 ( .A(n3969), .B(n3970), .Z(n3967) );
  NANDN U3474 ( .A(B[32]), .B(A[32]), .Z(n3970) );
  AND U3475 ( .A(n3971), .B(n3972), .Z(n3969) );
  NAND U3476 ( .A(n3973), .B(n3974), .Z(n3972) );
  NANDN U3477 ( .A(A[31]), .B(B[31]), .Z(n3974) );
  AND U3478 ( .A(n3975), .B(n3976), .Z(n3973) );
  NANDN U3479 ( .A(A[30]), .B(B[30]), .Z(n3976) );
  NAND U3480 ( .A(n3977), .B(n3978), .Z(n3975) );
  NANDN U3481 ( .A(B[30]), .B(A[30]), .Z(n3978) );
  AND U3482 ( .A(n3979), .B(n3980), .Z(n3977) );
  NAND U3483 ( .A(n3981), .B(n3982), .Z(n3980) );
  NANDN U3484 ( .A(A[29]), .B(B[29]), .Z(n3982) );
  AND U3485 ( .A(n3983), .B(n3984), .Z(n3981) );
  NANDN U3486 ( .A(A[28]), .B(B[28]), .Z(n3984) );
  NAND U3487 ( .A(n3985), .B(n3986), .Z(n3983) );
  NANDN U3488 ( .A(B[28]), .B(A[28]), .Z(n3986) );
  AND U3489 ( .A(n3987), .B(n3988), .Z(n3985) );
  NAND U3490 ( .A(n3989), .B(n3990), .Z(n3988) );
  NANDN U3491 ( .A(A[27]), .B(B[27]), .Z(n3990) );
  AND U3492 ( .A(n3991), .B(n3992), .Z(n3989) );
  NANDN U3493 ( .A(A[26]), .B(B[26]), .Z(n3992) );
  NAND U3494 ( .A(n3993), .B(n3994), .Z(n3991) );
  NANDN U3495 ( .A(B[26]), .B(A[26]), .Z(n3994) );
  AND U3496 ( .A(n3995), .B(n3996), .Z(n3993) );
  NAND U3497 ( .A(n3997), .B(n3998), .Z(n3996) );
  NANDN U3498 ( .A(A[25]), .B(B[25]), .Z(n3998) );
  AND U3499 ( .A(n3999), .B(n4000), .Z(n3997) );
  NANDN U3500 ( .A(A[24]), .B(B[24]), .Z(n4000) );
  NAND U3501 ( .A(n4001), .B(n4002), .Z(n3999) );
  NANDN U3502 ( .A(B[24]), .B(A[24]), .Z(n4002) );
  AND U3503 ( .A(n4003), .B(n4004), .Z(n4001) );
  NAND U3504 ( .A(n4005), .B(n4006), .Z(n4004) );
  NANDN U3505 ( .A(A[23]), .B(B[23]), .Z(n4006) );
  AND U3506 ( .A(n4007), .B(n4008), .Z(n4005) );
  NANDN U3507 ( .A(A[22]), .B(B[22]), .Z(n4008) );
  NAND U3508 ( .A(n4009), .B(n4010), .Z(n4007) );
  NANDN U3509 ( .A(B[22]), .B(A[22]), .Z(n4010) );
  AND U3510 ( .A(n4011), .B(n4012), .Z(n4009) );
  NAND U3511 ( .A(n4013), .B(n4014), .Z(n4012) );
  NANDN U3512 ( .A(A[21]), .B(B[21]), .Z(n4014) );
  AND U3513 ( .A(n4015), .B(n4016), .Z(n4013) );
  NANDN U3514 ( .A(A[20]), .B(B[20]), .Z(n4016) );
  NAND U3515 ( .A(n4017), .B(n4018), .Z(n4015) );
  NANDN U3516 ( .A(B[20]), .B(A[20]), .Z(n4018) );
  AND U3517 ( .A(n4019), .B(n4020), .Z(n4017) );
  NAND U3518 ( .A(n4021), .B(n4022), .Z(n4020) );
  NANDN U3519 ( .A(A[19]), .B(B[19]), .Z(n4022) );
  AND U3520 ( .A(n4023), .B(n4024), .Z(n4021) );
  NANDN U3521 ( .A(A[18]), .B(B[18]), .Z(n4024) );
  NAND U3522 ( .A(n4025), .B(n4026), .Z(n4023) );
  NANDN U3523 ( .A(B[18]), .B(A[18]), .Z(n4026) );
  AND U3524 ( .A(n4027), .B(n4028), .Z(n4025) );
  NAND U3525 ( .A(n4029), .B(n4030), .Z(n4028) );
  NANDN U3526 ( .A(A[17]), .B(B[17]), .Z(n4030) );
  AND U3527 ( .A(n4031), .B(n4032), .Z(n4029) );
  NANDN U3528 ( .A(A[16]), .B(B[16]), .Z(n4032) );
  NAND U3529 ( .A(n4033), .B(n4034), .Z(n4031) );
  NANDN U3530 ( .A(B[16]), .B(A[16]), .Z(n4034) );
  AND U3531 ( .A(n4035), .B(n4036), .Z(n4033) );
  NAND U3532 ( .A(n4037), .B(n4038), .Z(n4036) );
  NANDN U3533 ( .A(A[15]), .B(B[15]), .Z(n4038) );
  AND U3534 ( .A(n4039), .B(n4040), .Z(n4037) );
  NANDN U3535 ( .A(A[14]), .B(B[14]), .Z(n4040) );
  NAND U3536 ( .A(n4041), .B(n4042), .Z(n4039) );
  NANDN U3537 ( .A(B[14]), .B(A[14]), .Z(n4042) );
  AND U3538 ( .A(n4043), .B(n4044), .Z(n4041) );
  NAND U3539 ( .A(n4045), .B(n4046), .Z(n4044) );
  NANDN U3540 ( .A(A[13]), .B(B[13]), .Z(n4046) );
  AND U3541 ( .A(n4047), .B(n4048), .Z(n4045) );
  NANDN U3542 ( .A(A[12]), .B(B[12]), .Z(n4048) );
  NAND U3543 ( .A(n4049), .B(n4050), .Z(n4047) );
  NANDN U3544 ( .A(B[12]), .B(A[12]), .Z(n4050) );
  AND U3545 ( .A(n4051), .B(n4052), .Z(n4049) );
  NAND U3546 ( .A(n4053), .B(n4054), .Z(n4052) );
  NANDN U3547 ( .A(A[11]), .B(B[11]), .Z(n4054) );
  AND U3548 ( .A(n4055), .B(n4056), .Z(n4053) );
  NANDN U3549 ( .A(A[10]), .B(B[10]), .Z(n4056) );
  NAND U3550 ( .A(n4057), .B(n4058), .Z(n4055) );
  NANDN U3551 ( .A(B[9]), .B(A[9]), .Z(n4058) );
  AND U3552 ( .A(n4059), .B(n4060), .Z(n4057) );
  NAND U3553 ( .A(n4061), .B(n4062), .Z(n4060) );
  NANDN U3554 ( .A(A[9]), .B(B[9]), .Z(n4062) );
  AND U3555 ( .A(n4063), .B(n4064), .Z(n4061) );
  NANDN U3556 ( .A(A[8]), .B(B[8]), .Z(n4064) );
  NAND U3557 ( .A(n4065), .B(n4066), .Z(n4063) );
  NANDN U3558 ( .A(B[8]), .B(A[8]), .Z(n4066) );
  AND U3559 ( .A(n4067), .B(n4068), .Z(n4065) );
  NAND U3560 ( .A(n4069), .B(n4070), .Z(n4068) );
  NANDN U3561 ( .A(A[7]), .B(B[7]), .Z(n4070) );
  AND U3562 ( .A(n4071), .B(n4072), .Z(n4069) );
  NANDN U3563 ( .A(A[6]), .B(B[6]), .Z(n4072) );
  NAND U3564 ( .A(n4073), .B(n4074), .Z(n4071) );
  NANDN U3565 ( .A(B[6]), .B(A[6]), .Z(n4074) );
  AND U3566 ( .A(n4075), .B(n4076), .Z(n4073) );
  NAND U3567 ( .A(n4077), .B(n4078), .Z(n4076) );
  NANDN U3568 ( .A(A[5]), .B(B[5]), .Z(n4078) );
  AND U3569 ( .A(n4079), .B(n4080), .Z(n4077) );
  NANDN U3570 ( .A(A[4]), .B(B[4]), .Z(n4080) );
  NAND U3571 ( .A(n4081), .B(n4082), .Z(n4079) );
  NANDN U3572 ( .A(B[4]), .B(A[4]), .Z(n4082) );
  AND U3573 ( .A(n4083), .B(n4084), .Z(n4081) );
  NAND U3574 ( .A(n4085), .B(n4086), .Z(n4084) );
  NANDN U3575 ( .A(A[3]), .B(B[3]), .Z(n4086) );
  AND U3576 ( .A(n4087), .B(n4088), .Z(n4085) );
  NANDN U3577 ( .A(A[2]), .B(B[2]), .Z(n4088) );
  NAND U3578 ( .A(n4089), .B(n4090), .Z(n4087) );
  NANDN U3579 ( .A(B[2]), .B(A[2]), .Z(n4090) );
  AND U3580 ( .A(n4091), .B(n4092), .Z(n4089) );
  NANDN U3581 ( .A(B[1]), .B(n4093), .Z(n4092) );
  NANDN U3582 ( .A(A[1]), .B(n4094), .Z(n4093) );
  NANDN U3583 ( .A(n4094), .B(A[1]), .Z(n4091) );
  ANDN U3584 ( .B(B[0]), .A(A[0]), .Z(n4094) );
  NANDN U3585 ( .A(B[3]), .B(A[3]), .Z(n4083) );
  NANDN U3586 ( .A(B[5]), .B(A[5]), .Z(n4075) );
  NANDN U3587 ( .A(B[7]), .B(A[7]), .Z(n4067) );
  NANDN U3588 ( .A(B[10]), .B(A[10]), .Z(n4059) );
  NANDN U3589 ( .A(B[11]), .B(A[11]), .Z(n4051) );
  NANDN U3590 ( .A(B[13]), .B(A[13]), .Z(n4043) );
  NANDN U3591 ( .A(B[15]), .B(A[15]), .Z(n4035) );
  NANDN U3592 ( .A(B[17]), .B(A[17]), .Z(n4027) );
  NANDN U3593 ( .A(B[19]), .B(A[19]), .Z(n4019) );
  NANDN U3594 ( .A(B[21]), .B(A[21]), .Z(n4011) );
  NANDN U3595 ( .A(B[23]), .B(A[23]), .Z(n4003) );
  NANDN U3596 ( .A(B[25]), .B(A[25]), .Z(n3995) );
  NANDN U3597 ( .A(B[27]), .B(A[27]), .Z(n3987) );
  NANDN U3598 ( .A(B[29]), .B(A[29]), .Z(n3979) );
  NANDN U3599 ( .A(B[31]), .B(A[31]), .Z(n3971) );
  NANDN U3600 ( .A(B[33]), .B(A[33]), .Z(n3963) );
  NANDN U3601 ( .A(B[35]), .B(A[35]), .Z(n3955) );
  NANDN U3602 ( .A(B[37]), .B(A[37]), .Z(n3947) );
  NANDN U3603 ( .A(B[39]), .B(A[39]), .Z(n3939) );
  NANDN U3604 ( .A(B[41]), .B(A[41]), .Z(n3931) );
  NANDN U3605 ( .A(B[43]), .B(A[43]), .Z(n3923) );
  NANDN U3606 ( .A(B[45]), .B(A[45]), .Z(n3915) );
  NANDN U3607 ( .A(B[47]), .B(A[47]), .Z(n3907) );
  NANDN U3608 ( .A(B[49]), .B(A[49]), .Z(n3899) );
  NANDN U3609 ( .A(B[51]), .B(A[51]), .Z(n3891) );
  NANDN U3610 ( .A(B[53]), .B(A[53]), .Z(n3883) );
  NANDN U3611 ( .A(B[55]), .B(A[55]), .Z(n3875) );
  NANDN U3612 ( .A(B[57]), .B(A[57]), .Z(n3867) );
  NANDN U3613 ( .A(B[59]), .B(A[59]), .Z(n3859) );
  NANDN U3614 ( .A(B[61]), .B(A[61]), .Z(n3851) );
  NANDN U3615 ( .A(B[63]), .B(A[63]), .Z(n3843) );
  NANDN U3616 ( .A(B[65]), .B(A[65]), .Z(n3835) );
  NANDN U3617 ( .A(B[67]), .B(A[67]), .Z(n3827) );
  NANDN U3618 ( .A(B[69]), .B(A[69]), .Z(n3819) );
  NANDN U3619 ( .A(B[71]), .B(A[71]), .Z(n3811) );
  NANDN U3620 ( .A(B[73]), .B(A[73]), .Z(n3803) );
  NANDN U3621 ( .A(B[75]), .B(A[75]), .Z(n3795) );
  NANDN U3622 ( .A(B[77]), .B(A[77]), .Z(n3787) );
  NANDN U3623 ( .A(B[79]), .B(A[79]), .Z(n3779) );
  NANDN U3624 ( .A(B[81]), .B(A[81]), .Z(n3771) );
  NANDN U3625 ( .A(B[83]), .B(A[83]), .Z(n3763) );
  NANDN U3626 ( .A(B[85]), .B(A[85]), .Z(n3755) );
  NANDN U3627 ( .A(B[87]), .B(A[87]), .Z(n3747) );
  NANDN U3628 ( .A(B[89]), .B(A[89]), .Z(n3739) );
  NANDN U3629 ( .A(B[91]), .B(A[91]), .Z(n3731) );
  NANDN U3630 ( .A(B[93]), .B(A[93]), .Z(n3723) );
  NANDN U3631 ( .A(B[95]), .B(A[95]), .Z(n3715) );
  NANDN U3632 ( .A(B[97]), .B(A[97]), .Z(n3707) );
  NANDN U3633 ( .A(B[100]), .B(A[100]), .Z(n3699) );
  NANDN U3634 ( .A(B[101]), .B(A[101]), .Z(n3691) );
  NANDN U3635 ( .A(B[103]), .B(A[103]), .Z(n3683) );
  NANDN U3636 ( .A(B[105]), .B(A[105]), .Z(n3675) );
  NANDN U3637 ( .A(B[107]), .B(A[107]), .Z(n3667) );
  NANDN U3638 ( .A(B[109]), .B(A[109]), .Z(n3659) );
  NANDN U3639 ( .A(B[111]), .B(A[111]), .Z(n3651) );
  NANDN U3640 ( .A(B[113]), .B(A[113]), .Z(n3643) );
  NANDN U3641 ( .A(B[115]), .B(A[115]), .Z(n3635) );
  NANDN U3642 ( .A(B[117]), .B(A[117]), .Z(n3627) );
  NANDN U3643 ( .A(B[119]), .B(A[119]), .Z(n3619) );
  NANDN U3644 ( .A(B[121]), .B(A[121]), .Z(n3611) );
  NANDN U3645 ( .A(B[123]), .B(A[123]), .Z(n3603) );
  NANDN U3646 ( .A(B[125]), .B(A[125]), .Z(n3595) );
  NANDN U3647 ( .A(B[127]), .B(A[127]), .Z(n3587) );
  NANDN U3648 ( .A(B[129]), .B(A[129]), .Z(n3579) );
  NANDN U3649 ( .A(B[131]), .B(A[131]), .Z(n3571) );
  NANDN U3650 ( .A(B[133]), .B(A[133]), .Z(n3563) );
  NANDN U3651 ( .A(B[135]), .B(A[135]), .Z(n3555) );
  NANDN U3652 ( .A(B[137]), .B(A[137]), .Z(n3547) );
  NANDN U3653 ( .A(B[139]), .B(A[139]), .Z(n3539) );
  NANDN U3654 ( .A(B[141]), .B(A[141]), .Z(n3531) );
  NANDN U3655 ( .A(B[143]), .B(A[143]), .Z(n3523) );
  NANDN U3656 ( .A(B[145]), .B(A[145]), .Z(n3515) );
  NANDN U3657 ( .A(B[147]), .B(A[147]), .Z(n3507) );
  NANDN U3658 ( .A(B[149]), .B(A[149]), .Z(n3499) );
  NANDN U3659 ( .A(B[151]), .B(A[151]), .Z(n3491) );
  NANDN U3660 ( .A(B[153]), .B(A[153]), .Z(n3483) );
  NANDN U3661 ( .A(B[155]), .B(A[155]), .Z(n3475) );
  NANDN U3662 ( .A(B[157]), .B(A[157]), .Z(n3467) );
  NANDN U3663 ( .A(B[159]), .B(A[159]), .Z(n3459) );
  NANDN U3664 ( .A(B[161]), .B(A[161]), .Z(n3451) );
  NANDN U3665 ( .A(B[163]), .B(A[163]), .Z(n3443) );
  NANDN U3666 ( .A(B[165]), .B(A[165]), .Z(n3435) );
  NANDN U3667 ( .A(B[167]), .B(A[167]), .Z(n3427) );
  NANDN U3668 ( .A(B[169]), .B(A[169]), .Z(n3419) );
  NANDN U3669 ( .A(B[171]), .B(A[171]), .Z(n3411) );
  NANDN U3670 ( .A(B[173]), .B(A[173]), .Z(n3403) );
  NANDN U3671 ( .A(B[175]), .B(A[175]), .Z(n3395) );
  NANDN U3672 ( .A(B[177]), .B(A[177]), .Z(n3387) );
  NANDN U3673 ( .A(B[179]), .B(A[179]), .Z(n3379) );
  NANDN U3674 ( .A(B[181]), .B(A[181]), .Z(n3371) );
  NANDN U3675 ( .A(B[183]), .B(A[183]), .Z(n3363) );
  NANDN U3676 ( .A(B[185]), .B(A[185]), .Z(n3355) );
  NANDN U3677 ( .A(B[187]), .B(A[187]), .Z(n3347) );
  NANDN U3678 ( .A(B[189]), .B(A[189]), .Z(n3339) );
  NANDN U3679 ( .A(B[191]), .B(A[191]), .Z(n3331) );
  NANDN U3680 ( .A(B[193]), .B(A[193]), .Z(n3323) );
  NANDN U3681 ( .A(B[195]), .B(A[195]), .Z(n3315) );
  NANDN U3682 ( .A(B[197]), .B(A[197]), .Z(n3307) );
  NANDN U3683 ( .A(B[199]), .B(A[199]), .Z(n3299) );
  NANDN U3684 ( .A(B[201]), .B(A[201]), .Z(n3291) );
  NANDN U3685 ( .A(B[203]), .B(A[203]), .Z(n3283) );
  NANDN U3686 ( .A(B[205]), .B(A[205]), .Z(n3275) );
  NANDN U3687 ( .A(B[207]), .B(A[207]), .Z(n3267) );
  NANDN U3688 ( .A(B[209]), .B(A[209]), .Z(n3259) );
  NANDN U3689 ( .A(B[211]), .B(A[211]), .Z(n3251) );
  NANDN U3690 ( .A(B[213]), .B(A[213]), .Z(n3243) );
  NANDN U3691 ( .A(B[215]), .B(A[215]), .Z(n3235) );
  NANDN U3692 ( .A(B[217]), .B(A[217]), .Z(n3227) );
  NANDN U3693 ( .A(B[219]), .B(A[219]), .Z(n3219) );
  NANDN U3694 ( .A(B[221]), .B(A[221]), .Z(n3211) );
  NANDN U3695 ( .A(B[223]), .B(A[223]), .Z(n3203) );
  NANDN U3696 ( .A(B[225]), .B(A[225]), .Z(n3195) );
  NANDN U3697 ( .A(B[227]), .B(A[227]), .Z(n3187) );
  NANDN U3698 ( .A(B[229]), .B(A[229]), .Z(n3179) );
  NANDN U3699 ( .A(B[231]), .B(A[231]), .Z(n3171) );
  NANDN U3700 ( .A(B[233]), .B(A[233]), .Z(n3163) );
  NANDN U3701 ( .A(B[235]), .B(A[235]), .Z(n3155) );
  NANDN U3702 ( .A(B[237]), .B(A[237]), .Z(n3147) );
  NANDN U3703 ( .A(B[239]), .B(A[239]), .Z(n3139) );
  NANDN U3704 ( .A(B[241]), .B(A[241]), .Z(n3131) );
  NANDN U3705 ( .A(B[243]), .B(A[243]), .Z(n3123) );
  NANDN U3706 ( .A(B[245]), .B(A[245]), .Z(n3115) );
  NANDN U3707 ( .A(B[247]), .B(A[247]), .Z(n3107) );
  NANDN U3708 ( .A(B[249]), .B(A[249]), .Z(n3099) );
  NANDN U3709 ( .A(B[251]), .B(A[251]), .Z(n3091) );
  NANDN U3710 ( .A(B[253]), .B(A[253]), .Z(n3083) );
  NANDN U3711 ( .A(B[255]), .B(A[255]), .Z(n3075) );
  NANDN U3712 ( .A(B[257]), .B(A[257]), .Z(n3067) );
  NANDN U3713 ( .A(B[259]), .B(A[259]), .Z(n3059) );
  NANDN U3714 ( .A(B[261]), .B(A[261]), .Z(n3051) );
  NANDN U3715 ( .A(B[263]), .B(A[263]), .Z(n3043) );
  NANDN U3716 ( .A(B[265]), .B(A[265]), .Z(n3035) );
  NANDN U3717 ( .A(B[267]), .B(A[267]), .Z(n3027) );
  NANDN U3718 ( .A(B[269]), .B(A[269]), .Z(n3019) );
  NANDN U3719 ( .A(B[271]), .B(A[271]), .Z(n3011) );
  NANDN U3720 ( .A(B[273]), .B(A[273]), .Z(n3003) );
  NANDN U3721 ( .A(B[275]), .B(A[275]), .Z(n2995) );
  NANDN U3722 ( .A(B[277]), .B(A[277]), .Z(n2987) );
  NANDN U3723 ( .A(B[279]), .B(A[279]), .Z(n2979) );
  NANDN U3724 ( .A(B[281]), .B(A[281]), .Z(n2971) );
  NANDN U3725 ( .A(B[283]), .B(A[283]), .Z(n2963) );
  NANDN U3726 ( .A(B[285]), .B(A[285]), .Z(n2955) );
  NANDN U3727 ( .A(B[287]), .B(A[287]), .Z(n2947) );
  NANDN U3728 ( .A(B[289]), .B(A[289]), .Z(n2939) );
  NANDN U3729 ( .A(B[291]), .B(A[291]), .Z(n2931) );
  NANDN U3730 ( .A(B[293]), .B(A[293]), .Z(n2923) );
  NANDN U3731 ( .A(B[295]), .B(A[295]), .Z(n2915) );
  NANDN U3732 ( .A(B[297]), .B(A[297]), .Z(n2907) );
  NANDN U3733 ( .A(B[299]), .B(A[299]), .Z(n2899) );
  NANDN U3734 ( .A(B[301]), .B(A[301]), .Z(n2891) );
  NANDN U3735 ( .A(B[303]), .B(A[303]), .Z(n2883) );
  NANDN U3736 ( .A(B[305]), .B(A[305]), .Z(n2875) );
  NANDN U3737 ( .A(B[307]), .B(A[307]), .Z(n2867) );
  NANDN U3738 ( .A(B[309]), .B(A[309]), .Z(n2859) );
  NANDN U3739 ( .A(B[311]), .B(A[311]), .Z(n2851) );
  NANDN U3740 ( .A(B[313]), .B(A[313]), .Z(n2843) );
  NANDN U3741 ( .A(B[315]), .B(A[315]), .Z(n2835) );
  NANDN U3742 ( .A(B[317]), .B(A[317]), .Z(n2827) );
  NANDN U3743 ( .A(B[319]), .B(A[319]), .Z(n2819) );
  NANDN U3744 ( .A(B[321]), .B(A[321]), .Z(n2811) );
  NANDN U3745 ( .A(B[323]), .B(A[323]), .Z(n2803) );
  NANDN U3746 ( .A(B[325]), .B(A[325]), .Z(n2795) );
  NANDN U3747 ( .A(B[327]), .B(A[327]), .Z(n2787) );
  NANDN U3748 ( .A(B[329]), .B(A[329]), .Z(n2779) );
  NANDN U3749 ( .A(B[331]), .B(A[331]), .Z(n2771) );
  NANDN U3750 ( .A(B[333]), .B(A[333]), .Z(n2763) );
  NANDN U3751 ( .A(B[335]), .B(A[335]), .Z(n2755) );
  NANDN U3752 ( .A(B[337]), .B(A[337]), .Z(n2747) );
  NANDN U3753 ( .A(B[339]), .B(A[339]), .Z(n2739) );
  NANDN U3754 ( .A(B[341]), .B(A[341]), .Z(n2731) );
  NANDN U3755 ( .A(B[343]), .B(A[343]), .Z(n2723) );
  NANDN U3756 ( .A(B[345]), .B(A[345]), .Z(n2715) );
  NANDN U3757 ( .A(B[347]), .B(A[347]), .Z(n2707) );
  NANDN U3758 ( .A(B[349]), .B(A[349]), .Z(n2699) );
  NANDN U3759 ( .A(B[351]), .B(A[351]), .Z(n2691) );
  NANDN U3760 ( .A(B[353]), .B(A[353]), .Z(n2683) );
  NANDN U3761 ( .A(B[355]), .B(A[355]), .Z(n2675) );
  NANDN U3762 ( .A(B[357]), .B(A[357]), .Z(n2667) );
  NANDN U3763 ( .A(B[359]), .B(A[359]), .Z(n2659) );
  NANDN U3764 ( .A(B[361]), .B(A[361]), .Z(n2651) );
  NANDN U3765 ( .A(B[363]), .B(A[363]), .Z(n2643) );
  NANDN U3766 ( .A(B[365]), .B(A[365]), .Z(n2635) );
  NANDN U3767 ( .A(B[367]), .B(A[367]), .Z(n2627) );
  NANDN U3768 ( .A(B[369]), .B(A[369]), .Z(n2619) );
  NANDN U3769 ( .A(B[371]), .B(A[371]), .Z(n2611) );
  NANDN U3770 ( .A(B[373]), .B(A[373]), .Z(n2603) );
  NANDN U3771 ( .A(B[375]), .B(A[375]), .Z(n2595) );
  NANDN U3772 ( .A(B[377]), .B(A[377]), .Z(n2587) );
  NANDN U3773 ( .A(B[379]), .B(A[379]), .Z(n2579) );
  NANDN U3774 ( .A(B[381]), .B(A[381]), .Z(n2571) );
  NANDN U3775 ( .A(B[383]), .B(A[383]), .Z(n2563) );
  NANDN U3776 ( .A(B[385]), .B(A[385]), .Z(n2555) );
  NANDN U3777 ( .A(B[387]), .B(A[387]), .Z(n2547) );
  NANDN U3778 ( .A(B[389]), .B(A[389]), .Z(n2539) );
  NANDN U3779 ( .A(B[391]), .B(A[391]), .Z(n2531) );
  NANDN U3780 ( .A(B[393]), .B(A[393]), .Z(n2523) );
  NANDN U3781 ( .A(B[395]), .B(A[395]), .Z(n2515) );
  NANDN U3782 ( .A(B[397]), .B(A[397]), .Z(n2507) );
  NANDN U3783 ( .A(B[399]), .B(A[399]), .Z(n2499) );
  NANDN U3784 ( .A(B[401]), .B(A[401]), .Z(n2491) );
  NANDN U3785 ( .A(B[403]), .B(A[403]), .Z(n2483) );
  NANDN U3786 ( .A(B[405]), .B(A[405]), .Z(n2475) );
  NANDN U3787 ( .A(B[407]), .B(A[407]), .Z(n2467) );
  NANDN U3788 ( .A(B[409]), .B(A[409]), .Z(n2459) );
  NANDN U3789 ( .A(B[411]), .B(A[411]), .Z(n2451) );
  NANDN U3790 ( .A(B[413]), .B(A[413]), .Z(n2443) );
  NANDN U3791 ( .A(B[415]), .B(A[415]), .Z(n2435) );
  NANDN U3792 ( .A(B[417]), .B(A[417]), .Z(n2427) );
  NANDN U3793 ( .A(B[419]), .B(A[419]), .Z(n2419) );
  NANDN U3794 ( .A(B[421]), .B(A[421]), .Z(n2411) );
  NANDN U3795 ( .A(B[423]), .B(A[423]), .Z(n2403) );
  NANDN U3796 ( .A(B[425]), .B(A[425]), .Z(n2395) );
  NANDN U3797 ( .A(B[427]), .B(A[427]), .Z(n2387) );
  NANDN U3798 ( .A(B[429]), .B(A[429]), .Z(n2379) );
  NANDN U3799 ( .A(B[431]), .B(A[431]), .Z(n2371) );
  NANDN U3800 ( .A(B[433]), .B(A[433]), .Z(n2363) );
  NANDN U3801 ( .A(B[435]), .B(A[435]), .Z(n2355) );
  NANDN U3802 ( .A(B[437]), .B(A[437]), .Z(n2347) );
  NANDN U3803 ( .A(B[439]), .B(A[439]), .Z(n2339) );
  NANDN U3804 ( .A(B[441]), .B(A[441]), .Z(n2331) );
  NANDN U3805 ( .A(B[443]), .B(A[443]), .Z(n2323) );
  NANDN U3806 ( .A(B[445]), .B(A[445]), .Z(n2315) );
  NANDN U3807 ( .A(B[447]), .B(A[447]), .Z(n2307) );
  NANDN U3808 ( .A(B[449]), .B(A[449]), .Z(n2299) );
  NANDN U3809 ( .A(B[451]), .B(A[451]), .Z(n2291) );
  NANDN U3810 ( .A(B[453]), .B(A[453]), .Z(n2283) );
  NANDN U3811 ( .A(B[455]), .B(A[455]), .Z(n2275) );
  NANDN U3812 ( .A(B[457]), .B(A[457]), .Z(n2267) );
  NANDN U3813 ( .A(B[459]), .B(A[459]), .Z(n2259) );
  NANDN U3814 ( .A(B[461]), .B(A[461]), .Z(n2251) );
  NANDN U3815 ( .A(B[463]), .B(A[463]), .Z(n2243) );
  NANDN U3816 ( .A(B[465]), .B(A[465]), .Z(n2235) );
  NANDN U3817 ( .A(B[467]), .B(A[467]), .Z(n2227) );
  NANDN U3818 ( .A(B[469]), .B(A[469]), .Z(n2219) );
  NANDN U3819 ( .A(B[471]), .B(A[471]), .Z(n2211) );
  NANDN U3820 ( .A(B[473]), .B(A[473]), .Z(n2203) );
  NANDN U3821 ( .A(B[475]), .B(A[475]), .Z(n2195) );
  NANDN U3822 ( .A(B[477]), .B(A[477]), .Z(n2187) );
  NANDN U3823 ( .A(B[479]), .B(A[479]), .Z(n2179) );
  NANDN U3824 ( .A(B[481]), .B(A[481]), .Z(n2171) );
  NANDN U3825 ( .A(B[483]), .B(A[483]), .Z(n2163) );
  NANDN U3826 ( .A(B[485]), .B(A[485]), .Z(n2155) );
  NANDN U3827 ( .A(B[487]), .B(A[487]), .Z(n2147) );
  NANDN U3828 ( .A(B[489]), .B(A[489]), .Z(n2139) );
  NANDN U3829 ( .A(B[491]), .B(A[491]), .Z(n2131) );
  NANDN U3830 ( .A(B[493]), .B(A[493]), .Z(n2123) );
  NANDN U3831 ( .A(B[495]), .B(A[495]), .Z(n2115) );
  NANDN U3832 ( .A(B[497]), .B(A[497]), .Z(n2107) );
  NANDN U3833 ( .A(B[499]), .B(A[499]), .Z(n2099) );
  NANDN U3834 ( .A(B[501]), .B(A[501]), .Z(n2091) );
  NANDN U3835 ( .A(B[503]), .B(A[503]), .Z(n2083) );
  NANDN U3836 ( .A(B[505]), .B(A[505]), .Z(n2075) );
  NANDN U3837 ( .A(B[507]), .B(A[507]), .Z(n2067) );
  NANDN U3838 ( .A(B[509]), .B(A[509]), .Z(n2059) );
  NANDN U3839 ( .A(B[511]), .B(A[511]), .Z(n2051) );
  NANDN U3840 ( .A(B[513]), .B(A[513]), .Z(n2043) );
  NANDN U3841 ( .A(B[515]), .B(A[515]), .Z(n2035) );
  NANDN U3842 ( .A(B[517]), .B(A[517]), .Z(n2027) );
  NANDN U3843 ( .A(B[519]), .B(A[519]), .Z(n2019) );
  NANDN U3844 ( .A(B[521]), .B(A[521]), .Z(n2011) );
  NANDN U3845 ( .A(B[523]), .B(A[523]), .Z(n2003) );
  NANDN U3846 ( .A(B[525]), .B(A[525]), .Z(n1995) );
  NANDN U3847 ( .A(B[527]), .B(A[527]), .Z(n1987) );
  NANDN U3848 ( .A(B[529]), .B(A[529]), .Z(n1979) );
  NANDN U3849 ( .A(B[531]), .B(A[531]), .Z(n1971) );
  NANDN U3850 ( .A(B[533]), .B(A[533]), .Z(n1963) );
  NANDN U3851 ( .A(B[535]), .B(A[535]), .Z(n1955) );
  NANDN U3852 ( .A(B[537]), .B(A[537]), .Z(n1947) );
  NANDN U3853 ( .A(B[539]), .B(A[539]), .Z(n1939) );
  NANDN U3854 ( .A(B[541]), .B(A[541]), .Z(n1931) );
  NANDN U3855 ( .A(B[543]), .B(A[543]), .Z(n1923) );
  NANDN U3856 ( .A(B[545]), .B(A[545]), .Z(n1915) );
  NANDN U3857 ( .A(B[547]), .B(A[547]), .Z(n1907) );
  NANDN U3858 ( .A(B[549]), .B(A[549]), .Z(n1899) );
  NANDN U3859 ( .A(B[551]), .B(A[551]), .Z(n1891) );
  NANDN U3860 ( .A(B[553]), .B(A[553]), .Z(n1883) );
  NANDN U3861 ( .A(B[555]), .B(A[555]), .Z(n1875) );
  NANDN U3862 ( .A(B[557]), .B(A[557]), .Z(n1867) );
  NANDN U3863 ( .A(B[559]), .B(A[559]), .Z(n1859) );
  NANDN U3864 ( .A(B[561]), .B(A[561]), .Z(n1851) );
  NANDN U3865 ( .A(B[563]), .B(A[563]), .Z(n1843) );
  NANDN U3866 ( .A(B[565]), .B(A[565]), .Z(n1835) );
  NANDN U3867 ( .A(B[567]), .B(A[567]), .Z(n1827) );
  NANDN U3868 ( .A(B[569]), .B(A[569]), .Z(n1819) );
  NANDN U3869 ( .A(B[571]), .B(A[571]), .Z(n1811) );
  NANDN U3870 ( .A(B[573]), .B(A[573]), .Z(n1803) );
  NANDN U3871 ( .A(B[575]), .B(A[575]), .Z(n1795) );
  NANDN U3872 ( .A(B[577]), .B(A[577]), .Z(n1787) );
  NANDN U3873 ( .A(B[579]), .B(A[579]), .Z(n1779) );
  NANDN U3874 ( .A(B[581]), .B(A[581]), .Z(n1771) );
  NANDN U3875 ( .A(B[583]), .B(A[583]), .Z(n1763) );
  NANDN U3876 ( .A(B[585]), .B(A[585]), .Z(n1755) );
  NANDN U3877 ( .A(B[587]), .B(A[587]), .Z(n1747) );
  NANDN U3878 ( .A(B[589]), .B(A[589]), .Z(n1739) );
  NANDN U3879 ( .A(B[591]), .B(A[591]), .Z(n1731) );
  NANDN U3880 ( .A(B[593]), .B(A[593]), .Z(n1723) );
  NANDN U3881 ( .A(B[595]), .B(A[595]), .Z(n1715) );
  NANDN U3882 ( .A(B[597]), .B(A[597]), .Z(n1707) );
  NANDN U3883 ( .A(B[599]), .B(A[599]), .Z(n1699) );
  NANDN U3884 ( .A(B[601]), .B(A[601]), .Z(n1691) );
  NANDN U3885 ( .A(B[603]), .B(A[603]), .Z(n1683) );
  NANDN U3886 ( .A(B[605]), .B(A[605]), .Z(n1675) );
  NANDN U3887 ( .A(B[607]), .B(A[607]), .Z(n1667) );
  NANDN U3888 ( .A(B[609]), .B(A[609]), .Z(n1659) );
  NANDN U3889 ( .A(B[611]), .B(A[611]), .Z(n1651) );
  NANDN U3890 ( .A(B[613]), .B(A[613]), .Z(n1643) );
  NANDN U3891 ( .A(B[615]), .B(A[615]), .Z(n1635) );
  NANDN U3892 ( .A(B[617]), .B(A[617]), .Z(n1627) );
  NANDN U3893 ( .A(B[619]), .B(A[619]), .Z(n1619) );
  NANDN U3894 ( .A(B[621]), .B(A[621]), .Z(n1611) );
  NANDN U3895 ( .A(B[623]), .B(A[623]), .Z(n1603) );
  NANDN U3896 ( .A(B[625]), .B(A[625]), .Z(n1595) );
  NANDN U3897 ( .A(B[627]), .B(A[627]), .Z(n1587) );
  NANDN U3898 ( .A(B[629]), .B(A[629]), .Z(n1579) );
  NANDN U3899 ( .A(B[631]), .B(A[631]), .Z(n1571) );
  NANDN U3900 ( .A(B[633]), .B(A[633]), .Z(n1563) );
  NANDN U3901 ( .A(B[635]), .B(A[635]), .Z(n1555) );
  NANDN U3902 ( .A(B[637]), .B(A[637]), .Z(n1547) );
  NANDN U3903 ( .A(B[639]), .B(A[639]), .Z(n1539) );
  NANDN U3904 ( .A(B[641]), .B(A[641]), .Z(n1531) );
  NANDN U3905 ( .A(B[643]), .B(A[643]), .Z(n1523) );
  NANDN U3906 ( .A(B[645]), .B(A[645]), .Z(n1515) );
  NANDN U3907 ( .A(B[647]), .B(A[647]), .Z(n1507) );
  NANDN U3908 ( .A(B[649]), .B(A[649]), .Z(n1499) );
  NANDN U3909 ( .A(B[651]), .B(A[651]), .Z(n1491) );
  NANDN U3910 ( .A(B[653]), .B(A[653]), .Z(n1483) );
  NANDN U3911 ( .A(B[655]), .B(A[655]), .Z(n1475) );
  NANDN U3912 ( .A(B[657]), .B(A[657]), .Z(n1467) );
  NANDN U3913 ( .A(B[659]), .B(A[659]), .Z(n1459) );
  NANDN U3914 ( .A(B[661]), .B(A[661]), .Z(n1451) );
  NANDN U3915 ( .A(B[663]), .B(A[663]), .Z(n1443) );
  NANDN U3916 ( .A(B[665]), .B(A[665]), .Z(n1435) );
  NANDN U3917 ( .A(B[667]), .B(A[667]), .Z(n1427) );
  NANDN U3918 ( .A(B[669]), .B(A[669]), .Z(n1419) );
  NANDN U3919 ( .A(B[671]), .B(A[671]), .Z(n1411) );
  NANDN U3920 ( .A(B[673]), .B(A[673]), .Z(n1403) );
  NANDN U3921 ( .A(B[675]), .B(A[675]), .Z(n1395) );
  NANDN U3922 ( .A(B[677]), .B(A[677]), .Z(n1387) );
  NANDN U3923 ( .A(B[679]), .B(A[679]), .Z(n1379) );
  NANDN U3924 ( .A(B[681]), .B(A[681]), .Z(n1371) );
  NANDN U3925 ( .A(B[683]), .B(A[683]), .Z(n1363) );
  NANDN U3926 ( .A(B[685]), .B(A[685]), .Z(n1355) );
  NANDN U3927 ( .A(B[687]), .B(A[687]), .Z(n1347) );
  NANDN U3928 ( .A(B[689]), .B(A[689]), .Z(n1339) );
  NANDN U3929 ( .A(B[691]), .B(A[691]), .Z(n1331) );
  NANDN U3930 ( .A(B[693]), .B(A[693]), .Z(n1323) );
  NANDN U3931 ( .A(B[695]), .B(A[695]), .Z(n1315) );
  NANDN U3932 ( .A(B[697]), .B(A[697]), .Z(n1307) );
  NANDN U3933 ( .A(B[699]), .B(A[699]), .Z(n1299) );
  NANDN U3934 ( .A(B[701]), .B(A[701]), .Z(n1291) );
  NANDN U3935 ( .A(B[703]), .B(A[703]), .Z(n1283) );
  NANDN U3936 ( .A(B[705]), .B(A[705]), .Z(n1275) );
  NANDN U3937 ( .A(B[707]), .B(A[707]), .Z(n1267) );
  NANDN U3938 ( .A(B[709]), .B(A[709]), .Z(n1259) );
  NANDN U3939 ( .A(B[711]), .B(A[711]), .Z(n1251) );
  NANDN U3940 ( .A(B[713]), .B(A[713]), .Z(n1243) );
  NANDN U3941 ( .A(B[715]), .B(A[715]), .Z(n1235) );
  NANDN U3942 ( .A(B[717]), .B(A[717]), .Z(n1227) );
  NANDN U3943 ( .A(B[719]), .B(A[719]), .Z(n1219) );
  NANDN U3944 ( .A(B[721]), .B(A[721]), .Z(n1211) );
  NANDN U3945 ( .A(B[723]), .B(A[723]), .Z(n1203) );
  NANDN U3946 ( .A(B[725]), .B(A[725]), .Z(n1195) );
  NANDN U3947 ( .A(B[727]), .B(A[727]), .Z(n1187) );
  NANDN U3948 ( .A(B[729]), .B(A[729]), .Z(n1179) );
  NANDN U3949 ( .A(B[731]), .B(A[731]), .Z(n1171) );
  NANDN U3950 ( .A(B[733]), .B(A[733]), .Z(n1163) );
  NANDN U3951 ( .A(B[735]), .B(A[735]), .Z(n1155) );
  NANDN U3952 ( .A(B[737]), .B(A[737]), .Z(n1147) );
  NANDN U3953 ( .A(B[739]), .B(A[739]), .Z(n1139) );
  NANDN U3954 ( .A(B[741]), .B(A[741]), .Z(n1131) );
  NANDN U3955 ( .A(B[743]), .B(A[743]), .Z(n1123) );
  NANDN U3956 ( .A(B[745]), .B(A[745]), .Z(n1115) );
  NANDN U3957 ( .A(B[747]), .B(A[747]), .Z(n1107) );
  NANDN U3958 ( .A(B[749]), .B(A[749]), .Z(n1099) );
  NANDN U3959 ( .A(B[751]), .B(A[751]), .Z(n1091) );
  NANDN U3960 ( .A(B[753]), .B(A[753]), .Z(n1083) );
  NANDN U3961 ( .A(B[755]), .B(A[755]), .Z(n1075) );
  NANDN U3962 ( .A(B[757]), .B(A[757]), .Z(n1067) );
  NANDN U3963 ( .A(B[759]), .B(A[759]), .Z(n1059) );
  NANDN U3964 ( .A(B[761]), .B(A[761]), .Z(n1051) );
  NANDN U3965 ( .A(B[763]), .B(A[763]), .Z(n1043) );
  NANDN U3966 ( .A(B[765]), .B(A[765]), .Z(n1035) );
  NANDN U3967 ( .A(B[767]), .B(A[767]), .Z(n1027) );
  NANDN U3968 ( .A(B[769]), .B(A[769]), .Z(n1019) );
  NANDN U3969 ( .A(B[771]), .B(A[771]), .Z(n1011) );
  NANDN U3970 ( .A(B[773]), .B(A[773]), .Z(n1003) );
  NANDN U3971 ( .A(B[775]), .B(A[775]), .Z(n995) );
  NANDN U3972 ( .A(B[777]), .B(A[777]), .Z(n987) );
  NANDN U3973 ( .A(B[779]), .B(A[779]), .Z(n979) );
  NANDN U3974 ( .A(B[781]), .B(A[781]), .Z(n971) );
  NANDN U3975 ( .A(B[783]), .B(A[783]), .Z(n963) );
  NANDN U3976 ( .A(B[785]), .B(A[785]), .Z(n955) );
  NANDN U3977 ( .A(B[787]), .B(A[787]), .Z(n947) );
  NANDN U3978 ( .A(B[789]), .B(A[789]), .Z(n939) );
  NANDN U3979 ( .A(B[791]), .B(A[791]), .Z(n931) );
  NANDN U3980 ( .A(B[793]), .B(A[793]), .Z(n923) );
  NANDN U3981 ( .A(B[795]), .B(A[795]), .Z(n915) );
  NANDN U3982 ( .A(B[797]), .B(A[797]), .Z(n907) );
  NANDN U3983 ( .A(B[799]), .B(A[799]), .Z(n899) );
  NANDN U3984 ( .A(B[801]), .B(A[801]), .Z(n891) );
  NANDN U3985 ( .A(B[803]), .B(A[803]), .Z(n883) );
  NANDN U3986 ( .A(B[805]), .B(A[805]), .Z(n875) );
  NANDN U3987 ( .A(B[807]), .B(A[807]), .Z(n867) );
  NANDN U3988 ( .A(B[809]), .B(A[809]), .Z(n859) );
  NANDN U3989 ( .A(B[811]), .B(A[811]), .Z(n851) );
  NANDN U3990 ( .A(B[813]), .B(A[813]), .Z(n843) );
  NANDN U3991 ( .A(B[815]), .B(A[815]), .Z(n835) );
  NANDN U3992 ( .A(B[817]), .B(A[817]), .Z(n827) );
  NANDN U3993 ( .A(B[819]), .B(A[819]), .Z(n819) );
  NANDN U3994 ( .A(B[821]), .B(A[821]), .Z(n811) );
  NANDN U3995 ( .A(B[823]), .B(A[823]), .Z(n803) );
  NANDN U3996 ( .A(B[825]), .B(A[825]), .Z(n795) );
  NANDN U3997 ( .A(B[827]), .B(A[827]), .Z(n787) );
  NANDN U3998 ( .A(B[829]), .B(A[829]), .Z(n779) );
  NANDN U3999 ( .A(B[831]), .B(A[831]), .Z(n771) );
  NANDN U4000 ( .A(B[833]), .B(A[833]), .Z(n763) );
  NANDN U4001 ( .A(B[835]), .B(A[835]), .Z(n755) );
  NANDN U4002 ( .A(B[837]), .B(A[837]), .Z(n747) );
  NANDN U4003 ( .A(B[839]), .B(A[839]), .Z(n739) );
  NANDN U4004 ( .A(B[841]), .B(A[841]), .Z(n731) );
  NANDN U4005 ( .A(B[843]), .B(A[843]), .Z(n723) );
  NANDN U4006 ( .A(B[845]), .B(A[845]), .Z(n715) );
  NANDN U4007 ( .A(B[847]), .B(A[847]), .Z(n707) );
  NANDN U4008 ( .A(B[849]), .B(A[849]), .Z(n699) );
  NANDN U4009 ( .A(B[851]), .B(A[851]), .Z(n691) );
  NANDN U4010 ( .A(B[853]), .B(A[853]), .Z(n683) );
  NANDN U4011 ( .A(B[855]), .B(A[855]), .Z(n675) );
  NANDN U4012 ( .A(B[857]), .B(A[857]), .Z(n667) );
  NANDN U4013 ( .A(B[859]), .B(A[859]), .Z(n659) );
  NANDN U4014 ( .A(B[861]), .B(A[861]), .Z(n651) );
  NANDN U4015 ( .A(B[863]), .B(A[863]), .Z(n643) );
  NANDN U4016 ( .A(B[865]), .B(A[865]), .Z(n635) );
  NANDN U4017 ( .A(B[867]), .B(A[867]), .Z(n627) );
  NANDN U4018 ( .A(B[869]), .B(A[869]), .Z(n619) );
  NANDN U4019 ( .A(B[871]), .B(A[871]), .Z(n611) );
  NANDN U4020 ( .A(B[873]), .B(A[873]), .Z(n603) );
  NANDN U4021 ( .A(B[875]), .B(A[875]), .Z(n595) );
  NANDN U4022 ( .A(B[877]), .B(A[877]), .Z(n587) );
  NANDN U4023 ( .A(B[879]), .B(A[879]), .Z(n579) );
  NANDN U4024 ( .A(B[881]), .B(A[881]), .Z(n571) );
  NANDN U4025 ( .A(B[883]), .B(A[883]), .Z(n563) );
  NANDN U4026 ( .A(B[885]), .B(A[885]), .Z(n555) );
  NANDN U4027 ( .A(B[887]), .B(A[887]), .Z(n547) );
  NANDN U4028 ( .A(B[889]), .B(A[889]), .Z(n539) );
  NANDN U4029 ( .A(B[891]), .B(A[891]), .Z(n531) );
  NANDN U4030 ( .A(B[893]), .B(A[893]), .Z(n523) );
  NANDN U4031 ( .A(B[895]), .B(A[895]), .Z(n515) );
  NANDN U4032 ( .A(B[897]), .B(A[897]), .Z(n507) );
  NANDN U4033 ( .A(B[899]), .B(A[899]), .Z(n499) );
  NANDN U4034 ( .A(B[901]), .B(A[901]), .Z(n491) );
  NANDN U4035 ( .A(B[903]), .B(A[903]), .Z(n483) );
  NANDN U4036 ( .A(B[905]), .B(A[905]), .Z(n475) );
  NANDN U4037 ( .A(B[907]), .B(A[907]), .Z(n467) );
  NANDN U4038 ( .A(B[909]), .B(A[909]), .Z(n459) );
  NANDN U4039 ( .A(B[911]), .B(A[911]), .Z(n451) );
  NANDN U4040 ( .A(B[913]), .B(A[913]), .Z(n443) );
  NANDN U4041 ( .A(B[915]), .B(A[915]), .Z(n435) );
  NANDN U4042 ( .A(B[917]), .B(A[917]), .Z(n427) );
  NANDN U4043 ( .A(B[919]), .B(A[919]), .Z(n419) );
  NANDN U4044 ( .A(B[921]), .B(A[921]), .Z(n411) );
  NANDN U4045 ( .A(B[923]), .B(A[923]), .Z(n403) );
  NANDN U4046 ( .A(B[925]), .B(A[925]), .Z(n395) );
  NANDN U4047 ( .A(B[927]), .B(A[927]), .Z(n387) );
  NANDN U4048 ( .A(B[929]), .B(A[929]), .Z(n379) );
  NANDN U4049 ( .A(B[931]), .B(A[931]), .Z(n371) );
  NANDN U4050 ( .A(B[933]), .B(A[933]), .Z(n363) );
  NANDN U4051 ( .A(B[935]), .B(A[935]), .Z(n355) );
  NANDN U4052 ( .A(B[937]), .B(A[937]), .Z(n347) );
  NANDN U4053 ( .A(B[939]), .B(A[939]), .Z(n339) );
  NANDN U4054 ( .A(B[941]), .B(A[941]), .Z(n331) );
  NANDN U4055 ( .A(B[943]), .B(A[943]), .Z(n323) );
  NANDN U4056 ( .A(B[945]), .B(A[945]), .Z(n315) );
  NANDN U4057 ( .A(B[947]), .B(A[947]), .Z(n307) );
  NANDN U4058 ( .A(B[949]), .B(A[949]), .Z(n299) );
  NANDN U4059 ( .A(B[951]), .B(A[951]), .Z(n291) );
  NANDN U4060 ( .A(B[953]), .B(A[953]), .Z(n283) );
  NANDN U4061 ( .A(B[955]), .B(A[955]), .Z(n275) );
  NANDN U4062 ( .A(B[957]), .B(A[957]), .Z(n267) );
  NANDN U4063 ( .A(B[959]), .B(A[959]), .Z(n259) );
  NANDN U4064 ( .A(B[961]), .B(A[961]), .Z(n251) );
  NANDN U4065 ( .A(B[963]), .B(A[963]), .Z(n243) );
  NANDN U4066 ( .A(B[965]), .B(A[965]), .Z(n235) );
  NANDN U4067 ( .A(B[967]), .B(A[967]), .Z(n227) );
  NANDN U4068 ( .A(B[969]), .B(A[969]), .Z(n219) );
  NANDN U4069 ( .A(B[971]), .B(A[971]), .Z(n211) );
  NANDN U4070 ( .A(B[973]), .B(A[973]), .Z(n203) );
  NANDN U4071 ( .A(B[975]), .B(A[975]), .Z(n195) );
  NANDN U4072 ( .A(B[977]), .B(A[977]), .Z(n187) );
  NANDN U4073 ( .A(B[979]), .B(A[979]), .Z(n179) );
  NANDN U4074 ( .A(B[981]), .B(A[981]), .Z(n171) );
  NANDN U4075 ( .A(B[983]), .B(A[983]), .Z(n163) );
  NANDN U4076 ( .A(B[985]), .B(A[985]), .Z(n155) );
  NANDN U4077 ( .A(B[987]), .B(A[987]), .Z(n147) );
  NANDN U4078 ( .A(B[989]), .B(A[989]), .Z(n139) );
  NANDN U4079 ( .A(B[991]), .B(A[991]), .Z(n131) );
  NANDN U4080 ( .A(B[993]), .B(A[993]), .Z(n123) );
  NANDN U4081 ( .A(B[995]), .B(A[995]), .Z(n115) );
  NANDN U4082 ( .A(B[997]), .B(A[997]), .Z(n107) );
  NANDN U4083 ( .A(B[1000]), .B(A[1000]), .Z(n99) );
  NANDN U4084 ( .A(B[1001]), .B(A[1001]), .Z(n91) );
  NANDN U4085 ( .A(B[1003]), .B(A[1003]), .Z(n83) );
  NANDN U4086 ( .A(B[1005]), .B(A[1005]), .Z(n75) );
  NANDN U4087 ( .A(B[1007]), .B(A[1007]), .Z(n67) );
  NANDN U4088 ( .A(B[1009]), .B(A[1009]), .Z(n59) );
  NANDN U4089 ( .A(B[1011]), .B(A[1011]), .Z(n51) );
  NANDN U4090 ( .A(B[1013]), .B(A[1013]), .Z(n43) );
  NANDN U4091 ( .A(B[1015]), .B(A[1015]), .Z(n35) );
  NANDN U4092 ( .A(B[1017]), .B(A[1017]), .Z(n27) );
  NANDN U4093 ( .A(B[1019]), .B(A[1019]), .Z(n19) );
  NANDN U4094 ( .A(B[1021]), .B(A[1021]), .Z(n11) );
  NANDN U4095 ( .A(A[1023]), .B(B[1023]), .Z(n3) );
endmodule


module modmult_step_N1024_DW01_add_0 ( A, B, CI, SUM, CO );
  input [1025:0] A;
  input [1025:0] B;
  output [1025:0] SUM;
  input CI;
  output CO;
  wire   \B[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
         n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
         n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
         n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
         n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
         n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
         n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
         n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
         n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
         n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
         n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
         n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112;
  assign SUM[0] = \B[0] ;
  assign \B[0]  = B[0];

  XNOR U1 ( .A(n1), .B(n2), .Z(SUM[9]) );
  XNOR U2 ( .A(B[9]), .B(A[9]), .Z(n2) );
  XNOR U3 ( .A(n3), .B(n4), .Z(SUM[99]) );
  XNOR U4 ( .A(B[99]), .B(A[99]), .Z(n4) );
  XNOR U5 ( .A(n5), .B(n6), .Z(SUM[999]) );
  XNOR U6 ( .A(B[999]), .B(A[999]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[998]) );
  XNOR U8 ( .A(B[998]), .B(A[998]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[997]) );
  XNOR U10 ( .A(B[997]), .B(A[997]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[996]) );
  XNOR U12 ( .A(B[996]), .B(A[996]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[995]) );
  XNOR U14 ( .A(B[995]), .B(A[995]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(SUM[994]) );
  XNOR U16 ( .A(B[994]), .B(A[994]), .Z(n16) );
  XOR U17 ( .A(n17), .B(n18), .Z(SUM[993]) );
  XNOR U18 ( .A(B[993]), .B(A[993]), .Z(n18) );
  XOR U19 ( .A(n19), .B(n20), .Z(SUM[992]) );
  XNOR U20 ( .A(B[992]), .B(A[992]), .Z(n20) );
  XOR U21 ( .A(n21), .B(n22), .Z(SUM[991]) );
  XNOR U22 ( .A(B[991]), .B(A[991]), .Z(n22) );
  XOR U23 ( .A(n23), .B(n24), .Z(SUM[990]) );
  XNOR U24 ( .A(B[990]), .B(A[990]), .Z(n24) );
  XOR U25 ( .A(n25), .B(n26), .Z(SUM[98]) );
  XNOR U26 ( .A(B[98]), .B(A[98]), .Z(n26) );
  XOR U27 ( .A(n27), .B(n28), .Z(SUM[989]) );
  XNOR U28 ( .A(B[989]), .B(A[989]), .Z(n28) );
  XOR U29 ( .A(n29), .B(n30), .Z(SUM[988]) );
  XNOR U30 ( .A(B[988]), .B(A[988]), .Z(n30) );
  XOR U31 ( .A(n31), .B(n32), .Z(SUM[987]) );
  XNOR U32 ( .A(B[987]), .B(A[987]), .Z(n32) );
  XOR U33 ( .A(n33), .B(n34), .Z(SUM[986]) );
  XNOR U34 ( .A(B[986]), .B(A[986]), .Z(n34) );
  XOR U35 ( .A(n35), .B(n36), .Z(SUM[985]) );
  XNOR U36 ( .A(B[985]), .B(A[985]), .Z(n36) );
  XOR U37 ( .A(n37), .B(n38), .Z(SUM[984]) );
  XNOR U38 ( .A(B[984]), .B(A[984]), .Z(n38) );
  XOR U39 ( .A(n39), .B(n40), .Z(SUM[983]) );
  XNOR U40 ( .A(B[983]), .B(A[983]), .Z(n40) );
  XOR U41 ( .A(n41), .B(n42), .Z(SUM[982]) );
  XNOR U42 ( .A(B[982]), .B(A[982]), .Z(n42) );
  XOR U43 ( .A(n43), .B(n44), .Z(SUM[981]) );
  XNOR U44 ( .A(B[981]), .B(A[981]), .Z(n44) );
  XOR U45 ( .A(n45), .B(n46), .Z(SUM[980]) );
  XNOR U46 ( .A(B[980]), .B(A[980]), .Z(n46) );
  XOR U47 ( .A(n47), .B(n48), .Z(SUM[97]) );
  XNOR U48 ( .A(B[97]), .B(A[97]), .Z(n48) );
  XOR U49 ( .A(n49), .B(n50), .Z(SUM[979]) );
  XNOR U50 ( .A(B[979]), .B(A[979]), .Z(n50) );
  XOR U51 ( .A(n51), .B(n52), .Z(SUM[978]) );
  XNOR U52 ( .A(B[978]), .B(A[978]), .Z(n52) );
  XOR U53 ( .A(n53), .B(n54), .Z(SUM[977]) );
  XNOR U54 ( .A(B[977]), .B(A[977]), .Z(n54) );
  XOR U55 ( .A(n55), .B(n56), .Z(SUM[976]) );
  XNOR U56 ( .A(B[976]), .B(A[976]), .Z(n56) );
  XOR U57 ( .A(n57), .B(n58), .Z(SUM[975]) );
  XNOR U58 ( .A(B[975]), .B(A[975]), .Z(n58) );
  XOR U59 ( .A(n59), .B(n60), .Z(SUM[974]) );
  XNOR U60 ( .A(B[974]), .B(A[974]), .Z(n60) );
  XOR U61 ( .A(n61), .B(n62), .Z(SUM[973]) );
  XNOR U62 ( .A(B[973]), .B(A[973]), .Z(n62) );
  XOR U63 ( .A(n63), .B(n64), .Z(SUM[972]) );
  XNOR U64 ( .A(B[972]), .B(A[972]), .Z(n64) );
  XOR U65 ( .A(n65), .B(n66), .Z(SUM[971]) );
  XNOR U66 ( .A(B[971]), .B(A[971]), .Z(n66) );
  XOR U67 ( .A(n67), .B(n68), .Z(SUM[970]) );
  XNOR U68 ( .A(B[970]), .B(A[970]), .Z(n68) );
  XOR U69 ( .A(n69), .B(n70), .Z(SUM[96]) );
  XNOR U70 ( .A(B[96]), .B(A[96]), .Z(n70) );
  XOR U71 ( .A(n71), .B(n72), .Z(SUM[969]) );
  XNOR U72 ( .A(B[969]), .B(A[969]), .Z(n72) );
  XOR U73 ( .A(n73), .B(n74), .Z(SUM[968]) );
  XNOR U74 ( .A(B[968]), .B(A[968]), .Z(n74) );
  XOR U75 ( .A(n75), .B(n76), .Z(SUM[967]) );
  XNOR U76 ( .A(B[967]), .B(A[967]), .Z(n76) );
  XOR U77 ( .A(n77), .B(n78), .Z(SUM[966]) );
  XNOR U78 ( .A(B[966]), .B(A[966]), .Z(n78) );
  XOR U79 ( .A(n79), .B(n80), .Z(SUM[965]) );
  XNOR U80 ( .A(B[965]), .B(A[965]), .Z(n80) );
  XOR U81 ( .A(n81), .B(n82), .Z(SUM[964]) );
  XNOR U82 ( .A(B[964]), .B(A[964]), .Z(n82) );
  XOR U83 ( .A(n83), .B(n84), .Z(SUM[963]) );
  XNOR U84 ( .A(B[963]), .B(A[963]), .Z(n84) );
  XOR U85 ( .A(n85), .B(n86), .Z(SUM[962]) );
  XNOR U86 ( .A(B[962]), .B(A[962]), .Z(n86) );
  XOR U87 ( .A(n87), .B(n88), .Z(SUM[961]) );
  XNOR U88 ( .A(B[961]), .B(A[961]), .Z(n88) );
  XOR U89 ( .A(n89), .B(n90), .Z(SUM[960]) );
  XNOR U90 ( .A(B[960]), .B(A[960]), .Z(n90) );
  XOR U91 ( .A(n91), .B(n92), .Z(SUM[95]) );
  XNOR U92 ( .A(B[95]), .B(A[95]), .Z(n92) );
  XOR U93 ( .A(n93), .B(n94), .Z(SUM[959]) );
  XNOR U94 ( .A(B[959]), .B(A[959]), .Z(n94) );
  XOR U95 ( .A(n95), .B(n96), .Z(SUM[958]) );
  XNOR U96 ( .A(B[958]), .B(A[958]), .Z(n96) );
  XOR U97 ( .A(n97), .B(n98), .Z(SUM[957]) );
  XNOR U98 ( .A(B[957]), .B(A[957]), .Z(n98) );
  XOR U99 ( .A(n99), .B(n100), .Z(SUM[956]) );
  XNOR U100 ( .A(B[956]), .B(A[956]), .Z(n100) );
  XOR U101 ( .A(n101), .B(n102), .Z(SUM[955]) );
  XNOR U102 ( .A(B[955]), .B(A[955]), .Z(n102) );
  XOR U103 ( .A(n103), .B(n104), .Z(SUM[954]) );
  XNOR U104 ( .A(B[954]), .B(A[954]), .Z(n104) );
  XOR U105 ( .A(n105), .B(n106), .Z(SUM[953]) );
  XNOR U106 ( .A(B[953]), .B(A[953]), .Z(n106) );
  XOR U107 ( .A(n107), .B(n108), .Z(SUM[952]) );
  XNOR U108 ( .A(B[952]), .B(A[952]), .Z(n108) );
  XOR U109 ( .A(n109), .B(n110), .Z(SUM[951]) );
  XNOR U110 ( .A(B[951]), .B(A[951]), .Z(n110) );
  XOR U111 ( .A(n111), .B(n112), .Z(SUM[950]) );
  XNOR U112 ( .A(B[950]), .B(A[950]), .Z(n112) );
  XOR U113 ( .A(n113), .B(n114), .Z(SUM[94]) );
  XNOR U114 ( .A(B[94]), .B(A[94]), .Z(n114) );
  XOR U115 ( .A(n115), .B(n116), .Z(SUM[949]) );
  XNOR U116 ( .A(B[949]), .B(A[949]), .Z(n116) );
  XOR U117 ( .A(n117), .B(n118), .Z(SUM[948]) );
  XNOR U118 ( .A(B[948]), .B(A[948]), .Z(n118) );
  XOR U119 ( .A(n119), .B(n120), .Z(SUM[947]) );
  XNOR U120 ( .A(B[947]), .B(A[947]), .Z(n120) );
  XOR U121 ( .A(n121), .B(n122), .Z(SUM[946]) );
  XNOR U122 ( .A(B[946]), .B(A[946]), .Z(n122) );
  XOR U123 ( .A(n123), .B(n124), .Z(SUM[945]) );
  XNOR U124 ( .A(B[945]), .B(A[945]), .Z(n124) );
  XOR U125 ( .A(n125), .B(n126), .Z(SUM[944]) );
  XNOR U126 ( .A(B[944]), .B(A[944]), .Z(n126) );
  XOR U127 ( .A(n127), .B(n128), .Z(SUM[943]) );
  XNOR U128 ( .A(B[943]), .B(A[943]), .Z(n128) );
  XOR U129 ( .A(n129), .B(n130), .Z(SUM[942]) );
  XNOR U130 ( .A(B[942]), .B(A[942]), .Z(n130) );
  XOR U131 ( .A(n131), .B(n132), .Z(SUM[941]) );
  XNOR U132 ( .A(B[941]), .B(A[941]), .Z(n132) );
  XOR U133 ( .A(n133), .B(n134), .Z(SUM[940]) );
  XNOR U134 ( .A(B[940]), .B(A[940]), .Z(n134) );
  XOR U135 ( .A(n135), .B(n136), .Z(SUM[93]) );
  XNOR U136 ( .A(B[93]), .B(A[93]), .Z(n136) );
  XOR U137 ( .A(n137), .B(n138), .Z(SUM[939]) );
  XNOR U138 ( .A(B[939]), .B(A[939]), .Z(n138) );
  XOR U139 ( .A(n139), .B(n140), .Z(SUM[938]) );
  XNOR U140 ( .A(B[938]), .B(A[938]), .Z(n140) );
  XOR U141 ( .A(n141), .B(n142), .Z(SUM[937]) );
  XNOR U142 ( .A(B[937]), .B(A[937]), .Z(n142) );
  XOR U143 ( .A(n143), .B(n144), .Z(SUM[936]) );
  XNOR U144 ( .A(B[936]), .B(A[936]), .Z(n144) );
  XOR U145 ( .A(n145), .B(n146), .Z(SUM[935]) );
  XNOR U146 ( .A(B[935]), .B(A[935]), .Z(n146) );
  XOR U147 ( .A(n147), .B(n148), .Z(SUM[934]) );
  XNOR U148 ( .A(B[934]), .B(A[934]), .Z(n148) );
  XOR U149 ( .A(n149), .B(n150), .Z(SUM[933]) );
  XNOR U150 ( .A(B[933]), .B(A[933]), .Z(n150) );
  XOR U151 ( .A(n151), .B(n152), .Z(SUM[932]) );
  XNOR U152 ( .A(B[932]), .B(A[932]), .Z(n152) );
  XOR U153 ( .A(n153), .B(n154), .Z(SUM[931]) );
  XNOR U154 ( .A(B[931]), .B(A[931]), .Z(n154) );
  XOR U155 ( .A(n155), .B(n156), .Z(SUM[930]) );
  XNOR U156 ( .A(B[930]), .B(A[930]), .Z(n156) );
  XOR U157 ( .A(n157), .B(n158), .Z(SUM[92]) );
  XNOR U158 ( .A(B[92]), .B(A[92]), .Z(n158) );
  XOR U159 ( .A(n159), .B(n160), .Z(SUM[929]) );
  XNOR U160 ( .A(B[929]), .B(A[929]), .Z(n160) );
  XOR U161 ( .A(n161), .B(n162), .Z(SUM[928]) );
  XNOR U162 ( .A(B[928]), .B(A[928]), .Z(n162) );
  XOR U163 ( .A(n163), .B(n164), .Z(SUM[927]) );
  XNOR U164 ( .A(B[927]), .B(A[927]), .Z(n164) );
  XOR U165 ( .A(n165), .B(n166), .Z(SUM[926]) );
  XNOR U166 ( .A(B[926]), .B(A[926]), .Z(n166) );
  XOR U167 ( .A(n167), .B(n168), .Z(SUM[925]) );
  XNOR U168 ( .A(B[925]), .B(A[925]), .Z(n168) );
  XOR U169 ( .A(n169), .B(n170), .Z(SUM[924]) );
  XNOR U170 ( .A(B[924]), .B(A[924]), .Z(n170) );
  XOR U171 ( .A(n171), .B(n172), .Z(SUM[923]) );
  XNOR U172 ( .A(B[923]), .B(A[923]), .Z(n172) );
  XOR U173 ( .A(n173), .B(n174), .Z(SUM[922]) );
  XNOR U174 ( .A(B[922]), .B(A[922]), .Z(n174) );
  XOR U175 ( .A(n175), .B(n176), .Z(SUM[921]) );
  XNOR U176 ( .A(B[921]), .B(A[921]), .Z(n176) );
  XOR U177 ( .A(n177), .B(n178), .Z(SUM[920]) );
  XNOR U178 ( .A(B[920]), .B(A[920]), .Z(n178) );
  XOR U179 ( .A(n179), .B(n180), .Z(SUM[91]) );
  XNOR U180 ( .A(B[91]), .B(A[91]), .Z(n180) );
  XOR U181 ( .A(n181), .B(n182), .Z(SUM[919]) );
  XNOR U182 ( .A(B[919]), .B(A[919]), .Z(n182) );
  XOR U183 ( .A(n183), .B(n184), .Z(SUM[918]) );
  XNOR U184 ( .A(B[918]), .B(A[918]), .Z(n184) );
  XOR U185 ( .A(n185), .B(n186), .Z(SUM[917]) );
  XNOR U186 ( .A(B[917]), .B(A[917]), .Z(n186) );
  XOR U187 ( .A(n187), .B(n188), .Z(SUM[916]) );
  XNOR U188 ( .A(B[916]), .B(A[916]), .Z(n188) );
  XOR U189 ( .A(n189), .B(n190), .Z(SUM[915]) );
  XNOR U190 ( .A(B[915]), .B(A[915]), .Z(n190) );
  XOR U191 ( .A(n191), .B(n192), .Z(SUM[914]) );
  XNOR U192 ( .A(B[914]), .B(A[914]), .Z(n192) );
  XOR U193 ( .A(n193), .B(n194), .Z(SUM[913]) );
  XNOR U194 ( .A(B[913]), .B(A[913]), .Z(n194) );
  XOR U195 ( .A(n195), .B(n196), .Z(SUM[912]) );
  XNOR U196 ( .A(B[912]), .B(A[912]), .Z(n196) );
  XOR U197 ( .A(n197), .B(n198), .Z(SUM[911]) );
  XNOR U198 ( .A(B[911]), .B(A[911]), .Z(n198) );
  XOR U199 ( .A(n199), .B(n200), .Z(SUM[910]) );
  XNOR U200 ( .A(B[910]), .B(A[910]), .Z(n200) );
  XOR U201 ( .A(n201), .B(n202), .Z(SUM[90]) );
  XNOR U202 ( .A(B[90]), .B(A[90]), .Z(n202) );
  XOR U203 ( .A(n203), .B(n204), .Z(SUM[909]) );
  XNOR U204 ( .A(B[909]), .B(A[909]), .Z(n204) );
  XOR U205 ( .A(n205), .B(n206), .Z(SUM[908]) );
  XNOR U206 ( .A(B[908]), .B(A[908]), .Z(n206) );
  XOR U207 ( .A(n207), .B(n208), .Z(SUM[907]) );
  XNOR U208 ( .A(B[907]), .B(A[907]), .Z(n208) );
  XOR U209 ( .A(n209), .B(n210), .Z(SUM[906]) );
  XNOR U210 ( .A(B[906]), .B(A[906]), .Z(n210) );
  XOR U211 ( .A(n211), .B(n212), .Z(SUM[905]) );
  XNOR U212 ( .A(B[905]), .B(A[905]), .Z(n212) );
  XOR U213 ( .A(n213), .B(n214), .Z(SUM[904]) );
  XNOR U214 ( .A(B[904]), .B(A[904]), .Z(n214) );
  XOR U215 ( .A(n215), .B(n216), .Z(SUM[903]) );
  XNOR U216 ( .A(B[903]), .B(A[903]), .Z(n216) );
  XOR U217 ( .A(n217), .B(n218), .Z(SUM[902]) );
  XNOR U218 ( .A(B[902]), .B(A[902]), .Z(n218) );
  XOR U219 ( .A(n219), .B(n220), .Z(SUM[901]) );
  XNOR U220 ( .A(B[901]), .B(A[901]), .Z(n220) );
  XOR U221 ( .A(n221), .B(n222), .Z(SUM[900]) );
  XNOR U222 ( .A(B[900]), .B(A[900]), .Z(n222) );
  XOR U223 ( .A(n223), .B(n224), .Z(SUM[8]) );
  XNOR U224 ( .A(B[8]), .B(A[8]), .Z(n224) );
  XOR U225 ( .A(n225), .B(n226), .Z(SUM[89]) );
  XNOR U226 ( .A(B[89]), .B(A[89]), .Z(n226) );
  XOR U227 ( .A(n227), .B(n228), .Z(SUM[899]) );
  XNOR U228 ( .A(B[899]), .B(A[899]), .Z(n228) );
  XOR U229 ( .A(n229), .B(n230), .Z(SUM[898]) );
  XNOR U230 ( .A(B[898]), .B(A[898]), .Z(n230) );
  XOR U231 ( .A(n231), .B(n232), .Z(SUM[897]) );
  XNOR U232 ( .A(B[897]), .B(A[897]), .Z(n232) );
  XOR U233 ( .A(n233), .B(n234), .Z(SUM[896]) );
  XNOR U234 ( .A(B[896]), .B(A[896]), .Z(n234) );
  XOR U235 ( .A(n235), .B(n236), .Z(SUM[895]) );
  XNOR U236 ( .A(B[895]), .B(A[895]), .Z(n236) );
  XOR U237 ( .A(n237), .B(n238), .Z(SUM[894]) );
  XNOR U238 ( .A(B[894]), .B(A[894]), .Z(n238) );
  XOR U239 ( .A(n239), .B(n240), .Z(SUM[893]) );
  XNOR U240 ( .A(B[893]), .B(A[893]), .Z(n240) );
  XOR U241 ( .A(n241), .B(n242), .Z(SUM[892]) );
  XNOR U242 ( .A(B[892]), .B(A[892]), .Z(n242) );
  XOR U243 ( .A(n243), .B(n244), .Z(SUM[891]) );
  XNOR U244 ( .A(B[891]), .B(A[891]), .Z(n244) );
  XOR U245 ( .A(n245), .B(n246), .Z(SUM[890]) );
  XNOR U246 ( .A(B[890]), .B(A[890]), .Z(n246) );
  XOR U247 ( .A(n247), .B(n248), .Z(SUM[88]) );
  XNOR U248 ( .A(B[88]), .B(A[88]), .Z(n248) );
  XOR U249 ( .A(n249), .B(n250), .Z(SUM[889]) );
  XNOR U250 ( .A(B[889]), .B(A[889]), .Z(n250) );
  XOR U251 ( .A(n251), .B(n252), .Z(SUM[888]) );
  XNOR U252 ( .A(B[888]), .B(A[888]), .Z(n252) );
  XOR U253 ( .A(n253), .B(n254), .Z(SUM[887]) );
  XNOR U254 ( .A(B[887]), .B(A[887]), .Z(n254) );
  XOR U255 ( .A(n255), .B(n256), .Z(SUM[886]) );
  XNOR U256 ( .A(B[886]), .B(A[886]), .Z(n256) );
  XOR U257 ( .A(n257), .B(n258), .Z(SUM[885]) );
  XNOR U258 ( .A(B[885]), .B(A[885]), .Z(n258) );
  XOR U259 ( .A(n259), .B(n260), .Z(SUM[884]) );
  XNOR U260 ( .A(B[884]), .B(A[884]), .Z(n260) );
  XOR U261 ( .A(n261), .B(n262), .Z(SUM[883]) );
  XNOR U262 ( .A(B[883]), .B(A[883]), .Z(n262) );
  XOR U263 ( .A(n263), .B(n264), .Z(SUM[882]) );
  XNOR U264 ( .A(B[882]), .B(A[882]), .Z(n264) );
  XOR U265 ( .A(n265), .B(n266), .Z(SUM[881]) );
  XNOR U266 ( .A(B[881]), .B(A[881]), .Z(n266) );
  XOR U267 ( .A(n267), .B(n268), .Z(SUM[880]) );
  XNOR U268 ( .A(B[880]), .B(A[880]), .Z(n268) );
  XOR U269 ( .A(n269), .B(n270), .Z(SUM[87]) );
  XNOR U270 ( .A(B[87]), .B(A[87]), .Z(n270) );
  XOR U271 ( .A(n271), .B(n272), .Z(SUM[879]) );
  XNOR U272 ( .A(B[879]), .B(A[879]), .Z(n272) );
  XOR U273 ( .A(n273), .B(n274), .Z(SUM[878]) );
  XNOR U274 ( .A(B[878]), .B(A[878]), .Z(n274) );
  XOR U275 ( .A(n275), .B(n276), .Z(SUM[877]) );
  XNOR U276 ( .A(B[877]), .B(A[877]), .Z(n276) );
  XOR U277 ( .A(n277), .B(n278), .Z(SUM[876]) );
  XNOR U278 ( .A(B[876]), .B(A[876]), .Z(n278) );
  XOR U279 ( .A(n279), .B(n280), .Z(SUM[875]) );
  XNOR U280 ( .A(B[875]), .B(A[875]), .Z(n280) );
  XOR U281 ( .A(n281), .B(n282), .Z(SUM[874]) );
  XNOR U282 ( .A(B[874]), .B(A[874]), .Z(n282) );
  XOR U283 ( .A(n283), .B(n284), .Z(SUM[873]) );
  XNOR U284 ( .A(B[873]), .B(A[873]), .Z(n284) );
  XOR U285 ( .A(n285), .B(n286), .Z(SUM[872]) );
  XNOR U286 ( .A(B[872]), .B(A[872]), .Z(n286) );
  XOR U287 ( .A(n287), .B(n288), .Z(SUM[871]) );
  XNOR U288 ( .A(B[871]), .B(A[871]), .Z(n288) );
  XOR U289 ( .A(n289), .B(n290), .Z(SUM[870]) );
  XNOR U290 ( .A(B[870]), .B(A[870]), .Z(n290) );
  XOR U291 ( .A(n291), .B(n292), .Z(SUM[86]) );
  XNOR U292 ( .A(B[86]), .B(A[86]), .Z(n292) );
  XOR U293 ( .A(n293), .B(n294), .Z(SUM[869]) );
  XNOR U294 ( .A(B[869]), .B(A[869]), .Z(n294) );
  XOR U295 ( .A(n295), .B(n296), .Z(SUM[868]) );
  XNOR U296 ( .A(B[868]), .B(A[868]), .Z(n296) );
  XOR U297 ( .A(n297), .B(n298), .Z(SUM[867]) );
  XNOR U298 ( .A(B[867]), .B(A[867]), .Z(n298) );
  XOR U299 ( .A(n299), .B(n300), .Z(SUM[866]) );
  XNOR U300 ( .A(B[866]), .B(A[866]), .Z(n300) );
  XOR U301 ( .A(n301), .B(n302), .Z(SUM[865]) );
  XNOR U302 ( .A(B[865]), .B(A[865]), .Z(n302) );
  XOR U303 ( .A(n303), .B(n304), .Z(SUM[864]) );
  XNOR U304 ( .A(B[864]), .B(A[864]), .Z(n304) );
  XOR U305 ( .A(n305), .B(n306), .Z(SUM[863]) );
  XNOR U306 ( .A(B[863]), .B(A[863]), .Z(n306) );
  XOR U307 ( .A(n307), .B(n308), .Z(SUM[862]) );
  XNOR U308 ( .A(B[862]), .B(A[862]), .Z(n308) );
  XOR U309 ( .A(n309), .B(n310), .Z(SUM[861]) );
  XNOR U310 ( .A(B[861]), .B(A[861]), .Z(n310) );
  XOR U311 ( .A(n311), .B(n312), .Z(SUM[860]) );
  XNOR U312 ( .A(B[860]), .B(A[860]), .Z(n312) );
  XOR U313 ( .A(n313), .B(n314), .Z(SUM[85]) );
  XNOR U314 ( .A(B[85]), .B(A[85]), .Z(n314) );
  XOR U315 ( .A(n315), .B(n316), .Z(SUM[859]) );
  XNOR U316 ( .A(B[859]), .B(A[859]), .Z(n316) );
  XOR U317 ( .A(n317), .B(n318), .Z(SUM[858]) );
  XNOR U318 ( .A(B[858]), .B(A[858]), .Z(n318) );
  XOR U319 ( .A(n319), .B(n320), .Z(SUM[857]) );
  XNOR U320 ( .A(B[857]), .B(A[857]), .Z(n320) );
  XOR U321 ( .A(n321), .B(n322), .Z(SUM[856]) );
  XNOR U322 ( .A(B[856]), .B(A[856]), .Z(n322) );
  XOR U323 ( .A(n323), .B(n324), .Z(SUM[855]) );
  XNOR U324 ( .A(B[855]), .B(A[855]), .Z(n324) );
  XOR U325 ( .A(n325), .B(n326), .Z(SUM[854]) );
  XNOR U326 ( .A(B[854]), .B(A[854]), .Z(n326) );
  XOR U327 ( .A(n327), .B(n328), .Z(SUM[853]) );
  XNOR U328 ( .A(B[853]), .B(A[853]), .Z(n328) );
  XOR U329 ( .A(n329), .B(n330), .Z(SUM[852]) );
  XNOR U330 ( .A(B[852]), .B(A[852]), .Z(n330) );
  XOR U331 ( .A(n331), .B(n332), .Z(SUM[851]) );
  XNOR U332 ( .A(B[851]), .B(A[851]), .Z(n332) );
  XOR U333 ( .A(n333), .B(n334), .Z(SUM[850]) );
  XNOR U334 ( .A(B[850]), .B(A[850]), .Z(n334) );
  XOR U335 ( .A(n335), .B(n336), .Z(SUM[84]) );
  XNOR U336 ( .A(B[84]), .B(A[84]), .Z(n336) );
  XOR U337 ( .A(n337), .B(n338), .Z(SUM[849]) );
  XNOR U338 ( .A(B[849]), .B(A[849]), .Z(n338) );
  XOR U339 ( .A(n339), .B(n340), .Z(SUM[848]) );
  XNOR U340 ( .A(B[848]), .B(A[848]), .Z(n340) );
  XOR U341 ( .A(n341), .B(n342), .Z(SUM[847]) );
  XNOR U342 ( .A(B[847]), .B(A[847]), .Z(n342) );
  XOR U343 ( .A(n343), .B(n344), .Z(SUM[846]) );
  XNOR U344 ( .A(B[846]), .B(A[846]), .Z(n344) );
  XOR U345 ( .A(n345), .B(n346), .Z(SUM[845]) );
  XNOR U346 ( .A(B[845]), .B(A[845]), .Z(n346) );
  XOR U347 ( .A(n347), .B(n348), .Z(SUM[844]) );
  XNOR U348 ( .A(B[844]), .B(A[844]), .Z(n348) );
  XOR U349 ( .A(n349), .B(n350), .Z(SUM[843]) );
  XNOR U350 ( .A(B[843]), .B(A[843]), .Z(n350) );
  XOR U351 ( .A(n351), .B(n352), .Z(SUM[842]) );
  XNOR U352 ( .A(B[842]), .B(A[842]), .Z(n352) );
  XOR U353 ( .A(n353), .B(n354), .Z(SUM[841]) );
  XNOR U354 ( .A(B[841]), .B(A[841]), .Z(n354) );
  XOR U355 ( .A(n355), .B(n356), .Z(SUM[840]) );
  XNOR U356 ( .A(B[840]), .B(A[840]), .Z(n356) );
  XOR U357 ( .A(n357), .B(n358), .Z(SUM[83]) );
  XNOR U358 ( .A(B[83]), .B(A[83]), .Z(n358) );
  XOR U359 ( .A(n359), .B(n360), .Z(SUM[839]) );
  XNOR U360 ( .A(B[839]), .B(A[839]), .Z(n360) );
  XOR U361 ( .A(n361), .B(n362), .Z(SUM[838]) );
  XNOR U362 ( .A(B[838]), .B(A[838]), .Z(n362) );
  XOR U363 ( .A(n363), .B(n364), .Z(SUM[837]) );
  XNOR U364 ( .A(B[837]), .B(A[837]), .Z(n364) );
  XOR U365 ( .A(n365), .B(n366), .Z(SUM[836]) );
  XNOR U366 ( .A(B[836]), .B(A[836]), .Z(n366) );
  XOR U367 ( .A(n367), .B(n368), .Z(SUM[835]) );
  XNOR U368 ( .A(B[835]), .B(A[835]), .Z(n368) );
  XOR U369 ( .A(n369), .B(n370), .Z(SUM[834]) );
  XNOR U370 ( .A(B[834]), .B(A[834]), .Z(n370) );
  XOR U371 ( .A(n371), .B(n372), .Z(SUM[833]) );
  XNOR U372 ( .A(B[833]), .B(A[833]), .Z(n372) );
  XOR U373 ( .A(n373), .B(n374), .Z(SUM[832]) );
  XNOR U374 ( .A(B[832]), .B(A[832]), .Z(n374) );
  XOR U375 ( .A(n375), .B(n376), .Z(SUM[831]) );
  XNOR U376 ( .A(B[831]), .B(A[831]), .Z(n376) );
  XOR U377 ( .A(n377), .B(n378), .Z(SUM[830]) );
  XNOR U378 ( .A(B[830]), .B(A[830]), .Z(n378) );
  XOR U379 ( .A(n379), .B(n380), .Z(SUM[82]) );
  XNOR U380 ( .A(B[82]), .B(A[82]), .Z(n380) );
  XOR U381 ( .A(n381), .B(n382), .Z(SUM[829]) );
  XNOR U382 ( .A(B[829]), .B(A[829]), .Z(n382) );
  XOR U383 ( .A(n383), .B(n384), .Z(SUM[828]) );
  XNOR U384 ( .A(B[828]), .B(A[828]), .Z(n384) );
  XOR U385 ( .A(n385), .B(n386), .Z(SUM[827]) );
  XNOR U386 ( .A(B[827]), .B(A[827]), .Z(n386) );
  XOR U387 ( .A(n387), .B(n388), .Z(SUM[826]) );
  XNOR U388 ( .A(B[826]), .B(A[826]), .Z(n388) );
  XOR U389 ( .A(n389), .B(n390), .Z(SUM[825]) );
  XNOR U390 ( .A(B[825]), .B(A[825]), .Z(n390) );
  XOR U391 ( .A(n391), .B(n392), .Z(SUM[824]) );
  XNOR U392 ( .A(B[824]), .B(A[824]), .Z(n392) );
  XOR U393 ( .A(n393), .B(n394), .Z(SUM[823]) );
  XNOR U394 ( .A(B[823]), .B(A[823]), .Z(n394) );
  XOR U395 ( .A(n395), .B(n396), .Z(SUM[822]) );
  XNOR U396 ( .A(B[822]), .B(A[822]), .Z(n396) );
  XOR U397 ( .A(n397), .B(n398), .Z(SUM[821]) );
  XNOR U398 ( .A(B[821]), .B(A[821]), .Z(n398) );
  XOR U399 ( .A(n399), .B(n400), .Z(SUM[820]) );
  XNOR U400 ( .A(B[820]), .B(A[820]), .Z(n400) );
  XOR U401 ( .A(n401), .B(n402), .Z(SUM[81]) );
  XNOR U402 ( .A(B[81]), .B(A[81]), .Z(n402) );
  XOR U403 ( .A(n403), .B(n404), .Z(SUM[819]) );
  XNOR U404 ( .A(B[819]), .B(A[819]), .Z(n404) );
  XOR U405 ( .A(n405), .B(n406), .Z(SUM[818]) );
  XNOR U406 ( .A(B[818]), .B(A[818]), .Z(n406) );
  XOR U407 ( .A(n407), .B(n408), .Z(SUM[817]) );
  XNOR U408 ( .A(B[817]), .B(A[817]), .Z(n408) );
  XOR U409 ( .A(n409), .B(n410), .Z(SUM[816]) );
  XNOR U410 ( .A(B[816]), .B(A[816]), .Z(n410) );
  XOR U411 ( .A(n411), .B(n412), .Z(SUM[815]) );
  XNOR U412 ( .A(B[815]), .B(A[815]), .Z(n412) );
  XOR U413 ( .A(n413), .B(n414), .Z(SUM[814]) );
  XNOR U414 ( .A(B[814]), .B(A[814]), .Z(n414) );
  XOR U415 ( .A(n415), .B(n416), .Z(SUM[813]) );
  XNOR U416 ( .A(B[813]), .B(A[813]), .Z(n416) );
  XOR U417 ( .A(n417), .B(n418), .Z(SUM[812]) );
  XNOR U418 ( .A(B[812]), .B(A[812]), .Z(n418) );
  XOR U419 ( .A(n419), .B(n420), .Z(SUM[811]) );
  XNOR U420 ( .A(B[811]), .B(A[811]), .Z(n420) );
  XOR U421 ( .A(n421), .B(n422), .Z(SUM[810]) );
  XNOR U422 ( .A(B[810]), .B(A[810]), .Z(n422) );
  XOR U423 ( .A(n423), .B(n424), .Z(SUM[80]) );
  XNOR U424 ( .A(B[80]), .B(A[80]), .Z(n424) );
  XOR U425 ( .A(n425), .B(n426), .Z(SUM[809]) );
  XNOR U426 ( .A(B[809]), .B(A[809]), .Z(n426) );
  XOR U427 ( .A(n427), .B(n428), .Z(SUM[808]) );
  XNOR U428 ( .A(B[808]), .B(A[808]), .Z(n428) );
  XOR U429 ( .A(n429), .B(n430), .Z(SUM[807]) );
  XNOR U430 ( .A(B[807]), .B(A[807]), .Z(n430) );
  XOR U431 ( .A(n431), .B(n432), .Z(SUM[806]) );
  XNOR U432 ( .A(B[806]), .B(A[806]), .Z(n432) );
  XOR U433 ( .A(n433), .B(n434), .Z(SUM[805]) );
  XNOR U434 ( .A(B[805]), .B(A[805]), .Z(n434) );
  XOR U435 ( .A(n435), .B(n436), .Z(SUM[804]) );
  XNOR U436 ( .A(B[804]), .B(A[804]), .Z(n436) );
  XOR U437 ( .A(n437), .B(n438), .Z(SUM[803]) );
  XNOR U438 ( .A(B[803]), .B(A[803]), .Z(n438) );
  XOR U439 ( .A(n439), .B(n440), .Z(SUM[802]) );
  XNOR U440 ( .A(B[802]), .B(A[802]), .Z(n440) );
  XOR U441 ( .A(n441), .B(n442), .Z(SUM[801]) );
  XNOR U442 ( .A(B[801]), .B(A[801]), .Z(n442) );
  XOR U443 ( .A(n443), .B(n444), .Z(SUM[800]) );
  XNOR U444 ( .A(B[800]), .B(A[800]), .Z(n444) );
  XOR U445 ( .A(n445), .B(n446), .Z(SUM[7]) );
  XNOR U446 ( .A(B[7]), .B(A[7]), .Z(n446) );
  XOR U447 ( .A(n447), .B(n448), .Z(SUM[79]) );
  XNOR U448 ( .A(B[79]), .B(A[79]), .Z(n448) );
  XOR U449 ( .A(n449), .B(n450), .Z(SUM[799]) );
  XNOR U450 ( .A(B[799]), .B(A[799]), .Z(n450) );
  XOR U451 ( .A(n451), .B(n452), .Z(SUM[798]) );
  XNOR U452 ( .A(B[798]), .B(A[798]), .Z(n452) );
  XOR U453 ( .A(n453), .B(n454), .Z(SUM[797]) );
  XNOR U454 ( .A(B[797]), .B(A[797]), .Z(n454) );
  XOR U455 ( .A(n455), .B(n456), .Z(SUM[796]) );
  XNOR U456 ( .A(B[796]), .B(A[796]), .Z(n456) );
  XOR U457 ( .A(n457), .B(n458), .Z(SUM[795]) );
  XNOR U458 ( .A(B[795]), .B(A[795]), .Z(n458) );
  XOR U459 ( .A(n459), .B(n460), .Z(SUM[794]) );
  XNOR U460 ( .A(B[794]), .B(A[794]), .Z(n460) );
  XOR U461 ( .A(n461), .B(n462), .Z(SUM[793]) );
  XNOR U462 ( .A(B[793]), .B(A[793]), .Z(n462) );
  XOR U463 ( .A(n463), .B(n464), .Z(SUM[792]) );
  XNOR U464 ( .A(B[792]), .B(A[792]), .Z(n464) );
  XOR U465 ( .A(n465), .B(n466), .Z(SUM[791]) );
  XNOR U466 ( .A(B[791]), .B(A[791]), .Z(n466) );
  XOR U467 ( .A(n467), .B(n468), .Z(SUM[790]) );
  XNOR U468 ( .A(B[790]), .B(A[790]), .Z(n468) );
  XOR U469 ( .A(n469), .B(n470), .Z(SUM[78]) );
  XNOR U470 ( .A(B[78]), .B(A[78]), .Z(n470) );
  XOR U471 ( .A(n471), .B(n472), .Z(SUM[789]) );
  XNOR U472 ( .A(B[789]), .B(A[789]), .Z(n472) );
  XOR U473 ( .A(n473), .B(n474), .Z(SUM[788]) );
  XNOR U474 ( .A(B[788]), .B(A[788]), .Z(n474) );
  XOR U475 ( .A(n475), .B(n476), .Z(SUM[787]) );
  XNOR U476 ( .A(B[787]), .B(A[787]), .Z(n476) );
  XOR U477 ( .A(n477), .B(n478), .Z(SUM[786]) );
  XNOR U478 ( .A(B[786]), .B(A[786]), .Z(n478) );
  XOR U479 ( .A(n479), .B(n480), .Z(SUM[785]) );
  XNOR U480 ( .A(B[785]), .B(A[785]), .Z(n480) );
  XOR U481 ( .A(n481), .B(n482), .Z(SUM[784]) );
  XNOR U482 ( .A(B[784]), .B(A[784]), .Z(n482) );
  XOR U483 ( .A(n483), .B(n484), .Z(SUM[783]) );
  XNOR U484 ( .A(B[783]), .B(A[783]), .Z(n484) );
  XOR U485 ( .A(n485), .B(n486), .Z(SUM[782]) );
  XNOR U486 ( .A(B[782]), .B(A[782]), .Z(n486) );
  XOR U487 ( .A(n487), .B(n488), .Z(SUM[781]) );
  XNOR U488 ( .A(B[781]), .B(A[781]), .Z(n488) );
  XOR U489 ( .A(n489), .B(n490), .Z(SUM[780]) );
  XNOR U490 ( .A(B[780]), .B(A[780]), .Z(n490) );
  XOR U491 ( .A(n491), .B(n492), .Z(SUM[77]) );
  XNOR U492 ( .A(B[77]), .B(A[77]), .Z(n492) );
  XOR U493 ( .A(n493), .B(n494), .Z(SUM[779]) );
  XNOR U494 ( .A(B[779]), .B(A[779]), .Z(n494) );
  XOR U495 ( .A(n495), .B(n496), .Z(SUM[778]) );
  XNOR U496 ( .A(B[778]), .B(A[778]), .Z(n496) );
  XOR U497 ( .A(n497), .B(n498), .Z(SUM[777]) );
  XNOR U498 ( .A(B[777]), .B(A[777]), .Z(n498) );
  XOR U499 ( .A(n499), .B(n500), .Z(SUM[776]) );
  XNOR U500 ( .A(B[776]), .B(A[776]), .Z(n500) );
  XOR U501 ( .A(n501), .B(n502), .Z(SUM[775]) );
  XNOR U502 ( .A(B[775]), .B(A[775]), .Z(n502) );
  XOR U503 ( .A(n503), .B(n504), .Z(SUM[774]) );
  XNOR U504 ( .A(B[774]), .B(A[774]), .Z(n504) );
  XOR U505 ( .A(n505), .B(n506), .Z(SUM[773]) );
  XNOR U506 ( .A(B[773]), .B(A[773]), .Z(n506) );
  XOR U507 ( .A(n507), .B(n508), .Z(SUM[772]) );
  XNOR U508 ( .A(B[772]), .B(A[772]), .Z(n508) );
  XOR U509 ( .A(n509), .B(n510), .Z(SUM[771]) );
  XNOR U510 ( .A(B[771]), .B(A[771]), .Z(n510) );
  XOR U511 ( .A(n511), .B(n512), .Z(SUM[770]) );
  XNOR U512 ( .A(B[770]), .B(A[770]), .Z(n512) );
  XOR U513 ( .A(n513), .B(n514), .Z(SUM[76]) );
  XNOR U514 ( .A(B[76]), .B(A[76]), .Z(n514) );
  XOR U515 ( .A(n515), .B(n516), .Z(SUM[769]) );
  XNOR U516 ( .A(B[769]), .B(A[769]), .Z(n516) );
  XOR U517 ( .A(n517), .B(n518), .Z(SUM[768]) );
  XNOR U518 ( .A(B[768]), .B(A[768]), .Z(n518) );
  XOR U519 ( .A(n519), .B(n520), .Z(SUM[767]) );
  XNOR U520 ( .A(B[767]), .B(A[767]), .Z(n520) );
  XOR U521 ( .A(n521), .B(n522), .Z(SUM[766]) );
  XNOR U522 ( .A(B[766]), .B(A[766]), .Z(n522) );
  XOR U523 ( .A(n523), .B(n524), .Z(SUM[765]) );
  XNOR U524 ( .A(B[765]), .B(A[765]), .Z(n524) );
  XOR U525 ( .A(n525), .B(n526), .Z(SUM[764]) );
  XNOR U526 ( .A(B[764]), .B(A[764]), .Z(n526) );
  XOR U527 ( .A(n527), .B(n528), .Z(SUM[763]) );
  XNOR U528 ( .A(B[763]), .B(A[763]), .Z(n528) );
  XOR U529 ( .A(n529), .B(n530), .Z(SUM[762]) );
  XNOR U530 ( .A(B[762]), .B(A[762]), .Z(n530) );
  XOR U531 ( .A(n531), .B(n532), .Z(SUM[761]) );
  XNOR U532 ( .A(B[761]), .B(A[761]), .Z(n532) );
  XOR U533 ( .A(n533), .B(n534), .Z(SUM[760]) );
  XNOR U534 ( .A(B[760]), .B(A[760]), .Z(n534) );
  XOR U535 ( .A(n535), .B(n536), .Z(SUM[75]) );
  XNOR U536 ( .A(B[75]), .B(A[75]), .Z(n536) );
  XOR U537 ( .A(n537), .B(n538), .Z(SUM[759]) );
  XNOR U538 ( .A(B[759]), .B(A[759]), .Z(n538) );
  XOR U539 ( .A(n539), .B(n540), .Z(SUM[758]) );
  XNOR U540 ( .A(B[758]), .B(A[758]), .Z(n540) );
  XOR U541 ( .A(n541), .B(n542), .Z(SUM[757]) );
  XNOR U542 ( .A(B[757]), .B(A[757]), .Z(n542) );
  XOR U543 ( .A(n543), .B(n544), .Z(SUM[756]) );
  XNOR U544 ( .A(B[756]), .B(A[756]), .Z(n544) );
  XOR U545 ( .A(n545), .B(n546), .Z(SUM[755]) );
  XNOR U546 ( .A(B[755]), .B(A[755]), .Z(n546) );
  XOR U547 ( .A(n547), .B(n548), .Z(SUM[754]) );
  XNOR U548 ( .A(B[754]), .B(A[754]), .Z(n548) );
  XOR U549 ( .A(n549), .B(n550), .Z(SUM[753]) );
  XNOR U550 ( .A(B[753]), .B(A[753]), .Z(n550) );
  XOR U551 ( .A(n551), .B(n552), .Z(SUM[752]) );
  XNOR U552 ( .A(B[752]), .B(A[752]), .Z(n552) );
  XOR U553 ( .A(n553), .B(n554), .Z(SUM[751]) );
  XNOR U554 ( .A(B[751]), .B(A[751]), .Z(n554) );
  XOR U555 ( .A(n555), .B(n556), .Z(SUM[750]) );
  XNOR U556 ( .A(B[750]), .B(A[750]), .Z(n556) );
  XOR U557 ( .A(n557), .B(n558), .Z(SUM[74]) );
  XNOR U558 ( .A(B[74]), .B(A[74]), .Z(n558) );
  XOR U559 ( .A(n559), .B(n560), .Z(SUM[749]) );
  XNOR U560 ( .A(B[749]), .B(A[749]), .Z(n560) );
  XOR U561 ( .A(n561), .B(n562), .Z(SUM[748]) );
  XNOR U562 ( .A(B[748]), .B(A[748]), .Z(n562) );
  XOR U563 ( .A(n563), .B(n564), .Z(SUM[747]) );
  XNOR U564 ( .A(B[747]), .B(A[747]), .Z(n564) );
  XOR U565 ( .A(n565), .B(n566), .Z(SUM[746]) );
  XNOR U566 ( .A(B[746]), .B(A[746]), .Z(n566) );
  XOR U567 ( .A(n567), .B(n568), .Z(SUM[745]) );
  XNOR U568 ( .A(B[745]), .B(A[745]), .Z(n568) );
  XOR U569 ( .A(n569), .B(n570), .Z(SUM[744]) );
  XNOR U570 ( .A(B[744]), .B(A[744]), .Z(n570) );
  XOR U571 ( .A(n571), .B(n572), .Z(SUM[743]) );
  XNOR U572 ( .A(B[743]), .B(A[743]), .Z(n572) );
  XOR U573 ( .A(n573), .B(n574), .Z(SUM[742]) );
  XNOR U574 ( .A(B[742]), .B(A[742]), .Z(n574) );
  XOR U575 ( .A(n575), .B(n576), .Z(SUM[741]) );
  XNOR U576 ( .A(B[741]), .B(A[741]), .Z(n576) );
  XOR U577 ( .A(n577), .B(n578), .Z(SUM[740]) );
  XNOR U578 ( .A(B[740]), .B(A[740]), .Z(n578) );
  XOR U579 ( .A(n579), .B(n580), .Z(SUM[73]) );
  XNOR U580 ( .A(B[73]), .B(A[73]), .Z(n580) );
  XOR U581 ( .A(n581), .B(n582), .Z(SUM[739]) );
  XNOR U582 ( .A(B[739]), .B(A[739]), .Z(n582) );
  XOR U583 ( .A(n583), .B(n584), .Z(SUM[738]) );
  XNOR U584 ( .A(B[738]), .B(A[738]), .Z(n584) );
  XOR U585 ( .A(n585), .B(n586), .Z(SUM[737]) );
  XNOR U586 ( .A(B[737]), .B(A[737]), .Z(n586) );
  XOR U587 ( .A(n587), .B(n588), .Z(SUM[736]) );
  XNOR U588 ( .A(B[736]), .B(A[736]), .Z(n588) );
  XOR U589 ( .A(n589), .B(n590), .Z(SUM[735]) );
  XNOR U590 ( .A(B[735]), .B(A[735]), .Z(n590) );
  XOR U591 ( .A(n591), .B(n592), .Z(SUM[734]) );
  XNOR U592 ( .A(B[734]), .B(A[734]), .Z(n592) );
  XOR U593 ( .A(n593), .B(n594), .Z(SUM[733]) );
  XNOR U594 ( .A(B[733]), .B(A[733]), .Z(n594) );
  XOR U595 ( .A(n595), .B(n596), .Z(SUM[732]) );
  XNOR U596 ( .A(B[732]), .B(A[732]), .Z(n596) );
  XOR U597 ( .A(n597), .B(n598), .Z(SUM[731]) );
  XNOR U598 ( .A(B[731]), .B(A[731]), .Z(n598) );
  XOR U599 ( .A(n599), .B(n600), .Z(SUM[730]) );
  XNOR U600 ( .A(B[730]), .B(A[730]), .Z(n600) );
  XOR U601 ( .A(n601), .B(n602), .Z(SUM[72]) );
  XNOR U602 ( .A(B[72]), .B(A[72]), .Z(n602) );
  XOR U603 ( .A(n603), .B(n604), .Z(SUM[729]) );
  XNOR U604 ( .A(B[729]), .B(A[729]), .Z(n604) );
  XOR U605 ( .A(n605), .B(n606), .Z(SUM[728]) );
  XNOR U606 ( .A(B[728]), .B(A[728]), .Z(n606) );
  XOR U607 ( .A(n607), .B(n608), .Z(SUM[727]) );
  XNOR U608 ( .A(B[727]), .B(A[727]), .Z(n608) );
  XOR U609 ( .A(n609), .B(n610), .Z(SUM[726]) );
  XNOR U610 ( .A(B[726]), .B(A[726]), .Z(n610) );
  XOR U611 ( .A(n611), .B(n612), .Z(SUM[725]) );
  XNOR U612 ( .A(B[725]), .B(A[725]), .Z(n612) );
  XOR U613 ( .A(n613), .B(n614), .Z(SUM[724]) );
  XNOR U614 ( .A(B[724]), .B(A[724]), .Z(n614) );
  XOR U615 ( .A(n615), .B(n616), .Z(SUM[723]) );
  XNOR U616 ( .A(B[723]), .B(A[723]), .Z(n616) );
  XOR U617 ( .A(n617), .B(n618), .Z(SUM[722]) );
  XNOR U618 ( .A(B[722]), .B(A[722]), .Z(n618) );
  XOR U619 ( .A(n619), .B(n620), .Z(SUM[721]) );
  XNOR U620 ( .A(B[721]), .B(A[721]), .Z(n620) );
  XOR U621 ( .A(n621), .B(n622), .Z(SUM[720]) );
  XNOR U622 ( .A(B[720]), .B(A[720]), .Z(n622) );
  XOR U623 ( .A(n623), .B(n624), .Z(SUM[71]) );
  XNOR U624 ( .A(B[71]), .B(A[71]), .Z(n624) );
  XOR U625 ( .A(n625), .B(n626), .Z(SUM[719]) );
  XNOR U626 ( .A(B[719]), .B(A[719]), .Z(n626) );
  XOR U627 ( .A(n627), .B(n628), .Z(SUM[718]) );
  XNOR U628 ( .A(B[718]), .B(A[718]), .Z(n628) );
  XOR U629 ( .A(n629), .B(n630), .Z(SUM[717]) );
  XNOR U630 ( .A(B[717]), .B(A[717]), .Z(n630) );
  XOR U631 ( .A(n631), .B(n632), .Z(SUM[716]) );
  XNOR U632 ( .A(B[716]), .B(A[716]), .Z(n632) );
  XOR U633 ( .A(n633), .B(n634), .Z(SUM[715]) );
  XNOR U634 ( .A(B[715]), .B(A[715]), .Z(n634) );
  XOR U635 ( .A(n635), .B(n636), .Z(SUM[714]) );
  XNOR U636 ( .A(B[714]), .B(A[714]), .Z(n636) );
  XOR U637 ( .A(n637), .B(n638), .Z(SUM[713]) );
  XNOR U638 ( .A(B[713]), .B(A[713]), .Z(n638) );
  XOR U639 ( .A(n639), .B(n640), .Z(SUM[712]) );
  XNOR U640 ( .A(B[712]), .B(A[712]), .Z(n640) );
  XOR U641 ( .A(n641), .B(n642), .Z(SUM[711]) );
  XNOR U642 ( .A(B[711]), .B(A[711]), .Z(n642) );
  XOR U643 ( .A(n643), .B(n644), .Z(SUM[710]) );
  XNOR U644 ( .A(B[710]), .B(A[710]), .Z(n644) );
  XOR U645 ( .A(n645), .B(n646), .Z(SUM[70]) );
  XNOR U646 ( .A(B[70]), .B(A[70]), .Z(n646) );
  XOR U647 ( .A(n647), .B(n648), .Z(SUM[709]) );
  XNOR U648 ( .A(B[709]), .B(A[709]), .Z(n648) );
  XOR U649 ( .A(n649), .B(n650), .Z(SUM[708]) );
  XNOR U650 ( .A(B[708]), .B(A[708]), .Z(n650) );
  XOR U651 ( .A(n651), .B(n652), .Z(SUM[707]) );
  XNOR U652 ( .A(B[707]), .B(A[707]), .Z(n652) );
  XOR U653 ( .A(n653), .B(n654), .Z(SUM[706]) );
  XNOR U654 ( .A(B[706]), .B(A[706]), .Z(n654) );
  XOR U655 ( .A(n655), .B(n656), .Z(SUM[705]) );
  XNOR U656 ( .A(B[705]), .B(A[705]), .Z(n656) );
  XOR U657 ( .A(n657), .B(n658), .Z(SUM[704]) );
  XNOR U658 ( .A(B[704]), .B(A[704]), .Z(n658) );
  XOR U659 ( .A(n659), .B(n660), .Z(SUM[703]) );
  XNOR U660 ( .A(B[703]), .B(A[703]), .Z(n660) );
  XOR U661 ( .A(n661), .B(n662), .Z(SUM[702]) );
  XNOR U662 ( .A(B[702]), .B(A[702]), .Z(n662) );
  XOR U663 ( .A(n663), .B(n664), .Z(SUM[701]) );
  XNOR U664 ( .A(B[701]), .B(A[701]), .Z(n664) );
  XOR U665 ( .A(n665), .B(n666), .Z(SUM[700]) );
  XNOR U666 ( .A(B[700]), .B(A[700]), .Z(n666) );
  XOR U667 ( .A(n667), .B(n668), .Z(SUM[6]) );
  XNOR U668 ( .A(B[6]), .B(A[6]), .Z(n668) );
  XOR U669 ( .A(n669), .B(n670), .Z(SUM[69]) );
  XNOR U670 ( .A(B[69]), .B(A[69]), .Z(n670) );
  XOR U671 ( .A(n671), .B(n672), .Z(SUM[699]) );
  XNOR U672 ( .A(B[699]), .B(A[699]), .Z(n672) );
  XOR U673 ( .A(n673), .B(n674), .Z(SUM[698]) );
  XNOR U674 ( .A(B[698]), .B(A[698]), .Z(n674) );
  XOR U675 ( .A(n675), .B(n676), .Z(SUM[697]) );
  XNOR U676 ( .A(B[697]), .B(A[697]), .Z(n676) );
  XOR U677 ( .A(n677), .B(n678), .Z(SUM[696]) );
  XNOR U678 ( .A(B[696]), .B(A[696]), .Z(n678) );
  XOR U679 ( .A(n679), .B(n680), .Z(SUM[695]) );
  XNOR U680 ( .A(B[695]), .B(A[695]), .Z(n680) );
  XOR U681 ( .A(n681), .B(n682), .Z(SUM[694]) );
  XNOR U682 ( .A(B[694]), .B(A[694]), .Z(n682) );
  XOR U683 ( .A(n683), .B(n684), .Z(SUM[693]) );
  XNOR U684 ( .A(B[693]), .B(A[693]), .Z(n684) );
  XOR U685 ( .A(n685), .B(n686), .Z(SUM[692]) );
  XNOR U686 ( .A(B[692]), .B(A[692]), .Z(n686) );
  XOR U687 ( .A(n687), .B(n688), .Z(SUM[691]) );
  XNOR U688 ( .A(B[691]), .B(A[691]), .Z(n688) );
  XOR U689 ( .A(n689), .B(n690), .Z(SUM[690]) );
  XNOR U690 ( .A(B[690]), .B(A[690]), .Z(n690) );
  XOR U691 ( .A(n691), .B(n692), .Z(SUM[68]) );
  XNOR U692 ( .A(B[68]), .B(A[68]), .Z(n692) );
  XOR U693 ( .A(n693), .B(n694), .Z(SUM[689]) );
  XNOR U694 ( .A(B[689]), .B(A[689]), .Z(n694) );
  XOR U695 ( .A(n695), .B(n696), .Z(SUM[688]) );
  XNOR U696 ( .A(B[688]), .B(A[688]), .Z(n696) );
  XOR U697 ( .A(n697), .B(n698), .Z(SUM[687]) );
  XNOR U698 ( .A(B[687]), .B(A[687]), .Z(n698) );
  XOR U699 ( .A(n699), .B(n700), .Z(SUM[686]) );
  XNOR U700 ( .A(B[686]), .B(A[686]), .Z(n700) );
  XOR U701 ( .A(n701), .B(n702), .Z(SUM[685]) );
  XNOR U702 ( .A(B[685]), .B(A[685]), .Z(n702) );
  XOR U703 ( .A(n703), .B(n704), .Z(SUM[684]) );
  XNOR U704 ( .A(B[684]), .B(A[684]), .Z(n704) );
  XOR U705 ( .A(n705), .B(n706), .Z(SUM[683]) );
  XNOR U706 ( .A(B[683]), .B(A[683]), .Z(n706) );
  XOR U707 ( .A(n707), .B(n708), .Z(SUM[682]) );
  XNOR U708 ( .A(B[682]), .B(A[682]), .Z(n708) );
  XOR U709 ( .A(n709), .B(n710), .Z(SUM[681]) );
  XNOR U710 ( .A(B[681]), .B(A[681]), .Z(n710) );
  XOR U711 ( .A(n711), .B(n712), .Z(SUM[680]) );
  XNOR U712 ( .A(B[680]), .B(A[680]), .Z(n712) );
  XOR U713 ( .A(n713), .B(n714), .Z(SUM[67]) );
  XNOR U714 ( .A(B[67]), .B(A[67]), .Z(n714) );
  XOR U715 ( .A(n715), .B(n716), .Z(SUM[679]) );
  XNOR U716 ( .A(B[679]), .B(A[679]), .Z(n716) );
  XOR U717 ( .A(n717), .B(n718), .Z(SUM[678]) );
  XNOR U718 ( .A(B[678]), .B(A[678]), .Z(n718) );
  XOR U719 ( .A(n719), .B(n720), .Z(SUM[677]) );
  XNOR U720 ( .A(B[677]), .B(A[677]), .Z(n720) );
  XOR U721 ( .A(n721), .B(n722), .Z(SUM[676]) );
  XNOR U722 ( .A(B[676]), .B(A[676]), .Z(n722) );
  XOR U723 ( .A(n723), .B(n724), .Z(SUM[675]) );
  XNOR U724 ( .A(B[675]), .B(A[675]), .Z(n724) );
  XOR U725 ( .A(n725), .B(n726), .Z(SUM[674]) );
  XNOR U726 ( .A(B[674]), .B(A[674]), .Z(n726) );
  XOR U727 ( .A(n727), .B(n728), .Z(SUM[673]) );
  XNOR U728 ( .A(B[673]), .B(A[673]), .Z(n728) );
  XOR U729 ( .A(n729), .B(n730), .Z(SUM[672]) );
  XNOR U730 ( .A(B[672]), .B(A[672]), .Z(n730) );
  XOR U731 ( .A(n731), .B(n732), .Z(SUM[671]) );
  XNOR U732 ( .A(B[671]), .B(A[671]), .Z(n732) );
  XOR U733 ( .A(n733), .B(n734), .Z(SUM[670]) );
  XNOR U734 ( .A(B[670]), .B(A[670]), .Z(n734) );
  XOR U735 ( .A(n735), .B(n736), .Z(SUM[66]) );
  XNOR U736 ( .A(B[66]), .B(A[66]), .Z(n736) );
  XOR U737 ( .A(n737), .B(n738), .Z(SUM[669]) );
  XNOR U738 ( .A(B[669]), .B(A[669]), .Z(n738) );
  XOR U739 ( .A(n739), .B(n740), .Z(SUM[668]) );
  XNOR U740 ( .A(B[668]), .B(A[668]), .Z(n740) );
  XOR U741 ( .A(n741), .B(n742), .Z(SUM[667]) );
  XNOR U742 ( .A(B[667]), .B(A[667]), .Z(n742) );
  XOR U743 ( .A(n743), .B(n744), .Z(SUM[666]) );
  XNOR U744 ( .A(B[666]), .B(A[666]), .Z(n744) );
  XOR U745 ( .A(n745), .B(n746), .Z(SUM[665]) );
  XNOR U746 ( .A(B[665]), .B(A[665]), .Z(n746) );
  XOR U747 ( .A(n747), .B(n748), .Z(SUM[664]) );
  XNOR U748 ( .A(B[664]), .B(A[664]), .Z(n748) );
  XOR U749 ( .A(n749), .B(n750), .Z(SUM[663]) );
  XNOR U750 ( .A(B[663]), .B(A[663]), .Z(n750) );
  XOR U751 ( .A(n751), .B(n752), .Z(SUM[662]) );
  XNOR U752 ( .A(B[662]), .B(A[662]), .Z(n752) );
  XOR U753 ( .A(n753), .B(n754), .Z(SUM[661]) );
  XNOR U754 ( .A(B[661]), .B(A[661]), .Z(n754) );
  XOR U755 ( .A(n755), .B(n756), .Z(SUM[660]) );
  XNOR U756 ( .A(B[660]), .B(A[660]), .Z(n756) );
  XOR U757 ( .A(n757), .B(n758), .Z(SUM[65]) );
  XNOR U758 ( .A(B[65]), .B(A[65]), .Z(n758) );
  XOR U759 ( .A(n759), .B(n760), .Z(SUM[659]) );
  XNOR U760 ( .A(B[659]), .B(A[659]), .Z(n760) );
  XOR U761 ( .A(n761), .B(n762), .Z(SUM[658]) );
  XNOR U762 ( .A(B[658]), .B(A[658]), .Z(n762) );
  XOR U763 ( .A(n763), .B(n764), .Z(SUM[657]) );
  XNOR U764 ( .A(B[657]), .B(A[657]), .Z(n764) );
  XOR U765 ( .A(n765), .B(n766), .Z(SUM[656]) );
  XNOR U766 ( .A(B[656]), .B(A[656]), .Z(n766) );
  XOR U767 ( .A(n767), .B(n768), .Z(SUM[655]) );
  XNOR U768 ( .A(B[655]), .B(A[655]), .Z(n768) );
  XOR U769 ( .A(n769), .B(n770), .Z(SUM[654]) );
  XNOR U770 ( .A(B[654]), .B(A[654]), .Z(n770) );
  XOR U771 ( .A(n771), .B(n772), .Z(SUM[653]) );
  XNOR U772 ( .A(B[653]), .B(A[653]), .Z(n772) );
  XOR U773 ( .A(n773), .B(n774), .Z(SUM[652]) );
  XNOR U774 ( .A(B[652]), .B(A[652]), .Z(n774) );
  XOR U775 ( .A(n775), .B(n776), .Z(SUM[651]) );
  XNOR U776 ( .A(B[651]), .B(A[651]), .Z(n776) );
  XOR U777 ( .A(n777), .B(n778), .Z(SUM[650]) );
  XNOR U778 ( .A(B[650]), .B(A[650]), .Z(n778) );
  XOR U779 ( .A(n779), .B(n780), .Z(SUM[64]) );
  XNOR U780 ( .A(B[64]), .B(A[64]), .Z(n780) );
  XOR U781 ( .A(n781), .B(n782), .Z(SUM[649]) );
  XNOR U782 ( .A(B[649]), .B(A[649]), .Z(n782) );
  XOR U783 ( .A(n783), .B(n784), .Z(SUM[648]) );
  XNOR U784 ( .A(B[648]), .B(A[648]), .Z(n784) );
  XOR U785 ( .A(n785), .B(n786), .Z(SUM[647]) );
  XNOR U786 ( .A(B[647]), .B(A[647]), .Z(n786) );
  XOR U787 ( .A(n787), .B(n788), .Z(SUM[646]) );
  XNOR U788 ( .A(B[646]), .B(A[646]), .Z(n788) );
  XOR U789 ( .A(n789), .B(n790), .Z(SUM[645]) );
  XNOR U790 ( .A(B[645]), .B(A[645]), .Z(n790) );
  XOR U791 ( .A(n791), .B(n792), .Z(SUM[644]) );
  XNOR U792 ( .A(B[644]), .B(A[644]), .Z(n792) );
  XOR U793 ( .A(n793), .B(n794), .Z(SUM[643]) );
  XNOR U794 ( .A(B[643]), .B(A[643]), .Z(n794) );
  XOR U795 ( .A(n795), .B(n796), .Z(SUM[642]) );
  XNOR U796 ( .A(B[642]), .B(A[642]), .Z(n796) );
  XOR U797 ( .A(n797), .B(n798), .Z(SUM[641]) );
  XNOR U798 ( .A(B[641]), .B(A[641]), .Z(n798) );
  XOR U799 ( .A(n799), .B(n800), .Z(SUM[640]) );
  XNOR U800 ( .A(B[640]), .B(A[640]), .Z(n800) );
  XOR U801 ( .A(n801), .B(n802), .Z(SUM[63]) );
  XNOR U802 ( .A(B[63]), .B(A[63]), .Z(n802) );
  XOR U803 ( .A(n803), .B(n804), .Z(SUM[639]) );
  XNOR U804 ( .A(B[639]), .B(A[639]), .Z(n804) );
  XOR U805 ( .A(n805), .B(n806), .Z(SUM[638]) );
  XNOR U806 ( .A(B[638]), .B(A[638]), .Z(n806) );
  XOR U807 ( .A(n807), .B(n808), .Z(SUM[637]) );
  XNOR U808 ( .A(B[637]), .B(A[637]), .Z(n808) );
  XOR U809 ( .A(n809), .B(n810), .Z(SUM[636]) );
  XNOR U810 ( .A(B[636]), .B(A[636]), .Z(n810) );
  XOR U811 ( .A(n811), .B(n812), .Z(SUM[635]) );
  XNOR U812 ( .A(B[635]), .B(A[635]), .Z(n812) );
  XOR U813 ( .A(n813), .B(n814), .Z(SUM[634]) );
  XNOR U814 ( .A(B[634]), .B(A[634]), .Z(n814) );
  XOR U815 ( .A(n815), .B(n816), .Z(SUM[633]) );
  XNOR U816 ( .A(B[633]), .B(A[633]), .Z(n816) );
  XOR U817 ( .A(n817), .B(n818), .Z(SUM[632]) );
  XNOR U818 ( .A(B[632]), .B(A[632]), .Z(n818) );
  XOR U819 ( .A(n819), .B(n820), .Z(SUM[631]) );
  XNOR U820 ( .A(B[631]), .B(A[631]), .Z(n820) );
  XOR U821 ( .A(n821), .B(n822), .Z(SUM[630]) );
  XNOR U822 ( .A(B[630]), .B(A[630]), .Z(n822) );
  XOR U823 ( .A(n823), .B(n824), .Z(SUM[62]) );
  XNOR U824 ( .A(B[62]), .B(A[62]), .Z(n824) );
  XOR U825 ( .A(n825), .B(n826), .Z(SUM[629]) );
  XNOR U826 ( .A(B[629]), .B(A[629]), .Z(n826) );
  XOR U827 ( .A(n827), .B(n828), .Z(SUM[628]) );
  XNOR U828 ( .A(B[628]), .B(A[628]), .Z(n828) );
  XOR U829 ( .A(n829), .B(n830), .Z(SUM[627]) );
  XNOR U830 ( .A(B[627]), .B(A[627]), .Z(n830) );
  XOR U831 ( .A(n831), .B(n832), .Z(SUM[626]) );
  XNOR U832 ( .A(B[626]), .B(A[626]), .Z(n832) );
  XOR U833 ( .A(n833), .B(n834), .Z(SUM[625]) );
  XNOR U834 ( .A(B[625]), .B(A[625]), .Z(n834) );
  XOR U835 ( .A(n835), .B(n836), .Z(SUM[624]) );
  XNOR U836 ( .A(B[624]), .B(A[624]), .Z(n836) );
  XOR U837 ( .A(n837), .B(n838), .Z(SUM[623]) );
  XNOR U838 ( .A(B[623]), .B(A[623]), .Z(n838) );
  XOR U839 ( .A(n839), .B(n840), .Z(SUM[622]) );
  XNOR U840 ( .A(B[622]), .B(A[622]), .Z(n840) );
  XOR U841 ( .A(n841), .B(n842), .Z(SUM[621]) );
  XNOR U842 ( .A(B[621]), .B(A[621]), .Z(n842) );
  XOR U843 ( .A(n843), .B(n844), .Z(SUM[620]) );
  XNOR U844 ( .A(B[620]), .B(A[620]), .Z(n844) );
  XOR U845 ( .A(n845), .B(n846), .Z(SUM[61]) );
  XNOR U846 ( .A(B[61]), .B(A[61]), .Z(n846) );
  XOR U847 ( .A(n847), .B(n848), .Z(SUM[619]) );
  XNOR U848 ( .A(B[619]), .B(A[619]), .Z(n848) );
  XOR U849 ( .A(n849), .B(n850), .Z(SUM[618]) );
  XNOR U850 ( .A(B[618]), .B(A[618]), .Z(n850) );
  XOR U851 ( .A(n851), .B(n852), .Z(SUM[617]) );
  XNOR U852 ( .A(B[617]), .B(A[617]), .Z(n852) );
  XOR U853 ( .A(n853), .B(n854), .Z(SUM[616]) );
  XNOR U854 ( .A(B[616]), .B(A[616]), .Z(n854) );
  XOR U855 ( .A(n855), .B(n856), .Z(SUM[615]) );
  XNOR U856 ( .A(B[615]), .B(A[615]), .Z(n856) );
  XOR U857 ( .A(n857), .B(n858), .Z(SUM[614]) );
  XNOR U858 ( .A(B[614]), .B(A[614]), .Z(n858) );
  XOR U859 ( .A(n859), .B(n860), .Z(SUM[613]) );
  XNOR U860 ( .A(B[613]), .B(A[613]), .Z(n860) );
  XOR U861 ( .A(n861), .B(n862), .Z(SUM[612]) );
  XNOR U862 ( .A(B[612]), .B(A[612]), .Z(n862) );
  XOR U863 ( .A(n863), .B(n864), .Z(SUM[611]) );
  XNOR U864 ( .A(B[611]), .B(A[611]), .Z(n864) );
  XOR U865 ( .A(n865), .B(n866), .Z(SUM[610]) );
  XNOR U866 ( .A(B[610]), .B(A[610]), .Z(n866) );
  XOR U867 ( .A(n867), .B(n868), .Z(SUM[60]) );
  XNOR U868 ( .A(B[60]), .B(A[60]), .Z(n868) );
  XOR U869 ( .A(n869), .B(n870), .Z(SUM[609]) );
  XNOR U870 ( .A(B[609]), .B(A[609]), .Z(n870) );
  XOR U871 ( .A(n871), .B(n872), .Z(SUM[608]) );
  XNOR U872 ( .A(B[608]), .B(A[608]), .Z(n872) );
  XOR U873 ( .A(n873), .B(n874), .Z(SUM[607]) );
  XNOR U874 ( .A(B[607]), .B(A[607]), .Z(n874) );
  XOR U875 ( .A(n875), .B(n876), .Z(SUM[606]) );
  XNOR U876 ( .A(B[606]), .B(A[606]), .Z(n876) );
  XOR U877 ( .A(n877), .B(n878), .Z(SUM[605]) );
  XNOR U878 ( .A(B[605]), .B(A[605]), .Z(n878) );
  XOR U879 ( .A(n879), .B(n880), .Z(SUM[604]) );
  XNOR U880 ( .A(B[604]), .B(A[604]), .Z(n880) );
  XOR U881 ( .A(n881), .B(n882), .Z(SUM[603]) );
  XNOR U882 ( .A(B[603]), .B(A[603]), .Z(n882) );
  XOR U883 ( .A(n883), .B(n884), .Z(SUM[602]) );
  XNOR U884 ( .A(B[602]), .B(A[602]), .Z(n884) );
  XOR U885 ( .A(n885), .B(n886), .Z(SUM[601]) );
  XNOR U886 ( .A(B[601]), .B(A[601]), .Z(n886) );
  XOR U887 ( .A(n887), .B(n888), .Z(SUM[600]) );
  XNOR U888 ( .A(B[600]), .B(A[600]), .Z(n888) );
  XOR U889 ( .A(n889), .B(n890), .Z(SUM[5]) );
  XNOR U890 ( .A(B[5]), .B(A[5]), .Z(n890) );
  XOR U891 ( .A(n891), .B(n892), .Z(SUM[59]) );
  XNOR U892 ( .A(B[59]), .B(A[59]), .Z(n892) );
  XOR U893 ( .A(n893), .B(n894), .Z(SUM[599]) );
  XNOR U894 ( .A(B[599]), .B(A[599]), .Z(n894) );
  XOR U895 ( .A(n895), .B(n896), .Z(SUM[598]) );
  XNOR U896 ( .A(B[598]), .B(A[598]), .Z(n896) );
  XOR U897 ( .A(n897), .B(n898), .Z(SUM[597]) );
  XNOR U898 ( .A(B[597]), .B(A[597]), .Z(n898) );
  XOR U899 ( .A(n899), .B(n900), .Z(SUM[596]) );
  XNOR U900 ( .A(B[596]), .B(A[596]), .Z(n900) );
  XOR U901 ( .A(n901), .B(n902), .Z(SUM[595]) );
  XNOR U902 ( .A(B[595]), .B(A[595]), .Z(n902) );
  XOR U903 ( .A(n903), .B(n904), .Z(SUM[594]) );
  XNOR U904 ( .A(B[594]), .B(A[594]), .Z(n904) );
  XOR U905 ( .A(n905), .B(n906), .Z(SUM[593]) );
  XNOR U906 ( .A(B[593]), .B(A[593]), .Z(n906) );
  XOR U907 ( .A(n907), .B(n908), .Z(SUM[592]) );
  XNOR U908 ( .A(B[592]), .B(A[592]), .Z(n908) );
  XOR U909 ( .A(n909), .B(n910), .Z(SUM[591]) );
  XNOR U910 ( .A(B[591]), .B(A[591]), .Z(n910) );
  XOR U911 ( .A(n911), .B(n912), .Z(SUM[590]) );
  XNOR U912 ( .A(B[590]), .B(A[590]), .Z(n912) );
  XOR U913 ( .A(n913), .B(n914), .Z(SUM[58]) );
  XNOR U914 ( .A(B[58]), .B(A[58]), .Z(n914) );
  XOR U915 ( .A(n915), .B(n916), .Z(SUM[589]) );
  XNOR U916 ( .A(B[589]), .B(A[589]), .Z(n916) );
  XOR U917 ( .A(n917), .B(n918), .Z(SUM[588]) );
  XNOR U918 ( .A(B[588]), .B(A[588]), .Z(n918) );
  XOR U919 ( .A(n919), .B(n920), .Z(SUM[587]) );
  XNOR U920 ( .A(B[587]), .B(A[587]), .Z(n920) );
  XOR U921 ( .A(n921), .B(n922), .Z(SUM[586]) );
  XNOR U922 ( .A(B[586]), .B(A[586]), .Z(n922) );
  XOR U923 ( .A(n923), .B(n924), .Z(SUM[585]) );
  XNOR U924 ( .A(B[585]), .B(A[585]), .Z(n924) );
  XOR U925 ( .A(n925), .B(n926), .Z(SUM[584]) );
  XNOR U926 ( .A(B[584]), .B(A[584]), .Z(n926) );
  XOR U927 ( .A(n927), .B(n928), .Z(SUM[583]) );
  XNOR U928 ( .A(B[583]), .B(A[583]), .Z(n928) );
  XOR U929 ( .A(n929), .B(n930), .Z(SUM[582]) );
  XNOR U930 ( .A(B[582]), .B(A[582]), .Z(n930) );
  XOR U931 ( .A(n931), .B(n932), .Z(SUM[581]) );
  XNOR U932 ( .A(B[581]), .B(A[581]), .Z(n932) );
  XOR U933 ( .A(n933), .B(n934), .Z(SUM[580]) );
  XNOR U934 ( .A(B[580]), .B(A[580]), .Z(n934) );
  XOR U935 ( .A(n935), .B(n936), .Z(SUM[57]) );
  XNOR U936 ( .A(B[57]), .B(A[57]), .Z(n936) );
  XOR U937 ( .A(n937), .B(n938), .Z(SUM[579]) );
  XNOR U938 ( .A(B[579]), .B(A[579]), .Z(n938) );
  XOR U939 ( .A(n939), .B(n940), .Z(SUM[578]) );
  XNOR U940 ( .A(B[578]), .B(A[578]), .Z(n940) );
  XOR U941 ( .A(n941), .B(n942), .Z(SUM[577]) );
  XNOR U942 ( .A(B[577]), .B(A[577]), .Z(n942) );
  XOR U943 ( .A(n943), .B(n944), .Z(SUM[576]) );
  XNOR U944 ( .A(B[576]), .B(A[576]), .Z(n944) );
  XOR U945 ( .A(n945), .B(n946), .Z(SUM[575]) );
  XNOR U946 ( .A(B[575]), .B(A[575]), .Z(n946) );
  XOR U947 ( .A(n947), .B(n948), .Z(SUM[574]) );
  XNOR U948 ( .A(B[574]), .B(A[574]), .Z(n948) );
  XOR U949 ( .A(n949), .B(n950), .Z(SUM[573]) );
  XNOR U950 ( .A(B[573]), .B(A[573]), .Z(n950) );
  XOR U951 ( .A(n951), .B(n952), .Z(SUM[572]) );
  XNOR U952 ( .A(B[572]), .B(A[572]), .Z(n952) );
  XOR U953 ( .A(n953), .B(n954), .Z(SUM[571]) );
  XNOR U954 ( .A(B[571]), .B(A[571]), .Z(n954) );
  XOR U955 ( .A(n955), .B(n956), .Z(SUM[570]) );
  XNOR U956 ( .A(B[570]), .B(A[570]), .Z(n956) );
  XOR U957 ( .A(n957), .B(n958), .Z(SUM[56]) );
  XNOR U958 ( .A(B[56]), .B(A[56]), .Z(n958) );
  XOR U959 ( .A(n959), .B(n960), .Z(SUM[569]) );
  XNOR U960 ( .A(B[569]), .B(A[569]), .Z(n960) );
  XOR U961 ( .A(n961), .B(n962), .Z(SUM[568]) );
  XNOR U962 ( .A(B[568]), .B(A[568]), .Z(n962) );
  XOR U963 ( .A(n963), .B(n964), .Z(SUM[567]) );
  XNOR U964 ( .A(B[567]), .B(A[567]), .Z(n964) );
  XOR U965 ( .A(n965), .B(n966), .Z(SUM[566]) );
  XNOR U966 ( .A(B[566]), .B(A[566]), .Z(n966) );
  XOR U967 ( .A(n967), .B(n968), .Z(SUM[565]) );
  XNOR U968 ( .A(B[565]), .B(A[565]), .Z(n968) );
  XOR U969 ( .A(n969), .B(n970), .Z(SUM[564]) );
  XNOR U970 ( .A(B[564]), .B(A[564]), .Z(n970) );
  XOR U971 ( .A(n971), .B(n972), .Z(SUM[563]) );
  XNOR U972 ( .A(B[563]), .B(A[563]), .Z(n972) );
  XOR U973 ( .A(n973), .B(n974), .Z(SUM[562]) );
  XNOR U974 ( .A(B[562]), .B(A[562]), .Z(n974) );
  XOR U975 ( .A(n975), .B(n976), .Z(SUM[561]) );
  XNOR U976 ( .A(B[561]), .B(A[561]), .Z(n976) );
  XOR U977 ( .A(n977), .B(n978), .Z(SUM[560]) );
  XNOR U978 ( .A(B[560]), .B(A[560]), .Z(n978) );
  XOR U979 ( .A(n979), .B(n980), .Z(SUM[55]) );
  XNOR U980 ( .A(B[55]), .B(A[55]), .Z(n980) );
  XOR U981 ( .A(n981), .B(n982), .Z(SUM[559]) );
  XNOR U982 ( .A(B[559]), .B(A[559]), .Z(n982) );
  XOR U983 ( .A(n983), .B(n984), .Z(SUM[558]) );
  XNOR U984 ( .A(B[558]), .B(A[558]), .Z(n984) );
  XOR U985 ( .A(n985), .B(n986), .Z(SUM[557]) );
  XNOR U986 ( .A(B[557]), .B(A[557]), .Z(n986) );
  XOR U987 ( .A(n987), .B(n988), .Z(SUM[556]) );
  XNOR U988 ( .A(B[556]), .B(A[556]), .Z(n988) );
  XOR U989 ( .A(n989), .B(n990), .Z(SUM[555]) );
  XNOR U990 ( .A(B[555]), .B(A[555]), .Z(n990) );
  XOR U991 ( .A(n991), .B(n992), .Z(SUM[554]) );
  XNOR U992 ( .A(B[554]), .B(A[554]), .Z(n992) );
  XOR U993 ( .A(n993), .B(n994), .Z(SUM[553]) );
  XNOR U994 ( .A(B[553]), .B(A[553]), .Z(n994) );
  XOR U995 ( .A(n995), .B(n996), .Z(SUM[552]) );
  XNOR U996 ( .A(B[552]), .B(A[552]), .Z(n996) );
  XOR U997 ( .A(n997), .B(n998), .Z(SUM[551]) );
  XNOR U998 ( .A(B[551]), .B(A[551]), .Z(n998) );
  XOR U999 ( .A(n999), .B(n1000), .Z(SUM[550]) );
  XNOR U1000 ( .A(B[550]), .B(A[550]), .Z(n1000) );
  XOR U1001 ( .A(n1001), .B(n1002), .Z(SUM[54]) );
  XNOR U1002 ( .A(B[54]), .B(A[54]), .Z(n1002) );
  XOR U1003 ( .A(n1003), .B(n1004), .Z(SUM[549]) );
  XNOR U1004 ( .A(B[549]), .B(A[549]), .Z(n1004) );
  XOR U1005 ( .A(n1005), .B(n1006), .Z(SUM[548]) );
  XNOR U1006 ( .A(B[548]), .B(A[548]), .Z(n1006) );
  XOR U1007 ( .A(n1007), .B(n1008), .Z(SUM[547]) );
  XNOR U1008 ( .A(B[547]), .B(A[547]), .Z(n1008) );
  XOR U1009 ( .A(n1009), .B(n1010), .Z(SUM[546]) );
  XNOR U1010 ( .A(B[546]), .B(A[546]), .Z(n1010) );
  XOR U1011 ( .A(n1011), .B(n1012), .Z(SUM[545]) );
  XNOR U1012 ( .A(B[545]), .B(A[545]), .Z(n1012) );
  XOR U1013 ( .A(n1013), .B(n1014), .Z(SUM[544]) );
  XNOR U1014 ( .A(B[544]), .B(A[544]), .Z(n1014) );
  XOR U1015 ( .A(n1015), .B(n1016), .Z(SUM[543]) );
  XNOR U1016 ( .A(B[543]), .B(A[543]), .Z(n1016) );
  XOR U1017 ( .A(n1017), .B(n1018), .Z(SUM[542]) );
  XNOR U1018 ( .A(B[542]), .B(A[542]), .Z(n1018) );
  XOR U1019 ( .A(n1019), .B(n1020), .Z(SUM[541]) );
  XNOR U1020 ( .A(B[541]), .B(A[541]), .Z(n1020) );
  XOR U1021 ( .A(n1021), .B(n1022), .Z(SUM[540]) );
  XNOR U1022 ( .A(B[540]), .B(A[540]), .Z(n1022) );
  XOR U1023 ( .A(n1023), .B(n1024), .Z(SUM[53]) );
  XNOR U1024 ( .A(B[53]), .B(A[53]), .Z(n1024) );
  XOR U1025 ( .A(n1025), .B(n1026), .Z(SUM[539]) );
  XNOR U1026 ( .A(B[539]), .B(A[539]), .Z(n1026) );
  XOR U1027 ( .A(n1027), .B(n1028), .Z(SUM[538]) );
  XNOR U1028 ( .A(B[538]), .B(A[538]), .Z(n1028) );
  XOR U1029 ( .A(n1029), .B(n1030), .Z(SUM[537]) );
  XNOR U1030 ( .A(B[537]), .B(A[537]), .Z(n1030) );
  XOR U1031 ( .A(n1031), .B(n1032), .Z(SUM[536]) );
  XNOR U1032 ( .A(B[536]), .B(A[536]), .Z(n1032) );
  XOR U1033 ( .A(n1033), .B(n1034), .Z(SUM[535]) );
  XNOR U1034 ( .A(B[535]), .B(A[535]), .Z(n1034) );
  XOR U1035 ( .A(n1035), .B(n1036), .Z(SUM[534]) );
  XNOR U1036 ( .A(B[534]), .B(A[534]), .Z(n1036) );
  XOR U1037 ( .A(n1037), .B(n1038), .Z(SUM[533]) );
  XNOR U1038 ( .A(B[533]), .B(A[533]), .Z(n1038) );
  XOR U1039 ( .A(n1039), .B(n1040), .Z(SUM[532]) );
  XNOR U1040 ( .A(B[532]), .B(A[532]), .Z(n1040) );
  XOR U1041 ( .A(n1041), .B(n1042), .Z(SUM[531]) );
  XNOR U1042 ( .A(B[531]), .B(A[531]), .Z(n1042) );
  XOR U1043 ( .A(n1043), .B(n1044), .Z(SUM[530]) );
  XNOR U1044 ( .A(B[530]), .B(A[530]), .Z(n1044) );
  XOR U1045 ( .A(n1045), .B(n1046), .Z(SUM[52]) );
  XNOR U1046 ( .A(B[52]), .B(A[52]), .Z(n1046) );
  XOR U1047 ( .A(n1047), .B(n1048), .Z(SUM[529]) );
  XNOR U1048 ( .A(B[529]), .B(A[529]), .Z(n1048) );
  XOR U1049 ( .A(n1049), .B(n1050), .Z(SUM[528]) );
  XNOR U1050 ( .A(B[528]), .B(A[528]), .Z(n1050) );
  XOR U1051 ( .A(n1051), .B(n1052), .Z(SUM[527]) );
  XNOR U1052 ( .A(B[527]), .B(A[527]), .Z(n1052) );
  XOR U1053 ( .A(n1053), .B(n1054), .Z(SUM[526]) );
  XNOR U1054 ( .A(B[526]), .B(A[526]), .Z(n1054) );
  XOR U1055 ( .A(n1055), .B(n1056), .Z(SUM[525]) );
  XNOR U1056 ( .A(B[525]), .B(A[525]), .Z(n1056) );
  XOR U1057 ( .A(n1057), .B(n1058), .Z(SUM[524]) );
  XNOR U1058 ( .A(B[524]), .B(A[524]), .Z(n1058) );
  XOR U1059 ( .A(n1059), .B(n1060), .Z(SUM[523]) );
  XNOR U1060 ( .A(B[523]), .B(A[523]), .Z(n1060) );
  XOR U1061 ( .A(n1061), .B(n1062), .Z(SUM[522]) );
  XNOR U1062 ( .A(B[522]), .B(A[522]), .Z(n1062) );
  XOR U1063 ( .A(n1063), .B(n1064), .Z(SUM[521]) );
  XNOR U1064 ( .A(B[521]), .B(A[521]), .Z(n1064) );
  XOR U1065 ( .A(n1065), .B(n1066), .Z(SUM[520]) );
  XNOR U1066 ( .A(B[520]), .B(A[520]), .Z(n1066) );
  XOR U1067 ( .A(n1067), .B(n1068), .Z(SUM[51]) );
  XNOR U1068 ( .A(B[51]), .B(A[51]), .Z(n1068) );
  XOR U1069 ( .A(n1069), .B(n1070), .Z(SUM[519]) );
  XNOR U1070 ( .A(B[519]), .B(A[519]), .Z(n1070) );
  XOR U1071 ( .A(n1071), .B(n1072), .Z(SUM[518]) );
  XNOR U1072 ( .A(B[518]), .B(A[518]), .Z(n1072) );
  XOR U1073 ( .A(n1073), .B(n1074), .Z(SUM[517]) );
  XNOR U1074 ( .A(B[517]), .B(A[517]), .Z(n1074) );
  XOR U1075 ( .A(n1075), .B(n1076), .Z(SUM[516]) );
  XNOR U1076 ( .A(B[516]), .B(A[516]), .Z(n1076) );
  XOR U1077 ( .A(n1077), .B(n1078), .Z(SUM[515]) );
  XNOR U1078 ( .A(B[515]), .B(A[515]), .Z(n1078) );
  XOR U1079 ( .A(n1079), .B(n1080), .Z(SUM[514]) );
  XNOR U1080 ( .A(B[514]), .B(A[514]), .Z(n1080) );
  XOR U1081 ( .A(n1081), .B(n1082), .Z(SUM[513]) );
  XNOR U1082 ( .A(B[513]), .B(A[513]), .Z(n1082) );
  XOR U1083 ( .A(n1083), .B(n1084), .Z(SUM[512]) );
  XNOR U1084 ( .A(B[512]), .B(A[512]), .Z(n1084) );
  XOR U1085 ( .A(n1085), .B(n1086), .Z(SUM[511]) );
  XNOR U1086 ( .A(B[511]), .B(A[511]), .Z(n1086) );
  XOR U1087 ( .A(n1087), .B(n1088), .Z(SUM[510]) );
  XNOR U1088 ( .A(B[510]), .B(A[510]), .Z(n1088) );
  XOR U1089 ( .A(n1089), .B(n1090), .Z(SUM[50]) );
  XNOR U1090 ( .A(B[50]), .B(A[50]), .Z(n1090) );
  XOR U1091 ( .A(n1091), .B(n1092), .Z(SUM[509]) );
  XNOR U1092 ( .A(B[509]), .B(A[509]), .Z(n1092) );
  XOR U1093 ( .A(n1093), .B(n1094), .Z(SUM[508]) );
  XNOR U1094 ( .A(B[508]), .B(A[508]), .Z(n1094) );
  XOR U1095 ( .A(n1095), .B(n1096), .Z(SUM[507]) );
  XNOR U1096 ( .A(B[507]), .B(A[507]), .Z(n1096) );
  XOR U1097 ( .A(n1097), .B(n1098), .Z(SUM[506]) );
  XNOR U1098 ( .A(B[506]), .B(A[506]), .Z(n1098) );
  XOR U1099 ( .A(n1099), .B(n1100), .Z(SUM[505]) );
  XNOR U1100 ( .A(B[505]), .B(A[505]), .Z(n1100) );
  XOR U1101 ( .A(n1101), .B(n1102), .Z(SUM[504]) );
  XNOR U1102 ( .A(B[504]), .B(A[504]), .Z(n1102) );
  XOR U1103 ( .A(n1103), .B(n1104), .Z(SUM[503]) );
  XNOR U1104 ( .A(B[503]), .B(A[503]), .Z(n1104) );
  XOR U1105 ( .A(n1105), .B(n1106), .Z(SUM[502]) );
  XNOR U1106 ( .A(B[502]), .B(A[502]), .Z(n1106) );
  XOR U1107 ( .A(n1107), .B(n1108), .Z(SUM[501]) );
  XNOR U1108 ( .A(B[501]), .B(A[501]), .Z(n1108) );
  XOR U1109 ( .A(n1109), .B(n1110), .Z(SUM[500]) );
  XNOR U1110 ( .A(B[500]), .B(A[500]), .Z(n1110) );
  XOR U1111 ( .A(n1111), .B(n1112), .Z(SUM[4]) );
  XNOR U1112 ( .A(B[4]), .B(A[4]), .Z(n1112) );
  XOR U1113 ( .A(n1113), .B(n1114), .Z(SUM[49]) );
  XNOR U1114 ( .A(B[49]), .B(A[49]), .Z(n1114) );
  XOR U1115 ( .A(n1115), .B(n1116), .Z(SUM[499]) );
  XNOR U1116 ( .A(B[499]), .B(A[499]), .Z(n1116) );
  XOR U1117 ( .A(n1117), .B(n1118), .Z(SUM[498]) );
  XNOR U1118 ( .A(B[498]), .B(A[498]), .Z(n1118) );
  XOR U1119 ( .A(n1119), .B(n1120), .Z(SUM[497]) );
  XNOR U1120 ( .A(B[497]), .B(A[497]), .Z(n1120) );
  XOR U1121 ( .A(n1121), .B(n1122), .Z(SUM[496]) );
  XNOR U1122 ( .A(B[496]), .B(A[496]), .Z(n1122) );
  XOR U1123 ( .A(n1123), .B(n1124), .Z(SUM[495]) );
  XNOR U1124 ( .A(B[495]), .B(A[495]), .Z(n1124) );
  XOR U1125 ( .A(n1125), .B(n1126), .Z(SUM[494]) );
  XNOR U1126 ( .A(B[494]), .B(A[494]), .Z(n1126) );
  XOR U1127 ( .A(n1127), .B(n1128), .Z(SUM[493]) );
  XNOR U1128 ( .A(B[493]), .B(A[493]), .Z(n1128) );
  XOR U1129 ( .A(n1129), .B(n1130), .Z(SUM[492]) );
  XNOR U1130 ( .A(B[492]), .B(A[492]), .Z(n1130) );
  XOR U1131 ( .A(n1131), .B(n1132), .Z(SUM[491]) );
  XNOR U1132 ( .A(B[491]), .B(A[491]), .Z(n1132) );
  XOR U1133 ( .A(n1133), .B(n1134), .Z(SUM[490]) );
  XNOR U1134 ( .A(B[490]), .B(A[490]), .Z(n1134) );
  XOR U1135 ( .A(n1135), .B(n1136), .Z(SUM[48]) );
  XNOR U1136 ( .A(B[48]), .B(A[48]), .Z(n1136) );
  XOR U1137 ( .A(n1137), .B(n1138), .Z(SUM[489]) );
  XNOR U1138 ( .A(B[489]), .B(A[489]), .Z(n1138) );
  XOR U1139 ( .A(n1139), .B(n1140), .Z(SUM[488]) );
  XNOR U1140 ( .A(B[488]), .B(A[488]), .Z(n1140) );
  XOR U1141 ( .A(n1141), .B(n1142), .Z(SUM[487]) );
  XNOR U1142 ( .A(B[487]), .B(A[487]), .Z(n1142) );
  XOR U1143 ( .A(n1143), .B(n1144), .Z(SUM[486]) );
  XNOR U1144 ( .A(B[486]), .B(A[486]), .Z(n1144) );
  XOR U1145 ( .A(n1145), .B(n1146), .Z(SUM[485]) );
  XNOR U1146 ( .A(B[485]), .B(A[485]), .Z(n1146) );
  XOR U1147 ( .A(n1147), .B(n1148), .Z(SUM[484]) );
  XNOR U1148 ( .A(B[484]), .B(A[484]), .Z(n1148) );
  XOR U1149 ( .A(n1149), .B(n1150), .Z(SUM[483]) );
  XNOR U1150 ( .A(B[483]), .B(A[483]), .Z(n1150) );
  XOR U1151 ( .A(n1151), .B(n1152), .Z(SUM[482]) );
  XNOR U1152 ( .A(B[482]), .B(A[482]), .Z(n1152) );
  XOR U1153 ( .A(n1153), .B(n1154), .Z(SUM[481]) );
  XNOR U1154 ( .A(B[481]), .B(A[481]), .Z(n1154) );
  XOR U1155 ( .A(n1155), .B(n1156), .Z(SUM[480]) );
  XNOR U1156 ( .A(B[480]), .B(A[480]), .Z(n1156) );
  XOR U1157 ( .A(n1157), .B(n1158), .Z(SUM[47]) );
  XNOR U1158 ( .A(B[47]), .B(A[47]), .Z(n1158) );
  XOR U1159 ( .A(n1159), .B(n1160), .Z(SUM[479]) );
  XNOR U1160 ( .A(B[479]), .B(A[479]), .Z(n1160) );
  XOR U1161 ( .A(n1161), .B(n1162), .Z(SUM[478]) );
  XNOR U1162 ( .A(B[478]), .B(A[478]), .Z(n1162) );
  XOR U1163 ( .A(n1163), .B(n1164), .Z(SUM[477]) );
  XNOR U1164 ( .A(B[477]), .B(A[477]), .Z(n1164) );
  XOR U1165 ( .A(n1165), .B(n1166), .Z(SUM[476]) );
  XNOR U1166 ( .A(B[476]), .B(A[476]), .Z(n1166) );
  XOR U1167 ( .A(n1167), .B(n1168), .Z(SUM[475]) );
  XNOR U1168 ( .A(B[475]), .B(A[475]), .Z(n1168) );
  XOR U1169 ( .A(n1169), .B(n1170), .Z(SUM[474]) );
  XNOR U1170 ( .A(B[474]), .B(A[474]), .Z(n1170) );
  XOR U1171 ( .A(n1171), .B(n1172), .Z(SUM[473]) );
  XNOR U1172 ( .A(B[473]), .B(A[473]), .Z(n1172) );
  XOR U1173 ( .A(n1173), .B(n1174), .Z(SUM[472]) );
  XNOR U1174 ( .A(B[472]), .B(A[472]), .Z(n1174) );
  XOR U1175 ( .A(n1175), .B(n1176), .Z(SUM[471]) );
  XNOR U1176 ( .A(B[471]), .B(A[471]), .Z(n1176) );
  XOR U1177 ( .A(n1177), .B(n1178), .Z(SUM[470]) );
  XNOR U1178 ( .A(B[470]), .B(A[470]), .Z(n1178) );
  XOR U1179 ( .A(n1179), .B(n1180), .Z(SUM[46]) );
  XNOR U1180 ( .A(B[46]), .B(A[46]), .Z(n1180) );
  XOR U1181 ( .A(n1181), .B(n1182), .Z(SUM[469]) );
  XNOR U1182 ( .A(B[469]), .B(A[469]), .Z(n1182) );
  XOR U1183 ( .A(n1183), .B(n1184), .Z(SUM[468]) );
  XNOR U1184 ( .A(B[468]), .B(A[468]), .Z(n1184) );
  XOR U1185 ( .A(n1185), .B(n1186), .Z(SUM[467]) );
  XNOR U1186 ( .A(B[467]), .B(A[467]), .Z(n1186) );
  XOR U1187 ( .A(n1187), .B(n1188), .Z(SUM[466]) );
  XNOR U1188 ( .A(B[466]), .B(A[466]), .Z(n1188) );
  XOR U1189 ( .A(n1189), .B(n1190), .Z(SUM[465]) );
  XNOR U1190 ( .A(B[465]), .B(A[465]), .Z(n1190) );
  XOR U1191 ( .A(n1191), .B(n1192), .Z(SUM[464]) );
  XNOR U1192 ( .A(B[464]), .B(A[464]), .Z(n1192) );
  XOR U1193 ( .A(n1193), .B(n1194), .Z(SUM[463]) );
  XNOR U1194 ( .A(B[463]), .B(A[463]), .Z(n1194) );
  XOR U1195 ( .A(n1195), .B(n1196), .Z(SUM[462]) );
  XNOR U1196 ( .A(B[462]), .B(A[462]), .Z(n1196) );
  XOR U1197 ( .A(n1197), .B(n1198), .Z(SUM[461]) );
  XNOR U1198 ( .A(B[461]), .B(A[461]), .Z(n1198) );
  XOR U1199 ( .A(n1199), .B(n1200), .Z(SUM[460]) );
  XNOR U1200 ( .A(B[460]), .B(A[460]), .Z(n1200) );
  XOR U1201 ( .A(n1201), .B(n1202), .Z(SUM[45]) );
  XNOR U1202 ( .A(B[45]), .B(A[45]), .Z(n1202) );
  XOR U1203 ( .A(n1203), .B(n1204), .Z(SUM[459]) );
  XNOR U1204 ( .A(B[459]), .B(A[459]), .Z(n1204) );
  XOR U1205 ( .A(n1205), .B(n1206), .Z(SUM[458]) );
  XNOR U1206 ( .A(B[458]), .B(A[458]), .Z(n1206) );
  XOR U1207 ( .A(n1207), .B(n1208), .Z(SUM[457]) );
  XNOR U1208 ( .A(B[457]), .B(A[457]), .Z(n1208) );
  XOR U1209 ( .A(n1209), .B(n1210), .Z(SUM[456]) );
  XNOR U1210 ( .A(B[456]), .B(A[456]), .Z(n1210) );
  XOR U1211 ( .A(n1211), .B(n1212), .Z(SUM[455]) );
  XNOR U1212 ( .A(B[455]), .B(A[455]), .Z(n1212) );
  XOR U1213 ( .A(n1213), .B(n1214), .Z(SUM[454]) );
  XNOR U1214 ( .A(B[454]), .B(A[454]), .Z(n1214) );
  XOR U1215 ( .A(n1215), .B(n1216), .Z(SUM[453]) );
  XNOR U1216 ( .A(B[453]), .B(A[453]), .Z(n1216) );
  XOR U1217 ( .A(n1217), .B(n1218), .Z(SUM[452]) );
  XNOR U1218 ( .A(B[452]), .B(A[452]), .Z(n1218) );
  XOR U1219 ( .A(n1219), .B(n1220), .Z(SUM[451]) );
  XNOR U1220 ( .A(B[451]), .B(A[451]), .Z(n1220) );
  XOR U1221 ( .A(n1221), .B(n1222), .Z(SUM[450]) );
  XNOR U1222 ( .A(B[450]), .B(A[450]), .Z(n1222) );
  XOR U1223 ( .A(n1223), .B(n1224), .Z(SUM[44]) );
  XNOR U1224 ( .A(B[44]), .B(A[44]), .Z(n1224) );
  XOR U1225 ( .A(n1225), .B(n1226), .Z(SUM[449]) );
  XNOR U1226 ( .A(B[449]), .B(A[449]), .Z(n1226) );
  XOR U1227 ( .A(n1227), .B(n1228), .Z(SUM[448]) );
  XNOR U1228 ( .A(B[448]), .B(A[448]), .Z(n1228) );
  XOR U1229 ( .A(n1229), .B(n1230), .Z(SUM[447]) );
  XNOR U1230 ( .A(B[447]), .B(A[447]), .Z(n1230) );
  XOR U1231 ( .A(n1231), .B(n1232), .Z(SUM[446]) );
  XNOR U1232 ( .A(B[446]), .B(A[446]), .Z(n1232) );
  XOR U1233 ( .A(n1233), .B(n1234), .Z(SUM[445]) );
  XNOR U1234 ( .A(B[445]), .B(A[445]), .Z(n1234) );
  XOR U1235 ( .A(n1235), .B(n1236), .Z(SUM[444]) );
  XNOR U1236 ( .A(B[444]), .B(A[444]), .Z(n1236) );
  XOR U1237 ( .A(n1237), .B(n1238), .Z(SUM[443]) );
  XNOR U1238 ( .A(B[443]), .B(A[443]), .Z(n1238) );
  XOR U1239 ( .A(n1239), .B(n1240), .Z(SUM[442]) );
  XNOR U1240 ( .A(B[442]), .B(A[442]), .Z(n1240) );
  XOR U1241 ( .A(n1241), .B(n1242), .Z(SUM[441]) );
  XNOR U1242 ( .A(B[441]), .B(A[441]), .Z(n1242) );
  XOR U1243 ( .A(n1243), .B(n1244), .Z(SUM[440]) );
  XNOR U1244 ( .A(B[440]), .B(A[440]), .Z(n1244) );
  XOR U1245 ( .A(n1245), .B(n1246), .Z(SUM[43]) );
  XNOR U1246 ( .A(B[43]), .B(A[43]), .Z(n1246) );
  XOR U1247 ( .A(n1247), .B(n1248), .Z(SUM[439]) );
  XNOR U1248 ( .A(B[439]), .B(A[439]), .Z(n1248) );
  XOR U1249 ( .A(n1249), .B(n1250), .Z(SUM[438]) );
  XNOR U1250 ( .A(B[438]), .B(A[438]), .Z(n1250) );
  XOR U1251 ( .A(n1251), .B(n1252), .Z(SUM[437]) );
  XNOR U1252 ( .A(B[437]), .B(A[437]), .Z(n1252) );
  XOR U1253 ( .A(n1253), .B(n1254), .Z(SUM[436]) );
  XNOR U1254 ( .A(B[436]), .B(A[436]), .Z(n1254) );
  XOR U1255 ( .A(n1255), .B(n1256), .Z(SUM[435]) );
  XNOR U1256 ( .A(B[435]), .B(A[435]), .Z(n1256) );
  XOR U1257 ( .A(n1257), .B(n1258), .Z(SUM[434]) );
  XNOR U1258 ( .A(B[434]), .B(A[434]), .Z(n1258) );
  XOR U1259 ( .A(n1259), .B(n1260), .Z(SUM[433]) );
  XNOR U1260 ( .A(B[433]), .B(A[433]), .Z(n1260) );
  XOR U1261 ( .A(n1261), .B(n1262), .Z(SUM[432]) );
  XNOR U1262 ( .A(B[432]), .B(A[432]), .Z(n1262) );
  XOR U1263 ( .A(n1263), .B(n1264), .Z(SUM[431]) );
  XNOR U1264 ( .A(B[431]), .B(A[431]), .Z(n1264) );
  XOR U1265 ( .A(n1265), .B(n1266), .Z(SUM[430]) );
  XNOR U1266 ( .A(B[430]), .B(A[430]), .Z(n1266) );
  XOR U1267 ( .A(n1267), .B(n1268), .Z(SUM[42]) );
  XNOR U1268 ( .A(B[42]), .B(A[42]), .Z(n1268) );
  XOR U1269 ( .A(n1269), .B(n1270), .Z(SUM[429]) );
  XNOR U1270 ( .A(B[429]), .B(A[429]), .Z(n1270) );
  XOR U1271 ( .A(n1271), .B(n1272), .Z(SUM[428]) );
  XNOR U1272 ( .A(B[428]), .B(A[428]), .Z(n1272) );
  XOR U1273 ( .A(n1273), .B(n1274), .Z(SUM[427]) );
  XNOR U1274 ( .A(B[427]), .B(A[427]), .Z(n1274) );
  XOR U1275 ( .A(n1275), .B(n1276), .Z(SUM[426]) );
  XNOR U1276 ( .A(B[426]), .B(A[426]), .Z(n1276) );
  XOR U1277 ( .A(n1277), .B(n1278), .Z(SUM[425]) );
  XNOR U1278 ( .A(B[425]), .B(A[425]), .Z(n1278) );
  XOR U1279 ( .A(n1279), .B(n1280), .Z(SUM[424]) );
  XNOR U1280 ( .A(B[424]), .B(A[424]), .Z(n1280) );
  XOR U1281 ( .A(n1281), .B(n1282), .Z(SUM[423]) );
  XNOR U1282 ( .A(B[423]), .B(A[423]), .Z(n1282) );
  XOR U1283 ( .A(n1283), .B(n1284), .Z(SUM[422]) );
  XNOR U1284 ( .A(B[422]), .B(A[422]), .Z(n1284) );
  XOR U1285 ( .A(n1285), .B(n1286), .Z(SUM[421]) );
  XNOR U1286 ( .A(B[421]), .B(A[421]), .Z(n1286) );
  XOR U1287 ( .A(n1287), .B(n1288), .Z(SUM[420]) );
  XNOR U1288 ( .A(B[420]), .B(A[420]), .Z(n1288) );
  XOR U1289 ( .A(n1289), .B(n1290), .Z(SUM[41]) );
  XNOR U1290 ( .A(B[41]), .B(A[41]), .Z(n1290) );
  XOR U1291 ( .A(n1291), .B(n1292), .Z(SUM[419]) );
  XNOR U1292 ( .A(B[419]), .B(A[419]), .Z(n1292) );
  XOR U1293 ( .A(n1293), .B(n1294), .Z(SUM[418]) );
  XNOR U1294 ( .A(B[418]), .B(A[418]), .Z(n1294) );
  XOR U1295 ( .A(n1295), .B(n1296), .Z(SUM[417]) );
  XNOR U1296 ( .A(B[417]), .B(A[417]), .Z(n1296) );
  XOR U1297 ( .A(n1297), .B(n1298), .Z(SUM[416]) );
  XNOR U1298 ( .A(B[416]), .B(A[416]), .Z(n1298) );
  XOR U1299 ( .A(n1299), .B(n1300), .Z(SUM[415]) );
  XNOR U1300 ( .A(B[415]), .B(A[415]), .Z(n1300) );
  XOR U1301 ( .A(n1301), .B(n1302), .Z(SUM[414]) );
  XNOR U1302 ( .A(B[414]), .B(A[414]), .Z(n1302) );
  XOR U1303 ( .A(n1303), .B(n1304), .Z(SUM[413]) );
  XNOR U1304 ( .A(B[413]), .B(A[413]), .Z(n1304) );
  XOR U1305 ( .A(n1305), .B(n1306), .Z(SUM[412]) );
  XNOR U1306 ( .A(B[412]), .B(A[412]), .Z(n1306) );
  XOR U1307 ( .A(n1307), .B(n1308), .Z(SUM[411]) );
  XNOR U1308 ( .A(B[411]), .B(A[411]), .Z(n1308) );
  XOR U1309 ( .A(n1309), .B(n1310), .Z(SUM[410]) );
  XNOR U1310 ( .A(B[410]), .B(A[410]), .Z(n1310) );
  XOR U1311 ( .A(n1311), .B(n1312), .Z(SUM[40]) );
  XNOR U1312 ( .A(B[40]), .B(A[40]), .Z(n1312) );
  XOR U1313 ( .A(n1313), .B(n1314), .Z(SUM[409]) );
  XNOR U1314 ( .A(B[409]), .B(A[409]), .Z(n1314) );
  XOR U1315 ( .A(n1315), .B(n1316), .Z(SUM[408]) );
  XNOR U1316 ( .A(B[408]), .B(A[408]), .Z(n1316) );
  XOR U1317 ( .A(n1317), .B(n1318), .Z(SUM[407]) );
  XNOR U1318 ( .A(B[407]), .B(A[407]), .Z(n1318) );
  XOR U1319 ( .A(n1319), .B(n1320), .Z(SUM[406]) );
  XNOR U1320 ( .A(B[406]), .B(A[406]), .Z(n1320) );
  XOR U1321 ( .A(n1321), .B(n1322), .Z(SUM[405]) );
  XNOR U1322 ( .A(B[405]), .B(A[405]), .Z(n1322) );
  XOR U1323 ( .A(n1323), .B(n1324), .Z(SUM[404]) );
  XNOR U1324 ( .A(B[404]), .B(A[404]), .Z(n1324) );
  XOR U1325 ( .A(n1325), .B(n1326), .Z(SUM[403]) );
  XNOR U1326 ( .A(B[403]), .B(A[403]), .Z(n1326) );
  XOR U1327 ( .A(n1327), .B(n1328), .Z(SUM[402]) );
  XNOR U1328 ( .A(B[402]), .B(A[402]), .Z(n1328) );
  XOR U1329 ( .A(n1329), .B(n1330), .Z(SUM[401]) );
  XNOR U1330 ( .A(B[401]), .B(A[401]), .Z(n1330) );
  XOR U1331 ( .A(n1331), .B(n1332), .Z(SUM[400]) );
  XNOR U1332 ( .A(B[400]), .B(A[400]), .Z(n1332) );
  XOR U1333 ( .A(n1333), .B(n1334), .Z(SUM[3]) );
  XNOR U1334 ( .A(B[3]), .B(A[3]), .Z(n1334) );
  XOR U1335 ( .A(n1335), .B(n1336), .Z(SUM[39]) );
  XNOR U1336 ( .A(B[39]), .B(A[39]), .Z(n1336) );
  XOR U1337 ( .A(n1337), .B(n1338), .Z(SUM[399]) );
  XNOR U1338 ( .A(B[399]), .B(A[399]), .Z(n1338) );
  XOR U1339 ( .A(n1339), .B(n1340), .Z(SUM[398]) );
  XNOR U1340 ( .A(B[398]), .B(A[398]), .Z(n1340) );
  XOR U1341 ( .A(n1341), .B(n1342), .Z(SUM[397]) );
  XNOR U1342 ( .A(B[397]), .B(A[397]), .Z(n1342) );
  XOR U1343 ( .A(n1343), .B(n1344), .Z(SUM[396]) );
  XNOR U1344 ( .A(B[396]), .B(A[396]), .Z(n1344) );
  XOR U1345 ( .A(n1345), .B(n1346), .Z(SUM[395]) );
  XNOR U1346 ( .A(B[395]), .B(A[395]), .Z(n1346) );
  XOR U1347 ( .A(n1347), .B(n1348), .Z(SUM[394]) );
  XNOR U1348 ( .A(B[394]), .B(A[394]), .Z(n1348) );
  XOR U1349 ( .A(n1349), .B(n1350), .Z(SUM[393]) );
  XNOR U1350 ( .A(B[393]), .B(A[393]), .Z(n1350) );
  XOR U1351 ( .A(n1351), .B(n1352), .Z(SUM[392]) );
  XNOR U1352 ( .A(B[392]), .B(A[392]), .Z(n1352) );
  XOR U1353 ( .A(n1353), .B(n1354), .Z(SUM[391]) );
  XNOR U1354 ( .A(B[391]), .B(A[391]), .Z(n1354) );
  XOR U1355 ( .A(n1355), .B(n1356), .Z(SUM[390]) );
  XNOR U1356 ( .A(B[390]), .B(A[390]), .Z(n1356) );
  XOR U1357 ( .A(n1357), .B(n1358), .Z(SUM[38]) );
  XNOR U1358 ( .A(B[38]), .B(A[38]), .Z(n1358) );
  XOR U1359 ( .A(n1359), .B(n1360), .Z(SUM[389]) );
  XNOR U1360 ( .A(B[389]), .B(A[389]), .Z(n1360) );
  XOR U1361 ( .A(n1361), .B(n1362), .Z(SUM[388]) );
  XNOR U1362 ( .A(B[388]), .B(A[388]), .Z(n1362) );
  XOR U1363 ( .A(n1363), .B(n1364), .Z(SUM[387]) );
  XNOR U1364 ( .A(B[387]), .B(A[387]), .Z(n1364) );
  XOR U1365 ( .A(n1365), .B(n1366), .Z(SUM[386]) );
  XNOR U1366 ( .A(B[386]), .B(A[386]), .Z(n1366) );
  XOR U1367 ( .A(n1367), .B(n1368), .Z(SUM[385]) );
  XNOR U1368 ( .A(B[385]), .B(A[385]), .Z(n1368) );
  XOR U1369 ( .A(n1369), .B(n1370), .Z(SUM[384]) );
  XNOR U1370 ( .A(B[384]), .B(A[384]), .Z(n1370) );
  XOR U1371 ( .A(n1371), .B(n1372), .Z(SUM[383]) );
  XNOR U1372 ( .A(B[383]), .B(A[383]), .Z(n1372) );
  XOR U1373 ( .A(n1373), .B(n1374), .Z(SUM[382]) );
  XNOR U1374 ( .A(B[382]), .B(A[382]), .Z(n1374) );
  XOR U1375 ( .A(n1375), .B(n1376), .Z(SUM[381]) );
  XNOR U1376 ( .A(B[381]), .B(A[381]), .Z(n1376) );
  XOR U1377 ( .A(n1377), .B(n1378), .Z(SUM[380]) );
  XNOR U1378 ( .A(B[380]), .B(A[380]), .Z(n1378) );
  XOR U1379 ( .A(n1379), .B(n1380), .Z(SUM[37]) );
  XNOR U1380 ( .A(B[37]), .B(A[37]), .Z(n1380) );
  XOR U1381 ( .A(n1381), .B(n1382), .Z(SUM[379]) );
  XNOR U1382 ( .A(B[379]), .B(A[379]), .Z(n1382) );
  XOR U1383 ( .A(n1383), .B(n1384), .Z(SUM[378]) );
  XNOR U1384 ( .A(B[378]), .B(A[378]), .Z(n1384) );
  XOR U1385 ( .A(n1385), .B(n1386), .Z(SUM[377]) );
  XNOR U1386 ( .A(B[377]), .B(A[377]), .Z(n1386) );
  XOR U1387 ( .A(n1387), .B(n1388), .Z(SUM[376]) );
  XNOR U1388 ( .A(B[376]), .B(A[376]), .Z(n1388) );
  XOR U1389 ( .A(n1389), .B(n1390), .Z(SUM[375]) );
  XNOR U1390 ( .A(B[375]), .B(A[375]), .Z(n1390) );
  XOR U1391 ( .A(n1391), .B(n1392), .Z(SUM[374]) );
  XNOR U1392 ( .A(B[374]), .B(A[374]), .Z(n1392) );
  XOR U1393 ( .A(n1393), .B(n1394), .Z(SUM[373]) );
  XNOR U1394 ( .A(B[373]), .B(A[373]), .Z(n1394) );
  XOR U1395 ( .A(n1395), .B(n1396), .Z(SUM[372]) );
  XNOR U1396 ( .A(B[372]), .B(A[372]), .Z(n1396) );
  XOR U1397 ( .A(n1397), .B(n1398), .Z(SUM[371]) );
  XNOR U1398 ( .A(B[371]), .B(A[371]), .Z(n1398) );
  XOR U1399 ( .A(n1399), .B(n1400), .Z(SUM[370]) );
  XNOR U1400 ( .A(B[370]), .B(A[370]), .Z(n1400) );
  XOR U1401 ( .A(n1401), .B(n1402), .Z(SUM[36]) );
  XNOR U1402 ( .A(B[36]), .B(A[36]), .Z(n1402) );
  XOR U1403 ( .A(n1403), .B(n1404), .Z(SUM[369]) );
  XNOR U1404 ( .A(B[369]), .B(A[369]), .Z(n1404) );
  XOR U1405 ( .A(n1405), .B(n1406), .Z(SUM[368]) );
  XNOR U1406 ( .A(B[368]), .B(A[368]), .Z(n1406) );
  XOR U1407 ( .A(n1407), .B(n1408), .Z(SUM[367]) );
  XNOR U1408 ( .A(B[367]), .B(A[367]), .Z(n1408) );
  XOR U1409 ( .A(n1409), .B(n1410), .Z(SUM[366]) );
  XNOR U1410 ( .A(B[366]), .B(A[366]), .Z(n1410) );
  XOR U1411 ( .A(n1411), .B(n1412), .Z(SUM[365]) );
  XNOR U1412 ( .A(B[365]), .B(A[365]), .Z(n1412) );
  XOR U1413 ( .A(n1413), .B(n1414), .Z(SUM[364]) );
  XNOR U1414 ( .A(B[364]), .B(A[364]), .Z(n1414) );
  XOR U1415 ( .A(n1415), .B(n1416), .Z(SUM[363]) );
  XNOR U1416 ( .A(B[363]), .B(A[363]), .Z(n1416) );
  XOR U1417 ( .A(n1417), .B(n1418), .Z(SUM[362]) );
  XNOR U1418 ( .A(B[362]), .B(A[362]), .Z(n1418) );
  XOR U1419 ( .A(n1419), .B(n1420), .Z(SUM[361]) );
  XNOR U1420 ( .A(B[361]), .B(A[361]), .Z(n1420) );
  XOR U1421 ( .A(n1421), .B(n1422), .Z(SUM[360]) );
  XNOR U1422 ( .A(B[360]), .B(A[360]), .Z(n1422) );
  XOR U1423 ( .A(n1423), .B(n1424), .Z(SUM[35]) );
  XNOR U1424 ( .A(B[35]), .B(A[35]), .Z(n1424) );
  XOR U1425 ( .A(n1425), .B(n1426), .Z(SUM[359]) );
  XNOR U1426 ( .A(B[359]), .B(A[359]), .Z(n1426) );
  XOR U1427 ( .A(n1427), .B(n1428), .Z(SUM[358]) );
  XNOR U1428 ( .A(B[358]), .B(A[358]), .Z(n1428) );
  XOR U1429 ( .A(n1429), .B(n1430), .Z(SUM[357]) );
  XNOR U1430 ( .A(B[357]), .B(A[357]), .Z(n1430) );
  XOR U1431 ( .A(n1431), .B(n1432), .Z(SUM[356]) );
  XNOR U1432 ( .A(B[356]), .B(A[356]), .Z(n1432) );
  XOR U1433 ( .A(n1433), .B(n1434), .Z(SUM[355]) );
  XNOR U1434 ( .A(B[355]), .B(A[355]), .Z(n1434) );
  XOR U1435 ( .A(n1435), .B(n1436), .Z(SUM[354]) );
  XNOR U1436 ( .A(B[354]), .B(A[354]), .Z(n1436) );
  XOR U1437 ( .A(n1437), .B(n1438), .Z(SUM[353]) );
  XNOR U1438 ( .A(B[353]), .B(A[353]), .Z(n1438) );
  XOR U1439 ( .A(n1439), .B(n1440), .Z(SUM[352]) );
  XNOR U1440 ( .A(B[352]), .B(A[352]), .Z(n1440) );
  XOR U1441 ( .A(n1441), .B(n1442), .Z(SUM[351]) );
  XNOR U1442 ( .A(B[351]), .B(A[351]), .Z(n1442) );
  XOR U1443 ( .A(n1443), .B(n1444), .Z(SUM[350]) );
  XNOR U1444 ( .A(B[350]), .B(A[350]), .Z(n1444) );
  XOR U1445 ( .A(n1445), .B(n1446), .Z(SUM[34]) );
  XNOR U1446 ( .A(B[34]), .B(A[34]), .Z(n1446) );
  XOR U1447 ( .A(n1447), .B(n1448), .Z(SUM[349]) );
  XNOR U1448 ( .A(B[349]), .B(A[349]), .Z(n1448) );
  XOR U1449 ( .A(n1449), .B(n1450), .Z(SUM[348]) );
  XNOR U1450 ( .A(B[348]), .B(A[348]), .Z(n1450) );
  XOR U1451 ( .A(n1451), .B(n1452), .Z(SUM[347]) );
  XNOR U1452 ( .A(B[347]), .B(A[347]), .Z(n1452) );
  XOR U1453 ( .A(n1453), .B(n1454), .Z(SUM[346]) );
  XNOR U1454 ( .A(B[346]), .B(A[346]), .Z(n1454) );
  XOR U1455 ( .A(n1455), .B(n1456), .Z(SUM[345]) );
  XNOR U1456 ( .A(B[345]), .B(A[345]), .Z(n1456) );
  XOR U1457 ( .A(n1457), .B(n1458), .Z(SUM[344]) );
  XNOR U1458 ( .A(B[344]), .B(A[344]), .Z(n1458) );
  XOR U1459 ( .A(n1459), .B(n1460), .Z(SUM[343]) );
  XNOR U1460 ( .A(B[343]), .B(A[343]), .Z(n1460) );
  XOR U1461 ( .A(n1461), .B(n1462), .Z(SUM[342]) );
  XNOR U1462 ( .A(B[342]), .B(A[342]), .Z(n1462) );
  XOR U1463 ( .A(n1463), .B(n1464), .Z(SUM[341]) );
  XNOR U1464 ( .A(B[341]), .B(A[341]), .Z(n1464) );
  XOR U1465 ( .A(n1465), .B(n1466), .Z(SUM[340]) );
  XNOR U1466 ( .A(B[340]), .B(A[340]), .Z(n1466) );
  XOR U1467 ( .A(n1467), .B(n1468), .Z(SUM[33]) );
  XNOR U1468 ( .A(B[33]), .B(A[33]), .Z(n1468) );
  XOR U1469 ( .A(n1469), .B(n1470), .Z(SUM[339]) );
  XNOR U1470 ( .A(B[339]), .B(A[339]), .Z(n1470) );
  XOR U1471 ( .A(n1471), .B(n1472), .Z(SUM[338]) );
  XNOR U1472 ( .A(B[338]), .B(A[338]), .Z(n1472) );
  XOR U1473 ( .A(n1473), .B(n1474), .Z(SUM[337]) );
  XNOR U1474 ( .A(B[337]), .B(A[337]), .Z(n1474) );
  XOR U1475 ( .A(n1475), .B(n1476), .Z(SUM[336]) );
  XNOR U1476 ( .A(B[336]), .B(A[336]), .Z(n1476) );
  XOR U1477 ( .A(n1477), .B(n1478), .Z(SUM[335]) );
  XNOR U1478 ( .A(B[335]), .B(A[335]), .Z(n1478) );
  XOR U1479 ( .A(n1479), .B(n1480), .Z(SUM[334]) );
  XNOR U1480 ( .A(B[334]), .B(A[334]), .Z(n1480) );
  XOR U1481 ( .A(n1481), .B(n1482), .Z(SUM[333]) );
  XNOR U1482 ( .A(B[333]), .B(A[333]), .Z(n1482) );
  XOR U1483 ( .A(n1483), .B(n1484), .Z(SUM[332]) );
  XNOR U1484 ( .A(B[332]), .B(A[332]), .Z(n1484) );
  XOR U1485 ( .A(n1485), .B(n1486), .Z(SUM[331]) );
  XNOR U1486 ( .A(B[331]), .B(A[331]), .Z(n1486) );
  XOR U1487 ( .A(n1487), .B(n1488), .Z(SUM[330]) );
  XNOR U1488 ( .A(B[330]), .B(A[330]), .Z(n1488) );
  XOR U1489 ( .A(n1489), .B(n1490), .Z(SUM[32]) );
  XNOR U1490 ( .A(B[32]), .B(A[32]), .Z(n1490) );
  XOR U1491 ( .A(n1491), .B(n1492), .Z(SUM[329]) );
  XNOR U1492 ( .A(B[329]), .B(A[329]), .Z(n1492) );
  XOR U1493 ( .A(n1493), .B(n1494), .Z(SUM[328]) );
  XNOR U1494 ( .A(B[328]), .B(A[328]), .Z(n1494) );
  XOR U1495 ( .A(n1495), .B(n1496), .Z(SUM[327]) );
  XNOR U1496 ( .A(B[327]), .B(A[327]), .Z(n1496) );
  XOR U1497 ( .A(n1497), .B(n1498), .Z(SUM[326]) );
  XNOR U1498 ( .A(B[326]), .B(A[326]), .Z(n1498) );
  XOR U1499 ( .A(n1499), .B(n1500), .Z(SUM[325]) );
  XNOR U1500 ( .A(B[325]), .B(A[325]), .Z(n1500) );
  XOR U1501 ( .A(n1501), .B(n1502), .Z(SUM[324]) );
  XNOR U1502 ( .A(B[324]), .B(A[324]), .Z(n1502) );
  XOR U1503 ( .A(n1503), .B(n1504), .Z(SUM[323]) );
  XNOR U1504 ( .A(B[323]), .B(A[323]), .Z(n1504) );
  XOR U1505 ( .A(n1505), .B(n1506), .Z(SUM[322]) );
  XNOR U1506 ( .A(B[322]), .B(A[322]), .Z(n1506) );
  XOR U1507 ( .A(n1507), .B(n1508), .Z(SUM[321]) );
  XNOR U1508 ( .A(B[321]), .B(A[321]), .Z(n1508) );
  XOR U1509 ( .A(n1509), .B(n1510), .Z(SUM[320]) );
  XNOR U1510 ( .A(B[320]), .B(A[320]), .Z(n1510) );
  XOR U1511 ( .A(n1511), .B(n1512), .Z(SUM[31]) );
  XNOR U1512 ( .A(B[31]), .B(A[31]), .Z(n1512) );
  XOR U1513 ( .A(n1513), .B(n1514), .Z(SUM[319]) );
  XNOR U1514 ( .A(B[319]), .B(A[319]), .Z(n1514) );
  XOR U1515 ( .A(n1515), .B(n1516), .Z(SUM[318]) );
  XNOR U1516 ( .A(B[318]), .B(A[318]), .Z(n1516) );
  XOR U1517 ( .A(n1517), .B(n1518), .Z(SUM[317]) );
  XNOR U1518 ( .A(B[317]), .B(A[317]), .Z(n1518) );
  XOR U1519 ( .A(n1519), .B(n1520), .Z(SUM[316]) );
  XNOR U1520 ( .A(B[316]), .B(A[316]), .Z(n1520) );
  XOR U1521 ( .A(n1521), .B(n1522), .Z(SUM[315]) );
  XNOR U1522 ( .A(B[315]), .B(A[315]), .Z(n1522) );
  XOR U1523 ( .A(n1523), .B(n1524), .Z(SUM[314]) );
  XNOR U1524 ( .A(B[314]), .B(A[314]), .Z(n1524) );
  XOR U1525 ( .A(n1525), .B(n1526), .Z(SUM[313]) );
  XNOR U1526 ( .A(B[313]), .B(A[313]), .Z(n1526) );
  XOR U1527 ( .A(n1527), .B(n1528), .Z(SUM[312]) );
  XNOR U1528 ( .A(B[312]), .B(A[312]), .Z(n1528) );
  XOR U1529 ( .A(n1529), .B(n1530), .Z(SUM[311]) );
  XNOR U1530 ( .A(B[311]), .B(A[311]), .Z(n1530) );
  XOR U1531 ( .A(n1531), .B(n1532), .Z(SUM[310]) );
  XNOR U1532 ( .A(B[310]), .B(A[310]), .Z(n1532) );
  XOR U1533 ( .A(n1533), .B(n1534), .Z(SUM[30]) );
  XNOR U1534 ( .A(B[30]), .B(A[30]), .Z(n1534) );
  XOR U1535 ( .A(n1535), .B(n1536), .Z(SUM[309]) );
  XNOR U1536 ( .A(B[309]), .B(A[309]), .Z(n1536) );
  XOR U1537 ( .A(n1537), .B(n1538), .Z(SUM[308]) );
  XNOR U1538 ( .A(B[308]), .B(A[308]), .Z(n1538) );
  XOR U1539 ( .A(n1539), .B(n1540), .Z(SUM[307]) );
  XNOR U1540 ( .A(B[307]), .B(A[307]), .Z(n1540) );
  XOR U1541 ( .A(n1541), .B(n1542), .Z(SUM[306]) );
  XNOR U1542 ( .A(B[306]), .B(A[306]), .Z(n1542) );
  XOR U1543 ( .A(n1543), .B(n1544), .Z(SUM[305]) );
  XNOR U1544 ( .A(B[305]), .B(A[305]), .Z(n1544) );
  XOR U1545 ( .A(n1545), .B(n1546), .Z(SUM[304]) );
  XNOR U1546 ( .A(B[304]), .B(A[304]), .Z(n1546) );
  XOR U1547 ( .A(n1547), .B(n1548), .Z(SUM[303]) );
  XNOR U1548 ( .A(B[303]), .B(A[303]), .Z(n1548) );
  XOR U1549 ( .A(n1549), .B(n1550), .Z(SUM[302]) );
  XNOR U1550 ( .A(B[302]), .B(A[302]), .Z(n1550) );
  XOR U1551 ( .A(n1551), .B(n1552), .Z(SUM[301]) );
  XNOR U1552 ( .A(B[301]), .B(A[301]), .Z(n1552) );
  XOR U1553 ( .A(n1553), .B(n1554), .Z(SUM[300]) );
  XNOR U1554 ( .A(B[300]), .B(A[300]), .Z(n1554) );
  XOR U1555 ( .A(n1555), .B(n1556), .Z(SUM[2]) );
  XOR U1556 ( .A(B[2]), .B(A[2]), .Z(n1556) );
  XOR U1557 ( .A(n1557), .B(n1558), .Z(SUM[29]) );
  XNOR U1558 ( .A(B[29]), .B(A[29]), .Z(n1558) );
  XOR U1559 ( .A(n1559), .B(n1560), .Z(SUM[299]) );
  XNOR U1560 ( .A(B[299]), .B(A[299]), .Z(n1560) );
  XOR U1561 ( .A(n1561), .B(n1562), .Z(SUM[298]) );
  XNOR U1562 ( .A(B[298]), .B(A[298]), .Z(n1562) );
  XOR U1563 ( .A(n1563), .B(n1564), .Z(SUM[297]) );
  XNOR U1564 ( .A(B[297]), .B(A[297]), .Z(n1564) );
  XOR U1565 ( .A(n1565), .B(n1566), .Z(SUM[296]) );
  XNOR U1566 ( .A(B[296]), .B(A[296]), .Z(n1566) );
  XOR U1567 ( .A(n1567), .B(n1568), .Z(SUM[295]) );
  XNOR U1568 ( .A(B[295]), .B(A[295]), .Z(n1568) );
  XOR U1569 ( .A(n1569), .B(n1570), .Z(SUM[294]) );
  XNOR U1570 ( .A(B[294]), .B(A[294]), .Z(n1570) );
  XOR U1571 ( .A(n1571), .B(n1572), .Z(SUM[293]) );
  XNOR U1572 ( .A(B[293]), .B(A[293]), .Z(n1572) );
  XOR U1573 ( .A(n1573), .B(n1574), .Z(SUM[292]) );
  XNOR U1574 ( .A(B[292]), .B(A[292]), .Z(n1574) );
  XOR U1575 ( .A(n1575), .B(n1576), .Z(SUM[291]) );
  XNOR U1576 ( .A(B[291]), .B(A[291]), .Z(n1576) );
  XOR U1577 ( .A(n1577), .B(n1578), .Z(SUM[290]) );
  XNOR U1578 ( .A(B[290]), .B(A[290]), .Z(n1578) );
  XOR U1579 ( .A(n1579), .B(n1580), .Z(SUM[28]) );
  XNOR U1580 ( .A(B[28]), .B(A[28]), .Z(n1580) );
  XOR U1581 ( .A(n1581), .B(n1582), .Z(SUM[289]) );
  XNOR U1582 ( .A(B[289]), .B(A[289]), .Z(n1582) );
  XOR U1583 ( .A(n1583), .B(n1584), .Z(SUM[288]) );
  XNOR U1584 ( .A(B[288]), .B(A[288]), .Z(n1584) );
  XOR U1585 ( .A(n1585), .B(n1586), .Z(SUM[287]) );
  XNOR U1586 ( .A(B[287]), .B(A[287]), .Z(n1586) );
  XOR U1587 ( .A(n1587), .B(n1588), .Z(SUM[286]) );
  XNOR U1588 ( .A(B[286]), .B(A[286]), .Z(n1588) );
  XOR U1589 ( .A(n1589), .B(n1590), .Z(SUM[285]) );
  XNOR U1590 ( .A(B[285]), .B(A[285]), .Z(n1590) );
  XOR U1591 ( .A(n1591), .B(n1592), .Z(SUM[284]) );
  XNOR U1592 ( .A(B[284]), .B(A[284]), .Z(n1592) );
  XOR U1593 ( .A(n1593), .B(n1594), .Z(SUM[283]) );
  XNOR U1594 ( .A(B[283]), .B(A[283]), .Z(n1594) );
  XOR U1595 ( .A(n1595), .B(n1596), .Z(SUM[282]) );
  XNOR U1596 ( .A(B[282]), .B(A[282]), .Z(n1596) );
  XOR U1597 ( .A(n1597), .B(n1598), .Z(SUM[281]) );
  XNOR U1598 ( .A(B[281]), .B(A[281]), .Z(n1598) );
  XOR U1599 ( .A(n1599), .B(n1600), .Z(SUM[280]) );
  XNOR U1600 ( .A(B[280]), .B(A[280]), .Z(n1600) );
  XOR U1601 ( .A(n1601), .B(n1602), .Z(SUM[27]) );
  XNOR U1602 ( .A(B[27]), .B(A[27]), .Z(n1602) );
  XOR U1603 ( .A(n1603), .B(n1604), .Z(SUM[279]) );
  XNOR U1604 ( .A(B[279]), .B(A[279]), .Z(n1604) );
  XOR U1605 ( .A(n1605), .B(n1606), .Z(SUM[278]) );
  XNOR U1606 ( .A(B[278]), .B(A[278]), .Z(n1606) );
  XOR U1607 ( .A(n1607), .B(n1608), .Z(SUM[277]) );
  XNOR U1608 ( .A(B[277]), .B(A[277]), .Z(n1608) );
  XOR U1609 ( .A(n1609), .B(n1610), .Z(SUM[276]) );
  XNOR U1610 ( .A(B[276]), .B(A[276]), .Z(n1610) );
  XOR U1611 ( .A(n1611), .B(n1612), .Z(SUM[275]) );
  XNOR U1612 ( .A(B[275]), .B(A[275]), .Z(n1612) );
  XOR U1613 ( .A(n1613), .B(n1614), .Z(SUM[274]) );
  XNOR U1614 ( .A(B[274]), .B(A[274]), .Z(n1614) );
  XOR U1615 ( .A(n1615), .B(n1616), .Z(SUM[273]) );
  XNOR U1616 ( .A(B[273]), .B(A[273]), .Z(n1616) );
  XOR U1617 ( .A(n1617), .B(n1618), .Z(SUM[272]) );
  XNOR U1618 ( .A(B[272]), .B(A[272]), .Z(n1618) );
  XOR U1619 ( .A(n1619), .B(n1620), .Z(SUM[271]) );
  XNOR U1620 ( .A(B[271]), .B(A[271]), .Z(n1620) );
  XOR U1621 ( .A(n1621), .B(n1622), .Z(SUM[270]) );
  XNOR U1622 ( .A(B[270]), .B(A[270]), .Z(n1622) );
  XOR U1623 ( .A(n1623), .B(n1624), .Z(SUM[26]) );
  XNOR U1624 ( .A(B[26]), .B(A[26]), .Z(n1624) );
  XOR U1625 ( .A(n1625), .B(n1626), .Z(SUM[269]) );
  XNOR U1626 ( .A(B[269]), .B(A[269]), .Z(n1626) );
  XOR U1627 ( .A(n1627), .B(n1628), .Z(SUM[268]) );
  XNOR U1628 ( .A(B[268]), .B(A[268]), .Z(n1628) );
  XOR U1629 ( .A(n1629), .B(n1630), .Z(SUM[267]) );
  XNOR U1630 ( .A(B[267]), .B(A[267]), .Z(n1630) );
  XOR U1631 ( .A(n1631), .B(n1632), .Z(SUM[266]) );
  XNOR U1632 ( .A(B[266]), .B(A[266]), .Z(n1632) );
  XOR U1633 ( .A(n1633), .B(n1634), .Z(SUM[265]) );
  XNOR U1634 ( .A(B[265]), .B(A[265]), .Z(n1634) );
  XOR U1635 ( .A(n1635), .B(n1636), .Z(SUM[264]) );
  XNOR U1636 ( .A(B[264]), .B(A[264]), .Z(n1636) );
  XOR U1637 ( .A(n1637), .B(n1638), .Z(SUM[263]) );
  XNOR U1638 ( .A(B[263]), .B(A[263]), .Z(n1638) );
  XOR U1639 ( .A(n1639), .B(n1640), .Z(SUM[262]) );
  XNOR U1640 ( .A(B[262]), .B(A[262]), .Z(n1640) );
  XOR U1641 ( .A(n1641), .B(n1642), .Z(SUM[261]) );
  XNOR U1642 ( .A(B[261]), .B(A[261]), .Z(n1642) );
  XOR U1643 ( .A(n1643), .B(n1644), .Z(SUM[260]) );
  XNOR U1644 ( .A(B[260]), .B(A[260]), .Z(n1644) );
  XOR U1645 ( .A(n1645), .B(n1646), .Z(SUM[25]) );
  XNOR U1646 ( .A(B[25]), .B(A[25]), .Z(n1646) );
  XOR U1647 ( .A(n1647), .B(n1648), .Z(SUM[259]) );
  XNOR U1648 ( .A(B[259]), .B(A[259]), .Z(n1648) );
  XOR U1649 ( .A(n1649), .B(n1650), .Z(SUM[258]) );
  XNOR U1650 ( .A(B[258]), .B(A[258]), .Z(n1650) );
  XOR U1651 ( .A(n1651), .B(n1652), .Z(SUM[257]) );
  XNOR U1652 ( .A(B[257]), .B(A[257]), .Z(n1652) );
  XOR U1653 ( .A(n1653), .B(n1654), .Z(SUM[256]) );
  XNOR U1654 ( .A(B[256]), .B(A[256]), .Z(n1654) );
  XOR U1655 ( .A(n1655), .B(n1656), .Z(SUM[255]) );
  XNOR U1656 ( .A(B[255]), .B(A[255]), .Z(n1656) );
  XOR U1657 ( .A(n1657), .B(n1658), .Z(SUM[254]) );
  XNOR U1658 ( .A(B[254]), .B(A[254]), .Z(n1658) );
  XOR U1659 ( .A(n1659), .B(n1660), .Z(SUM[253]) );
  XNOR U1660 ( .A(B[253]), .B(A[253]), .Z(n1660) );
  XOR U1661 ( .A(n1661), .B(n1662), .Z(SUM[252]) );
  XNOR U1662 ( .A(B[252]), .B(A[252]), .Z(n1662) );
  XOR U1663 ( .A(n1663), .B(n1664), .Z(SUM[251]) );
  XNOR U1664 ( .A(B[251]), .B(A[251]), .Z(n1664) );
  XOR U1665 ( .A(n1665), .B(n1666), .Z(SUM[250]) );
  XNOR U1666 ( .A(B[250]), .B(A[250]), .Z(n1666) );
  XOR U1667 ( .A(n1667), .B(n1668), .Z(SUM[24]) );
  XNOR U1668 ( .A(B[24]), .B(A[24]), .Z(n1668) );
  XOR U1669 ( .A(n1669), .B(n1670), .Z(SUM[249]) );
  XNOR U1670 ( .A(B[249]), .B(A[249]), .Z(n1670) );
  XOR U1671 ( .A(n1671), .B(n1672), .Z(SUM[248]) );
  XNOR U1672 ( .A(B[248]), .B(A[248]), .Z(n1672) );
  XOR U1673 ( .A(n1673), .B(n1674), .Z(SUM[247]) );
  XNOR U1674 ( .A(B[247]), .B(A[247]), .Z(n1674) );
  XOR U1675 ( .A(n1675), .B(n1676), .Z(SUM[246]) );
  XNOR U1676 ( .A(B[246]), .B(A[246]), .Z(n1676) );
  XOR U1677 ( .A(n1677), .B(n1678), .Z(SUM[245]) );
  XNOR U1678 ( .A(B[245]), .B(A[245]), .Z(n1678) );
  XOR U1679 ( .A(n1679), .B(n1680), .Z(SUM[244]) );
  XNOR U1680 ( .A(B[244]), .B(A[244]), .Z(n1680) );
  XOR U1681 ( .A(n1681), .B(n1682), .Z(SUM[243]) );
  XNOR U1682 ( .A(B[243]), .B(A[243]), .Z(n1682) );
  XOR U1683 ( .A(n1683), .B(n1684), .Z(SUM[242]) );
  XNOR U1684 ( .A(B[242]), .B(A[242]), .Z(n1684) );
  XOR U1685 ( .A(n1685), .B(n1686), .Z(SUM[241]) );
  XNOR U1686 ( .A(B[241]), .B(A[241]), .Z(n1686) );
  XOR U1687 ( .A(n1687), .B(n1688), .Z(SUM[240]) );
  XNOR U1688 ( .A(B[240]), .B(A[240]), .Z(n1688) );
  XOR U1689 ( .A(n1689), .B(n1690), .Z(SUM[23]) );
  XNOR U1690 ( .A(B[23]), .B(A[23]), .Z(n1690) );
  XOR U1691 ( .A(n1691), .B(n1692), .Z(SUM[239]) );
  XNOR U1692 ( .A(B[239]), .B(A[239]), .Z(n1692) );
  XOR U1693 ( .A(n1693), .B(n1694), .Z(SUM[238]) );
  XNOR U1694 ( .A(B[238]), .B(A[238]), .Z(n1694) );
  XOR U1695 ( .A(n1695), .B(n1696), .Z(SUM[237]) );
  XNOR U1696 ( .A(B[237]), .B(A[237]), .Z(n1696) );
  XOR U1697 ( .A(n1697), .B(n1698), .Z(SUM[236]) );
  XNOR U1698 ( .A(B[236]), .B(A[236]), .Z(n1698) );
  XOR U1699 ( .A(n1699), .B(n1700), .Z(SUM[235]) );
  XNOR U1700 ( .A(B[235]), .B(A[235]), .Z(n1700) );
  XOR U1701 ( .A(n1701), .B(n1702), .Z(SUM[234]) );
  XNOR U1702 ( .A(B[234]), .B(A[234]), .Z(n1702) );
  XOR U1703 ( .A(n1703), .B(n1704), .Z(SUM[233]) );
  XNOR U1704 ( .A(B[233]), .B(A[233]), .Z(n1704) );
  XOR U1705 ( .A(n1705), .B(n1706), .Z(SUM[232]) );
  XNOR U1706 ( .A(B[232]), .B(A[232]), .Z(n1706) );
  XOR U1707 ( .A(n1707), .B(n1708), .Z(SUM[231]) );
  XNOR U1708 ( .A(B[231]), .B(A[231]), .Z(n1708) );
  XOR U1709 ( .A(n1709), .B(n1710), .Z(SUM[230]) );
  XNOR U1710 ( .A(B[230]), .B(A[230]), .Z(n1710) );
  XOR U1711 ( .A(n1711), .B(n1712), .Z(SUM[22]) );
  XNOR U1712 ( .A(B[22]), .B(A[22]), .Z(n1712) );
  XOR U1713 ( .A(n1713), .B(n1714), .Z(SUM[229]) );
  XNOR U1714 ( .A(B[229]), .B(A[229]), .Z(n1714) );
  XOR U1715 ( .A(n1715), .B(n1716), .Z(SUM[228]) );
  XNOR U1716 ( .A(B[228]), .B(A[228]), .Z(n1716) );
  XOR U1717 ( .A(n1717), .B(n1718), .Z(SUM[227]) );
  XNOR U1718 ( .A(B[227]), .B(A[227]), .Z(n1718) );
  XOR U1719 ( .A(n1719), .B(n1720), .Z(SUM[226]) );
  XNOR U1720 ( .A(B[226]), .B(A[226]), .Z(n1720) );
  XOR U1721 ( .A(n1721), .B(n1722), .Z(SUM[225]) );
  XNOR U1722 ( .A(B[225]), .B(A[225]), .Z(n1722) );
  XOR U1723 ( .A(n1723), .B(n1724), .Z(SUM[224]) );
  XNOR U1724 ( .A(B[224]), .B(A[224]), .Z(n1724) );
  XOR U1725 ( .A(n1725), .B(n1726), .Z(SUM[223]) );
  XNOR U1726 ( .A(B[223]), .B(A[223]), .Z(n1726) );
  XOR U1727 ( .A(n1727), .B(n1728), .Z(SUM[222]) );
  XNOR U1728 ( .A(B[222]), .B(A[222]), .Z(n1728) );
  XOR U1729 ( .A(n1729), .B(n1730), .Z(SUM[221]) );
  XNOR U1730 ( .A(B[221]), .B(A[221]), .Z(n1730) );
  XOR U1731 ( .A(n1731), .B(n1732), .Z(SUM[220]) );
  XNOR U1732 ( .A(B[220]), .B(A[220]), .Z(n1732) );
  XOR U1733 ( .A(n1733), .B(n1734), .Z(SUM[21]) );
  XNOR U1734 ( .A(B[21]), .B(A[21]), .Z(n1734) );
  XOR U1735 ( .A(n1735), .B(n1736), .Z(SUM[219]) );
  XNOR U1736 ( .A(B[219]), .B(A[219]), .Z(n1736) );
  XOR U1737 ( .A(n1737), .B(n1738), .Z(SUM[218]) );
  XNOR U1738 ( .A(B[218]), .B(A[218]), .Z(n1738) );
  XOR U1739 ( .A(n1739), .B(n1740), .Z(SUM[217]) );
  XNOR U1740 ( .A(B[217]), .B(A[217]), .Z(n1740) );
  XOR U1741 ( .A(n1741), .B(n1742), .Z(SUM[216]) );
  XNOR U1742 ( .A(B[216]), .B(A[216]), .Z(n1742) );
  XOR U1743 ( .A(n1743), .B(n1744), .Z(SUM[215]) );
  XNOR U1744 ( .A(B[215]), .B(A[215]), .Z(n1744) );
  XOR U1745 ( .A(n1745), .B(n1746), .Z(SUM[214]) );
  XNOR U1746 ( .A(B[214]), .B(A[214]), .Z(n1746) );
  XOR U1747 ( .A(n1747), .B(n1748), .Z(SUM[213]) );
  XNOR U1748 ( .A(B[213]), .B(A[213]), .Z(n1748) );
  XOR U1749 ( .A(n1749), .B(n1750), .Z(SUM[212]) );
  XNOR U1750 ( .A(B[212]), .B(A[212]), .Z(n1750) );
  XOR U1751 ( .A(n1751), .B(n1752), .Z(SUM[211]) );
  XNOR U1752 ( .A(B[211]), .B(A[211]), .Z(n1752) );
  XOR U1753 ( .A(n1753), .B(n1754), .Z(SUM[210]) );
  XNOR U1754 ( .A(B[210]), .B(A[210]), .Z(n1754) );
  XOR U1755 ( .A(n1755), .B(n1756), .Z(SUM[20]) );
  XNOR U1756 ( .A(B[20]), .B(A[20]), .Z(n1756) );
  XOR U1757 ( .A(n1757), .B(n1758), .Z(SUM[209]) );
  XNOR U1758 ( .A(B[209]), .B(A[209]), .Z(n1758) );
  XOR U1759 ( .A(n1759), .B(n1760), .Z(SUM[208]) );
  XNOR U1760 ( .A(B[208]), .B(A[208]), .Z(n1760) );
  XOR U1761 ( .A(n1761), .B(n1762), .Z(SUM[207]) );
  XNOR U1762 ( .A(B[207]), .B(A[207]), .Z(n1762) );
  XOR U1763 ( .A(n1763), .B(n1764), .Z(SUM[206]) );
  XNOR U1764 ( .A(B[206]), .B(A[206]), .Z(n1764) );
  XOR U1765 ( .A(n1765), .B(n1766), .Z(SUM[205]) );
  XNOR U1766 ( .A(B[205]), .B(A[205]), .Z(n1766) );
  XOR U1767 ( .A(n1767), .B(n1768), .Z(SUM[204]) );
  XNOR U1768 ( .A(B[204]), .B(A[204]), .Z(n1768) );
  XOR U1769 ( .A(n1769), .B(n1770), .Z(SUM[203]) );
  XNOR U1770 ( .A(B[203]), .B(A[203]), .Z(n1770) );
  XOR U1771 ( .A(n1771), .B(n1772), .Z(SUM[202]) );
  XNOR U1772 ( .A(B[202]), .B(A[202]), .Z(n1772) );
  XOR U1773 ( .A(n1773), .B(n1774), .Z(SUM[201]) );
  XNOR U1774 ( .A(B[201]), .B(A[201]), .Z(n1774) );
  XOR U1775 ( .A(n1775), .B(n1776), .Z(SUM[200]) );
  XNOR U1776 ( .A(B[200]), .B(A[200]), .Z(n1776) );
  XOR U1777 ( .A(B[1]), .B(A[1]), .Z(SUM[1]) );
  XOR U1778 ( .A(n1777), .B(n1778), .Z(SUM[19]) );
  XNOR U1779 ( .A(B[19]), .B(A[19]), .Z(n1778) );
  XOR U1780 ( .A(n1779), .B(n1780), .Z(SUM[199]) );
  XNOR U1781 ( .A(B[199]), .B(A[199]), .Z(n1780) );
  XOR U1782 ( .A(n1781), .B(n1782), .Z(SUM[198]) );
  XNOR U1783 ( .A(B[198]), .B(A[198]), .Z(n1782) );
  XOR U1784 ( .A(n1783), .B(n1784), .Z(SUM[197]) );
  XNOR U1785 ( .A(B[197]), .B(A[197]), .Z(n1784) );
  XOR U1786 ( .A(n1785), .B(n1786), .Z(SUM[196]) );
  XNOR U1787 ( .A(B[196]), .B(A[196]), .Z(n1786) );
  XOR U1788 ( .A(n1787), .B(n1788), .Z(SUM[195]) );
  XNOR U1789 ( .A(B[195]), .B(A[195]), .Z(n1788) );
  XOR U1790 ( .A(n1789), .B(n1790), .Z(SUM[194]) );
  XNOR U1791 ( .A(B[194]), .B(A[194]), .Z(n1790) );
  XOR U1792 ( .A(n1791), .B(n1792), .Z(SUM[193]) );
  XNOR U1793 ( .A(B[193]), .B(A[193]), .Z(n1792) );
  XOR U1794 ( .A(n1793), .B(n1794), .Z(SUM[192]) );
  XNOR U1795 ( .A(B[192]), .B(A[192]), .Z(n1794) );
  XOR U1796 ( .A(n1795), .B(n1796), .Z(SUM[191]) );
  XNOR U1797 ( .A(B[191]), .B(A[191]), .Z(n1796) );
  XOR U1798 ( .A(n1797), .B(n1798), .Z(SUM[190]) );
  XNOR U1799 ( .A(B[190]), .B(A[190]), .Z(n1798) );
  XOR U1800 ( .A(n1799), .B(n1800), .Z(SUM[18]) );
  XNOR U1801 ( .A(B[18]), .B(A[18]), .Z(n1800) );
  XOR U1802 ( .A(n1801), .B(n1802), .Z(SUM[189]) );
  XNOR U1803 ( .A(B[189]), .B(A[189]), .Z(n1802) );
  XOR U1804 ( .A(n1803), .B(n1804), .Z(SUM[188]) );
  XNOR U1805 ( .A(B[188]), .B(A[188]), .Z(n1804) );
  XOR U1806 ( .A(n1805), .B(n1806), .Z(SUM[187]) );
  XNOR U1807 ( .A(B[187]), .B(A[187]), .Z(n1806) );
  XOR U1808 ( .A(n1807), .B(n1808), .Z(SUM[186]) );
  XNOR U1809 ( .A(B[186]), .B(A[186]), .Z(n1808) );
  XOR U1810 ( .A(n1809), .B(n1810), .Z(SUM[185]) );
  XNOR U1811 ( .A(B[185]), .B(A[185]), .Z(n1810) );
  XOR U1812 ( .A(n1811), .B(n1812), .Z(SUM[184]) );
  XNOR U1813 ( .A(B[184]), .B(A[184]), .Z(n1812) );
  XOR U1814 ( .A(n1813), .B(n1814), .Z(SUM[183]) );
  XNOR U1815 ( .A(B[183]), .B(A[183]), .Z(n1814) );
  XOR U1816 ( .A(n1815), .B(n1816), .Z(SUM[182]) );
  XNOR U1817 ( .A(B[182]), .B(A[182]), .Z(n1816) );
  XOR U1818 ( .A(n1817), .B(n1818), .Z(SUM[181]) );
  XNOR U1819 ( .A(B[181]), .B(A[181]), .Z(n1818) );
  XOR U1820 ( .A(n1819), .B(n1820), .Z(SUM[180]) );
  XNOR U1821 ( .A(B[180]), .B(A[180]), .Z(n1820) );
  XOR U1822 ( .A(n1821), .B(n1822), .Z(SUM[17]) );
  XNOR U1823 ( .A(B[17]), .B(A[17]), .Z(n1822) );
  XOR U1824 ( .A(n1823), .B(n1824), .Z(SUM[179]) );
  XNOR U1825 ( .A(B[179]), .B(A[179]), .Z(n1824) );
  XOR U1826 ( .A(n1825), .B(n1826), .Z(SUM[178]) );
  XNOR U1827 ( .A(B[178]), .B(A[178]), .Z(n1826) );
  XOR U1828 ( .A(n1827), .B(n1828), .Z(SUM[177]) );
  XNOR U1829 ( .A(B[177]), .B(A[177]), .Z(n1828) );
  XOR U1830 ( .A(n1829), .B(n1830), .Z(SUM[176]) );
  XNOR U1831 ( .A(B[176]), .B(A[176]), .Z(n1830) );
  XOR U1832 ( .A(n1831), .B(n1832), .Z(SUM[175]) );
  XNOR U1833 ( .A(B[175]), .B(A[175]), .Z(n1832) );
  XOR U1834 ( .A(n1833), .B(n1834), .Z(SUM[174]) );
  XNOR U1835 ( .A(B[174]), .B(A[174]), .Z(n1834) );
  XOR U1836 ( .A(n1835), .B(n1836), .Z(SUM[173]) );
  XNOR U1837 ( .A(B[173]), .B(A[173]), .Z(n1836) );
  XOR U1838 ( .A(n1837), .B(n1838), .Z(SUM[172]) );
  XNOR U1839 ( .A(B[172]), .B(A[172]), .Z(n1838) );
  XOR U1840 ( .A(n1839), .B(n1840), .Z(SUM[171]) );
  XNOR U1841 ( .A(B[171]), .B(A[171]), .Z(n1840) );
  XOR U1842 ( .A(n1841), .B(n1842), .Z(SUM[170]) );
  XNOR U1843 ( .A(B[170]), .B(A[170]), .Z(n1842) );
  XOR U1844 ( .A(n1843), .B(n1844), .Z(SUM[16]) );
  XNOR U1845 ( .A(B[16]), .B(A[16]), .Z(n1844) );
  XOR U1846 ( .A(n1845), .B(n1846), .Z(SUM[169]) );
  XNOR U1847 ( .A(B[169]), .B(A[169]), .Z(n1846) );
  XOR U1848 ( .A(n1847), .B(n1848), .Z(SUM[168]) );
  XNOR U1849 ( .A(B[168]), .B(A[168]), .Z(n1848) );
  XOR U1850 ( .A(n1849), .B(n1850), .Z(SUM[167]) );
  XNOR U1851 ( .A(B[167]), .B(A[167]), .Z(n1850) );
  XOR U1852 ( .A(n1851), .B(n1852), .Z(SUM[166]) );
  XNOR U1853 ( .A(B[166]), .B(A[166]), .Z(n1852) );
  XOR U1854 ( .A(n1853), .B(n1854), .Z(SUM[165]) );
  XNOR U1855 ( .A(B[165]), .B(A[165]), .Z(n1854) );
  XOR U1856 ( .A(n1855), .B(n1856), .Z(SUM[164]) );
  XNOR U1857 ( .A(B[164]), .B(A[164]), .Z(n1856) );
  XOR U1858 ( .A(n1857), .B(n1858), .Z(SUM[163]) );
  XNOR U1859 ( .A(B[163]), .B(A[163]), .Z(n1858) );
  XOR U1860 ( .A(n1859), .B(n1860), .Z(SUM[162]) );
  XNOR U1861 ( .A(B[162]), .B(A[162]), .Z(n1860) );
  XOR U1862 ( .A(n1861), .B(n1862), .Z(SUM[161]) );
  XNOR U1863 ( .A(B[161]), .B(A[161]), .Z(n1862) );
  XOR U1864 ( .A(n1863), .B(n1864), .Z(SUM[160]) );
  XNOR U1865 ( .A(B[160]), .B(A[160]), .Z(n1864) );
  XOR U1866 ( .A(n1865), .B(n1866), .Z(SUM[15]) );
  XNOR U1867 ( .A(B[15]), .B(A[15]), .Z(n1866) );
  XOR U1868 ( .A(n1867), .B(n1868), .Z(SUM[159]) );
  XNOR U1869 ( .A(B[159]), .B(A[159]), .Z(n1868) );
  XOR U1870 ( .A(n1869), .B(n1870), .Z(SUM[158]) );
  XNOR U1871 ( .A(B[158]), .B(A[158]), .Z(n1870) );
  XOR U1872 ( .A(n1871), .B(n1872), .Z(SUM[157]) );
  XNOR U1873 ( .A(B[157]), .B(A[157]), .Z(n1872) );
  XOR U1874 ( .A(n1873), .B(n1874), .Z(SUM[156]) );
  XNOR U1875 ( .A(B[156]), .B(A[156]), .Z(n1874) );
  XOR U1876 ( .A(n1875), .B(n1876), .Z(SUM[155]) );
  XNOR U1877 ( .A(B[155]), .B(A[155]), .Z(n1876) );
  XOR U1878 ( .A(n1877), .B(n1878), .Z(SUM[154]) );
  XNOR U1879 ( .A(B[154]), .B(A[154]), .Z(n1878) );
  XOR U1880 ( .A(n1879), .B(n1880), .Z(SUM[153]) );
  XNOR U1881 ( .A(B[153]), .B(A[153]), .Z(n1880) );
  XOR U1882 ( .A(n1881), .B(n1882), .Z(SUM[152]) );
  XNOR U1883 ( .A(B[152]), .B(A[152]), .Z(n1882) );
  XOR U1884 ( .A(n1883), .B(n1884), .Z(SUM[151]) );
  XNOR U1885 ( .A(B[151]), .B(A[151]), .Z(n1884) );
  XOR U1886 ( .A(n1885), .B(n1886), .Z(SUM[150]) );
  XNOR U1887 ( .A(B[150]), .B(A[150]), .Z(n1886) );
  XOR U1888 ( .A(n1887), .B(n1888), .Z(SUM[14]) );
  XNOR U1889 ( .A(B[14]), .B(A[14]), .Z(n1888) );
  XOR U1890 ( .A(n1889), .B(n1890), .Z(SUM[149]) );
  XNOR U1891 ( .A(B[149]), .B(A[149]), .Z(n1890) );
  XOR U1892 ( .A(n1891), .B(n1892), .Z(SUM[148]) );
  XNOR U1893 ( .A(B[148]), .B(A[148]), .Z(n1892) );
  XOR U1894 ( .A(n1893), .B(n1894), .Z(SUM[147]) );
  XNOR U1895 ( .A(B[147]), .B(A[147]), .Z(n1894) );
  XOR U1896 ( .A(n1895), .B(n1896), .Z(SUM[146]) );
  XNOR U1897 ( .A(B[146]), .B(A[146]), .Z(n1896) );
  XOR U1898 ( .A(n1897), .B(n1898), .Z(SUM[145]) );
  XNOR U1899 ( .A(B[145]), .B(A[145]), .Z(n1898) );
  XOR U1900 ( .A(n1899), .B(n1900), .Z(SUM[144]) );
  XNOR U1901 ( .A(B[144]), .B(A[144]), .Z(n1900) );
  XOR U1902 ( .A(n1901), .B(n1902), .Z(SUM[143]) );
  XNOR U1903 ( .A(B[143]), .B(A[143]), .Z(n1902) );
  XOR U1904 ( .A(n1903), .B(n1904), .Z(SUM[142]) );
  XNOR U1905 ( .A(B[142]), .B(A[142]), .Z(n1904) );
  XOR U1906 ( .A(n1905), .B(n1906), .Z(SUM[141]) );
  XNOR U1907 ( .A(B[141]), .B(A[141]), .Z(n1906) );
  XOR U1908 ( .A(n1907), .B(n1908), .Z(SUM[140]) );
  XNOR U1909 ( .A(B[140]), .B(A[140]), .Z(n1908) );
  XOR U1910 ( .A(n1909), .B(n1910), .Z(SUM[13]) );
  XNOR U1911 ( .A(B[13]), .B(A[13]), .Z(n1910) );
  XOR U1912 ( .A(n1911), .B(n1912), .Z(SUM[139]) );
  XNOR U1913 ( .A(B[139]), .B(A[139]), .Z(n1912) );
  XOR U1914 ( .A(n1913), .B(n1914), .Z(SUM[138]) );
  XNOR U1915 ( .A(B[138]), .B(A[138]), .Z(n1914) );
  XOR U1916 ( .A(n1915), .B(n1916), .Z(SUM[137]) );
  XNOR U1917 ( .A(B[137]), .B(A[137]), .Z(n1916) );
  XOR U1918 ( .A(n1917), .B(n1918), .Z(SUM[136]) );
  XNOR U1919 ( .A(B[136]), .B(A[136]), .Z(n1918) );
  XOR U1920 ( .A(n1919), .B(n1920), .Z(SUM[135]) );
  XNOR U1921 ( .A(B[135]), .B(A[135]), .Z(n1920) );
  XOR U1922 ( .A(n1921), .B(n1922), .Z(SUM[134]) );
  XNOR U1923 ( .A(B[134]), .B(A[134]), .Z(n1922) );
  XOR U1924 ( .A(n1923), .B(n1924), .Z(SUM[133]) );
  XNOR U1925 ( .A(B[133]), .B(A[133]), .Z(n1924) );
  XOR U1926 ( .A(n1925), .B(n1926), .Z(SUM[132]) );
  XNOR U1927 ( .A(B[132]), .B(A[132]), .Z(n1926) );
  XOR U1928 ( .A(n1927), .B(n1928), .Z(SUM[131]) );
  XNOR U1929 ( .A(B[131]), .B(A[131]), .Z(n1928) );
  XOR U1930 ( .A(n1929), .B(n1930), .Z(SUM[130]) );
  XNOR U1931 ( .A(B[130]), .B(A[130]), .Z(n1930) );
  XOR U1932 ( .A(n1931), .B(n1932), .Z(SUM[12]) );
  XNOR U1933 ( .A(B[12]), .B(A[12]), .Z(n1932) );
  XOR U1934 ( .A(n1933), .B(n1934), .Z(SUM[129]) );
  XNOR U1935 ( .A(B[129]), .B(A[129]), .Z(n1934) );
  XOR U1936 ( .A(n1935), .B(n1936), .Z(SUM[128]) );
  XNOR U1937 ( .A(B[128]), .B(A[128]), .Z(n1936) );
  XOR U1938 ( .A(n1937), .B(n1938), .Z(SUM[127]) );
  XNOR U1939 ( .A(B[127]), .B(A[127]), .Z(n1938) );
  XOR U1940 ( .A(n1939), .B(n1940), .Z(SUM[126]) );
  XNOR U1941 ( .A(B[126]), .B(A[126]), .Z(n1940) );
  XOR U1942 ( .A(n1941), .B(n1942), .Z(SUM[125]) );
  XNOR U1943 ( .A(B[125]), .B(A[125]), .Z(n1942) );
  XOR U1944 ( .A(n1943), .B(n1944), .Z(SUM[124]) );
  XNOR U1945 ( .A(B[124]), .B(A[124]), .Z(n1944) );
  XOR U1946 ( .A(n1945), .B(n1946), .Z(SUM[123]) );
  XNOR U1947 ( .A(B[123]), .B(A[123]), .Z(n1946) );
  XOR U1948 ( .A(n1947), .B(n1948), .Z(SUM[122]) );
  XNOR U1949 ( .A(B[122]), .B(A[122]), .Z(n1948) );
  XOR U1950 ( .A(n1949), .B(n1950), .Z(SUM[121]) );
  XNOR U1951 ( .A(B[121]), .B(A[121]), .Z(n1950) );
  XOR U1952 ( .A(n1951), .B(n1952), .Z(SUM[120]) );
  XNOR U1953 ( .A(B[120]), .B(A[120]), .Z(n1952) );
  XOR U1954 ( .A(n1953), .B(n1954), .Z(SUM[11]) );
  XNOR U1955 ( .A(B[11]), .B(A[11]), .Z(n1954) );
  XOR U1956 ( .A(n1955), .B(n1956), .Z(SUM[119]) );
  XNOR U1957 ( .A(B[119]), .B(A[119]), .Z(n1956) );
  XOR U1958 ( .A(n1957), .B(n1958), .Z(SUM[118]) );
  XNOR U1959 ( .A(B[118]), .B(A[118]), .Z(n1958) );
  XOR U1960 ( .A(n1959), .B(n1960), .Z(SUM[117]) );
  XNOR U1961 ( .A(B[117]), .B(A[117]), .Z(n1960) );
  XOR U1962 ( .A(n1961), .B(n1962), .Z(SUM[116]) );
  XNOR U1963 ( .A(B[116]), .B(A[116]), .Z(n1962) );
  XOR U1964 ( .A(n1963), .B(n1964), .Z(SUM[115]) );
  XNOR U1965 ( .A(B[115]), .B(A[115]), .Z(n1964) );
  XOR U1966 ( .A(n1965), .B(n1966), .Z(SUM[114]) );
  XNOR U1967 ( .A(B[114]), .B(A[114]), .Z(n1966) );
  XOR U1968 ( .A(n1967), .B(n1968), .Z(SUM[113]) );
  XNOR U1969 ( .A(B[113]), .B(A[113]), .Z(n1968) );
  XOR U1970 ( .A(n1969), .B(n1970), .Z(SUM[112]) );
  XNOR U1971 ( .A(B[112]), .B(A[112]), .Z(n1970) );
  XOR U1972 ( .A(n1971), .B(n1972), .Z(SUM[111]) );
  XNOR U1973 ( .A(B[111]), .B(A[111]), .Z(n1972) );
  XOR U1974 ( .A(n1973), .B(n1974), .Z(SUM[110]) );
  XNOR U1975 ( .A(B[110]), .B(A[110]), .Z(n1974) );
  XOR U1976 ( .A(n1975), .B(n1976), .Z(SUM[10]) );
  XNOR U1977 ( .A(B[10]), .B(A[10]), .Z(n1976) );
  XOR U1978 ( .A(n1977), .B(n1978), .Z(SUM[109]) );
  XNOR U1979 ( .A(B[109]), .B(A[109]), .Z(n1978) );
  XOR U1980 ( .A(n1979), .B(n1980), .Z(SUM[108]) );
  XNOR U1981 ( .A(B[108]), .B(A[108]), .Z(n1980) );
  XOR U1982 ( .A(n1981), .B(n1982), .Z(SUM[107]) );
  XNOR U1983 ( .A(B[107]), .B(A[107]), .Z(n1982) );
  XOR U1984 ( .A(n1983), .B(n1984), .Z(SUM[106]) );
  XNOR U1985 ( .A(B[106]), .B(A[106]), .Z(n1984) );
  XOR U1986 ( .A(n1985), .B(n1986), .Z(SUM[105]) );
  XNOR U1987 ( .A(B[105]), .B(A[105]), .Z(n1986) );
  XOR U1988 ( .A(n1987), .B(n1988), .Z(SUM[104]) );
  XNOR U1989 ( .A(B[104]), .B(A[104]), .Z(n1988) );
  XOR U1990 ( .A(n1989), .B(n1990), .Z(SUM[103]) );
  XNOR U1991 ( .A(B[103]), .B(A[103]), .Z(n1990) );
  XOR U1992 ( .A(n1991), .B(n1992), .Z(SUM[102]) );
  XNOR U1993 ( .A(B[102]), .B(A[102]), .Z(n1992) );
  XOR U1994 ( .A(A[1025]), .B(n1993), .Z(SUM[1025]) );
  AND U1995 ( .A(A[1024]), .B(n1994), .Z(n1993) );
  XOR U1996 ( .A(A[1024]), .B(n1994), .Z(SUM[1024]) );
  NAND U1997 ( .A(n1995), .B(n1996), .Z(n1994) );
  NAND U1998 ( .A(B[1023]), .B(n1997), .Z(n1996) );
  NANDN U1999 ( .A(A[1023]), .B(n1998), .Z(n1997) );
  NANDN U2000 ( .A(n1998), .B(A[1023]), .Z(n1995) );
  XOR U2001 ( .A(n1998), .B(n1999), .Z(SUM[1023]) );
  XNOR U2002 ( .A(B[1023]), .B(A[1023]), .Z(n1999) );
  AND U2003 ( .A(n2000), .B(n2001), .Z(n1998) );
  NAND U2004 ( .A(B[1022]), .B(n2002), .Z(n2001) );
  NANDN U2005 ( .A(A[1022]), .B(n2003), .Z(n2002) );
  NANDN U2006 ( .A(n2003), .B(A[1022]), .Z(n2000) );
  XOR U2007 ( .A(n2003), .B(n2004), .Z(SUM[1022]) );
  XNOR U2008 ( .A(B[1022]), .B(A[1022]), .Z(n2004) );
  AND U2009 ( .A(n2005), .B(n2006), .Z(n2003) );
  NAND U2010 ( .A(B[1021]), .B(n2007), .Z(n2006) );
  NANDN U2011 ( .A(A[1021]), .B(n2008), .Z(n2007) );
  NANDN U2012 ( .A(n2008), .B(A[1021]), .Z(n2005) );
  XOR U2013 ( .A(n2008), .B(n2009), .Z(SUM[1021]) );
  XNOR U2014 ( .A(B[1021]), .B(A[1021]), .Z(n2009) );
  AND U2015 ( .A(n2010), .B(n2011), .Z(n2008) );
  NAND U2016 ( .A(B[1020]), .B(n2012), .Z(n2011) );
  NANDN U2017 ( .A(A[1020]), .B(n2013), .Z(n2012) );
  NANDN U2018 ( .A(n2013), .B(A[1020]), .Z(n2010) );
  XOR U2019 ( .A(n2013), .B(n2014), .Z(SUM[1020]) );
  XNOR U2020 ( .A(B[1020]), .B(A[1020]), .Z(n2014) );
  AND U2021 ( .A(n2015), .B(n2016), .Z(n2013) );
  NAND U2022 ( .A(B[1019]), .B(n2017), .Z(n2016) );
  NANDN U2023 ( .A(A[1019]), .B(n2018), .Z(n2017) );
  NANDN U2024 ( .A(n2018), .B(A[1019]), .Z(n2015) );
  XOR U2025 ( .A(n2019), .B(n2020), .Z(SUM[101]) );
  XNOR U2026 ( .A(B[101]), .B(A[101]), .Z(n2020) );
  XOR U2027 ( .A(n2018), .B(n2021), .Z(SUM[1019]) );
  XNOR U2028 ( .A(B[1019]), .B(A[1019]), .Z(n2021) );
  AND U2029 ( .A(n2022), .B(n2023), .Z(n2018) );
  NAND U2030 ( .A(B[1018]), .B(n2024), .Z(n2023) );
  NANDN U2031 ( .A(A[1018]), .B(n2025), .Z(n2024) );
  NANDN U2032 ( .A(n2025), .B(A[1018]), .Z(n2022) );
  XOR U2033 ( .A(n2025), .B(n2026), .Z(SUM[1018]) );
  XNOR U2034 ( .A(B[1018]), .B(A[1018]), .Z(n2026) );
  AND U2035 ( .A(n2027), .B(n2028), .Z(n2025) );
  NAND U2036 ( .A(B[1017]), .B(n2029), .Z(n2028) );
  NANDN U2037 ( .A(A[1017]), .B(n2030), .Z(n2029) );
  NANDN U2038 ( .A(n2030), .B(A[1017]), .Z(n2027) );
  XOR U2039 ( .A(n2030), .B(n2031), .Z(SUM[1017]) );
  XNOR U2040 ( .A(B[1017]), .B(A[1017]), .Z(n2031) );
  AND U2041 ( .A(n2032), .B(n2033), .Z(n2030) );
  NAND U2042 ( .A(B[1016]), .B(n2034), .Z(n2033) );
  NANDN U2043 ( .A(A[1016]), .B(n2035), .Z(n2034) );
  NANDN U2044 ( .A(n2035), .B(A[1016]), .Z(n2032) );
  XOR U2045 ( .A(n2035), .B(n2036), .Z(SUM[1016]) );
  XNOR U2046 ( .A(B[1016]), .B(A[1016]), .Z(n2036) );
  AND U2047 ( .A(n2037), .B(n2038), .Z(n2035) );
  NAND U2048 ( .A(B[1015]), .B(n2039), .Z(n2038) );
  NANDN U2049 ( .A(A[1015]), .B(n2040), .Z(n2039) );
  NANDN U2050 ( .A(n2040), .B(A[1015]), .Z(n2037) );
  XOR U2051 ( .A(n2040), .B(n2041), .Z(SUM[1015]) );
  XNOR U2052 ( .A(B[1015]), .B(A[1015]), .Z(n2041) );
  AND U2053 ( .A(n2042), .B(n2043), .Z(n2040) );
  NAND U2054 ( .A(B[1014]), .B(n2044), .Z(n2043) );
  NANDN U2055 ( .A(A[1014]), .B(n2045), .Z(n2044) );
  NANDN U2056 ( .A(n2045), .B(A[1014]), .Z(n2042) );
  XOR U2057 ( .A(n2045), .B(n2046), .Z(SUM[1014]) );
  XNOR U2058 ( .A(B[1014]), .B(A[1014]), .Z(n2046) );
  AND U2059 ( .A(n2047), .B(n2048), .Z(n2045) );
  NAND U2060 ( .A(B[1013]), .B(n2049), .Z(n2048) );
  NANDN U2061 ( .A(A[1013]), .B(n2050), .Z(n2049) );
  NANDN U2062 ( .A(n2050), .B(A[1013]), .Z(n2047) );
  XOR U2063 ( .A(n2050), .B(n2051), .Z(SUM[1013]) );
  XNOR U2064 ( .A(B[1013]), .B(A[1013]), .Z(n2051) );
  AND U2065 ( .A(n2052), .B(n2053), .Z(n2050) );
  NAND U2066 ( .A(B[1012]), .B(n2054), .Z(n2053) );
  NANDN U2067 ( .A(A[1012]), .B(n2055), .Z(n2054) );
  NANDN U2068 ( .A(n2055), .B(A[1012]), .Z(n2052) );
  XOR U2069 ( .A(n2055), .B(n2056), .Z(SUM[1012]) );
  XNOR U2070 ( .A(B[1012]), .B(A[1012]), .Z(n2056) );
  AND U2071 ( .A(n2057), .B(n2058), .Z(n2055) );
  NAND U2072 ( .A(B[1011]), .B(n2059), .Z(n2058) );
  NANDN U2073 ( .A(A[1011]), .B(n2060), .Z(n2059) );
  NANDN U2074 ( .A(n2060), .B(A[1011]), .Z(n2057) );
  XOR U2075 ( .A(n2060), .B(n2061), .Z(SUM[1011]) );
  XNOR U2076 ( .A(B[1011]), .B(A[1011]), .Z(n2061) );
  AND U2077 ( .A(n2062), .B(n2063), .Z(n2060) );
  NAND U2078 ( .A(B[1010]), .B(n2064), .Z(n2063) );
  NANDN U2079 ( .A(A[1010]), .B(n2065), .Z(n2064) );
  NANDN U2080 ( .A(n2065), .B(A[1010]), .Z(n2062) );
  XOR U2081 ( .A(n2065), .B(n2066), .Z(SUM[1010]) );
  XNOR U2082 ( .A(B[1010]), .B(A[1010]), .Z(n2066) );
  AND U2083 ( .A(n2067), .B(n2068), .Z(n2065) );
  NAND U2084 ( .A(B[1009]), .B(n2069), .Z(n2068) );
  NANDN U2085 ( .A(A[1009]), .B(n2070), .Z(n2069) );
  NANDN U2086 ( .A(n2070), .B(A[1009]), .Z(n2067) );
  XOR U2087 ( .A(n2071), .B(n2072), .Z(SUM[100]) );
  XNOR U2088 ( .A(B[100]), .B(A[100]), .Z(n2072) );
  XOR U2089 ( .A(n2070), .B(n2073), .Z(SUM[1009]) );
  XNOR U2090 ( .A(B[1009]), .B(A[1009]), .Z(n2073) );
  AND U2091 ( .A(n2074), .B(n2075), .Z(n2070) );
  NAND U2092 ( .A(B[1008]), .B(n2076), .Z(n2075) );
  NANDN U2093 ( .A(A[1008]), .B(n2077), .Z(n2076) );
  NANDN U2094 ( .A(n2077), .B(A[1008]), .Z(n2074) );
  XOR U2095 ( .A(n2077), .B(n2078), .Z(SUM[1008]) );
  XNOR U2096 ( .A(B[1008]), .B(A[1008]), .Z(n2078) );
  AND U2097 ( .A(n2079), .B(n2080), .Z(n2077) );
  NAND U2098 ( .A(B[1007]), .B(n2081), .Z(n2080) );
  NANDN U2099 ( .A(A[1007]), .B(n2082), .Z(n2081) );
  NANDN U2100 ( .A(n2082), .B(A[1007]), .Z(n2079) );
  XOR U2101 ( .A(n2082), .B(n2083), .Z(SUM[1007]) );
  XNOR U2102 ( .A(B[1007]), .B(A[1007]), .Z(n2083) );
  AND U2103 ( .A(n2084), .B(n2085), .Z(n2082) );
  NAND U2104 ( .A(B[1006]), .B(n2086), .Z(n2085) );
  NANDN U2105 ( .A(A[1006]), .B(n2087), .Z(n2086) );
  NANDN U2106 ( .A(n2087), .B(A[1006]), .Z(n2084) );
  XOR U2107 ( .A(n2087), .B(n2088), .Z(SUM[1006]) );
  XNOR U2108 ( .A(B[1006]), .B(A[1006]), .Z(n2088) );
  AND U2109 ( .A(n2089), .B(n2090), .Z(n2087) );
  NAND U2110 ( .A(B[1005]), .B(n2091), .Z(n2090) );
  NANDN U2111 ( .A(A[1005]), .B(n2092), .Z(n2091) );
  NANDN U2112 ( .A(n2092), .B(A[1005]), .Z(n2089) );
  XOR U2113 ( .A(n2092), .B(n2093), .Z(SUM[1005]) );
  XNOR U2114 ( .A(B[1005]), .B(A[1005]), .Z(n2093) );
  AND U2115 ( .A(n2094), .B(n2095), .Z(n2092) );
  NAND U2116 ( .A(B[1004]), .B(n2096), .Z(n2095) );
  NANDN U2117 ( .A(A[1004]), .B(n2097), .Z(n2096) );
  NANDN U2118 ( .A(n2097), .B(A[1004]), .Z(n2094) );
  XOR U2119 ( .A(n2097), .B(n2098), .Z(SUM[1004]) );
  XNOR U2120 ( .A(B[1004]), .B(A[1004]), .Z(n2098) );
  AND U2121 ( .A(n2099), .B(n2100), .Z(n2097) );
  NAND U2122 ( .A(B[1003]), .B(n2101), .Z(n2100) );
  NANDN U2123 ( .A(A[1003]), .B(n2102), .Z(n2101) );
  NANDN U2124 ( .A(n2102), .B(A[1003]), .Z(n2099) );
  XOR U2125 ( .A(n2102), .B(n2103), .Z(SUM[1003]) );
  XNOR U2126 ( .A(B[1003]), .B(A[1003]), .Z(n2103) );
  AND U2127 ( .A(n2104), .B(n2105), .Z(n2102) );
  NAND U2128 ( .A(B[1002]), .B(n2106), .Z(n2105) );
  NANDN U2129 ( .A(A[1002]), .B(n2107), .Z(n2106) );
  NANDN U2130 ( .A(n2107), .B(A[1002]), .Z(n2104) );
  XOR U2131 ( .A(n2107), .B(n2108), .Z(SUM[1002]) );
  XNOR U2132 ( .A(B[1002]), .B(A[1002]), .Z(n2108) );
  AND U2133 ( .A(n2109), .B(n2110), .Z(n2107) );
  NAND U2134 ( .A(B[1001]), .B(n2111), .Z(n2110) );
  NANDN U2135 ( .A(A[1001]), .B(n2112), .Z(n2111) );
  NANDN U2136 ( .A(n2112), .B(A[1001]), .Z(n2109) );
  XOR U2137 ( .A(n2112), .B(n2113), .Z(SUM[1001]) );
  XNOR U2138 ( .A(B[1001]), .B(A[1001]), .Z(n2113) );
  AND U2139 ( .A(n2114), .B(n2115), .Z(n2112) );
  NAND U2140 ( .A(B[1000]), .B(n2116), .Z(n2115) );
  NANDN U2141 ( .A(A[1000]), .B(n2117), .Z(n2116) );
  NANDN U2142 ( .A(n2117), .B(A[1000]), .Z(n2114) );
  XOR U2143 ( .A(n2117), .B(n2118), .Z(SUM[1000]) );
  XNOR U2144 ( .A(B[1000]), .B(A[1000]), .Z(n2118) );
  AND U2145 ( .A(n2119), .B(n2120), .Z(n2117) );
  NAND U2146 ( .A(B[999]), .B(n2121), .Z(n2120) );
  OR U2147 ( .A(n5), .B(A[999]), .Z(n2121) );
  NAND U2148 ( .A(A[999]), .B(n5), .Z(n2119) );
  NAND U2149 ( .A(n2122), .B(n2123), .Z(n5) );
  NAND U2150 ( .A(B[998]), .B(n2124), .Z(n2123) );
  NANDN U2151 ( .A(A[998]), .B(n7), .Z(n2124) );
  NANDN U2152 ( .A(n7), .B(A[998]), .Z(n2122) );
  AND U2153 ( .A(n2125), .B(n2126), .Z(n7) );
  NAND U2154 ( .A(B[997]), .B(n2127), .Z(n2126) );
  NANDN U2155 ( .A(A[997]), .B(n9), .Z(n2127) );
  NANDN U2156 ( .A(n9), .B(A[997]), .Z(n2125) );
  AND U2157 ( .A(n2128), .B(n2129), .Z(n9) );
  NAND U2158 ( .A(B[996]), .B(n2130), .Z(n2129) );
  NANDN U2159 ( .A(A[996]), .B(n11), .Z(n2130) );
  NANDN U2160 ( .A(n11), .B(A[996]), .Z(n2128) );
  AND U2161 ( .A(n2131), .B(n2132), .Z(n11) );
  NAND U2162 ( .A(B[995]), .B(n2133), .Z(n2132) );
  NANDN U2163 ( .A(A[995]), .B(n13), .Z(n2133) );
  NANDN U2164 ( .A(n13), .B(A[995]), .Z(n2131) );
  AND U2165 ( .A(n2134), .B(n2135), .Z(n13) );
  NAND U2166 ( .A(B[994]), .B(n2136), .Z(n2135) );
  NANDN U2167 ( .A(A[994]), .B(n15), .Z(n2136) );
  NANDN U2168 ( .A(n15), .B(A[994]), .Z(n2134) );
  AND U2169 ( .A(n2137), .B(n2138), .Z(n15) );
  NAND U2170 ( .A(B[993]), .B(n2139), .Z(n2138) );
  NANDN U2171 ( .A(A[993]), .B(n17), .Z(n2139) );
  NANDN U2172 ( .A(n17), .B(A[993]), .Z(n2137) );
  AND U2173 ( .A(n2140), .B(n2141), .Z(n17) );
  NAND U2174 ( .A(B[992]), .B(n2142), .Z(n2141) );
  NANDN U2175 ( .A(A[992]), .B(n19), .Z(n2142) );
  NANDN U2176 ( .A(n19), .B(A[992]), .Z(n2140) );
  AND U2177 ( .A(n2143), .B(n2144), .Z(n19) );
  NAND U2178 ( .A(B[991]), .B(n2145), .Z(n2144) );
  NANDN U2179 ( .A(A[991]), .B(n21), .Z(n2145) );
  NANDN U2180 ( .A(n21), .B(A[991]), .Z(n2143) );
  AND U2181 ( .A(n2146), .B(n2147), .Z(n21) );
  NAND U2182 ( .A(B[990]), .B(n2148), .Z(n2147) );
  NANDN U2183 ( .A(A[990]), .B(n23), .Z(n2148) );
  NANDN U2184 ( .A(n23), .B(A[990]), .Z(n2146) );
  AND U2185 ( .A(n2149), .B(n2150), .Z(n23) );
  NAND U2186 ( .A(B[989]), .B(n2151), .Z(n2150) );
  NANDN U2187 ( .A(A[989]), .B(n27), .Z(n2151) );
  NANDN U2188 ( .A(n27), .B(A[989]), .Z(n2149) );
  AND U2189 ( .A(n2152), .B(n2153), .Z(n27) );
  NAND U2190 ( .A(B[988]), .B(n2154), .Z(n2153) );
  NANDN U2191 ( .A(A[988]), .B(n29), .Z(n2154) );
  NANDN U2192 ( .A(n29), .B(A[988]), .Z(n2152) );
  AND U2193 ( .A(n2155), .B(n2156), .Z(n29) );
  NAND U2194 ( .A(B[987]), .B(n2157), .Z(n2156) );
  NANDN U2195 ( .A(A[987]), .B(n31), .Z(n2157) );
  NANDN U2196 ( .A(n31), .B(A[987]), .Z(n2155) );
  AND U2197 ( .A(n2158), .B(n2159), .Z(n31) );
  NAND U2198 ( .A(B[986]), .B(n2160), .Z(n2159) );
  NANDN U2199 ( .A(A[986]), .B(n33), .Z(n2160) );
  NANDN U2200 ( .A(n33), .B(A[986]), .Z(n2158) );
  AND U2201 ( .A(n2161), .B(n2162), .Z(n33) );
  NAND U2202 ( .A(B[985]), .B(n2163), .Z(n2162) );
  NANDN U2203 ( .A(A[985]), .B(n35), .Z(n2163) );
  NANDN U2204 ( .A(n35), .B(A[985]), .Z(n2161) );
  AND U2205 ( .A(n2164), .B(n2165), .Z(n35) );
  NAND U2206 ( .A(B[984]), .B(n2166), .Z(n2165) );
  NANDN U2207 ( .A(A[984]), .B(n37), .Z(n2166) );
  NANDN U2208 ( .A(n37), .B(A[984]), .Z(n2164) );
  AND U2209 ( .A(n2167), .B(n2168), .Z(n37) );
  NAND U2210 ( .A(B[983]), .B(n2169), .Z(n2168) );
  NANDN U2211 ( .A(A[983]), .B(n39), .Z(n2169) );
  NANDN U2212 ( .A(n39), .B(A[983]), .Z(n2167) );
  AND U2213 ( .A(n2170), .B(n2171), .Z(n39) );
  NAND U2214 ( .A(B[982]), .B(n2172), .Z(n2171) );
  NANDN U2215 ( .A(A[982]), .B(n41), .Z(n2172) );
  NANDN U2216 ( .A(n41), .B(A[982]), .Z(n2170) );
  AND U2217 ( .A(n2173), .B(n2174), .Z(n41) );
  NAND U2218 ( .A(B[981]), .B(n2175), .Z(n2174) );
  NANDN U2219 ( .A(A[981]), .B(n43), .Z(n2175) );
  NANDN U2220 ( .A(n43), .B(A[981]), .Z(n2173) );
  AND U2221 ( .A(n2176), .B(n2177), .Z(n43) );
  NAND U2222 ( .A(B[980]), .B(n2178), .Z(n2177) );
  NANDN U2223 ( .A(A[980]), .B(n45), .Z(n2178) );
  NANDN U2224 ( .A(n45), .B(A[980]), .Z(n2176) );
  AND U2225 ( .A(n2179), .B(n2180), .Z(n45) );
  NAND U2226 ( .A(B[979]), .B(n2181), .Z(n2180) );
  NANDN U2227 ( .A(A[979]), .B(n49), .Z(n2181) );
  NANDN U2228 ( .A(n49), .B(A[979]), .Z(n2179) );
  AND U2229 ( .A(n2182), .B(n2183), .Z(n49) );
  NAND U2230 ( .A(B[978]), .B(n2184), .Z(n2183) );
  NANDN U2231 ( .A(A[978]), .B(n51), .Z(n2184) );
  NANDN U2232 ( .A(n51), .B(A[978]), .Z(n2182) );
  AND U2233 ( .A(n2185), .B(n2186), .Z(n51) );
  NAND U2234 ( .A(B[977]), .B(n2187), .Z(n2186) );
  NANDN U2235 ( .A(A[977]), .B(n53), .Z(n2187) );
  NANDN U2236 ( .A(n53), .B(A[977]), .Z(n2185) );
  AND U2237 ( .A(n2188), .B(n2189), .Z(n53) );
  NAND U2238 ( .A(B[976]), .B(n2190), .Z(n2189) );
  NANDN U2239 ( .A(A[976]), .B(n55), .Z(n2190) );
  NANDN U2240 ( .A(n55), .B(A[976]), .Z(n2188) );
  AND U2241 ( .A(n2191), .B(n2192), .Z(n55) );
  NAND U2242 ( .A(B[975]), .B(n2193), .Z(n2192) );
  NANDN U2243 ( .A(A[975]), .B(n57), .Z(n2193) );
  NANDN U2244 ( .A(n57), .B(A[975]), .Z(n2191) );
  AND U2245 ( .A(n2194), .B(n2195), .Z(n57) );
  NAND U2246 ( .A(B[974]), .B(n2196), .Z(n2195) );
  NANDN U2247 ( .A(A[974]), .B(n59), .Z(n2196) );
  NANDN U2248 ( .A(n59), .B(A[974]), .Z(n2194) );
  AND U2249 ( .A(n2197), .B(n2198), .Z(n59) );
  NAND U2250 ( .A(B[973]), .B(n2199), .Z(n2198) );
  NANDN U2251 ( .A(A[973]), .B(n61), .Z(n2199) );
  NANDN U2252 ( .A(n61), .B(A[973]), .Z(n2197) );
  AND U2253 ( .A(n2200), .B(n2201), .Z(n61) );
  NAND U2254 ( .A(B[972]), .B(n2202), .Z(n2201) );
  NANDN U2255 ( .A(A[972]), .B(n63), .Z(n2202) );
  NANDN U2256 ( .A(n63), .B(A[972]), .Z(n2200) );
  AND U2257 ( .A(n2203), .B(n2204), .Z(n63) );
  NAND U2258 ( .A(B[971]), .B(n2205), .Z(n2204) );
  NANDN U2259 ( .A(A[971]), .B(n65), .Z(n2205) );
  NANDN U2260 ( .A(n65), .B(A[971]), .Z(n2203) );
  AND U2261 ( .A(n2206), .B(n2207), .Z(n65) );
  NAND U2262 ( .A(B[970]), .B(n2208), .Z(n2207) );
  NANDN U2263 ( .A(A[970]), .B(n67), .Z(n2208) );
  NANDN U2264 ( .A(n67), .B(A[970]), .Z(n2206) );
  AND U2265 ( .A(n2209), .B(n2210), .Z(n67) );
  NAND U2266 ( .A(B[969]), .B(n2211), .Z(n2210) );
  NANDN U2267 ( .A(A[969]), .B(n71), .Z(n2211) );
  NANDN U2268 ( .A(n71), .B(A[969]), .Z(n2209) );
  AND U2269 ( .A(n2212), .B(n2213), .Z(n71) );
  NAND U2270 ( .A(B[968]), .B(n2214), .Z(n2213) );
  NANDN U2271 ( .A(A[968]), .B(n73), .Z(n2214) );
  NANDN U2272 ( .A(n73), .B(A[968]), .Z(n2212) );
  AND U2273 ( .A(n2215), .B(n2216), .Z(n73) );
  NAND U2274 ( .A(B[967]), .B(n2217), .Z(n2216) );
  NANDN U2275 ( .A(A[967]), .B(n75), .Z(n2217) );
  NANDN U2276 ( .A(n75), .B(A[967]), .Z(n2215) );
  AND U2277 ( .A(n2218), .B(n2219), .Z(n75) );
  NAND U2278 ( .A(B[966]), .B(n2220), .Z(n2219) );
  NANDN U2279 ( .A(A[966]), .B(n77), .Z(n2220) );
  NANDN U2280 ( .A(n77), .B(A[966]), .Z(n2218) );
  AND U2281 ( .A(n2221), .B(n2222), .Z(n77) );
  NAND U2282 ( .A(B[965]), .B(n2223), .Z(n2222) );
  NANDN U2283 ( .A(A[965]), .B(n79), .Z(n2223) );
  NANDN U2284 ( .A(n79), .B(A[965]), .Z(n2221) );
  AND U2285 ( .A(n2224), .B(n2225), .Z(n79) );
  NAND U2286 ( .A(B[964]), .B(n2226), .Z(n2225) );
  NANDN U2287 ( .A(A[964]), .B(n81), .Z(n2226) );
  NANDN U2288 ( .A(n81), .B(A[964]), .Z(n2224) );
  AND U2289 ( .A(n2227), .B(n2228), .Z(n81) );
  NAND U2290 ( .A(B[963]), .B(n2229), .Z(n2228) );
  NANDN U2291 ( .A(A[963]), .B(n83), .Z(n2229) );
  NANDN U2292 ( .A(n83), .B(A[963]), .Z(n2227) );
  AND U2293 ( .A(n2230), .B(n2231), .Z(n83) );
  NAND U2294 ( .A(B[962]), .B(n2232), .Z(n2231) );
  NANDN U2295 ( .A(A[962]), .B(n85), .Z(n2232) );
  NANDN U2296 ( .A(n85), .B(A[962]), .Z(n2230) );
  AND U2297 ( .A(n2233), .B(n2234), .Z(n85) );
  NAND U2298 ( .A(B[961]), .B(n2235), .Z(n2234) );
  NANDN U2299 ( .A(A[961]), .B(n87), .Z(n2235) );
  NANDN U2300 ( .A(n87), .B(A[961]), .Z(n2233) );
  AND U2301 ( .A(n2236), .B(n2237), .Z(n87) );
  NAND U2302 ( .A(B[960]), .B(n2238), .Z(n2237) );
  NANDN U2303 ( .A(A[960]), .B(n89), .Z(n2238) );
  NANDN U2304 ( .A(n89), .B(A[960]), .Z(n2236) );
  AND U2305 ( .A(n2239), .B(n2240), .Z(n89) );
  NAND U2306 ( .A(B[959]), .B(n2241), .Z(n2240) );
  NANDN U2307 ( .A(A[959]), .B(n93), .Z(n2241) );
  NANDN U2308 ( .A(n93), .B(A[959]), .Z(n2239) );
  AND U2309 ( .A(n2242), .B(n2243), .Z(n93) );
  NAND U2310 ( .A(B[958]), .B(n2244), .Z(n2243) );
  NANDN U2311 ( .A(A[958]), .B(n95), .Z(n2244) );
  NANDN U2312 ( .A(n95), .B(A[958]), .Z(n2242) );
  AND U2313 ( .A(n2245), .B(n2246), .Z(n95) );
  NAND U2314 ( .A(B[957]), .B(n2247), .Z(n2246) );
  NANDN U2315 ( .A(A[957]), .B(n97), .Z(n2247) );
  NANDN U2316 ( .A(n97), .B(A[957]), .Z(n2245) );
  AND U2317 ( .A(n2248), .B(n2249), .Z(n97) );
  NAND U2318 ( .A(B[956]), .B(n2250), .Z(n2249) );
  NANDN U2319 ( .A(A[956]), .B(n99), .Z(n2250) );
  NANDN U2320 ( .A(n99), .B(A[956]), .Z(n2248) );
  AND U2321 ( .A(n2251), .B(n2252), .Z(n99) );
  NAND U2322 ( .A(B[955]), .B(n2253), .Z(n2252) );
  NANDN U2323 ( .A(A[955]), .B(n101), .Z(n2253) );
  NANDN U2324 ( .A(n101), .B(A[955]), .Z(n2251) );
  AND U2325 ( .A(n2254), .B(n2255), .Z(n101) );
  NAND U2326 ( .A(B[954]), .B(n2256), .Z(n2255) );
  NANDN U2327 ( .A(A[954]), .B(n103), .Z(n2256) );
  NANDN U2328 ( .A(n103), .B(A[954]), .Z(n2254) );
  AND U2329 ( .A(n2257), .B(n2258), .Z(n103) );
  NAND U2330 ( .A(B[953]), .B(n2259), .Z(n2258) );
  NANDN U2331 ( .A(A[953]), .B(n105), .Z(n2259) );
  NANDN U2332 ( .A(n105), .B(A[953]), .Z(n2257) );
  AND U2333 ( .A(n2260), .B(n2261), .Z(n105) );
  NAND U2334 ( .A(B[952]), .B(n2262), .Z(n2261) );
  NANDN U2335 ( .A(A[952]), .B(n107), .Z(n2262) );
  NANDN U2336 ( .A(n107), .B(A[952]), .Z(n2260) );
  AND U2337 ( .A(n2263), .B(n2264), .Z(n107) );
  NAND U2338 ( .A(B[951]), .B(n2265), .Z(n2264) );
  NANDN U2339 ( .A(A[951]), .B(n109), .Z(n2265) );
  NANDN U2340 ( .A(n109), .B(A[951]), .Z(n2263) );
  AND U2341 ( .A(n2266), .B(n2267), .Z(n109) );
  NAND U2342 ( .A(B[950]), .B(n2268), .Z(n2267) );
  NANDN U2343 ( .A(A[950]), .B(n111), .Z(n2268) );
  NANDN U2344 ( .A(n111), .B(A[950]), .Z(n2266) );
  AND U2345 ( .A(n2269), .B(n2270), .Z(n111) );
  NAND U2346 ( .A(B[949]), .B(n2271), .Z(n2270) );
  NANDN U2347 ( .A(A[949]), .B(n115), .Z(n2271) );
  NANDN U2348 ( .A(n115), .B(A[949]), .Z(n2269) );
  AND U2349 ( .A(n2272), .B(n2273), .Z(n115) );
  NAND U2350 ( .A(B[948]), .B(n2274), .Z(n2273) );
  NANDN U2351 ( .A(A[948]), .B(n117), .Z(n2274) );
  NANDN U2352 ( .A(n117), .B(A[948]), .Z(n2272) );
  AND U2353 ( .A(n2275), .B(n2276), .Z(n117) );
  NAND U2354 ( .A(B[947]), .B(n2277), .Z(n2276) );
  NANDN U2355 ( .A(A[947]), .B(n119), .Z(n2277) );
  NANDN U2356 ( .A(n119), .B(A[947]), .Z(n2275) );
  AND U2357 ( .A(n2278), .B(n2279), .Z(n119) );
  NAND U2358 ( .A(B[946]), .B(n2280), .Z(n2279) );
  NANDN U2359 ( .A(A[946]), .B(n121), .Z(n2280) );
  NANDN U2360 ( .A(n121), .B(A[946]), .Z(n2278) );
  AND U2361 ( .A(n2281), .B(n2282), .Z(n121) );
  NAND U2362 ( .A(B[945]), .B(n2283), .Z(n2282) );
  NANDN U2363 ( .A(A[945]), .B(n123), .Z(n2283) );
  NANDN U2364 ( .A(n123), .B(A[945]), .Z(n2281) );
  AND U2365 ( .A(n2284), .B(n2285), .Z(n123) );
  NAND U2366 ( .A(B[944]), .B(n2286), .Z(n2285) );
  NANDN U2367 ( .A(A[944]), .B(n125), .Z(n2286) );
  NANDN U2368 ( .A(n125), .B(A[944]), .Z(n2284) );
  AND U2369 ( .A(n2287), .B(n2288), .Z(n125) );
  NAND U2370 ( .A(B[943]), .B(n2289), .Z(n2288) );
  NANDN U2371 ( .A(A[943]), .B(n127), .Z(n2289) );
  NANDN U2372 ( .A(n127), .B(A[943]), .Z(n2287) );
  AND U2373 ( .A(n2290), .B(n2291), .Z(n127) );
  NAND U2374 ( .A(B[942]), .B(n2292), .Z(n2291) );
  NANDN U2375 ( .A(A[942]), .B(n129), .Z(n2292) );
  NANDN U2376 ( .A(n129), .B(A[942]), .Z(n2290) );
  AND U2377 ( .A(n2293), .B(n2294), .Z(n129) );
  NAND U2378 ( .A(B[941]), .B(n2295), .Z(n2294) );
  NANDN U2379 ( .A(A[941]), .B(n131), .Z(n2295) );
  NANDN U2380 ( .A(n131), .B(A[941]), .Z(n2293) );
  AND U2381 ( .A(n2296), .B(n2297), .Z(n131) );
  NAND U2382 ( .A(B[940]), .B(n2298), .Z(n2297) );
  NANDN U2383 ( .A(A[940]), .B(n133), .Z(n2298) );
  NANDN U2384 ( .A(n133), .B(A[940]), .Z(n2296) );
  AND U2385 ( .A(n2299), .B(n2300), .Z(n133) );
  NAND U2386 ( .A(B[939]), .B(n2301), .Z(n2300) );
  NANDN U2387 ( .A(A[939]), .B(n137), .Z(n2301) );
  NANDN U2388 ( .A(n137), .B(A[939]), .Z(n2299) );
  AND U2389 ( .A(n2302), .B(n2303), .Z(n137) );
  NAND U2390 ( .A(B[938]), .B(n2304), .Z(n2303) );
  NANDN U2391 ( .A(A[938]), .B(n139), .Z(n2304) );
  NANDN U2392 ( .A(n139), .B(A[938]), .Z(n2302) );
  AND U2393 ( .A(n2305), .B(n2306), .Z(n139) );
  NAND U2394 ( .A(B[937]), .B(n2307), .Z(n2306) );
  NANDN U2395 ( .A(A[937]), .B(n141), .Z(n2307) );
  NANDN U2396 ( .A(n141), .B(A[937]), .Z(n2305) );
  AND U2397 ( .A(n2308), .B(n2309), .Z(n141) );
  NAND U2398 ( .A(B[936]), .B(n2310), .Z(n2309) );
  NANDN U2399 ( .A(A[936]), .B(n143), .Z(n2310) );
  NANDN U2400 ( .A(n143), .B(A[936]), .Z(n2308) );
  AND U2401 ( .A(n2311), .B(n2312), .Z(n143) );
  NAND U2402 ( .A(B[935]), .B(n2313), .Z(n2312) );
  NANDN U2403 ( .A(A[935]), .B(n145), .Z(n2313) );
  NANDN U2404 ( .A(n145), .B(A[935]), .Z(n2311) );
  AND U2405 ( .A(n2314), .B(n2315), .Z(n145) );
  NAND U2406 ( .A(B[934]), .B(n2316), .Z(n2315) );
  NANDN U2407 ( .A(A[934]), .B(n147), .Z(n2316) );
  NANDN U2408 ( .A(n147), .B(A[934]), .Z(n2314) );
  AND U2409 ( .A(n2317), .B(n2318), .Z(n147) );
  NAND U2410 ( .A(B[933]), .B(n2319), .Z(n2318) );
  NANDN U2411 ( .A(A[933]), .B(n149), .Z(n2319) );
  NANDN U2412 ( .A(n149), .B(A[933]), .Z(n2317) );
  AND U2413 ( .A(n2320), .B(n2321), .Z(n149) );
  NAND U2414 ( .A(B[932]), .B(n2322), .Z(n2321) );
  NANDN U2415 ( .A(A[932]), .B(n151), .Z(n2322) );
  NANDN U2416 ( .A(n151), .B(A[932]), .Z(n2320) );
  AND U2417 ( .A(n2323), .B(n2324), .Z(n151) );
  NAND U2418 ( .A(B[931]), .B(n2325), .Z(n2324) );
  NANDN U2419 ( .A(A[931]), .B(n153), .Z(n2325) );
  NANDN U2420 ( .A(n153), .B(A[931]), .Z(n2323) );
  AND U2421 ( .A(n2326), .B(n2327), .Z(n153) );
  NAND U2422 ( .A(B[930]), .B(n2328), .Z(n2327) );
  NANDN U2423 ( .A(A[930]), .B(n155), .Z(n2328) );
  NANDN U2424 ( .A(n155), .B(A[930]), .Z(n2326) );
  AND U2425 ( .A(n2329), .B(n2330), .Z(n155) );
  NAND U2426 ( .A(B[929]), .B(n2331), .Z(n2330) );
  NANDN U2427 ( .A(A[929]), .B(n159), .Z(n2331) );
  NANDN U2428 ( .A(n159), .B(A[929]), .Z(n2329) );
  AND U2429 ( .A(n2332), .B(n2333), .Z(n159) );
  NAND U2430 ( .A(B[928]), .B(n2334), .Z(n2333) );
  NANDN U2431 ( .A(A[928]), .B(n161), .Z(n2334) );
  NANDN U2432 ( .A(n161), .B(A[928]), .Z(n2332) );
  AND U2433 ( .A(n2335), .B(n2336), .Z(n161) );
  NAND U2434 ( .A(B[927]), .B(n2337), .Z(n2336) );
  NANDN U2435 ( .A(A[927]), .B(n163), .Z(n2337) );
  NANDN U2436 ( .A(n163), .B(A[927]), .Z(n2335) );
  AND U2437 ( .A(n2338), .B(n2339), .Z(n163) );
  NAND U2438 ( .A(B[926]), .B(n2340), .Z(n2339) );
  NANDN U2439 ( .A(A[926]), .B(n165), .Z(n2340) );
  NANDN U2440 ( .A(n165), .B(A[926]), .Z(n2338) );
  AND U2441 ( .A(n2341), .B(n2342), .Z(n165) );
  NAND U2442 ( .A(B[925]), .B(n2343), .Z(n2342) );
  NANDN U2443 ( .A(A[925]), .B(n167), .Z(n2343) );
  NANDN U2444 ( .A(n167), .B(A[925]), .Z(n2341) );
  AND U2445 ( .A(n2344), .B(n2345), .Z(n167) );
  NAND U2446 ( .A(B[924]), .B(n2346), .Z(n2345) );
  NANDN U2447 ( .A(A[924]), .B(n169), .Z(n2346) );
  NANDN U2448 ( .A(n169), .B(A[924]), .Z(n2344) );
  AND U2449 ( .A(n2347), .B(n2348), .Z(n169) );
  NAND U2450 ( .A(B[923]), .B(n2349), .Z(n2348) );
  NANDN U2451 ( .A(A[923]), .B(n171), .Z(n2349) );
  NANDN U2452 ( .A(n171), .B(A[923]), .Z(n2347) );
  AND U2453 ( .A(n2350), .B(n2351), .Z(n171) );
  NAND U2454 ( .A(B[922]), .B(n2352), .Z(n2351) );
  NANDN U2455 ( .A(A[922]), .B(n173), .Z(n2352) );
  NANDN U2456 ( .A(n173), .B(A[922]), .Z(n2350) );
  AND U2457 ( .A(n2353), .B(n2354), .Z(n173) );
  NAND U2458 ( .A(B[921]), .B(n2355), .Z(n2354) );
  NANDN U2459 ( .A(A[921]), .B(n175), .Z(n2355) );
  NANDN U2460 ( .A(n175), .B(A[921]), .Z(n2353) );
  AND U2461 ( .A(n2356), .B(n2357), .Z(n175) );
  NAND U2462 ( .A(B[920]), .B(n2358), .Z(n2357) );
  NANDN U2463 ( .A(A[920]), .B(n177), .Z(n2358) );
  NANDN U2464 ( .A(n177), .B(A[920]), .Z(n2356) );
  AND U2465 ( .A(n2359), .B(n2360), .Z(n177) );
  NAND U2466 ( .A(B[919]), .B(n2361), .Z(n2360) );
  NANDN U2467 ( .A(A[919]), .B(n181), .Z(n2361) );
  NANDN U2468 ( .A(n181), .B(A[919]), .Z(n2359) );
  AND U2469 ( .A(n2362), .B(n2363), .Z(n181) );
  NAND U2470 ( .A(B[918]), .B(n2364), .Z(n2363) );
  NANDN U2471 ( .A(A[918]), .B(n183), .Z(n2364) );
  NANDN U2472 ( .A(n183), .B(A[918]), .Z(n2362) );
  AND U2473 ( .A(n2365), .B(n2366), .Z(n183) );
  NAND U2474 ( .A(B[917]), .B(n2367), .Z(n2366) );
  NANDN U2475 ( .A(A[917]), .B(n185), .Z(n2367) );
  NANDN U2476 ( .A(n185), .B(A[917]), .Z(n2365) );
  AND U2477 ( .A(n2368), .B(n2369), .Z(n185) );
  NAND U2478 ( .A(B[916]), .B(n2370), .Z(n2369) );
  NANDN U2479 ( .A(A[916]), .B(n187), .Z(n2370) );
  NANDN U2480 ( .A(n187), .B(A[916]), .Z(n2368) );
  AND U2481 ( .A(n2371), .B(n2372), .Z(n187) );
  NAND U2482 ( .A(B[915]), .B(n2373), .Z(n2372) );
  NANDN U2483 ( .A(A[915]), .B(n189), .Z(n2373) );
  NANDN U2484 ( .A(n189), .B(A[915]), .Z(n2371) );
  AND U2485 ( .A(n2374), .B(n2375), .Z(n189) );
  NAND U2486 ( .A(B[914]), .B(n2376), .Z(n2375) );
  NANDN U2487 ( .A(A[914]), .B(n191), .Z(n2376) );
  NANDN U2488 ( .A(n191), .B(A[914]), .Z(n2374) );
  AND U2489 ( .A(n2377), .B(n2378), .Z(n191) );
  NAND U2490 ( .A(B[913]), .B(n2379), .Z(n2378) );
  NANDN U2491 ( .A(A[913]), .B(n193), .Z(n2379) );
  NANDN U2492 ( .A(n193), .B(A[913]), .Z(n2377) );
  AND U2493 ( .A(n2380), .B(n2381), .Z(n193) );
  NAND U2494 ( .A(B[912]), .B(n2382), .Z(n2381) );
  NANDN U2495 ( .A(A[912]), .B(n195), .Z(n2382) );
  NANDN U2496 ( .A(n195), .B(A[912]), .Z(n2380) );
  AND U2497 ( .A(n2383), .B(n2384), .Z(n195) );
  NAND U2498 ( .A(B[911]), .B(n2385), .Z(n2384) );
  NANDN U2499 ( .A(A[911]), .B(n197), .Z(n2385) );
  NANDN U2500 ( .A(n197), .B(A[911]), .Z(n2383) );
  AND U2501 ( .A(n2386), .B(n2387), .Z(n197) );
  NAND U2502 ( .A(B[910]), .B(n2388), .Z(n2387) );
  NANDN U2503 ( .A(A[910]), .B(n199), .Z(n2388) );
  NANDN U2504 ( .A(n199), .B(A[910]), .Z(n2386) );
  AND U2505 ( .A(n2389), .B(n2390), .Z(n199) );
  NAND U2506 ( .A(B[909]), .B(n2391), .Z(n2390) );
  NANDN U2507 ( .A(A[909]), .B(n203), .Z(n2391) );
  NANDN U2508 ( .A(n203), .B(A[909]), .Z(n2389) );
  AND U2509 ( .A(n2392), .B(n2393), .Z(n203) );
  NAND U2510 ( .A(B[908]), .B(n2394), .Z(n2393) );
  NANDN U2511 ( .A(A[908]), .B(n205), .Z(n2394) );
  NANDN U2512 ( .A(n205), .B(A[908]), .Z(n2392) );
  AND U2513 ( .A(n2395), .B(n2396), .Z(n205) );
  NAND U2514 ( .A(B[907]), .B(n2397), .Z(n2396) );
  NANDN U2515 ( .A(A[907]), .B(n207), .Z(n2397) );
  NANDN U2516 ( .A(n207), .B(A[907]), .Z(n2395) );
  AND U2517 ( .A(n2398), .B(n2399), .Z(n207) );
  NAND U2518 ( .A(B[906]), .B(n2400), .Z(n2399) );
  NANDN U2519 ( .A(A[906]), .B(n209), .Z(n2400) );
  NANDN U2520 ( .A(n209), .B(A[906]), .Z(n2398) );
  AND U2521 ( .A(n2401), .B(n2402), .Z(n209) );
  NAND U2522 ( .A(B[905]), .B(n2403), .Z(n2402) );
  NANDN U2523 ( .A(A[905]), .B(n211), .Z(n2403) );
  NANDN U2524 ( .A(n211), .B(A[905]), .Z(n2401) );
  AND U2525 ( .A(n2404), .B(n2405), .Z(n211) );
  NAND U2526 ( .A(B[904]), .B(n2406), .Z(n2405) );
  NANDN U2527 ( .A(A[904]), .B(n213), .Z(n2406) );
  NANDN U2528 ( .A(n213), .B(A[904]), .Z(n2404) );
  AND U2529 ( .A(n2407), .B(n2408), .Z(n213) );
  NAND U2530 ( .A(B[903]), .B(n2409), .Z(n2408) );
  NANDN U2531 ( .A(A[903]), .B(n215), .Z(n2409) );
  NANDN U2532 ( .A(n215), .B(A[903]), .Z(n2407) );
  AND U2533 ( .A(n2410), .B(n2411), .Z(n215) );
  NAND U2534 ( .A(B[902]), .B(n2412), .Z(n2411) );
  NANDN U2535 ( .A(A[902]), .B(n217), .Z(n2412) );
  NANDN U2536 ( .A(n217), .B(A[902]), .Z(n2410) );
  AND U2537 ( .A(n2413), .B(n2414), .Z(n217) );
  NAND U2538 ( .A(B[901]), .B(n2415), .Z(n2414) );
  NANDN U2539 ( .A(A[901]), .B(n219), .Z(n2415) );
  NANDN U2540 ( .A(n219), .B(A[901]), .Z(n2413) );
  AND U2541 ( .A(n2416), .B(n2417), .Z(n219) );
  NAND U2542 ( .A(B[900]), .B(n2418), .Z(n2417) );
  NANDN U2543 ( .A(A[900]), .B(n221), .Z(n2418) );
  NANDN U2544 ( .A(n221), .B(A[900]), .Z(n2416) );
  AND U2545 ( .A(n2419), .B(n2420), .Z(n221) );
  NAND U2546 ( .A(B[899]), .B(n2421), .Z(n2420) );
  NANDN U2547 ( .A(A[899]), .B(n227), .Z(n2421) );
  NANDN U2548 ( .A(n227), .B(A[899]), .Z(n2419) );
  AND U2549 ( .A(n2422), .B(n2423), .Z(n227) );
  NAND U2550 ( .A(B[898]), .B(n2424), .Z(n2423) );
  NANDN U2551 ( .A(A[898]), .B(n229), .Z(n2424) );
  NANDN U2552 ( .A(n229), .B(A[898]), .Z(n2422) );
  AND U2553 ( .A(n2425), .B(n2426), .Z(n229) );
  NAND U2554 ( .A(B[897]), .B(n2427), .Z(n2426) );
  NANDN U2555 ( .A(A[897]), .B(n231), .Z(n2427) );
  NANDN U2556 ( .A(n231), .B(A[897]), .Z(n2425) );
  AND U2557 ( .A(n2428), .B(n2429), .Z(n231) );
  NAND U2558 ( .A(B[896]), .B(n2430), .Z(n2429) );
  NANDN U2559 ( .A(A[896]), .B(n233), .Z(n2430) );
  NANDN U2560 ( .A(n233), .B(A[896]), .Z(n2428) );
  AND U2561 ( .A(n2431), .B(n2432), .Z(n233) );
  NAND U2562 ( .A(B[895]), .B(n2433), .Z(n2432) );
  NANDN U2563 ( .A(A[895]), .B(n235), .Z(n2433) );
  NANDN U2564 ( .A(n235), .B(A[895]), .Z(n2431) );
  AND U2565 ( .A(n2434), .B(n2435), .Z(n235) );
  NAND U2566 ( .A(B[894]), .B(n2436), .Z(n2435) );
  NANDN U2567 ( .A(A[894]), .B(n237), .Z(n2436) );
  NANDN U2568 ( .A(n237), .B(A[894]), .Z(n2434) );
  AND U2569 ( .A(n2437), .B(n2438), .Z(n237) );
  NAND U2570 ( .A(B[893]), .B(n2439), .Z(n2438) );
  NANDN U2571 ( .A(A[893]), .B(n239), .Z(n2439) );
  NANDN U2572 ( .A(n239), .B(A[893]), .Z(n2437) );
  AND U2573 ( .A(n2440), .B(n2441), .Z(n239) );
  NAND U2574 ( .A(B[892]), .B(n2442), .Z(n2441) );
  NANDN U2575 ( .A(A[892]), .B(n241), .Z(n2442) );
  NANDN U2576 ( .A(n241), .B(A[892]), .Z(n2440) );
  AND U2577 ( .A(n2443), .B(n2444), .Z(n241) );
  NAND U2578 ( .A(B[891]), .B(n2445), .Z(n2444) );
  NANDN U2579 ( .A(A[891]), .B(n243), .Z(n2445) );
  NANDN U2580 ( .A(n243), .B(A[891]), .Z(n2443) );
  AND U2581 ( .A(n2446), .B(n2447), .Z(n243) );
  NAND U2582 ( .A(B[890]), .B(n2448), .Z(n2447) );
  NANDN U2583 ( .A(A[890]), .B(n245), .Z(n2448) );
  NANDN U2584 ( .A(n245), .B(A[890]), .Z(n2446) );
  AND U2585 ( .A(n2449), .B(n2450), .Z(n245) );
  NAND U2586 ( .A(B[889]), .B(n2451), .Z(n2450) );
  NANDN U2587 ( .A(A[889]), .B(n249), .Z(n2451) );
  NANDN U2588 ( .A(n249), .B(A[889]), .Z(n2449) );
  AND U2589 ( .A(n2452), .B(n2453), .Z(n249) );
  NAND U2590 ( .A(B[888]), .B(n2454), .Z(n2453) );
  NANDN U2591 ( .A(A[888]), .B(n251), .Z(n2454) );
  NANDN U2592 ( .A(n251), .B(A[888]), .Z(n2452) );
  AND U2593 ( .A(n2455), .B(n2456), .Z(n251) );
  NAND U2594 ( .A(B[887]), .B(n2457), .Z(n2456) );
  NANDN U2595 ( .A(A[887]), .B(n253), .Z(n2457) );
  NANDN U2596 ( .A(n253), .B(A[887]), .Z(n2455) );
  AND U2597 ( .A(n2458), .B(n2459), .Z(n253) );
  NAND U2598 ( .A(B[886]), .B(n2460), .Z(n2459) );
  NANDN U2599 ( .A(A[886]), .B(n255), .Z(n2460) );
  NANDN U2600 ( .A(n255), .B(A[886]), .Z(n2458) );
  AND U2601 ( .A(n2461), .B(n2462), .Z(n255) );
  NAND U2602 ( .A(B[885]), .B(n2463), .Z(n2462) );
  NANDN U2603 ( .A(A[885]), .B(n257), .Z(n2463) );
  NANDN U2604 ( .A(n257), .B(A[885]), .Z(n2461) );
  AND U2605 ( .A(n2464), .B(n2465), .Z(n257) );
  NAND U2606 ( .A(B[884]), .B(n2466), .Z(n2465) );
  NANDN U2607 ( .A(A[884]), .B(n259), .Z(n2466) );
  NANDN U2608 ( .A(n259), .B(A[884]), .Z(n2464) );
  AND U2609 ( .A(n2467), .B(n2468), .Z(n259) );
  NAND U2610 ( .A(B[883]), .B(n2469), .Z(n2468) );
  NANDN U2611 ( .A(A[883]), .B(n261), .Z(n2469) );
  NANDN U2612 ( .A(n261), .B(A[883]), .Z(n2467) );
  AND U2613 ( .A(n2470), .B(n2471), .Z(n261) );
  NAND U2614 ( .A(B[882]), .B(n2472), .Z(n2471) );
  NANDN U2615 ( .A(A[882]), .B(n263), .Z(n2472) );
  NANDN U2616 ( .A(n263), .B(A[882]), .Z(n2470) );
  AND U2617 ( .A(n2473), .B(n2474), .Z(n263) );
  NAND U2618 ( .A(B[881]), .B(n2475), .Z(n2474) );
  NANDN U2619 ( .A(A[881]), .B(n265), .Z(n2475) );
  NANDN U2620 ( .A(n265), .B(A[881]), .Z(n2473) );
  AND U2621 ( .A(n2476), .B(n2477), .Z(n265) );
  NAND U2622 ( .A(B[880]), .B(n2478), .Z(n2477) );
  NANDN U2623 ( .A(A[880]), .B(n267), .Z(n2478) );
  NANDN U2624 ( .A(n267), .B(A[880]), .Z(n2476) );
  AND U2625 ( .A(n2479), .B(n2480), .Z(n267) );
  NAND U2626 ( .A(B[879]), .B(n2481), .Z(n2480) );
  NANDN U2627 ( .A(A[879]), .B(n271), .Z(n2481) );
  NANDN U2628 ( .A(n271), .B(A[879]), .Z(n2479) );
  AND U2629 ( .A(n2482), .B(n2483), .Z(n271) );
  NAND U2630 ( .A(B[878]), .B(n2484), .Z(n2483) );
  NANDN U2631 ( .A(A[878]), .B(n273), .Z(n2484) );
  NANDN U2632 ( .A(n273), .B(A[878]), .Z(n2482) );
  AND U2633 ( .A(n2485), .B(n2486), .Z(n273) );
  NAND U2634 ( .A(B[877]), .B(n2487), .Z(n2486) );
  NANDN U2635 ( .A(A[877]), .B(n275), .Z(n2487) );
  NANDN U2636 ( .A(n275), .B(A[877]), .Z(n2485) );
  AND U2637 ( .A(n2488), .B(n2489), .Z(n275) );
  NAND U2638 ( .A(B[876]), .B(n2490), .Z(n2489) );
  NANDN U2639 ( .A(A[876]), .B(n277), .Z(n2490) );
  NANDN U2640 ( .A(n277), .B(A[876]), .Z(n2488) );
  AND U2641 ( .A(n2491), .B(n2492), .Z(n277) );
  NAND U2642 ( .A(B[875]), .B(n2493), .Z(n2492) );
  NANDN U2643 ( .A(A[875]), .B(n279), .Z(n2493) );
  NANDN U2644 ( .A(n279), .B(A[875]), .Z(n2491) );
  AND U2645 ( .A(n2494), .B(n2495), .Z(n279) );
  NAND U2646 ( .A(B[874]), .B(n2496), .Z(n2495) );
  NANDN U2647 ( .A(A[874]), .B(n281), .Z(n2496) );
  NANDN U2648 ( .A(n281), .B(A[874]), .Z(n2494) );
  AND U2649 ( .A(n2497), .B(n2498), .Z(n281) );
  NAND U2650 ( .A(B[873]), .B(n2499), .Z(n2498) );
  NANDN U2651 ( .A(A[873]), .B(n283), .Z(n2499) );
  NANDN U2652 ( .A(n283), .B(A[873]), .Z(n2497) );
  AND U2653 ( .A(n2500), .B(n2501), .Z(n283) );
  NAND U2654 ( .A(B[872]), .B(n2502), .Z(n2501) );
  NANDN U2655 ( .A(A[872]), .B(n285), .Z(n2502) );
  NANDN U2656 ( .A(n285), .B(A[872]), .Z(n2500) );
  AND U2657 ( .A(n2503), .B(n2504), .Z(n285) );
  NAND U2658 ( .A(B[871]), .B(n2505), .Z(n2504) );
  NANDN U2659 ( .A(A[871]), .B(n287), .Z(n2505) );
  NANDN U2660 ( .A(n287), .B(A[871]), .Z(n2503) );
  AND U2661 ( .A(n2506), .B(n2507), .Z(n287) );
  NAND U2662 ( .A(B[870]), .B(n2508), .Z(n2507) );
  NANDN U2663 ( .A(A[870]), .B(n289), .Z(n2508) );
  NANDN U2664 ( .A(n289), .B(A[870]), .Z(n2506) );
  AND U2665 ( .A(n2509), .B(n2510), .Z(n289) );
  NAND U2666 ( .A(B[869]), .B(n2511), .Z(n2510) );
  NANDN U2667 ( .A(A[869]), .B(n293), .Z(n2511) );
  NANDN U2668 ( .A(n293), .B(A[869]), .Z(n2509) );
  AND U2669 ( .A(n2512), .B(n2513), .Z(n293) );
  NAND U2670 ( .A(B[868]), .B(n2514), .Z(n2513) );
  NANDN U2671 ( .A(A[868]), .B(n295), .Z(n2514) );
  NANDN U2672 ( .A(n295), .B(A[868]), .Z(n2512) );
  AND U2673 ( .A(n2515), .B(n2516), .Z(n295) );
  NAND U2674 ( .A(B[867]), .B(n2517), .Z(n2516) );
  NANDN U2675 ( .A(A[867]), .B(n297), .Z(n2517) );
  NANDN U2676 ( .A(n297), .B(A[867]), .Z(n2515) );
  AND U2677 ( .A(n2518), .B(n2519), .Z(n297) );
  NAND U2678 ( .A(B[866]), .B(n2520), .Z(n2519) );
  NANDN U2679 ( .A(A[866]), .B(n299), .Z(n2520) );
  NANDN U2680 ( .A(n299), .B(A[866]), .Z(n2518) );
  AND U2681 ( .A(n2521), .B(n2522), .Z(n299) );
  NAND U2682 ( .A(B[865]), .B(n2523), .Z(n2522) );
  NANDN U2683 ( .A(A[865]), .B(n301), .Z(n2523) );
  NANDN U2684 ( .A(n301), .B(A[865]), .Z(n2521) );
  AND U2685 ( .A(n2524), .B(n2525), .Z(n301) );
  NAND U2686 ( .A(B[864]), .B(n2526), .Z(n2525) );
  NANDN U2687 ( .A(A[864]), .B(n303), .Z(n2526) );
  NANDN U2688 ( .A(n303), .B(A[864]), .Z(n2524) );
  AND U2689 ( .A(n2527), .B(n2528), .Z(n303) );
  NAND U2690 ( .A(B[863]), .B(n2529), .Z(n2528) );
  NANDN U2691 ( .A(A[863]), .B(n305), .Z(n2529) );
  NANDN U2692 ( .A(n305), .B(A[863]), .Z(n2527) );
  AND U2693 ( .A(n2530), .B(n2531), .Z(n305) );
  NAND U2694 ( .A(B[862]), .B(n2532), .Z(n2531) );
  NANDN U2695 ( .A(A[862]), .B(n307), .Z(n2532) );
  NANDN U2696 ( .A(n307), .B(A[862]), .Z(n2530) );
  AND U2697 ( .A(n2533), .B(n2534), .Z(n307) );
  NAND U2698 ( .A(B[861]), .B(n2535), .Z(n2534) );
  NANDN U2699 ( .A(A[861]), .B(n309), .Z(n2535) );
  NANDN U2700 ( .A(n309), .B(A[861]), .Z(n2533) );
  AND U2701 ( .A(n2536), .B(n2537), .Z(n309) );
  NAND U2702 ( .A(B[860]), .B(n2538), .Z(n2537) );
  NANDN U2703 ( .A(A[860]), .B(n311), .Z(n2538) );
  NANDN U2704 ( .A(n311), .B(A[860]), .Z(n2536) );
  AND U2705 ( .A(n2539), .B(n2540), .Z(n311) );
  NAND U2706 ( .A(B[859]), .B(n2541), .Z(n2540) );
  NANDN U2707 ( .A(A[859]), .B(n315), .Z(n2541) );
  NANDN U2708 ( .A(n315), .B(A[859]), .Z(n2539) );
  AND U2709 ( .A(n2542), .B(n2543), .Z(n315) );
  NAND U2710 ( .A(B[858]), .B(n2544), .Z(n2543) );
  NANDN U2711 ( .A(A[858]), .B(n317), .Z(n2544) );
  NANDN U2712 ( .A(n317), .B(A[858]), .Z(n2542) );
  AND U2713 ( .A(n2545), .B(n2546), .Z(n317) );
  NAND U2714 ( .A(B[857]), .B(n2547), .Z(n2546) );
  NANDN U2715 ( .A(A[857]), .B(n319), .Z(n2547) );
  NANDN U2716 ( .A(n319), .B(A[857]), .Z(n2545) );
  AND U2717 ( .A(n2548), .B(n2549), .Z(n319) );
  NAND U2718 ( .A(B[856]), .B(n2550), .Z(n2549) );
  NANDN U2719 ( .A(A[856]), .B(n321), .Z(n2550) );
  NANDN U2720 ( .A(n321), .B(A[856]), .Z(n2548) );
  AND U2721 ( .A(n2551), .B(n2552), .Z(n321) );
  NAND U2722 ( .A(B[855]), .B(n2553), .Z(n2552) );
  NANDN U2723 ( .A(A[855]), .B(n323), .Z(n2553) );
  NANDN U2724 ( .A(n323), .B(A[855]), .Z(n2551) );
  AND U2725 ( .A(n2554), .B(n2555), .Z(n323) );
  NAND U2726 ( .A(B[854]), .B(n2556), .Z(n2555) );
  NANDN U2727 ( .A(A[854]), .B(n325), .Z(n2556) );
  NANDN U2728 ( .A(n325), .B(A[854]), .Z(n2554) );
  AND U2729 ( .A(n2557), .B(n2558), .Z(n325) );
  NAND U2730 ( .A(B[853]), .B(n2559), .Z(n2558) );
  NANDN U2731 ( .A(A[853]), .B(n327), .Z(n2559) );
  NANDN U2732 ( .A(n327), .B(A[853]), .Z(n2557) );
  AND U2733 ( .A(n2560), .B(n2561), .Z(n327) );
  NAND U2734 ( .A(B[852]), .B(n2562), .Z(n2561) );
  NANDN U2735 ( .A(A[852]), .B(n329), .Z(n2562) );
  NANDN U2736 ( .A(n329), .B(A[852]), .Z(n2560) );
  AND U2737 ( .A(n2563), .B(n2564), .Z(n329) );
  NAND U2738 ( .A(B[851]), .B(n2565), .Z(n2564) );
  NANDN U2739 ( .A(A[851]), .B(n331), .Z(n2565) );
  NANDN U2740 ( .A(n331), .B(A[851]), .Z(n2563) );
  AND U2741 ( .A(n2566), .B(n2567), .Z(n331) );
  NAND U2742 ( .A(B[850]), .B(n2568), .Z(n2567) );
  NANDN U2743 ( .A(A[850]), .B(n333), .Z(n2568) );
  NANDN U2744 ( .A(n333), .B(A[850]), .Z(n2566) );
  AND U2745 ( .A(n2569), .B(n2570), .Z(n333) );
  NAND U2746 ( .A(B[849]), .B(n2571), .Z(n2570) );
  NANDN U2747 ( .A(A[849]), .B(n337), .Z(n2571) );
  NANDN U2748 ( .A(n337), .B(A[849]), .Z(n2569) );
  AND U2749 ( .A(n2572), .B(n2573), .Z(n337) );
  NAND U2750 ( .A(B[848]), .B(n2574), .Z(n2573) );
  NANDN U2751 ( .A(A[848]), .B(n339), .Z(n2574) );
  NANDN U2752 ( .A(n339), .B(A[848]), .Z(n2572) );
  AND U2753 ( .A(n2575), .B(n2576), .Z(n339) );
  NAND U2754 ( .A(B[847]), .B(n2577), .Z(n2576) );
  NANDN U2755 ( .A(A[847]), .B(n341), .Z(n2577) );
  NANDN U2756 ( .A(n341), .B(A[847]), .Z(n2575) );
  AND U2757 ( .A(n2578), .B(n2579), .Z(n341) );
  NAND U2758 ( .A(B[846]), .B(n2580), .Z(n2579) );
  NANDN U2759 ( .A(A[846]), .B(n343), .Z(n2580) );
  NANDN U2760 ( .A(n343), .B(A[846]), .Z(n2578) );
  AND U2761 ( .A(n2581), .B(n2582), .Z(n343) );
  NAND U2762 ( .A(B[845]), .B(n2583), .Z(n2582) );
  NANDN U2763 ( .A(A[845]), .B(n345), .Z(n2583) );
  NANDN U2764 ( .A(n345), .B(A[845]), .Z(n2581) );
  AND U2765 ( .A(n2584), .B(n2585), .Z(n345) );
  NAND U2766 ( .A(B[844]), .B(n2586), .Z(n2585) );
  NANDN U2767 ( .A(A[844]), .B(n347), .Z(n2586) );
  NANDN U2768 ( .A(n347), .B(A[844]), .Z(n2584) );
  AND U2769 ( .A(n2587), .B(n2588), .Z(n347) );
  NAND U2770 ( .A(B[843]), .B(n2589), .Z(n2588) );
  NANDN U2771 ( .A(A[843]), .B(n349), .Z(n2589) );
  NANDN U2772 ( .A(n349), .B(A[843]), .Z(n2587) );
  AND U2773 ( .A(n2590), .B(n2591), .Z(n349) );
  NAND U2774 ( .A(B[842]), .B(n2592), .Z(n2591) );
  NANDN U2775 ( .A(A[842]), .B(n351), .Z(n2592) );
  NANDN U2776 ( .A(n351), .B(A[842]), .Z(n2590) );
  AND U2777 ( .A(n2593), .B(n2594), .Z(n351) );
  NAND U2778 ( .A(B[841]), .B(n2595), .Z(n2594) );
  NANDN U2779 ( .A(A[841]), .B(n353), .Z(n2595) );
  NANDN U2780 ( .A(n353), .B(A[841]), .Z(n2593) );
  AND U2781 ( .A(n2596), .B(n2597), .Z(n353) );
  NAND U2782 ( .A(B[840]), .B(n2598), .Z(n2597) );
  NANDN U2783 ( .A(A[840]), .B(n355), .Z(n2598) );
  NANDN U2784 ( .A(n355), .B(A[840]), .Z(n2596) );
  AND U2785 ( .A(n2599), .B(n2600), .Z(n355) );
  NAND U2786 ( .A(B[839]), .B(n2601), .Z(n2600) );
  NANDN U2787 ( .A(A[839]), .B(n359), .Z(n2601) );
  NANDN U2788 ( .A(n359), .B(A[839]), .Z(n2599) );
  AND U2789 ( .A(n2602), .B(n2603), .Z(n359) );
  NAND U2790 ( .A(B[838]), .B(n2604), .Z(n2603) );
  NANDN U2791 ( .A(A[838]), .B(n361), .Z(n2604) );
  NANDN U2792 ( .A(n361), .B(A[838]), .Z(n2602) );
  AND U2793 ( .A(n2605), .B(n2606), .Z(n361) );
  NAND U2794 ( .A(B[837]), .B(n2607), .Z(n2606) );
  NANDN U2795 ( .A(A[837]), .B(n363), .Z(n2607) );
  NANDN U2796 ( .A(n363), .B(A[837]), .Z(n2605) );
  AND U2797 ( .A(n2608), .B(n2609), .Z(n363) );
  NAND U2798 ( .A(B[836]), .B(n2610), .Z(n2609) );
  NANDN U2799 ( .A(A[836]), .B(n365), .Z(n2610) );
  NANDN U2800 ( .A(n365), .B(A[836]), .Z(n2608) );
  AND U2801 ( .A(n2611), .B(n2612), .Z(n365) );
  NAND U2802 ( .A(B[835]), .B(n2613), .Z(n2612) );
  NANDN U2803 ( .A(A[835]), .B(n367), .Z(n2613) );
  NANDN U2804 ( .A(n367), .B(A[835]), .Z(n2611) );
  AND U2805 ( .A(n2614), .B(n2615), .Z(n367) );
  NAND U2806 ( .A(B[834]), .B(n2616), .Z(n2615) );
  NANDN U2807 ( .A(A[834]), .B(n369), .Z(n2616) );
  NANDN U2808 ( .A(n369), .B(A[834]), .Z(n2614) );
  AND U2809 ( .A(n2617), .B(n2618), .Z(n369) );
  NAND U2810 ( .A(B[833]), .B(n2619), .Z(n2618) );
  NANDN U2811 ( .A(A[833]), .B(n371), .Z(n2619) );
  NANDN U2812 ( .A(n371), .B(A[833]), .Z(n2617) );
  AND U2813 ( .A(n2620), .B(n2621), .Z(n371) );
  NAND U2814 ( .A(B[832]), .B(n2622), .Z(n2621) );
  NANDN U2815 ( .A(A[832]), .B(n373), .Z(n2622) );
  NANDN U2816 ( .A(n373), .B(A[832]), .Z(n2620) );
  AND U2817 ( .A(n2623), .B(n2624), .Z(n373) );
  NAND U2818 ( .A(B[831]), .B(n2625), .Z(n2624) );
  NANDN U2819 ( .A(A[831]), .B(n375), .Z(n2625) );
  NANDN U2820 ( .A(n375), .B(A[831]), .Z(n2623) );
  AND U2821 ( .A(n2626), .B(n2627), .Z(n375) );
  NAND U2822 ( .A(B[830]), .B(n2628), .Z(n2627) );
  NANDN U2823 ( .A(A[830]), .B(n377), .Z(n2628) );
  NANDN U2824 ( .A(n377), .B(A[830]), .Z(n2626) );
  AND U2825 ( .A(n2629), .B(n2630), .Z(n377) );
  NAND U2826 ( .A(B[829]), .B(n2631), .Z(n2630) );
  NANDN U2827 ( .A(A[829]), .B(n381), .Z(n2631) );
  NANDN U2828 ( .A(n381), .B(A[829]), .Z(n2629) );
  AND U2829 ( .A(n2632), .B(n2633), .Z(n381) );
  NAND U2830 ( .A(B[828]), .B(n2634), .Z(n2633) );
  NANDN U2831 ( .A(A[828]), .B(n383), .Z(n2634) );
  NANDN U2832 ( .A(n383), .B(A[828]), .Z(n2632) );
  AND U2833 ( .A(n2635), .B(n2636), .Z(n383) );
  NAND U2834 ( .A(B[827]), .B(n2637), .Z(n2636) );
  NANDN U2835 ( .A(A[827]), .B(n385), .Z(n2637) );
  NANDN U2836 ( .A(n385), .B(A[827]), .Z(n2635) );
  AND U2837 ( .A(n2638), .B(n2639), .Z(n385) );
  NAND U2838 ( .A(B[826]), .B(n2640), .Z(n2639) );
  NANDN U2839 ( .A(A[826]), .B(n387), .Z(n2640) );
  NANDN U2840 ( .A(n387), .B(A[826]), .Z(n2638) );
  AND U2841 ( .A(n2641), .B(n2642), .Z(n387) );
  NAND U2842 ( .A(B[825]), .B(n2643), .Z(n2642) );
  NANDN U2843 ( .A(A[825]), .B(n389), .Z(n2643) );
  NANDN U2844 ( .A(n389), .B(A[825]), .Z(n2641) );
  AND U2845 ( .A(n2644), .B(n2645), .Z(n389) );
  NAND U2846 ( .A(B[824]), .B(n2646), .Z(n2645) );
  NANDN U2847 ( .A(A[824]), .B(n391), .Z(n2646) );
  NANDN U2848 ( .A(n391), .B(A[824]), .Z(n2644) );
  AND U2849 ( .A(n2647), .B(n2648), .Z(n391) );
  NAND U2850 ( .A(B[823]), .B(n2649), .Z(n2648) );
  NANDN U2851 ( .A(A[823]), .B(n393), .Z(n2649) );
  NANDN U2852 ( .A(n393), .B(A[823]), .Z(n2647) );
  AND U2853 ( .A(n2650), .B(n2651), .Z(n393) );
  NAND U2854 ( .A(B[822]), .B(n2652), .Z(n2651) );
  NANDN U2855 ( .A(A[822]), .B(n395), .Z(n2652) );
  NANDN U2856 ( .A(n395), .B(A[822]), .Z(n2650) );
  AND U2857 ( .A(n2653), .B(n2654), .Z(n395) );
  NAND U2858 ( .A(B[821]), .B(n2655), .Z(n2654) );
  NANDN U2859 ( .A(A[821]), .B(n397), .Z(n2655) );
  NANDN U2860 ( .A(n397), .B(A[821]), .Z(n2653) );
  AND U2861 ( .A(n2656), .B(n2657), .Z(n397) );
  NAND U2862 ( .A(B[820]), .B(n2658), .Z(n2657) );
  NANDN U2863 ( .A(A[820]), .B(n399), .Z(n2658) );
  NANDN U2864 ( .A(n399), .B(A[820]), .Z(n2656) );
  AND U2865 ( .A(n2659), .B(n2660), .Z(n399) );
  NAND U2866 ( .A(B[819]), .B(n2661), .Z(n2660) );
  NANDN U2867 ( .A(A[819]), .B(n403), .Z(n2661) );
  NANDN U2868 ( .A(n403), .B(A[819]), .Z(n2659) );
  AND U2869 ( .A(n2662), .B(n2663), .Z(n403) );
  NAND U2870 ( .A(B[818]), .B(n2664), .Z(n2663) );
  NANDN U2871 ( .A(A[818]), .B(n405), .Z(n2664) );
  NANDN U2872 ( .A(n405), .B(A[818]), .Z(n2662) );
  AND U2873 ( .A(n2665), .B(n2666), .Z(n405) );
  NAND U2874 ( .A(B[817]), .B(n2667), .Z(n2666) );
  NANDN U2875 ( .A(A[817]), .B(n407), .Z(n2667) );
  NANDN U2876 ( .A(n407), .B(A[817]), .Z(n2665) );
  AND U2877 ( .A(n2668), .B(n2669), .Z(n407) );
  NAND U2878 ( .A(B[816]), .B(n2670), .Z(n2669) );
  NANDN U2879 ( .A(A[816]), .B(n409), .Z(n2670) );
  NANDN U2880 ( .A(n409), .B(A[816]), .Z(n2668) );
  AND U2881 ( .A(n2671), .B(n2672), .Z(n409) );
  NAND U2882 ( .A(B[815]), .B(n2673), .Z(n2672) );
  NANDN U2883 ( .A(A[815]), .B(n411), .Z(n2673) );
  NANDN U2884 ( .A(n411), .B(A[815]), .Z(n2671) );
  AND U2885 ( .A(n2674), .B(n2675), .Z(n411) );
  NAND U2886 ( .A(B[814]), .B(n2676), .Z(n2675) );
  NANDN U2887 ( .A(A[814]), .B(n413), .Z(n2676) );
  NANDN U2888 ( .A(n413), .B(A[814]), .Z(n2674) );
  AND U2889 ( .A(n2677), .B(n2678), .Z(n413) );
  NAND U2890 ( .A(B[813]), .B(n2679), .Z(n2678) );
  NANDN U2891 ( .A(A[813]), .B(n415), .Z(n2679) );
  NANDN U2892 ( .A(n415), .B(A[813]), .Z(n2677) );
  AND U2893 ( .A(n2680), .B(n2681), .Z(n415) );
  NAND U2894 ( .A(B[812]), .B(n2682), .Z(n2681) );
  NANDN U2895 ( .A(A[812]), .B(n417), .Z(n2682) );
  NANDN U2896 ( .A(n417), .B(A[812]), .Z(n2680) );
  AND U2897 ( .A(n2683), .B(n2684), .Z(n417) );
  NAND U2898 ( .A(B[811]), .B(n2685), .Z(n2684) );
  NANDN U2899 ( .A(A[811]), .B(n419), .Z(n2685) );
  NANDN U2900 ( .A(n419), .B(A[811]), .Z(n2683) );
  AND U2901 ( .A(n2686), .B(n2687), .Z(n419) );
  NAND U2902 ( .A(B[810]), .B(n2688), .Z(n2687) );
  NANDN U2903 ( .A(A[810]), .B(n421), .Z(n2688) );
  NANDN U2904 ( .A(n421), .B(A[810]), .Z(n2686) );
  AND U2905 ( .A(n2689), .B(n2690), .Z(n421) );
  NAND U2906 ( .A(B[809]), .B(n2691), .Z(n2690) );
  NANDN U2907 ( .A(A[809]), .B(n425), .Z(n2691) );
  NANDN U2908 ( .A(n425), .B(A[809]), .Z(n2689) );
  AND U2909 ( .A(n2692), .B(n2693), .Z(n425) );
  NAND U2910 ( .A(B[808]), .B(n2694), .Z(n2693) );
  NANDN U2911 ( .A(A[808]), .B(n427), .Z(n2694) );
  NANDN U2912 ( .A(n427), .B(A[808]), .Z(n2692) );
  AND U2913 ( .A(n2695), .B(n2696), .Z(n427) );
  NAND U2914 ( .A(B[807]), .B(n2697), .Z(n2696) );
  NANDN U2915 ( .A(A[807]), .B(n429), .Z(n2697) );
  NANDN U2916 ( .A(n429), .B(A[807]), .Z(n2695) );
  AND U2917 ( .A(n2698), .B(n2699), .Z(n429) );
  NAND U2918 ( .A(B[806]), .B(n2700), .Z(n2699) );
  NANDN U2919 ( .A(A[806]), .B(n431), .Z(n2700) );
  NANDN U2920 ( .A(n431), .B(A[806]), .Z(n2698) );
  AND U2921 ( .A(n2701), .B(n2702), .Z(n431) );
  NAND U2922 ( .A(B[805]), .B(n2703), .Z(n2702) );
  NANDN U2923 ( .A(A[805]), .B(n433), .Z(n2703) );
  NANDN U2924 ( .A(n433), .B(A[805]), .Z(n2701) );
  AND U2925 ( .A(n2704), .B(n2705), .Z(n433) );
  NAND U2926 ( .A(B[804]), .B(n2706), .Z(n2705) );
  NANDN U2927 ( .A(A[804]), .B(n435), .Z(n2706) );
  NANDN U2928 ( .A(n435), .B(A[804]), .Z(n2704) );
  AND U2929 ( .A(n2707), .B(n2708), .Z(n435) );
  NAND U2930 ( .A(B[803]), .B(n2709), .Z(n2708) );
  NANDN U2931 ( .A(A[803]), .B(n437), .Z(n2709) );
  NANDN U2932 ( .A(n437), .B(A[803]), .Z(n2707) );
  AND U2933 ( .A(n2710), .B(n2711), .Z(n437) );
  NAND U2934 ( .A(B[802]), .B(n2712), .Z(n2711) );
  NANDN U2935 ( .A(A[802]), .B(n439), .Z(n2712) );
  NANDN U2936 ( .A(n439), .B(A[802]), .Z(n2710) );
  AND U2937 ( .A(n2713), .B(n2714), .Z(n439) );
  NAND U2938 ( .A(B[801]), .B(n2715), .Z(n2714) );
  NANDN U2939 ( .A(A[801]), .B(n441), .Z(n2715) );
  NANDN U2940 ( .A(n441), .B(A[801]), .Z(n2713) );
  AND U2941 ( .A(n2716), .B(n2717), .Z(n441) );
  NAND U2942 ( .A(B[800]), .B(n2718), .Z(n2717) );
  NANDN U2943 ( .A(A[800]), .B(n443), .Z(n2718) );
  NANDN U2944 ( .A(n443), .B(A[800]), .Z(n2716) );
  AND U2945 ( .A(n2719), .B(n2720), .Z(n443) );
  NAND U2946 ( .A(B[799]), .B(n2721), .Z(n2720) );
  NANDN U2947 ( .A(A[799]), .B(n449), .Z(n2721) );
  NANDN U2948 ( .A(n449), .B(A[799]), .Z(n2719) );
  AND U2949 ( .A(n2722), .B(n2723), .Z(n449) );
  NAND U2950 ( .A(B[798]), .B(n2724), .Z(n2723) );
  NANDN U2951 ( .A(A[798]), .B(n451), .Z(n2724) );
  NANDN U2952 ( .A(n451), .B(A[798]), .Z(n2722) );
  AND U2953 ( .A(n2725), .B(n2726), .Z(n451) );
  NAND U2954 ( .A(B[797]), .B(n2727), .Z(n2726) );
  NANDN U2955 ( .A(A[797]), .B(n453), .Z(n2727) );
  NANDN U2956 ( .A(n453), .B(A[797]), .Z(n2725) );
  AND U2957 ( .A(n2728), .B(n2729), .Z(n453) );
  NAND U2958 ( .A(B[796]), .B(n2730), .Z(n2729) );
  NANDN U2959 ( .A(A[796]), .B(n455), .Z(n2730) );
  NANDN U2960 ( .A(n455), .B(A[796]), .Z(n2728) );
  AND U2961 ( .A(n2731), .B(n2732), .Z(n455) );
  NAND U2962 ( .A(B[795]), .B(n2733), .Z(n2732) );
  NANDN U2963 ( .A(A[795]), .B(n457), .Z(n2733) );
  NANDN U2964 ( .A(n457), .B(A[795]), .Z(n2731) );
  AND U2965 ( .A(n2734), .B(n2735), .Z(n457) );
  NAND U2966 ( .A(B[794]), .B(n2736), .Z(n2735) );
  NANDN U2967 ( .A(A[794]), .B(n459), .Z(n2736) );
  NANDN U2968 ( .A(n459), .B(A[794]), .Z(n2734) );
  AND U2969 ( .A(n2737), .B(n2738), .Z(n459) );
  NAND U2970 ( .A(B[793]), .B(n2739), .Z(n2738) );
  NANDN U2971 ( .A(A[793]), .B(n461), .Z(n2739) );
  NANDN U2972 ( .A(n461), .B(A[793]), .Z(n2737) );
  AND U2973 ( .A(n2740), .B(n2741), .Z(n461) );
  NAND U2974 ( .A(B[792]), .B(n2742), .Z(n2741) );
  NANDN U2975 ( .A(A[792]), .B(n463), .Z(n2742) );
  NANDN U2976 ( .A(n463), .B(A[792]), .Z(n2740) );
  AND U2977 ( .A(n2743), .B(n2744), .Z(n463) );
  NAND U2978 ( .A(B[791]), .B(n2745), .Z(n2744) );
  NANDN U2979 ( .A(A[791]), .B(n465), .Z(n2745) );
  NANDN U2980 ( .A(n465), .B(A[791]), .Z(n2743) );
  AND U2981 ( .A(n2746), .B(n2747), .Z(n465) );
  NAND U2982 ( .A(B[790]), .B(n2748), .Z(n2747) );
  NANDN U2983 ( .A(A[790]), .B(n467), .Z(n2748) );
  NANDN U2984 ( .A(n467), .B(A[790]), .Z(n2746) );
  AND U2985 ( .A(n2749), .B(n2750), .Z(n467) );
  NAND U2986 ( .A(B[789]), .B(n2751), .Z(n2750) );
  NANDN U2987 ( .A(A[789]), .B(n471), .Z(n2751) );
  NANDN U2988 ( .A(n471), .B(A[789]), .Z(n2749) );
  AND U2989 ( .A(n2752), .B(n2753), .Z(n471) );
  NAND U2990 ( .A(B[788]), .B(n2754), .Z(n2753) );
  NANDN U2991 ( .A(A[788]), .B(n473), .Z(n2754) );
  NANDN U2992 ( .A(n473), .B(A[788]), .Z(n2752) );
  AND U2993 ( .A(n2755), .B(n2756), .Z(n473) );
  NAND U2994 ( .A(B[787]), .B(n2757), .Z(n2756) );
  NANDN U2995 ( .A(A[787]), .B(n475), .Z(n2757) );
  NANDN U2996 ( .A(n475), .B(A[787]), .Z(n2755) );
  AND U2997 ( .A(n2758), .B(n2759), .Z(n475) );
  NAND U2998 ( .A(B[786]), .B(n2760), .Z(n2759) );
  NANDN U2999 ( .A(A[786]), .B(n477), .Z(n2760) );
  NANDN U3000 ( .A(n477), .B(A[786]), .Z(n2758) );
  AND U3001 ( .A(n2761), .B(n2762), .Z(n477) );
  NAND U3002 ( .A(B[785]), .B(n2763), .Z(n2762) );
  NANDN U3003 ( .A(A[785]), .B(n479), .Z(n2763) );
  NANDN U3004 ( .A(n479), .B(A[785]), .Z(n2761) );
  AND U3005 ( .A(n2764), .B(n2765), .Z(n479) );
  NAND U3006 ( .A(B[784]), .B(n2766), .Z(n2765) );
  NANDN U3007 ( .A(A[784]), .B(n481), .Z(n2766) );
  NANDN U3008 ( .A(n481), .B(A[784]), .Z(n2764) );
  AND U3009 ( .A(n2767), .B(n2768), .Z(n481) );
  NAND U3010 ( .A(B[783]), .B(n2769), .Z(n2768) );
  NANDN U3011 ( .A(A[783]), .B(n483), .Z(n2769) );
  NANDN U3012 ( .A(n483), .B(A[783]), .Z(n2767) );
  AND U3013 ( .A(n2770), .B(n2771), .Z(n483) );
  NAND U3014 ( .A(B[782]), .B(n2772), .Z(n2771) );
  NANDN U3015 ( .A(A[782]), .B(n485), .Z(n2772) );
  NANDN U3016 ( .A(n485), .B(A[782]), .Z(n2770) );
  AND U3017 ( .A(n2773), .B(n2774), .Z(n485) );
  NAND U3018 ( .A(B[781]), .B(n2775), .Z(n2774) );
  NANDN U3019 ( .A(A[781]), .B(n487), .Z(n2775) );
  NANDN U3020 ( .A(n487), .B(A[781]), .Z(n2773) );
  AND U3021 ( .A(n2776), .B(n2777), .Z(n487) );
  NAND U3022 ( .A(B[780]), .B(n2778), .Z(n2777) );
  NANDN U3023 ( .A(A[780]), .B(n489), .Z(n2778) );
  NANDN U3024 ( .A(n489), .B(A[780]), .Z(n2776) );
  AND U3025 ( .A(n2779), .B(n2780), .Z(n489) );
  NAND U3026 ( .A(B[779]), .B(n2781), .Z(n2780) );
  NANDN U3027 ( .A(A[779]), .B(n493), .Z(n2781) );
  NANDN U3028 ( .A(n493), .B(A[779]), .Z(n2779) );
  AND U3029 ( .A(n2782), .B(n2783), .Z(n493) );
  NAND U3030 ( .A(B[778]), .B(n2784), .Z(n2783) );
  NANDN U3031 ( .A(A[778]), .B(n495), .Z(n2784) );
  NANDN U3032 ( .A(n495), .B(A[778]), .Z(n2782) );
  AND U3033 ( .A(n2785), .B(n2786), .Z(n495) );
  NAND U3034 ( .A(B[777]), .B(n2787), .Z(n2786) );
  NANDN U3035 ( .A(A[777]), .B(n497), .Z(n2787) );
  NANDN U3036 ( .A(n497), .B(A[777]), .Z(n2785) );
  AND U3037 ( .A(n2788), .B(n2789), .Z(n497) );
  NAND U3038 ( .A(B[776]), .B(n2790), .Z(n2789) );
  NANDN U3039 ( .A(A[776]), .B(n499), .Z(n2790) );
  NANDN U3040 ( .A(n499), .B(A[776]), .Z(n2788) );
  AND U3041 ( .A(n2791), .B(n2792), .Z(n499) );
  NAND U3042 ( .A(B[775]), .B(n2793), .Z(n2792) );
  NANDN U3043 ( .A(A[775]), .B(n501), .Z(n2793) );
  NANDN U3044 ( .A(n501), .B(A[775]), .Z(n2791) );
  AND U3045 ( .A(n2794), .B(n2795), .Z(n501) );
  NAND U3046 ( .A(B[774]), .B(n2796), .Z(n2795) );
  NANDN U3047 ( .A(A[774]), .B(n503), .Z(n2796) );
  NANDN U3048 ( .A(n503), .B(A[774]), .Z(n2794) );
  AND U3049 ( .A(n2797), .B(n2798), .Z(n503) );
  NAND U3050 ( .A(B[773]), .B(n2799), .Z(n2798) );
  NANDN U3051 ( .A(A[773]), .B(n505), .Z(n2799) );
  NANDN U3052 ( .A(n505), .B(A[773]), .Z(n2797) );
  AND U3053 ( .A(n2800), .B(n2801), .Z(n505) );
  NAND U3054 ( .A(B[772]), .B(n2802), .Z(n2801) );
  NANDN U3055 ( .A(A[772]), .B(n507), .Z(n2802) );
  NANDN U3056 ( .A(n507), .B(A[772]), .Z(n2800) );
  AND U3057 ( .A(n2803), .B(n2804), .Z(n507) );
  NAND U3058 ( .A(B[771]), .B(n2805), .Z(n2804) );
  NANDN U3059 ( .A(A[771]), .B(n509), .Z(n2805) );
  NANDN U3060 ( .A(n509), .B(A[771]), .Z(n2803) );
  AND U3061 ( .A(n2806), .B(n2807), .Z(n509) );
  NAND U3062 ( .A(B[770]), .B(n2808), .Z(n2807) );
  NANDN U3063 ( .A(A[770]), .B(n511), .Z(n2808) );
  NANDN U3064 ( .A(n511), .B(A[770]), .Z(n2806) );
  AND U3065 ( .A(n2809), .B(n2810), .Z(n511) );
  NAND U3066 ( .A(B[769]), .B(n2811), .Z(n2810) );
  NANDN U3067 ( .A(A[769]), .B(n515), .Z(n2811) );
  NANDN U3068 ( .A(n515), .B(A[769]), .Z(n2809) );
  AND U3069 ( .A(n2812), .B(n2813), .Z(n515) );
  NAND U3070 ( .A(B[768]), .B(n2814), .Z(n2813) );
  NANDN U3071 ( .A(A[768]), .B(n517), .Z(n2814) );
  NANDN U3072 ( .A(n517), .B(A[768]), .Z(n2812) );
  AND U3073 ( .A(n2815), .B(n2816), .Z(n517) );
  NAND U3074 ( .A(B[767]), .B(n2817), .Z(n2816) );
  NANDN U3075 ( .A(A[767]), .B(n519), .Z(n2817) );
  NANDN U3076 ( .A(n519), .B(A[767]), .Z(n2815) );
  AND U3077 ( .A(n2818), .B(n2819), .Z(n519) );
  NAND U3078 ( .A(B[766]), .B(n2820), .Z(n2819) );
  NANDN U3079 ( .A(A[766]), .B(n521), .Z(n2820) );
  NANDN U3080 ( .A(n521), .B(A[766]), .Z(n2818) );
  AND U3081 ( .A(n2821), .B(n2822), .Z(n521) );
  NAND U3082 ( .A(B[765]), .B(n2823), .Z(n2822) );
  NANDN U3083 ( .A(A[765]), .B(n523), .Z(n2823) );
  NANDN U3084 ( .A(n523), .B(A[765]), .Z(n2821) );
  AND U3085 ( .A(n2824), .B(n2825), .Z(n523) );
  NAND U3086 ( .A(B[764]), .B(n2826), .Z(n2825) );
  NANDN U3087 ( .A(A[764]), .B(n525), .Z(n2826) );
  NANDN U3088 ( .A(n525), .B(A[764]), .Z(n2824) );
  AND U3089 ( .A(n2827), .B(n2828), .Z(n525) );
  NAND U3090 ( .A(B[763]), .B(n2829), .Z(n2828) );
  NANDN U3091 ( .A(A[763]), .B(n527), .Z(n2829) );
  NANDN U3092 ( .A(n527), .B(A[763]), .Z(n2827) );
  AND U3093 ( .A(n2830), .B(n2831), .Z(n527) );
  NAND U3094 ( .A(B[762]), .B(n2832), .Z(n2831) );
  NANDN U3095 ( .A(A[762]), .B(n529), .Z(n2832) );
  NANDN U3096 ( .A(n529), .B(A[762]), .Z(n2830) );
  AND U3097 ( .A(n2833), .B(n2834), .Z(n529) );
  NAND U3098 ( .A(B[761]), .B(n2835), .Z(n2834) );
  NANDN U3099 ( .A(A[761]), .B(n531), .Z(n2835) );
  NANDN U3100 ( .A(n531), .B(A[761]), .Z(n2833) );
  AND U3101 ( .A(n2836), .B(n2837), .Z(n531) );
  NAND U3102 ( .A(B[760]), .B(n2838), .Z(n2837) );
  NANDN U3103 ( .A(A[760]), .B(n533), .Z(n2838) );
  NANDN U3104 ( .A(n533), .B(A[760]), .Z(n2836) );
  AND U3105 ( .A(n2839), .B(n2840), .Z(n533) );
  NAND U3106 ( .A(B[759]), .B(n2841), .Z(n2840) );
  NANDN U3107 ( .A(A[759]), .B(n537), .Z(n2841) );
  NANDN U3108 ( .A(n537), .B(A[759]), .Z(n2839) );
  AND U3109 ( .A(n2842), .B(n2843), .Z(n537) );
  NAND U3110 ( .A(B[758]), .B(n2844), .Z(n2843) );
  NANDN U3111 ( .A(A[758]), .B(n539), .Z(n2844) );
  NANDN U3112 ( .A(n539), .B(A[758]), .Z(n2842) );
  AND U3113 ( .A(n2845), .B(n2846), .Z(n539) );
  NAND U3114 ( .A(B[757]), .B(n2847), .Z(n2846) );
  NANDN U3115 ( .A(A[757]), .B(n541), .Z(n2847) );
  NANDN U3116 ( .A(n541), .B(A[757]), .Z(n2845) );
  AND U3117 ( .A(n2848), .B(n2849), .Z(n541) );
  NAND U3118 ( .A(B[756]), .B(n2850), .Z(n2849) );
  NANDN U3119 ( .A(A[756]), .B(n543), .Z(n2850) );
  NANDN U3120 ( .A(n543), .B(A[756]), .Z(n2848) );
  AND U3121 ( .A(n2851), .B(n2852), .Z(n543) );
  NAND U3122 ( .A(B[755]), .B(n2853), .Z(n2852) );
  NANDN U3123 ( .A(A[755]), .B(n545), .Z(n2853) );
  NANDN U3124 ( .A(n545), .B(A[755]), .Z(n2851) );
  AND U3125 ( .A(n2854), .B(n2855), .Z(n545) );
  NAND U3126 ( .A(B[754]), .B(n2856), .Z(n2855) );
  NANDN U3127 ( .A(A[754]), .B(n547), .Z(n2856) );
  NANDN U3128 ( .A(n547), .B(A[754]), .Z(n2854) );
  AND U3129 ( .A(n2857), .B(n2858), .Z(n547) );
  NAND U3130 ( .A(B[753]), .B(n2859), .Z(n2858) );
  NANDN U3131 ( .A(A[753]), .B(n549), .Z(n2859) );
  NANDN U3132 ( .A(n549), .B(A[753]), .Z(n2857) );
  AND U3133 ( .A(n2860), .B(n2861), .Z(n549) );
  NAND U3134 ( .A(B[752]), .B(n2862), .Z(n2861) );
  NANDN U3135 ( .A(A[752]), .B(n551), .Z(n2862) );
  NANDN U3136 ( .A(n551), .B(A[752]), .Z(n2860) );
  AND U3137 ( .A(n2863), .B(n2864), .Z(n551) );
  NAND U3138 ( .A(B[751]), .B(n2865), .Z(n2864) );
  NANDN U3139 ( .A(A[751]), .B(n553), .Z(n2865) );
  NANDN U3140 ( .A(n553), .B(A[751]), .Z(n2863) );
  AND U3141 ( .A(n2866), .B(n2867), .Z(n553) );
  NAND U3142 ( .A(B[750]), .B(n2868), .Z(n2867) );
  NANDN U3143 ( .A(A[750]), .B(n555), .Z(n2868) );
  NANDN U3144 ( .A(n555), .B(A[750]), .Z(n2866) );
  AND U3145 ( .A(n2869), .B(n2870), .Z(n555) );
  NAND U3146 ( .A(B[749]), .B(n2871), .Z(n2870) );
  NANDN U3147 ( .A(A[749]), .B(n559), .Z(n2871) );
  NANDN U3148 ( .A(n559), .B(A[749]), .Z(n2869) );
  AND U3149 ( .A(n2872), .B(n2873), .Z(n559) );
  NAND U3150 ( .A(B[748]), .B(n2874), .Z(n2873) );
  NANDN U3151 ( .A(A[748]), .B(n561), .Z(n2874) );
  NANDN U3152 ( .A(n561), .B(A[748]), .Z(n2872) );
  AND U3153 ( .A(n2875), .B(n2876), .Z(n561) );
  NAND U3154 ( .A(B[747]), .B(n2877), .Z(n2876) );
  NANDN U3155 ( .A(A[747]), .B(n563), .Z(n2877) );
  NANDN U3156 ( .A(n563), .B(A[747]), .Z(n2875) );
  AND U3157 ( .A(n2878), .B(n2879), .Z(n563) );
  NAND U3158 ( .A(B[746]), .B(n2880), .Z(n2879) );
  NANDN U3159 ( .A(A[746]), .B(n565), .Z(n2880) );
  NANDN U3160 ( .A(n565), .B(A[746]), .Z(n2878) );
  AND U3161 ( .A(n2881), .B(n2882), .Z(n565) );
  NAND U3162 ( .A(B[745]), .B(n2883), .Z(n2882) );
  NANDN U3163 ( .A(A[745]), .B(n567), .Z(n2883) );
  NANDN U3164 ( .A(n567), .B(A[745]), .Z(n2881) );
  AND U3165 ( .A(n2884), .B(n2885), .Z(n567) );
  NAND U3166 ( .A(B[744]), .B(n2886), .Z(n2885) );
  NANDN U3167 ( .A(A[744]), .B(n569), .Z(n2886) );
  NANDN U3168 ( .A(n569), .B(A[744]), .Z(n2884) );
  AND U3169 ( .A(n2887), .B(n2888), .Z(n569) );
  NAND U3170 ( .A(B[743]), .B(n2889), .Z(n2888) );
  NANDN U3171 ( .A(A[743]), .B(n571), .Z(n2889) );
  NANDN U3172 ( .A(n571), .B(A[743]), .Z(n2887) );
  AND U3173 ( .A(n2890), .B(n2891), .Z(n571) );
  NAND U3174 ( .A(B[742]), .B(n2892), .Z(n2891) );
  NANDN U3175 ( .A(A[742]), .B(n573), .Z(n2892) );
  NANDN U3176 ( .A(n573), .B(A[742]), .Z(n2890) );
  AND U3177 ( .A(n2893), .B(n2894), .Z(n573) );
  NAND U3178 ( .A(B[741]), .B(n2895), .Z(n2894) );
  NANDN U3179 ( .A(A[741]), .B(n575), .Z(n2895) );
  NANDN U3180 ( .A(n575), .B(A[741]), .Z(n2893) );
  AND U3181 ( .A(n2896), .B(n2897), .Z(n575) );
  NAND U3182 ( .A(B[740]), .B(n2898), .Z(n2897) );
  NANDN U3183 ( .A(A[740]), .B(n577), .Z(n2898) );
  NANDN U3184 ( .A(n577), .B(A[740]), .Z(n2896) );
  AND U3185 ( .A(n2899), .B(n2900), .Z(n577) );
  NAND U3186 ( .A(B[739]), .B(n2901), .Z(n2900) );
  NANDN U3187 ( .A(A[739]), .B(n581), .Z(n2901) );
  NANDN U3188 ( .A(n581), .B(A[739]), .Z(n2899) );
  AND U3189 ( .A(n2902), .B(n2903), .Z(n581) );
  NAND U3190 ( .A(B[738]), .B(n2904), .Z(n2903) );
  NANDN U3191 ( .A(A[738]), .B(n583), .Z(n2904) );
  NANDN U3192 ( .A(n583), .B(A[738]), .Z(n2902) );
  AND U3193 ( .A(n2905), .B(n2906), .Z(n583) );
  NAND U3194 ( .A(B[737]), .B(n2907), .Z(n2906) );
  NANDN U3195 ( .A(A[737]), .B(n585), .Z(n2907) );
  NANDN U3196 ( .A(n585), .B(A[737]), .Z(n2905) );
  AND U3197 ( .A(n2908), .B(n2909), .Z(n585) );
  NAND U3198 ( .A(B[736]), .B(n2910), .Z(n2909) );
  NANDN U3199 ( .A(A[736]), .B(n587), .Z(n2910) );
  NANDN U3200 ( .A(n587), .B(A[736]), .Z(n2908) );
  AND U3201 ( .A(n2911), .B(n2912), .Z(n587) );
  NAND U3202 ( .A(B[735]), .B(n2913), .Z(n2912) );
  NANDN U3203 ( .A(A[735]), .B(n589), .Z(n2913) );
  NANDN U3204 ( .A(n589), .B(A[735]), .Z(n2911) );
  AND U3205 ( .A(n2914), .B(n2915), .Z(n589) );
  NAND U3206 ( .A(B[734]), .B(n2916), .Z(n2915) );
  NANDN U3207 ( .A(A[734]), .B(n591), .Z(n2916) );
  NANDN U3208 ( .A(n591), .B(A[734]), .Z(n2914) );
  AND U3209 ( .A(n2917), .B(n2918), .Z(n591) );
  NAND U3210 ( .A(B[733]), .B(n2919), .Z(n2918) );
  NANDN U3211 ( .A(A[733]), .B(n593), .Z(n2919) );
  NANDN U3212 ( .A(n593), .B(A[733]), .Z(n2917) );
  AND U3213 ( .A(n2920), .B(n2921), .Z(n593) );
  NAND U3214 ( .A(B[732]), .B(n2922), .Z(n2921) );
  NANDN U3215 ( .A(A[732]), .B(n595), .Z(n2922) );
  NANDN U3216 ( .A(n595), .B(A[732]), .Z(n2920) );
  AND U3217 ( .A(n2923), .B(n2924), .Z(n595) );
  NAND U3218 ( .A(B[731]), .B(n2925), .Z(n2924) );
  NANDN U3219 ( .A(A[731]), .B(n597), .Z(n2925) );
  NANDN U3220 ( .A(n597), .B(A[731]), .Z(n2923) );
  AND U3221 ( .A(n2926), .B(n2927), .Z(n597) );
  NAND U3222 ( .A(B[730]), .B(n2928), .Z(n2927) );
  NANDN U3223 ( .A(A[730]), .B(n599), .Z(n2928) );
  NANDN U3224 ( .A(n599), .B(A[730]), .Z(n2926) );
  AND U3225 ( .A(n2929), .B(n2930), .Z(n599) );
  NAND U3226 ( .A(B[729]), .B(n2931), .Z(n2930) );
  NANDN U3227 ( .A(A[729]), .B(n603), .Z(n2931) );
  NANDN U3228 ( .A(n603), .B(A[729]), .Z(n2929) );
  AND U3229 ( .A(n2932), .B(n2933), .Z(n603) );
  NAND U3230 ( .A(B[728]), .B(n2934), .Z(n2933) );
  NANDN U3231 ( .A(A[728]), .B(n605), .Z(n2934) );
  NANDN U3232 ( .A(n605), .B(A[728]), .Z(n2932) );
  AND U3233 ( .A(n2935), .B(n2936), .Z(n605) );
  NAND U3234 ( .A(B[727]), .B(n2937), .Z(n2936) );
  NANDN U3235 ( .A(A[727]), .B(n607), .Z(n2937) );
  NANDN U3236 ( .A(n607), .B(A[727]), .Z(n2935) );
  AND U3237 ( .A(n2938), .B(n2939), .Z(n607) );
  NAND U3238 ( .A(B[726]), .B(n2940), .Z(n2939) );
  NANDN U3239 ( .A(A[726]), .B(n609), .Z(n2940) );
  NANDN U3240 ( .A(n609), .B(A[726]), .Z(n2938) );
  AND U3241 ( .A(n2941), .B(n2942), .Z(n609) );
  NAND U3242 ( .A(B[725]), .B(n2943), .Z(n2942) );
  NANDN U3243 ( .A(A[725]), .B(n611), .Z(n2943) );
  NANDN U3244 ( .A(n611), .B(A[725]), .Z(n2941) );
  AND U3245 ( .A(n2944), .B(n2945), .Z(n611) );
  NAND U3246 ( .A(B[724]), .B(n2946), .Z(n2945) );
  NANDN U3247 ( .A(A[724]), .B(n613), .Z(n2946) );
  NANDN U3248 ( .A(n613), .B(A[724]), .Z(n2944) );
  AND U3249 ( .A(n2947), .B(n2948), .Z(n613) );
  NAND U3250 ( .A(B[723]), .B(n2949), .Z(n2948) );
  NANDN U3251 ( .A(A[723]), .B(n615), .Z(n2949) );
  NANDN U3252 ( .A(n615), .B(A[723]), .Z(n2947) );
  AND U3253 ( .A(n2950), .B(n2951), .Z(n615) );
  NAND U3254 ( .A(B[722]), .B(n2952), .Z(n2951) );
  NANDN U3255 ( .A(A[722]), .B(n617), .Z(n2952) );
  NANDN U3256 ( .A(n617), .B(A[722]), .Z(n2950) );
  AND U3257 ( .A(n2953), .B(n2954), .Z(n617) );
  NAND U3258 ( .A(B[721]), .B(n2955), .Z(n2954) );
  NANDN U3259 ( .A(A[721]), .B(n619), .Z(n2955) );
  NANDN U3260 ( .A(n619), .B(A[721]), .Z(n2953) );
  AND U3261 ( .A(n2956), .B(n2957), .Z(n619) );
  NAND U3262 ( .A(B[720]), .B(n2958), .Z(n2957) );
  NANDN U3263 ( .A(A[720]), .B(n621), .Z(n2958) );
  NANDN U3264 ( .A(n621), .B(A[720]), .Z(n2956) );
  AND U3265 ( .A(n2959), .B(n2960), .Z(n621) );
  NAND U3266 ( .A(B[719]), .B(n2961), .Z(n2960) );
  NANDN U3267 ( .A(A[719]), .B(n625), .Z(n2961) );
  NANDN U3268 ( .A(n625), .B(A[719]), .Z(n2959) );
  AND U3269 ( .A(n2962), .B(n2963), .Z(n625) );
  NAND U3270 ( .A(B[718]), .B(n2964), .Z(n2963) );
  NANDN U3271 ( .A(A[718]), .B(n627), .Z(n2964) );
  NANDN U3272 ( .A(n627), .B(A[718]), .Z(n2962) );
  AND U3273 ( .A(n2965), .B(n2966), .Z(n627) );
  NAND U3274 ( .A(B[717]), .B(n2967), .Z(n2966) );
  NANDN U3275 ( .A(A[717]), .B(n629), .Z(n2967) );
  NANDN U3276 ( .A(n629), .B(A[717]), .Z(n2965) );
  AND U3277 ( .A(n2968), .B(n2969), .Z(n629) );
  NAND U3278 ( .A(B[716]), .B(n2970), .Z(n2969) );
  NANDN U3279 ( .A(A[716]), .B(n631), .Z(n2970) );
  NANDN U3280 ( .A(n631), .B(A[716]), .Z(n2968) );
  AND U3281 ( .A(n2971), .B(n2972), .Z(n631) );
  NAND U3282 ( .A(B[715]), .B(n2973), .Z(n2972) );
  NANDN U3283 ( .A(A[715]), .B(n633), .Z(n2973) );
  NANDN U3284 ( .A(n633), .B(A[715]), .Z(n2971) );
  AND U3285 ( .A(n2974), .B(n2975), .Z(n633) );
  NAND U3286 ( .A(B[714]), .B(n2976), .Z(n2975) );
  NANDN U3287 ( .A(A[714]), .B(n635), .Z(n2976) );
  NANDN U3288 ( .A(n635), .B(A[714]), .Z(n2974) );
  AND U3289 ( .A(n2977), .B(n2978), .Z(n635) );
  NAND U3290 ( .A(B[713]), .B(n2979), .Z(n2978) );
  NANDN U3291 ( .A(A[713]), .B(n637), .Z(n2979) );
  NANDN U3292 ( .A(n637), .B(A[713]), .Z(n2977) );
  AND U3293 ( .A(n2980), .B(n2981), .Z(n637) );
  NAND U3294 ( .A(B[712]), .B(n2982), .Z(n2981) );
  NANDN U3295 ( .A(A[712]), .B(n639), .Z(n2982) );
  NANDN U3296 ( .A(n639), .B(A[712]), .Z(n2980) );
  AND U3297 ( .A(n2983), .B(n2984), .Z(n639) );
  NAND U3298 ( .A(B[711]), .B(n2985), .Z(n2984) );
  NANDN U3299 ( .A(A[711]), .B(n641), .Z(n2985) );
  NANDN U3300 ( .A(n641), .B(A[711]), .Z(n2983) );
  AND U3301 ( .A(n2986), .B(n2987), .Z(n641) );
  NAND U3302 ( .A(B[710]), .B(n2988), .Z(n2987) );
  NANDN U3303 ( .A(A[710]), .B(n643), .Z(n2988) );
  NANDN U3304 ( .A(n643), .B(A[710]), .Z(n2986) );
  AND U3305 ( .A(n2989), .B(n2990), .Z(n643) );
  NAND U3306 ( .A(B[709]), .B(n2991), .Z(n2990) );
  NANDN U3307 ( .A(A[709]), .B(n647), .Z(n2991) );
  NANDN U3308 ( .A(n647), .B(A[709]), .Z(n2989) );
  AND U3309 ( .A(n2992), .B(n2993), .Z(n647) );
  NAND U3310 ( .A(B[708]), .B(n2994), .Z(n2993) );
  NANDN U3311 ( .A(A[708]), .B(n649), .Z(n2994) );
  NANDN U3312 ( .A(n649), .B(A[708]), .Z(n2992) );
  AND U3313 ( .A(n2995), .B(n2996), .Z(n649) );
  NAND U3314 ( .A(B[707]), .B(n2997), .Z(n2996) );
  NANDN U3315 ( .A(A[707]), .B(n651), .Z(n2997) );
  NANDN U3316 ( .A(n651), .B(A[707]), .Z(n2995) );
  AND U3317 ( .A(n2998), .B(n2999), .Z(n651) );
  NAND U3318 ( .A(B[706]), .B(n3000), .Z(n2999) );
  NANDN U3319 ( .A(A[706]), .B(n653), .Z(n3000) );
  NANDN U3320 ( .A(n653), .B(A[706]), .Z(n2998) );
  AND U3321 ( .A(n3001), .B(n3002), .Z(n653) );
  NAND U3322 ( .A(B[705]), .B(n3003), .Z(n3002) );
  NANDN U3323 ( .A(A[705]), .B(n655), .Z(n3003) );
  NANDN U3324 ( .A(n655), .B(A[705]), .Z(n3001) );
  AND U3325 ( .A(n3004), .B(n3005), .Z(n655) );
  NAND U3326 ( .A(B[704]), .B(n3006), .Z(n3005) );
  NANDN U3327 ( .A(A[704]), .B(n657), .Z(n3006) );
  NANDN U3328 ( .A(n657), .B(A[704]), .Z(n3004) );
  AND U3329 ( .A(n3007), .B(n3008), .Z(n657) );
  NAND U3330 ( .A(B[703]), .B(n3009), .Z(n3008) );
  NANDN U3331 ( .A(A[703]), .B(n659), .Z(n3009) );
  NANDN U3332 ( .A(n659), .B(A[703]), .Z(n3007) );
  AND U3333 ( .A(n3010), .B(n3011), .Z(n659) );
  NAND U3334 ( .A(B[702]), .B(n3012), .Z(n3011) );
  NANDN U3335 ( .A(A[702]), .B(n661), .Z(n3012) );
  NANDN U3336 ( .A(n661), .B(A[702]), .Z(n3010) );
  AND U3337 ( .A(n3013), .B(n3014), .Z(n661) );
  NAND U3338 ( .A(B[701]), .B(n3015), .Z(n3014) );
  NANDN U3339 ( .A(A[701]), .B(n663), .Z(n3015) );
  NANDN U3340 ( .A(n663), .B(A[701]), .Z(n3013) );
  AND U3341 ( .A(n3016), .B(n3017), .Z(n663) );
  NAND U3342 ( .A(B[700]), .B(n3018), .Z(n3017) );
  NANDN U3343 ( .A(A[700]), .B(n665), .Z(n3018) );
  NANDN U3344 ( .A(n665), .B(A[700]), .Z(n3016) );
  AND U3345 ( .A(n3019), .B(n3020), .Z(n665) );
  NAND U3346 ( .A(B[699]), .B(n3021), .Z(n3020) );
  NANDN U3347 ( .A(A[699]), .B(n671), .Z(n3021) );
  NANDN U3348 ( .A(n671), .B(A[699]), .Z(n3019) );
  AND U3349 ( .A(n3022), .B(n3023), .Z(n671) );
  NAND U3350 ( .A(B[698]), .B(n3024), .Z(n3023) );
  NANDN U3351 ( .A(A[698]), .B(n673), .Z(n3024) );
  NANDN U3352 ( .A(n673), .B(A[698]), .Z(n3022) );
  AND U3353 ( .A(n3025), .B(n3026), .Z(n673) );
  NAND U3354 ( .A(B[697]), .B(n3027), .Z(n3026) );
  NANDN U3355 ( .A(A[697]), .B(n675), .Z(n3027) );
  NANDN U3356 ( .A(n675), .B(A[697]), .Z(n3025) );
  AND U3357 ( .A(n3028), .B(n3029), .Z(n675) );
  NAND U3358 ( .A(B[696]), .B(n3030), .Z(n3029) );
  NANDN U3359 ( .A(A[696]), .B(n677), .Z(n3030) );
  NANDN U3360 ( .A(n677), .B(A[696]), .Z(n3028) );
  AND U3361 ( .A(n3031), .B(n3032), .Z(n677) );
  NAND U3362 ( .A(B[695]), .B(n3033), .Z(n3032) );
  NANDN U3363 ( .A(A[695]), .B(n679), .Z(n3033) );
  NANDN U3364 ( .A(n679), .B(A[695]), .Z(n3031) );
  AND U3365 ( .A(n3034), .B(n3035), .Z(n679) );
  NAND U3366 ( .A(B[694]), .B(n3036), .Z(n3035) );
  NANDN U3367 ( .A(A[694]), .B(n681), .Z(n3036) );
  NANDN U3368 ( .A(n681), .B(A[694]), .Z(n3034) );
  AND U3369 ( .A(n3037), .B(n3038), .Z(n681) );
  NAND U3370 ( .A(B[693]), .B(n3039), .Z(n3038) );
  NANDN U3371 ( .A(A[693]), .B(n683), .Z(n3039) );
  NANDN U3372 ( .A(n683), .B(A[693]), .Z(n3037) );
  AND U3373 ( .A(n3040), .B(n3041), .Z(n683) );
  NAND U3374 ( .A(B[692]), .B(n3042), .Z(n3041) );
  NANDN U3375 ( .A(A[692]), .B(n685), .Z(n3042) );
  NANDN U3376 ( .A(n685), .B(A[692]), .Z(n3040) );
  AND U3377 ( .A(n3043), .B(n3044), .Z(n685) );
  NAND U3378 ( .A(B[691]), .B(n3045), .Z(n3044) );
  NANDN U3379 ( .A(A[691]), .B(n687), .Z(n3045) );
  NANDN U3380 ( .A(n687), .B(A[691]), .Z(n3043) );
  AND U3381 ( .A(n3046), .B(n3047), .Z(n687) );
  NAND U3382 ( .A(B[690]), .B(n3048), .Z(n3047) );
  NANDN U3383 ( .A(A[690]), .B(n689), .Z(n3048) );
  NANDN U3384 ( .A(n689), .B(A[690]), .Z(n3046) );
  AND U3385 ( .A(n3049), .B(n3050), .Z(n689) );
  NAND U3386 ( .A(B[689]), .B(n3051), .Z(n3050) );
  NANDN U3387 ( .A(A[689]), .B(n693), .Z(n3051) );
  NANDN U3388 ( .A(n693), .B(A[689]), .Z(n3049) );
  AND U3389 ( .A(n3052), .B(n3053), .Z(n693) );
  NAND U3390 ( .A(B[688]), .B(n3054), .Z(n3053) );
  NANDN U3391 ( .A(A[688]), .B(n695), .Z(n3054) );
  NANDN U3392 ( .A(n695), .B(A[688]), .Z(n3052) );
  AND U3393 ( .A(n3055), .B(n3056), .Z(n695) );
  NAND U3394 ( .A(B[687]), .B(n3057), .Z(n3056) );
  NANDN U3395 ( .A(A[687]), .B(n697), .Z(n3057) );
  NANDN U3396 ( .A(n697), .B(A[687]), .Z(n3055) );
  AND U3397 ( .A(n3058), .B(n3059), .Z(n697) );
  NAND U3398 ( .A(B[686]), .B(n3060), .Z(n3059) );
  NANDN U3399 ( .A(A[686]), .B(n699), .Z(n3060) );
  NANDN U3400 ( .A(n699), .B(A[686]), .Z(n3058) );
  AND U3401 ( .A(n3061), .B(n3062), .Z(n699) );
  NAND U3402 ( .A(B[685]), .B(n3063), .Z(n3062) );
  NANDN U3403 ( .A(A[685]), .B(n701), .Z(n3063) );
  NANDN U3404 ( .A(n701), .B(A[685]), .Z(n3061) );
  AND U3405 ( .A(n3064), .B(n3065), .Z(n701) );
  NAND U3406 ( .A(B[684]), .B(n3066), .Z(n3065) );
  NANDN U3407 ( .A(A[684]), .B(n703), .Z(n3066) );
  NANDN U3408 ( .A(n703), .B(A[684]), .Z(n3064) );
  AND U3409 ( .A(n3067), .B(n3068), .Z(n703) );
  NAND U3410 ( .A(B[683]), .B(n3069), .Z(n3068) );
  NANDN U3411 ( .A(A[683]), .B(n705), .Z(n3069) );
  NANDN U3412 ( .A(n705), .B(A[683]), .Z(n3067) );
  AND U3413 ( .A(n3070), .B(n3071), .Z(n705) );
  NAND U3414 ( .A(B[682]), .B(n3072), .Z(n3071) );
  NANDN U3415 ( .A(A[682]), .B(n707), .Z(n3072) );
  NANDN U3416 ( .A(n707), .B(A[682]), .Z(n3070) );
  AND U3417 ( .A(n3073), .B(n3074), .Z(n707) );
  NAND U3418 ( .A(B[681]), .B(n3075), .Z(n3074) );
  NANDN U3419 ( .A(A[681]), .B(n709), .Z(n3075) );
  NANDN U3420 ( .A(n709), .B(A[681]), .Z(n3073) );
  AND U3421 ( .A(n3076), .B(n3077), .Z(n709) );
  NAND U3422 ( .A(B[680]), .B(n3078), .Z(n3077) );
  NANDN U3423 ( .A(A[680]), .B(n711), .Z(n3078) );
  NANDN U3424 ( .A(n711), .B(A[680]), .Z(n3076) );
  AND U3425 ( .A(n3079), .B(n3080), .Z(n711) );
  NAND U3426 ( .A(B[679]), .B(n3081), .Z(n3080) );
  NANDN U3427 ( .A(A[679]), .B(n715), .Z(n3081) );
  NANDN U3428 ( .A(n715), .B(A[679]), .Z(n3079) );
  AND U3429 ( .A(n3082), .B(n3083), .Z(n715) );
  NAND U3430 ( .A(B[678]), .B(n3084), .Z(n3083) );
  NANDN U3431 ( .A(A[678]), .B(n717), .Z(n3084) );
  NANDN U3432 ( .A(n717), .B(A[678]), .Z(n3082) );
  AND U3433 ( .A(n3085), .B(n3086), .Z(n717) );
  NAND U3434 ( .A(B[677]), .B(n3087), .Z(n3086) );
  NANDN U3435 ( .A(A[677]), .B(n719), .Z(n3087) );
  NANDN U3436 ( .A(n719), .B(A[677]), .Z(n3085) );
  AND U3437 ( .A(n3088), .B(n3089), .Z(n719) );
  NAND U3438 ( .A(B[676]), .B(n3090), .Z(n3089) );
  NANDN U3439 ( .A(A[676]), .B(n721), .Z(n3090) );
  NANDN U3440 ( .A(n721), .B(A[676]), .Z(n3088) );
  AND U3441 ( .A(n3091), .B(n3092), .Z(n721) );
  NAND U3442 ( .A(B[675]), .B(n3093), .Z(n3092) );
  NANDN U3443 ( .A(A[675]), .B(n723), .Z(n3093) );
  NANDN U3444 ( .A(n723), .B(A[675]), .Z(n3091) );
  AND U3445 ( .A(n3094), .B(n3095), .Z(n723) );
  NAND U3446 ( .A(B[674]), .B(n3096), .Z(n3095) );
  NANDN U3447 ( .A(A[674]), .B(n725), .Z(n3096) );
  NANDN U3448 ( .A(n725), .B(A[674]), .Z(n3094) );
  AND U3449 ( .A(n3097), .B(n3098), .Z(n725) );
  NAND U3450 ( .A(B[673]), .B(n3099), .Z(n3098) );
  NANDN U3451 ( .A(A[673]), .B(n727), .Z(n3099) );
  NANDN U3452 ( .A(n727), .B(A[673]), .Z(n3097) );
  AND U3453 ( .A(n3100), .B(n3101), .Z(n727) );
  NAND U3454 ( .A(B[672]), .B(n3102), .Z(n3101) );
  NANDN U3455 ( .A(A[672]), .B(n729), .Z(n3102) );
  NANDN U3456 ( .A(n729), .B(A[672]), .Z(n3100) );
  AND U3457 ( .A(n3103), .B(n3104), .Z(n729) );
  NAND U3458 ( .A(B[671]), .B(n3105), .Z(n3104) );
  NANDN U3459 ( .A(A[671]), .B(n731), .Z(n3105) );
  NANDN U3460 ( .A(n731), .B(A[671]), .Z(n3103) );
  AND U3461 ( .A(n3106), .B(n3107), .Z(n731) );
  NAND U3462 ( .A(B[670]), .B(n3108), .Z(n3107) );
  NANDN U3463 ( .A(A[670]), .B(n733), .Z(n3108) );
  NANDN U3464 ( .A(n733), .B(A[670]), .Z(n3106) );
  AND U3465 ( .A(n3109), .B(n3110), .Z(n733) );
  NAND U3466 ( .A(B[669]), .B(n3111), .Z(n3110) );
  NANDN U3467 ( .A(A[669]), .B(n737), .Z(n3111) );
  NANDN U3468 ( .A(n737), .B(A[669]), .Z(n3109) );
  AND U3469 ( .A(n3112), .B(n3113), .Z(n737) );
  NAND U3470 ( .A(B[668]), .B(n3114), .Z(n3113) );
  NANDN U3471 ( .A(A[668]), .B(n739), .Z(n3114) );
  NANDN U3472 ( .A(n739), .B(A[668]), .Z(n3112) );
  AND U3473 ( .A(n3115), .B(n3116), .Z(n739) );
  NAND U3474 ( .A(B[667]), .B(n3117), .Z(n3116) );
  NANDN U3475 ( .A(A[667]), .B(n741), .Z(n3117) );
  NANDN U3476 ( .A(n741), .B(A[667]), .Z(n3115) );
  AND U3477 ( .A(n3118), .B(n3119), .Z(n741) );
  NAND U3478 ( .A(B[666]), .B(n3120), .Z(n3119) );
  NANDN U3479 ( .A(A[666]), .B(n743), .Z(n3120) );
  NANDN U3480 ( .A(n743), .B(A[666]), .Z(n3118) );
  AND U3481 ( .A(n3121), .B(n3122), .Z(n743) );
  NAND U3482 ( .A(B[665]), .B(n3123), .Z(n3122) );
  NANDN U3483 ( .A(A[665]), .B(n745), .Z(n3123) );
  NANDN U3484 ( .A(n745), .B(A[665]), .Z(n3121) );
  AND U3485 ( .A(n3124), .B(n3125), .Z(n745) );
  NAND U3486 ( .A(B[664]), .B(n3126), .Z(n3125) );
  NANDN U3487 ( .A(A[664]), .B(n747), .Z(n3126) );
  NANDN U3488 ( .A(n747), .B(A[664]), .Z(n3124) );
  AND U3489 ( .A(n3127), .B(n3128), .Z(n747) );
  NAND U3490 ( .A(B[663]), .B(n3129), .Z(n3128) );
  NANDN U3491 ( .A(A[663]), .B(n749), .Z(n3129) );
  NANDN U3492 ( .A(n749), .B(A[663]), .Z(n3127) );
  AND U3493 ( .A(n3130), .B(n3131), .Z(n749) );
  NAND U3494 ( .A(B[662]), .B(n3132), .Z(n3131) );
  NANDN U3495 ( .A(A[662]), .B(n751), .Z(n3132) );
  NANDN U3496 ( .A(n751), .B(A[662]), .Z(n3130) );
  AND U3497 ( .A(n3133), .B(n3134), .Z(n751) );
  NAND U3498 ( .A(B[661]), .B(n3135), .Z(n3134) );
  NANDN U3499 ( .A(A[661]), .B(n753), .Z(n3135) );
  NANDN U3500 ( .A(n753), .B(A[661]), .Z(n3133) );
  AND U3501 ( .A(n3136), .B(n3137), .Z(n753) );
  NAND U3502 ( .A(B[660]), .B(n3138), .Z(n3137) );
  NANDN U3503 ( .A(A[660]), .B(n755), .Z(n3138) );
  NANDN U3504 ( .A(n755), .B(A[660]), .Z(n3136) );
  AND U3505 ( .A(n3139), .B(n3140), .Z(n755) );
  NAND U3506 ( .A(B[659]), .B(n3141), .Z(n3140) );
  NANDN U3507 ( .A(A[659]), .B(n759), .Z(n3141) );
  NANDN U3508 ( .A(n759), .B(A[659]), .Z(n3139) );
  AND U3509 ( .A(n3142), .B(n3143), .Z(n759) );
  NAND U3510 ( .A(B[658]), .B(n3144), .Z(n3143) );
  NANDN U3511 ( .A(A[658]), .B(n761), .Z(n3144) );
  NANDN U3512 ( .A(n761), .B(A[658]), .Z(n3142) );
  AND U3513 ( .A(n3145), .B(n3146), .Z(n761) );
  NAND U3514 ( .A(B[657]), .B(n3147), .Z(n3146) );
  NANDN U3515 ( .A(A[657]), .B(n763), .Z(n3147) );
  NANDN U3516 ( .A(n763), .B(A[657]), .Z(n3145) );
  AND U3517 ( .A(n3148), .B(n3149), .Z(n763) );
  NAND U3518 ( .A(B[656]), .B(n3150), .Z(n3149) );
  NANDN U3519 ( .A(A[656]), .B(n765), .Z(n3150) );
  NANDN U3520 ( .A(n765), .B(A[656]), .Z(n3148) );
  AND U3521 ( .A(n3151), .B(n3152), .Z(n765) );
  NAND U3522 ( .A(B[655]), .B(n3153), .Z(n3152) );
  NANDN U3523 ( .A(A[655]), .B(n767), .Z(n3153) );
  NANDN U3524 ( .A(n767), .B(A[655]), .Z(n3151) );
  AND U3525 ( .A(n3154), .B(n3155), .Z(n767) );
  NAND U3526 ( .A(B[654]), .B(n3156), .Z(n3155) );
  NANDN U3527 ( .A(A[654]), .B(n769), .Z(n3156) );
  NANDN U3528 ( .A(n769), .B(A[654]), .Z(n3154) );
  AND U3529 ( .A(n3157), .B(n3158), .Z(n769) );
  NAND U3530 ( .A(B[653]), .B(n3159), .Z(n3158) );
  NANDN U3531 ( .A(A[653]), .B(n771), .Z(n3159) );
  NANDN U3532 ( .A(n771), .B(A[653]), .Z(n3157) );
  AND U3533 ( .A(n3160), .B(n3161), .Z(n771) );
  NAND U3534 ( .A(B[652]), .B(n3162), .Z(n3161) );
  NANDN U3535 ( .A(A[652]), .B(n773), .Z(n3162) );
  NANDN U3536 ( .A(n773), .B(A[652]), .Z(n3160) );
  AND U3537 ( .A(n3163), .B(n3164), .Z(n773) );
  NAND U3538 ( .A(B[651]), .B(n3165), .Z(n3164) );
  NANDN U3539 ( .A(A[651]), .B(n775), .Z(n3165) );
  NANDN U3540 ( .A(n775), .B(A[651]), .Z(n3163) );
  AND U3541 ( .A(n3166), .B(n3167), .Z(n775) );
  NAND U3542 ( .A(B[650]), .B(n3168), .Z(n3167) );
  NANDN U3543 ( .A(A[650]), .B(n777), .Z(n3168) );
  NANDN U3544 ( .A(n777), .B(A[650]), .Z(n3166) );
  AND U3545 ( .A(n3169), .B(n3170), .Z(n777) );
  NAND U3546 ( .A(B[649]), .B(n3171), .Z(n3170) );
  NANDN U3547 ( .A(A[649]), .B(n781), .Z(n3171) );
  NANDN U3548 ( .A(n781), .B(A[649]), .Z(n3169) );
  AND U3549 ( .A(n3172), .B(n3173), .Z(n781) );
  NAND U3550 ( .A(B[648]), .B(n3174), .Z(n3173) );
  NANDN U3551 ( .A(A[648]), .B(n783), .Z(n3174) );
  NANDN U3552 ( .A(n783), .B(A[648]), .Z(n3172) );
  AND U3553 ( .A(n3175), .B(n3176), .Z(n783) );
  NAND U3554 ( .A(B[647]), .B(n3177), .Z(n3176) );
  NANDN U3555 ( .A(A[647]), .B(n785), .Z(n3177) );
  NANDN U3556 ( .A(n785), .B(A[647]), .Z(n3175) );
  AND U3557 ( .A(n3178), .B(n3179), .Z(n785) );
  NAND U3558 ( .A(B[646]), .B(n3180), .Z(n3179) );
  NANDN U3559 ( .A(A[646]), .B(n787), .Z(n3180) );
  NANDN U3560 ( .A(n787), .B(A[646]), .Z(n3178) );
  AND U3561 ( .A(n3181), .B(n3182), .Z(n787) );
  NAND U3562 ( .A(B[645]), .B(n3183), .Z(n3182) );
  NANDN U3563 ( .A(A[645]), .B(n789), .Z(n3183) );
  NANDN U3564 ( .A(n789), .B(A[645]), .Z(n3181) );
  AND U3565 ( .A(n3184), .B(n3185), .Z(n789) );
  NAND U3566 ( .A(B[644]), .B(n3186), .Z(n3185) );
  NANDN U3567 ( .A(A[644]), .B(n791), .Z(n3186) );
  NANDN U3568 ( .A(n791), .B(A[644]), .Z(n3184) );
  AND U3569 ( .A(n3187), .B(n3188), .Z(n791) );
  NAND U3570 ( .A(B[643]), .B(n3189), .Z(n3188) );
  NANDN U3571 ( .A(A[643]), .B(n793), .Z(n3189) );
  NANDN U3572 ( .A(n793), .B(A[643]), .Z(n3187) );
  AND U3573 ( .A(n3190), .B(n3191), .Z(n793) );
  NAND U3574 ( .A(B[642]), .B(n3192), .Z(n3191) );
  NANDN U3575 ( .A(A[642]), .B(n795), .Z(n3192) );
  NANDN U3576 ( .A(n795), .B(A[642]), .Z(n3190) );
  AND U3577 ( .A(n3193), .B(n3194), .Z(n795) );
  NAND U3578 ( .A(B[641]), .B(n3195), .Z(n3194) );
  NANDN U3579 ( .A(A[641]), .B(n797), .Z(n3195) );
  NANDN U3580 ( .A(n797), .B(A[641]), .Z(n3193) );
  AND U3581 ( .A(n3196), .B(n3197), .Z(n797) );
  NAND U3582 ( .A(B[640]), .B(n3198), .Z(n3197) );
  NANDN U3583 ( .A(A[640]), .B(n799), .Z(n3198) );
  NANDN U3584 ( .A(n799), .B(A[640]), .Z(n3196) );
  AND U3585 ( .A(n3199), .B(n3200), .Z(n799) );
  NAND U3586 ( .A(B[639]), .B(n3201), .Z(n3200) );
  NANDN U3587 ( .A(A[639]), .B(n803), .Z(n3201) );
  NANDN U3588 ( .A(n803), .B(A[639]), .Z(n3199) );
  AND U3589 ( .A(n3202), .B(n3203), .Z(n803) );
  NAND U3590 ( .A(B[638]), .B(n3204), .Z(n3203) );
  NANDN U3591 ( .A(A[638]), .B(n805), .Z(n3204) );
  NANDN U3592 ( .A(n805), .B(A[638]), .Z(n3202) );
  AND U3593 ( .A(n3205), .B(n3206), .Z(n805) );
  NAND U3594 ( .A(B[637]), .B(n3207), .Z(n3206) );
  NANDN U3595 ( .A(A[637]), .B(n807), .Z(n3207) );
  NANDN U3596 ( .A(n807), .B(A[637]), .Z(n3205) );
  AND U3597 ( .A(n3208), .B(n3209), .Z(n807) );
  NAND U3598 ( .A(B[636]), .B(n3210), .Z(n3209) );
  NANDN U3599 ( .A(A[636]), .B(n809), .Z(n3210) );
  NANDN U3600 ( .A(n809), .B(A[636]), .Z(n3208) );
  AND U3601 ( .A(n3211), .B(n3212), .Z(n809) );
  NAND U3602 ( .A(B[635]), .B(n3213), .Z(n3212) );
  NANDN U3603 ( .A(A[635]), .B(n811), .Z(n3213) );
  NANDN U3604 ( .A(n811), .B(A[635]), .Z(n3211) );
  AND U3605 ( .A(n3214), .B(n3215), .Z(n811) );
  NAND U3606 ( .A(B[634]), .B(n3216), .Z(n3215) );
  NANDN U3607 ( .A(A[634]), .B(n813), .Z(n3216) );
  NANDN U3608 ( .A(n813), .B(A[634]), .Z(n3214) );
  AND U3609 ( .A(n3217), .B(n3218), .Z(n813) );
  NAND U3610 ( .A(B[633]), .B(n3219), .Z(n3218) );
  NANDN U3611 ( .A(A[633]), .B(n815), .Z(n3219) );
  NANDN U3612 ( .A(n815), .B(A[633]), .Z(n3217) );
  AND U3613 ( .A(n3220), .B(n3221), .Z(n815) );
  NAND U3614 ( .A(B[632]), .B(n3222), .Z(n3221) );
  NANDN U3615 ( .A(A[632]), .B(n817), .Z(n3222) );
  NANDN U3616 ( .A(n817), .B(A[632]), .Z(n3220) );
  AND U3617 ( .A(n3223), .B(n3224), .Z(n817) );
  NAND U3618 ( .A(B[631]), .B(n3225), .Z(n3224) );
  NANDN U3619 ( .A(A[631]), .B(n819), .Z(n3225) );
  NANDN U3620 ( .A(n819), .B(A[631]), .Z(n3223) );
  AND U3621 ( .A(n3226), .B(n3227), .Z(n819) );
  NAND U3622 ( .A(B[630]), .B(n3228), .Z(n3227) );
  NANDN U3623 ( .A(A[630]), .B(n821), .Z(n3228) );
  NANDN U3624 ( .A(n821), .B(A[630]), .Z(n3226) );
  AND U3625 ( .A(n3229), .B(n3230), .Z(n821) );
  NAND U3626 ( .A(B[629]), .B(n3231), .Z(n3230) );
  NANDN U3627 ( .A(A[629]), .B(n825), .Z(n3231) );
  NANDN U3628 ( .A(n825), .B(A[629]), .Z(n3229) );
  AND U3629 ( .A(n3232), .B(n3233), .Z(n825) );
  NAND U3630 ( .A(B[628]), .B(n3234), .Z(n3233) );
  NANDN U3631 ( .A(A[628]), .B(n827), .Z(n3234) );
  NANDN U3632 ( .A(n827), .B(A[628]), .Z(n3232) );
  AND U3633 ( .A(n3235), .B(n3236), .Z(n827) );
  NAND U3634 ( .A(B[627]), .B(n3237), .Z(n3236) );
  NANDN U3635 ( .A(A[627]), .B(n829), .Z(n3237) );
  NANDN U3636 ( .A(n829), .B(A[627]), .Z(n3235) );
  AND U3637 ( .A(n3238), .B(n3239), .Z(n829) );
  NAND U3638 ( .A(B[626]), .B(n3240), .Z(n3239) );
  NANDN U3639 ( .A(A[626]), .B(n831), .Z(n3240) );
  NANDN U3640 ( .A(n831), .B(A[626]), .Z(n3238) );
  AND U3641 ( .A(n3241), .B(n3242), .Z(n831) );
  NAND U3642 ( .A(B[625]), .B(n3243), .Z(n3242) );
  NANDN U3643 ( .A(A[625]), .B(n833), .Z(n3243) );
  NANDN U3644 ( .A(n833), .B(A[625]), .Z(n3241) );
  AND U3645 ( .A(n3244), .B(n3245), .Z(n833) );
  NAND U3646 ( .A(B[624]), .B(n3246), .Z(n3245) );
  NANDN U3647 ( .A(A[624]), .B(n835), .Z(n3246) );
  NANDN U3648 ( .A(n835), .B(A[624]), .Z(n3244) );
  AND U3649 ( .A(n3247), .B(n3248), .Z(n835) );
  NAND U3650 ( .A(B[623]), .B(n3249), .Z(n3248) );
  NANDN U3651 ( .A(A[623]), .B(n837), .Z(n3249) );
  NANDN U3652 ( .A(n837), .B(A[623]), .Z(n3247) );
  AND U3653 ( .A(n3250), .B(n3251), .Z(n837) );
  NAND U3654 ( .A(B[622]), .B(n3252), .Z(n3251) );
  NANDN U3655 ( .A(A[622]), .B(n839), .Z(n3252) );
  NANDN U3656 ( .A(n839), .B(A[622]), .Z(n3250) );
  AND U3657 ( .A(n3253), .B(n3254), .Z(n839) );
  NAND U3658 ( .A(B[621]), .B(n3255), .Z(n3254) );
  NANDN U3659 ( .A(A[621]), .B(n841), .Z(n3255) );
  NANDN U3660 ( .A(n841), .B(A[621]), .Z(n3253) );
  AND U3661 ( .A(n3256), .B(n3257), .Z(n841) );
  NAND U3662 ( .A(B[620]), .B(n3258), .Z(n3257) );
  NANDN U3663 ( .A(A[620]), .B(n843), .Z(n3258) );
  NANDN U3664 ( .A(n843), .B(A[620]), .Z(n3256) );
  AND U3665 ( .A(n3259), .B(n3260), .Z(n843) );
  NAND U3666 ( .A(B[619]), .B(n3261), .Z(n3260) );
  NANDN U3667 ( .A(A[619]), .B(n847), .Z(n3261) );
  NANDN U3668 ( .A(n847), .B(A[619]), .Z(n3259) );
  AND U3669 ( .A(n3262), .B(n3263), .Z(n847) );
  NAND U3670 ( .A(B[618]), .B(n3264), .Z(n3263) );
  NANDN U3671 ( .A(A[618]), .B(n849), .Z(n3264) );
  NANDN U3672 ( .A(n849), .B(A[618]), .Z(n3262) );
  AND U3673 ( .A(n3265), .B(n3266), .Z(n849) );
  NAND U3674 ( .A(B[617]), .B(n3267), .Z(n3266) );
  NANDN U3675 ( .A(A[617]), .B(n851), .Z(n3267) );
  NANDN U3676 ( .A(n851), .B(A[617]), .Z(n3265) );
  AND U3677 ( .A(n3268), .B(n3269), .Z(n851) );
  NAND U3678 ( .A(B[616]), .B(n3270), .Z(n3269) );
  NANDN U3679 ( .A(A[616]), .B(n853), .Z(n3270) );
  NANDN U3680 ( .A(n853), .B(A[616]), .Z(n3268) );
  AND U3681 ( .A(n3271), .B(n3272), .Z(n853) );
  NAND U3682 ( .A(B[615]), .B(n3273), .Z(n3272) );
  NANDN U3683 ( .A(A[615]), .B(n855), .Z(n3273) );
  NANDN U3684 ( .A(n855), .B(A[615]), .Z(n3271) );
  AND U3685 ( .A(n3274), .B(n3275), .Z(n855) );
  NAND U3686 ( .A(B[614]), .B(n3276), .Z(n3275) );
  NANDN U3687 ( .A(A[614]), .B(n857), .Z(n3276) );
  NANDN U3688 ( .A(n857), .B(A[614]), .Z(n3274) );
  AND U3689 ( .A(n3277), .B(n3278), .Z(n857) );
  NAND U3690 ( .A(B[613]), .B(n3279), .Z(n3278) );
  NANDN U3691 ( .A(A[613]), .B(n859), .Z(n3279) );
  NANDN U3692 ( .A(n859), .B(A[613]), .Z(n3277) );
  AND U3693 ( .A(n3280), .B(n3281), .Z(n859) );
  NAND U3694 ( .A(B[612]), .B(n3282), .Z(n3281) );
  NANDN U3695 ( .A(A[612]), .B(n861), .Z(n3282) );
  NANDN U3696 ( .A(n861), .B(A[612]), .Z(n3280) );
  AND U3697 ( .A(n3283), .B(n3284), .Z(n861) );
  NAND U3698 ( .A(B[611]), .B(n3285), .Z(n3284) );
  NANDN U3699 ( .A(A[611]), .B(n863), .Z(n3285) );
  NANDN U3700 ( .A(n863), .B(A[611]), .Z(n3283) );
  AND U3701 ( .A(n3286), .B(n3287), .Z(n863) );
  NAND U3702 ( .A(B[610]), .B(n3288), .Z(n3287) );
  NANDN U3703 ( .A(A[610]), .B(n865), .Z(n3288) );
  NANDN U3704 ( .A(n865), .B(A[610]), .Z(n3286) );
  AND U3705 ( .A(n3289), .B(n3290), .Z(n865) );
  NAND U3706 ( .A(B[609]), .B(n3291), .Z(n3290) );
  NANDN U3707 ( .A(A[609]), .B(n869), .Z(n3291) );
  NANDN U3708 ( .A(n869), .B(A[609]), .Z(n3289) );
  AND U3709 ( .A(n3292), .B(n3293), .Z(n869) );
  NAND U3710 ( .A(B[608]), .B(n3294), .Z(n3293) );
  NANDN U3711 ( .A(A[608]), .B(n871), .Z(n3294) );
  NANDN U3712 ( .A(n871), .B(A[608]), .Z(n3292) );
  AND U3713 ( .A(n3295), .B(n3296), .Z(n871) );
  NAND U3714 ( .A(B[607]), .B(n3297), .Z(n3296) );
  NANDN U3715 ( .A(A[607]), .B(n873), .Z(n3297) );
  NANDN U3716 ( .A(n873), .B(A[607]), .Z(n3295) );
  AND U3717 ( .A(n3298), .B(n3299), .Z(n873) );
  NAND U3718 ( .A(B[606]), .B(n3300), .Z(n3299) );
  NANDN U3719 ( .A(A[606]), .B(n875), .Z(n3300) );
  NANDN U3720 ( .A(n875), .B(A[606]), .Z(n3298) );
  AND U3721 ( .A(n3301), .B(n3302), .Z(n875) );
  NAND U3722 ( .A(B[605]), .B(n3303), .Z(n3302) );
  NANDN U3723 ( .A(A[605]), .B(n877), .Z(n3303) );
  NANDN U3724 ( .A(n877), .B(A[605]), .Z(n3301) );
  AND U3725 ( .A(n3304), .B(n3305), .Z(n877) );
  NAND U3726 ( .A(B[604]), .B(n3306), .Z(n3305) );
  NANDN U3727 ( .A(A[604]), .B(n879), .Z(n3306) );
  NANDN U3728 ( .A(n879), .B(A[604]), .Z(n3304) );
  AND U3729 ( .A(n3307), .B(n3308), .Z(n879) );
  NAND U3730 ( .A(B[603]), .B(n3309), .Z(n3308) );
  NANDN U3731 ( .A(A[603]), .B(n881), .Z(n3309) );
  NANDN U3732 ( .A(n881), .B(A[603]), .Z(n3307) );
  AND U3733 ( .A(n3310), .B(n3311), .Z(n881) );
  NAND U3734 ( .A(B[602]), .B(n3312), .Z(n3311) );
  NANDN U3735 ( .A(A[602]), .B(n883), .Z(n3312) );
  NANDN U3736 ( .A(n883), .B(A[602]), .Z(n3310) );
  AND U3737 ( .A(n3313), .B(n3314), .Z(n883) );
  NAND U3738 ( .A(B[601]), .B(n3315), .Z(n3314) );
  NANDN U3739 ( .A(A[601]), .B(n885), .Z(n3315) );
  NANDN U3740 ( .A(n885), .B(A[601]), .Z(n3313) );
  AND U3741 ( .A(n3316), .B(n3317), .Z(n885) );
  NAND U3742 ( .A(B[600]), .B(n3318), .Z(n3317) );
  NANDN U3743 ( .A(A[600]), .B(n887), .Z(n3318) );
  NANDN U3744 ( .A(n887), .B(A[600]), .Z(n3316) );
  AND U3745 ( .A(n3319), .B(n3320), .Z(n887) );
  NAND U3746 ( .A(B[599]), .B(n3321), .Z(n3320) );
  NANDN U3747 ( .A(A[599]), .B(n893), .Z(n3321) );
  NANDN U3748 ( .A(n893), .B(A[599]), .Z(n3319) );
  AND U3749 ( .A(n3322), .B(n3323), .Z(n893) );
  NAND U3750 ( .A(B[598]), .B(n3324), .Z(n3323) );
  NANDN U3751 ( .A(A[598]), .B(n895), .Z(n3324) );
  NANDN U3752 ( .A(n895), .B(A[598]), .Z(n3322) );
  AND U3753 ( .A(n3325), .B(n3326), .Z(n895) );
  NAND U3754 ( .A(B[597]), .B(n3327), .Z(n3326) );
  NANDN U3755 ( .A(A[597]), .B(n897), .Z(n3327) );
  NANDN U3756 ( .A(n897), .B(A[597]), .Z(n3325) );
  AND U3757 ( .A(n3328), .B(n3329), .Z(n897) );
  NAND U3758 ( .A(B[596]), .B(n3330), .Z(n3329) );
  NANDN U3759 ( .A(A[596]), .B(n899), .Z(n3330) );
  NANDN U3760 ( .A(n899), .B(A[596]), .Z(n3328) );
  AND U3761 ( .A(n3331), .B(n3332), .Z(n899) );
  NAND U3762 ( .A(B[595]), .B(n3333), .Z(n3332) );
  NANDN U3763 ( .A(A[595]), .B(n901), .Z(n3333) );
  NANDN U3764 ( .A(n901), .B(A[595]), .Z(n3331) );
  AND U3765 ( .A(n3334), .B(n3335), .Z(n901) );
  NAND U3766 ( .A(B[594]), .B(n3336), .Z(n3335) );
  NANDN U3767 ( .A(A[594]), .B(n903), .Z(n3336) );
  NANDN U3768 ( .A(n903), .B(A[594]), .Z(n3334) );
  AND U3769 ( .A(n3337), .B(n3338), .Z(n903) );
  NAND U3770 ( .A(B[593]), .B(n3339), .Z(n3338) );
  NANDN U3771 ( .A(A[593]), .B(n905), .Z(n3339) );
  NANDN U3772 ( .A(n905), .B(A[593]), .Z(n3337) );
  AND U3773 ( .A(n3340), .B(n3341), .Z(n905) );
  NAND U3774 ( .A(B[592]), .B(n3342), .Z(n3341) );
  NANDN U3775 ( .A(A[592]), .B(n907), .Z(n3342) );
  NANDN U3776 ( .A(n907), .B(A[592]), .Z(n3340) );
  AND U3777 ( .A(n3343), .B(n3344), .Z(n907) );
  NAND U3778 ( .A(B[591]), .B(n3345), .Z(n3344) );
  NANDN U3779 ( .A(A[591]), .B(n909), .Z(n3345) );
  NANDN U3780 ( .A(n909), .B(A[591]), .Z(n3343) );
  AND U3781 ( .A(n3346), .B(n3347), .Z(n909) );
  NAND U3782 ( .A(B[590]), .B(n3348), .Z(n3347) );
  NANDN U3783 ( .A(A[590]), .B(n911), .Z(n3348) );
  NANDN U3784 ( .A(n911), .B(A[590]), .Z(n3346) );
  AND U3785 ( .A(n3349), .B(n3350), .Z(n911) );
  NAND U3786 ( .A(B[589]), .B(n3351), .Z(n3350) );
  NANDN U3787 ( .A(A[589]), .B(n915), .Z(n3351) );
  NANDN U3788 ( .A(n915), .B(A[589]), .Z(n3349) );
  AND U3789 ( .A(n3352), .B(n3353), .Z(n915) );
  NAND U3790 ( .A(B[588]), .B(n3354), .Z(n3353) );
  NANDN U3791 ( .A(A[588]), .B(n917), .Z(n3354) );
  NANDN U3792 ( .A(n917), .B(A[588]), .Z(n3352) );
  AND U3793 ( .A(n3355), .B(n3356), .Z(n917) );
  NAND U3794 ( .A(B[587]), .B(n3357), .Z(n3356) );
  NANDN U3795 ( .A(A[587]), .B(n919), .Z(n3357) );
  NANDN U3796 ( .A(n919), .B(A[587]), .Z(n3355) );
  AND U3797 ( .A(n3358), .B(n3359), .Z(n919) );
  NAND U3798 ( .A(B[586]), .B(n3360), .Z(n3359) );
  NANDN U3799 ( .A(A[586]), .B(n921), .Z(n3360) );
  NANDN U3800 ( .A(n921), .B(A[586]), .Z(n3358) );
  AND U3801 ( .A(n3361), .B(n3362), .Z(n921) );
  NAND U3802 ( .A(B[585]), .B(n3363), .Z(n3362) );
  NANDN U3803 ( .A(A[585]), .B(n923), .Z(n3363) );
  NANDN U3804 ( .A(n923), .B(A[585]), .Z(n3361) );
  AND U3805 ( .A(n3364), .B(n3365), .Z(n923) );
  NAND U3806 ( .A(B[584]), .B(n3366), .Z(n3365) );
  NANDN U3807 ( .A(A[584]), .B(n925), .Z(n3366) );
  NANDN U3808 ( .A(n925), .B(A[584]), .Z(n3364) );
  AND U3809 ( .A(n3367), .B(n3368), .Z(n925) );
  NAND U3810 ( .A(B[583]), .B(n3369), .Z(n3368) );
  NANDN U3811 ( .A(A[583]), .B(n927), .Z(n3369) );
  NANDN U3812 ( .A(n927), .B(A[583]), .Z(n3367) );
  AND U3813 ( .A(n3370), .B(n3371), .Z(n927) );
  NAND U3814 ( .A(B[582]), .B(n3372), .Z(n3371) );
  NANDN U3815 ( .A(A[582]), .B(n929), .Z(n3372) );
  NANDN U3816 ( .A(n929), .B(A[582]), .Z(n3370) );
  AND U3817 ( .A(n3373), .B(n3374), .Z(n929) );
  NAND U3818 ( .A(B[581]), .B(n3375), .Z(n3374) );
  NANDN U3819 ( .A(A[581]), .B(n931), .Z(n3375) );
  NANDN U3820 ( .A(n931), .B(A[581]), .Z(n3373) );
  AND U3821 ( .A(n3376), .B(n3377), .Z(n931) );
  NAND U3822 ( .A(B[580]), .B(n3378), .Z(n3377) );
  NANDN U3823 ( .A(A[580]), .B(n933), .Z(n3378) );
  NANDN U3824 ( .A(n933), .B(A[580]), .Z(n3376) );
  AND U3825 ( .A(n3379), .B(n3380), .Z(n933) );
  NAND U3826 ( .A(B[579]), .B(n3381), .Z(n3380) );
  NANDN U3827 ( .A(A[579]), .B(n937), .Z(n3381) );
  NANDN U3828 ( .A(n937), .B(A[579]), .Z(n3379) );
  AND U3829 ( .A(n3382), .B(n3383), .Z(n937) );
  NAND U3830 ( .A(B[578]), .B(n3384), .Z(n3383) );
  NANDN U3831 ( .A(A[578]), .B(n939), .Z(n3384) );
  NANDN U3832 ( .A(n939), .B(A[578]), .Z(n3382) );
  AND U3833 ( .A(n3385), .B(n3386), .Z(n939) );
  NAND U3834 ( .A(B[577]), .B(n3387), .Z(n3386) );
  NANDN U3835 ( .A(A[577]), .B(n941), .Z(n3387) );
  NANDN U3836 ( .A(n941), .B(A[577]), .Z(n3385) );
  AND U3837 ( .A(n3388), .B(n3389), .Z(n941) );
  NAND U3838 ( .A(B[576]), .B(n3390), .Z(n3389) );
  NANDN U3839 ( .A(A[576]), .B(n943), .Z(n3390) );
  NANDN U3840 ( .A(n943), .B(A[576]), .Z(n3388) );
  AND U3841 ( .A(n3391), .B(n3392), .Z(n943) );
  NAND U3842 ( .A(B[575]), .B(n3393), .Z(n3392) );
  NANDN U3843 ( .A(A[575]), .B(n945), .Z(n3393) );
  NANDN U3844 ( .A(n945), .B(A[575]), .Z(n3391) );
  AND U3845 ( .A(n3394), .B(n3395), .Z(n945) );
  NAND U3846 ( .A(B[574]), .B(n3396), .Z(n3395) );
  NANDN U3847 ( .A(A[574]), .B(n947), .Z(n3396) );
  NANDN U3848 ( .A(n947), .B(A[574]), .Z(n3394) );
  AND U3849 ( .A(n3397), .B(n3398), .Z(n947) );
  NAND U3850 ( .A(B[573]), .B(n3399), .Z(n3398) );
  NANDN U3851 ( .A(A[573]), .B(n949), .Z(n3399) );
  NANDN U3852 ( .A(n949), .B(A[573]), .Z(n3397) );
  AND U3853 ( .A(n3400), .B(n3401), .Z(n949) );
  NAND U3854 ( .A(B[572]), .B(n3402), .Z(n3401) );
  NANDN U3855 ( .A(A[572]), .B(n951), .Z(n3402) );
  NANDN U3856 ( .A(n951), .B(A[572]), .Z(n3400) );
  AND U3857 ( .A(n3403), .B(n3404), .Z(n951) );
  NAND U3858 ( .A(B[571]), .B(n3405), .Z(n3404) );
  NANDN U3859 ( .A(A[571]), .B(n953), .Z(n3405) );
  NANDN U3860 ( .A(n953), .B(A[571]), .Z(n3403) );
  AND U3861 ( .A(n3406), .B(n3407), .Z(n953) );
  NAND U3862 ( .A(B[570]), .B(n3408), .Z(n3407) );
  NANDN U3863 ( .A(A[570]), .B(n955), .Z(n3408) );
  NANDN U3864 ( .A(n955), .B(A[570]), .Z(n3406) );
  AND U3865 ( .A(n3409), .B(n3410), .Z(n955) );
  NAND U3866 ( .A(B[569]), .B(n3411), .Z(n3410) );
  NANDN U3867 ( .A(A[569]), .B(n959), .Z(n3411) );
  NANDN U3868 ( .A(n959), .B(A[569]), .Z(n3409) );
  AND U3869 ( .A(n3412), .B(n3413), .Z(n959) );
  NAND U3870 ( .A(B[568]), .B(n3414), .Z(n3413) );
  NANDN U3871 ( .A(A[568]), .B(n961), .Z(n3414) );
  NANDN U3872 ( .A(n961), .B(A[568]), .Z(n3412) );
  AND U3873 ( .A(n3415), .B(n3416), .Z(n961) );
  NAND U3874 ( .A(B[567]), .B(n3417), .Z(n3416) );
  NANDN U3875 ( .A(A[567]), .B(n963), .Z(n3417) );
  NANDN U3876 ( .A(n963), .B(A[567]), .Z(n3415) );
  AND U3877 ( .A(n3418), .B(n3419), .Z(n963) );
  NAND U3878 ( .A(B[566]), .B(n3420), .Z(n3419) );
  NANDN U3879 ( .A(A[566]), .B(n965), .Z(n3420) );
  NANDN U3880 ( .A(n965), .B(A[566]), .Z(n3418) );
  AND U3881 ( .A(n3421), .B(n3422), .Z(n965) );
  NAND U3882 ( .A(B[565]), .B(n3423), .Z(n3422) );
  NANDN U3883 ( .A(A[565]), .B(n967), .Z(n3423) );
  NANDN U3884 ( .A(n967), .B(A[565]), .Z(n3421) );
  AND U3885 ( .A(n3424), .B(n3425), .Z(n967) );
  NAND U3886 ( .A(B[564]), .B(n3426), .Z(n3425) );
  NANDN U3887 ( .A(A[564]), .B(n969), .Z(n3426) );
  NANDN U3888 ( .A(n969), .B(A[564]), .Z(n3424) );
  AND U3889 ( .A(n3427), .B(n3428), .Z(n969) );
  NAND U3890 ( .A(B[563]), .B(n3429), .Z(n3428) );
  NANDN U3891 ( .A(A[563]), .B(n971), .Z(n3429) );
  NANDN U3892 ( .A(n971), .B(A[563]), .Z(n3427) );
  AND U3893 ( .A(n3430), .B(n3431), .Z(n971) );
  NAND U3894 ( .A(B[562]), .B(n3432), .Z(n3431) );
  NANDN U3895 ( .A(A[562]), .B(n973), .Z(n3432) );
  NANDN U3896 ( .A(n973), .B(A[562]), .Z(n3430) );
  AND U3897 ( .A(n3433), .B(n3434), .Z(n973) );
  NAND U3898 ( .A(B[561]), .B(n3435), .Z(n3434) );
  NANDN U3899 ( .A(A[561]), .B(n975), .Z(n3435) );
  NANDN U3900 ( .A(n975), .B(A[561]), .Z(n3433) );
  AND U3901 ( .A(n3436), .B(n3437), .Z(n975) );
  NAND U3902 ( .A(B[560]), .B(n3438), .Z(n3437) );
  NANDN U3903 ( .A(A[560]), .B(n977), .Z(n3438) );
  NANDN U3904 ( .A(n977), .B(A[560]), .Z(n3436) );
  AND U3905 ( .A(n3439), .B(n3440), .Z(n977) );
  NAND U3906 ( .A(B[559]), .B(n3441), .Z(n3440) );
  NANDN U3907 ( .A(A[559]), .B(n981), .Z(n3441) );
  NANDN U3908 ( .A(n981), .B(A[559]), .Z(n3439) );
  AND U3909 ( .A(n3442), .B(n3443), .Z(n981) );
  NAND U3910 ( .A(B[558]), .B(n3444), .Z(n3443) );
  NANDN U3911 ( .A(A[558]), .B(n983), .Z(n3444) );
  NANDN U3912 ( .A(n983), .B(A[558]), .Z(n3442) );
  AND U3913 ( .A(n3445), .B(n3446), .Z(n983) );
  NAND U3914 ( .A(B[557]), .B(n3447), .Z(n3446) );
  NANDN U3915 ( .A(A[557]), .B(n985), .Z(n3447) );
  NANDN U3916 ( .A(n985), .B(A[557]), .Z(n3445) );
  AND U3917 ( .A(n3448), .B(n3449), .Z(n985) );
  NAND U3918 ( .A(B[556]), .B(n3450), .Z(n3449) );
  NANDN U3919 ( .A(A[556]), .B(n987), .Z(n3450) );
  NANDN U3920 ( .A(n987), .B(A[556]), .Z(n3448) );
  AND U3921 ( .A(n3451), .B(n3452), .Z(n987) );
  NAND U3922 ( .A(B[555]), .B(n3453), .Z(n3452) );
  NANDN U3923 ( .A(A[555]), .B(n989), .Z(n3453) );
  NANDN U3924 ( .A(n989), .B(A[555]), .Z(n3451) );
  AND U3925 ( .A(n3454), .B(n3455), .Z(n989) );
  NAND U3926 ( .A(B[554]), .B(n3456), .Z(n3455) );
  NANDN U3927 ( .A(A[554]), .B(n991), .Z(n3456) );
  NANDN U3928 ( .A(n991), .B(A[554]), .Z(n3454) );
  AND U3929 ( .A(n3457), .B(n3458), .Z(n991) );
  NAND U3930 ( .A(B[553]), .B(n3459), .Z(n3458) );
  NANDN U3931 ( .A(A[553]), .B(n993), .Z(n3459) );
  NANDN U3932 ( .A(n993), .B(A[553]), .Z(n3457) );
  AND U3933 ( .A(n3460), .B(n3461), .Z(n993) );
  NAND U3934 ( .A(B[552]), .B(n3462), .Z(n3461) );
  NANDN U3935 ( .A(A[552]), .B(n995), .Z(n3462) );
  NANDN U3936 ( .A(n995), .B(A[552]), .Z(n3460) );
  AND U3937 ( .A(n3463), .B(n3464), .Z(n995) );
  NAND U3938 ( .A(B[551]), .B(n3465), .Z(n3464) );
  NANDN U3939 ( .A(A[551]), .B(n997), .Z(n3465) );
  NANDN U3940 ( .A(n997), .B(A[551]), .Z(n3463) );
  AND U3941 ( .A(n3466), .B(n3467), .Z(n997) );
  NAND U3942 ( .A(B[550]), .B(n3468), .Z(n3467) );
  NANDN U3943 ( .A(A[550]), .B(n999), .Z(n3468) );
  NANDN U3944 ( .A(n999), .B(A[550]), .Z(n3466) );
  AND U3945 ( .A(n3469), .B(n3470), .Z(n999) );
  NAND U3946 ( .A(B[549]), .B(n3471), .Z(n3470) );
  NANDN U3947 ( .A(A[549]), .B(n1003), .Z(n3471) );
  NANDN U3948 ( .A(n1003), .B(A[549]), .Z(n3469) );
  AND U3949 ( .A(n3472), .B(n3473), .Z(n1003) );
  NAND U3950 ( .A(B[548]), .B(n3474), .Z(n3473) );
  NANDN U3951 ( .A(A[548]), .B(n1005), .Z(n3474) );
  NANDN U3952 ( .A(n1005), .B(A[548]), .Z(n3472) );
  AND U3953 ( .A(n3475), .B(n3476), .Z(n1005) );
  NAND U3954 ( .A(B[547]), .B(n3477), .Z(n3476) );
  NANDN U3955 ( .A(A[547]), .B(n1007), .Z(n3477) );
  NANDN U3956 ( .A(n1007), .B(A[547]), .Z(n3475) );
  AND U3957 ( .A(n3478), .B(n3479), .Z(n1007) );
  NAND U3958 ( .A(B[546]), .B(n3480), .Z(n3479) );
  NANDN U3959 ( .A(A[546]), .B(n1009), .Z(n3480) );
  NANDN U3960 ( .A(n1009), .B(A[546]), .Z(n3478) );
  AND U3961 ( .A(n3481), .B(n3482), .Z(n1009) );
  NAND U3962 ( .A(B[545]), .B(n3483), .Z(n3482) );
  NANDN U3963 ( .A(A[545]), .B(n1011), .Z(n3483) );
  NANDN U3964 ( .A(n1011), .B(A[545]), .Z(n3481) );
  AND U3965 ( .A(n3484), .B(n3485), .Z(n1011) );
  NAND U3966 ( .A(B[544]), .B(n3486), .Z(n3485) );
  NANDN U3967 ( .A(A[544]), .B(n1013), .Z(n3486) );
  NANDN U3968 ( .A(n1013), .B(A[544]), .Z(n3484) );
  AND U3969 ( .A(n3487), .B(n3488), .Z(n1013) );
  NAND U3970 ( .A(B[543]), .B(n3489), .Z(n3488) );
  NANDN U3971 ( .A(A[543]), .B(n1015), .Z(n3489) );
  NANDN U3972 ( .A(n1015), .B(A[543]), .Z(n3487) );
  AND U3973 ( .A(n3490), .B(n3491), .Z(n1015) );
  NAND U3974 ( .A(B[542]), .B(n3492), .Z(n3491) );
  NANDN U3975 ( .A(A[542]), .B(n1017), .Z(n3492) );
  NANDN U3976 ( .A(n1017), .B(A[542]), .Z(n3490) );
  AND U3977 ( .A(n3493), .B(n3494), .Z(n1017) );
  NAND U3978 ( .A(B[541]), .B(n3495), .Z(n3494) );
  NANDN U3979 ( .A(A[541]), .B(n1019), .Z(n3495) );
  NANDN U3980 ( .A(n1019), .B(A[541]), .Z(n3493) );
  AND U3981 ( .A(n3496), .B(n3497), .Z(n1019) );
  NAND U3982 ( .A(B[540]), .B(n3498), .Z(n3497) );
  NANDN U3983 ( .A(A[540]), .B(n1021), .Z(n3498) );
  NANDN U3984 ( .A(n1021), .B(A[540]), .Z(n3496) );
  AND U3985 ( .A(n3499), .B(n3500), .Z(n1021) );
  NAND U3986 ( .A(B[539]), .B(n3501), .Z(n3500) );
  NANDN U3987 ( .A(A[539]), .B(n1025), .Z(n3501) );
  NANDN U3988 ( .A(n1025), .B(A[539]), .Z(n3499) );
  AND U3989 ( .A(n3502), .B(n3503), .Z(n1025) );
  NAND U3990 ( .A(B[538]), .B(n3504), .Z(n3503) );
  NANDN U3991 ( .A(A[538]), .B(n1027), .Z(n3504) );
  NANDN U3992 ( .A(n1027), .B(A[538]), .Z(n3502) );
  AND U3993 ( .A(n3505), .B(n3506), .Z(n1027) );
  NAND U3994 ( .A(B[537]), .B(n3507), .Z(n3506) );
  NANDN U3995 ( .A(A[537]), .B(n1029), .Z(n3507) );
  NANDN U3996 ( .A(n1029), .B(A[537]), .Z(n3505) );
  AND U3997 ( .A(n3508), .B(n3509), .Z(n1029) );
  NAND U3998 ( .A(B[536]), .B(n3510), .Z(n3509) );
  NANDN U3999 ( .A(A[536]), .B(n1031), .Z(n3510) );
  NANDN U4000 ( .A(n1031), .B(A[536]), .Z(n3508) );
  AND U4001 ( .A(n3511), .B(n3512), .Z(n1031) );
  NAND U4002 ( .A(B[535]), .B(n3513), .Z(n3512) );
  NANDN U4003 ( .A(A[535]), .B(n1033), .Z(n3513) );
  NANDN U4004 ( .A(n1033), .B(A[535]), .Z(n3511) );
  AND U4005 ( .A(n3514), .B(n3515), .Z(n1033) );
  NAND U4006 ( .A(B[534]), .B(n3516), .Z(n3515) );
  NANDN U4007 ( .A(A[534]), .B(n1035), .Z(n3516) );
  NANDN U4008 ( .A(n1035), .B(A[534]), .Z(n3514) );
  AND U4009 ( .A(n3517), .B(n3518), .Z(n1035) );
  NAND U4010 ( .A(B[533]), .B(n3519), .Z(n3518) );
  NANDN U4011 ( .A(A[533]), .B(n1037), .Z(n3519) );
  NANDN U4012 ( .A(n1037), .B(A[533]), .Z(n3517) );
  AND U4013 ( .A(n3520), .B(n3521), .Z(n1037) );
  NAND U4014 ( .A(B[532]), .B(n3522), .Z(n3521) );
  NANDN U4015 ( .A(A[532]), .B(n1039), .Z(n3522) );
  NANDN U4016 ( .A(n1039), .B(A[532]), .Z(n3520) );
  AND U4017 ( .A(n3523), .B(n3524), .Z(n1039) );
  NAND U4018 ( .A(B[531]), .B(n3525), .Z(n3524) );
  NANDN U4019 ( .A(A[531]), .B(n1041), .Z(n3525) );
  NANDN U4020 ( .A(n1041), .B(A[531]), .Z(n3523) );
  AND U4021 ( .A(n3526), .B(n3527), .Z(n1041) );
  NAND U4022 ( .A(B[530]), .B(n3528), .Z(n3527) );
  NANDN U4023 ( .A(A[530]), .B(n1043), .Z(n3528) );
  NANDN U4024 ( .A(n1043), .B(A[530]), .Z(n3526) );
  AND U4025 ( .A(n3529), .B(n3530), .Z(n1043) );
  NAND U4026 ( .A(B[529]), .B(n3531), .Z(n3530) );
  NANDN U4027 ( .A(A[529]), .B(n1047), .Z(n3531) );
  NANDN U4028 ( .A(n1047), .B(A[529]), .Z(n3529) );
  AND U4029 ( .A(n3532), .B(n3533), .Z(n1047) );
  NAND U4030 ( .A(B[528]), .B(n3534), .Z(n3533) );
  NANDN U4031 ( .A(A[528]), .B(n1049), .Z(n3534) );
  NANDN U4032 ( .A(n1049), .B(A[528]), .Z(n3532) );
  AND U4033 ( .A(n3535), .B(n3536), .Z(n1049) );
  NAND U4034 ( .A(B[527]), .B(n3537), .Z(n3536) );
  NANDN U4035 ( .A(A[527]), .B(n1051), .Z(n3537) );
  NANDN U4036 ( .A(n1051), .B(A[527]), .Z(n3535) );
  AND U4037 ( .A(n3538), .B(n3539), .Z(n1051) );
  NAND U4038 ( .A(B[526]), .B(n3540), .Z(n3539) );
  NANDN U4039 ( .A(A[526]), .B(n1053), .Z(n3540) );
  NANDN U4040 ( .A(n1053), .B(A[526]), .Z(n3538) );
  AND U4041 ( .A(n3541), .B(n3542), .Z(n1053) );
  NAND U4042 ( .A(B[525]), .B(n3543), .Z(n3542) );
  NANDN U4043 ( .A(A[525]), .B(n1055), .Z(n3543) );
  NANDN U4044 ( .A(n1055), .B(A[525]), .Z(n3541) );
  AND U4045 ( .A(n3544), .B(n3545), .Z(n1055) );
  NAND U4046 ( .A(B[524]), .B(n3546), .Z(n3545) );
  NANDN U4047 ( .A(A[524]), .B(n1057), .Z(n3546) );
  NANDN U4048 ( .A(n1057), .B(A[524]), .Z(n3544) );
  AND U4049 ( .A(n3547), .B(n3548), .Z(n1057) );
  NAND U4050 ( .A(B[523]), .B(n3549), .Z(n3548) );
  NANDN U4051 ( .A(A[523]), .B(n1059), .Z(n3549) );
  NANDN U4052 ( .A(n1059), .B(A[523]), .Z(n3547) );
  AND U4053 ( .A(n3550), .B(n3551), .Z(n1059) );
  NAND U4054 ( .A(B[522]), .B(n3552), .Z(n3551) );
  NANDN U4055 ( .A(A[522]), .B(n1061), .Z(n3552) );
  NANDN U4056 ( .A(n1061), .B(A[522]), .Z(n3550) );
  AND U4057 ( .A(n3553), .B(n3554), .Z(n1061) );
  NAND U4058 ( .A(B[521]), .B(n3555), .Z(n3554) );
  NANDN U4059 ( .A(A[521]), .B(n1063), .Z(n3555) );
  NANDN U4060 ( .A(n1063), .B(A[521]), .Z(n3553) );
  AND U4061 ( .A(n3556), .B(n3557), .Z(n1063) );
  NAND U4062 ( .A(B[520]), .B(n3558), .Z(n3557) );
  NANDN U4063 ( .A(A[520]), .B(n1065), .Z(n3558) );
  NANDN U4064 ( .A(n1065), .B(A[520]), .Z(n3556) );
  AND U4065 ( .A(n3559), .B(n3560), .Z(n1065) );
  NAND U4066 ( .A(B[519]), .B(n3561), .Z(n3560) );
  NANDN U4067 ( .A(A[519]), .B(n1069), .Z(n3561) );
  NANDN U4068 ( .A(n1069), .B(A[519]), .Z(n3559) );
  AND U4069 ( .A(n3562), .B(n3563), .Z(n1069) );
  NAND U4070 ( .A(B[518]), .B(n3564), .Z(n3563) );
  NANDN U4071 ( .A(A[518]), .B(n1071), .Z(n3564) );
  NANDN U4072 ( .A(n1071), .B(A[518]), .Z(n3562) );
  AND U4073 ( .A(n3565), .B(n3566), .Z(n1071) );
  NAND U4074 ( .A(B[517]), .B(n3567), .Z(n3566) );
  NANDN U4075 ( .A(A[517]), .B(n1073), .Z(n3567) );
  NANDN U4076 ( .A(n1073), .B(A[517]), .Z(n3565) );
  AND U4077 ( .A(n3568), .B(n3569), .Z(n1073) );
  NAND U4078 ( .A(B[516]), .B(n3570), .Z(n3569) );
  NANDN U4079 ( .A(A[516]), .B(n1075), .Z(n3570) );
  NANDN U4080 ( .A(n1075), .B(A[516]), .Z(n3568) );
  AND U4081 ( .A(n3571), .B(n3572), .Z(n1075) );
  NAND U4082 ( .A(B[515]), .B(n3573), .Z(n3572) );
  NANDN U4083 ( .A(A[515]), .B(n1077), .Z(n3573) );
  NANDN U4084 ( .A(n1077), .B(A[515]), .Z(n3571) );
  AND U4085 ( .A(n3574), .B(n3575), .Z(n1077) );
  NAND U4086 ( .A(B[514]), .B(n3576), .Z(n3575) );
  NANDN U4087 ( .A(A[514]), .B(n1079), .Z(n3576) );
  NANDN U4088 ( .A(n1079), .B(A[514]), .Z(n3574) );
  AND U4089 ( .A(n3577), .B(n3578), .Z(n1079) );
  NAND U4090 ( .A(B[513]), .B(n3579), .Z(n3578) );
  NANDN U4091 ( .A(A[513]), .B(n1081), .Z(n3579) );
  NANDN U4092 ( .A(n1081), .B(A[513]), .Z(n3577) );
  AND U4093 ( .A(n3580), .B(n3581), .Z(n1081) );
  NAND U4094 ( .A(B[512]), .B(n3582), .Z(n3581) );
  NANDN U4095 ( .A(A[512]), .B(n1083), .Z(n3582) );
  NANDN U4096 ( .A(n1083), .B(A[512]), .Z(n3580) );
  AND U4097 ( .A(n3583), .B(n3584), .Z(n1083) );
  NAND U4098 ( .A(B[511]), .B(n3585), .Z(n3584) );
  NANDN U4099 ( .A(A[511]), .B(n1085), .Z(n3585) );
  NANDN U4100 ( .A(n1085), .B(A[511]), .Z(n3583) );
  AND U4101 ( .A(n3586), .B(n3587), .Z(n1085) );
  NAND U4102 ( .A(B[510]), .B(n3588), .Z(n3587) );
  NANDN U4103 ( .A(A[510]), .B(n1087), .Z(n3588) );
  NANDN U4104 ( .A(n1087), .B(A[510]), .Z(n3586) );
  AND U4105 ( .A(n3589), .B(n3590), .Z(n1087) );
  NAND U4106 ( .A(B[509]), .B(n3591), .Z(n3590) );
  NANDN U4107 ( .A(A[509]), .B(n1091), .Z(n3591) );
  NANDN U4108 ( .A(n1091), .B(A[509]), .Z(n3589) );
  AND U4109 ( .A(n3592), .B(n3593), .Z(n1091) );
  NAND U4110 ( .A(B[508]), .B(n3594), .Z(n3593) );
  NANDN U4111 ( .A(A[508]), .B(n1093), .Z(n3594) );
  NANDN U4112 ( .A(n1093), .B(A[508]), .Z(n3592) );
  AND U4113 ( .A(n3595), .B(n3596), .Z(n1093) );
  NAND U4114 ( .A(B[507]), .B(n3597), .Z(n3596) );
  NANDN U4115 ( .A(A[507]), .B(n1095), .Z(n3597) );
  NANDN U4116 ( .A(n1095), .B(A[507]), .Z(n3595) );
  AND U4117 ( .A(n3598), .B(n3599), .Z(n1095) );
  NAND U4118 ( .A(B[506]), .B(n3600), .Z(n3599) );
  NANDN U4119 ( .A(A[506]), .B(n1097), .Z(n3600) );
  NANDN U4120 ( .A(n1097), .B(A[506]), .Z(n3598) );
  AND U4121 ( .A(n3601), .B(n3602), .Z(n1097) );
  NAND U4122 ( .A(B[505]), .B(n3603), .Z(n3602) );
  NANDN U4123 ( .A(A[505]), .B(n1099), .Z(n3603) );
  NANDN U4124 ( .A(n1099), .B(A[505]), .Z(n3601) );
  AND U4125 ( .A(n3604), .B(n3605), .Z(n1099) );
  NAND U4126 ( .A(B[504]), .B(n3606), .Z(n3605) );
  NANDN U4127 ( .A(A[504]), .B(n1101), .Z(n3606) );
  NANDN U4128 ( .A(n1101), .B(A[504]), .Z(n3604) );
  AND U4129 ( .A(n3607), .B(n3608), .Z(n1101) );
  NAND U4130 ( .A(B[503]), .B(n3609), .Z(n3608) );
  NANDN U4131 ( .A(A[503]), .B(n1103), .Z(n3609) );
  NANDN U4132 ( .A(n1103), .B(A[503]), .Z(n3607) );
  AND U4133 ( .A(n3610), .B(n3611), .Z(n1103) );
  NAND U4134 ( .A(B[502]), .B(n3612), .Z(n3611) );
  NANDN U4135 ( .A(A[502]), .B(n1105), .Z(n3612) );
  NANDN U4136 ( .A(n1105), .B(A[502]), .Z(n3610) );
  AND U4137 ( .A(n3613), .B(n3614), .Z(n1105) );
  NAND U4138 ( .A(B[501]), .B(n3615), .Z(n3614) );
  NANDN U4139 ( .A(A[501]), .B(n1107), .Z(n3615) );
  NANDN U4140 ( .A(n1107), .B(A[501]), .Z(n3613) );
  AND U4141 ( .A(n3616), .B(n3617), .Z(n1107) );
  NAND U4142 ( .A(B[500]), .B(n3618), .Z(n3617) );
  NANDN U4143 ( .A(A[500]), .B(n1109), .Z(n3618) );
  NANDN U4144 ( .A(n1109), .B(A[500]), .Z(n3616) );
  AND U4145 ( .A(n3619), .B(n3620), .Z(n1109) );
  NAND U4146 ( .A(B[499]), .B(n3621), .Z(n3620) );
  NANDN U4147 ( .A(A[499]), .B(n1115), .Z(n3621) );
  NANDN U4148 ( .A(n1115), .B(A[499]), .Z(n3619) );
  AND U4149 ( .A(n3622), .B(n3623), .Z(n1115) );
  NAND U4150 ( .A(B[498]), .B(n3624), .Z(n3623) );
  NANDN U4151 ( .A(A[498]), .B(n1117), .Z(n3624) );
  NANDN U4152 ( .A(n1117), .B(A[498]), .Z(n3622) );
  AND U4153 ( .A(n3625), .B(n3626), .Z(n1117) );
  NAND U4154 ( .A(B[497]), .B(n3627), .Z(n3626) );
  NANDN U4155 ( .A(A[497]), .B(n1119), .Z(n3627) );
  NANDN U4156 ( .A(n1119), .B(A[497]), .Z(n3625) );
  AND U4157 ( .A(n3628), .B(n3629), .Z(n1119) );
  NAND U4158 ( .A(B[496]), .B(n3630), .Z(n3629) );
  NANDN U4159 ( .A(A[496]), .B(n1121), .Z(n3630) );
  NANDN U4160 ( .A(n1121), .B(A[496]), .Z(n3628) );
  AND U4161 ( .A(n3631), .B(n3632), .Z(n1121) );
  NAND U4162 ( .A(B[495]), .B(n3633), .Z(n3632) );
  NANDN U4163 ( .A(A[495]), .B(n1123), .Z(n3633) );
  NANDN U4164 ( .A(n1123), .B(A[495]), .Z(n3631) );
  AND U4165 ( .A(n3634), .B(n3635), .Z(n1123) );
  NAND U4166 ( .A(B[494]), .B(n3636), .Z(n3635) );
  NANDN U4167 ( .A(A[494]), .B(n1125), .Z(n3636) );
  NANDN U4168 ( .A(n1125), .B(A[494]), .Z(n3634) );
  AND U4169 ( .A(n3637), .B(n3638), .Z(n1125) );
  NAND U4170 ( .A(B[493]), .B(n3639), .Z(n3638) );
  NANDN U4171 ( .A(A[493]), .B(n1127), .Z(n3639) );
  NANDN U4172 ( .A(n1127), .B(A[493]), .Z(n3637) );
  AND U4173 ( .A(n3640), .B(n3641), .Z(n1127) );
  NAND U4174 ( .A(B[492]), .B(n3642), .Z(n3641) );
  NANDN U4175 ( .A(A[492]), .B(n1129), .Z(n3642) );
  NANDN U4176 ( .A(n1129), .B(A[492]), .Z(n3640) );
  AND U4177 ( .A(n3643), .B(n3644), .Z(n1129) );
  NAND U4178 ( .A(B[491]), .B(n3645), .Z(n3644) );
  NANDN U4179 ( .A(A[491]), .B(n1131), .Z(n3645) );
  NANDN U4180 ( .A(n1131), .B(A[491]), .Z(n3643) );
  AND U4181 ( .A(n3646), .B(n3647), .Z(n1131) );
  NAND U4182 ( .A(B[490]), .B(n3648), .Z(n3647) );
  NANDN U4183 ( .A(A[490]), .B(n1133), .Z(n3648) );
  NANDN U4184 ( .A(n1133), .B(A[490]), .Z(n3646) );
  AND U4185 ( .A(n3649), .B(n3650), .Z(n1133) );
  NAND U4186 ( .A(B[489]), .B(n3651), .Z(n3650) );
  NANDN U4187 ( .A(A[489]), .B(n1137), .Z(n3651) );
  NANDN U4188 ( .A(n1137), .B(A[489]), .Z(n3649) );
  AND U4189 ( .A(n3652), .B(n3653), .Z(n1137) );
  NAND U4190 ( .A(B[488]), .B(n3654), .Z(n3653) );
  NANDN U4191 ( .A(A[488]), .B(n1139), .Z(n3654) );
  NANDN U4192 ( .A(n1139), .B(A[488]), .Z(n3652) );
  AND U4193 ( .A(n3655), .B(n3656), .Z(n1139) );
  NAND U4194 ( .A(B[487]), .B(n3657), .Z(n3656) );
  NANDN U4195 ( .A(A[487]), .B(n1141), .Z(n3657) );
  NANDN U4196 ( .A(n1141), .B(A[487]), .Z(n3655) );
  AND U4197 ( .A(n3658), .B(n3659), .Z(n1141) );
  NAND U4198 ( .A(B[486]), .B(n3660), .Z(n3659) );
  NANDN U4199 ( .A(A[486]), .B(n1143), .Z(n3660) );
  NANDN U4200 ( .A(n1143), .B(A[486]), .Z(n3658) );
  AND U4201 ( .A(n3661), .B(n3662), .Z(n1143) );
  NAND U4202 ( .A(B[485]), .B(n3663), .Z(n3662) );
  NANDN U4203 ( .A(A[485]), .B(n1145), .Z(n3663) );
  NANDN U4204 ( .A(n1145), .B(A[485]), .Z(n3661) );
  AND U4205 ( .A(n3664), .B(n3665), .Z(n1145) );
  NAND U4206 ( .A(B[484]), .B(n3666), .Z(n3665) );
  NANDN U4207 ( .A(A[484]), .B(n1147), .Z(n3666) );
  NANDN U4208 ( .A(n1147), .B(A[484]), .Z(n3664) );
  AND U4209 ( .A(n3667), .B(n3668), .Z(n1147) );
  NAND U4210 ( .A(B[483]), .B(n3669), .Z(n3668) );
  NANDN U4211 ( .A(A[483]), .B(n1149), .Z(n3669) );
  NANDN U4212 ( .A(n1149), .B(A[483]), .Z(n3667) );
  AND U4213 ( .A(n3670), .B(n3671), .Z(n1149) );
  NAND U4214 ( .A(B[482]), .B(n3672), .Z(n3671) );
  NANDN U4215 ( .A(A[482]), .B(n1151), .Z(n3672) );
  NANDN U4216 ( .A(n1151), .B(A[482]), .Z(n3670) );
  AND U4217 ( .A(n3673), .B(n3674), .Z(n1151) );
  NAND U4218 ( .A(B[481]), .B(n3675), .Z(n3674) );
  NANDN U4219 ( .A(A[481]), .B(n1153), .Z(n3675) );
  NANDN U4220 ( .A(n1153), .B(A[481]), .Z(n3673) );
  AND U4221 ( .A(n3676), .B(n3677), .Z(n1153) );
  NAND U4222 ( .A(B[480]), .B(n3678), .Z(n3677) );
  NANDN U4223 ( .A(A[480]), .B(n1155), .Z(n3678) );
  NANDN U4224 ( .A(n1155), .B(A[480]), .Z(n3676) );
  AND U4225 ( .A(n3679), .B(n3680), .Z(n1155) );
  NAND U4226 ( .A(B[479]), .B(n3681), .Z(n3680) );
  NANDN U4227 ( .A(A[479]), .B(n1159), .Z(n3681) );
  NANDN U4228 ( .A(n1159), .B(A[479]), .Z(n3679) );
  AND U4229 ( .A(n3682), .B(n3683), .Z(n1159) );
  NAND U4230 ( .A(B[478]), .B(n3684), .Z(n3683) );
  NANDN U4231 ( .A(A[478]), .B(n1161), .Z(n3684) );
  NANDN U4232 ( .A(n1161), .B(A[478]), .Z(n3682) );
  AND U4233 ( .A(n3685), .B(n3686), .Z(n1161) );
  NAND U4234 ( .A(B[477]), .B(n3687), .Z(n3686) );
  NANDN U4235 ( .A(A[477]), .B(n1163), .Z(n3687) );
  NANDN U4236 ( .A(n1163), .B(A[477]), .Z(n3685) );
  AND U4237 ( .A(n3688), .B(n3689), .Z(n1163) );
  NAND U4238 ( .A(B[476]), .B(n3690), .Z(n3689) );
  NANDN U4239 ( .A(A[476]), .B(n1165), .Z(n3690) );
  NANDN U4240 ( .A(n1165), .B(A[476]), .Z(n3688) );
  AND U4241 ( .A(n3691), .B(n3692), .Z(n1165) );
  NAND U4242 ( .A(B[475]), .B(n3693), .Z(n3692) );
  NANDN U4243 ( .A(A[475]), .B(n1167), .Z(n3693) );
  NANDN U4244 ( .A(n1167), .B(A[475]), .Z(n3691) );
  AND U4245 ( .A(n3694), .B(n3695), .Z(n1167) );
  NAND U4246 ( .A(B[474]), .B(n3696), .Z(n3695) );
  NANDN U4247 ( .A(A[474]), .B(n1169), .Z(n3696) );
  NANDN U4248 ( .A(n1169), .B(A[474]), .Z(n3694) );
  AND U4249 ( .A(n3697), .B(n3698), .Z(n1169) );
  NAND U4250 ( .A(B[473]), .B(n3699), .Z(n3698) );
  NANDN U4251 ( .A(A[473]), .B(n1171), .Z(n3699) );
  NANDN U4252 ( .A(n1171), .B(A[473]), .Z(n3697) );
  AND U4253 ( .A(n3700), .B(n3701), .Z(n1171) );
  NAND U4254 ( .A(B[472]), .B(n3702), .Z(n3701) );
  NANDN U4255 ( .A(A[472]), .B(n1173), .Z(n3702) );
  NANDN U4256 ( .A(n1173), .B(A[472]), .Z(n3700) );
  AND U4257 ( .A(n3703), .B(n3704), .Z(n1173) );
  NAND U4258 ( .A(B[471]), .B(n3705), .Z(n3704) );
  NANDN U4259 ( .A(A[471]), .B(n1175), .Z(n3705) );
  NANDN U4260 ( .A(n1175), .B(A[471]), .Z(n3703) );
  AND U4261 ( .A(n3706), .B(n3707), .Z(n1175) );
  NAND U4262 ( .A(B[470]), .B(n3708), .Z(n3707) );
  NANDN U4263 ( .A(A[470]), .B(n1177), .Z(n3708) );
  NANDN U4264 ( .A(n1177), .B(A[470]), .Z(n3706) );
  AND U4265 ( .A(n3709), .B(n3710), .Z(n1177) );
  NAND U4266 ( .A(B[469]), .B(n3711), .Z(n3710) );
  NANDN U4267 ( .A(A[469]), .B(n1181), .Z(n3711) );
  NANDN U4268 ( .A(n1181), .B(A[469]), .Z(n3709) );
  AND U4269 ( .A(n3712), .B(n3713), .Z(n1181) );
  NAND U4270 ( .A(B[468]), .B(n3714), .Z(n3713) );
  NANDN U4271 ( .A(A[468]), .B(n1183), .Z(n3714) );
  NANDN U4272 ( .A(n1183), .B(A[468]), .Z(n3712) );
  AND U4273 ( .A(n3715), .B(n3716), .Z(n1183) );
  NAND U4274 ( .A(B[467]), .B(n3717), .Z(n3716) );
  NANDN U4275 ( .A(A[467]), .B(n1185), .Z(n3717) );
  NANDN U4276 ( .A(n1185), .B(A[467]), .Z(n3715) );
  AND U4277 ( .A(n3718), .B(n3719), .Z(n1185) );
  NAND U4278 ( .A(B[466]), .B(n3720), .Z(n3719) );
  NANDN U4279 ( .A(A[466]), .B(n1187), .Z(n3720) );
  NANDN U4280 ( .A(n1187), .B(A[466]), .Z(n3718) );
  AND U4281 ( .A(n3721), .B(n3722), .Z(n1187) );
  NAND U4282 ( .A(B[465]), .B(n3723), .Z(n3722) );
  NANDN U4283 ( .A(A[465]), .B(n1189), .Z(n3723) );
  NANDN U4284 ( .A(n1189), .B(A[465]), .Z(n3721) );
  AND U4285 ( .A(n3724), .B(n3725), .Z(n1189) );
  NAND U4286 ( .A(B[464]), .B(n3726), .Z(n3725) );
  NANDN U4287 ( .A(A[464]), .B(n1191), .Z(n3726) );
  NANDN U4288 ( .A(n1191), .B(A[464]), .Z(n3724) );
  AND U4289 ( .A(n3727), .B(n3728), .Z(n1191) );
  NAND U4290 ( .A(B[463]), .B(n3729), .Z(n3728) );
  NANDN U4291 ( .A(A[463]), .B(n1193), .Z(n3729) );
  NANDN U4292 ( .A(n1193), .B(A[463]), .Z(n3727) );
  AND U4293 ( .A(n3730), .B(n3731), .Z(n1193) );
  NAND U4294 ( .A(B[462]), .B(n3732), .Z(n3731) );
  NANDN U4295 ( .A(A[462]), .B(n1195), .Z(n3732) );
  NANDN U4296 ( .A(n1195), .B(A[462]), .Z(n3730) );
  AND U4297 ( .A(n3733), .B(n3734), .Z(n1195) );
  NAND U4298 ( .A(B[461]), .B(n3735), .Z(n3734) );
  NANDN U4299 ( .A(A[461]), .B(n1197), .Z(n3735) );
  NANDN U4300 ( .A(n1197), .B(A[461]), .Z(n3733) );
  AND U4301 ( .A(n3736), .B(n3737), .Z(n1197) );
  NAND U4302 ( .A(B[460]), .B(n3738), .Z(n3737) );
  NANDN U4303 ( .A(A[460]), .B(n1199), .Z(n3738) );
  NANDN U4304 ( .A(n1199), .B(A[460]), .Z(n3736) );
  AND U4305 ( .A(n3739), .B(n3740), .Z(n1199) );
  NAND U4306 ( .A(B[459]), .B(n3741), .Z(n3740) );
  NANDN U4307 ( .A(A[459]), .B(n1203), .Z(n3741) );
  NANDN U4308 ( .A(n1203), .B(A[459]), .Z(n3739) );
  AND U4309 ( .A(n3742), .B(n3743), .Z(n1203) );
  NAND U4310 ( .A(B[458]), .B(n3744), .Z(n3743) );
  NANDN U4311 ( .A(A[458]), .B(n1205), .Z(n3744) );
  NANDN U4312 ( .A(n1205), .B(A[458]), .Z(n3742) );
  AND U4313 ( .A(n3745), .B(n3746), .Z(n1205) );
  NAND U4314 ( .A(B[457]), .B(n3747), .Z(n3746) );
  NANDN U4315 ( .A(A[457]), .B(n1207), .Z(n3747) );
  NANDN U4316 ( .A(n1207), .B(A[457]), .Z(n3745) );
  AND U4317 ( .A(n3748), .B(n3749), .Z(n1207) );
  NAND U4318 ( .A(B[456]), .B(n3750), .Z(n3749) );
  NANDN U4319 ( .A(A[456]), .B(n1209), .Z(n3750) );
  NANDN U4320 ( .A(n1209), .B(A[456]), .Z(n3748) );
  AND U4321 ( .A(n3751), .B(n3752), .Z(n1209) );
  NAND U4322 ( .A(B[455]), .B(n3753), .Z(n3752) );
  NANDN U4323 ( .A(A[455]), .B(n1211), .Z(n3753) );
  NANDN U4324 ( .A(n1211), .B(A[455]), .Z(n3751) );
  AND U4325 ( .A(n3754), .B(n3755), .Z(n1211) );
  NAND U4326 ( .A(B[454]), .B(n3756), .Z(n3755) );
  NANDN U4327 ( .A(A[454]), .B(n1213), .Z(n3756) );
  NANDN U4328 ( .A(n1213), .B(A[454]), .Z(n3754) );
  AND U4329 ( .A(n3757), .B(n3758), .Z(n1213) );
  NAND U4330 ( .A(B[453]), .B(n3759), .Z(n3758) );
  NANDN U4331 ( .A(A[453]), .B(n1215), .Z(n3759) );
  NANDN U4332 ( .A(n1215), .B(A[453]), .Z(n3757) );
  AND U4333 ( .A(n3760), .B(n3761), .Z(n1215) );
  NAND U4334 ( .A(B[452]), .B(n3762), .Z(n3761) );
  NANDN U4335 ( .A(A[452]), .B(n1217), .Z(n3762) );
  NANDN U4336 ( .A(n1217), .B(A[452]), .Z(n3760) );
  AND U4337 ( .A(n3763), .B(n3764), .Z(n1217) );
  NAND U4338 ( .A(B[451]), .B(n3765), .Z(n3764) );
  NANDN U4339 ( .A(A[451]), .B(n1219), .Z(n3765) );
  NANDN U4340 ( .A(n1219), .B(A[451]), .Z(n3763) );
  AND U4341 ( .A(n3766), .B(n3767), .Z(n1219) );
  NAND U4342 ( .A(B[450]), .B(n3768), .Z(n3767) );
  NANDN U4343 ( .A(A[450]), .B(n1221), .Z(n3768) );
  NANDN U4344 ( .A(n1221), .B(A[450]), .Z(n3766) );
  AND U4345 ( .A(n3769), .B(n3770), .Z(n1221) );
  NAND U4346 ( .A(B[449]), .B(n3771), .Z(n3770) );
  NANDN U4347 ( .A(A[449]), .B(n1225), .Z(n3771) );
  NANDN U4348 ( .A(n1225), .B(A[449]), .Z(n3769) );
  AND U4349 ( .A(n3772), .B(n3773), .Z(n1225) );
  NAND U4350 ( .A(B[448]), .B(n3774), .Z(n3773) );
  NANDN U4351 ( .A(A[448]), .B(n1227), .Z(n3774) );
  NANDN U4352 ( .A(n1227), .B(A[448]), .Z(n3772) );
  AND U4353 ( .A(n3775), .B(n3776), .Z(n1227) );
  NAND U4354 ( .A(B[447]), .B(n3777), .Z(n3776) );
  NANDN U4355 ( .A(A[447]), .B(n1229), .Z(n3777) );
  NANDN U4356 ( .A(n1229), .B(A[447]), .Z(n3775) );
  AND U4357 ( .A(n3778), .B(n3779), .Z(n1229) );
  NAND U4358 ( .A(B[446]), .B(n3780), .Z(n3779) );
  NANDN U4359 ( .A(A[446]), .B(n1231), .Z(n3780) );
  NANDN U4360 ( .A(n1231), .B(A[446]), .Z(n3778) );
  AND U4361 ( .A(n3781), .B(n3782), .Z(n1231) );
  NAND U4362 ( .A(B[445]), .B(n3783), .Z(n3782) );
  NANDN U4363 ( .A(A[445]), .B(n1233), .Z(n3783) );
  NANDN U4364 ( .A(n1233), .B(A[445]), .Z(n3781) );
  AND U4365 ( .A(n3784), .B(n3785), .Z(n1233) );
  NAND U4366 ( .A(B[444]), .B(n3786), .Z(n3785) );
  NANDN U4367 ( .A(A[444]), .B(n1235), .Z(n3786) );
  NANDN U4368 ( .A(n1235), .B(A[444]), .Z(n3784) );
  AND U4369 ( .A(n3787), .B(n3788), .Z(n1235) );
  NAND U4370 ( .A(B[443]), .B(n3789), .Z(n3788) );
  NANDN U4371 ( .A(A[443]), .B(n1237), .Z(n3789) );
  NANDN U4372 ( .A(n1237), .B(A[443]), .Z(n3787) );
  AND U4373 ( .A(n3790), .B(n3791), .Z(n1237) );
  NAND U4374 ( .A(B[442]), .B(n3792), .Z(n3791) );
  NANDN U4375 ( .A(A[442]), .B(n1239), .Z(n3792) );
  NANDN U4376 ( .A(n1239), .B(A[442]), .Z(n3790) );
  AND U4377 ( .A(n3793), .B(n3794), .Z(n1239) );
  NAND U4378 ( .A(B[441]), .B(n3795), .Z(n3794) );
  NANDN U4379 ( .A(A[441]), .B(n1241), .Z(n3795) );
  NANDN U4380 ( .A(n1241), .B(A[441]), .Z(n3793) );
  AND U4381 ( .A(n3796), .B(n3797), .Z(n1241) );
  NAND U4382 ( .A(B[440]), .B(n3798), .Z(n3797) );
  NANDN U4383 ( .A(A[440]), .B(n1243), .Z(n3798) );
  NANDN U4384 ( .A(n1243), .B(A[440]), .Z(n3796) );
  AND U4385 ( .A(n3799), .B(n3800), .Z(n1243) );
  NAND U4386 ( .A(B[439]), .B(n3801), .Z(n3800) );
  NANDN U4387 ( .A(A[439]), .B(n1247), .Z(n3801) );
  NANDN U4388 ( .A(n1247), .B(A[439]), .Z(n3799) );
  AND U4389 ( .A(n3802), .B(n3803), .Z(n1247) );
  NAND U4390 ( .A(B[438]), .B(n3804), .Z(n3803) );
  NANDN U4391 ( .A(A[438]), .B(n1249), .Z(n3804) );
  NANDN U4392 ( .A(n1249), .B(A[438]), .Z(n3802) );
  AND U4393 ( .A(n3805), .B(n3806), .Z(n1249) );
  NAND U4394 ( .A(B[437]), .B(n3807), .Z(n3806) );
  NANDN U4395 ( .A(A[437]), .B(n1251), .Z(n3807) );
  NANDN U4396 ( .A(n1251), .B(A[437]), .Z(n3805) );
  AND U4397 ( .A(n3808), .B(n3809), .Z(n1251) );
  NAND U4398 ( .A(B[436]), .B(n3810), .Z(n3809) );
  NANDN U4399 ( .A(A[436]), .B(n1253), .Z(n3810) );
  NANDN U4400 ( .A(n1253), .B(A[436]), .Z(n3808) );
  AND U4401 ( .A(n3811), .B(n3812), .Z(n1253) );
  NAND U4402 ( .A(B[435]), .B(n3813), .Z(n3812) );
  NANDN U4403 ( .A(A[435]), .B(n1255), .Z(n3813) );
  NANDN U4404 ( .A(n1255), .B(A[435]), .Z(n3811) );
  AND U4405 ( .A(n3814), .B(n3815), .Z(n1255) );
  NAND U4406 ( .A(B[434]), .B(n3816), .Z(n3815) );
  NANDN U4407 ( .A(A[434]), .B(n1257), .Z(n3816) );
  NANDN U4408 ( .A(n1257), .B(A[434]), .Z(n3814) );
  AND U4409 ( .A(n3817), .B(n3818), .Z(n1257) );
  NAND U4410 ( .A(B[433]), .B(n3819), .Z(n3818) );
  NANDN U4411 ( .A(A[433]), .B(n1259), .Z(n3819) );
  NANDN U4412 ( .A(n1259), .B(A[433]), .Z(n3817) );
  AND U4413 ( .A(n3820), .B(n3821), .Z(n1259) );
  NAND U4414 ( .A(B[432]), .B(n3822), .Z(n3821) );
  NANDN U4415 ( .A(A[432]), .B(n1261), .Z(n3822) );
  NANDN U4416 ( .A(n1261), .B(A[432]), .Z(n3820) );
  AND U4417 ( .A(n3823), .B(n3824), .Z(n1261) );
  NAND U4418 ( .A(B[431]), .B(n3825), .Z(n3824) );
  NANDN U4419 ( .A(A[431]), .B(n1263), .Z(n3825) );
  NANDN U4420 ( .A(n1263), .B(A[431]), .Z(n3823) );
  AND U4421 ( .A(n3826), .B(n3827), .Z(n1263) );
  NAND U4422 ( .A(B[430]), .B(n3828), .Z(n3827) );
  NANDN U4423 ( .A(A[430]), .B(n1265), .Z(n3828) );
  NANDN U4424 ( .A(n1265), .B(A[430]), .Z(n3826) );
  AND U4425 ( .A(n3829), .B(n3830), .Z(n1265) );
  NAND U4426 ( .A(B[429]), .B(n3831), .Z(n3830) );
  NANDN U4427 ( .A(A[429]), .B(n1269), .Z(n3831) );
  NANDN U4428 ( .A(n1269), .B(A[429]), .Z(n3829) );
  AND U4429 ( .A(n3832), .B(n3833), .Z(n1269) );
  NAND U4430 ( .A(B[428]), .B(n3834), .Z(n3833) );
  NANDN U4431 ( .A(A[428]), .B(n1271), .Z(n3834) );
  NANDN U4432 ( .A(n1271), .B(A[428]), .Z(n3832) );
  AND U4433 ( .A(n3835), .B(n3836), .Z(n1271) );
  NAND U4434 ( .A(B[427]), .B(n3837), .Z(n3836) );
  NANDN U4435 ( .A(A[427]), .B(n1273), .Z(n3837) );
  NANDN U4436 ( .A(n1273), .B(A[427]), .Z(n3835) );
  AND U4437 ( .A(n3838), .B(n3839), .Z(n1273) );
  NAND U4438 ( .A(B[426]), .B(n3840), .Z(n3839) );
  NANDN U4439 ( .A(A[426]), .B(n1275), .Z(n3840) );
  NANDN U4440 ( .A(n1275), .B(A[426]), .Z(n3838) );
  AND U4441 ( .A(n3841), .B(n3842), .Z(n1275) );
  NAND U4442 ( .A(B[425]), .B(n3843), .Z(n3842) );
  NANDN U4443 ( .A(A[425]), .B(n1277), .Z(n3843) );
  NANDN U4444 ( .A(n1277), .B(A[425]), .Z(n3841) );
  AND U4445 ( .A(n3844), .B(n3845), .Z(n1277) );
  NAND U4446 ( .A(B[424]), .B(n3846), .Z(n3845) );
  NANDN U4447 ( .A(A[424]), .B(n1279), .Z(n3846) );
  NANDN U4448 ( .A(n1279), .B(A[424]), .Z(n3844) );
  AND U4449 ( .A(n3847), .B(n3848), .Z(n1279) );
  NAND U4450 ( .A(B[423]), .B(n3849), .Z(n3848) );
  NANDN U4451 ( .A(A[423]), .B(n1281), .Z(n3849) );
  NANDN U4452 ( .A(n1281), .B(A[423]), .Z(n3847) );
  AND U4453 ( .A(n3850), .B(n3851), .Z(n1281) );
  NAND U4454 ( .A(B[422]), .B(n3852), .Z(n3851) );
  NANDN U4455 ( .A(A[422]), .B(n1283), .Z(n3852) );
  NANDN U4456 ( .A(n1283), .B(A[422]), .Z(n3850) );
  AND U4457 ( .A(n3853), .B(n3854), .Z(n1283) );
  NAND U4458 ( .A(B[421]), .B(n3855), .Z(n3854) );
  NANDN U4459 ( .A(A[421]), .B(n1285), .Z(n3855) );
  NANDN U4460 ( .A(n1285), .B(A[421]), .Z(n3853) );
  AND U4461 ( .A(n3856), .B(n3857), .Z(n1285) );
  NAND U4462 ( .A(B[420]), .B(n3858), .Z(n3857) );
  NANDN U4463 ( .A(A[420]), .B(n1287), .Z(n3858) );
  NANDN U4464 ( .A(n1287), .B(A[420]), .Z(n3856) );
  AND U4465 ( .A(n3859), .B(n3860), .Z(n1287) );
  NAND U4466 ( .A(B[419]), .B(n3861), .Z(n3860) );
  NANDN U4467 ( .A(A[419]), .B(n1291), .Z(n3861) );
  NANDN U4468 ( .A(n1291), .B(A[419]), .Z(n3859) );
  AND U4469 ( .A(n3862), .B(n3863), .Z(n1291) );
  NAND U4470 ( .A(B[418]), .B(n3864), .Z(n3863) );
  NANDN U4471 ( .A(A[418]), .B(n1293), .Z(n3864) );
  NANDN U4472 ( .A(n1293), .B(A[418]), .Z(n3862) );
  AND U4473 ( .A(n3865), .B(n3866), .Z(n1293) );
  NAND U4474 ( .A(B[417]), .B(n3867), .Z(n3866) );
  NANDN U4475 ( .A(A[417]), .B(n1295), .Z(n3867) );
  NANDN U4476 ( .A(n1295), .B(A[417]), .Z(n3865) );
  AND U4477 ( .A(n3868), .B(n3869), .Z(n1295) );
  NAND U4478 ( .A(B[416]), .B(n3870), .Z(n3869) );
  NANDN U4479 ( .A(A[416]), .B(n1297), .Z(n3870) );
  NANDN U4480 ( .A(n1297), .B(A[416]), .Z(n3868) );
  AND U4481 ( .A(n3871), .B(n3872), .Z(n1297) );
  NAND U4482 ( .A(B[415]), .B(n3873), .Z(n3872) );
  NANDN U4483 ( .A(A[415]), .B(n1299), .Z(n3873) );
  NANDN U4484 ( .A(n1299), .B(A[415]), .Z(n3871) );
  AND U4485 ( .A(n3874), .B(n3875), .Z(n1299) );
  NAND U4486 ( .A(B[414]), .B(n3876), .Z(n3875) );
  NANDN U4487 ( .A(A[414]), .B(n1301), .Z(n3876) );
  NANDN U4488 ( .A(n1301), .B(A[414]), .Z(n3874) );
  AND U4489 ( .A(n3877), .B(n3878), .Z(n1301) );
  NAND U4490 ( .A(B[413]), .B(n3879), .Z(n3878) );
  NANDN U4491 ( .A(A[413]), .B(n1303), .Z(n3879) );
  NANDN U4492 ( .A(n1303), .B(A[413]), .Z(n3877) );
  AND U4493 ( .A(n3880), .B(n3881), .Z(n1303) );
  NAND U4494 ( .A(B[412]), .B(n3882), .Z(n3881) );
  NANDN U4495 ( .A(A[412]), .B(n1305), .Z(n3882) );
  NANDN U4496 ( .A(n1305), .B(A[412]), .Z(n3880) );
  AND U4497 ( .A(n3883), .B(n3884), .Z(n1305) );
  NAND U4498 ( .A(B[411]), .B(n3885), .Z(n3884) );
  NANDN U4499 ( .A(A[411]), .B(n1307), .Z(n3885) );
  NANDN U4500 ( .A(n1307), .B(A[411]), .Z(n3883) );
  AND U4501 ( .A(n3886), .B(n3887), .Z(n1307) );
  NAND U4502 ( .A(B[410]), .B(n3888), .Z(n3887) );
  NANDN U4503 ( .A(A[410]), .B(n1309), .Z(n3888) );
  NANDN U4504 ( .A(n1309), .B(A[410]), .Z(n3886) );
  AND U4505 ( .A(n3889), .B(n3890), .Z(n1309) );
  NAND U4506 ( .A(B[409]), .B(n3891), .Z(n3890) );
  NANDN U4507 ( .A(A[409]), .B(n1313), .Z(n3891) );
  NANDN U4508 ( .A(n1313), .B(A[409]), .Z(n3889) );
  AND U4509 ( .A(n3892), .B(n3893), .Z(n1313) );
  NAND U4510 ( .A(B[408]), .B(n3894), .Z(n3893) );
  NANDN U4511 ( .A(A[408]), .B(n1315), .Z(n3894) );
  NANDN U4512 ( .A(n1315), .B(A[408]), .Z(n3892) );
  AND U4513 ( .A(n3895), .B(n3896), .Z(n1315) );
  NAND U4514 ( .A(B[407]), .B(n3897), .Z(n3896) );
  NANDN U4515 ( .A(A[407]), .B(n1317), .Z(n3897) );
  NANDN U4516 ( .A(n1317), .B(A[407]), .Z(n3895) );
  AND U4517 ( .A(n3898), .B(n3899), .Z(n1317) );
  NAND U4518 ( .A(B[406]), .B(n3900), .Z(n3899) );
  NANDN U4519 ( .A(A[406]), .B(n1319), .Z(n3900) );
  NANDN U4520 ( .A(n1319), .B(A[406]), .Z(n3898) );
  AND U4521 ( .A(n3901), .B(n3902), .Z(n1319) );
  NAND U4522 ( .A(B[405]), .B(n3903), .Z(n3902) );
  NANDN U4523 ( .A(A[405]), .B(n1321), .Z(n3903) );
  NANDN U4524 ( .A(n1321), .B(A[405]), .Z(n3901) );
  AND U4525 ( .A(n3904), .B(n3905), .Z(n1321) );
  NAND U4526 ( .A(B[404]), .B(n3906), .Z(n3905) );
  NANDN U4527 ( .A(A[404]), .B(n1323), .Z(n3906) );
  NANDN U4528 ( .A(n1323), .B(A[404]), .Z(n3904) );
  AND U4529 ( .A(n3907), .B(n3908), .Z(n1323) );
  NAND U4530 ( .A(B[403]), .B(n3909), .Z(n3908) );
  NANDN U4531 ( .A(A[403]), .B(n1325), .Z(n3909) );
  NANDN U4532 ( .A(n1325), .B(A[403]), .Z(n3907) );
  AND U4533 ( .A(n3910), .B(n3911), .Z(n1325) );
  NAND U4534 ( .A(B[402]), .B(n3912), .Z(n3911) );
  NANDN U4535 ( .A(A[402]), .B(n1327), .Z(n3912) );
  NANDN U4536 ( .A(n1327), .B(A[402]), .Z(n3910) );
  AND U4537 ( .A(n3913), .B(n3914), .Z(n1327) );
  NAND U4538 ( .A(B[401]), .B(n3915), .Z(n3914) );
  NANDN U4539 ( .A(A[401]), .B(n1329), .Z(n3915) );
  NANDN U4540 ( .A(n1329), .B(A[401]), .Z(n3913) );
  AND U4541 ( .A(n3916), .B(n3917), .Z(n1329) );
  NAND U4542 ( .A(B[400]), .B(n3918), .Z(n3917) );
  NANDN U4543 ( .A(A[400]), .B(n1331), .Z(n3918) );
  NANDN U4544 ( .A(n1331), .B(A[400]), .Z(n3916) );
  AND U4545 ( .A(n3919), .B(n3920), .Z(n1331) );
  NAND U4546 ( .A(B[399]), .B(n3921), .Z(n3920) );
  NANDN U4547 ( .A(A[399]), .B(n1337), .Z(n3921) );
  NANDN U4548 ( .A(n1337), .B(A[399]), .Z(n3919) );
  AND U4549 ( .A(n3922), .B(n3923), .Z(n1337) );
  NAND U4550 ( .A(B[398]), .B(n3924), .Z(n3923) );
  NANDN U4551 ( .A(A[398]), .B(n1339), .Z(n3924) );
  NANDN U4552 ( .A(n1339), .B(A[398]), .Z(n3922) );
  AND U4553 ( .A(n3925), .B(n3926), .Z(n1339) );
  NAND U4554 ( .A(B[397]), .B(n3927), .Z(n3926) );
  NANDN U4555 ( .A(A[397]), .B(n1341), .Z(n3927) );
  NANDN U4556 ( .A(n1341), .B(A[397]), .Z(n3925) );
  AND U4557 ( .A(n3928), .B(n3929), .Z(n1341) );
  NAND U4558 ( .A(B[396]), .B(n3930), .Z(n3929) );
  NANDN U4559 ( .A(A[396]), .B(n1343), .Z(n3930) );
  NANDN U4560 ( .A(n1343), .B(A[396]), .Z(n3928) );
  AND U4561 ( .A(n3931), .B(n3932), .Z(n1343) );
  NAND U4562 ( .A(B[395]), .B(n3933), .Z(n3932) );
  NANDN U4563 ( .A(A[395]), .B(n1345), .Z(n3933) );
  NANDN U4564 ( .A(n1345), .B(A[395]), .Z(n3931) );
  AND U4565 ( .A(n3934), .B(n3935), .Z(n1345) );
  NAND U4566 ( .A(B[394]), .B(n3936), .Z(n3935) );
  NANDN U4567 ( .A(A[394]), .B(n1347), .Z(n3936) );
  NANDN U4568 ( .A(n1347), .B(A[394]), .Z(n3934) );
  AND U4569 ( .A(n3937), .B(n3938), .Z(n1347) );
  NAND U4570 ( .A(B[393]), .B(n3939), .Z(n3938) );
  NANDN U4571 ( .A(A[393]), .B(n1349), .Z(n3939) );
  NANDN U4572 ( .A(n1349), .B(A[393]), .Z(n3937) );
  AND U4573 ( .A(n3940), .B(n3941), .Z(n1349) );
  NAND U4574 ( .A(B[392]), .B(n3942), .Z(n3941) );
  NANDN U4575 ( .A(A[392]), .B(n1351), .Z(n3942) );
  NANDN U4576 ( .A(n1351), .B(A[392]), .Z(n3940) );
  AND U4577 ( .A(n3943), .B(n3944), .Z(n1351) );
  NAND U4578 ( .A(B[391]), .B(n3945), .Z(n3944) );
  NANDN U4579 ( .A(A[391]), .B(n1353), .Z(n3945) );
  NANDN U4580 ( .A(n1353), .B(A[391]), .Z(n3943) );
  AND U4581 ( .A(n3946), .B(n3947), .Z(n1353) );
  NAND U4582 ( .A(B[390]), .B(n3948), .Z(n3947) );
  NANDN U4583 ( .A(A[390]), .B(n1355), .Z(n3948) );
  NANDN U4584 ( .A(n1355), .B(A[390]), .Z(n3946) );
  AND U4585 ( .A(n3949), .B(n3950), .Z(n1355) );
  NAND U4586 ( .A(B[389]), .B(n3951), .Z(n3950) );
  NANDN U4587 ( .A(A[389]), .B(n1359), .Z(n3951) );
  NANDN U4588 ( .A(n1359), .B(A[389]), .Z(n3949) );
  AND U4589 ( .A(n3952), .B(n3953), .Z(n1359) );
  NAND U4590 ( .A(B[388]), .B(n3954), .Z(n3953) );
  NANDN U4591 ( .A(A[388]), .B(n1361), .Z(n3954) );
  NANDN U4592 ( .A(n1361), .B(A[388]), .Z(n3952) );
  AND U4593 ( .A(n3955), .B(n3956), .Z(n1361) );
  NAND U4594 ( .A(B[387]), .B(n3957), .Z(n3956) );
  NANDN U4595 ( .A(A[387]), .B(n1363), .Z(n3957) );
  NANDN U4596 ( .A(n1363), .B(A[387]), .Z(n3955) );
  AND U4597 ( .A(n3958), .B(n3959), .Z(n1363) );
  NAND U4598 ( .A(B[386]), .B(n3960), .Z(n3959) );
  NANDN U4599 ( .A(A[386]), .B(n1365), .Z(n3960) );
  NANDN U4600 ( .A(n1365), .B(A[386]), .Z(n3958) );
  AND U4601 ( .A(n3961), .B(n3962), .Z(n1365) );
  NAND U4602 ( .A(B[385]), .B(n3963), .Z(n3962) );
  NANDN U4603 ( .A(A[385]), .B(n1367), .Z(n3963) );
  NANDN U4604 ( .A(n1367), .B(A[385]), .Z(n3961) );
  AND U4605 ( .A(n3964), .B(n3965), .Z(n1367) );
  NAND U4606 ( .A(B[384]), .B(n3966), .Z(n3965) );
  NANDN U4607 ( .A(A[384]), .B(n1369), .Z(n3966) );
  NANDN U4608 ( .A(n1369), .B(A[384]), .Z(n3964) );
  AND U4609 ( .A(n3967), .B(n3968), .Z(n1369) );
  NAND U4610 ( .A(B[383]), .B(n3969), .Z(n3968) );
  NANDN U4611 ( .A(A[383]), .B(n1371), .Z(n3969) );
  NANDN U4612 ( .A(n1371), .B(A[383]), .Z(n3967) );
  AND U4613 ( .A(n3970), .B(n3971), .Z(n1371) );
  NAND U4614 ( .A(B[382]), .B(n3972), .Z(n3971) );
  NANDN U4615 ( .A(A[382]), .B(n1373), .Z(n3972) );
  NANDN U4616 ( .A(n1373), .B(A[382]), .Z(n3970) );
  AND U4617 ( .A(n3973), .B(n3974), .Z(n1373) );
  NAND U4618 ( .A(B[381]), .B(n3975), .Z(n3974) );
  NANDN U4619 ( .A(A[381]), .B(n1375), .Z(n3975) );
  NANDN U4620 ( .A(n1375), .B(A[381]), .Z(n3973) );
  AND U4621 ( .A(n3976), .B(n3977), .Z(n1375) );
  NAND U4622 ( .A(B[380]), .B(n3978), .Z(n3977) );
  NANDN U4623 ( .A(A[380]), .B(n1377), .Z(n3978) );
  NANDN U4624 ( .A(n1377), .B(A[380]), .Z(n3976) );
  AND U4625 ( .A(n3979), .B(n3980), .Z(n1377) );
  NAND U4626 ( .A(B[379]), .B(n3981), .Z(n3980) );
  NANDN U4627 ( .A(A[379]), .B(n1381), .Z(n3981) );
  NANDN U4628 ( .A(n1381), .B(A[379]), .Z(n3979) );
  AND U4629 ( .A(n3982), .B(n3983), .Z(n1381) );
  NAND U4630 ( .A(B[378]), .B(n3984), .Z(n3983) );
  NANDN U4631 ( .A(A[378]), .B(n1383), .Z(n3984) );
  NANDN U4632 ( .A(n1383), .B(A[378]), .Z(n3982) );
  AND U4633 ( .A(n3985), .B(n3986), .Z(n1383) );
  NAND U4634 ( .A(B[377]), .B(n3987), .Z(n3986) );
  NANDN U4635 ( .A(A[377]), .B(n1385), .Z(n3987) );
  NANDN U4636 ( .A(n1385), .B(A[377]), .Z(n3985) );
  AND U4637 ( .A(n3988), .B(n3989), .Z(n1385) );
  NAND U4638 ( .A(B[376]), .B(n3990), .Z(n3989) );
  NANDN U4639 ( .A(A[376]), .B(n1387), .Z(n3990) );
  NANDN U4640 ( .A(n1387), .B(A[376]), .Z(n3988) );
  AND U4641 ( .A(n3991), .B(n3992), .Z(n1387) );
  NAND U4642 ( .A(B[375]), .B(n3993), .Z(n3992) );
  NANDN U4643 ( .A(A[375]), .B(n1389), .Z(n3993) );
  NANDN U4644 ( .A(n1389), .B(A[375]), .Z(n3991) );
  AND U4645 ( .A(n3994), .B(n3995), .Z(n1389) );
  NAND U4646 ( .A(B[374]), .B(n3996), .Z(n3995) );
  NANDN U4647 ( .A(A[374]), .B(n1391), .Z(n3996) );
  NANDN U4648 ( .A(n1391), .B(A[374]), .Z(n3994) );
  AND U4649 ( .A(n3997), .B(n3998), .Z(n1391) );
  NAND U4650 ( .A(B[373]), .B(n3999), .Z(n3998) );
  NANDN U4651 ( .A(A[373]), .B(n1393), .Z(n3999) );
  NANDN U4652 ( .A(n1393), .B(A[373]), .Z(n3997) );
  AND U4653 ( .A(n4000), .B(n4001), .Z(n1393) );
  NAND U4654 ( .A(B[372]), .B(n4002), .Z(n4001) );
  NANDN U4655 ( .A(A[372]), .B(n1395), .Z(n4002) );
  NANDN U4656 ( .A(n1395), .B(A[372]), .Z(n4000) );
  AND U4657 ( .A(n4003), .B(n4004), .Z(n1395) );
  NAND U4658 ( .A(B[371]), .B(n4005), .Z(n4004) );
  NANDN U4659 ( .A(A[371]), .B(n1397), .Z(n4005) );
  NANDN U4660 ( .A(n1397), .B(A[371]), .Z(n4003) );
  AND U4661 ( .A(n4006), .B(n4007), .Z(n1397) );
  NAND U4662 ( .A(B[370]), .B(n4008), .Z(n4007) );
  NANDN U4663 ( .A(A[370]), .B(n1399), .Z(n4008) );
  NANDN U4664 ( .A(n1399), .B(A[370]), .Z(n4006) );
  AND U4665 ( .A(n4009), .B(n4010), .Z(n1399) );
  NAND U4666 ( .A(B[369]), .B(n4011), .Z(n4010) );
  NANDN U4667 ( .A(A[369]), .B(n1403), .Z(n4011) );
  NANDN U4668 ( .A(n1403), .B(A[369]), .Z(n4009) );
  AND U4669 ( .A(n4012), .B(n4013), .Z(n1403) );
  NAND U4670 ( .A(B[368]), .B(n4014), .Z(n4013) );
  NANDN U4671 ( .A(A[368]), .B(n1405), .Z(n4014) );
  NANDN U4672 ( .A(n1405), .B(A[368]), .Z(n4012) );
  AND U4673 ( .A(n4015), .B(n4016), .Z(n1405) );
  NAND U4674 ( .A(B[367]), .B(n4017), .Z(n4016) );
  NANDN U4675 ( .A(A[367]), .B(n1407), .Z(n4017) );
  NANDN U4676 ( .A(n1407), .B(A[367]), .Z(n4015) );
  AND U4677 ( .A(n4018), .B(n4019), .Z(n1407) );
  NAND U4678 ( .A(B[366]), .B(n4020), .Z(n4019) );
  NANDN U4679 ( .A(A[366]), .B(n1409), .Z(n4020) );
  NANDN U4680 ( .A(n1409), .B(A[366]), .Z(n4018) );
  AND U4681 ( .A(n4021), .B(n4022), .Z(n1409) );
  NAND U4682 ( .A(B[365]), .B(n4023), .Z(n4022) );
  NANDN U4683 ( .A(A[365]), .B(n1411), .Z(n4023) );
  NANDN U4684 ( .A(n1411), .B(A[365]), .Z(n4021) );
  AND U4685 ( .A(n4024), .B(n4025), .Z(n1411) );
  NAND U4686 ( .A(B[364]), .B(n4026), .Z(n4025) );
  NANDN U4687 ( .A(A[364]), .B(n1413), .Z(n4026) );
  NANDN U4688 ( .A(n1413), .B(A[364]), .Z(n4024) );
  AND U4689 ( .A(n4027), .B(n4028), .Z(n1413) );
  NAND U4690 ( .A(B[363]), .B(n4029), .Z(n4028) );
  NANDN U4691 ( .A(A[363]), .B(n1415), .Z(n4029) );
  NANDN U4692 ( .A(n1415), .B(A[363]), .Z(n4027) );
  AND U4693 ( .A(n4030), .B(n4031), .Z(n1415) );
  NAND U4694 ( .A(B[362]), .B(n4032), .Z(n4031) );
  NANDN U4695 ( .A(A[362]), .B(n1417), .Z(n4032) );
  NANDN U4696 ( .A(n1417), .B(A[362]), .Z(n4030) );
  AND U4697 ( .A(n4033), .B(n4034), .Z(n1417) );
  NAND U4698 ( .A(B[361]), .B(n4035), .Z(n4034) );
  NANDN U4699 ( .A(A[361]), .B(n1419), .Z(n4035) );
  NANDN U4700 ( .A(n1419), .B(A[361]), .Z(n4033) );
  AND U4701 ( .A(n4036), .B(n4037), .Z(n1419) );
  NAND U4702 ( .A(B[360]), .B(n4038), .Z(n4037) );
  NANDN U4703 ( .A(A[360]), .B(n1421), .Z(n4038) );
  NANDN U4704 ( .A(n1421), .B(A[360]), .Z(n4036) );
  AND U4705 ( .A(n4039), .B(n4040), .Z(n1421) );
  NAND U4706 ( .A(B[359]), .B(n4041), .Z(n4040) );
  NANDN U4707 ( .A(A[359]), .B(n1425), .Z(n4041) );
  NANDN U4708 ( .A(n1425), .B(A[359]), .Z(n4039) );
  AND U4709 ( .A(n4042), .B(n4043), .Z(n1425) );
  NAND U4710 ( .A(B[358]), .B(n4044), .Z(n4043) );
  NANDN U4711 ( .A(A[358]), .B(n1427), .Z(n4044) );
  NANDN U4712 ( .A(n1427), .B(A[358]), .Z(n4042) );
  AND U4713 ( .A(n4045), .B(n4046), .Z(n1427) );
  NAND U4714 ( .A(B[357]), .B(n4047), .Z(n4046) );
  NANDN U4715 ( .A(A[357]), .B(n1429), .Z(n4047) );
  NANDN U4716 ( .A(n1429), .B(A[357]), .Z(n4045) );
  AND U4717 ( .A(n4048), .B(n4049), .Z(n1429) );
  NAND U4718 ( .A(B[356]), .B(n4050), .Z(n4049) );
  NANDN U4719 ( .A(A[356]), .B(n1431), .Z(n4050) );
  NANDN U4720 ( .A(n1431), .B(A[356]), .Z(n4048) );
  AND U4721 ( .A(n4051), .B(n4052), .Z(n1431) );
  NAND U4722 ( .A(B[355]), .B(n4053), .Z(n4052) );
  NANDN U4723 ( .A(A[355]), .B(n1433), .Z(n4053) );
  NANDN U4724 ( .A(n1433), .B(A[355]), .Z(n4051) );
  AND U4725 ( .A(n4054), .B(n4055), .Z(n1433) );
  NAND U4726 ( .A(B[354]), .B(n4056), .Z(n4055) );
  NANDN U4727 ( .A(A[354]), .B(n1435), .Z(n4056) );
  NANDN U4728 ( .A(n1435), .B(A[354]), .Z(n4054) );
  AND U4729 ( .A(n4057), .B(n4058), .Z(n1435) );
  NAND U4730 ( .A(B[353]), .B(n4059), .Z(n4058) );
  NANDN U4731 ( .A(A[353]), .B(n1437), .Z(n4059) );
  NANDN U4732 ( .A(n1437), .B(A[353]), .Z(n4057) );
  AND U4733 ( .A(n4060), .B(n4061), .Z(n1437) );
  NAND U4734 ( .A(B[352]), .B(n4062), .Z(n4061) );
  NANDN U4735 ( .A(A[352]), .B(n1439), .Z(n4062) );
  NANDN U4736 ( .A(n1439), .B(A[352]), .Z(n4060) );
  AND U4737 ( .A(n4063), .B(n4064), .Z(n1439) );
  NAND U4738 ( .A(B[351]), .B(n4065), .Z(n4064) );
  NANDN U4739 ( .A(A[351]), .B(n1441), .Z(n4065) );
  NANDN U4740 ( .A(n1441), .B(A[351]), .Z(n4063) );
  AND U4741 ( .A(n4066), .B(n4067), .Z(n1441) );
  NAND U4742 ( .A(B[350]), .B(n4068), .Z(n4067) );
  NANDN U4743 ( .A(A[350]), .B(n1443), .Z(n4068) );
  NANDN U4744 ( .A(n1443), .B(A[350]), .Z(n4066) );
  AND U4745 ( .A(n4069), .B(n4070), .Z(n1443) );
  NAND U4746 ( .A(B[349]), .B(n4071), .Z(n4070) );
  NANDN U4747 ( .A(A[349]), .B(n1447), .Z(n4071) );
  NANDN U4748 ( .A(n1447), .B(A[349]), .Z(n4069) );
  AND U4749 ( .A(n4072), .B(n4073), .Z(n1447) );
  NAND U4750 ( .A(B[348]), .B(n4074), .Z(n4073) );
  NANDN U4751 ( .A(A[348]), .B(n1449), .Z(n4074) );
  NANDN U4752 ( .A(n1449), .B(A[348]), .Z(n4072) );
  AND U4753 ( .A(n4075), .B(n4076), .Z(n1449) );
  NAND U4754 ( .A(B[347]), .B(n4077), .Z(n4076) );
  NANDN U4755 ( .A(A[347]), .B(n1451), .Z(n4077) );
  NANDN U4756 ( .A(n1451), .B(A[347]), .Z(n4075) );
  AND U4757 ( .A(n4078), .B(n4079), .Z(n1451) );
  NAND U4758 ( .A(B[346]), .B(n4080), .Z(n4079) );
  NANDN U4759 ( .A(A[346]), .B(n1453), .Z(n4080) );
  NANDN U4760 ( .A(n1453), .B(A[346]), .Z(n4078) );
  AND U4761 ( .A(n4081), .B(n4082), .Z(n1453) );
  NAND U4762 ( .A(B[345]), .B(n4083), .Z(n4082) );
  NANDN U4763 ( .A(A[345]), .B(n1455), .Z(n4083) );
  NANDN U4764 ( .A(n1455), .B(A[345]), .Z(n4081) );
  AND U4765 ( .A(n4084), .B(n4085), .Z(n1455) );
  NAND U4766 ( .A(B[344]), .B(n4086), .Z(n4085) );
  NANDN U4767 ( .A(A[344]), .B(n1457), .Z(n4086) );
  NANDN U4768 ( .A(n1457), .B(A[344]), .Z(n4084) );
  AND U4769 ( .A(n4087), .B(n4088), .Z(n1457) );
  NAND U4770 ( .A(B[343]), .B(n4089), .Z(n4088) );
  NANDN U4771 ( .A(A[343]), .B(n1459), .Z(n4089) );
  NANDN U4772 ( .A(n1459), .B(A[343]), .Z(n4087) );
  AND U4773 ( .A(n4090), .B(n4091), .Z(n1459) );
  NAND U4774 ( .A(B[342]), .B(n4092), .Z(n4091) );
  NANDN U4775 ( .A(A[342]), .B(n1461), .Z(n4092) );
  NANDN U4776 ( .A(n1461), .B(A[342]), .Z(n4090) );
  AND U4777 ( .A(n4093), .B(n4094), .Z(n1461) );
  NAND U4778 ( .A(B[341]), .B(n4095), .Z(n4094) );
  NANDN U4779 ( .A(A[341]), .B(n1463), .Z(n4095) );
  NANDN U4780 ( .A(n1463), .B(A[341]), .Z(n4093) );
  AND U4781 ( .A(n4096), .B(n4097), .Z(n1463) );
  NAND U4782 ( .A(B[340]), .B(n4098), .Z(n4097) );
  NANDN U4783 ( .A(A[340]), .B(n1465), .Z(n4098) );
  NANDN U4784 ( .A(n1465), .B(A[340]), .Z(n4096) );
  AND U4785 ( .A(n4099), .B(n4100), .Z(n1465) );
  NAND U4786 ( .A(B[339]), .B(n4101), .Z(n4100) );
  NANDN U4787 ( .A(A[339]), .B(n1469), .Z(n4101) );
  NANDN U4788 ( .A(n1469), .B(A[339]), .Z(n4099) );
  AND U4789 ( .A(n4102), .B(n4103), .Z(n1469) );
  NAND U4790 ( .A(B[338]), .B(n4104), .Z(n4103) );
  NANDN U4791 ( .A(A[338]), .B(n1471), .Z(n4104) );
  NANDN U4792 ( .A(n1471), .B(A[338]), .Z(n4102) );
  AND U4793 ( .A(n4105), .B(n4106), .Z(n1471) );
  NAND U4794 ( .A(B[337]), .B(n4107), .Z(n4106) );
  NANDN U4795 ( .A(A[337]), .B(n1473), .Z(n4107) );
  NANDN U4796 ( .A(n1473), .B(A[337]), .Z(n4105) );
  AND U4797 ( .A(n4108), .B(n4109), .Z(n1473) );
  NAND U4798 ( .A(B[336]), .B(n4110), .Z(n4109) );
  NANDN U4799 ( .A(A[336]), .B(n1475), .Z(n4110) );
  NANDN U4800 ( .A(n1475), .B(A[336]), .Z(n4108) );
  AND U4801 ( .A(n4111), .B(n4112), .Z(n1475) );
  NAND U4802 ( .A(B[335]), .B(n4113), .Z(n4112) );
  NANDN U4803 ( .A(A[335]), .B(n1477), .Z(n4113) );
  NANDN U4804 ( .A(n1477), .B(A[335]), .Z(n4111) );
  AND U4805 ( .A(n4114), .B(n4115), .Z(n1477) );
  NAND U4806 ( .A(B[334]), .B(n4116), .Z(n4115) );
  NANDN U4807 ( .A(A[334]), .B(n1479), .Z(n4116) );
  NANDN U4808 ( .A(n1479), .B(A[334]), .Z(n4114) );
  AND U4809 ( .A(n4117), .B(n4118), .Z(n1479) );
  NAND U4810 ( .A(B[333]), .B(n4119), .Z(n4118) );
  NANDN U4811 ( .A(A[333]), .B(n1481), .Z(n4119) );
  NANDN U4812 ( .A(n1481), .B(A[333]), .Z(n4117) );
  AND U4813 ( .A(n4120), .B(n4121), .Z(n1481) );
  NAND U4814 ( .A(B[332]), .B(n4122), .Z(n4121) );
  NANDN U4815 ( .A(A[332]), .B(n1483), .Z(n4122) );
  NANDN U4816 ( .A(n1483), .B(A[332]), .Z(n4120) );
  AND U4817 ( .A(n4123), .B(n4124), .Z(n1483) );
  NAND U4818 ( .A(B[331]), .B(n4125), .Z(n4124) );
  NANDN U4819 ( .A(A[331]), .B(n1485), .Z(n4125) );
  NANDN U4820 ( .A(n1485), .B(A[331]), .Z(n4123) );
  AND U4821 ( .A(n4126), .B(n4127), .Z(n1485) );
  NAND U4822 ( .A(B[330]), .B(n4128), .Z(n4127) );
  NANDN U4823 ( .A(A[330]), .B(n1487), .Z(n4128) );
  NANDN U4824 ( .A(n1487), .B(A[330]), .Z(n4126) );
  AND U4825 ( .A(n4129), .B(n4130), .Z(n1487) );
  NAND U4826 ( .A(B[329]), .B(n4131), .Z(n4130) );
  NANDN U4827 ( .A(A[329]), .B(n1491), .Z(n4131) );
  NANDN U4828 ( .A(n1491), .B(A[329]), .Z(n4129) );
  AND U4829 ( .A(n4132), .B(n4133), .Z(n1491) );
  NAND U4830 ( .A(B[328]), .B(n4134), .Z(n4133) );
  NANDN U4831 ( .A(A[328]), .B(n1493), .Z(n4134) );
  NANDN U4832 ( .A(n1493), .B(A[328]), .Z(n4132) );
  AND U4833 ( .A(n4135), .B(n4136), .Z(n1493) );
  NAND U4834 ( .A(B[327]), .B(n4137), .Z(n4136) );
  NANDN U4835 ( .A(A[327]), .B(n1495), .Z(n4137) );
  NANDN U4836 ( .A(n1495), .B(A[327]), .Z(n4135) );
  AND U4837 ( .A(n4138), .B(n4139), .Z(n1495) );
  NAND U4838 ( .A(B[326]), .B(n4140), .Z(n4139) );
  NANDN U4839 ( .A(A[326]), .B(n1497), .Z(n4140) );
  NANDN U4840 ( .A(n1497), .B(A[326]), .Z(n4138) );
  AND U4841 ( .A(n4141), .B(n4142), .Z(n1497) );
  NAND U4842 ( .A(B[325]), .B(n4143), .Z(n4142) );
  NANDN U4843 ( .A(A[325]), .B(n1499), .Z(n4143) );
  NANDN U4844 ( .A(n1499), .B(A[325]), .Z(n4141) );
  AND U4845 ( .A(n4144), .B(n4145), .Z(n1499) );
  NAND U4846 ( .A(B[324]), .B(n4146), .Z(n4145) );
  NANDN U4847 ( .A(A[324]), .B(n1501), .Z(n4146) );
  NANDN U4848 ( .A(n1501), .B(A[324]), .Z(n4144) );
  AND U4849 ( .A(n4147), .B(n4148), .Z(n1501) );
  NAND U4850 ( .A(B[323]), .B(n4149), .Z(n4148) );
  NANDN U4851 ( .A(A[323]), .B(n1503), .Z(n4149) );
  NANDN U4852 ( .A(n1503), .B(A[323]), .Z(n4147) );
  AND U4853 ( .A(n4150), .B(n4151), .Z(n1503) );
  NAND U4854 ( .A(B[322]), .B(n4152), .Z(n4151) );
  NANDN U4855 ( .A(A[322]), .B(n1505), .Z(n4152) );
  NANDN U4856 ( .A(n1505), .B(A[322]), .Z(n4150) );
  AND U4857 ( .A(n4153), .B(n4154), .Z(n1505) );
  NAND U4858 ( .A(B[321]), .B(n4155), .Z(n4154) );
  NANDN U4859 ( .A(A[321]), .B(n1507), .Z(n4155) );
  NANDN U4860 ( .A(n1507), .B(A[321]), .Z(n4153) );
  AND U4861 ( .A(n4156), .B(n4157), .Z(n1507) );
  NAND U4862 ( .A(B[320]), .B(n4158), .Z(n4157) );
  NANDN U4863 ( .A(A[320]), .B(n1509), .Z(n4158) );
  NANDN U4864 ( .A(n1509), .B(A[320]), .Z(n4156) );
  AND U4865 ( .A(n4159), .B(n4160), .Z(n1509) );
  NAND U4866 ( .A(B[319]), .B(n4161), .Z(n4160) );
  NANDN U4867 ( .A(A[319]), .B(n1513), .Z(n4161) );
  NANDN U4868 ( .A(n1513), .B(A[319]), .Z(n4159) );
  AND U4869 ( .A(n4162), .B(n4163), .Z(n1513) );
  NAND U4870 ( .A(B[318]), .B(n4164), .Z(n4163) );
  NANDN U4871 ( .A(A[318]), .B(n1515), .Z(n4164) );
  NANDN U4872 ( .A(n1515), .B(A[318]), .Z(n4162) );
  AND U4873 ( .A(n4165), .B(n4166), .Z(n1515) );
  NAND U4874 ( .A(B[317]), .B(n4167), .Z(n4166) );
  NANDN U4875 ( .A(A[317]), .B(n1517), .Z(n4167) );
  NANDN U4876 ( .A(n1517), .B(A[317]), .Z(n4165) );
  AND U4877 ( .A(n4168), .B(n4169), .Z(n1517) );
  NAND U4878 ( .A(B[316]), .B(n4170), .Z(n4169) );
  NANDN U4879 ( .A(A[316]), .B(n1519), .Z(n4170) );
  NANDN U4880 ( .A(n1519), .B(A[316]), .Z(n4168) );
  AND U4881 ( .A(n4171), .B(n4172), .Z(n1519) );
  NAND U4882 ( .A(B[315]), .B(n4173), .Z(n4172) );
  NANDN U4883 ( .A(A[315]), .B(n1521), .Z(n4173) );
  NANDN U4884 ( .A(n1521), .B(A[315]), .Z(n4171) );
  AND U4885 ( .A(n4174), .B(n4175), .Z(n1521) );
  NAND U4886 ( .A(B[314]), .B(n4176), .Z(n4175) );
  NANDN U4887 ( .A(A[314]), .B(n1523), .Z(n4176) );
  NANDN U4888 ( .A(n1523), .B(A[314]), .Z(n4174) );
  AND U4889 ( .A(n4177), .B(n4178), .Z(n1523) );
  NAND U4890 ( .A(B[313]), .B(n4179), .Z(n4178) );
  NANDN U4891 ( .A(A[313]), .B(n1525), .Z(n4179) );
  NANDN U4892 ( .A(n1525), .B(A[313]), .Z(n4177) );
  AND U4893 ( .A(n4180), .B(n4181), .Z(n1525) );
  NAND U4894 ( .A(B[312]), .B(n4182), .Z(n4181) );
  NANDN U4895 ( .A(A[312]), .B(n1527), .Z(n4182) );
  NANDN U4896 ( .A(n1527), .B(A[312]), .Z(n4180) );
  AND U4897 ( .A(n4183), .B(n4184), .Z(n1527) );
  NAND U4898 ( .A(B[311]), .B(n4185), .Z(n4184) );
  NANDN U4899 ( .A(A[311]), .B(n1529), .Z(n4185) );
  NANDN U4900 ( .A(n1529), .B(A[311]), .Z(n4183) );
  AND U4901 ( .A(n4186), .B(n4187), .Z(n1529) );
  NAND U4902 ( .A(B[310]), .B(n4188), .Z(n4187) );
  NANDN U4903 ( .A(A[310]), .B(n1531), .Z(n4188) );
  NANDN U4904 ( .A(n1531), .B(A[310]), .Z(n4186) );
  AND U4905 ( .A(n4189), .B(n4190), .Z(n1531) );
  NAND U4906 ( .A(B[309]), .B(n4191), .Z(n4190) );
  NANDN U4907 ( .A(A[309]), .B(n1535), .Z(n4191) );
  NANDN U4908 ( .A(n1535), .B(A[309]), .Z(n4189) );
  AND U4909 ( .A(n4192), .B(n4193), .Z(n1535) );
  NAND U4910 ( .A(B[308]), .B(n4194), .Z(n4193) );
  NANDN U4911 ( .A(A[308]), .B(n1537), .Z(n4194) );
  NANDN U4912 ( .A(n1537), .B(A[308]), .Z(n4192) );
  AND U4913 ( .A(n4195), .B(n4196), .Z(n1537) );
  NAND U4914 ( .A(B[307]), .B(n4197), .Z(n4196) );
  NANDN U4915 ( .A(A[307]), .B(n1539), .Z(n4197) );
  NANDN U4916 ( .A(n1539), .B(A[307]), .Z(n4195) );
  AND U4917 ( .A(n4198), .B(n4199), .Z(n1539) );
  NAND U4918 ( .A(B[306]), .B(n4200), .Z(n4199) );
  NANDN U4919 ( .A(A[306]), .B(n1541), .Z(n4200) );
  NANDN U4920 ( .A(n1541), .B(A[306]), .Z(n4198) );
  AND U4921 ( .A(n4201), .B(n4202), .Z(n1541) );
  NAND U4922 ( .A(B[305]), .B(n4203), .Z(n4202) );
  NANDN U4923 ( .A(A[305]), .B(n1543), .Z(n4203) );
  NANDN U4924 ( .A(n1543), .B(A[305]), .Z(n4201) );
  AND U4925 ( .A(n4204), .B(n4205), .Z(n1543) );
  NAND U4926 ( .A(B[304]), .B(n4206), .Z(n4205) );
  NANDN U4927 ( .A(A[304]), .B(n1545), .Z(n4206) );
  NANDN U4928 ( .A(n1545), .B(A[304]), .Z(n4204) );
  AND U4929 ( .A(n4207), .B(n4208), .Z(n1545) );
  NAND U4930 ( .A(B[303]), .B(n4209), .Z(n4208) );
  NANDN U4931 ( .A(A[303]), .B(n1547), .Z(n4209) );
  NANDN U4932 ( .A(n1547), .B(A[303]), .Z(n4207) );
  AND U4933 ( .A(n4210), .B(n4211), .Z(n1547) );
  NAND U4934 ( .A(B[302]), .B(n4212), .Z(n4211) );
  NANDN U4935 ( .A(A[302]), .B(n1549), .Z(n4212) );
  NANDN U4936 ( .A(n1549), .B(A[302]), .Z(n4210) );
  AND U4937 ( .A(n4213), .B(n4214), .Z(n1549) );
  NAND U4938 ( .A(B[301]), .B(n4215), .Z(n4214) );
  NANDN U4939 ( .A(A[301]), .B(n1551), .Z(n4215) );
  NANDN U4940 ( .A(n1551), .B(A[301]), .Z(n4213) );
  AND U4941 ( .A(n4216), .B(n4217), .Z(n1551) );
  NAND U4942 ( .A(B[300]), .B(n4218), .Z(n4217) );
  NANDN U4943 ( .A(A[300]), .B(n1553), .Z(n4218) );
  NANDN U4944 ( .A(n1553), .B(A[300]), .Z(n4216) );
  AND U4945 ( .A(n4219), .B(n4220), .Z(n1553) );
  NAND U4946 ( .A(B[299]), .B(n4221), .Z(n4220) );
  NANDN U4947 ( .A(A[299]), .B(n1559), .Z(n4221) );
  NANDN U4948 ( .A(n1559), .B(A[299]), .Z(n4219) );
  AND U4949 ( .A(n4222), .B(n4223), .Z(n1559) );
  NAND U4950 ( .A(B[298]), .B(n4224), .Z(n4223) );
  NANDN U4951 ( .A(A[298]), .B(n1561), .Z(n4224) );
  NANDN U4952 ( .A(n1561), .B(A[298]), .Z(n4222) );
  AND U4953 ( .A(n4225), .B(n4226), .Z(n1561) );
  NAND U4954 ( .A(B[297]), .B(n4227), .Z(n4226) );
  NANDN U4955 ( .A(A[297]), .B(n1563), .Z(n4227) );
  NANDN U4956 ( .A(n1563), .B(A[297]), .Z(n4225) );
  AND U4957 ( .A(n4228), .B(n4229), .Z(n1563) );
  NAND U4958 ( .A(B[296]), .B(n4230), .Z(n4229) );
  NANDN U4959 ( .A(A[296]), .B(n1565), .Z(n4230) );
  NANDN U4960 ( .A(n1565), .B(A[296]), .Z(n4228) );
  AND U4961 ( .A(n4231), .B(n4232), .Z(n1565) );
  NAND U4962 ( .A(B[295]), .B(n4233), .Z(n4232) );
  NANDN U4963 ( .A(A[295]), .B(n1567), .Z(n4233) );
  NANDN U4964 ( .A(n1567), .B(A[295]), .Z(n4231) );
  AND U4965 ( .A(n4234), .B(n4235), .Z(n1567) );
  NAND U4966 ( .A(B[294]), .B(n4236), .Z(n4235) );
  NANDN U4967 ( .A(A[294]), .B(n1569), .Z(n4236) );
  NANDN U4968 ( .A(n1569), .B(A[294]), .Z(n4234) );
  AND U4969 ( .A(n4237), .B(n4238), .Z(n1569) );
  NAND U4970 ( .A(B[293]), .B(n4239), .Z(n4238) );
  NANDN U4971 ( .A(A[293]), .B(n1571), .Z(n4239) );
  NANDN U4972 ( .A(n1571), .B(A[293]), .Z(n4237) );
  AND U4973 ( .A(n4240), .B(n4241), .Z(n1571) );
  NAND U4974 ( .A(B[292]), .B(n4242), .Z(n4241) );
  NANDN U4975 ( .A(A[292]), .B(n1573), .Z(n4242) );
  NANDN U4976 ( .A(n1573), .B(A[292]), .Z(n4240) );
  AND U4977 ( .A(n4243), .B(n4244), .Z(n1573) );
  NAND U4978 ( .A(B[291]), .B(n4245), .Z(n4244) );
  NANDN U4979 ( .A(A[291]), .B(n1575), .Z(n4245) );
  NANDN U4980 ( .A(n1575), .B(A[291]), .Z(n4243) );
  AND U4981 ( .A(n4246), .B(n4247), .Z(n1575) );
  NAND U4982 ( .A(B[290]), .B(n4248), .Z(n4247) );
  NANDN U4983 ( .A(A[290]), .B(n1577), .Z(n4248) );
  NANDN U4984 ( .A(n1577), .B(A[290]), .Z(n4246) );
  AND U4985 ( .A(n4249), .B(n4250), .Z(n1577) );
  NAND U4986 ( .A(B[289]), .B(n4251), .Z(n4250) );
  NANDN U4987 ( .A(A[289]), .B(n1581), .Z(n4251) );
  NANDN U4988 ( .A(n1581), .B(A[289]), .Z(n4249) );
  AND U4989 ( .A(n4252), .B(n4253), .Z(n1581) );
  NAND U4990 ( .A(B[288]), .B(n4254), .Z(n4253) );
  NANDN U4991 ( .A(A[288]), .B(n1583), .Z(n4254) );
  NANDN U4992 ( .A(n1583), .B(A[288]), .Z(n4252) );
  AND U4993 ( .A(n4255), .B(n4256), .Z(n1583) );
  NAND U4994 ( .A(B[287]), .B(n4257), .Z(n4256) );
  NANDN U4995 ( .A(A[287]), .B(n1585), .Z(n4257) );
  NANDN U4996 ( .A(n1585), .B(A[287]), .Z(n4255) );
  AND U4997 ( .A(n4258), .B(n4259), .Z(n1585) );
  NAND U4998 ( .A(B[286]), .B(n4260), .Z(n4259) );
  NANDN U4999 ( .A(A[286]), .B(n1587), .Z(n4260) );
  NANDN U5000 ( .A(n1587), .B(A[286]), .Z(n4258) );
  AND U5001 ( .A(n4261), .B(n4262), .Z(n1587) );
  NAND U5002 ( .A(B[285]), .B(n4263), .Z(n4262) );
  NANDN U5003 ( .A(A[285]), .B(n1589), .Z(n4263) );
  NANDN U5004 ( .A(n1589), .B(A[285]), .Z(n4261) );
  AND U5005 ( .A(n4264), .B(n4265), .Z(n1589) );
  NAND U5006 ( .A(B[284]), .B(n4266), .Z(n4265) );
  NANDN U5007 ( .A(A[284]), .B(n1591), .Z(n4266) );
  NANDN U5008 ( .A(n1591), .B(A[284]), .Z(n4264) );
  AND U5009 ( .A(n4267), .B(n4268), .Z(n1591) );
  NAND U5010 ( .A(B[283]), .B(n4269), .Z(n4268) );
  NANDN U5011 ( .A(A[283]), .B(n1593), .Z(n4269) );
  NANDN U5012 ( .A(n1593), .B(A[283]), .Z(n4267) );
  AND U5013 ( .A(n4270), .B(n4271), .Z(n1593) );
  NAND U5014 ( .A(B[282]), .B(n4272), .Z(n4271) );
  NANDN U5015 ( .A(A[282]), .B(n1595), .Z(n4272) );
  NANDN U5016 ( .A(n1595), .B(A[282]), .Z(n4270) );
  AND U5017 ( .A(n4273), .B(n4274), .Z(n1595) );
  NAND U5018 ( .A(B[281]), .B(n4275), .Z(n4274) );
  NANDN U5019 ( .A(A[281]), .B(n1597), .Z(n4275) );
  NANDN U5020 ( .A(n1597), .B(A[281]), .Z(n4273) );
  AND U5021 ( .A(n4276), .B(n4277), .Z(n1597) );
  NAND U5022 ( .A(B[280]), .B(n4278), .Z(n4277) );
  NANDN U5023 ( .A(A[280]), .B(n1599), .Z(n4278) );
  NANDN U5024 ( .A(n1599), .B(A[280]), .Z(n4276) );
  AND U5025 ( .A(n4279), .B(n4280), .Z(n1599) );
  NAND U5026 ( .A(B[279]), .B(n4281), .Z(n4280) );
  NANDN U5027 ( .A(A[279]), .B(n1603), .Z(n4281) );
  NANDN U5028 ( .A(n1603), .B(A[279]), .Z(n4279) );
  AND U5029 ( .A(n4282), .B(n4283), .Z(n1603) );
  NAND U5030 ( .A(B[278]), .B(n4284), .Z(n4283) );
  NANDN U5031 ( .A(A[278]), .B(n1605), .Z(n4284) );
  NANDN U5032 ( .A(n1605), .B(A[278]), .Z(n4282) );
  AND U5033 ( .A(n4285), .B(n4286), .Z(n1605) );
  NAND U5034 ( .A(B[277]), .B(n4287), .Z(n4286) );
  NANDN U5035 ( .A(A[277]), .B(n1607), .Z(n4287) );
  NANDN U5036 ( .A(n1607), .B(A[277]), .Z(n4285) );
  AND U5037 ( .A(n4288), .B(n4289), .Z(n1607) );
  NAND U5038 ( .A(B[276]), .B(n4290), .Z(n4289) );
  NANDN U5039 ( .A(A[276]), .B(n1609), .Z(n4290) );
  NANDN U5040 ( .A(n1609), .B(A[276]), .Z(n4288) );
  AND U5041 ( .A(n4291), .B(n4292), .Z(n1609) );
  NAND U5042 ( .A(B[275]), .B(n4293), .Z(n4292) );
  NANDN U5043 ( .A(A[275]), .B(n1611), .Z(n4293) );
  NANDN U5044 ( .A(n1611), .B(A[275]), .Z(n4291) );
  AND U5045 ( .A(n4294), .B(n4295), .Z(n1611) );
  NAND U5046 ( .A(B[274]), .B(n4296), .Z(n4295) );
  NANDN U5047 ( .A(A[274]), .B(n1613), .Z(n4296) );
  NANDN U5048 ( .A(n1613), .B(A[274]), .Z(n4294) );
  AND U5049 ( .A(n4297), .B(n4298), .Z(n1613) );
  NAND U5050 ( .A(B[273]), .B(n4299), .Z(n4298) );
  NANDN U5051 ( .A(A[273]), .B(n1615), .Z(n4299) );
  NANDN U5052 ( .A(n1615), .B(A[273]), .Z(n4297) );
  AND U5053 ( .A(n4300), .B(n4301), .Z(n1615) );
  NAND U5054 ( .A(B[272]), .B(n4302), .Z(n4301) );
  NANDN U5055 ( .A(A[272]), .B(n1617), .Z(n4302) );
  NANDN U5056 ( .A(n1617), .B(A[272]), .Z(n4300) );
  AND U5057 ( .A(n4303), .B(n4304), .Z(n1617) );
  NAND U5058 ( .A(B[271]), .B(n4305), .Z(n4304) );
  NANDN U5059 ( .A(A[271]), .B(n1619), .Z(n4305) );
  NANDN U5060 ( .A(n1619), .B(A[271]), .Z(n4303) );
  AND U5061 ( .A(n4306), .B(n4307), .Z(n1619) );
  NAND U5062 ( .A(B[270]), .B(n4308), .Z(n4307) );
  NANDN U5063 ( .A(A[270]), .B(n1621), .Z(n4308) );
  NANDN U5064 ( .A(n1621), .B(A[270]), .Z(n4306) );
  AND U5065 ( .A(n4309), .B(n4310), .Z(n1621) );
  NAND U5066 ( .A(B[269]), .B(n4311), .Z(n4310) );
  NANDN U5067 ( .A(A[269]), .B(n1625), .Z(n4311) );
  NANDN U5068 ( .A(n1625), .B(A[269]), .Z(n4309) );
  AND U5069 ( .A(n4312), .B(n4313), .Z(n1625) );
  NAND U5070 ( .A(B[268]), .B(n4314), .Z(n4313) );
  NANDN U5071 ( .A(A[268]), .B(n1627), .Z(n4314) );
  NANDN U5072 ( .A(n1627), .B(A[268]), .Z(n4312) );
  AND U5073 ( .A(n4315), .B(n4316), .Z(n1627) );
  NAND U5074 ( .A(B[267]), .B(n4317), .Z(n4316) );
  NANDN U5075 ( .A(A[267]), .B(n1629), .Z(n4317) );
  NANDN U5076 ( .A(n1629), .B(A[267]), .Z(n4315) );
  AND U5077 ( .A(n4318), .B(n4319), .Z(n1629) );
  NAND U5078 ( .A(B[266]), .B(n4320), .Z(n4319) );
  NANDN U5079 ( .A(A[266]), .B(n1631), .Z(n4320) );
  NANDN U5080 ( .A(n1631), .B(A[266]), .Z(n4318) );
  AND U5081 ( .A(n4321), .B(n4322), .Z(n1631) );
  NAND U5082 ( .A(B[265]), .B(n4323), .Z(n4322) );
  NANDN U5083 ( .A(A[265]), .B(n1633), .Z(n4323) );
  NANDN U5084 ( .A(n1633), .B(A[265]), .Z(n4321) );
  AND U5085 ( .A(n4324), .B(n4325), .Z(n1633) );
  NAND U5086 ( .A(B[264]), .B(n4326), .Z(n4325) );
  NANDN U5087 ( .A(A[264]), .B(n1635), .Z(n4326) );
  NANDN U5088 ( .A(n1635), .B(A[264]), .Z(n4324) );
  AND U5089 ( .A(n4327), .B(n4328), .Z(n1635) );
  NAND U5090 ( .A(B[263]), .B(n4329), .Z(n4328) );
  NANDN U5091 ( .A(A[263]), .B(n1637), .Z(n4329) );
  NANDN U5092 ( .A(n1637), .B(A[263]), .Z(n4327) );
  AND U5093 ( .A(n4330), .B(n4331), .Z(n1637) );
  NAND U5094 ( .A(B[262]), .B(n4332), .Z(n4331) );
  NANDN U5095 ( .A(A[262]), .B(n1639), .Z(n4332) );
  NANDN U5096 ( .A(n1639), .B(A[262]), .Z(n4330) );
  AND U5097 ( .A(n4333), .B(n4334), .Z(n1639) );
  NAND U5098 ( .A(B[261]), .B(n4335), .Z(n4334) );
  NANDN U5099 ( .A(A[261]), .B(n1641), .Z(n4335) );
  NANDN U5100 ( .A(n1641), .B(A[261]), .Z(n4333) );
  AND U5101 ( .A(n4336), .B(n4337), .Z(n1641) );
  NAND U5102 ( .A(B[260]), .B(n4338), .Z(n4337) );
  NANDN U5103 ( .A(A[260]), .B(n1643), .Z(n4338) );
  NANDN U5104 ( .A(n1643), .B(A[260]), .Z(n4336) );
  AND U5105 ( .A(n4339), .B(n4340), .Z(n1643) );
  NAND U5106 ( .A(B[259]), .B(n4341), .Z(n4340) );
  NANDN U5107 ( .A(A[259]), .B(n1647), .Z(n4341) );
  NANDN U5108 ( .A(n1647), .B(A[259]), .Z(n4339) );
  AND U5109 ( .A(n4342), .B(n4343), .Z(n1647) );
  NAND U5110 ( .A(B[258]), .B(n4344), .Z(n4343) );
  NANDN U5111 ( .A(A[258]), .B(n1649), .Z(n4344) );
  NANDN U5112 ( .A(n1649), .B(A[258]), .Z(n4342) );
  AND U5113 ( .A(n4345), .B(n4346), .Z(n1649) );
  NAND U5114 ( .A(B[257]), .B(n4347), .Z(n4346) );
  NANDN U5115 ( .A(A[257]), .B(n1651), .Z(n4347) );
  NANDN U5116 ( .A(n1651), .B(A[257]), .Z(n4345) );
  AND U5117 ( .A(n4348), .B(n4349), .Z(n1651) );
  NAND U5118 ( .A(B[256]), .B(n4350), .Z(n4349) );
  NANDN U5119 ( .A(A[256]), .B(n1653), .Z(n4350) );
  NANDN U5120 ( .A(n1653), .B(A[256]), .Z(n4348) );
  AND U5121 ( .A(n4351), .B(n4352), .Z(n1653) );
  NAND U5122 ( .A(B[255]), .B(n4353), .Z(n4352) );
  NANDN U5123 ( .A(A[255]), .B(n1655), .Z(n4353) );
  NANDN U5124 ( .A(n1655), .B(A[255]), .Z(n4351) );
  AND U5125 ( .A(n4354), .B(n4355), .Z(n1655) );
  NAND U5126 ( .A(B[254]), .B(n4356), .Z(n4355) );
  NANDN U5127 ( .A(A[254]), .B(n1657), .Z(n4356) );
  NANDN U5128 ( .A(n1657), .B(A[254]), .Z(n4354) );
  AND U5129 ( .A(n4357), .B(n4358), .Z(n1657) );
  NAND U5130 ( .A(B[253]), .B(n4359), .Z(n4358) );
  NANDN U5131 ( .A(A[253]), .B(n1659), .Z(n4359) );
  NANDN U5132 ( .A(n1659), .B(A[253]), .Z(n4357) );
  AND U5133 ( .A(n4360), .B(n4361), .Z(n1659) );
  NAND U5134 ( .A(B[252]), .B(n4362), .Z(n4361) );
  NANDN U5135 ( .A(A[252]), .B(n1661), .Z(n4362) );
  NANDN U5136 ( .A(n1661), .B(A[252]), .Z(n4360) );
  AND U5137 ( .A(n4363), .B(n4364), .Z(n1661) );
  NAND U5138 ( .A(B[251]), .B(n4365), .Z(n4364) );
  NANDN U5139 ( .A(A[251]), .B(n1663), .Z(n4365) );
  NANDN U5140 ( .A(n1663), .B(A[251]), .Z(n4363) );
  AND U5141 ( .A(n4366), .B(n4367), .Z(n1663) );
  NAND U5142 ( .A(B[250]), .B(n4368), .Z(n4367) );
  NANDN U5143 ( .A(A[250]), .B(n1665), .Z(n4368) );
  NANDN U5144 ( .A(n1665), .B(A[250]), .Z(n4366) );
  AND U5145 ( .A(n4369), .B(n4370), .Z(n1665) );
  NAND U5146 ( .A(B[249]), .B(n4371), .Z(n4370) );
  NANDN U5147 ( .A(A[249]), .B(n1669), .Z(n4371) );
  NANDN U5148 ( .A(n1669), .B(A[249]), .Z(n4369) );
  AND U5149 ( .A(n4372), .B(n4373), .Z(n1669) );
  NAND U5150 ( .A(B[248]), .B(n4374), .Z(n4373) );
  NANDN U5151 ( .A(A[248]), .B(n1671), .Z(n4374) );
  NANDN U5152 ( .A(n1671), .B(A[248]), .Z(n4372) );
  AND U5153 ( .A(n4375), .B(n4376), .Z(n1671) );
  NAND U5154 ( .A(B[247]), .B(n4377), .Z(n4376) );
  NANDN U5155 ( .A(A[247]), .B(n1673), .Z(n4377) );
  NANDN U5156 ( .A(n1673), .B(A[247]), .Z(n4375) );
  AND U5157 ( .A(n4378), .B(n4379), .Z(n1673) );
  NAND U5158 ( .A(B[246]), .B(n4380), .Z(n4379) );
  NANDN U5159 ( .A(A[246]), .B(n1675), .Z(n4380) );
  NANDN U5160 ( .A(n1675), .B(A[246]), .Z(n4378) );
  AND U5161 ( .A(n4381), .B(n4382), .Z(n1675) );
  NAND U5162 ( .A(B[245]), .B(n4383), .Z(n4382) );
  NANDN U5163 ( .A(A[245]), .B(n1677), .Z(n4383) );
  NANDN U5164 ( .A(n1677), .B(A[245]), .Z(n4381) );
  AND U5165 ( .A(n4384), .B(n4385), .Z(n1677) );
  NAND U5166 ( .A(B[244]), .B(n4386), .Z(n4385) );
  NANDN U5167 ( .A(A[244]), .B(n1679), .Z(n4386) );
  NANDN U5168 ( .A(n1679), .B(A[244]), .Z(n4384) );
  AND U5169 ( .A(n4387), .B(n4388), .Z(n1679) );
  NAND U5170 ( .A(B[243]), .B(n4389), .Z(n4388) );
  NANDN U5171 ( .A(A[243]), .B(n1681), .Z(n4389) );
  NANDN U5172 ( .A(n1681), .B(A[243]), .Z(n4387) );
  AND U5173 ( .A(n4390), .B(n4391), .Z(n1681) );
  NAND U5174 ( .A(B[242]), .B(n4392), .Z(n4391) );
  NANDN U5175 ( .A(A[242]), .B(n1683), .Z(n4392) );
  NANDN U5176 ( .A(n1683), .B(A[242]), .Z(n4390) );
  AND U5177 ( .A(n4393), .B(n4394), .Z(n1683) );
  NAND U5178 ( .A(B[241]), .B(n4395), .Z(n4394) );
  NANDN U5179 ( .A(A[241]), .B(n1685), .Z(n4395) );
  NANDN U5180 ( .A(n1685), .B(A[241]), .Z(n4393) );
  AND U5181 ( .A(n4396), .B(n4397), .Z(n1685) );
  NAND U5182 ( .A(B[240]), .B(n4398), .Z(n4397) );
  NANDN U5183 ( .A(A[240]), .B(n1687), .Z(n4398) );
  NANDN U5184 ( .A(n1687), .B(A[240]), .Z(n4396) );
  AND U5185 ( .A(n4399), .B(n4400), .Z(n1687) );
  NAND U5186 ( .A(B[239]), .B(n4401), .Z(n4400) );
  NANDN U5187 ( .A(A[239]), .B(n1691), .Z(n4401) );
  NANDN U5188 ( .A(n1691), .B(A[239]), .Z(n4399) );
  AND U5189 ( .A(n4402), .B(n4403), .Z(n1691) );
  NAND U5190 ( .A(B[238]), .B(n4404), .Z(n4403) );
  NANDN U5191 ( .A(A[238]), .B(n1693), .Z(n4404) );
  NANDN U5192 ( .A(n1693), .B(A[238]), .Z(n4402) );
  AND U5193 ( .A(n4405), .B(n4406), .Z(n1693) );
  NAND U5194 ( .A(B[237]), .B(n4407), .Z(n4406) );
  NANDN U5195 ( .A(A[237]), .B(n1695), .Z(n4407) );
  NANDN U5196 ( .A(n1695), .B(A[237]), .Z(n4405) );
  AND U5197 ( .A(n4408), .B(n4409), .Z(n1695) );
  NAND U5198 ( .A(B[236]), .B(n4410), .Z(n4409) );
  NANDN U5199 ( .A(A[236]), .B(n1697), .Z(n4410) );
  NANDN U5200 ( .A(n1697), .B(A[236]), .Z(n4408) );
  AND U5201 ( .A(n4411), .B(n4412), .Z(n1697) );
  NAND U5202 ( .A(B[235]), .B(n4413), .Z(n4412) );
  NANDN U5203 ( .A(A[235]), .B(n1699), .Z(n4413) );
  NANDN U5204 ( .A(n1699), .B(A[235]), .Z(n4411) );
  AND U5205 ( .A(n4414), .B(n4415), .Z(n1699) );
  NAND U5206 ( .A(B[234]), .B(n4416), .Z(n4415) );
  NANDN U5207 ( .A(A[234]), .B(n1701), .Z(n4416) );
  NANDN U5208 ( .A(n1701), .B(A[234]), .Z(n4414) );
  AND U5209 ( .A(n4417), .B(n4418), .Z(n1701) );
  NAND U5210 ( .A(B[233]), .B(n4419), .Z(n4418) );
  NANDN U5211 ( .A(A[233]), .B(n1703), .Z(n4419) );
  NANDN U5212 ( .A(n1703), .B(A[233]), .Z(n4417) );
  AND U5213 ( .A(n4420), .B(n4421), .Z(n1703) );
  NAND U5214 ( .A(B[232]), .B(n4422), .Z(n4421) );
  NANDN U5215 ( .A(A[232]), .B(n1705), .Z(n4422) );
  NANDN U5216 ( .A(n1705), .B(A[232]), .Z(n4420) );
  AND U5217 ( .A(n4423), .B(n4424), .Z(n1705) );
  NAND U5218 ( .A(B[231]), .B(n4425), .Z(n4424) );
  NANDN U5219 ( .A(A[231]), .B(n1707), .Z(n4425) );
  NANDN U5220 ( .A(n1707), .B(A[231]), .Z(n4423) );
  AND U5221 ( .A(n4426), .B(n4427), .Z(n1707) );
  NAND U5222 ( .A(B[230]), .B(n4428), .Z(n4427) );
  NANDN U5223 ( .A(A[230]), .B(n1709), .Z(n4428) );
  NANDN U5224 ( .A(n1709), .B(A[230]), .Z(n4426) );
  AND U5225 ( .A(n4429), .B(n4430), .Z(n1709) );
  NAND U5226 ( .A(B[229]), .B(n4431), .Z(n4430) );
  NANDN U5227 ( .A(A[229]), .B(n1713), .Z(n4431) );
  NANDN U5228 ( .A(n1713), .B(A[229]), .Z(n4429) );
  AND U5229 ( .A(n4432), .B(n4433), .Z(n1713) );
  NAND U5230 ( .A(B[228]), .B(n4434), .Z(n4433) );
  NANDN U5231 ( .A(A[228]), .B(n1715), .Z(n4434) );
  NANDN U5232 ( .A(n1715), .B(A[228]), .Z(n4432) );
  AND U5233 ( .A(n4435), .B(n4436), .Z(n1715) );
  NAND U5234 ( .A(B[227]), .B(n4437), .Z(n4436) );
  NANDN U5235 ( .A(A[227]), .B(n1717), .Z(n4437) );
  NANDN U5236 ( .A(n1717), .B(A[227]), .Z(n4435) );
  AND U5237 ( .A(n4438), .B(n4439), .Z(n1717) );
  NAND U5238 ( .A(B[226]), .B(n4440), .Z(n4439) );
  NANDN U5239 ( .A(A[226]), .B(n1719), .Z(n4440) );
  NANDN U5240 ( .A(n1719), .B(A[226]), .Z(n4438) );
  AND U5241 ( .A(n4441), .B(n4442), .Z(n1719) );
  NAND U5242 ( .A(B[225]), .B(n4443), .Z(n4442) );
  NANDN U5243 ( .A(A[225]), .B(n1721), .Z(n4443) );
  NANDN U5244 ( .A(n1721), .B(A[225]), .Z(n4441) );
  AND U5245 ( .A(n4444), .B(n4445), .Z(n1721) );
  NAND U5246 ( .A(B[224]), .B(n4446), .Z(n4445) );
  NANDN U5247 ( .A(A[224]), .B(n1723), .Z(n4446) );
  NANDN U5248 ( .A(n1723), .B(A[224]), .Z(n4444) );
  AND U5249 ( .A(n4447), .B(n4448), .Z(n1723) );
  NAND U5250 ( .A(B[223]), .B(n4449), .Z(n4448) );
  NANDN U5251 ( .A(A[223]), .B(n1725), .Z(n4449) );
  NANDN U5252 ( .A(n1725), .B(A[223]), .Z(n4447) );
  AND U5253 ( .A(n4450), .B(n4451), .Z(n1725) );
  NAND U5254 ( .A(B[222]), .B(n4452), .Z(n4451) );
  NANDN U5255 ( .A(A[222]), .B(n1727), .Z(n4452) );
  NANDN U5256 ( .A(n1727), .B(A[222]), .Z(n4450) );
  AND U5257 ( .A(n4453), .B(n4454), .Z(n1727) );
  NAND U5258 ( .A(B[221]), .B(n4455), .Z(n4454) );
  NANDN U5259 ( .A(A[221]), .B(n1729), .Z(n4455) );
  NANDN U5260 ( .A(n1729), .B(A[221]), .Z(n4453) );
  AND U5261 ( .A(n4456), .B(n4457), .Z(n1729) );
  NAND U5262 ( .A(B[220]), .B(n4458), .Z(n4457) );
  NANDN U5263 ( .A(A[220]), .B(n1731), .Z(n4458) );
  NANDN U5264 ( .A(n1731), .B(A[220]), .Z(n4456) );
  AND U5265 ( .A(n4459), .B(n4460), .Z(n1731) );
  NAND U5266 ( .A(B[219]), .B(n4461), .Z(n4460) );
  NANDN U5267 ( .A(A[219]), .B(n1735), .Z(n4461) );
  NANDN U5268 ( .A(n1735), .B(A[219]), .Z(n4459) );
  AND U5269 ( .A(n4462), .B(n4463), .Z(n1735) );
  NAND U5270 ( .A(B[218]), .B(n4464), .Z(n4463) );
  NANDN U5271 ( .A(A[218]), .B(n1737), .Z(n4464) );
  NANDN U5272 ( .A(n1737), .B(A[218]), .Z(n4462) );
  AND U5273 ( .A(n4465), .B(n4466), .Z(n1737) );
  NAND U5274 ( .A(B[217]), .B(n4467), .Z(n4466) );
  NANDN U5275 ( .A(A[217]), .B(n1739), .Z(n4467) );
  NANDN U5276 ( .A(n1739), .B(A[217]), .Z(n4465) );
  AND U5277 ( .A(n4468), .B(n4469), .Z(n1739) );
  NAND U5278 ( .A(B[216]), .B(n4470), .Z(n4469) );
  NANDN U5279 ( .A(A[216]), .B(n1741), .Z(n4470) );
  NANDN U5280 ( .A(n1741), .B(A[216]), .Z(n4468) );
  AND U5281 ( .A(n4471), .B(n4472), .Z(n1741) );
  NAND U5282 ( .A(B[215]), .B(n4473), .Z(n4472) );
  NANDN U5283 ( .A(A[215]), .B(n1743), .Z(n4473) );
  NANDN U5284 ( .A(n1743), .B(A[215]), .Z(n4471) );
  AND U5285 ( .A(n4474), .B(n4475), .Z(n1743) );
  NAND U5286 ( .A(B[214]), .B(n4476), .Z(n4475) );
  NANDN U5287 ( .A(A[214]), .B(n1745), .Z(n4476) );
  NANDN U5288 ( .A(n1745), .B(A[214]), .Z(n4474) );
  AND U5289 ( .A(n4477), .B(n4478), .Z(n1745) );
  NAND U5290 ( .A(B[213]), .B(n4479), .Z(n4478) );
  NANDN U5291 ( .A(A[213]), .B(n1747), .Z(n4479) );
  NANDN U5292 ( .A(n1747), .B(A[213]), .Z(n4477) );
  AND U5293 ( .A(n4480), .B(n4481), .Z(n1747) );
  NAND U5294 ( .A(B[212]), .B(n4482), .Z(n4481) );
  NANDN U5295 ( .A(A[212]), .B(n1749), .Z(n4482) );
  NANDN U5296 ( .A(n1749), .B(A[212]), .Z(n4480) );
  AND U5297 ( .A(n4483), .B(n4484), .Z(n1749) );
  NAND U5298 ( .A(B[211]), .B(n4485), .Z(n4484) );
  NANDN U5299 ( .A(A[211]), .B(n1751), .Z(n4485) );
  NANDN U5300 ( .A(n1751), .B(A[211]), .Z(n4483) );
  AND U5301 ( .A(n4486), .B(n4487), .Z(n1751) );
  NAND U5302 ( .A(B[210]), .B(n4488), .Z(n4487) );
  NANDN U5303 ( .A(A[210]), .B(n1753), .Z(n4488) );
  NANDN U5304 ( .A(n1753), .B(A[210]), .Z(n4486) );
  AND U5305 ( .A(n4489), .B(n4490), .Z(n1753) );
  NAND U5306 ( .A(B[209]), .B(n4491), .Z(n4490) );
  NANDN U5307 ( .A(A[209]), .B(n1757), .Z(n4491) );
  NANDN U5308 ( .A(n1757), .B(A[209]), .Z(n4489) );
  AND U5309 ( .A(n4492), .B(n4493), .Z(n1757) );
  NAND U5310 ( .A(B[208]), .B(n4494), .Z(n4493) );
  NANDN U5311 ( .A(A[208]), .B(n1759), .Z(n4494) );
  NANDN U5312 ( .A(n1759), .B(A[208]), .Z(n4492) );
  AND U5313 ( .A(n4495), .B(n4496), .Z(n1759) );
  NAND U5314 ( .A(B[207]), .B(n4497), .Z(n4496) );
  NANDN U5315 ( .A(A[207]), .B(n1761), .Z(n4497) );
  NANDN U5316 ( .A(n1761), .B(A[207]), .Z(n4495) );
  AND U5317 ( .A(n4498), .B(n4499), .Z(n1761) );
  NAND U5318 ( .A(B[206]), .B(n4500), .Z(n4499) );
  NANDN U5319 ( .A(A[206]), .B(n1763), .Z(n4500) );
  NANDN U5320 ( .A(n1763), .B(A[206]), .Z(n4498) );
  AND U5321 ( .A(n4501), .B(n4502), .Z(n1763) );
  NAND U5322 ( .A(B[205]), .B(n4503), .Z(n4502) );
  NANDN U5323 ( .A(A[205]), .B(n1765), .Z(n4503) );
  NANDN U5324 ( .A(n1765), .B(A[205]), .Z(n4501) );
  AND U5325 ( .A(n4504), .B(n4505), .Z(n1765) );
  NAND U5326 ( .A(B[204]), .B(n4506), .Z(n4505) );
  NANDN U5327 ( .A(A[204]), .B(n1767), .Z(n4506) );
  NANDN U5328 ( .A(n1767), .B(A[204]), .Z(n4504) );
  AND U5329 ( .A(n4507), .B(n4508), .Z(n1767) );
  NAND U5330 ( .A(B[203]), .B(n4509), .Z(n4508) );
  NANDN U5331 ( .A(A[203]), .B(n1769), .Z(n4509) );
  NANDN U5332 ( .A(n1769), .B(A[203]), .Z(n4507) );
  AND U5333 ( .A(n4510), .B(n4511), .Z(n1769) );
  NAND U5334 ( .A(B[202]), .B(n4512), .Z(n4511) );
  NANDN U5335 ( .A(A[202]), .B(n1771), .Z(n4512) );
  NANDN U5336 ( .A(n1771), .B(A[202]), .Z(n4510) );
  AND U5337 ( .A(n4513), .B(n4514), .Z(n1771) );
  NAND U5338 ( .A(B[201]), .B(n4515), .Z(n4514) );
  NANDN U5339 ( .A(A[201]), .B(n1773), .Z(n4515) );
  NANDN U5340 ( .A(n1773), .B(A[201]), .Z(n4513) );
  AND U5341 ( .A(n4516), .B(n4517), .Z(n1773) );
  NAND U5342 ( .A(B[200]), .B(n4518), .Z(n4517) );
  NANDN U5343 ( .A(A[200]), .B(n1775), .Z(n4518) );
  NANDN U5344 ( .A(n1775), .B(A[200]), .Z(n4516) );
  AND U5345 ( .A(n4519), .B(n4520), .Z(n1775) );
  NAND U5346 ( .A(B[199]), .B(n4521), .Z(n4520) );
  NANDN U5347 ( .A(A[199]), .B(n1779), .Z(n4521) );
  NANDN U5348 ( .A(n1779), .B(A[199]), .Z(n4519) );
  AND U5349 ( .A(n4522), .B(n4523), .Z(n1779) );
  NAND U5350 ( .A(B[198]), .B(n4524), .Z(n4523) );
  NANDN U5351 ( .A(A[198]), .B(n1781), .Z(n4524) );
  NANDN U5352 ( .A(n1781), .B(A[198]), .Z(n4522) );
  AND U5353 ( .A(n4525), .B(n4526), .Z(n1781) );
  NAND U5354 ( .A(B[197]), .B(n4527), .Z(n4526) );
  NANDN U5355 ( .A(A[197]), .B(n1783), .Z(n4527) );
  NANDN U5356 ( .A(n1783), .B(A[197]), .Z(n4525) );
  AND U5357 ( .A(n4528), .B(n4529), .Z(n1783) );
  NAND U5358 ( .A(B[196]), .B(n4530), .Z(n4529) );
  NANDN U5359 ( .A(A[196]), .B(n1785), .Z(n4530) );
  NANDN U5360 ( .A(n1785), .B(A[196]), .Z(n4528) );
  AND U5361 ( .A(n4531), .B(n4532), .Z(n1785) );
  NAND U5362 ( .A(B[195]), .B(n4533), .Z(n4532) );
  NANDN U5363 ( .A(A[195]), .B(n1787), .Z(n4533) );
  NANDN U5364 ( .A(n1787), .B(A[195]), .Z(n4531) );
  AND U5365 ( .A(n4534), .B(n4535), .Z(n1787) );
  NAND U5366 ( .A(B[194]), .B(n4536), .Z(n4535) );
  NANDN U5367 ( .A(A[194]), .B(n1789), .Z(n4536) );
  NANDN U5368 ( .A(n1789), .B(A[194]), .Z(n4534) );
  AND U5369 ( .A(n4537), .B(n4538), .Z(n1789) );
  NAND U5370 ( .A(B[193]), .B(n4539), .Z(n4538) );
  NANDN U5371 ( .A(A[193]), .B(n1791), .Z(n4539) );
  NANDN U5372 ( .A(n1791), .B(A[193]), .Z(n4537) );
  AND U5373 ( .A(n4540), .B(n4541), .Z(n1791) );
  NAND U5374 ( .A(B[192]), .B(n4542), .Z(n4541) );
  NANDN U5375 ( .A(A[192]), .B(n1793), .Z(n4542) );
  NANDN U5376 ( .A(n1793), .B(A[192]), .Z(n4540) );
  AND U5377 ( .A(n4543), .B(n4544), .Z(n1793) );
  NAND U5378 ( .A(B[191]), .B(n4545), .Z(n4544) );
  NANDN U5379 ( .A(A[191]), .B(n1795), .Z(n4545) );
  NANDN U5380 ( .A(n1795), .B(A[191]), .Z(n4543) );
  AND U5381 ( .A(n4546), .B(n4547), .Z(n1795) );
  NAND U5382 ( .A(B[190]), .B(n4548), .Z(n4547) );
  NANDN U5383 ( .A(A[190]), .B(n1797), .Z(n4548) );
  NANDN U5384 ( .A(n1797), .B(A[190]), .Z(n4546) );
  AND U5385 ( .A(n4549), .B(n4550), .Z(n1797) );
  NAND U5386 ( .A(B[189]), .B(n4551), .Z(n4550) );
  NANDN U5387 ( .A(A[189]), .B(n1801), .Z(n4551) );
  NANDN U5388 ( .A(n1801), .B(A[189]), .Z(n4549) );
  AND U5389 ( .A(n4552), .B(n4553), .Z(n1801) );
  NAND U5390 ( .A(B[188]), .B(n4554), .Z(n4553) );
  NANDN U5391 ( .A(A[188]), .B(n1803), .Z(n4554) );
  NANDN U5392 ( .A(n1803), .B(A[188]), .Z(n4552) );
  AND U5393 ( .A(n4555), .B(n4556), .Z(n1803) );
  NAND U5394 ( .A(B[187]), .B(n4557), .Z(n4556) );
  NANDN U5395 ( .A(A[187]), .B(n1805), .Z(n4557) );
  NANDN U5396 ( .A(n1805), .B(A[187]), .Z(n4555) );
  AND U5397 ( .A(n4558), .B(n4559), .Z(n1805) );
  NAND U5398 ( .A(B[186]), .B(n4560), .Z(n4559) );
  NANDN U5399 ( .A(A[186]), .B(n1807), .Z(n4560) );
  NANDN U5400 ( .A(n1807), .B(A[186]), .Z(n4558) );
  AND U5401 ( .A(n4561), .B(n4562), .Z(n1807) );
  NAND U5402 ( .A(B[185]), .B(n4563), .Z(n4562) );
  NANDN U5403 ( .A(A[185]), .B(n1809), .Z(n4563) );
  NANDN U5404 ( .A(n1809), .B(A[185]), .Z(n4561) );
  AND U5405 ( .A(n4564), .B(n4565), .Z(n1809) );
  NAND U5406 ( .A(B[184]), .B(n4566), .Z(n4565) );
  NANDN U5407 ( .A(A[184]), .B(n1811), .Z(n4566) );
  NANDN U5408 ( .A(n1811), .B(A[184]), .Z(n4564) );
  AND U5409 ( .A(n4567), .B(n4568), .Z(n1811) );
  NAND U5410 ( .A(B[183]), .B(n4569), .Z(n4568) );
  NANDN U5411 ( .A(A[183]), .B(n1813), .Z(n4569) );
  NANDN U5412 ( .A(n1813), .B(A[183]), .Z(n4567) );
  AND U5413 ( .A(n4570), .B(n4571), .Z(n1813) );
  NAND U5414 ( .A(B[182]), .B(n4572), .Z(n4571) );
  NANDN U5415 ( .A(A[182]), .B(n1815), .Z(n4572) );
  NANDN U5416 ( .A(n1815), .B(A[182]), .Z(n4570) );
  AND U5417 ( .A(n4573), .B(n4574), .Z(n1815) );
  NAND U5418 ( .A(B[181]), .B(n4575), .Z(n4574) );
  NANDN U5419 ( .A(A[181]), .B(n1817), .Z(n4575) );
  NANDN U5420 ( .A(n1817), .B(A[181]), .Z(n4573) );
  AND U5421 ( .A(n4576), .B(n4577), .Z(n1817) );
  NAND U5422 ( .A(B[180]), .B(n4578), .Z(n4577) );
  NANDN U5423 ( .A(A[180]), .B(n1819), .Z(n4578) );
  NANDN U5424 ( .A(n1819), .B(A[180]), .Z(n4576) );
  AND U5425 ( .A(n4579), .B(n4580), .Z(n1819) );
  NAND U5426 ( .A(B[179]), .B(n4581), .Z(n4580) );
  NANDN U5427 ( .A(A[179]), .B(n1823), .Z(n4581) );
  NANDN U5428 ( .A(n1823), .B(A[179]), .Z(n4579) );
  AND U5429 ( .A(n4582), .B(n4583), .Z(n1823) );
  NAND U5430 ( .A(B[178]), .B(n4584), .Z(n4583) );
  NANDN U5431 ( .A(A[178]), .B(n1825), .Z(n4584) );
  NANDN U5432 ( .A(n1825), .B(A[178]), .Z(n4582) );
  AND U5433 ( .A(n4585), .B(n4586), .Z(n1825) );
  NAND U5434 ( .A(B[177]), .B(n4587), .Z(n4586) );
  NANDN U5435 ( .A(A[177]), .B(n1827), .Z(n4587) );
  NANDN U5436 ( .A(n1827), .B(A[177]), .Z(n4585) );
  AND U5437 ( .A(n4588), .B(n4589), .Z(n1827) );
  NAND U5438 ( .A(B[176]), .B(n4590), .Z(n4589) );
  NANDN U5439 ( .A(A[176]), .B(n1829), .Z(n4590) );
  NANDN U5440 ( .A(n1829), .B(A[176]), .Z(n4588) );
  AND U5441 ( .A(n4591), .B(n4592), .Z(n1829) );
  NAND U5442 ( .A(B[175]), .B(n4593), .Z(n4592) );
  NANDN U5443 ( .A(A[175]), .B(n1831), .Z(n4593) );
  NANDN U5444 ( .A(n1831), .B(A[175]), .Z(n4591) );
  AND U5445 ( .A(n4594), .B(n4595), .Z(n1831) );
  NAND U5446 ( .A(B[174]), .B(n4596), .Z(n4595) );
  NANDN U5447 ( .A(A[174]), .B(n1833), .Z(n4596) );
  NANDN U5448 ( .A(n1833), .B(A[174]), .Z(n4594) );
  AND U5449 ( .A(n4597), .B(n4598), .Z(n1833) );
  NAND U5450 ( .A(B[173]), .B(n4599), .Z(n4598) );
  NANDN U5451 ( .A(A[173]), .B(n1835), .Z(n4599) );
  NANDN U5452 ( .A(n1835), .B(A[173]), .Z(n4597) );
  AND U5453 ( .A(n4600), .B(n4601), .Z(n1835) );
  NAND U5454 ( .A(B[172]), .B(n4602), .Z(n4601) );
  NANDN U5455 ( .A(A[172]), .B(n1837), .Z(n4602) );
  NANDN U5456 ( .A(n1837), .B(A[172]), .Z(n4600) );
  AND U5457 ( .A(n4603), .B(n4604), .Z(n1837) );
  NAND U5458 ( .A(B[171]), .B(n4605), .Z(n4604) );
  NANDN U5459 ( .A(A[171]), .B(n1839), .Z(n4605) );
  NANDN U5460 ( .A(n1839), .B(A[171]), .Z(n4603) );
  AND U5461 ( .A(n4606), .B(n4607), .Z(n1839) );
  NAND U5462 ( .A(B[170]), .B(n4608), .Z(n4607) );
  NANDN U5463 ( .A(A[170]), .B(n1841), .Z(n4608) );
  NANDN U5464 ( .A(n1841), .B(A[170]), .Z(n4606) );
  AND U5465 ( .A(n4609), .B(n4610), .Z(n1841) );
  NAND U5466 ( .A(B[169]), .B(n4611), .Z(n4610) );
  NANDN U5467 ( .A(A[169]), .B(n1845), .Z(n4611) );
  NANDN U5468 ( .A(n1845), .B(A[169]), .Z(n4609) );
  AND U5469 ( .A(n4612), .B(n4613), .Z(n1845) );
  NAND U5470 ( .A(B[168]), .B(n4614), .Z(n4613) );
  NANDN U5471 ( .A(A[168]), .B(n1847), .Z(n4614) );
  NANDN U5472 ( .A(n1847), .B(A[168]), .Z(n4612) );
  AND U5473 ( .A(n4615), .B(n4616), .Z(n1847) );
  NAND U5474 ( .A(B[167]), .B(n4617), .Z(n4616) );
  NANDN U5475 ( .A(A[167]), .B(n1849), .Z(n4617) );
  NANDN U5476 ( .A(n1849), .B(A[167]), .Z(n4615) );
  AND U5477 ( .A(n4618), .B(n4619), .Z(n1849) );
  NAND U5478 ( .A(B[166]), .B(n4620), .Z(n4619) );
  NANDN U5479 ( .A(A[166]), .B(n1851), .Z(n4620) );
  NANDN U5480 ( .A(n1851), .B(A[166]), .Z(n4618) );
  AND U5481 ( .A(n4621), .B(n4622), .Z(n1851) );
  NAND U5482 ( .A(B[165]), .B(n4623), .Z(n4622) );
  NANDN U5483 ( .A(A[165]), .B(n1853), .Z(n4623) );
  NANDN U5484 ( .A(n1853), .B(A[165]), .Z(n4621) );
  AND U5485 ( .A(n4624), .B(n4625), .Z(n1853) );
  NAND U5486 ( .A(B[164]), .B(n4626), .Z(n4625) );
  NANDN U5487 ( .A(A[164]), .B(n1855), .Z(n4626) );
  NANDN U5488 ( .A(n1855), .B(A[164]), .Z(n4624) );
  AND U5489 ( .A(n4627), .B(n4628), .Z(n1855) );
  NAND U5490 ( .A(B[163]), .B(n4629), .Z(n4628) );
  NANDN U5491 ( .A(A[163]), .B(n1857), .Z(n4629) );
  NANDN U5492 ( .A(n1857), .B(A[163]), .Z(n4627) );
  AND U5493 ( .A(n4630), .B(n4631), .Z(n1857) );
  NAND U5494 ( .A(B[162]), .B(n4632), .Z(n4631) );
  NANDN U5495 ( .A(A[162]), .B(n1859), .Z(n4632) );
  NANDN U5496 ( .A(n1859), .B(A[162]), .Z(n4630) );
  AND U5497 ( .A(n4633), .B(n4634), .Z(n1859) );
  NAND U5498 ( .A(B[161]), .B(n4635), .Z(n4634) );
  NANDN U5499 ( .A(A[161]), .B(n1861), .Z(n4635) );
  NANDN U5500 ( .A(n1861), .B(A[161]), .Z(n4633) );
  AND U5501 ( .A(n4636), .B(n4637), .Z(n1861) );
  NAND U5502 ( .A(B[160]), .B(n4638), .Z(n4637) );
  NANDN U5503 ( .A(A[160]), .B(n1863), .Z(n4638) );
  NANDN U5504 ( .A(n1863), .B(A[160]), .Z(n4636) );
  AND U5505 ( .A(n4639), .B(n4640), .Z(n1863) );
  NAND U5506 ( .A(B[159]), .B(n4641), .Z(n4640) );
  NANDN U5507 ( .A(A[159]), .B(n1867), .Z(n4641) );
  NANDN U5508 ( .A(n1867), .B(A[159]), .Z(n4639) );
  AND U5509 ( .A(n4642), .B(n4643), .Z(n1867) );
  NAND U5510 ( .A(B[158]), .B(n4644), .Z(n4643) );
  NANDN U5511 ( .A(A[158]), .B(n1869), .Z(n4644) );
  NANDN U5512 ( .A(n1869), .B(A[158]), .Z(n4642) );
  AND U5513 ( .A(n4645), .B(n4646), .Z(n1869) );
  NAND U5514 ( .A(B[157]), .B(n4647), .Z(n4646) );
  NANDN U5515 ( .A(A[157]), .B(n1871), .Z(n4647) );
  NANDN U5516 ( .A(n1871), .B(A[157]), .Z(n4645) );
  AND U5517 ( .A(n4648), .B(n4649), .Z(n1871) );
  NAND U5518 ( .A(B[156]), .B(n4650), .Z(n4649) );
  NANDN U5519 ( .A(A[156]), .B(n1873), .Z(n4650) );
  NANDN U5520 ( .A(n1873), .B(A[156]), .Z(n4648) );
  AND U5521 ( .A(n4651), .B(n4652), .Z(n1873) );
  NAND U5522 ( .A(B[155]), .B(n4653), .Z(n4652) );
  NANDN U5523 ( .A(A[155]), .B(n1875), .Z(n4653) );
  NANDN U5524 ( .A(n1875), .B(A[155]), .Z(n4651) );
  AND U5525 ( .A(n4654), .B(n4655), .Z(n1875) );
  NAND U5526 ( .A(B[154]), .B(n4656), .Z(n4655) );
  NANDN U5527 ( .A(A[154]), .B(n1877), .Z(n4656) );
  NANDN U5528 ( .A(n1877), .B(A[154]), .Z(n4654) );
  AND U5529 ( .A(n4657), .B(n4658), .Z(n1877) );
  NAND U5530 ( .A(B[153]), .B(n4659), .Z(n4658) );
  NANDN U5531 ( .A(A[153]), .B(n1879), .Z(n4659) );
  NANDN U5532 ( .A(n1879), .B(A[153]), .Z(n4657) );
  AND U5533 ( .A(n4660), .B(n4661), .Z(n1879) );
  NAND U5534 ( .A(B[152]), .B(n4662), .Z(n4661) );
  NANDN U5535 ( .A(A[152]), .B(n1881), .Z(n4662) );
  NANDN U5536 ( .A(n1881), .B(A[152]), .Z(n4660) );
  AND U5537 ( .A(n4663), .B(n4664), .Z(n1881) );
  NAND U5538 ( .A(B[151]), .B(n4665), .Z(n4664) );
  NANDN U5539 ( .A(A[151]), .B(n1883), .Z(n4665) );
  NANDN U5540 ( .A(n1883), .B(A[151]), .Z(n4663) );
  AND U5541 ( .A(n4666), .B(n4667), .Z(n1883) );
  NAND U5542 ( .A(B[150]), .B(n4668), .Z(n4667) );
  NANDN U5543 ( .A(A[150]), .B(n1885), .Z(n4668) );
  NANDN U5544 ( .A(n1885), .B(A[150]), .Z(n4666) );
  AND U5545 ( .A(n4669), .B(n4670), .Z(n1885) );
  NAND U5546 ( .A(B[149]), .B(n4671), .Z(n4670) );
  NANDN U5547 ( .A(A[149]), .B(n1889), .Z(n4671) );
  NANDN U5548 ( .A(n1889), .B(A[149]), .Z(n4669) );
  AND U5549 ( .A(n4672), .B(n4673), .Z(n1889) );
  NAND U5550 ( .A(B[148]), .B(n4674), .Z(n4673) );
  NANDN U5551 ( .A(A[148]), .B(n1891), .Z(n4674) );
  NANDN U5552 ( .A(n1891), .B(A[148]), .Z(n4672) );
  AND U5553 ( .A(n4675), .B(n4676), .Z(n1891) );
  NAND U5554 ( .A(B[147]), .B(n4677), .Z(n4676) );
  NANDN U5555 ( .A(A[147]), .B(n1893), .Z(n4677) );
  NANDN U5556 ( .A(n1893), .B(A[147]), .Z(n4675) );
  AND U5557 ( .A(n4678), .B(n4679), .Z(n1893) );
  NAND U5558 ( .A(B[146]), .B(n4680), .Z(n4679) );
  NANDN U5559 ( .A(A[146]), .B(n1895), .Z(n4680) );
  NANDN U5560 ( .A(n1895), .B(A[146]), .Z(n4678) );
  AND U5561 ( .A(n4681), .B(n4682), .Z(n1895) );
  NAND U5562 ( .A(B[145]), .B(n4683), .Z(n4682) );
  NANDN U5563 ( .A(A[145]), .B(n1897), .Z(n4683) );
  NANDN U5564 ( .A(n1897), .B(A[145]), .Z(n4681) );
  AND U5565 ( .A(n4684), .B(n4685), .Z(n1897) );
  NAND U5566 ( .A(B[144]), .B(n4686), .Z(n4685) );
  NANDN U5567 ( .A(A[144]), .B(n1899), .Z(n4686) );
  NANDN U5568 ( .A(n1899), .B(A[144]), .Z(n4684) );
  AND U5569 ( .A(n4687), .B(n4688), .Z(n1899) );
  NAND U5570 ( .A(B[143]), .B(n4689), .Z(n4688) );
  NANDN U5571 ( .A(A[143]), .B(n1901), .Z(n4689) );
  NANDN U5572 ( .A(n1901), .B(A[143]), .Z(n4687) );
  AND U5573 ( .A(n4690), .B(n4691), .Z(n1901) );
  NAND U5574 ( .A(B[142]), .B(n4692), .Z(n4691) );
  NANDN U5575 ( .A(A[142]), .B(n1903), .Z(n4692) );
  NANDN U5576 ( .A(n1903), .B(A[142]), .Z(n4690) );
  AND U5577 ( .A(n4693), .B(n4694), .Z(n1903) );
  NAND U5578 ( .A(B[141]), .B(n4695), .Z(n4694) );
  NANDN U5579 ( .A(A[141]), .B(n1905), .Z(n4695) );
  NANDN U5580 ( .A(n1905), .B(A[141]), .Z(n4693) );
  AND U5581 ( .A(n4696), .B(n4697), .Z(n1905) );
  NAND U5582 ( .A(B[140]), .B(n4698), .Z(n4697) );
  NANDN U5583 ( .A(A[140]), .B(n1907), .Z(n4698) );
  NANDN U5584 ( .A(n1907), .B(A[140]), .Z(n4696) );
  AND U5585 ( .A(n4699), .B(n4700), .Z(n1907) );
  NAND U5586 ( .A(B[139]), .B(n4701), .Z(n4700) );
  NANDN U5587 ( .A(A[139]), .B(n1911), .Z(n4701) );
  NANDN U5588 ( .A(n1911), .B(A[139]), .Z(n4699) );
  AND U5589 ( .A(n4702), .B(n4703), .Z(n1911) );
  NAND U5590 ( .A(B[138]), .B(n4704), .Z(n4703) );
  NANDN U5591 ( .A(A[138]), .B(n1913), .Z(n4704) );
  NANDN U5592 ( .A(n1913), .B(A[138]), .Z(n4702) );
  AND U5593 ( .A(n4705), .B(n4706), .Z(n1913) );
  NAND U5594 ( .A(B[137]), .B(n4707), .Z(n4706) );
  NANDN U5595 ( .A(A[137]), .B(n1915), .Z(n4707) );
  NANDN U5596 ( .A(n1915), .B(A[137]), .Z(n4705) );
  AND U5597 ( .A(n4708), .B(n4709), .Z(n1915) );
  NAND U5598 ( .A(B[136]), .B(n4710), .Z(n4709) );
  NANDN U5599 ( .A(A[136]), .B(n1917), .Z(n4710) );
  NANDN U5600 ( .A(n1917), .B(A[136]), .Z(n4708) );
  AND U5601 ( .A(n4711), .B(n4712), .Z(n1917) );
  NAND U5602 ( .A(B[135]), .B(n4713), .Z(n4712) );
  NANDN U5603 ( .A(A[135]), .B(n1919), .Z(n4713) );
  NANDN U5604 ( .A(n1919), .B(A[135]), .Z(n4711) );
  AND U5605 ( .A(n4714), .B(n4715), .Z(n1919) );
  NAND U5606 ( .A(B[134]), .B(n4716), .Z(n4715) );
  NANDN U5607 ( .A(A[134]), .B(n1921), .Z(n4716) );
  NANDN U5608 ( .A(n1921), .B(A[134]), .Z(n4714) );
  AND U5609 ( .A(n4717), .B(n4718), .Z(n1921) );
  NAND U5610 ( .A(B[133]), .B(n4719), .Z(n4718) );
  NANDN U5611 ( .A(A[133]), .B(n1923), .Z(n4719) );
  NANDN U5612 ( .A(n1923), .B(A[133]), .Z(n4717) );
  AND U5613 ( .A(n4720), .B(n4721), .Z(n1923) );
  NAND U5614 ( .A(B[132]), .B(n4722), .Z(n4721) );
  NANDN U5615 ( .A(A[132]), .B(n1925), .Z(n4722) );
  NANDN U5616 ( .A(n1925), .B(A[132]), .Z(n4720) );
  AND U5617 ( .A(n4723), .B(n4724), .Z(n1925) );
  NAND U5618 ( .A(B[131]), .B(n4725), .Z(n4724) );
  NANDN U5619 ( .A(A[131]), .B(n1927), .Z(n4725) );
  NANDN U5620 ( .A(n1927), .B(A[131]), .Z(n4723) );
  AND U5621 ( .A(n4726), .B(n4727), .Z(n1927) );
  NAND U5622 ( .A(B[130]), .B(n4728), .Z(n4727) );
  NANDN U5623 ( .A(A[130]), .B(n1929), .Z(n4728) );
  NANDN U5624 ( .A(n1929), .B(A[130]), .Z(n4726) );
  AND U5625 ( .A(n4729), .B(n4730), .Z(n1929) );
  NAND U5626 ( .A(B[129]), .B(n4731), .Z(n4730) );
  NANDN U5627 ( .A(A[129]), .B(n1933), .Z(n4731) );
  NANDN U5628 ( .A(n1933), .B(A[129]), .Z(n4729) );
  AND U5629 ( .A(n4732), .B(n4733), .Z(n1933) );
  NAND U5630 ( .A(B[128]), .B(n4734), .Z(n4733) );
  NANDN U5631 ( .A(A[128]), .B(n1935), .Z(n4734) );
  NANDN U5632 ( .A(n1935), .B(A[128]), .Z(n4732) );
  AND U5633 ( .A(n4735), .B(n4736), .Z(n1935) );
  NAND U5634 ( .A(B[127]), .B(n4737), .Z(n4736) );
  NANDN U5635 ( .A(A[127]), .B(n1937), .Z(n4737) );
  NANDN U5636 ( .A(n1937), .B(A[127]), .Z(n4735) );
  AND U5637 ( .A(n4738), .B(n4739), .Z(n1937) );
  NAND U5638 ( .A(B[126]), .B(n4740), .Z(n4739) );
  NANDN U5639 ( .A(A[126]), .B(n1939), .Z(n4740) );
  NANDN U5640 ( .A(n1939), .B(A[126]), .Z(n4738) );
  AND U5641 ( .A(n4741), .B(n4742), .Z(n1939) );
  NAND U5642 ( .A(B[125]), .B(n4743), .Z(n4742) );
  NANDN U5643 ( .A(A[125]), .B(n1941), .Z(n4743) );
  NANDN U5644 ( .A(n1941), .B(A[125]), .Z(n4741) );
  AND U5645 ( .A(n4744), .B(n4745), .Z(n1941) );
  NAND U5646 ( .A(B[124]), .B(n4746), .Z(n4745) );
  NANDN U5647 ( .A(A[124]), .B(n1943), .Z(n4746) );
  NANDN U5648 ( .A(n1943), .B(A[124]), .Z(n4744) );
  AND U5649 ( .A(n4747), .B(n4748), .Z(n1943) );
  NAND U5650 ( .A(B[123]), .B(n4749), .Z(n4748) );
  NANDN U5651 ( .A(A[123]), .B(n1945), .Z(n4749) );
  NANDN U5652 ( .A(n1945), .B(A[123]), .Z(n4747) );
  AND U5653 ( .A(n4750), .B(n4751), .Z(n1945) );
  NAND U5654 ( .A(B[122]), .B(n4752), .Z(n4751) );
  NANDN U5655 ( .A(A[122]), .B(n1947), .Z(n4752) );
  NANDN U5656 ( .A(n1947), .B(A[122]), .Z(n4750) );
  AND U5657 ( .A(n4753), .B(n4754), .Z(n1947) );
  NAND U5658 ( .A(B[121]), .B(n4755), .Z(n4754) );
  NANDN U5659 ( .A(A[121]), .B(n1949), .Z(n4755) );
  NANDN U5660 ( .A(n1949), .B(A[121]), .Z(n4753) );
  AND U5661 ( .A(n4756), .B(n4757), .Z(n1949) );
  NAND U5662 ( .A(B[120]), .B(n4758), .Z(n4757) );
  NANDN U5663 ( .A(A[120]), .B(n1951), .Z(n4758) );
  NANDN U5664 ( .A(n1951), .B(A[120]), .Z(n4756) );
  AND U5665 ( .A(n4759), .B(n4760), .Z(n1951) );
  NAND U5666 ( .A(B[119]), .B(n4761), .Z(n4760) );
  NANDN U5667 ( .A(A[119]), .B(n1955), .Z(n4761) );
  NANDN U5668 ( .A(n1955), .B(A[119]), .Z(n4759) );
  AND U5669 ( .A(n4762), .B(n4763), .Z(n1955) );
  NAND U5670 ( .A(B[118]), .B(n4764), .Z(n4763) );
  NANDN U5671 ( .A(A[118]), .B(n1957), .Z(n4764) );
  NANDN U5672 ( .A(n1957), .B(A[118]), .Z(n4762) );
  AND U5673 ( .A(n4765), .B(n4766), .Z(n1957) );
  NAND U5674 ( .A(B[117]), .B(n4767), .Z(n4766) );
  NANDN U5675 ( .A(A[117]), .B(n1959), .Z(n4767) );
  NANDN U5676 ( .A(n1959), .B(A[117]), .Z(n4765) );
  AND U5677 ( .A(n4768), .B(n4769), .Z(n1959) );
  NAND U5678 ( .A(B[116]), .B(n4770), .Z(n4769) );
  NANDN U5679 ( .A(A[116]), .B(n1961), .Z(n4770) );
  NANDN U5680 ( .A(n1961), .B(A[116]), .Z(n4768) );
  AND U5681 ( .A(n4771), .B(n4772), .Z(n1961) );
  NAND U5682 ( .A(B[115]), .B(n4773), .Z(n4772) );
  NANDN U5683 ( .A(A[115]), .B(n1963), .Z(n4773) );
  NANDN U5684 ( .A(n1963), .B(A[115]), .Z(n4771) );
  AND U5685 ( .A(n4774), .B(n4775), .Z(n1963) );
  NAND U5686 ( .A(B[114]), .B(n4776), .Z(n4775) );
  NANDN U5687 ( .A(A[114]), .B(n1965), .Z(n4776) );
  NANDN U5688 ( .A(n1965), .B(A[114]), .Z(n4774) );
  AND U5689 ( .A(n4777), .B(n4778), .Z(n1965) );
  NAND U5690 ( .A(B[113]), .B(n4779), .Z(n4778) );
  NANDN U5691 ( .A(A[113]), .B(n1967), .Z(n4779) );
  NANDN U5692 ( .A(n1967), .B(A[113]), .Z(n4777) );
  AND U5693 ( .A(n4780), .B(n4781), .Z(n1967) );
  NAND U5694 ( .A(B[112]), .B(n4782), .Z(n4781) );
  NANDN U5695 ( .A(A[112]), .B(n1969), .Z(n4782) );
  NANDN U5696 ( .A(n1969), .B(A[112]), .Z(n4780) );
  AND U5697 ( .A(n4783), .B(n4784), .Z(n1969) );
  NAND U5698 ( .A(B[111]), .B(n4785), .Z(n4784) );
  NANDN U5699 ( .A(A[111]), .B(n1971), .Z(n4785) );
  NANDN U5700 ( .A(n1971), .B(A[111]), .Z(n4783) );
  AND U5701 ( .A(n4786), .B(n4787), .Z(n1971) );
  NAND U5702 ( .A(B[110]), .B(n4788), .Z(n4787) );
  NANDN U5703 ( .A(A[110]), .B(n1973), .Z(n4788) );
  NANDN U5704 ( .A(n1973), .B(A[110]), .Z(n4786) );
  AND U5705 ( .A(n4789), .B(n4790), .Z(n1973) );
  NAND U5706 ( .A(B[109]), .B(n4791), .Z(n4790) );
  NANDN U5707 ( .A(A[109]), .B(n1977), .Z(n4791) );
  NANDN U5708 ( .A(n1977), .B(A[109]), .Z(n4789) );
  AND U5709 ( .A(n4792), .B(n4793), .Z(n1977) );
  NAND U5710 ( .A(B[108]), .B(n4794), .Z(n4793) );
  NANDN U5711 ( .A(A[108]), .B(n1979), .Z(n4794) );
  NANDN U5712 ( .A(n1979), .B(A[108]), .Z(n4792) );
  AND U5713 ( .A(n4795), .B(n4796), .Z(n1979) );
  NAND U5714 ( .A(B[107]), .B(n4797), .Z(n4796) );
  NANDN U5715 ( .A(A[107]), .B(n1981), .Z(n4797) );
  NANDN U5716 ( .A(n1981), .B(A[107]), .Z(n4795) );
  AND U5717 ( .A(n4798), .B(n4799), .Z(n1981) );
  NAND U5718 ( .A(B[106]), .B(n4800), .Z(n4799) );
  NANDN U5719 ( .A(A[106]), .B(n1983), .Z(n4800) );
  NANDN U5720 ( .A(n1983), .B(A[106]), .Z(n4798) );
  AND U5721 ( .A(n4801), .B(n4802), .Z(n1983) );
  NAND U5722 ( .A(B[105]), .B(n4803), .Z(n4802) );
  NANDN U5723 ( .A(A[105]), .B(n1985), .Z(n4803) );
  NANDN U5724 ( .A(n1985), .B(A[105]), .Z(n4801) );
  AND U5725 ( .A(n4804), .B(n4805), .Z(n1985) );
  NAND U5726 ( .A(B[104]), .B(n4806), .Z(n4805) );
  NANDN U5727 ( .A(A[104]), .B(n1987), .Z(n4806) );
  NANDN U5728 ( .A(n1987), .B(A[104]), .Z(n4804) );
  AND U5729 ( .A(n4807), .B(n4808), .Z(n1987) );
  NAND U5730 ( .A(B[103]), .B(n4809), .Z(n4808) );
  NANDN U5731 ( .A(A[103]), .B(n1989), .Z(n4809) );
  NANDN U5732 ( .A(n1989), .B(A[103]), .Z(n4807) );
  AND U5733 ( .A(n4810), .B(n4811), .Z(n1989) );
  NAND U5734 ( .A(B[102]), .B(n4812), .Z(n4811) );
  NANDN U5735 ( .A(A[102]), .B(n1991), .Z(n4812) );
  NANDN U5736 ( .A(n1991), .B(A[102]), .Z(n4810) );
  AND U5737 ( .A(n4813), .B(n4814), .Z(n1991) );
  NAND U5738 ( .A(B[101]), .B(n4815), .Z(n4814) );
  NANDN U5739 ( .A(A[101]), .B(n2019), .Z(n4815) );
  NANDN U5740 ( .A(n2019), .B(A[101]), .Z(n4813) );
  AND U5741 ( .A(n4816), .B(n4817), .Z(n2019) );
  NAND U5742 ( .A(B[100]), .B(n4818), .Z(n4817) );
  NANDN U5743 ( .A(A[100]), .B(n2071), .Z(n4818) );
  NANDN U5744 ( .A(n2071), .B(A[100]), .Z(n4816) );
  AND U5745 ( .A(n4819), .B(n4820), .Z(n2071) );
  NAND U5746 ( .A(B[99]), .B(n4821), .Z(n4820) );
  OR U5747 ( .A(n3), .B(A[99]), .Z(n4821) );
  NAND U5748 ( .A(A[99]), .B(n3), .Z(n4819) );
  NAND U5749 ( .A(n4822), .B(n4823), .Z(n3) );
  NAND U5750 ( .A(B[98]), .B(n4824), .Z(n4823) );
  NANDN U5751 ( .A(A[98]), .B(n25), .Z(n4824) );
  NANDN U5752 ( .A(n25), .B(A[98]), .Z(n4822) );
  AND U5753 ( .A(n4825), .B(n4826), .Z(n25) );
  NAND U5754 ( .A(B[97]), .B(n4827), .Z(n4826) );
  NANDN U5755 ( .A(A[97]), .B(n47), .Z(n4827) );
  NANDN U5756 ( .A(n47), .B(A[97]), .Z(n4825) );
  AND U5757 ( .A(n4828), .B(n4829), .Z(n47) );
  NAND U5758 ( .A(B[96]), .B(n4830), .Z(n4829) );
  NANDN U5759 ( .A(A[96]), .B(n69), .Z(n4830) );
  NANDN U5760 ( .A(n69), .B(A[96]), .Z(n4828) );
  AND U5761 ( .A(n4831), .B(n4832), .Z(n69) );
  NAND U5762 ( .A(B[95]), .B(n4833), .Z(n4832) );
  NANDN U5763 ( .A(A[95]), .B(n91), .Z(n4833) );
  NANDN U5764 ( .A(n91), .B(A[95]), .Z(n4831) );
  AND U5765 ( .A(n4834), .B(n4835), .Z(n91) );
  NAND U5766 ( .A(B[94]), .B(n4836), .Z(n4835) );
  NANDN U5767 ( .A(A[94]), .B(n113), .Z(n4836) );
  NANDN U5768 ( .A(n113), .B(A[94]), .Z(n4834) );
  AND U5769 ( .A(n4837), .B(n4838), .Z(n113) );
  NAND U5770 ( .A(B[93]), .B(n4839), .Z(n4838) );
  NANDN U5771 ( .A(A[93]), .B(n135), .Z(n4839) );
  NANDN U5772 ( .A(n135), .B(A[93]), .Z(n4837) );
  AND U5773 ( .A(n4840), .B(n4841), .Z(n135) );
  NAND U5774 ( .A(B[92]), .B(n4842), .Z(n4841) );
  NANDN U5775 ( .A(A[92]), .B(n157), .Z(n4842) );
  NANDN U5776 ( .A(n157), .B(A[92]), .Z(n4840) );
  AND U5777 ( .A(n4843), .B(n4844), .Z(n157) );
  NAND U5778 ( .A(B[91]), .B(n4845), .Z(n4844) );
  NANDN U5779 ( .A(A[91]), .B(n179), .Z(n4845) );
  NANDN U5780 ( .A(n179), .B(A[91]), .Z(n4843) );
  AND U5781 ( .A(n4846), .B(n4847), .Z(n179) );
  NAND U5782 ( .A(B[90]), .B(n4848), .Z(n4847) );
  NANDN U5783 ( .A(A[90]), .B(n201), .Z(n4848) );
  NANDN U5784 ( .A(n201), .B(A[90]), .Z(n4846) );
  AND U5785 ( .A(n4849), .B(n4850), .Z(n201) );
  NAND U5786 ( .A(B[89]), .B(n4851), .Z(n4850) );
  NANDN U5787 ( .A(A[89]), .B(n225), .Z(n4851) );
  NANDN U5788 ( .A(n225), .B(A[89]), .Z(n4849) );
  AND U5789 ( .A(n4852), .B(n4853), .Z(n225) );
  NAND U5790 ( .A(B[88]), .B(n4854), .Z(n4853) );
  NANDN U5791 ( .A(A[88]), .B(n247), .Z(n4854) );
  NANDN U5792 ( .A(n247), .B(A[88]), .Z(n4852) );
  AND U5793 ( .A(n4855), .B(n4856), .Z(n247) );
  NAND U5794 ( .A(B[87]), .B(n4857), .Z(n4856) );
  NANDN U5795 ( .A(A[87]), .B(n269), .Z(n4857) );
  NANDN U5796 ( .A(n269), .B(A[87]), .Z(n4855) );
  AND U5797 ( .A(n4858), .B(n4859), .Z(n269) );
  NAND U5798 ( .A(B[86]), .B(n4860), .Z(n4859) );
  NANDN U5799 ( .A(A[86]), .B(n291), .Z(n4860) );
  NANDN U5800 ( .A(n291), .B(A[86]), .Z(n4858) );
  AND U5801 ( .A(n4861), .B(n4862), .Z(n291) );
  NAND U5802 ( .A(B[85]), .B(n4863), .Z(n4862) );
  NANDN U5803 ( .A(A[85]), .B(n313), .Z(n4863) );
  NANDN U5804 ( .A(n313), .B(A[85]), .Z(n4861) );
  AND U5805 ( .A(n4864), .B(n4865), .Z(n313) );
  NAND U5806 ( .A(B[84]), .B(n4866), .Z(n4865) );
  NANDN U5807 ( .A(A[84]), .B(n335), .Z(n4866) );
  NANDN U5808 ( .A(n335), .B(A[84]), .Z(n4864) );
  AND U5809 ( .A(n4867), .B(n4868), .Z(n335) );
  NAND U5810 ( .A(B[83]), .B(n4869), .Z(n4868) );
  NANDN U5811 ( .A(A[83]), .B(n357), .Z(n4869) );
  NANDN U5812 ( .A(n357), .B(A[83]), .Z(n4867) );
  AND U5813 ( .A(n4870), .B(n4871), .Z(n357) );
  NAND U5814 ( .A(B[82]), .B(n4872), .Z(n4871) );
  NANDN U5815 ( .A(A[82]), .B(n379), .Z(n4872) );
  NANDN U5816 ( .A(n379), .B(A[82]), .Z(n4870) );
  AND U5817 ( .A(n4873), .B(n4874), .Z(n379) );
  NAND U5818 ( .A(B[81]), .B(n4875), .Z(n4874) );
  NANDN U5819 ( .A(A[81]), .B(n401), .Z(n4875) );
  NANDN U5820 ( .A(n401), .B(A[81]), .Z(n4873) );
  AND U5821 ( .A(n4876), .B(n4877), .Z(n401) );
  NAND U5822 ( .A(B[80]), .B(n4878), .Z(n4877) );
  NANDN U5823 ( .A(A[80]), .B(n423), .Z(n4878) );
  NANDN U5824 ( .A(n423), .B(A[80]), .Z(n4876) );
  AND U5825 ( .A(n4879), .B(n4880), .Z(n423) );
  NAND U5826 ( .A(B[79]), .B(n4881), .Z(n4880) );
  NANDN U5827 ( .A(A[79]), .B(n447), .Z(n4881) );
  NANDN U5828 ( .A(n447), .B(A[79]), .Z(n4879) );
  AND U5829 ( .A(n4882), .B(n4883), .Z(n447) );
  NAND U5830 ( .A(B[78]), .B(n4884), .Z(n4883) );
  NANDN U5831 ( .A(A[78]), .B(n469), .Z(n4884) );
  NANDN U5832 ( .A(n469), .B(A[78]), .Z(n4882) );
  AND U5833 ( .A(n4885), .B(n4886), .Z(n469) );
  NAND U5834 ( .A(B[77]), .B(n4887), .Z(n4886) );
  NANDN U5835 ( .A(A[77]), .B(n491), .Z(n4887) );
  NANDN U5836 ( .A(n491), .B(A[77]), .Z(n4885) );
  AND U5837 ( .A(n4888), .B(n4889), .Z(n491) );
  NAND U5838 ( .A(B[76]), .B(n4890), .Z(n4889) );
  NANDN U5839 ( .A(A[76]), .B(n513), .Z(n4890) );
  NANDN U5840 ( .A(n513), .B(A[76]), .Z(n4888) );
  AND U5841 ( .A(n4891), .B(n4892), .Z(n513) );
  NAND U5842 ( .A(B[75]), .B(n4893), .Z(n4892) );
  NANDN U5843 ( .A(A[75]), .B(n535), .Z(n4893) );
  NANDN U5844 ( .A(n535), .B(A[75]), .Z(n4891) );
  AND U5845 ( .A(n4894), .B(n4895), .Z(n535) );
  NAND U5846 ( .A(B[74]), .B(n4896), .Z(n4895) );
  NANDN U5847 ( .A(A[74]), .B(n557), .Z(n4896) );
  NANDN U5848 ( .A(n557), .B(A[74]), .Z(n4894) );
  AND U5849 ( .A(n4897), .B(n4898), .Z(n557) );
  NAND U5850 ( .A(B[73]), .B(n4899), .Z(n4898) );
  NANDN U5851 ( .A(A[73]), .B(n579), .Z(n4899) );
  NANDN U5852 ( .A(n579), .B(A[73]), .Z(n4897) );
  AND U5853 ( .A(n4900), .B(n4901), .Z(n579) );
  NAND U5854 ( .A(B[72]), .B(n4902), .Z(n4901) );
  NANDN U5855 ( .A(A[72]), .B(n601), .Z(n4902) );
  NANDN U5856 ( .A(n601), .B(A[72]), .Z(n4900) );
  AND U5857 ( .A(n4903), .B(n4904), .Z(n601) );
  NAND U5858 ( .A(B[71]), .B(n4905), .Z(n4904) );
  NANDN U5859 ( .A(A[71]), .B(n623), .Z(n4905) );
  NANDN U5860 ( .A(n623), .B(A[71]), .Z(n4903) );
  AND U5861 ( .A(n4906), .B(n4907), .Z(n623) );
  NAND U5862 ( .A(B[70]), .B(n4908), .Z(n4907) );
  NANDN U5863 ( .A(A[70]), .B(n645), .Z(n4908) );
  NANDN U5864 ( .A(n645), .B(A[70]), .Z(n4906) );
  AND U5865 ( .A(n4909), .B(n4910), .Z(n645) );
  NAND U5866 ( .A(B[69]), .B(n4911), .Z(n4910) );
  NANDN U5867 ( .A(A[69]), .B(n669), .Z(n4911) );
  NANDN U5868 ( .A(n669), .B(A[69]), .Z(n4909) );
  AND U5869 ( .A(n4912), .B(n4913), .Z(n669) );
  NAND U5870 ( .A(B[68]), .B(n4914), .Z(n4913) );
  NANDN U5871 ( .A(A[68]), .B(n691), .Z(n4914) );
  NANDN U5872 ( .A(n691), .B(A[68]), .Z(n4912) );
  AND U5873 ( .A(n4915), .B(n4916), .Z(n691) );
  NAND U5874 ( .A(B[67]), .B(n4917), .Z(n4916) );
  NANDN U5875 ( .A(A[67]), .B(n713), .Z(n4917) );
  NANDN U5876 ( .A(n713), .B(A[67]), .Z(n4915) );
  AND U5877 ( .A(n4918), .B(n4919), .Z(n713) );
  NAND U5878 ( .A(B[66]), .B(n4920), .Z(n4919) );
  NANDN U5879 ( .A(A[66]), .B(n735), .Z(n4920) );
  NANDN U5880 ( .A(n735), .B(A[66]), .Z(n4918) );
  AND U5881 ( .A(n4921), .B(n4922), .Z(n735) );
  NAND U5882 ( .A(B[65]), .B(n4923), .Z(n4922) );
  NANDN U5883 ( .A(A[65]), .B(n757), .Z(n4923) );
  NANDN U5884 ( .A(n757), .B(A[65]), .Z(n4921) );
  AND U5885 ( .A(n4924), .B(n4925), .Z(n757) );
  NAND U5886 ( .A(B[64]), .B(n4926), .Z(n4925) );
  NANDN U5887 ( .A(A[64]), .B(n779), .Z(n4926) );
  NANDN U5888 ( .A(n779), .B(A[64]), .Z(n4924) );
  AND U5889 ( .A(n4927), .B(n4928), .Z(n779) );
  NAND U5890 ( .A(B[63]), .B(n4929), .Z(n4928) );
  NANDN U5891 ( .A(A[63]), .B(n801), .Z(n4929) );
  NANDN U5892 ( .A(n801), .B(A[63]), .Z(n4927) );
  AND U5893 ( .A(n4930), .B(n4931), .Z(n801) );
  NAND U5894 ( .A(B[62]), .B(n4932), .Z(n4931) );
  NANDN U5895 ( .A(A[62]), .B(n823), .Z(n4932) );
  NANDN U5896 ( .A(n823), .B(A[62]), .Z(n4930) );
  AND U5897 ( .A(n4933), .B(n4934), .Z(n823) );
  NAND U5898 ( .A(B[61]), .B(n4935), .Z(n4934) );
  NANDN U5899 ( .A(A[61]), .B(n845), .Z(n4935) );
  NANDN U5900 ( .A(n845), .B(A[61]), .Z(n4933) );
  AND U5901 ( .A(n4936), .B(n4937), .Z(n845) );
  NAND U5902 ( .A(B[60]), .B(n4938), .Z(n4937) );
  NANDN U5903 ( .A(A[60]), .B(n867), .Z(n4938) );
  NANDN U5904 ( .A(n867), .B(A[60]), .Z(n4936) );
  AND U5905 ( .A(n4939), .B(n4940), .Z(n867) );
  NAND U5906 ( .A(B[59]), .B(n4941), .Z(n4940) );
  NANDN U5907 ( .A(A[59]), .B(n891), .Z(n4941) );
  NANDN U5908 ( .A(n891), .B(A[59]), .Z(n4939) );
  AND U5909 ( .A(n4942), .B(n4943), .Z(n891) );
  NAND U5910 ( .A(B[58]), .B(n4944), .Z(n4943) );
  NANDN U5911 ( .A(A[58]), .B(n913), .Z(n4944) );
  NANDN U5912 ( .A(n913), .B(A[58]), .Z(n4942) );
  AND U5913 ( .A(n4945), .B(n4946), .Z(n913) );
  NAND U5914 ( .A(B[57]), .B(n4947), .Z(n4946) );
  NANDN U5915 ( .A(A[57]), .B(n935), .Z(n4947) );
  NANDN U5916 ( .A(n935), .B(A[57]), .Z(n4945) );
  AND U5917 ( .A(n4948), .B(n4949), .Z(n935) );
  NAND U5918 ( .A(B[56]), .B(n4950), .Z(n4949) );
  NANDN U5919 ( .A(A[56]), .B(n957), .Z(n4950) );
  NANDN U5920 ( .A(n957), .B(A[56]), .Z(n4948) );
  AND U5921 ( .A(n4951), .B(n4952), .Z(n957) );
  NAND U5922 ( .A(B[55]), .B(n4953), .Z(n4952) );
  NANDN U5923 ( .A(A[55]), .B(n979), .Z(n4953) );
  NANDN U5924 ( .A(n979), .B(A[55]), .Z(n4951) );
  AND U5925 ( .A(n4954), .B(n4955), .Z(n979) );
  NAND U5926 ( .A(B[54]), .B(n4956), .Z(n4955) );
  NANDN U5927 ( .A(A[54]), .B(n1001), .Z(n4956) );
  NANDN U5928 ( .A(n1001), .B(A[54]), .Z(n4954) );
  AND U5929 ( .A(n4957), .B(n4958), .Z(n1001) );
  NAND U5930 ( .A(B[53]), .B(n4959), .Z(n4958) );
  NANDN U5931 ( .A(A[53]), .B(n1023), .Z(n4959) );
  NANDN U5932 ( .A(n1023), .B(A[53]), .Z(n4957) );
  AND U5933 ( .A(n4960), .B(n4961), .Z(n1023) );
  NAND U5934 ( .A(B[52]), .B(n4962), .Z(n4961) );
  NANDN U5935 ( .A(A[52]), .B(n1045), .Z(n4962) );
  NANDN U5936 ( .A(n1045), .B(A[52]), .Z(n4960) );
  AND U5937 ( .A(n4963), .B(n4964), .Z(n1045) );
  NAND U5938 ( .A(B[51]), .B(n4965), .Z(n4964) );
  NANDN U5939 ( .A(A[51]), .B(n1067), .Z(n4965) );
  NANDN U5940 ( .A(n1067), .B(A[51]), .Z(n4963) );
  AND U5941 ( .A(n4966), .B(n4967), .Z(n1067) );
  NAND U5942 ( .A(B[50]), .B(n4968), .Z(n4967) );
  NANDN U5943 ( .A(A[50]), .B(n1089), .Z(n4968) );
  NANDN U5944 ( .A(n1089), .B(A[50]), .Z(n4966) );
  AND U5945 ( .A(n4969), .B(n4970), .Z(n1089) );
  NAND U5946 ( .A(B[49]), .B(n4971), .Z(n4970) );
  NANDN U5947 ( .A(A[49]), .B(n1113), .Z(n4971) );
  NANDN U5948 ( .A(n1113), .B(A[49]), .Z(n4969) );
  AND U5949 ( .A(n4972), .B(n4973), .Z(n1113) );
  NAND U5950 ( .A(B[48]), .B(n4974), .Z(n4973) );
  NANDN U5951 ( .A(A[48]), .B(n1135), .Z(n4974) );
  NANDN U5952 ( .A(n1135), .B(A[48]), .Z(n4972) );
  AND U5953 ( .A(n4975), .B(n4976), .Z(n1135) );
  NAND U5954 ( .A(B[47]), .B(n4977), .Z(n4976) );
  NANDN U5955 ( .A(A[47]), .B(n1157), .Z(n4977) );
  NANDN U5956 ( .A(n1157), .B(A[47]), .Z(n4975) );
  AND U5957 ( .A(n4978), .B(n4979), .Z(n1157) );
  NAND U5958 ( .A(B[46]), .B(n4980), .Z(n4979) );
  NANDN U5959 ( .A(A[46]), .B(n1179), .Z(n4980) );
  NANDN U5960 ( .A(n1179), .B(A[46]), .Z(n4978) );
  AND U5961 ( .A(n4981), .B(n4982), .Z(n1179) );
  NAND U5962 ( .A(B[45]), .B(n4983), .Z(n4982) );
  NANDN U5963 ( .A(A[45]), .B(n1201), .Z(n4983) );
  NANDN U5964 ( .A(n1201), .B(A[45]), .Z(n4981) );
  AND U5965 ( .A(n4984), .B(n4985), .Z(n1201) );
  NAND U5966 ( .A(B[44]), .B(n4986), .Z(n4985) );
  NANDN U5967 ( .A(A[44]), .B(n1223), .Z(n4986) );
  NANDN U5968 ( .A(n1223), .B(A[44]), .Z(n4984) );
  AND U5969 ( .A(n4987), .B(n4988), .Z(n1223) );
  NAND U5970 ( .A(B[43]), .B(n4989), .Z(n4988) );
  NANDN U5971 ( .A(A[43]), .B(n1245), .Z(n4989) );
  NANDN U5972 ( .A(n1245), .B(A[43]), .Z(n4987) );
  AND U5973 ( .A(n4990), .B(n4991), .Z(n1245) );
  NAND U5974 ( .A(B[42]), .B(n4992), .Z(n4991) );
  NANDN U5975 ( .A(A[42]), .B(n1267), .Z(n4992) );
  NANDN U5976 ( .A(n1267), .B(A[42]), .Z(n4990) );
  AND U5977 ( .A(n4993), .B(n4994), .Z(n1267) );
  NAND U5978 ( .A(B[41]), .B(n4995), .Z(n4994) );
  NANDN U5979 ( .A(A[41]), .B(n1289), .Z(n4995) );
  NANDN U5980 ( .A(n1289), .B(A[41]), .Z(n4993) );
  AND U5981 ( .A(n4996), .B(n4997), .Z(n1289) );
  NAND U5982 ( .A(B[40]), .B(n4998), .Z(n4997) );
  NANDN U5983 ( .A(A[40]), .B(n1311), .Z(n4998) );
  NANDN U5984 ( .A(n1311), .B(A[40]), .Z(n4996) );
  AND U5985 ( .A(n4999), .B(n5000), .Z(n1311) );
  NAND U5986 ( .A(B[39]), .B(n5001), .Z(n5000) );
  NANDN U5987 ( .A(A[39]), .B(n1335), .Z(n5001) );
  NANDN U5988 ( .A(n1335), .B(A[39]), .Z(n4999) );
  AND U5989 ( .A(n5002), .B(n5003), .Z(n1335) );
  NAND U5990 ( .A(B[38]), .B(n5004), .Z(n5003) );
  NANDN U5991 ( .A(A[38]), .B(n1357), .Z(n5004) );
  NANDN U5992 ( .A(n1357), .B(A[38]), .Z(n5002) );
  AND U5993 ( .A(n5005), .B(n5006), .Z(n1357) );
  NAND U5994 ( .A(B[37]), .B(n5007), .Z(n5006) );
  NANDN U5995 ( .A(A[37]), .B(n1379), .Z(n5007) );
  NANDN U5996 ( .A(n1379), .B(A[37]), .Z(n5005) );
  AND U5997 ( .A(n5008), .B(n5009), .Z(n1379) );
  NAND U5998 ( .A(B[36]), .B(n5010), .Z(n5009) );
  NANDN U5999 ( .A(A[36]), .B(n1401), .Z(n5010) );
  NANDN U6000 ( .A(n1401), .B(A[36]), .Z(n5008) );
  AND U6001 ( .A(n5011), .B(n5012), .Z(n1401) );
  NAND U6002 ( .A(B[35]), .B(n5013), .Z(n5012) );
  NANDN U6003 ( .A(A[35]), .B(n1423), .Z(n5013) );
  NANDN U6004 ( .A(n1423), .B(A[35]), .Z(n5011) );
  AND U6005 ( .A(n5014), .B(n5015), .Z(n1423) );
  NAND U6006 ( .A(B[34]), .B(n5016), .Z(n5015) );
  NANDN U6007 ( .A(A[34]), .B(n1445), .Z(n5016) );
  NANDN U6008 ( .A(n1445), .B(A[34]), .Z(n5014) );
  AND U6009 ( .A(n5017), .B(n5018), .Z(n1445) );
  NAND U6010 ( .A(B[33]), .B(n5019), .Z(n5018) );
  NANDN U6011 ( .A(A[33]), .B(n1467), .Z(n5019) );
  NANDN U6012 ( .A(n1467), .B(A[33]), .Z(n5017) );
  AND U6013 ( .A(n5020), .B(n5021), .Z(n1467) );
  NAND U6014 ( .A(B[32]), .B(n5022), .Z(n5021) );
  NANDN U6015 ( .A(A[32]), .B(n1489), .Z(n5022) );
  NANDN U6016 ( .A(n1489), .B(A[32]), .Z(n5020) );
  AND U6017 ( .A(n5023), .B(n5024), .Z(n1489) );
  NAND U6018 ( .A(B[31]), .B(n5025), .Z(n5024) );
  NANDN U6019 ( .A(A[31]), .B(n1511), .Z(n5025) );
  NANDN U6020 ( .A(n1511), .B(A[31]), .Z(n5023) );
  AND U6021 ( .A(n5026), .B(n5027), .Z(n1511) );
  NAND U6022 ( .A(B[30]), .B(n5028), .Z(n5027) );
  NANDN U6023 ( .A(A[30]), .B(n1533), .Z(n5028) );
  NANDN U6024 ( .A(n1533), .B(A[30]), .Z(n5026) );
  AND U6025 ( .A(n5029), .B(n5030), .Z(n1533) );
  NAND U6026 ( .A(B[29]), .B(n5031), .Z(n5030) );
  NANDN U6027 ( .A(A[29]), .B(n1557), .Z(n5031) );
  NANDN U6028 ( .A(n1557), .B(A[29]), .Z(n5029) );
  AND U6029 ( .A(n5032), .B(n5033), .Z(n1557) );
  NAND U6030 ( .A(B[28]), .B(n5034), .Z(n5033) );
  NANDN U6031 ( .A(A[28]), .B(n1579), .Z(n5034) );
  NANDN U6032 ( .A(n1579), .B(A[28]), .Z(n5032) );
  AND U6033 ( .A(n5035), .B(n5036), .Z(n1579) );
  NAND U6034 ( .A(B[27]), .B(n5037), .Z(n5036) );
  NANDN U6035 ( .A(A[27]), .B(n1601), .Z(n5037) );
  NANDN U6036 ( .A(n1601), .B(A[27]), .Z(n5035) );
  AND U6037 ( .A(n5038), .B(n5039), .Z(n1601) );
  NAND U6038 ( .A(B[26]), .B(n5040), .Z(n5039) );
  NANDN U6039 ( .A(A[26]), .B(n1623), .Z(n5040) );
  NANDN U6040 ( .A(n1623), .B(A[26]), .Z(n5038) );
  AND U6041 ( .A(n5041), .B(n5042), .Z(n1623) );
  NAND U6042 ( .A(B[25]), .B(n5043), .Z(n5042) );
  NANDN U6043 ( .A(A[25]), .B(n1645), .Z(n5043) );
  NANDN U6044 ( .A(n1645), .B(A[25]), .Z(n5041) );
  AND U6045 ( .A(n5044), .B(n5045), .Z(n1645) );
  NAND U6046 ( .A(B[24]), .B(n5046), .Z(n5045) );
  NANDN U6047 ( .A(A[24]), .B(n1667), .Z(n5046) );
  NANDN U6048 ( .A(n1667), .B(A[24]), .Z(n5044) );
  AND U6049 ( .A(n5047), .B(n5048), .Z(n1667) );
  NAND U6050 ( .A(B[23]), .B(n5049), .Z(n5048) );
  NANDN U6051 ( .A(A[23]), .B(n1689), .Z(n5049) );
  NANDN U6052 ( .A(n1689), .B(A[23]), .Z(n5047) );
  AND U6053 ( .A(n5050), .B(n5051), .Z(n1689) );
  NAND U6054 ( .A(B[22]), .B(n5052), .Z(n5051) );
  NANDN U6055 ( .A(A[22]), .B(n1711), .Z(n5052) );
  NANDN U6056 ( .A(n1711), .B(A[22]), .Z(n5050) );
  AND U6057 ( .A(n5053), .B(n5054), .Z(n1711) );
  NAND U6058 ( .A(B[21]), .B(n5055), .Z(n5054) );
  NANDN U6059 ( .A(A[21]), .B(n1733), .Z(n5055) );
  NANDN U6060 ( .A(n1733), .B(A[21]), .Z(n5053) );
  AND U6061 ( .A(n5056), .B(n5057), .Z(n1733) );
  NAND U6062 ( .A(B[20]), .B(n5058), .Z(n5057) );
  NANDN U6063 ( .A(A[20]), .B(n1755), .Z(n5058) );
  NANDN U6064 ( .A(n1755), .B(A[20]), .Z(n5056) );
  AND U6065 ( .A(n5059), .B(n5060), .Z(n1755) );
  NAND U6066 ( .A(B[19]), .B(n5061), .Z(n5060) );
  NANDN U6067 ( .A(A[19]), .B(n1777), .Z(n5061) );
  NANDN U6068 ( .A(n1777), .B(A[19]), .Z(n5059) );
  AND U6069 ( .A(n5062), .B(n5063), .Z(n1777) );
  NAND U6070 ( .A(B[18]), .B(n5064), .Z(n5063) );
  NANDN U6071 ( .A(A[18]), .B(n1799), .Z(n5064) );
  NANDN U6072 ( .A(n1799), .B(A[18]), .Z(n5062) );
  AND U6073 ( .A(n5065), .B(n5066), .Z(n1799) );
  NAND U6074 ( .A(B[17]), .B(n5067), .Z(n5066) );
  NANDN U6075 ( .A(A[17]), .B(n1821), .Z(n5067) );
  NANDN U6076 ( .A(n1821), .B(A[17]), .Z(n5065) );
  AND U6077 ( .A(n5068), .B(n5069), .Z(n1821) );
  NAND U6078 ( .A(B[16]), .B(n5070), .Z(n5069) );
  NANDN U6079 ( .A(A[16]), .B(n1843), .Z(n5070) );
  NANDN U6080 ( .A(n1843), .B(A[16]), .Z(n5068) );
  AND U6081 ( .A(n5071), .B(n5072), .Z(n1843) );
  NAND U6082 ( .A(B[15]), .B(n5073), .Z(n5072) );
  NANDN U6083 ( .A(A[15]), .B(n1865), .Z(n5073) );
  NANDN U6084 ( .A(n1865), .B(A[15]), .Z(n5071) );
  AND U6085 ( .A(n5074), .B(n5075), .Z(n1865) );
  NAND U6086 ( .A(B[14]), .B(n5076), .Z(n5075) );
  NANDN U6087 ( .A(A[14]), .B(n1887), .Z(n5076) );
  NANDN U6088 ( .A(n1887), .B(A[14]), .Z(n5074) );
  AND U6089 ( .A(n5077), .B(n5078), .Z(n1887) );
  NAND U6090 ( .A(B[13]), .B(n5079), .Z(n5078) );
  NANDN U6091 ( .A(A[13]), .B(n1909), .Z(n5079) );
  NANDN U6092 ( .A(n1909), .B(A[13]), .Z(n5077) );
  AND U6093 ( .A(n5080), .B(n5081), .Z(n1909) );
  NAND U6094 ( .A(B[12]), .B(n5082), .Z(n5081) );
  NANDN U6095 ( .A(A[12]), .B(n1931), .Z(n5082) );
  NANDN U6096 ( .A(n1931), .B(A[12]), .Z(n5080) );
  AND U6097 ( .A(n5083), .B(n5084), .Z(n1931) );
  NAND U6098 ( .A(B[11]), .B(n5085), .Z(n5084) );
  NANDN U6099 ( .A(A[11]), .B(n1953), .Z(n5085) );
  NANDN U6100 ( .A(n1953), .B(A[11]), .Z(n5083) );
  AND U6101 ( .A(n5086), .B(n5087), .Z(n1953) );
  NAND U6102 ( .A(B[10]), .B(n5088), .Z(n5087) );
  NANDN U6103 ( .A(A[10]), .B(n1975), .Z(n5088) );
  NANDN U6104 ( .A(n1975), .B(A[10]), .Z(n5086) );
  AND U6105 ( .A(n5089), .B(n5090), .Z(n1975) );
  NAND U6106 ( .A(B[9]), .B(n5091), .Z(n5090) );
  OR U6107 ( .A(n1), .B(A[9]), .Z(n5091) );
  NAND U6108 ( .A(A[9]), .B(n1), .Z(n5089) );
  NAND U6109 ( .A(n5092), .B(n5093), .Z(n1) );
  NAND U6110 ( .A(B[8]), .B(n5094), .Z(n5093) );
  NANDN U6111 ( .A(A[8]), .B(n223), .Z(n5094) );
  NANDN U6112 ( .A(n223), .B(A[8]), .Z(n5092) );
  AND U6113 ( .A(n5095), .B(n5096), .Z(n223) );
  NAND U6114 ( .A(B[7]), .B(n5097), .Z(n5096) );
  NANDN U6115 ( .A(A[7]), .B(n445), .Z(n5097) );
  NANDN U6116 ( .A(n445), .B(A[7]), .Z(n5095) );
  AND U6117 ( .A(n5098), .B(n5099), .Z(n445) );
  NAND U6118 ( .A(B[6]), .B(n5100), .Z(n5099) );
  NANDN U6119 ( .A(A[6]), .B(n667), .Z(n5100) );
  NANDN U6120 ( .A(n667), .B(A[6]), .Z(n5098) );
  AND U6121 ( .A(n5101), .B(n5102), .Z(n667) );
  NAND U6122 ( .A(B[5]), .B(n5103), .Z(n5102) );
  NANDN U6123 ( .A(A[5]), .B(n889), .Z(n5103) );
  NANDN U6124 ( .A(n889), .B(A[5]), .Z(n5101) );
  AND U6125 ( .A(n5104), .B(n5105), .Z(n889) );
  NAND U6126 ( .A(B[4]), .B(n5106), .Z(n5105) );
  NANDN U6127 ( .A(A[4]), .B(n1111), .Z(n5106) );
  NANDN U6128 ( .A(n1111), .B(A[4]), .Z(n5104) );
  AND U6129 ( .A(n5107), .B(n5108), .Z(n1111) );
  NAND U6130 ( .A(B[3]), .B(n5109), .Z(n5108) );
  NANDN U6131 ( .A(A[3]), .B(n1333), .Z(n5109) );
  NANDN U6132 ( .A(n1333), .B(A[3]), .Z(n5107) );
  AND U6133 ( .A(n5110), .B(n5111), .Z(n1333) );
  NAND U6134 ( .A(B[2]), .B(n5112), .Z(n5111) );
  OR U6135 ( .A(n1555), .B(A[2]), .Z(n5112) );
  NAND U6136 ( .A(A[2]), .B(n1555), .Z(n5110) );
  AND U6137 ( .A(B[1]), .B(A[1]), .Z(n1555) );
endmodule


module modmult_step_N1024 ( xregN_1, y, n, zin, zout );
  input [1023:0] y;
  input [1023:0] n;
  input [1025:0] zin;
  output [1025:0] zout;
  input xregN_1;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74,
         N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88,
         N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101,
         N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112,
         N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, N123,
         N124, N125, N126, N127, N128, N129, N130, N131, N132, N133, N134,
         N135, N136, N137, N138, N139, N140, N141, N142, N143, N144, N145,
         N146, N147, N148, N149, N150, N151, N152, N153, N154, N155, N156,
         N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167,
         N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178,
         N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189,
         N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200,
         N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211,
         N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, N222,
         N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233,
         N234, N235, N236, N237, N238, N239, N240, N241, N242, N243, N244,
         N245, N246, N247, N248, N249, N250, N251, N252, N253, N254, N255,
         N256, N257, N258, N259, N260, N261, N262, N263, N264, N265, N266,
         N267, N268, N269, N270, N271, N272, N273, N274, N275, N276, N277,
         N278, N279, N280, N281, N282, N283, N284, N285, N286, N287, N288,
         N289, N290, N291, N292, N293, N294, N295, N296, N297, N298, N299,
         N300, N301, N302, N303, N304, N305, N306, N307, N308, N309, N310,
         N311, N312, N313, N314, N315, N316, N317, N318, N319, N320, N321,
         N322, N323, N324, N325, N326, N327, N328, N329, N330, N331, N332,
         N333, N334, N335, N336, N337, N338, N339, N340, N341, N342, N343,
         N344, N345, N346, N347, N348, N349, N350, N351, N352, N353, N354,
         N355, N356, N357, N358, N359, N360, N361, N362, N363, N364, N365,
         N366, N367, N368, N369, N370, N371, N372, N373, N374, N375, N376,
         N377, N378, N379, N380, N381, N382, N383, N384, N385, N386, N387,
         N388, N389, N390, N391, N392, N393, N394, N395, N396, N397, N398,
         N399, N400, N401, N402, N403, N404, N405, N406, N407, N408, N409,
         N410, N411, N412, N413, N414, N415, N416, N417, N418, N419, N420,
         N421, N422, N423, N424, N425, N426, N427, N428, N429, N430, N431,
         N432, N433, N434, N435, N436, N437, N438, N439, N440, N441, N442,
         N443, N444, N445, N446, N447, N448, N449, N450, N451, N452, N453,
         N454, N455, N456, N457, N458, N459, N460, N461, N462, N463, N464,
         N465, N466, N467, N468, N469, N470, N471, N472, N473, N474, N475,
         N476, N477, N478, N479, N480, N481, N482, N483, N484, N485, N486,
         N487, N488, N489, N490, N491, N492, N493, N494, N495, N496, N497,
         N498, N499, N500, N501, N502, N503, N504, N505, N506, N507, N508,
         N509, N510, N511, N512, N513, N514, N515, N516, N517, N518, N519,
         N520, N521, N522, N523, N524, N525, N526, N527, N528, N529, N530,
         N531, N532, N533, N534, N535, N536, N537, N538, N539, N540, N541,
         N542, N543, N544, N545, N546, N547, N548, N549, N550, N551, N552,
         N553, N554, N555, N556, N557, N558, N559, N560, N561, N562, N563,
         N564, N565, N566, N567, N568, N569, N570, N571, N572, N573, N574,
         N575, N576, N577, N578, N579, N580, N581, N582, N583, N584, N585,
         N586, N587, N588, N589, N590, N591, N592, N593, N594, N595, N596,
         N597, N598, N599, N600, N601, N602, N603, N604, N605, N606, N607,
         N608, N609, N610, N611, N612, N613, N614, N615, N616, N617, N618,
         N619, N620, N621, N622, N623, N624, N625, N626, N627, N628, N629,
         N630, N631, N632, N633, N634, N635, N636, N637, N638, N639, N640,
         N641, N642, N643, N644, N645, N646, N647, N648, N649, N650, N651,
         N652, N653, N654, N655, N656, N657, N658, N659, N660, N661, N662,
         N663, N664, N665, N666, N667, N668, N669, N670, N671, N672, N673,
         N674, N675, N676, N677, N678, N679, N680, N681, N682, N683, N684,
         N685, N686, N687, N688, N689, N690, N691, N692, N693, N694, N695,
         N696, N697, N698, N699, N700, N701, N702, N703, N704, N705, N706,
         N707, N708, N709, N710, N711, N712, N713, N714, N715, N716, N717,
         N718, N719, N720, N721, N722, N723, N724, N725, N726, N727, N728,
         N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739,
         N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750,
         N751, N752, N753, N754, N755, N756, N757, N758, N759, N760, N761,
         N762, N763, N764, N765, N766, N767, N768, N769, N770, N771, N772,
         N773, N774, N775, N776, N777, N778, N779, N780, N781, N782, N783,
         N784, N785, N786, N787, N788, N789, N790, N791, N792, N793, N794,
         N795, N796, N797, N798, N799, N800, N801, N802, N803, N804, N805,
         N806, N807, N808, N809, N810, N811, N812, N813, N814, N815, N816,
         N817, N818, N819, N820, N821, N822, N823, N824, N825, N826, N827,
         N828, N829, N830, N831, N832, N833, N834, N835, N836, N837, N838,
         N839, N840, N841, N842, N843, N844, N845, N846, N847, N848, N849,
         N850, N851, N852, N853, N854, N855, N856, N857, N858, N859, N860,
         N861, N862, N863, N864, N865, N866, N867, N868, N869, N870, N871,
         N872, N873, N874, N875, N876, N877, N878, N879, N880, N881, N882,
         N883, N884, N885, N886, N887, N888, N889, N890, N891, N892, N893,
         N894, N895, N896, N897, N898, N899, N900, N901, N902, N903, N904,
         N905, N906, N907, N908, N909, N910, N911, N912, N913, N914, N915,
         N916, N917, N918, N919, N920, N921, N922, N923, N924, N925, N926,
         N927, N928, N929, N930, N931, N932, N933, N934, N935, N936, N937,
         N938, N939, N940, N941, N942, N943, N944, N945, N946, N947, N948,
         N949, N950, N951, N952, N953, N954, N955, N956, N957, N958, N959,
         N960, N961, N962, N963, N964, N965, N966, N967, N968, N969, N970,
         N971, N972, N973, N974, N975, N976, N977, N978, N979, N980, N981,
         N982, N983, N984, N985, N986, N987, N988, N989, N990, N991, N992,
         N993, N994, N995, N996, N997, N998, N999, N1000, N1001, N1002, N1003,
         N1004, N1005, N1006, N1007, N1008, N1009, N1010, N1011, N1012, N1013,
         N1014, N1015, N1016, N1017, N1018, N1019, N1020, N1021, N1022, N1023,
         N1024, N1025, N1026, N1027, N1028, N1029, N1030, N1032, N1033, N1034,
         N1035, N1036, N1037, N1038, N1039, N1040, N1041, N1042, N1043, N1044,
         N1045, N1046, N1047, N1048, N1049, N1050, N1051, N1052, N1053, N1054,
         N1055, N1056, N1057, N1058, N1059, N1060, N1061, N1062, N1063, N1064,
         N1065, N1066, N1067, N1068, N1069, N1070, N1071, N1072, N1073, N1074,
         N1075, N1076, N1077, N1078, N1079, N1080, N1081, N1082, N1083, N1084,
         N1085, N1086, N1087, N1088, N1089, N1090, N1091, N1092, N1093, N1094,
         N1095, N1096, N1097, N1098, N1099, N1100, N1101, N1102, N1103, N1104,
         N1105, N1106, N1107, N1108, N1109, N1110, N1111, N1112, N1113, N1114,
         N1115, N1116, N1117, N1118, N1119, N1120, N1121, N1122, N1123, N1124,
         N1125, N1126, N1127, N1128, N1129, N1130, N1131, N1132, N1133, N1134,
         N1135, N1136, N1137, N1138, N1139, N1140, N1141, N1142, N1143, N1144,
         N1145, N1146, N1147, N1148, N1149, N1150, N1151, N1152, N1153, N1154,
         N1155, N1156, N1157, N1158, N1159, N1160, N1161, N1162, N1163, N1164,
         N1165, N1166, N1167, N1168, N1169, N1170, N1171, N1172, N1173, N1174,
         N1175, N1176, N1177, N1178, N1179, N1180, N1181, N1182, N1183, N1184,
         N1185, N1186, N1187, N1188, N1189, N1190, N1191, N1192, N1193, N1194,
         N1195, N1196, N1197, N1198, N1199, N1200, N1201, N1202, N1203, N1204,
         N1205, N1206, N1207, N1208, N1209, N1210, N1211, N1212, N1213, N1214,
         N1215, N1216, N1217, N1218, N1219, N1220, N1221, N1222, N1223, N1224,
         N1225, N1226, N1227, N1228, N1229, N1230, N1231, N1232, N1233, N1234,
         N1235, N1236, N1237, N1238, N1239, N1240, N1241, N1242, N1243, N1244,
         N1245, N1246, N1247, N1248, N1249, N1250, N1251, N1252, N1253, N1254,
         N1255, N1256, N1257, N1258, N1259, N1260, N1261, N1262, N1263, N1264,
         N1265, N1266, N1267, N1268, N1269, N1270, N1271, N1272, N1273, N1274,
         N1275, N1276, N1277, N1278, N1279, N1280, N1281, N1282, N1283, N1284,
         N1285, N1286, N1287, N1288, N1289, N1290, N1291, N1292, N1293, N1294,
         N1295, N1296, N1297, N1298, N1299, N1300, N1301, N1302, N1303, N1304,
         N1305, N1306, N1307, N1308, N1309, N1310, N1311, N1312, N1313, N1314,
         N1315, N1316, N1317, N1318, N1319, N1320, N1321, N1322, N1323, N1324,
         N1325, N1326, N1327, N1328, N1329, N1330, N1331, N1332, N1333, N1334,
         N1335, N1336, N1337, N1338, N1339, N1340, N1341, N1342, N1343, N1344,
         N1345, N1346, N1347, N1348, N1349, N1350, N1351, N1352, N1353, N1354,
         N1355, N1356, N1357, N1358, N1359, N1360, N1361, N1362, N1363, N1364,
         N1365, N1366, N1367, N1368, N1369, N1370, N1371, N1372, N1373, N1374,
         N1375, N1376, N1377, N1378, N1379, N1380, N1381, N1382, N1383, N1384,
         N1385, N1386, N1387, N1388, N1389, N1390, N1391, N1392, N1393, N1394,
         N1395, N1396, N1397, N1398, N1399, N1400, N1401, N1402, N1403, N1404,
         N1405, N1406, N1407, N1408, N1409, N1410, N1411, N1412, N1413, N1414,
         N1415, N1416, N1417, N1418, N1419, N1420, N1421, N1422, N1423, N1424,
         N1425, N1426, N1427, N1428, N1429, N1430, N1431, N1432, N1433, N1434,
         N1435, N1436, N1437, N1438, N1439, N1440, N1441, N1442, N1443, N1444,
         N1445, N1446, N1447, N1448, N1449, N1450, N1451, N1452, N1453, N1454,
         N1455, N1456, N1457, N1458, N1459, N1460, N1461, N1462, N1463, N1464,
         N1465, N1466, N1467, N1468, N1469, N1470, N1471, N1472, N1473, N1474,
         N1475, N1476, N1477, N1478, N1479, N1480, N1481, N1482, N1483, N1484,
         N1485, N1486, N1487, N1488, N1489, N1490, N1491, N1492, N1493, N1494,
         N1495, N1496, N1497, N1498, N1499, N1500, N1501, N1502, N1503, N1504,
         N1505, N1506, N1507, N1508, N1509, N1510, N1511, N1512, N1513, N1514,
         N1515, N1516, N1517, N1518, N1519, N1520, N1521, N1522, N1523, N1524,
         N1525, N1526, N1527, N1528, N1529, N1530, N1531, N1532, N1533, N1534,
         N1535, N1536, N1537, N1538, N1539, N1540, N1541, N1542, N1543, N1544,
         N1545, N1546, N1547, N1548, N1549, N1550, N1551, N1552, N1553, N1554,
         N1555, N1556, N1557, N1558, N1559, N1560, N1561, N1562, N1563, N1564,
         N1565, N1566, N1567, N1568, N1569, N1570, N1571, N1572, N1573, N1574,
         N1575, N1576, N1577, N1578, N1579, N1580, N1581, N1582, N1583, N1584,
         N1585, N1586, N1587, N1588, N1589, N1590, N1591, N1592, N1593, N1594,
         N1595, N1596, N1597, N1598, N1599, N1600, N1601, N1602, N1603, N1604,
         N1605, N1606, N1607, N1608, N1609, N1610, N1611, N1612, N1613, N1614,
         N1615, N1616, N1617, N1618, N1619, N1620, N1621, N1622, N1623, N1624,
         N1625, N1626, N1627, N1628, N1629, N1630, N1631, N1632, N1633, N1634,
         N1635, N1636, N1637, N1638, N1639, N1640, N1641, N1642, N1643, N1644,
         N1645, N1646, N1647, N1648, N1649, N1650, N1651, N1652, N1653, N1654,
         N1655, N1656, N1657, N1658, N1659, N1660, N1661, N1662, N1663, N1664,
         N1665, N1666, N1667, N1668, N1669, N1670, N1671, N1672, N1673, N1674,
         N1675, N1676, N1677, N1678, N1679, N1680, N1681, N1682, N1683, N1684,
         N1685, N1686, N1687, N1688, N1689, N1690, N1691, N1692, N1693, N1694,
         N1695, N1696, N1697, N1698, N1699, N1700, N1701, N1702, N1703, N1704,
         N1705, N1706, N1707, N1708, N1709, N1710, N1711, N1712, N1713, N1714,
         N1715, N1716, N1717, N1718, N1719, N1720, N1721, N1722, N1723, N1724,
         N1725, N1726, N1727, N1728, N1729, N1730, N1731, N1732, N1733, N1734,
         N1735, N1736, N1737, N1738, N1739, N1740, N1741, N1742, N1743, N1744,
         N1745, N1746, N1747, N1748, N1749, N1750, N1751, N1752, N1753, N1754,
         N1755, N1756, N1757, N1758, N1759, N1760, N1761, N1762, N1763, N1764,
         N1765, N1766, N1767, N1768, N1769, N1770, N1771, N1772, N1773, N1774,
         N1775, N1776, N1777, N1778, N1779, N1780, N1781, N1782, N1783, N1784,
         N1785, N1786, N1787, N1788, N1789, N1790, N1791, N1792, N1793, N1794,
         N1795, N1796, N1797, N1798, N1799, N1800, N1801, N1802, N1803, N1804,
         N1805, N1806, N1807, N1808, N1809, N1810, N1811, N1812, N1813, N1814,
         N1815, N1816, N1817, N1818, N1819, N1820, N1821, N1822, N1823, N1824,
         N1825, N1826, N1827, N1828, N1829, N1830, N1831, N1832, N1833, N1834,
         N1835, N1836, N1837, N1838, N1839, N1840, N1841, N1842, N1843, N1844,
         N1845, N1846, N1847, N1848, N1849, N1850, N1851, N1852, N1853, N1854,
         N1855, N1856, N1857, N1858, N1859, N1860, N1861, N1862, N1863, N1864,
         N1865, N1866, N1867, N1868, N1869, N1870, N1871, N1872, N1873, N1874,
         N1875, N1876, N1877, N1878, N1879, N1880, N1881, N1882, N1883, N1884,
         N1885, N1886, N1887, N1888, N1889, N1890, N1891, N1892, N1893, N1894,
         N1895, N1896, N1897, N1898, N1899, N1900, N1901, N1902, N1903, N1904,
         N1905, N1906, N1907, N1908, N1909, N1910, N1911, N1912, N1913, N1914,
         N1915, N1916, N1917, N1918, N1919, N1920, N1921, N1922, N1923, N1924,
         N1925, N1926, N1927, N1928, N1929, N1930, N1931, N1932, N1933, N1934,
         N1935, N1936, N1937, N1938, N1939, N1940, N1941, N1942, N1943, N1944,
         N1945, N1946, N1947, N1948, N1949, N1950, N1951, N1952, N1953, N1954,
         N1955, N1956, N1957, N1958, N1959, N1960, N1961, N1962, N1963, N1964,
         N1965, N1966, N1967, N1968, N1969, N1970, N1971, N1972, N1973, N1974,
         N1975, N1976, N1977, N1978, N1979, N1980, N1981, N1982, N1983, N1984,
         N1985, N1986, N1987, N1988, N1989, N1990, N1991, N1992, N1993, N1994,
         N1995, N1996, N1997, N1998, N1999, N2000, N2001, N2002, N2003, N2004,
         N2005, N2006, N2007, N2008, N2009, N2010, N2011, N2012, N2013, N2014,
         N2015, N2016, N2017, N2018, N2019, N2020, N2021, N2022, N2023, N2024,
         N2025, N2026, N2027, N2028, N2029, N2030, N2031, N2032, N2033, N2034,
         N2035, N2036, N2037, N2038, N2039, N2040, N2041, N2042, N2043, N2044,
         N2045, N2046, N2047, N2048, N2049, N2050, N2051, N2052, N2053, N2054,
         N2055, N2056, N2057, N3084, N3083, N3082, N3081, N3080, N3079, N3078,
         N3077, N3076, N3075, N3074, N3073, N3072, N3071, N3070, N3069, N3068,
         N3067, N3066, N3065, N3064, N3063, N3062, N3061, N3060, N3059, N3058,
         N3057, N3056, N3055, N3054, N3053, N3052, N3051, N3050, N3049, N3048,
         N3047, N3046, N3045, N3044, N3043, N3042, N3041, N3040, N3039, N3038,
         N3037, N3036, N3035, N3034, N3033, N3032, N3031, N3030, N3029, N3028,
         N3027, N3026, N3025, N3024, N3023, N3022, N3021, N3020, N3019, N3018,
         N3017, N3016, N3015, N3014, N3013, N3012, N3011, N3010, N3009, N3008,
         N3007, N3006, N3005, N3004, N3003, N3002, N3001, N3000, N2999, N2998,
         N2997, N2996, N2995, N2994, N2993, N2992, N2991, N2990, N2989, N2988,
         N2987, N2986, N2985, N2984, N2983, N2982, N2981, N2980, N2979, N2978,
         N2977, N2976, N2975, N2974, N2973, N2972, N2971, N2970, N2969, N2968,
         N2967, N2966, N2965, N2964, N2963, N2962, N2961, N2960, N2959, N2958,
         N2957, N2956, N2955, N2954, N2953, N2952, N2951, N2950, N2949, N2948,
         N2947, N2946, N2945, N2944, N2943, N2942, N2941, N2940, N2939, N2938,
         N2937, N2936, N2935, N2934, N2933, N2932, N2931, N2930, N2929, N2928,
         N2927, N2926, N2925, N2924, N2923, N2922, N2921, N2920, N2919, N2918,
         N2917, N2916, N2915, N2914, N2913, N2912, N2911, N2910, N2909, N2908,
         N2907, N2906, N2905, N2904, N2903, N2902, N2901, N2900, N2899, N2898,
         N2897, N2896, N2895, N2894, N2893, N2892, N2891, N2890, N2889, N2888,
         N2887, N2886, N2885, N2884, N2883, N2882, N2881, N2880, N2879, N2878,
         N2877, N2876, N2875, N2874, N2873, N2872, N2871, N2870, N2869, N2868,
         N2867, N2866, N2865, N2864, N2863, N2862, N2861, N2860, N2859, N2858,
         N2857, N2856, N2855, N2854, N2853, N2852, N2851, N2850, N2849, N2848,
         N2847, N2846, N2845, N2844, N2843, N2842, N2841, N2840, N2839, N2838,
         N2837, N2836, N2835, N2834, N2833, N2832, N2831, N2830, N2829, N2828,
         N2827, N2826, N2825, N2824, N2823, N2822, N2821, N2820, N2819, N2818,
         N2817, N2816, N2815, N2814, N2813, N2812, N2811, N2810, N2809, N2808,
         N2807, N2806, N2805, N2804, N2803, N2802, N2801, N2800, N2799, N2798,
         N2797, N2796, N2795, N2794, N2793, N2792, N2791, N2790, N2789, N2788,
         N2787, N2786, N2785, N2784, N2783, N2782, N2781, N2780, N2779, N2778,
         N2777, N2776, N2775, N2774, N2773, N2772, N2771, N2770, N2769, N2768,
         N2767, N2766, N2765, N2764, N2763, N2762, N2761, N2760, N2759, N2758,
         N2757, N2756, N2755, N2754, N2753, N2752, N2751, N2750, N2749, N2748,
         N2747, N2746, N2745, N2744, N2743, N2742, N2741, N2740, N2739, N2738,
         N2737, N2736, N2735, N2734, N2733, N2732, N2731, N2730, N2729, N2728,
         N2727, N2726, N2725, N2724, N2723, N2722, N2721, N2720, N2719, N2718,
         N2717, N2716, N2715, N2714, N2713, N2712, N2711, N2710, N2709, N2708,
         N2707, N2706, N2705, N2704, N2703, N2702, N2701, N2700, N2699, N2698,
         N2697, N2696, N2695, N2694, N2693, N2692, N2691, N2690, N2689, N2688,
         N2687, N2686, N2685, N2684, N2683, N2682, N2681, N2680, N2679, N2678,
         N2677, N2676, N2675, N2674, N2673, N2672, N2671, N2670, N2669, N2668,
         N2667, N2666, N2665, N2664, N2663, N2662, N2661, N2660, N2659, N2658,
         N2657, N2656, N2655, N2654, N2653, N2652, N2651, N2650, N2649, N2648,
         N2647, N2646, N2645, N2644, N2643, N2642, N2641, N2640, N2639, N2638,
         N2637, N2636, N2635, N2634, N2633, N2632, N2631, N2630, N2629, N2628,
         N2627, N2626, N2625, N2624, N2623, N2622, N2621, N2620, N2619, N2618,
         N2617, N2616, N2615, N2614, N2613, N2612, N2611, N2610, N2609, N2608,
         N2607, N2606, N2605, N2604, N2603, N2602, N2601, N2600, N2599, N2598,
         N2597, N2596, N2595, N2594, N2593, N2592, N2591, N2590, N2589, N2588,
         N2587, N2586, N2585, N2584, N2583, N2582, N2581, N2580, N2579, N2578,
         N2577, N2576, N2575, N2574, N2573, N2572, N2571, N2570, N2569, N2568,
         N2567, N2566, N2565, N2564, N2563, N2562, N2561, N2560, N2559, N2558,
         N2557, N2556, N2555, N2554, N2553, N2552, N2551, N2550, N2549, N2548,
         N2547, N2546, N2545, N2544, N2543, N2542, N2541, N2540, N2539, N2538,
         N2537, N2536, N2535, N2534, N2533, N2532, N2531, N2530, N2529, N2528,
         N2527, N2526, N2525, N2524, N2523, N2522, N2521, N2520, N2519, N2518,
         N2517, N2516, N2515, N2514, N2513, N2512, N2511, N2510, N2509, N2508,
         N2507, N2506, N2505, N2504, N2503, N2502, N2501, N2500, N2499, N2498,
         N2497, N2496, N2495, N2494, N2493, N2492, N2491, N2490, N2489, N2488,
         N2487, N2486, N2485, N2484, N2483, N2482, N2481, N2480, N2479, N2478,
         N2477, N2476, N2475, N2474, N2473, N2472, N2471, N2470, N2469, N2468,
         N2467, N2466, N2465, N2464, N2463, N2462, N2461, N2460, N2459, N2458,
         N2457, N2456, N2455, N2454, N2453, N2452, N2451, N2450, N2449, N2448,
         N2447, N2446, N2445, N2444, N2443, N2442, N2441, N2440, N2439, N2438,
         N2437, N2436, N2435, N2434, N2433, N2432, N2431, N2430, N2429, N2428,
         N2427, N2426, N2425, N2424, N2423, N2422, N2421, N2420, N2419, N2418,
         N2417, N2416, N2415, N2414, N2413, N2412, N2411, N2410, N2409, N2408,
         N2407, N2406, N2405, N2404, N2403, N2402, N2401, N2400, N2399, N2398,
         N2397, N2396, N2395, N2394, N2393, N2392, N2391, N2390, N2389, N2388,
         N2387, N2386, N2385, N2384, N2383, N2382, N2381, N2380, N2379, N2378,
         N2377, N2376, N2375, N2374, N2373, N2372, N2371, N2370, N2369, N2368,
         N2367, N2366, N2365, N2364, N2363, N2362, N2361, N2360, N2359, N2358,
         N2357, N2356, N2355, N2354, N2353, N2352, N2351, N2350, N2349, N2348,
         N2347, N2346, N2345, N2344, N2343, N2342, N2341, N2340, N2339, N2338,
         N2337, N2336, N2335, N2334, N2333, N2332, N2331, N2330, N2329, N2328,
         N2327, N2326, N2325, N2324, N2323, N2322, N2321, N2320, N2319, N2318,
         N2317, N2316, N2315, N2314, N2313, N2312, N2311, N2310, N2309, N2308,
         N2307, N2306, N2305, N2304, N2303, N2302, N2301, N2300, N2299, N2298,
         N2297, N2296, N2295, N2294, N2293, N2292, N2291, N2290, N2289, N2288,
         N2287, N2286, N2285, N2284, N2283, N2282, N2281, N2280, N2279, N2278,
         N2277, N2276, N2275, N2274, N2273, N2272, N2271, N2270, N2269, N2268,
         N2267, N2266, N2265, N2264, N2263, N2262, N2261, N2260, N2259, N2258,
         N2257, N2256, N2255, N2254, N2253, N2252, N2251, N2250, N2249, N2248,
         N2247, N2246, N2245, N2244, N2243, N2242, N2241, N2240, N2239, N2238,
         N2237, N2236, N2235, N2234, N2233, N2232, N2231, N2230, N2229, N2228,
         N2227, N2226, N2225, N2224, N2223, N2222, N2221, N2220, N2219, N2218,
         N2217, N2216, N2215, N2214, N2213, N2212, N2211, N2210, N2209, N2208,
         N2207, N2206, N2205, N2204, N2203, N2202, N2201, N2200, N2199, N2198,
         N2197, N2196, N2195, N2194, N2193, N2192, N2191, N2190, N2189, N2188,
         N2187, N2186, N2185, N2184, N2183, N2182, N2181, N2180, N2179, N2178,
         N2177, N2176, N2175, N2174, N2173, N2172, N2171, N2170, N2169, N2168,
         N2167, N2166, N2165, N2164, N2163, N2162, N2161, N2160, N2159, N2158,
         N2157, N2156, N2155, N2154, N2153, N2152, N2151, N2150, N2149, N2148,
         N2147, N2146, N2145, N2144, N2143, N2142, N2141, N2140, N2139, N2138,
         N2137, N2136, N2135, N2134, N2133, N2132, N2131, N2130, N2129, N2128,
         N2127, N2126, N2125, N2124, N2123, N2122, N2121, N2120, N2119, N2118,
         N2117, N2116, N2115, N2114, N2113, N2112, N2111, N2110, N2109, N2108,
         N2107, N2106, N2105, N2104, N2103, N2102, N2101, N2100, N2099, N2098,
         N2097, N2096, N2095, N2094, N2093, N2092, N2091, N2090, N2089, N2088,
         N2087, N2086, N2085, N2084, N2083, N2082, N2081, N2080, N2079, N2078,
         N2077, N2076, N2075, N2074, N2073, N2072, N2071, N2070, N2069, N2068,
         N2067, N2066, N2065, N2064, N2063, N2062, N2061, N2058, n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
         n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
         n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
         n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
         n4110, n4111;
  wire   [1025:0] z2;
  wire   [1025:0] z3;
  wire   SYNOPSYS_UNCONNECTED__0;

  modmult_step_N1024_DW01_sub_0 sub_129_aco ( .A(z3), .B({1'b0, 1'b0, N3084, 
        N3083, N3082, N3081, N3080, N3079, N3078, N3077, N3076, N3075, N3074, 
        N3073, N3072, N3071, N3070, N3069, N3068, N3067, N3066, N3065, N3064, 
        N3063, N3062, N3061, N3060, N3059, N3058, N3057, N3056, N3055, N3054, 
        N3053, N3052, N3051, N3050, N3049, N3048, N3047, N3046, N3045, N3044, 
        N3043, N3042, N3041, N3040, N3039, N3038, N3037, N3036, N3035, N3034, 
        N3033, N3032, N3031, N3030, N3029, N3028, N3027, N3026, N3025, N3024, 
        N3023, N3022, N3021, N3020, N3019, N3018, N3017, N3016, N3015, N3014, 
        N3013, N3012, N3011, N3010, N3009, N3008, N3007, N3006, N3005, N3004, 
        N3003, N3002, N3001, N3000, N2999, N2998, N2997, N2996, N2995, N2994, 
        N2993, N2992, N2991, N2990, N2989, N2988, N2987, N2986, N2985, N2984, 
        N2983, N2982, N2981, N2980, N2979, N2978, N2977, N2976, N2975, N2974, 
        N2973, N2972, N2971, N2970, N2969, N2968, N2967, N2966, N2965, N2964, 
        N2963, N2962, N2961, N2960, N2959, N2958, N2957, N2956, N2955, N2954, 
        N2953, N2952, N2951, N2950, N2949, N2948, N2947, N2946, N2945, N2944, 
        N2943, N2942, N2941, N2940, N2939, N2938, N2937, N2936, N2935, N2934, 
        N2933, N2932, N2931, N2930, N2929, N2928, N2927, N2926, N2925, N2924, 
        N2923, N2922, N2921, N2920, N2919, N2918, N2917, N2916, N2915, N2914, 
        N2913, N2912, N2911, N2910, N2909, N2908, N2907, N2906, N2905, N2904, 
        N2903, N2902, N2901, N2900, N2899, N2898, N2897, N2896, N2895, N2894, 
        N2893, N2892, N2891, N2890, N2889, N2888, N2887, N2886, N2885, N2884, 
        N2883, N2882, N2881, N2880, N2879, N2878, N2877, N2876, N2875, N2874, 
        N2873, N2872, N2871, N2870, N2869, N2868, N2867, N2866, N2865, N2864, 
        N2863, N2862, N2861, N2860, N2859, N2858, N2857, N2856, N2855, N2854, 
        N2853, N2852, N2851, N2850, N2849, N2848, N2847, N2846, N2845, N2844, 
        N2843, N2842, N2841, N2840, N2839, N2838, N2837, N2836, N2835, N2834, 
        N2833, N2832, N2831, N2830, N2829, N2828, N2827, N2826, N2825, N2824, 
        N2823, N2822, N2821, N2820, N2819, N2818, N2817, N2816, N2815, N2814, 
        N2813, N2812, N2811, N2810, N2809, N2808, N2807, N2806, N2805, N2804, 
        N2803, N2802, N2801, N2800, N2799, N2798, N2797, N2796, N2795, N2794, 
        N2793, N2792, N2791, N2790, N2789, N2788, N2787, N2786, N2785, N2784, 
        N2783, N2782, N2781, N2780, N2779, N2778, N2777, N2776, N2775, N2774, 
        N2773, N2772, N2771, N2770, N2769, N2768, N2767, N2766, N2765, N2764, 
        N2763, N2762, N2761, N2760, N2759, N2758, N2757, N2756, N2755, N2754, 
        N2753, N2752, N2751, N2750, N2749, N2748, N2747, N2746, N2745, N2744, 
        N2743, N2742, N2741, N2740, N2739, N2738, N2737, N2736, N2735, N2734, 
        N2733, N2732, N2731, N2730, N2729, N2728, N2727, N2726, N2725, N2724, 
        N2723, N2722, N2721, N2720, N2719, N2718, N2717, N2716, N2715, N2714, 
        N2713, N2712, N2711, N2710, N2709, N2708, N2707, N2706, N2705, N2704, 
        N2703, N2702, N2701, N2700, N2699, N2698, N2697, N2696, N2695, N2694, 
        N2693, N2692, N2691, N2690, N2689, N2688, N2687, N2686, N2685, N2684, 
        N2683, N2682, N2681, N2680, N2679, N2678, N2677, N2676, N2675, N2674, 
        N2673, N2672, N2671, N2670, N2669, N2668, N2667, N2666, N2665, N2664, 
        N2663, N2662, N2661, N2660, N2659, N2658, N2657, N2656, N2655, N2654, 
        N2653, N2652, N2651, N2650, N2649, N2648, N2647, N2646, N2645, N2644, 
        N2643, N2642, N2641, N2640, N2639, N2638, N2637, N2636, N2635, N2634, 
        N2633, N2632, N2631, N2630, N2629, N2628, N2627, N2626, N2625, N2624, 
        N2623, N2622, N2621, N2620, N2619, N2618, N2617, N2616, N2615, N2614, 
        N2613, N2612, N2611, N2610, N2609, N2608, N2607, N2606, N2605, N2604, 
        N2603, N2602, N2601, N2600, N2599, N2598, N2597, N2596, N2595, N2594, 
        N2593, N2592, N2591, N2590, N2589, N2588, N2587, N2586, N2585, N2584, 
        N2583, N2582, N2581, N2580, N2579, N2578, N2577, N2576, N2575, N2574, 
        N2573, N2572, N2571, N2570, N2569, N2568, N2567, N2566, N2565, N2564, 
        N2563, N2562, N2561, N2560, N2559, N2558, N2557, N2556, N2555, N2554, 
        N2553, N2552, N2551, N2550, N2549, N2548, N2547, N2546, N2545, N2544, 
        N2543, N2542, N2541, N2540, N2539, N2538, N2537, N2536, N2535, N2534, 
        N2533, N2532, N2531, N2530, N2529, N2528, N2527, N2526, N2525, N2524, 
        N2523, N2522, N2521, N2520, N2519, N2518, N2517, N2516, N2515, N2514, 
        N2513, N2512, N2511, N2510, N2509, N2508, N2507, N2506, N2505, N2504, 
        N2503, N2502, N2501, N2500, N2499, N2498, N2497, N2496, N2495, N2494, 
        N2493, N2492, N2491, N2490, N2489, N2488, N2487, N2486, N2485, N2484, 
        N2483, N2482, N2481, N2480, N2479, N2478, N2477, N2476, N2475, N2474, 
        N2473, N2472, N2471, N2470, N2469, N2468, N2467, N2466, N2465, N2464, 
        N2463, N2462, N2461, N2460, N2459, N2458, N2457, N2456, N2455, N2454, 
        N2453, N2452, N2451, N2450, N2449, N2448, N2447, N2446, N2445, N2444, 
        N2443, N2442, N2441, N2440, N2439, N2438, N2437, N2436, N2435, N2434, 
        N2433, N2432, N2431, N2430, N2429, N2428, N2427, N2426, N2425, N2424, 
        N2423, N2422, N2421, N2420, N2419, N2418, N2417, N2416, N2415, N2414, 
        N2413, N2412, N2411, N2410, N2409, N2408, N2407, N2406, N2405, N2404, 
        N2403, N2402, N2401, N2400, N2399, N2398, N2397, N2396, N2395, N2394, 
        N2393, N2392, N2391, N2390, N2389, N2388, N2387, N2386, N2385, N2384, 
        N2383, N2382, N2381, N2380, N2379, N2378, N2377, N2376, N2375, N2374, 
        N2373, N2372, N2371, N2370, N2369, N2368, N2367, N2366, N2365, N2364, 
        N2363, N2362, N2361, N2360, N2359, N2358, N2357, N2356, N2355, N2354, 
        N2353, N2352, N2351, N2350, N2349, N2348, N2347, N2346, N2345, N2344, 
        N2343, N2342, N2341, N2340, N2339, N2338, N2337, N2336, N2335, N2334, 
        N2333, N2332, N2331, N2330, N2329, N2328, N2327, N2326, N2325, N2324, 
        N2323, N2322, N2321, N2320, N2319, N2318, N2317, N2316, N2315, N2314, 
        N2313, N2312, N2311, N2310, N2309, N2308, N2307, N2306, N2305, N2304, 
        N2303, N2302, N2301, N2300, N2299, N2298, N2297, N2296, N2295, N2294, 
        N2293, N2292, N2291, N2290, N2289, N2288, N2287, N2286, N2285, N2284, 
        N2283, N2282, N2281, N2280, N2279, N2278, N2277, N2276, N2275, N2274, 
        N2273, N2272, N2271, N2270, N2269, N2268, N2267, N2266, N2265, N2264, 
        N2263, N2262, N2261, N2260, N2259, N2258, N2257, N2256, N2255, N2254, 
        N2253, N2252, N2251, N2250, N2249, N2248, N2247, N2246, N2245, N2244, 
        N2243, N2242, N2241, N2240, N2239, N2238, N2237, N2236, N2235, N2234, 
        N2233, N2232, N2231, N2230, N2229, N2228, N2227, N2226, N2225, N2224, 
        N2223, N2222, N2221, N2220, N2219, N2218, N2217, N2216, N2215, N2214, 
        N2213, N2212, N2211, N2210, N2209, N2208, N2207, N2206, N2205, N2204, 
        N2203, N2202, N2201, N2200, N2199, N2198, N2197, N2196, N2195, N2194, 
        N2193, N2192, N2191, N2190, N2189, N2188, N2187, N2186, N2185, N2184, 
        N2183, N2182, N2181, N2180, N2179, N2178, N2177, N2176, N2175, N2174, 
        N2173, N2172, N2171, N2170, N2169, N2168, N2167, N2166, N2165, N2164, 
        N2163, N2162, N2161, N2160, N2159, N2158, N2157, N2156, N2155, N2154, 
        N2153, N2152, N2151, N2150, N2149, N2148, N2147, N2146, N2145, N2144, 
        N2143, N2142, N2141, N2140, N2139, N2138, N2137, N2136, N2135, N2134, 
        N2133, N2132, N2131, N2130, N2129, N2128, N2127, N2126, N2125, N2124, 
        N2123, N2122, N2121, N2120, N2119, N2118, N2117, N2116, N2115, N2114, 
        N2113, N2112, N2111, N2110, N2109, N2108, N2107, N2106, N2105, N2104, 
        N2103, N2102, N2101, N2100, N2099, N2098, N2097, N2096, N2095, N2094, 
        N2093, N2092, N2091, N2090, N2089, N2088, N2087, N2086, N2085, N2084, 
        N2083, N2082, N2081, N2080, N2079, N2078, N2077, N2076, N2075, N2074, 
        N2073, N2072, N2071, N2070, N2069, N2068, N2067, N2066, N2065, N2064, 
        N2063, N2062, N2061}), .CI(1'b0), .DIFF(zout) );
  modmult_step_N1024_DW02_mult_0 mult_sub_129_aco ( .A(n), .B(N2058), .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__0, N3084, N3083, N3082, N3081, N3080, N3079, 
        N3078, N3077, N3076, N3075, N3074, N3073, N3072, N3071, N3070, N3069, 
        N3068, N3067, N3066, N3065, N3064, N3063, N3062, N3061, N3060, N3059, 
        N3058, N3057, N3056, N3055, N3054, N3053, N3052, N3051, N3050, N3049, 
        N3048, N3047, N3046, N3045, N3044, N3043, N3042, N3041, N3040, N3039, 
        N3038, N3037, N3036, N3035, N3034, N3033, N3032, N3031, N3030, N3029, 
        N3028, N3027, N3026, N3025, N3024, N3023, N3022, N3021, N3020, N3019, 
        N3018, N3017, N3016, N3015, N3014, N3013, N3012, N3011, N3010, N3009, 
        N3008, N3007, N3006, N3005, N3004, N3003, N3002, N3001, N3000, N2999, 
        N2998, N2997, N2996, N2995, N2994, N2993, N2992, N2991, N2990, N2989, 
        N2988, N2987, N2986, N2985, N2984, N2983, N2982, N2981, N2980, N2979, 
        N2978, N2977, N2976, N2975, N2974, N2973, N2972, N2971, N2970, N2969, 
        N2968, N2967, N2966, N2965, N2964, N2963, N2962, N2961, N2960, N2959, 
        N2958, N2957, N2956, N2955, N2954, N2953, N2952, N2951, N2950, N2949, 
        N2948, N2947, N2946, N2945, N2944, N2943, N2942, N2941, N2940, N2939, 
        N2938, N2937, N2936, N2935, N2934, N2933, N2932, N2931, N2930, N2929, 
        N2928, N2927, N2926, N2925, N2924, N2923, N2922, N2921, N2920, N2919, 
        N2918, N2917, N2916, N2915, N2914, N2913, N2912, N2911, N2910, N2909, 
        N2908, N2907, N2906, N2905, N2904, N2903, N2902, N2901, N2900, N2899, 
        N2898, N2897, N2896, N2895, N2894, N2893, N2892, N2891, N2890, N2889, 
        N2888, N2887, N2886, N2885, N2884, N2883, N2882, N2881, N2880, N2879, 
        N2878, N2877, N2876, N2875, N2874, N2873, N2872, N2871, N2870, N2869, 
        N2868, N2867, N2866, N2865, N2864, N2863, N2862, N2861, N2860, N2859, 
        N2858, N2857, N2856, N2855, N2854, N2853, N2852, N2851, N2850, N2849, 
        N2848, N2847, N2846, N2845, N2844, N2843, N2842, N2841, N2840, N2839, 
        N2838, N2837, N2836, N2835, N2834, N2833, N2832, N2831, N2830, N2829, 
        N2828, N2827, N2826, N2825, N2824, N2823, N2822, N2821, N2820, N2819, 
        N2818, N2817, N2816, N2815, N2814, N2813, N2812, N2811, N2810, N2809, 
        N2808, N2807, N2806, N2805, N2804, N2803, N2802, N2801, N2800, N2799, 
        N2798, N2797, N2796, N2795, N2794, N2793, N2792, N2791, N2790, N2789, 
        N2788, N2787, N2786, N2785, N2784, N2783, N2782, N2781, N2780, N2779, 
        N2778, N2777, N2776, N2775, N2774, N2773, N2772, N2771, N2770, N2769, 
        N2768, N2767, N2766, N2765, N2764, N2763, N2762, N2761, N2760, N2759, 
        N2758, N2757, N2756, N2755, N2754, N2753, N2752, N2751, N2750, N2749, 
        N2748, N2747, N2746, N2745, N2744, N2743, N2742, N2741, N2740, N2739, 
        N2738, N2737, N2736, N2735, N2734, N2733, N2732, N2731, N2730, N2729, 
        N2728, N2727, N2726, N2725, N2724, N2723, N2722, N2721, N2720, N2719, 
        N2718, N2717, N2716, N2715, N2714, N2713, N2712, N2711, N2710, N2709, 
        N2708, N2707, N2706, N2705, N2704, N2703, N2702, N2701, N2700, N2699, 
        N2698, N2697, N2696, N2695, N2694, N2693, N2692, N2691, N2690, N2689, 
        N2688, N2687, N2686, N2685, N2684, N2683, N2682, N2681, N2680, N2679, 
        N2678, N2677, N2676, N2675, N2674, N2673, N2672, N2671, N2670, N2669, 
        N2668, N2667, N2666, N2665, N2664, N2663, N2662, N2661, N2660, N2659, 
        N2658, N2657, N2656, N2655, N2654, N2653, N2652, N2651, N2650, N2649, 
        N2648, N2647, N2646, N2645, N2644, N2643, N2642, N2641, N2640, N2639, 
        N2638, N2637, N2636, N2635, N2634, N2633, N2632, N2631, N2630, N2629, 
        N2628, N2627, N2626, N2625, N2624, N2623, N2622, N2621, N2620, N2619, 
        N2618, N2617, N2616, N2615, N2614, N2613, N2612, N2611, N2610, N2609, 
        N2608, N2607, N2606, N2605, N2604, N2603, N2602, N2601, N2600, N2599, 
        N2598, N2597, N2596, N2595, N2594, N2593, N2592, N2591, N2590, N2589, 
        N2588, N2587, N2586, N2585, N2584, N2583, N2582, N2581, N2580, N2579, 
        N2578, N2577, N2576, N2575, N2574, N2573, N2572, N2571, N2570, N2569, 
        N2568, N2567, N2566, N2565, N2564, N2563, N2562, N2561, N2560, N2559, 
        N2558, N2557, N2556, N2555, N2554, N2553, N2552, N2551, N2550, N2549, 
        N2548, N2547, N2546, N2545, N2544, N2543, N2542, N2541, N2540, N2539, 
        N2538, N2537, N2536, N2535, N2534, N2533, N2532, N2531, N2530, N2529, 
        N2528, N2527, N2526, N2525, N2524, N2523, N2522, N2521, N2520, N2519, 
        N2518, N2517, N2516, N2515, N2514, N2513, N2512, N2511, N2510, N2509, 
        N2508, N2507, N2506, N2505, N2504, N2503, N2502, N2501, N2500, N2499, 
        N2498, N2497, N2496, N2495, N2494, N2493, N2492, N2491, N2490, N2489, 
        N2488, N2487, N2486, N2485, N2484, N2483, N2482, N2481, N2480, N2479, 
        N2478, N2477, N2476, N2475, N2474, N2473, N2472, N2471, N2470, N2469, 
        N2468, N2467, N2466, N2465, N2464, N2463, N2462, N2461, N2460, N2459, 
        N2458, N2457, N2456, N2455, N2454, N2453, N2452, N2451, N2450, N2449, 
        N2448, N2447, N2446, N2445, N2444, N2443, N2442, N2441, N2440, N2439, 
        N2438, N2437, N2436, N2435, N2434, N2433, N2432, N2431, N2430, N2429, 
        N2428, N2427, N2426, N2425, N2424, N2423, N2422, N2421, N2420, N2419, 
        N2418, N2417, N2416, N2415, N2414, N2413, N2412, N2411, N2410, N2409, 
        N2408, N2407, N2406, N2405, N2404, N2403, N2402, N2401, N2400, N2399, 
        N2398, N2397, N2396, N2395, N2394, N2393, N2392, N2391, N2390, N2389, 
        N2388, N2387, N2386, N2385, N2384, N2383, N2382, N2381, N2380, N2379, 
        N2378, N2377, N2376, N2375, N2374, N2373, N2372, N2371, N2370, N2369, 
        N2368, N2367, N2366, N2365, N2364, N2363, N2362, N2361, N2360, N2359, 
        N2358, N2357, N2356, N2355, N2354, N2353, N2352, N2351, N2350, N2349, 
        N2348, N2347, N2346, N2345, N2344, N2343, N2342, N2341, N2340, N2339, 
        N2338, N2337, N2336, N2335, N2334, N2333, N2332, N2331, N2330, N2329, 
        N2328, N2327, N2326, N2325, N2324, N2323, N2322, N2321, N2320, N2319, 
        N2318, N2317, N2316, N2315, N2314, N2313, N2312, N2311, N2310, N2309, 
        N2308, N2307, N2306, N2305, N2304, N2303, N2302, N2301, N2300, N2299, 
        N2298, N2297, N2296, N2295, N2294, N2293, N2292, N2291, N2290, N2289, 
        N2288, N2287, N2286, N2285, N2284, N2283, N2282, N2281, N2280, N2279, 
        N2278, N2277, N2276, N2275, N2274, N2273, N2272, N2271, N2270, N2269, 
        N2268, N2267, N2266, N2265, N2264, N2263, N2262, N2261, N2260, N2259, 
        N2258, N2257, N2256, N2255, N2254, N2253, N2252, N2251, N2250, N2249, 
        N2248, N2247, N2246, N2245, N2244, N2243, N2242, N2241, N2240, N2239, 
        N2238, N2237, N2236, N2235, N2234, N2233, N2232, N2231, N2230, N2229, 
        N2228, N2227, N2226, N2225, N2224, N2223, N2222, N2221, N2220, N2219, 
        N2218, N2217, N2216, N2215, N2214, N2213, N2212, N2211, N2210, N2209, 
        N2208, N2207, N2206, N2205, N2204, N2203, N2202, N2201, N2200, N2199, 
        N2198, N2197, N2196, N2195, N2194, N2193, N2192, N2191, N2190, N2189, 
        N2188, N2187, N2186, N2185, N2184, N2183, N2182, N2181, N2180, N2179, 
        N2178, N2177, N2176, N2175, N2174, N2173, N2172, N2171, N2170, N2169, 
        N2168, N2167, N2166, N2165, N2164, N2163, N2162, N2161, N2160, N2159, 
        N2158, N2157, N2156, N2155, N2154, N2153, N2152, N2151, N2150, N2149, 
        N2148, N2147, N2146, N2145, N2144, N2143, N2142, N2141, N2140, N2139, 
        N2138, N2137, N2136, N2135, N2134, N2133, N2132, N2131, N2130, N2129, 
        N2128, N2127, N2126, N2125, N2124, N2123, N2122, N2121, N2120, N2119, 
        N2118, N2117, N2116, N2115, N2114, N2113, N2112, N2111, N2110, N2109, 
        N2108, N2107, N2106, N2105, N2104, N2103, N2102, N2101, N2100, N2099, 
        N2098, N2097, N2096, N2095, N2094, N2093, N2092, N2091, N2090, N2089, 
        N2088, N2087, N2086, N2085, N2084, N2083, N2082, N2081, N2080, N2079, 
        N2078, N2077, N2076, N2075, N2074, N2073, N2072, N2071, N2070, N2069, 
        N2068, N2067, N2066, N2065, N2064, N2063, N2062, N2061}) );
  modmult_step_N1024_DW01_cmp2_0 gte_128 ( .A({1'b0, 1'b0, n}), .B(z3), .LEQ(
        1'b1), .TC(1'b0), .LT_LE(N2058) );
  modmult_step_N1024_DW01_sub_1 sub_124 ( .A(z2), .B({1'b0, 1'b0, n}), .CI(
        1'b0), .DIFF({N2057, N2056, N2055, N2054, N2053, N2052, N2051, N2050, 
        N2049, N2048, N2047, N2046, N2045, N2044, N2043, N2042, N2041, N2040, 
        N2039, N2038, N2037, N2036, N2035, N2034, N2033, N2032, N2031, N2030, 
        N2029, N2028, N2027, N2026, N2025, N2024, N2023, N2022, N2021, N2020, 
        N2019, N2018, N2017, N2016, N2015, N2014, N2013, N2012, N2011, N2010, 
        N2009, N2008, N2007, N2006, N2005, N2004, N2003, N2002, N2001, N2000, 
        N1999, N1998, N1997, N1996, N1995, N1994, N1993, N1992, N1991, N1990, 
        N1989, N1988, N1987, N1986, N1985, N1984, N1983, N1982, N1981, N1980, 
        N1979, N1978, N1977, N1976, N1975, N1974, N1973, N1972, N1971, N1970, 
        N1969, N1968, N1967, N1966, N1965, N1964, N1963, N1962, N1961, N1960, 
        N1959, N1958, N1957, N1956, N1955, N1954, N1953, N1952, N1951, N1950, 
        N1949, N1948, N1947, N1946, N1945, N1944, N1943, N1942, N1941, N1940, 
        N1939, N1938, N1937, N1936, N1935, N1934, N1933, N1932, N1931, N1930, 
        N1929, N1928, N1927, N1926, N1925, N1924, N1923, N1922, N1921, N1920, 
        N1919, N1918, N1917, N1916, N1915, N1914, N1913, N1912, N1911, N1910, 
        N1909, N1908, N1907, N1906, N1905, N1904, N1903, N1902, N1901, N1900, 
        N1899, N1898, N1897, N1896, N1895, N1894, N1893, N1892, N1891, N1890, 
        N1889, N1888, N1887, N1886, N1885, N1884, N1883, N1882, N1881, N1880, 
        N1879, N1878, N1877, N1876, N1875, N1874, N1873, N1872, N1871, N1870, 
        N1869, N1868, N1867, N1866, N1865, N1864, N1863, N1862, N1861, N1860, 
        N1859, N1858, N1857, N1856, N1855, N1854, N1853, N1852, N1851, N1850, 
        N1849, N1848, N1847, N1846, N1845, N1844, N1843, N1842, N1841, N1840, 
        N1839, N1838, N1837, N1836, N1835, N1834, N1833, N1832, N1831, N1830, 
        N1829, N1828, N1827, N1826, N1825, N1824, N1823, N1822, N1821, N1820, 
        N1819, N1818, N1817, N1816, N1815, N1814, N1813, N1812, N1811, N1810, 
        N1809, N1808, N1807, N1806, N1805, N1804, N1803, N1802, N1801, N1800, 
        N1799, N1798, N1797, N1796, N1795, N1794, N1793, N1792, N1791, N1790, 
        N1789, N1788, N1787, N1786, N1785, N1784, N1783, N1782, N1781, N1780, 
        N1779, N1778, N1777, N1776, N1775, N1774, N1773, N1772, N1771, N1770, 
        N1769, N1768, N1767, N1766, N1765, N1764, N1763, N1762, N1761, N1760, 
        N1759, N1758, N1757, N1756, N1755, N1754, N1753, N1752, N1751, N1750, 
        N1749, N1748, N1747, N1746, N1745, N1744, N1743, N1742, N1741, N1740, 
        N1739, N1738, N1737, N1736, N1735, N1734, N1733, N1732, N1731, N1730, 
        N1729, N1728, N1727, N1726, N1725, N1724, N1723, N1722, N1721, N1720, 
        N1719, N1718, N1717, N1716, N1715, N1714, N1713, N1712, N1711, N1710, 
        N1709, N1708, N1707, N1706, N1705, N1704, N1703, N1702, N1701, N1700, 
        N1699, N1698, N1697, N1696, N1695, N1694, N1693, N1692, N1691, N1690, 
        N1689, N1688, N1687, N1686, N1685, N1684, N1683, N1682, N1681, N1680, 
        N1679, N1678, N1677, N1676, N1675, N1674, N1673, N1672, N1671, N1670, 
        N1669, N1668, N1667, N1666, N1665, N1664, N1663, N1662, N1661, N1660, 
        N1659, N1658, N1657, N1656, N1655, N1654, N1653, N1652, N1651, N1650, 
        N1649, N1648, N1647, N1646, N1645, N1644, N1643, N1642, N1641, N1640, 
        N1639, N1638, N1637, N1636, N1635, N1634, N1633, N1632, N1631, N1630, 
        N1629, N1628, N1627, N1626, N1625, N1624, N1623, N1622, N1621, N1620, 
        N1619, N1618, N1617, N1616, N1615, N1614, N1613, N1612, N1611, N1610, 
        N1609, N1608, N1607, N1606, N1605, N1604, N1603, N1602, N1601, N1600, 
        N1599, N1598, N1597, N1596, N1595, N1594, N1593, N1592, N1591, N1590, 
        N1589, N1588, N1587, N1586, N1585, N1584, N1583, N1582, N1581, N1580, 
        N1579, N1578, N1577, N1576, N1575, N1574, N1573, N1572, N1571, N1570, 
        N1569, N1568, N1567, N1566, N1565, N1564, N1563, N1562, N1561, N1560, 
        N1559, N1558, N1557, N1556, N1555, N1554, N1553, N1552, N1551, N1550, 
        N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, 
        N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, 
        N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, 
        N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, 
        N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, 
        N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, 
        N1489, N1488, N1487, N1486, N1485, N1484, N1483, N1482, N1481, N1480, 
        N1479, N1478, N1477, N1476, N1475, N1474, N1473, N1472, N1471, N1470, 
        N1469, N1468, N1467, N1466, N1465, N1464, N1463, N1462, N1461, N1460, 
        N1459, N1458, N1457, N1456, N1455, N1454, N1453, N1452, N1451, N1450, 
        N1449, N1448, N1447, N1446, N1445, N1444, N1443, N1442, N1441, N1440, 
        N1439, N1438, N1437, N1436, N1435, N1434, N1433, N1432, N1431, N1430, 
        N1429, N1428, N1427, N1426, N1425, N1424, N1423, N1422, N1421, N1420, 
        N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, 
        N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, 
        N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, 
        N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, 
        N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, 
        N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, 
        N1359, N1358, N1357, N1356, N1355, N1354, N1353, N1352, N1351, N1350, 
        N1349, N1348, N1347, N1346, N1345, N1344, N1343, N1342, N1341, N1340, 
        N1339, N1338, N1337, N1336, N1335, N1334, N1333, N1332, N1331, N1330, 
        N1329, N1328, N1327, N1326, N1325, N1324, N1323, N1322, N1321, N1320, 
        N1319, N1318, N1317, N1316, N1315, N1314, N1313, N1312, N1311, N1310, 
        N1309, N1308, N1307, N1306, N1305, N1304, N1303, N1302, N1301, N1300, 
        N1299, N1298, N1297, N1296, N1295, N1294, N1293, N1292, N1291, N1290, 
        N1289, N1288, N1287, N1286, N1285, N1284, N1283, N1282, N1281, N1280, 
        N1279, N1278, N1277, N1276, N1275, N1274, N1273, N1272, N1271, N1270, 
        N1269, N1268, N1267, N1266, N1265, N1264, N1263, N1262, N1261, N1260, 
        N1259, N1258, N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250, 
        N1249, N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1240, 
        N1239, N1238, N1237, N1236, N1235, N1234, N1233, N1232, N1231, N1230, 
        N1229, N1228, N1227, N1226, N1225, N1224, N1223, N1222, N1221, N1220, 
        N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, 
        N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, 
        N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, 
        N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, 
        N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, 
        N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161, N1160, 
        N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, 
        N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, 
        N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, 
        N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, 
        N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, 
        N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, 
        N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, 
        N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, 
        N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, 
        N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, 
        N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, 
        N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, 
        N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032}) );
  modmult_step_N1024_DW01_cmp2_1 gt_123 ( .A({1'b0, 1'b0, n}), .B(z2), .LEQ(
        1'b0), .TC(1'b0), .LT_LE(N1030) );
  modmult_step_N1024_DW01_add_0 add_119 ( .A({zin[1024:0], 1'b0}), .B({1'b0, 
        1'b0, y}), .CI(1'b0), .SUM({N1029, N1028, N1027, N1026, N1025, N1024, 
        N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, 
        N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, 
        N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, 
        N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, 
        N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, 
        N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, 
        N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, 
        N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, 
        N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, 
        N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, 
        N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, 
        N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, 
        N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, 
        N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, 
        N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, 
        N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, 
        N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, 
        N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, 
        N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, 
        N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, 
        N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, 
        N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, 
        N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, 
        N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, 
        N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, 
        N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, 
        N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, 
        N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, 
        N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, 
        N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, 
        N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, 
        N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, 
        N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, 
        N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, 
        N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, 
        N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, 
        N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, 
        N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, 
        N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, 
        N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, 
        N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, 
        N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, 
        N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, 
        N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, 
        N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, 
        N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, 
        N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, 
        N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, 
        N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, 
        N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, 
        N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, 
        N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, 
        N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, 
        N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, 
        N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, 
        N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, 
        N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, 
        N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, 
        N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, 
        N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, 
        N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, 
        N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, 
        N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, 
        N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, 
        N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, 
        N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, 
        N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, 
        N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, 
        N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, 
        N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, 
        N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, 
        N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, 
        N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, 
        N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, 
        N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, 
        N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, 
        N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, 
        N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, 
        N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, 
        N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, 
        N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, 
        N6, N5, N4}) );
  NAND U5 ( .A(n1), .B(n2), .Z(z3[9]) );
  NANDN U6 ( .A(N1030), .B(z2[9]), .Z(n2) );
  NANDN U7 ( .A(n3), .B(N1041), .Z(n1) );
  NAND U8 ( .A(n4), .B(n5), .Z(z3[99]) );
  NANDN U9 ( .A(N1030), .B(z2[99]), .Z(n5) );
  NANDN U10 ( .A(n3), .B(N1131), .Z(n4) );
  NAND U11 ( .A(n6), .B(n7), .Z(z3[999]) );
  NANDN U17 ( .A(N1030), .B(z2[999]), .Z(n7) );
  NANDN U18 ( .A(n3), .B(N2031), .Z(n6) );
  NAND U19 ( .A(n8), .B(n9), .Z(z3[998]) );
  NANDN U20 ( .A(N1030), .B(z2[998]), .Z(n9) );
  NANDN U21 ( .A(n3), .B(N2030), .Z(n8) );
  NAND U22 ( .A(n10), .B(n11), .Z(z3[997]) );
  NANDN U23 ( .A(N1030), .B(z2[997]), .Z(n11) );
  NANDN U24 ( .A(n3), .B(N2029), .Z(n10) );
  NAND U25 ( .A(n12), .B(n13), .Z(z3[996]) );
  NANDN U26 ( .A(N1030), .B(z2[996]), .Z(n13) );
  NANDN U27 ( .A(n3), .B(N2028), .Z(n12) );
  NAND U28 ( .A(n14), .B(n23), .Z(z3[995]) );
  NANDN U29 ( .A(N1030), .B(z2[995]), .Z(n23) );
  NANDN U30 ( .A(n3), .B(N2027), .Z(n14) );
  NAND U31 ( .A(n24), .B(n25), .Z(z3[994]) );
  NANDN U32 ( .A(N1030), .B(z2[994]), .Z(n25) );
  NANDN U33 ( .A(n3), .B(N2026), .Z(n24) );
  NAND U34 ( .A(n26), .B(n27), .Z(z3[993]) );
  NANDN U35 ( .A(N1030), .B(z2[993]), .Z(n27) );
  NANDN U36 ( .A(n3), .B(N2025), .Z(n26) );
  NAND U37 ( .A(n28), .B(n29), .Z(z3[992]) );
  NANDN U38 ( .A(N1030), .B(z2[992]), .Z(n29) );
  NANDN U39 ( .A(n3), .B(N2024), .Z(n28) );
  NAND U40 ( .A(n30), .B(n31), .Z(z3[991]) );
  NANDN U41 ( .A(N1030), .B(z2[991]), .Z(n31) );
  NANDN U42 ( .A(n3), .B(N2023), .Z(n30) );
  NAND U43 ( .A(n32), .B(n33), .Z(z3[990]) );
  NANDN U44 ( .A(N1030), .B(z2[990]), .Z(n33) );
  NANDN U45 ( .A(n3), .B(N2022), .Z(n32) );
  NAND U46 ( .A(n34), .B(n35), .Z(z3[98]) );
  NANDN U47 ( .A(N1030), .B(z2[98]), .Z(n35) );
  NANDN U48 ( .A(n3), .B(N1130), .Z(n34) );
  NAND U49 ( .A(n36), .B(n37), .Z(z3[989]) );
  NANDN U50 ( .A(N1030), .B(z2[989]), .Z(n37) );
  NANDN U51 ( .A(n3), .B(N2021), .Z(n36) );
  NAND U52 ( .A(n38), .B(n39), .Z(z3[988]) );
  NANDN U53 ( .A(N1030), .B(z2[988]), .Z(n39) );
  NANDN U54 ( .A(n3), .B(N2020), .Z(n38) );
  NAND U55 ( .A(n40), .B(n41), .Z(z3[987]) );
  NANDN U56 ( .A(N1030), .B(z2[987]), .Z(n41) );
  NANDN U57 ( .A(n3), .B(N2019), .Z(n40) );
  NAND U58 ( .A(n42), .B(n43), .Z(z3[986]) );
  NANDN U59 ( .A(N1030), .B(z2[986]), .Z(n43) );
  NANDN U60 ( .A(n3), .B(N2018), .Z(n42) );
  NAND U61 ( .A(n44), .B(n45), .Z(z3[985]) );
  NANDN U62 ( .A(N1030), .B(z2[985]), .Z(n45) );
  NANDN U63 ( .A(n3), .B(N2017), .Z(n44) );
  NAND U64 ( .A(n46), .B(n47), .Z(z3[984]) );
  NANDN U65 ( .A(N1030), .B(z2[984]), .Z(n47) );
  NANDN U66 ( .A(n3), .B(N2016), .Z(n46) );
  NAND U67 ( .A(n48), .B(n49), .Z(z3[983]) );
  NANDN U68 ( .A(N1030), .B(z2[983]), .Z(n49) );
  NANDN U69 ( .A(n3), .B(N2015), .Z(n48) );
  NAND U70 ( .A(n50), .B(n51), .Z(z3[982]) );
  NANDN U71 ( .A(N1030), .B(z2[982]), .Z(n51) );
  NANDN U72 ( .A(n3), .B(N2014), .Z(n50) );
  NAND U73 ( .A(n52), .B(n53), .Z(z3[981]) );
  NANDN U74 ( .A(N1030), .B(z2[981]), .Z(n53) );
  NANDN U75 ( .A(n3), .B(N2013), .Z(n52) );
  NAND U76 ( .A(n54), .B(n55), .Z(z3[980]) );
  NANDN U77 ( .A(N1030), .B(z2[980]), .Z(n55) );
  NANDN U78 ( .A(n3), .B(N2012), .Z(n54) );
  NAND U79 ( .A(n56), .B(n57), .Z(z3[97]) );
  NANDN U80 ( .A(N1030), .B(z2[97]), .Z(n57) );
  NANDN U81 ( .A(n3), .B(N1129), .Z(n56) );
  NAND U82 ( .A(n58), .B(n59), .Z(z3[979]) );
  NANDN U83 ( .A(N1030), .B(z2[979]), .Z(n59) );
  NANDN U84 ( .A(n3), .B(N2011), .Z(n58) );
  NAND U85 ( .A(n60), .B(n61), .Z(z3[978]) );
  NANDN U86 ( .A(N1030), .B(z2[978]), .Z(n61) );
  NANDN U87 ( .A(n3), .B(N2010), .Z(n60) );
  NAND U88 ( .A(n62), .B(n63), .Z(z3[977]) );
  NANDN U89 ( .A(N1030), .B(z2[977]), .Z(n63) );
  NANDN U90 ( .A(n3), .B(N2009), .Z(n62) );
  NAND U91 ( .A(n64), .B(n65), .Z(z3[976]) );
  NANDN U92 ( .A(N1030), .B(z2[976]), .Z(n65) );
  NANDN U93 ( .A(n3), .B(N2008), .Z(n64) );
  NAND U94 ( .A(n66), .B(n67), .Z(z3[975]) );
  NANDN U95 ( .A(N1030), .B(z2[975]), .Z(n67) );
  NANDN U96 ( .A(n3), .B(N2007), .Z(n66) );
  NAND U97 ( .A(n68), .B(n69), .Z(z3[974]) );
  NANDN U98 ( .A(N1030), .B(z2[974]), .Z(n69) );
  NANDN U99 ( .A(n3), .B(N2006), .Z(n68) );
  NAND U100 ( .A(n70), .B(n71), .Z(z3[973]) );
  NANDN U101 ( .A(N1030), .B(z2[973]), .Z(n71) );
  NANDN U102 ( .A(n3), .B(N2005), .Z(n70) );
  NAND U103 ( .A(n72), .B(n73), .Z(z3[972]) );
  NANDN U104 ( .A(N1030), .B(z2[972]), .Z(n73) );
  NANDN U105 ( .A(n3), .B(N2004), .Z(n72) );
  NAND U106 ( .A(n74), .B(n75), .Z(z3[971]) );
  NANDN U107 ( .A(N1030), .B(z2[971]), .Z(n75) );
  NANDN U108 ( .A(n3), .B(N2003), .Z(n74) );
  NAND U109 ( .A(n76), .B(n77), .Z(z3[970]) );
  NANDN U110 ( .A(N1030), .B(z2[970]), .Z(n77) );
  NANDN U111 ( .A(n3), .B(N2002), .Z(n76) );
  NAND U112 ( .A(n78), .B(n79), .Z(z3[96]) );
  NANDN U113 ( .A(N1030), .B(z2[96]), .Z(n79) );
  NANDN U114 ( .A(n3), .B(N1128), .Z(n78) );
  NAND U115 ( .A(n80), .B(n81), .Z(z3[969]) );
  NANDN U116 ( .A(N1030), .B(z2[969]), .Z(n81) );
  NANDN U117 ( .A(n3), .B(N2001), .Z(n80) );
  NAND U118 ( .A(n82), .B(n83), .Z(z3[968]) );
  NANDN U119 ( .A(N1030), .B(z2[968]), .Z(n83) );
  NANDN U120 ( .A(n3), .B(N2000), .Z(n82) );
  NAND U121 ( .A(n84), .B(n85), .Z(z3[967]) );
  NANDN U122 ( .A(N1030), .B(z2[967]), .Z(n85) );
  NANDN U123 ( .A(n3), .B(N1999), .Z(n84) );
  NAND U124 ( .A(n86), .B(n87), .Z(z3[966]) );
  NANDN U125 ( .A(N1030), .B(z2[966]), .Z(n87) );
  NANDN U126 ( .A(n3), .B(N1998), .Z(n86) );
  NAND U127 ( .A(n88), .B(n89), .Z(z3[965]) );
  NANDN U128 ( .A(N1030), .B(z2[965]), .Z(n89) );
  NANDN U129 ( .A(n3), .B(N1997), .Z(n88) );
  NAND U130 ( .A(n90), .B(n91), .Z(z3[964]) );
  NANDN U131 ( .A(N1030), .B(z2[964]), .Z(n91) );
  NANDN U132 ( .A(n3), .B(N1996), .Z(n90) );
  NAND U133 ( .A(n92), .B(n93), .Z(z3[963]) );
  NANDN U134 ( .A(N1030), .B(z2[963]), .Z(n93) );
  NANDN U135 ( .A(n3), .B(N1995), .Z(n92) );
  NAND U136 ( .A(n94), .B(n95), .Z(z3[962]) );
  NANDN U137 ( .A(N1030), .B(z2[962]), .Z(n95) );
  NANDN U138 ( .A(n3), .B(N1994), .Z(n94) );
  NAND U139 ( .A(n96), .B(n97), .Z(z3[961]) );
  NANDN U140 ( .A(N1030), .B(z2[961]), .Z(n97) );
  NANDN U141 ( .A(n3), .B(N1993), .Z(n96) );
  NAND U142 ( .A(n98), .B(n99), .Z(z3[960]) );
  NANDN U143 ( .A(N1030), .B(z2[960]), .Z(n99) );
  NANDN U144 ( .A(n3), .B(N1992), .Z(n98) );
  NAND U145 ( .A(n100), .B(n101), .Z(z3[95]) );
  NANDN U146 ( .A(N1030), .B(z2[95]), .Z(n101) );
  NANDN U147 ( .A(n3), .B(N1127), .Z(n100) );
  NAND U148 ( .A(n102), .B(n103), .Z(z3[959]) );
  NANDN U149 ( .A(N1030), .B(z2[959]), .Z(n103) );
  NANDN U150 ( .A(n3), .B(N1991), .Z(n102) );
  NAND U151 ( .A(n104), .B(n105), .Z(z3[958]) );
  NANDN U152 ( .A(N1030), .B(z2[958]), .Z(n105) );
  NANDN U153 ( .A(n3), .B(N1990), .Z(n104) );
  NAND U154 ( .A(n106), .B(n107), .Z(z3[957]) );
  NANDN U155 ( .A(N1030), .B(z2[957]), .Z(n107) );
  NANDN U156 ( .A(n3), .B(N1989), .Z(n106) );
  NAND U157 ( .A(n108), .B(n109), .Z(z3[956]) );
  NANDN U158 ( .A(N1030), .B(z2[956]), .Z(n109) );
  NANDN U159 ( .A(n3), .B(N1988), .Z(n108) );
  NAND U160 ( .A(n110), .B(n111), .Z(z3[955]) );
  NANDN U161 ( .A(N1030), .B(z2[955]), .Z(n111) );
  NANDN U162 ( .A(n3), .B(N1987), .Z(n110) );
  NAND U163 ( .A(n112), .B(n113), .Z(z3[954]) );
  NANDN U164 ( .A(N1030), .B(z2[954]), .Z(n113) );
  NANDN U165 ( .A(n3), .B(N1986), .Z(n112) );
  NAND U166 ( .A(n114), .B(n115), .Z(z3[953]) );
  NANDN U167 ( .A(N1030), .B(z2[953]), .Z(n115) );
  NANDN U168 ( .A(n3), .B(N1985), .Z(n114) );
  NAND U169 ( .A(n116), .B(n117), .Z(z3[952]) );
  NANDN U170 ( .A(N1030), .B(z2[952]), .Z(n117) );
  NANDN U171 ( .A(n3), .B(N1984), .Z(n116) );
  NAND U172 ( .A(n118), .B(n119), .Z(z3[951]) );
  NANDN U173 ( .A(N1030), .B(z2[951]), .Z(n119) );
  NANDN U174 ( .A(n3), .B(N1983), .Z(n118) );
  NAND U175 ( .A(n120), .B(n121), .Z(z3[950]) );
  NANDN U176 ( .A(N1030), .B(z2[950]), .Z(n121) );
  NANDN U177 ( .A(n3), .B(N1982), .Z(n120) );
  NAND U178 ( .A(n122), .B(n123), .Z(z3[94]) );
  NANDN U179 ( .A(N1030), .B(z2[94]), .Z(n123) );
  NANDN U180 ( .A(n3), .B(N1126), .Z(n122) );
  NAND U181 ( .A(n124), .B(n125), .Z(z3[949]) );
  NANDN U182 ( .A(N1030), .B(z2[949]), .Z(n125) );
  NANDN U183 ( .A(n3), .B(N1981), .Z(n124) );
  NAND U184 ( .A(n126), .B(n127), .Z(z3[948]) );
  NANDN U185 ( .A(N1030), .B(z2[948]), .Z(n127) );
  NANDN U186 ( .A(n3), .B(N1980), .Z(n126) );
  NAND U187 ( .A(n128), .B(n129), .Z(z3[947]) );
  NANDN U188 ( .A(N1030), .B(z2[947]), .Z(n129) );
  NANDN U189 ( .A(n3), .B(N1979), .Z(n128) );
  NAND U190 ( .A(n130), .B(n131), .Z(z3[946]) );
  NANDN U191 ( .A(N1030), .B(z2[946]), .Z(n131) );
  NANDN U192 ( .A(n3), .B(N1978), .Z(n130) );
  NAND U193 ( .A(n132), .B(n133), .Z(z3[945]) );
  NANDN U194 ( .A(N1030), .B(z2[945]), .Z(n133) );
  NANDN U195 ( .A(n3), .B(N1977), .Z(n132) );
  NAND U196 ( .A(n134), .B(n135), .Z(z3[944]) );
  NANDN U197 ( .A(N1030), .B(z2[944]), .Z(n135) );
  NANDN U198 ( .A(n3), .B(N1976), .Z(n134) );
  NAND U199 ( .A(n136), .B(n137), .Z(z3[943]) );
  NANDN U200 ( .A(N1030), .B(z2[943]), .Z(n137) );
  NANDN U201 ( .A(n3), .B(N1975), .Z(n136) );
  NAND U202 ( .A(n138), .B(n139), .Z(z3[942]) );
  NANDN U203 ( .A(N1030), .B(z2[942]), .Z(n139) );
  NANDN U204 ( .A(n3), .B(N1974), .Z(n138) );
  NAND U205 ( .A(n140), .B(n141), .Z(z3[941]) );
  NANDN U206 ( .A(N1030), .B(z2[941]), .Z(n141) );
  NANDN U207 ( .A(n3), .B(N1973), .Z(n140) );
  NAND U208 ( .A(n142), .B(n143), .Z(z3[940]) );
  NANDN U209 ( .A(N1030), .B(z2[940]), .Z(n143) );
  NANDN U210 ( .A(n3), .B(N1972), .Z(n142) );
  NAND U211 ( .A(n144), .B(n145), .Z(z3[93]) );
  NANDN U212 ( .A(N1030), .B(z2[93]), .Z(n145) );
  NANDN U213 ( .A(n3), .B(N1125), .Z(n144) );
  NAND U214 ( .A(n146), .B(n147), .Z(z3[939]) );
  NANDN U215 ( .A(N1030), .B(z2[939]), .Z(n147) );
  NANDN U216 ( .A(n3), .B(N1971), .Z(n146) );
  NAND U217 ( .A(n148), .B(n149), .Z(z3[938]) );
  NANDN U218 ( .A(N1030), .B(z2[938]), .Z(n149) );
  NANDN U219 ( .A(n3), .B(N1970), .Z(n148) );
  NAND U220 ( .A(n150), .B(n151), .Z(z3[937]) );
  NANDN U221 ( .A(N1030), .B(z2[937]), .Z(n151) );
  NANDN U222 ( .A(n3), .B(N1969), .Z(n150) );
  NAND U223 ( .A(n152), .B(n153), .Z(z3[936]) );
  NANDN U224 ( .A(N1030), .B(z2[936]), .Z(n153) );
  NANDN U225 ( .A(n3), .B(N1968), .Z(n152) );
  NAND U226 ( .A(n154), .B(n155), .Z(z3[935]) );
  NANDN U227 ( .A(N1030), .B(z2[935]), .Z(n155) );
  NANDN U228 ( .A(n3), .B(N1967), .Z(n154) );
  NAND U229 ( .A(n156), .B(n157), .Z(z3[934]) );
  NANDN U230 ( .A(N1030), .B(z2[934]), .Z(n157) );
  NANDN U231 ( .A(n3), .B(N1966), .Z(n156) );
  NAND U232 ( .A(n158), .B(n159), .Z(z3[933]) );
  NANDN U233 ( .A(N1030), .B(z2[933]), .Z(n159) );
  NANDN U234 ( .A(n3), .B(N1965), .Z(n158) );
  NAND U235 ( .A(n160), .B(n161), .Z(z3[932]) );
  NANDN U236 ( .A(N1030), .B(z2[932]), .Z(n161) );
  NANDN U237 ( .A(n3), .B(N1964), .Z(n160) );
  NAND U238 ( .A(n162), .B(n163), .Z(z3[931]) );
  NANDN U239 ( .A(N1030), .B(z2[931]), .Z(n163) );
  NANDN U240 ( .A(n3), .B(N1963), .Z(n162) );
  NAND U241 ( .A(n164), .B(n165), .Z(z3[930]) );
  NANDN U242 ( .A(N1030), .B(z2[930]), .Z(n165) );
  NANDN U243 ( .A(n3), .B(N1962), .Z(n164) );
  NAND U244 ( .A(n166), .B(n167), .Z(z3[92]) );
  NANDN U245 ( .A(N1030), .B(z2[92]), .Z(n167) );
  NANDN U246 ( .A(n3), .B(N1124), .Z(n166) );
  NAND U247 ( .A(n168), .B(n169), .Z(z3[929]) );
  NANDN U248 ( .A(N1030), .B(z2[929]), .Z(n169) );
  NANDN U249 ( .A(n3), .B(N1961), .Z(n168) );
  NAND U250 ( .A(n170), .B(n171), .Z(z3[928]) );
  NANDN U251 ( .A(N1030), .B(z2[928]), .Z(n171) );
  NANDN U252 ( .A(n3), .B(N1960), .Z(n170) );
  NAND U253 ( .A(n172), .B(n173), .Z(z3[927]) );
  NANDN U254 ( .A(N1030), .B(z2[927]), .Z(n173) );
  NANDN U255 ( .A(n3), .B(N1959), .Z(n172) );
  NAND U256 ( .A(n174), .B(n175), .Z(z3[926]) );
  NANDN U257 ( .A(N1030), .B(z2[926]), .Z(n175) );
  NANDN U258 ( .A(n3), .B(N1958), .Z(n174) );
  NAND U259 ( .A(n176), .B(n177), .Z(z3[925]) );
  NANDN U260 ( .A(N1030), .B(z2[925]), .Z(n177) );
  NANDN U261 ( .A(n3), .B(N1957), .Z(n176) );
  NAND U262 ( .A(n178), .B(n179), .Z(z3[924]) );
  NANDN U263 ( .A(N1030), .B(z2[924]), .Z(n179) );
  NANDN U264 ( .A(n3), .B(N1956), .Z(n178) );
  NAND U265 ( .A(n180), .B(n181), .Z(z3[923]) );
  NANDN U266 ( .A(N1030), .B(z2[923]), .Z(n181) );
  NANDN U267 ( .A(n3), .B(N1955), .Z(n180) );
  NAND U268 ( .A(n182), .B(n183), .Z(z3[922]) );
  NANDN U269 ( .A(N1030), .B(z2[922]), .Z(n183) );
  NANDN U270 ( .A(n3), .B(N1954), .Z(n182) );
  NAND U271 ( .A(n184), .B(n185), .Z(z3[921]) );
  NANDN U272 ( .A(N1030), .B(z2[921]), .Z(n185) );
  NANDN U273 ( .A(n3), .B(N1953), .Z(n184) );
  NAND U274 ( .A(n186), .B(n187), .Z(z3[920]) );
  NANDN U275 ( .A(N1030), .B(z2[920]), .Z(n187) );
  NANDN U276 ( .A(n3), .B(N1952), .Z(n186) );
  NAND U277 ( .A(n188), .B(n189), .Z(z3[91]) );
  NANDN U278 ( .A(N1030), .B(z2[91]), .Z(n189) );
  NANDN U279 ( .A(n3), .B(N1123), .Z(n188) );
  NAND U280 ( .A(n190), .B(n191), .Z(z3[919]) );
  NANDN U281 ( .A(N1030), .B(z2[919]), .Z(n191) );
  NANDN U282 ( .A(n3), .B(N1951), .Z(n190) );
  NAND U283 ( .A(n192), .B(n193), .Z(z3[918]) );
  NANDN U284 ( .A(N1030), .B(z2[918]), .Z(n193) );
  NANDN U285 ( .A(n3), .B(N1950), .Z(n192) );
  NAND U286 ( .A(n194), .B(n195), .Z(z3[917]) );
  NANDN U287 ( .A(N1030), .B(z2[917]), .Z(n195) );
  NANDN U288 ( .A(n3), .B(N1949), .Z(n194) );
  NAND U289 ( .A(n196), .B(n197), .Z(z3[916]) );
  NANDN U290 ( .A(N1030), .B(z2[916]), .Z(n197) );
  NANDN U291 ( .A(n3), .B(N1948), .Z(n196) );
  NAND U292 ( .A(n198), .B(n199), .Z(z3[915]) );
  NANDN U293 ( .A(N1030), .B(z2[915]), .Z(n199) );
  NANDN U294 ( .A(n3), .B(N1947), .Z(n198) );
  NAND U295 ( .A(n200), .B(n201), .Z(z3[914]) );
  NANDN U296 ( .A(N1030), .B(z2[914]), .Z(n201) );
  NANDN U297 ( .A(n3), .B(N1946), .Z(n200) );
  NAND U298 ( .A(n202), .B(n203), .Z(z3[913]) );
  NANDN U299 ( .A(N1030), .B(z2[913]), .Z(n203) );
  NANDN U300 ( .A(n3), .B(N1945), .Z(n202) );
  NAND U301 ( .A(n204), .B(n205), .Z(z3[912]) );
  NANDN U302 ( .A(N1030), .B(z2[912]), .Z(n205) );
  NANDN U303 ( .A(n3), .B(N1944), .Z(n204) );
  NAND U304 ( .A(n206), .B(n207), .Z(z3[911]) );
  NANDN U305 ( .A(N1030), .B(z2[911]), .Z(n207) );
  NANDN U306 ( .A(n3), .B(N1943), .Z(n206) );
  NAND U307 ( .A(n208), .B(n209), .Z(z3[910]) );
  NANDN U308 ( .A(N1030), .B(z2[910]), .Z(n209) );
  NANDN U309 ( .A(n3), .B(N1942), .Z(n208) );
  NAND U310 ( .A(n210), .B(n211), .Z(z3[90]) );
  NANDN U311 ( .A(N1030), .B(z2[90]), .Z(n211) );
  NANDN U312 ( .A(n3), .B(N1122), .Z(n210) );
  NAND U313 ( .A(n212), .B(n213), .Z(z3[909]) );
  NANDN U314 ( .A(N1030), .B(z2[909]), .Z(n213) );
  NANDN U315 ( .A(n3), .B(N1941), .Z(n212) );
  NAND U316 ( .A(n214), .B(n215), .Z(z3[908]) );
  NANDN U317 ( .A(N1030), .B(z2[908]), .Z(n215) );
  NANDN U318 ( .A(n3), .B(N1940), .Z(n214) );
  NAND U319 ( .A(n216), .B(n217), .Z(z3[907]) );
  NANDN U320 ( .A(N1030), .B(z2[907]), .Z(n217) );
  NANDN U321 ( .A(n3), .B(N1939), .Z(n216) );
  NAND U322 ( .A(n218), .B(n219), .Z(z3[906]) );
  NANDN U323 ( .A(N1030), .B(z2[906]), .Z(n219) );
  NANDN U324 ( .A(n3), .B(N1938), .Z(n218) );
  NAND U325 ( .A(n220), .B(n221), .Z(z3[905]) );
  NANDN U326 ( .A(N1030), .B(z2[905]), .Z(n221) );
  NANDN U327 ( .A(n3), .B(N1937), .Z(n220) );
  NAND U328 ( .A(n222), .B(n223), .Z(z3[904]) );
  NANDN U329 ( .A(N1030), .B(z2[904]), .Z(n223) );
  NANDN U330 ( .A(n3), .B(N1936), .Z(n222) );
  NAND U331 ( .A(n224), .B(n225), .Z(z3[903]) );
  NANDN U332 ( .A(N1030), .B(z2[903]), .Z(n225) );
  NANDN U333 ( .A(n3), .B(N1935), .Z(n224) );
  NAND U334 ( .A(n226), .B(n227), .Z(z3[902]) );
  NANDN U335 ( .A(N1030), .B(z2[902]), .Z(n227) );
  NANDN U336 ( .A(n3), .B(N1934), .Z(n226) );
  NAND U337 ( .A(n228), .B(n229), .Z(z3[901]) );
  NANDN U338 ( .A(N1030), .B(z2[901]), .Z(n229) );
  NANDN U339 ( .A(n3), .B(N1933), .Z(n228) );
  NAND U340 ( .A(n230), .B(n231), .Z(z3[900]) );
  NANDN U341 ( .A(N1030), .B(z2[900]), .Z(n231) );
  NANDN U342 ( .A(n3), .B(N1932), .Z(n230) );
  NAND U343 ( .A(n232), .B(n233), .Z(z3[8]) );
  NANDN U344 ( .A(N1030), .B(z2[8]), .Z(n233) );
  NANDN U345 ( .A(n3), .B(N1040), .Z(n232) );
  NAND U346 ( .A(n234), .B(n235), .Z(z3[89]) );
  NANDN U347 ( .A(N1030), .B(z2[89]), .Z(n235) );
  NANDN U348 ( .A(n3), .B(N1121), .Z(n234) );
  NAND U349 ( .A(n236), .B(n237), .Z(z3[899]) );
  NANDN U350 ( .A(N1030), .B(z2[899]), .Z(n237) );
  NANDN U351 ( .A(n3), .B(N1931), .Z(n236) );
  NAND U352 ( .A(n238), .B(n239), .Z(z3[898]) );
  NANDN U353 ( .A(N1030), .B(z2[898]), .Z(n239) );
  NANDN U354 ( .A(n3), .B(N1930), .Z(n238) );
  NAND U355 ( .A(n240), .B(n241), .Z(z3[897]) );
  NANDN U356 ( .A(N1030), .B(z2[897]), .Z(n241) );
  NANDN U357 ( .A(n3), .B(N1929), .Z(n240) );
  NAND U358 ( .A(n242), .B(n243), .Z(z3[896]) );
  NANDN U359 ( .A(N1030), .B(z2[896]), .Z(n243) );
  NANDN U360 ( .A(n3), .B(N1928), .Z(n242) );
  NAND U361 ( .A(n244), .B(n245), .Z(z3[895]) );
  NANDN U362 ( .A(N1030), .B(z2[895]), .Z(n245) );
  NANDN U363 ( .A(n3), .B(N1927), .Z(n244) );
  NAND U364 ( .A(n246), .B(n247), .Z(z3[894]) );
  NANDN U365 ( .A(N1030), .B(z2[894]), .Z(n247) );
  NANDN U366 ( .A(n3), .B(N1926), .Z(n246) );
  NAND U367 ( .A(n248), .B(n249), .Z(z3[893]) );
  NANDN U368 ( .A(N1030), .B(z2[893]), .Z(n249) );
  NANDN U369 ( .A(n3), .B(N1925), .Z(n248) );
  NAND U370 ( .A(n250), .B(n251), .Z(z3[892]) );
  NANDN U371 ( .A(N1030), .B(z2[892]), .Z(n251) );
  NANDN U372 ( .A(n3), .B(N1924), .Z(n250) );
  NAND U373 ( .A(n252), .B(n253), .Z(z3[891]) );
  NANDN U374 ( .A(N1030), .B(z2[891]), .Z(n253) );
  NANDN U375 ( .A(n3), .B(N1923), .Z(n252) );
  NAND U376 ( .A(n254), .B(n255), .Z(z3[890]) );
  NANDN U377 ( .A(N1030), .B(z2[890]), .Z(n255) );
  NANDN U378 ( .A(n3), .B(N1922), .Z(n254) );
  NAND U379 ( .A(n256), .B(n257), .Z(z3[88]) );
  NANDN U380 ( .A(N1030), .B(z2[88]), .Z(n257) );
  NANDN U381 ( .A(n3), .B(N1120), .Z(n256) );
  NAND U382 ( .A(n258), .B(n259), .Z(z3[889]) );
  NANDN U383 ( .A(N1030), .B(z2[889]), .Z(n259) );
  NANDN U384 ( .A(n3), .B(N1921), .Z(n258) );
  NAND U385 ( .A(n260), .B(n261), .Z(z3[888]) );
  NANDN U386 ( .A(N1030), .B(z2[888]), .Z(n261) );
  NANDN U387 ( .A(n3), .B(N1920), .Z(n260) );
  NAND U388 ( .A(n262), .B(n263), .Z(z3[887]) );
  NANDN U389 ( .A(N1030), .B(z2[887]), .Z(n263) );
  NANDN U390 ( .A(n3), .B(N1919), .Z(n262) );
  NAND U391 ( .A(n264), .B(n265), .Z(z3[886]) );
  NANDN U392 ( .A(N1030), .B(z2[886]), .Z(n265) );
  NANDN U393 ( .A(n3), .B(N1918), .Z(n264) );
  NAND U394 ( .A(n266), .B(n267), .Z(z3[885]) );
  NANDN U395 ( .A(N1030), .B(z2[885]), .Z(n267) );
  NANDN U396 ( .A(n3), .B(N1917), .Z(n266) );
  NAND U397 ( .A(n268), .B(n269), .Z(z3[884]) );
  NANDN U398 ( .A(N1030), .B(z2[884]), .Z(n269) );
  NANDN U399 ( .A(n3), .B(N1916), .Z(n268) );
  NAND U400 ( .A(n270), .B(n271), .Z(z3[883]) );
  NANDN U401 ( .A(N1030), .B(z2[883]), .Z(n271) );
  NANDN U402 ( .A(n3), .B(N1915), .Z(n270) );
  NAND U403 ( .A(n272), .B(n273), .Z(z3[882]) );
  NANDN U404 ( .A(N1030), .B(z2[882]), .Z(n273) );
  NANDN U405 ( .A(n3), .B(N1914), .Z(n272) );
  NAND U406 ( .A(n274), .B(n275), .Z(z3[881]) );
  NANDN U407 ( .A(N1030), .B(z2[881]), .Z(n275) );
  NANDN U408 ( .A(n3), .B(N1913), .Z(n274) );
  NAND U409 ( .A(n276), .B(n277), .Z(z3[880]) );
  NANDN U410 ( .A(N1030), .B(z2[880]), .Z(n277) );
  NANDN U411 ( .A(n3), .B(N1912), .Z(n276) );
  NAND U412 ( .A(n278), .B(n279), .Z(z3[87]) );
  NANDN U413 ( .A(N1030), .B(z2[87]), .Z(n279) );
  NANDN U414 ( .A(n3), .B(N1119), .Z(n278) );
  NAND U415 ( .A(n280), .B(n281), .Z(z3[879]) );
  NANDN U416 ( .A(N1030), .B(z2[879]), .Z(n281) );
  NANDN U417 ( .A(n3), .B(N1911), .Z(n280) );
  NAND U418 ( .A(n282), .B(n283), .Z(z3[878]) );
  NANDN U419 ( .A(N1030), .B(z2[878]), .Z(n283) );
  NANDN U420 ( .A(n3), .B(N1910), .Z(n282) );
  NAND U421 ( .A(n284), .B(n285), .Z(z3[877]) );
  NANDN U422 ( .A(N1030), .B(z2[877]), .Z(n285) );
  NANDN U423 ( .A(n3), .B(N1909), .Z(n284) );
  NAND U424 ( .A(n286), .B(n287), .Z(z3[876]) );
  NANDN U425 ( .A(N1030), .B(z2[876]), .Z(n287) );
  NANDN U426 ( .A(n3), .B(N1908), .Z(n286) );
  NAND U427 ( .A(n288), .B(n289), .Z(z3[875]) );
  NANDN U428 ( .A(N1030), .B(z2[875]), .Z(n289) );
  NANDN U429 ( .A(n3), .B(N1907), .Z(n288) );
  NAND U430 ( .A(n290), .B(n291), .Z(z3[874]) );
  NANDN U431 ( .A(N1030), .B(z2[874]), .Z(n291) );
  NANDN U432 ( .A(n3), .B(N1906), .Z(n290) );
  NAND U433 ( .A(n292), .B(n293), .Z(z3[873]) );
  NANDN U434 ( .A(N1030), .B(z2[873]), .Z(n293) );
  NANDN U435 ( .A(n3), .B(N1905), .Z(n292) );
  NAND U436 ( .A(n294), .B(n295), .Z(z3[872]) );
  NANDN U437 ( .A(N1030), .B(z2[872]), .Z(n295) );
  NANDN U438 ( .A(n3), .B(N1904), .Z(n294) );
  NAND U439 ( .A(n296), .B(n297), .Z(z3[871]) );
  NANDN U440 ( .A(N1030), .B(z2[871]), .Z(n297) );
  NANDN U441 ( .A(n3), .B(N1903), .Z(n296) );
  NAND U442 ( .A(n298), .B(n299), .Z(z3[870]) );
  NANDN U443 ( .A(N1030), .B(z2[870]), .Z(n299) );
  NANDN U444 ( .A(n3), .B(N1902), .Z(n298) );
  NAND U445 ( .A(n300), .B(n301), .Z(z3[86]) );
  NANDN U446 ( .A(N1030), .B(z2[86]), .Z(n301) );
  NANDN U447 ( .A(n3), .B(N1118), .Z(n300) );
  NAND U448 ( .A(n302), .B(n303), .Z(z3[869]) );
  NANDN U449 ( .A(N1030), .B(z2[869]), .Z(n303) );
  NANDN U450 ( .A(n3), .B(N1901), .Z(n302) );
  NAND U451 ( .A(n304), .B(n305), .Z(z3[868]) );
  NANDN U452 ( .A(N1030), .B(z2[868]), .Z(n305) );
  NANDN U453 ( .A(n3), .B(N1900), .Z(n304) );
  NAND U454 ( .A(n306), .B(n307), .Z(z3[867]) );
  NANDN U455 ( .A(N1030), .B(z2[867]), .Z(n307) );
  NANDN U456 ( .A(n3), .B(N1899), .Z(n306) );
  NAND U457 ( .A(n308), .B(n309), .Z(z3[866]) );
  NANDN U458 ( .A(N1030), .B(z2[866]), .Z(n309) );
  NANDN U459 ( .A(n3), .B(N1898), .Z(n308) );
  NAND U460 ( .A(n310), .B(n311), .Z(z3[865]) );
  NANDN U461 ( .A(N1030), .B(z2[865]), .Z(n311) );
  NANDN U462 ( .A(n3), .B(N1897), .Z(n310) );
  NAND U463 ( .A(n312), .B(n313), .Z(z3[864]) );
  NANDN U464 ( .A(N1030), .B(z2[864]), .Z(n313) );
  NANDN U465 ( .A(n3), .B(N1896), .Z(n312) );
  NAND U466 ( .A(n314), .B(n315), .Z(z3[863]) );
  NANDN U467 ( .A(N1030), .B(z2[863]), .Z(n315) );
  NANDN U468 ( .A(n3), .B(N1895), .Z(n314) );
  NAND U469 ( .A(n316), .B(n317), .Z(z3[862]) );
  NANDN U470 ( .A(N1030), .B(z2[862]), .Z(n317) );
  NANDN U471 ( .A(n3), .B(N1894), .Z(n316) );
  NAND U472 ( .A(n318), .B(n319), .Z(z3[861]) );
  NANDN U473 ( .A(N1030), .B(z2[861]), .Z(n319) );
  NANDN U474 ( .A(n3), .B(N1893), .Z(n318) );
  NAND U475 ( .A(n320), .B(n321), .Z(z3[860]) );
  NANDN U476 ( .A(N1030), .B(z2[860]), .Z(n321) );
  NANDN U477 ( .A(n3), .B(N1892), .Z(n320) );
  NAND U478 ( .A(n322), .B(n323), .Z(z3[85]) );
  NANDN U479 ( .A(N1030), .B(z2[85]), .Z(n323) );
  NANDN U480 ( .A(n3), .B(N1117), .Z(n322) );
  NAND U481 ( .A(n324), .B(n325), .Z(z3[859]) );
  NANDN U482 ( .A(N1030), .B(z2[859]), .Z(n325) );
  NANDN U483 ( .A(n3), .B(N1891), .Z(n324) );
  NAND U484 ( .A(n326), .B(n327), .Z(z3[858]) );
  NANDN U485 ( .A(N1030), .B(z2[858]), .Z(n327) );
  NANDN U486 ( .A(n3), .B(N1890), .Z(n326) );
  NAND U487 ( .A(n328), .B(n329), .Z(z3[857]) );
  NANDN U488 ( .A(N1030), .B(z2[857]), .Z(n329) );
  NANDN U489 ( .A(n3), .B(N1889), .Z(n328) );
  NAND U490 ( .A(n330), .B(n331), .Z(z3[856]) );
  NANDN U491 ( .A(N1030), .B(z2[856]), .Z(n331) );
  NANDN U492 ( .A(n3), .B(N1888), .Z(n330) );
  NAND U493 ( .A(n332), .B(n333), .Z(z3[855]) );
  NANDN U494 ( .A(N1030), .B(z2[855]), .Z(n333) );
  NANDN U495 ( .A(n3), .B(N1887), .Z(n332) );
  NAND U496 ( .A(n334), .B(n335), .Z(z3[854]) );
  NANDN U497 ( .A(N1030), .B(z2[854]), .Z(n335) );
  NANDN U498 ( .A(n3), .B(N1886), .Z(n334) );
  NAND U499 ( .A(n336), .B(n337), .Z(z3[853]) );
  NANDN U500 ( .A(N1030), .B(z2[853]), .Z(n337) );
  NANDN U501 ( .A(n3), .B(N1885), .Z(n336) );
  NAND U502 ( .A(n338), .B(n339), .Z(z3[852]) );
  NANDN U503 ( .A(N1030), .B(z2[852]), .Z(n339) );
  NANDN U504 ( .A(n3), .B(N1884), .Z(n338) );
  NAND U505 ( .A(n340), .B(n341), .Z(z3[851]) );
  NANDN U506 ( .A(N1030), .B(z2[851]), .Z(n341) );
  NANDN U507 ( .A(n3), .B(N1883), .Z(n340) );
  NAND U508 ( .A(n342), .B(n343), .Z(z3[850]) );
  NANDN U509 ( .A(N1030), .B(z2[850]), .Z(n343) );
  NANDN U510 ( .A(n3), .B(N1882), .Z(n342) );
  NAND U511 ( .A(n344), .B(n345), .Z(z3[84]) );
  NANDN U512 ( .A(N1030), .B(z2[84]), .Z(n345) );
  NANDN U513 ( .A(n3), .B(N1116), .Z(n344) );
  NAND U514 ( .A(n346), .B(n347), .Z(z3[849]) );
  NANDN U515 ( .A(N1030), .B(z2[849]), .Z(n347) );
  NANDN U516 ( .A(n3), .B(N1881), .Z(n346) );
  NAND U517 ( .A(n348), .B(n349), .Z(z3[848]) );
  NANDN U518 ( .A(N1030), .B(z2[848]), .Z(n349) );
  NANDN U519 ( .A(n3), .B(N1880), .Z(n348) );
  NAND U520 ( .A(n350), .B(n351), .Z(z3[847]) );
  NANDN U521 ( .A(N1030), .B(z2[847]), .Z(n351) );
  NANDN U522 ( .A(n3), .B(N1879), .Z(n350) );
  NAND U523 ( .A(n352), .B(n353), .Z(z3[846]) );
  NANDN U524 ( .A(N1030), .B(z2[846]), .Z(n353) );
  NANDN U525 ( .A(n3), .B(N1878), .Z(n352) );
  NAND U526 ( .A(n354), .B(n355), .Z(z3[845]) );
  NANDN U527 ( .A(N1030), .B(z2[845]), .Z(n355) );
  NANDN U528 ( .A(n3), .B(N1877), .Z(n354) );
  NAND U529 ( .A(n356), .B(n357), .Z(z3[844]) );
  NANDN U530 ( .A(N1030), .B(z2[844]), .Z(n357) );
  NANDN U531 ( .A(n3), .B(N1876), .Z(n356) );
  NAND U532 ( .A(n358), .B(n359), .Z(z3[843]) );
  NANDN U533 ( .A(N1030), .B(z2[843]), .Z(n359) );
  NANDN U534 ( .A(n3), .B(N1875), .Z(n358) );
  NAND U535 ( .A(n360), .B(n361), .Z(z3[842]) );
  NANDN U536 ( .A(N1030), .B(z2[842]), .Z(n361) );
  NANDN U537 ( .A(n3), .B(N1874), .Z(n360) );
  NAND U538 ( .A(n362), .B(n363), .Z(z3[841]) );
  NANDN U539 ( .A(N1030), .B(z2[841]), .Z(n363) );
  NANDN U540 ( .A(n3), .B(N1873), .Z(n362) );
  NAND U541 ( .A(n364), .B(n365), .Z(z3[840]) );
  NANDN U542 ( .A(N1030), .B(z2[840]), .Z(n365) );
  NANDN U543 ( .A(n3), .B(N1872), .Z(n364) );
  NAND U544 ( .A(n366), .B(n367), .Z(z3[83]) );
  NANDN U545 ( .A(N1030), .B(z2[83]), .Z(n367) );
  NANDN U546 ( .A(n3), .B(N1115), .Z(n366) );
  NAND U547 ( .A(n368), .B(n369), .Z(z3[839]) );
  NANDN U548 ( .A(N1030), .B(z2[839]), .Z(n369) );
  NANDN U549 ( .A(n3), .B(N1871), .Z(n368) );
  NAND U550 ( .A(n370), .B(n371), .Z(z3[838]) );
  NANDN U551 ( .A(N1030), .B(z2[838]), .Z(n371) );
  NANDN U552 ( .A(n3), .B(N1870), .Z(n370) );
  NAND U553 ( .A(n372), .B(n373), .Z(z3[837]) );
  NANDN U554 ( .A(N1030), .B(z2[837]), .Z(n373) );
  NANDN U555 ( .A(n3), .B(N1869), .Z(n372) );
  NAND U556 ( .A(n374), .B(n375), .Z(z3[836]) );
  NANDN U557 ( .A(N1030), .B(z2[836]), .Z(n375) );
  NANDN U558 ( .A(n3), .B(N1868), .Z(n374) );
  NAND U559 ( .A(n376), .B(n377), .Z(z3[835]) );
  NANDN U560 ( .A(N1030), .B(z2[835]), .Z(n377) );
  NANDN U561 ( .A(n3), .B(N1867), .Z(n376) );
  NAND U562 ( .A(n378), .B(n379), .Z(z3[834]) );
  NANDN U563 ( .A(N1030), .B(z2[834]), .Z(n379) );
  NANDN U564 ( .A(n3), .B(N1866), .Z(n378) );
  NAND U565 ( .A(n380), .B(n381), .Z(z3[833]) );
  NANDN U566 ( .A(N1030), .B(z2[833]), .Z(n381) );
  NANDN U567 ( .A(n3), .B(N1865), .Z(n380) );
  NAND U568 ( .A(n382), .B(n383), .Z(z3[832]) );
  NANDN U569 ( .A(N1030), .B(z2[832]), .Z(n383) );
  NANDN U570 ( .A(n3), .B(N1864), .Z(n382) );
  NAND U571 ( .A(n384), .B(n385), .Z(z3[831]) );
  NANDN U572 ( .A(N1030), .B(z2[831]), .Z(n385) );
  NANDN U573 ( .A(n3), .B(N1863), .Z(n384) );
  NAND U574 ( .A(n386), .B(n387), .Z(z3[830]) );
  NANDN U575 ( .A(N1030), .B(z2[830]), .Z(n387) );
  NANDN U576 ( .A(n3), .B(N1862), .Z(n386) );
  NAND U577 ( .A(n388), .B(n389), .Z(z3[82]) );
  NANDN U578 ( .A(N1030), .B(z2[82]), .Z(n389) );
  NANDN U579 ( .A(n3), .B(N1114), .Z(n388) );
  NAND U580 ( .A(n390), .B(n391), .Z(z3[829]) );
  NANDN U581 ( .A(N1030), .B(z2[829]), .Z(n391) );
  NANDN U582 ( .A(n3), .B(N1861), .Z(n390) );
  NAND U583 ( .A(n392), .B(n393), .Z(z3[828]) );
  NANDN U584 ( .A(N1030), .B(z2[828]), .Z(n393) );
  NANDN U585 ( .A(n3), .B(N1860), .Z(n392) );
  NAND U586 ( .A(n394), .B(n395), .Z(z3[827]) );
  NANDN U587 ( .A(N1030), .B(z2[827]), .Z(n395) );
  NANDN U588 ( .A(n3), .B(N1859), .Z(n394) );
  NAND U589 ( .A(n396), .B(n397), .Z(z3[826]) );
  NANDN U590 ( .A(N1030), .B(z2[826]), .Z(n397) );
  NANDN U591 ( .A(n3), .B(N1858), .Z(n396) );
  NAND U592 ( .A(n398), .B(n399), .Z(z3[825]) );
  NANDN U593 ( .A(N1030), .B(z2[825]), .Z(n399) );
  NANDN U594 ( .A(n3), .B(N1857), .Z(n398) );
  NAND U595 ( .A(n400), .B(n401), .Z(z3[824]) );
  NANDN U596 ( .A(N1030), .B(z2[824]), .Z(n401) );
  NANDN U597 ( .A(n3), .B(N1856), .Z(n400) );
  NAND U598 ( .A(n402), .B(n403), .Z(z3[823]) );
  NANDN U599 ( .A(N1030), .B(z2[823]), .Z(n403) );
  NANDN U600 ( .A(n3), .B(N1855), .Z(n402) );
  NAND U601 ( .A(n404), .B(n405), .Z(z3[822]) );
  NANDN U602 ( .A(N1030), .B(z2[822]), .Z(n405) );
  NANDN U603 ( .A(n3), .B(N1854), .Z(n404) );
  NAND U604 ( .A(n406), .B(n407), .Z(z3[821]) );
  NANDN U605 ( .A(N1030), .B(z2[821]), .Z(n407) );
  NANDN U606 ( .A(n3), .B(N1853), .Z(n406) );
  NAND U607 ( .A(n408), .B(n409), .Z(z3[820]) );
  NANDN U608 ( .A(N1030), .B(z2[820]), .Z(n409) );
  NANDN U609 ( .A(n3), .B(N1852), .Z(n408) );
  NAND U610 ( .A(n410), .B(n411), .Z(z3[81]) );
  NANDN U611 ( .A(N1030), .B(z2[81]), .Z(n411) );
  NANDN U612 ( .A(n3), .B(N1113), .Z(n410) );
  NAND U613 ( .A(n412), .B(n413), .Z(z3[819]) );
  NANDN U614 ( .A(N1030), .B(z2[819]), .Z(n413) );
  NANDN U615 ( .A(n3), .B(N1851), .Z(n412) );
  NAND U616 ( .A(n414), .B(n415), .Z(z3[818]) );
  NANDN U617 ( .A(N1030), .B(z2[818]), .Z(n415) );
  NANDN U618 ( .A(n3), .B(N1850), .Z(n414) );
  NAND U619 ( .A(n416), .B(n417), .Z(z3[817]) );
  NANDN U620 ( .A(N1030), .B(z2[817]), .Z(n417) );
  NANDN U621 ( .A(n3), .B(N1849), .Z(n416) );
  NAND U622 ( .A(n418), .B(n419), .Z(z3[816]) );
  NANDN U623 ( .A(N1030), .B(z2[816]), .Z(n419) );
  NANDN U624 ( .A(n3), .B(N1848), .Z(n418) );
  NAND U625 ( .A(n420), .B(n421), .Z(z3[815]) );
  NANDN U626 ( .A(N1030), .B(z2[815]), .Z(n421) );
  NANDN U627 ( .A(n3), .B(N1847), .Z(n420) );
  NAND U628 ( .A(n422), .B(n423), .Z(z3[814]) );
  NANDN U629 ( .A(N1030), .B(z2[814]), .Z(n423) );
  NANDN U630 ( .A(n3), .B(N1846), .Z(n422) );
  NAND U631 ( .A(n424), .B(n425), .Z(z3[813]) );
  NANDN U632 ( .A(N1030), .B(z2[813]), .Z(n425) );
  NANDN U633 ( .A(n3), .B(N1845), .Z(n424) );
  NAND U634 ( .A(n426), .B(n427), .Z(z3[812]) );
  NANDN U635 ( .A(N1030), .B(z2[812]), .Z(n427) );
  NANDN U636 ( .A(n3), .B(N1844), .Z(n426) );
  NAND U637 ( .A(n428), .B(n429), .Z(z3[811]) );
  NANDN U638 ( .A(N1030), .B(z2[811]), .Z(n429) );
  NANDN U639 ( .A(n3), .B(N1843), .Z(n428) );
  NAND U640 ( .A(n430), .B(n431), .Z(z3[810]) );
  NANDN U641 ( .A(N1030), .B(z2[810]), .Z(n431) );
  NANDN U642 ( .A(n3), .B(N1842), .Z(n430) );
  NAND U643 ( .A(n432), .B(n433), .Z(z3[80]) );
  NANDN U644 ( .A(N1030), .B(z2[80]), .Z(n433) );
  NANDN U645 ( .A(n3), .B(N1112), .Z(n432) );
  NAND U646 ( .A(n434), .B(n435), .Z(z3[809]) );
  NANDN U647 ( .A(N1030), .B(z2[809]), .Z(n435) );
  NANDN U648 ( .A(n3), .B(N1841), .Z(n434) );
  NAND U649 ( .A(n436), .B(n437), .Z(z3[808]) );
  NANDN U650 ( .A(N1030), .B(z2[808]), .Z(n437) );
  NANDN U651 ( .A(n3), .B(N1840), .Z(n436) );
  NAND U652 ( .A(n438), .B(n439), .Z(z3[807]) );
  NANDN U653 ( .A(N1030), .B(z2[807]), .Z(n439) );
  NANDN U654 ( .A(n3), .B(N1839), .Z(n438) );
  NAND U655 ( .A(n440), .B(n441), .Z(z3[806]) );
  NANDN U656 ( .A(N1030), .B(z2[806]), .Z(n441) );
  NANDN U657 ( .A(n3), .B(N1838), .Z(n440) );
  NAND U658 ( .A(n442), .B(n443), .Z(z3[805]) );
  NANDN U659 ( .A(N1030), .B(z2[805]), .Z(n443) );
  NANDN U660 ( .A(n3), .B(N1837), .Z(n442) );
  NAND U661 ( .A(n444), .B(n445), .Z(z3[804]) );
  NANDN U662 ( .A(N1030), .B(z2[804]), .Z(n445) );
  NANDN U663 ( .A(n3), .B(N1836), .Z(n444) );
  NAND U664 ( .A(n446), .B(n447), .Z(z3[803]) );
  NANDN U665 ( .A(N1030), .B(z2[803]), .Z(n447) );
  NANDN U666 ( .A(n3), .B(N1835), .Z(n446) );
  NAND U667 ( .A(n448), .B(n449), .Z(z3[802]) );
  NANDN U668 ( .A(N1030), .B(z2[802]), .Z(n449) );
  NANDN U669 ( .A(n3), .B(N1834), .Z(n448) );
  NAND U670 ( .A(n450), .B(n451), .Z(z3[801]) );
  NANDN U671 ( .A(N1030), .B(z2[801]), .Z(n451) );
  NANDN U672 ( .A(n3), .B(N1833), .Z(n450) );
  NAND U673 ( .A(n452), .B(n453), .Z(z3[800]) );
  NANDN U674 ( .A(N1030), .B(z2[800]), .Z(n453) );
  NANDN U675 ( .A(n3), .B(N1832), .Z(n452) );
  NAND U676 ( .A(n454), .B(n455), .Z(z3[7]) );
  NANDN U677 ( .A(N1030), .B(z2[7]), .Z(n455) );
  NANDN U678 ( .A(n3), .B(N1039), .Z(n454) );
  NAND U679 ( .A(n456), .B(n457), .Z(z3[79]) );
  NANDN U680 ( .A(N1030), .B(z2[79]), .Z(n457) );
  NANDN U681 ( .A(n3), .B(N1111), .Z(n456) );
  NAND U682 ( .A(n458), .B(n459), .Z(z3[799]) );
  NANDN U683 ( .A(N1030), .B(z2[799]), .Z(n459) );
  NANDN U684 ( .A(n3), .B(N1831), .Z(n458) );
  NAND U685 ( .A(n460), .B(n461), .Z(z3[798]) );
  NANDN U686 ( .A(N1030), .B(z2[798]), .Z(n461) );
  NANDN U687 ( .A(n3), .B(N1830), .Z(n460) );
  NAND U688 ( .A(n462), .B(n463), .Z(z3[797]) );
  NANDN U689 ( .A(N1030), .B(z2[797]), .Z(n463) );
  NANDN U690 ( .A(n3), .B(N1829), .Z(n462) );
  NAND U691 ( .A(n464), .B(n465), .Z(z3[796]) );
  NANDN U692 ( .A(N1030), .B(z2[796]), .Z(n465) );
  NANDN U693 ( .A(n3), .B(N1828), .Z(n464) );
  NAND U694 ( .A(n466), .B(n467), .Z(z3[795]) );
  NANDN U695 ( .A(N1030), .B(z2[795]), .Z(n467) );
  NANDN U696 ( .A(n3), .B(N1827), .Z(n466) );
  NAND U697 ( .A(n468), .B(n469), .Z(z3[794]) );
  NANDN U698 ( .A(N1030), .B(z2[794]), .Z(n469) );
  NANDN U699 ( .A(n3), .B(N1826), .Z(n468) );
  NAND U700 ( .A(n470), .B(n471), .Z(z3[793]) );
  NANDN U701 ( .A(N1030), .B(z2[793]), .Z(n471) );
  NANDN U702 ( .A(n3), .B(N1825), .Z(n470) );
  NAND U703 ( .A(n472), .B(n473), .Z(z3[792]) );
  NANDN U704 ( .A(N1030), .B(z2[792]), .Z(n473) );
  NANDN U705 ( .A(n3), .B(N1824), .Z(n472) );
  NAND U706 ( .A(n474), .B(n475), .Z(z3[791]) );
  NANDN U707 ( .A(N1030), .B(z2[791]), .Z(n475) );
  NANDN U708 ( .A(n3), .B(N1823), .Z(n474) );
  NAND U709 ( .A(n476), .B(n477), .Z(z3[790]) );
  NANDN U710 ( .A(N1030), .B(z2[790]), .Z(n477) );
  NANDN U711 ( .A(n3), .B(N1822), .Z(n476) );
  NAND U712 ( .A(n478), .B(n479), .Z(z3[78]) );
  NANDN U713 ( .A(N1030), .B(z2[78]), .Z(n479) );
  NANDN U714 ( .A(n3), .B(N1110), .Z(n478) );
  NAND U715 ( .A(n480), .B(n481), .Z(z3[789]) );
  NANDN U716 ( .A(N1030), .B(z2[789]), .Z(n481) );
  NANDN U717 ( .A(n3), .B(N1821), .Z(n480) );
  NAND U718 ( .A(n482), .B(n483), .Z(z3[788]) );
  NANDN U719 ( .A(N1030), .B(z2[788]), .Z(n483) );
  NANDN U720 ( .A(n3), .B(N1820), .Z(n482) );
  NAND U721 ( .A(n484), .B(n485), .Z(z3[787]) );
  NANDN U722 ( .A(N1030), .B(z2[787]), .Z(n485) );
  NANDN U723 ( .A(n3), .B(N1819), .Z(n484) );
  NAND U724 ( .A(n486), .B(n487), .Z(z3[786]) );
  NANDN U725 ( .A(N1030), .B(z2[786]), .Z(n487) );
  NANDN U726 ( .A(n3), .B(N1818), .Z(n486) );
  NAND U727 ( .A(n488), .B(n489), .Z(z3[785]) );
  NANDN U728 ( .A(N1030), .B(z2[785]), .Z(n489) );
  NANDN U729 ( .A(n3), .B(N1817), .Z(n488) );
  NAND U730 ( .A(n490), .B(n491), .Z(z3[784]) );
  NANDN U731 ( .A(N1030), .B(z2[784]), .Z(n491) );
  NANDN U732 ( .A(n3), .B(N1816), .Z(n490) );
  NAND U733 ( .A(n492), .B(n493), .Z(z3[783]) );
  NANDN U734 ( .A(N1030), .B(z2[783]), .Z(n493) );
  NANDN U735 ( .A(n3), .B(N1815), .Z(n492) );
  NAND U736 ( .A(n494), .B(n495), .Z(z3[782]) );
  NANDN U737 ( .A(N1030), .B(z2[782]), .Z(n495) );
  NANDN U738 ( .A(n3), .B(N1814), .Z(n494) );
  NAND U739 ( .A(n496), .B(n497), .Z(z3[781]) );
  NANDN U740 ( .A(N1030), .B(z2[781]), .Z(n497) );
  NANDN U741 ( .A(n3), .B(N1813), .Z(n496) );
  NAND U742 ( .A(n498), .B(n499), .Z(z3[780]) );
  NANDN U743 ( .A(N1030), .B(z2[780]), .Z(n499) );
  NANDN U744 ( .A(n3), .B(N1812), .Z(n498) );
  NAND U745 ( .A(n500), .B(n501), .Z(z3[77]) );
  NANDN U746 ( .A(N1030), .B(z2[77]), .Z(n501) );
  NANDN U747 ( .A(n3), .B(N1109), .Z(n500) );
  NAND U748 ( .A(n502), .B(n503), .Z(z3[779]) );
  NANDN U749 ( .A(N1030), .B(z2[779]), .Z(n503) );
  NANDN U750 ( .A(n3), .B(N1811), .Z(n502) );
  NAND U751 ( .A(n504), .B(n505), .Z(z3[778]) );
  NANDN U752 ( .A(N1030), .B(z2[778]), .Z(n505) );
  NANDN U753 ( .A(n3), .B(N1810), .Z(n504) );
  NAND U754 ( .A(n506), .B(n507), .Z(z3[777]) );
  NANDN U755 ( .A(N1030), .B(z2[777]), .Z(n507) );
  NANDN U756 ( .A(n3), .B(N1809), .Z(n506) );
  NAND U757 ( .A(n508), .B(n509), .Z(z3[776]) );
  NANDN U758 ( .A(N1030), .B(z2[776]), .Z(n509) );
  NANDN U759 ( .A(n3), .B(N1808), .Z(n508) );
  NAND U760 ( .A(n510), .B(n511), .Z(z3[775]) );
  NANDN U761 ( .A(N1030), .B(z2[775]), .Z(n511) );
  NANDN U762 ( .A(n3), .B(N1807), .Z(n510) );
  NAND U763 ( .A(n512), .B(n513), .Z(z3[774]) );
  NANDN U764 ( .A(N1030), .B(z2[774]), .Z(n513) );
  NANDN U765 ( .A(n3), .B(N1806), .Z(n512) );
  NAND U766 ( .A(n514), .B(n515), .Z(z3[773]) );
  NANDN U767 ( .A(N1030), .B(z2[773]), .Z(n515) );
  NANDN U768 ( .A(n3), .B(N1805), .Z(n514) );
  NAND U769 ( .A(n516), .B(n517), .Z(z3[772]) );
  NANDN U770 ( .A(N1030), .B(z2[772]), .Z(n517) );
  NANDN U771 ( .A(n3), .B(N1804), .Z(n516) );
  NAND U772 ( .A(n518), .B(n519), .Z(z3[771]) );
  NANDN U773 ( .A(N1030), .B(z2[771]), .Z(n519) );
  NANDN U774 ( .A(n3), .B(N1803), .Z(n518) );
  NAND U775 ( .A(n520), .B(n521), .Z(z3[770]) );
  NANDN U776 ( .A(N1030), .B(z2[770]), .Z(n521) );
  NANDN U777 ( .A(n3), .B(N1802), .Z(n520) );
  NAND U778 ( .A(n522), .B(n523), .Z(z3[76]) );
  NANDN U779 ( .A(N1030), .B(z2[76]), .Z(n523) );
  NANDN U780 ( .A(n3), .B(N1108), .Z(n522) );
  NAND U781 ( .A(n524), .B(n525), .Z(z3[769]) );
  NANDN U782 ( .A(N1030), .B(z2[769]), .Z(n525) );
  NANDN U783 ( .A(n3), .B(N1801), .Z(n524) );
  NAND U784 ( .A(n526), .B(n527), .Z(z3[768]) );
  NANDN U785 ( .A(N1030), .B(z2[768]), .Z(n527) );
  NANDN U786 ( .A(n3), .B(N1800), .Z(n526) );
  NAND U787 ( .A(n528), .B(n529), .Z(z3[767]) );
  NANDN U788 ( .A(N1030), .B(z2[767]), .Z(n529) );
  NANDN U789 ( .A(n3), .B(N1799), .Z(n528) );
  NAND U790 ( .A(n530), .B(n531), .Z(z3[766]) );
  NANDN U791 ( .A(N1030), .B(z2[766]), .Z(n531) );
  NANDN U792 ( .A(n3), .B(N1798), .Z(n530) );
  NAND U793 ( .A(n532), .B(n533), .Z(z3[765]) );
  NANDN U794 ( .A(N1030), .B(z2[765]), .Z(n533) );
  NANDN U795 ( .A(n3), .B(N1797), .Z(n532) );
  NAND U796 ( .A(n534), .B(n535), .Z(z3[764]) );
  NANDN U797 ( .A(N1030), .B(z2[764]), .Z(n535) );
  NANDN U798 ( .A(n3), .B(N1796), .Z(n534) );
  NAND U799 ( .A(n536), .B(n537), .Z(z3[763]) );
  NANDN U800 ( .A(N1030), .B(z2[763]), .Z(n537) );
  NANDN U801 ( .A(n3), .B(N1795), .Z(n536) );
  NAND U802 ( .A(n538), .B(n539), .Z(z3[762]) );
  NANDN U803 ( .A(N1030), .B(z2[762]), .Z(n539) );
  NANDN U804 ( .A(n3), .B(N1794), .Z(n538) );
  NAND U805 ( .A(n540), .B(n541), .Z(z3[761]) );
  NANDN U806 ( .A(N1030), .B(z2[761]), .Z(n541) );
  NANDN U807 ( .A(n3), .B(N1793), .Z(n540) );
  NAND U808 ( .A(n542), .B(n543), .Z(z3[760]) );
  NANDN U809 ( .A(N1030), .B(z2[760]), .Z(n543) );
  NANDN U810 ( .A(n3), .B(N1792), .Z(n542) );
  NAND U811 ( .A(n544), .B(n545), .Z(z3[75]) );
  NANDN U812 ( .A(N1030), .B(z2[75]), .Z(n545) );
  NANDN U813 ( .A(n3), .B(N1107), .Z(n544) );
  NAND U814 ( .A(n546), .B(n547), .Z(z3[759]) );
  NANDN U815 ( .A(N1030), .B(z2[759]), .Z(n547) );
  NANDN U816 ( .A(n3), .B(N1791), .Z(n546) );
  NAND U817 ( .A(n548), .B(n549), .Z(z3[758]) );
  NANDN U818 ( .A(N1030), .B(z2[758]), .Z(n549) );
  NANDN U819 ( .A(n3), .B(N1790), .Z(n548) );
  NAND U820 ( .A(n550), .B(n551), .Z(z3[757]) );
  NANDN U821 ( .A(N1030), .B(z2[757]), .Z(n551) );
  NANDN U822 ( .A(n3), .B(N1789), .Z(n550) );
  NAND U823 ( .A(n552), .B(n553), .Z(z3[756]) );
  NANDN U824 ( .A(N1030), .B(z2[756]), .Z(n553) );
  NANDN U825 ( .A(n3), .B(N1788), .Z(n552) );
  NAND U826 ( .A(n554), .B(n555), .Z(z3[755]) );
  NANDN U827 ( .A(N1030), .B(z2[755]), .Z(n555) );
  NANDN U828 ( .A(n3), .B(N1787), .Z(n554) );
  NAND U829 ( .A(n556), .B(n557), .Z(z3[754]) );
  NANDN U830 ( .A(N1030), .B(z2[754]), .Z(n557) );
  NANDN U831 ( .A(n3), .B(N1786), .Z(n556) );
  NAND U832 ( .A(n558), .B(n559), .Z(z3[753]) );
  NANDN U833 ( .A(N1030), .B(z2[753]), .Z(n559) );
  NANDN U834 ( .A(n3), .B(N1785), .Z(n558) );
  NAND U835 ( .A(n560), .B(n561), .Z(z3[752]) );
  NANDN U836 ( .A(N1030), .B(z2[752]), .Z(n561) );
  NANDN U837 ( .A(n3), .B(N1784), .Z(n560) );
  NAND U838 ( .A(n562), .B(n563), .Z(z3[751]) );
  NANDN U839 ( .A(N1030), .B(z2[751]), .Z(n563) );
  NANDN U840 ( .A(n3), .B(N1783), .Z(n562) );
  NAND U841 ( .A(n564), .B(n565), .Z(z3[750]) );
  NANDN U842 ( .A(N1030), .B(z2[750]), .Z(n565) );
  NANDN U843 ( .A(n3), .B(N1782), .Z(n564) );
  NAND U844 ( .A(n566), .B(n567), .Z(z3[74]) );
  NANDN U845 ( .A(N1030), .B(z2[74]), .Z(n567) );
  NANDN U846 ( .A(n3), .B(N1106), .Z(n566) );
  NAND U847 ( .A(n568), .B(n569), .Z(z3[749]) );
  NANDN U848 ( .A(N1030), .B(z2[749]), .Z(n569) );
  NANDN U849 ( .A(n3), .B(N1781), .Z(n568) );
  NAND U850 ( .A(n570), .B(n571), .Z(z3[748]) );
  NANDN U851 ( .A(N1030), .B(z2[748]), .Z(n571) );
  NANDN U852 ( .A(n3), .B(N1780), .Z(n570) );
  NAND U853 ( .A(n572), .B(n573), .Z(z3[747]) );
  NANDN U854 ( .A(N1030), .B(z2[747]), .Z(n573) );
  NANDN U855 ( .A(n3), .B(N1779), .Z(n572) );
  NAND U856 ( .A(n574), .B(n575), .Z(z3[746]) );
  NANDN U857 ( .A(N1030), .B(z2[746]), .Z(n575) );
  NANDN U858 ( .A(n3), .B(N1778), .Z(n574) );
  NAND U859 ( .A(n576), .B(n577), .Z(z3[745]) );
  NANDN U860 ( .A(N1030), .B(z2[745]), .Z(n577) );
  NANDN U861 ( .A(n3), .B(N1777), .Z(n576) );
  NAND U862 ( .A(n578), .B(n579), .Z(z3[744]) );
  NANDN U863 ( .A(N1030), .B(z2[744]), .Z(n579) );
  NANDN U864 ( .A(n3), .B(N1776), .Z(n578) );
  NAND U865 ( .A(n580), .B(n581), .Z(z3[743]) );
  NANDN U866 ( .A(N1030), .B(z2[743]), .Z(n581) );
  NANDN U867 ( .A(n3), .B(N1775), .Z(n580) );
  NAND U868 ( .A(n582), .B(n583), .Z(z3[742]) );
  NANDN U869 ( .A(N1030), .B(z2[742]), .Z(n583) );
  NANDN U870 ( .A(n3), .B(N1774), .Z(n582) );
  NAND U871 ( .A(n584), .B(n585), .Z(z3[741]) );
  NANDN U872 ( .A(N1030), .B(z2[741]), .Z(n585) );
  NANDN U873 ( .A(n3), .B(N1773), .Z(n584) );
  NAND U874 ( .A(n586), .B(n587), .Z(z3[740]) );
  NANDN U875 ( .A(N1030), .B(z2[740]), .Z(n587) );
  NANDN U876 ( .A(n3), .B(N1772), .Z(n586) );
  NAND U877 ( .A(n588), .B(n589), .Z(z3[73]) );
  NANDN U878 ( .A(N1030), .B(z2[73]), .Z(n589) );
  NANDN U879 ( .A(n3), .B(N1105), .Z(n588) );
  NAND U880 ( .A(n590), .B(n591), .Z(z3[739]) );
  NANDN U881 ( .A(N1030), .B(z2[739]), .Z(n591) );
  NANDN U882 ( .A(n3), .B(N1771), .Z(n590) );
  NAND U883 ( .A(n592), .B(n593), .Z(z3[738]) );
  NANDN U884 ( .A(N1030), .B(z2[738]), .Z(n593) );
  NANDN U885 ( .A(n3), .B(N1770), .Z(n592) );
  NAND U886 ( .A(n594), .B(n595), .Z(z3[737]) );
  NANDN U887 ( .A(N1030), .B(z2[737]), .Z(n595) );
  NANDN U888 ( .A(n3), .B(N1769), .Z(n594) );
  NAND U889 ( .A(n596), .B(n597), .Z(z3[736]) );
  NANDN U890 ( .A(N1030), .B(z2[736]), .Z(n597) );
  NANDN U891 ( .A(n3), .B(N1768), .Z(n596) );
  NAND U892 ( .A(n598), .B(n599), .Z(z3[735]) );
  NANDN U893 ( .A(N1030), .B(z2[735]), .Z(n599) );
  NANDN U894 ( .A(n3), .B(N1767), .Z(n598) );
  NAND U895 ( .A(n600), .B(n601), .Z(z3[734]) );
  NANDN U896 ( .A(N1030), .B(z2[734]), .Z(n601) );
  NANDN U897 ( .A(n3), .B(N1766), .Z(n600) );
  NAND U898 ( .A(n602), .B(n603), .Z(z3[733]) );
  NANDN U899 ( .A(N1030), .B(z2[733]), .Z(n603) );
  NANDN U900 ( .A(n3), .B(N1765), .Z(n602) );
  NAND U901 ( .A(n604), .B(n605), .Z(z3[732]) );
  NANDN U902 ( .A(N1030), .B(z2[732]), .Z(n605) );
  NANDN U903 ( .A(n3), .B(N1764), .Z(n604) );
  NAND U904 ( .A(n606), .B(n607), .Z(z3[731]) );
  NANDN U905 ( .A(N1030), .B(z2[731]), .Z(n607) );
  NANDN U906 ( .A(n3), .B(N1763), .Z(n606) );
  NAND U907 ( .A(n608), .B(n609), .Z(z3[730]) );
  NANDN U908 ( .A(N1030), .B(z2[730]), .Z(n609) );
  NANDN U909 ( .A(n3), .B(N1762), .Z(n608) );
  NAND U910 ( .A(n610), .B(n611), .Z(z3[72]) );
  NANDN U911 ( .A(N1030), .B(z2[72]), .Z(n611) );
  NANDN U912 ( .A(n3), .B(N1104), .Z(n610) );
  NAND U913 ( .A(n612), .B(n613), .Z(z3[729]) );
  NANDN U914 ( .A(N1030), .B(z2[729]), .Z(n613) );
  NANDN U915 ( .A(n3), .B(N1761), .Z(n612) );
  NAND U916 ( .A(n614), .B(n615), .Z(z3[728]) );
  NANDN U917 ( .A(N1030), .B(z2[728]), .Z(n615) );
  NANDN U918 ( .A(n3), .B(N1760), .Z(n614) );
  NAND U919 ( .A(n616), .B(n617), .Z(z3[727]) );
  NANDN U920 ( .A(N1030), .B(z2[727]), .Z(n617) );
  NANDN U921 ( .A(n3), .B(N1759), .Z(n616) );
  NAND U922 ( .A(n618), .B(n619), .Z(z3[726]) );
  NANDN U923 ( .A(N1030), .B(z2[726]), .Z(n619) );
  NANDN U924 ( .A(n3), .B(N1758), .Z(n618) );
  NAND U925 ( .A(n620), .B(n621), .Z(z3[725]) );
  NANDN U926 ( .A(N1030), .B(z2[725]), .Z(n621) );
  NANDN U927 ( .A(n3), .B(N1757), .Z(n620) );
  NAND U928 ( .A(n622), .B(n623), .Z(z3[724]) );
  NANDN U929 ( .A(N1030), .B(z2[724]), .Z(n623) );
  NANDN U930 ( .A(n3), .B(N1756), .Z(n622) );
  NAND U931 ( .A(n624), .B(n625), .Z(z3[723]) );
  NANDN U932 ( .A(N1030), .B(z2[723]), .Z(n625) );
  NANDN U933 ( .A(n3), .B(N1755), .Z(n624) );
  NAND U934 ( .A(n626), .B(n627), .Z(z3[722]) );
  NANDN U935 ( .A(N1030), .B(z2[722]), .Z(n627) );
  NANDN U936 ( .A(n3), .B(N1754), .Z(n626) );
  NAND U937 ( .A(n628), .B(n629), .Z(z3[721]) );
  NANDN U938 ( .A(N1030), .B(z2[721]), .Z(n629) );
  NANDN U939 ( .A(n3), .B(N1753), .Z(n628) );
  NAND U940 ( .A(n630), .B(n631), .Z(z3[720]) );
  NANDN U941 ( .A(N1030), .B(z2[720]), .Z(n631) );
  NANDN U942 ( .A(n3), .B(N1752), .Z(n630) );
  NAND U943 ( .A(n632), .B(n633), .Z(z3[71]) );
  NANDN U944 ( .A(N1030), .B(z2[71]), .Z(n633) );
  NANDN U945 ( .A(n3), .B(N1103), .Z(n632) );
  NAND U946 ( .A(n634), .B(n635), .Z(z3[719]) );
  NANDN U947 ( .A(N1030), .B(z2[719]), .Z(n635) );
  NANDN U948 ( .A(n3), .B(N1751), .Z(n634) );
  NAND U949 ( .A(n636), .B(n637), .Z(z3[718]) );
  NANDN U950 ( .A(N1030), .B(z2[718]), .Z(n637) );
  NANDN U951 ( .A(n3), .B(N1750), .Z(n636) );
  NAND U952 ( .A(n638), .B(n639), .Z(z3[717]) );
  NANDN U953 ( .A(N1030), .B(z2[717]), .Z(n639) );
  NANDN U954 ( .A(n3), .B(N1749), .Z(n638) );
  NAND U955 ( .A(n640), .B(n641), .Z(z3[716]) );
  NANDN U956 ( .A(N1030), .B(z2[716]), .Z(n641) );
  NANDN U957 ( .A(n3), .B(N1748), .Z(n640) );
  NAND U958 ( .A(n642), .B(n643), .Z(z3[715]) );
  NANDN U959 ( .A(N1030), .B(z2[715]), .Z(n643) );
  NANDN U960 ( .A(n3), .B(N1747), .Z(n642) );
  NAND U961 ( .A(n644), .B(n645), .Z(z3[714]) );
  NANDN U962 ( .A(N1030), .B(z2[714]), .Z(n645) );
  NANDN U963 ( .A(n3), .B(N1746), .Z(n644) );
  NAND U964 ( .A(n646), .B(n647), .Z(z3[713]) );
  NANDN U965 ( .A(N1030), .B(z2[713]), .Z(n647) );
  NANDN U966 ( .A(n3), .B(N1745), .Z(n646) );
  NAND U967 ( .A(n648), .B(n649), .Z(z3[712]) );
  NANDN U968 ( .A(N1030), .B(z2[712]), .Z(n649) );
  NANDN U969 ( .A(n3), .B(N1744), .Z(n648) );
  NAND U970 ( .A(n650), .B(n651), .Z(z3[711]) );
  NANDN U971 ( .A(N1030), .B(z2[711]), .Z(n651) );
  NANDN U972 ( .A(n3), .B(N1743), .Z(n650) );
  NAND U973 ( .A(n652), .B(n653), .Z(z3[710]) );
  NANDN U974 ( .A(N1030), .B(z2[710]), .Z(n653) );
  NANDN U975 ( .A(n3), .B(N1742), .Z(n652) );
  NAND U976 ( .A(n654), .B(n655), .Z(z3[70]) );
  NANDN U977 ( .A(N1030), .B(z2[70]), .Z(n655) );
  NANDN U978 ( .A(n3), .B(N1102), .Z(n654) );
  NAND U979 ( .A(n656), .B(n657), .Z(z3[709]) );
  NANDN U980 ( .A(N1030), .B(z2[709]), .Z(n657) );
  NANDN U981 ( .A(n3), .B(N1741), .Z(n656) );
  NAND U982 ( .A(n658), .B(n659), .Z(z3[708]) );
  NANDN U983 ( .A(N1030), .B(z2[708]), .Z(n659) );
  NANDN U984 ( .A(n3), .B(N1740), .Z(n658) );
  NAND U985 ( .A(n660), .B(n661), .Z(z3[707]) );
  NANDN U986 ( .A(N1030), .B(z2[707]), .Z(n661) );
  NANDN U987 ( .A(n3), .B(N1739), .Z(n660) );
  NAND U988 ( .A(n662), .B(n663), .Z(z3[706]) );
  NANDN U989 ( .A(N1030), .B(z2[706]), .Z(n663) );
  NANDN U990 ( .A(n3), .B(N1738), .Z(n662) );
  NAND U991 ( .A(n664), .B(n665), .Z(z3[705]) );
  NANDN U992 ( .A(N1030), .B(z2[705]), .Z(n665) );
  NANDN U993 ( .A(n3), .B(N1737), .Z(n664) );
  NAND U994 ( .A(n666), .B(n667), .Z(z3[704]) );
  NANDN U995 ( .A(N1030), .B(z2[704]), .Z(n667) );
  NANDN U996 ( .A(n3), .B(N1736), .Z(n666) );
  NAND U997 ( .A(n668), .B(n669), .Z(z3[703]) );
  NANDN U998 ( .A(N1030), .B(z2[703]), .Z(n669) );
  NANDN U999 ( .A(n3), .B(N1735), .Z(n668) );
  NAND U1000 ( .A(n670), .B(n671), .Z(z3[702]) );
  NANDN U1001 ( .A(N1030), .B(z2[702]), .Z(n671) );
  NANDN U1002 ( .A(n3), .B(N1734), .Z(n670) );
  NAND U1003 ( .A(n672), .B(n673), .Z(z3[701]) );
  NANDN U1004 ( .A(N1030), .B(z2[701]), .Z(n673) );
  NANDN U1005 ( .A(n3), .B(N1733), .Z(n672) );
  NAND U1006 ( .A(n674), .B(n675), .Z(z3[700]) );
  NANDN U1007 ( .A(N1030), .B(z2[700]), .Z(n675) );
  NANDN U1008 ( .A(n3), .B(N1732), .Z(n674) );
  NAND U1009 ( .A(n676), .B(n677), .Z(z3[6]) );
  NANDN U1010 ( .A(N1030), .B(z2[6]), .Z(n677) );
  NANDN U1011 ( .A(n3), .B(N1038), .Z(n676) );
  NAND U1012 ( .A(n678), .B(n679), .Z(z3[69]) );
  NANDN U1013 ( .A(N1030), .B(z2[69]), .Z(n679) );
  NANDN U1014 ( .A(n3), .B(N1101), .Z(n678) );
  NAND U1015 ( .A(n680), .B(n681), .Z(z3[699]) );
  NANDN U1016 ( .A(N1030), .B(z2[699]), .Z(n681) );
  NANDN U1017 ( .A(n3), .B(N1731), .Z(n680) );
  NAND U1018 ( .A(n682), .B(n683), .Z(z3[698]) );
  NANDN U1019 ( .A(N1030), .B(z2[698]), .Z(n683) );
  NANDN U1020 ( .A(n3), .B(N1730), .Z(n682) );
  NAND U1021 ( .A(n684), .B(n685), .Z(z3[697]) );
  NANDN U1022 ( .A(N1030), .B(z2[697]), .Z(n685) );
  NANDN U1023 ( .A(n3), .B(N1729), .Z(n684) );
  NAND U1024 ( .A(n686), .B(n687), .Z(z3[696]) );
  NANDN U1025 ( .A(N1030), .B(z2[696]), .Z(n687) );
  NANDN U1026 ( .A(n3), .B(N1728), .Z(n686) );
  NAND U1027 ( .A(n688), .B(n689), .Z(z3[695]) );
  NANDN U1028 ( .A(N1030), .B(z2[695]), .Z(n689) );
  NANDN U1029 ( .A(n3), .B(N1727), .Z(n688) );
  NAND U1030 ( .A(n690), .B(n691), .Z(z3[694]) );
  NANDN U1031 ( .A(N1030), .B(z2[694]), .Z(n691) );
  NANDN U1032 ( .A(n3), .B(N1726), .Z(n690) );
  NAND U1033 ( .A(n692), .B(n693), .Z(z3[693]) );
  NANDN U1034 ( .A(N1030), .B(z2[693]), .Z(n693) );
  NANDN U1035 ( .A(n3), .B(N1725), .Z(n692) );
  NAND U1036 ( .A(n694), .B(n695), .Z(z3[692]) );
  NANDN U1037 ( .A(N1030), .B(z2[692]), .Z(n695) );
  NANDN U1038 ( .A(n3), .B(N1724), .Z(n694) );
  NAND U1039 ( .A(n696), .B(n697), .Z(z3[691]) );
  NANDN U1040 ( .A(N1030), .B(z2[691]), .Z(n697) );
  NANDN U1041 ( .A(n3), .B(N1723), .Z(n696) );
  NAND U1042 ( .A(n698), .B(n699), .Z(z3[690]) );
  NANDN U1043 ( .A(N1030), .B(z2[690]), .Z(n699) );
  NANDN U1044 ( .A(n3), .B(N1722), .Z(n698) );
  NAND U1045 ( .A(n700), .B(n701), .Z(z3[68]) );
  NANDN U1046 ( .A(N1030), .B(z2[68]), .Z(n701) );
  NANDN U1047 ( .A(n3), .B(N1100), .Z(n700) );
  NAND U1048 ( .A(n702), .B(n703), .Z(z3[689]) );
  NANDN U1049 ( .A(N1030), .B(z2[689]), .Z(n703) );
  NANDN U1050 ( .A(n3), .B(N1721), .Z(n702) );
  NAND U1051 ( .A(n704), .B(n705), .Z(z3[688]) );
  NANDN U1052 ( .A(N1030), .B(z2[688]), .Z(n705) );
  NANDN U1053 ( .A(n3), .B(N1720), .Z(n704) );
  NAND U1054 ( .A(n706), .B(n707), .Z(z3[687]) );
  NANDN U1055 ( .A(N1030), .B(z2[687]), .Z(n707) );
  NANDN U1056 ( .A(n3), .B(N1719), .Z(n706) );
  NAND U1057 ( .A(n708), .B(n709), .Z(z3[686]) );
  NANDN U1058 ( .A(N1030), .B(z2[686]), .Z(n709) );
  NANDN U1059 ( .A(n3), .B(N1718), .Z(n708) );
  NAND U1060 ( .A(n710), .B(n711), .Z(z3[685]) );
  NANDN U1061 ( .A(N1030), .B(z2[685]), .Z(n711) );
  NANDN U1062 ( .A(n3), .B(N1717), .Z(n710) );
  NAND U1063 ( .A(n712), .B(n713), .Z(z3[684]) );
  NANDN U1064 ( .A(N1030), .B(z2[684]), .Z(n713) );
  NANDN U1065 ( .A(n3), .B(N1716), .Z(n712) );
  NAND U1066 ( .A(n714), .B(n715), .Z(z3[683]) );
  NANDN U1067 ( .A(N1030), .B(z2[683]), .Z(n715) );
  NANDN U1068 ( .A(n3), .B(N1715), .Z(n714) );
  NAND U1069 ( .A(n716), .B(n717), .Z(z3[682]) );
  NANDN U1070 ( .A(N1030), .B(z2[682]), .Z(n717) );
  NANDN U1071 ( .A(n3), .B(N1714), .Z(n716) );
  NAND U1072 ( .A(n718), .B(n719), .Z(z3[681]) );
  NANDN U1073 ( .A(N1030), .B(z2[681]), .Z(n719) );
  NANDN U1074 ( .A(n3), .B(N1713), .Z(n718) );
  NAND U1075 ( .A(n720), .B(n721), .Z(z3[680]) );
  NANDN U1076 ( .A(N1030), .B(z2[680]), .Z(n721) );
  NANDN U1077 ( .A(n3), .B(N1712), .Z(n720) );
  NAND U1078 ( .A(n722), .B(n723), .Z(z3[67]) );
  NANDN U1079 ( .A(N1030), .B(z2[67]), .Z(n723) );
  NANDN U1080 ( .A(n3), .B(N1099), .Z(n722) );
  NAND U1081 ( .A(n724), .B(n725), .Z(z3[679]) );
  NANDN U1082 ( .A(N1030), .B(z2[679]), .Z(n725) );
  NANDN U1083 ( .A(n3), .B(N1711), .Z(n724) );
  NAND U1084 ( .A(n726), .B(n727), .Z(z3[678]) );
  NANDN U1085 ( .A(N1030), .B(z2[678]), .Z(n727) );
  NANDN U1086 ( .A(n3), .B(N1710), .Z(n726) );
  NAND U1087 ( .A(n728), .B(n729), .Z(z3[677]) );
  NANDN U1088 ( .A(N1030), .B(z2[677]), .Z(n729) );
  NANDN U1089 ( .A(n3), .B(N1709), .Z(n728) );
  NAND U1090 ( .A(n730), .B(n731), .Z(z3[676]) );
  NANDN U1091 ( .A(N1030), .B(z2[676]), .Z(n731) );
  NANDN U1092 ( .A(n3), .B(N1708), .Z(n730) );
  NAND U1093 ( .A(n732), .B(n733), .Z(z3[675]) );
  NANDN U1094 ( .A(N1030), .B(z2[675]), .Z(n733) );
  NANDN U1095 ( .A(n3), .B(N1707), .Z(n732) );
  NAND U1096 ( .A(n734), .B(n735), .Z(z3[674]) );
  NANDN U1097 ( .A(N1030), .B(z2[674]), .Z(n735) );
  NANDN U1098 ( .A(n3), .B(N1706), .Z(n734) );
  NAND U1099 ( .A(n736), .B(n737), .Z(z3[673]) );
  NANDN U1100 ( .A(N1030), .B(z2[673]), .Z(n737) );
  NANDN U1101 ( .A(n3), .B(N1705), .Z(n736) );
  NAND U1102 ( .A(n738), .B(n739), .Z(z3[672]) );
  NANDN U1103 ( .A(N1030), .B(z2[672]), .Z(n739) );
  NANDN U1104 ( .A(n3), .B(N1704), .Z(n738) );
  NAND U1105 ( .A(n740), .B(n741), .Z(z3[671]) );
  NANDN U1106 ( .A(N1030), .B(z2[671]), .Z(n741) );
  NANDN U1107 ( .A(n3), .B(N1703), .Z(n740) );
  NAND U1108 ( .A(n742), .B(n743), .Z(z3[670]) );
  NANDN U1109 ( .A(N1030), .B(z2[670]), .Z(n743) );
  NANDN U1110 ( .A(n3), .B(N1702), .Z(n742) );
  NAND U1111 ( .A(n744), .B(n745), .Z(z3[66]) );
  NANDN U1112 ( .A(N1030), .B(z2[66]), .Z(n745) );
  NANDN U1113 ( .A(n3), .B(N1098), .Z(n744) );
  NAND U1114 ( .A(n746), .B(n747), .Z(z3[669]) );
  NANDN U1115 ( .A(N1030), .B(z2[669]), .Z(n747) );
  NANDN U1116 ( .A(n3), .B(N1701), .Z(n746) );
  NAND U1117 ( .A(n748), .B(n749), .Z(z3[668]) );
  NANDN U1118 ( .A(N1030), .B(z2[668]), .Z(n749) );
  NANDN U1119 ( .A(n3), .B(N1700), .Z(n748) );
  NAND U1120 ( .A(n750), .B(n751), .Z(z3[667]) );
  NANDN U1121 ( .A(N1030), .B(z2[667]), .Z(n751) );
  NANDN U1122 ( .A(n3), .B(N1699), .Z(n750) );
  NAND U1123 ( .A(n752), .B(n753), .Z(z3[666]) );
  NANDN U1124 ( .A(N1030), .B(z2[666]), .Z(n753) );
  NANDN U1125 ( .A(n3), .B(N1698), .Z(n752) );
  NAND U1126 ( .A(n754), .B(n755), .Z(z3[665]) );
  NANDN U1127 ( .A(N1030), .B(z2[665]), .Z(n755) );
  NANDN U1128 ( .A(n3), .B(N1697), .Z(n754) );
  NAND U1129 ( .A(n756), .B(n757), .Z(z3[664]) );
  NANDN U1130 ( .A(N1030), .B(z2[664]), .Z(n757) );
  NANDN U1131 ( .A(n3), .B(N1696), .Z(n756) );
  NAND U1132 ( .A(n758), .B(n759), .Z(z3[663]) );
  NANDN U1133 ( .A(N1030), .B(z2[663]), .Z(n759) );
  NANDN U1134 ( .A(n3), .B(N1695), .Z(n758) );
  NAND U1135 ( .A(n760), .B(n761), .Z(z3[662]) );
  NANDN U1136 ( .A(N1030), .B(z2[662]), .Z(n761) );
  NANDN U1137 ( .A(n3), .B(N1694), .Z(n760) );
  NAND U1138 ( .A(n762), .B(n763), .Z(z3[661]) );
  NANDN U1139 ( .A(N1030), .B(z2[661]), .Z(n763) );
  NANDN U1140 ( .A(n3), .B(N1693), .Z(n762) );
  NAND U1141 ( .A(n764), .B(n765), .Z(z3[660]) );
  NANDN U1142 ( .A(N1030), .B(z2[660]), .Z(n765) );
  NANDN U1143 ( .A(n3), .B(N1692), .Z(n764) );
  NAND U1144 ( .A(n766), .B(n767), .Z(z3[65]) );
  NANDN U1145 ( .A(N1030), .B(z2[65]), .Z(n767) );
  NANDN U1146 ( .A(n3), .B(N1097), .Z(n766) );
  NAND U1147 ( .A(n768), .B(n769), .Z(z3[659]) );
  NANDN U1148 ( .A(N1030), .B(z2[659]), .Z(n769) );
  NANDN U1149 ( .A(n3), .B(N1691), .Z(n768) );
  NAND U1150 ( .A(n770), .B(n771), .Z(z3[658]) );
  NANDN U1151 ( .A(N1030), .B(z2[658]), .Z(n771) );
  NANDN U1152 ( .A(n3), .B(N1690), .Z(n770) );
  NAND U1153 ( .A(n772), .B(n773), .Z(z3[657]) );
  NANDN U1154 ( .A(N1030), .B(z2[657]), .Z(n773) );
  NANDN U1155 ( .A(n3), .B(N1689), .Z(n772) );
  NAND U1156 ( .A(n774), .B(n775), .Z(z3[656]) );
  NANDN U1157 ( .A(N1030), .B(z2[656]), .Z(n775) );
  NANDN U1158 ( .A(n3), .B(N1688), .Z(n774) );
  NAND U1159 ( .A(n776), .B(n777), .Z(z3[655]) );
  NANDN U1160 ( .A(N1030), .B(z2[655]), .Z(n777) );
  NANDN U1161 ( .A(n3), .B(N1687), .Z(n776) );
  NAND U1162 ( .A(n778), .B(n779), .Z(z3[654]) );
  NANDN U1163 ( .A(N1030), .B(z2[654]), .Z(n779) );
  NANDN U1164 ( .A(n3), .B(N1686), .Z(n778) );
  NAND U1165 ( .A(n780), .B(n781), .Z(z3[653]) );
  NANDN U1166 ( .A(N1030), .B(z2[653]), .Z(n781) );
  NANDN U1167 ( .A(n3), .B(N1685), .Z(n780) );
  NAND U1168 ( .A(n782), .B(n783), .Z(z3[652]) );
  NANDN U1169 ( .A(N1030), .B(z2[652]), .Z(n783) );
  NANDN U1170 ( .A(n3), .B(N1684), .Z(n782) );
  NAND U1171 ( .A(n784), .B(n785), .Z(z3[651]) );
  NANDN U1172 ( .A(N1030), .B(z2[651]), .Z(n785) );
  NANDN U1173 ( .A(n3), .B(N1683), .Z(n784) );
  NAND U1174 ( .A(n786), .B(n787), .Z(z3[650]) );
  NANDN U1175 ( .A(N1030), .B(z2[650]), .Z(n787) );
  NANDN U1176 ( .A(n3), .B(N1682), .Z(n786) );
  NAND U1177 ( .A(n788), .B(n789), .Z(z3[64]) );
  NANDN U1178 ( .A(N1030), .B(z2[64]), .Z(n789) );
  NANDN U1179 ( .A(n3), .B(N1096), .Z(n788) );
  NAND U1180 ( .A(n790), .B(n791), .Z(z3[649]) );
  NANDN U1181 ( .A(N1030), .B(z2[649]), .Z(n791) );
  NANDN U1182 ( .A(n3), .B(N1681), .Z(n790) );
  NAND U1183 ( .A(n792), .B(n793), .Z(z3[648]) );
  NANDN U1184 ( .A(N1030), .B(z2[648]), .Z(n793) );
  NANDN U1185 ( .A(n3), .B(N1680), .Z(n792) );
  NAND U1186 ( .A(n794), .B(n795), .Z(z3[647]) );
  NANDN U1187 ( .A(N1030), .B(z2[647]), .Z(n795) );
  NANDN U1188 ( .A(n3), .B(N1679), .Z(n794) );
  NAND U1189 ( .A(n796), .B(n797), .Z(z3[646]) );
  NANDN U1190 ( .A(N1030), .B(z2[646]), .Z(n797) );
  NANDN U1191 ( .A(n3), .B(N1678), .Z(n796) );
  NAND U1192 ( .A(n798), .B(n799), .Z(z3[645]) );
  NANDN U1193 ( .A(N1030), .B(z2[645]), .Z(n799) );
  NANDN U1194 ( .A(n3), .B(N1677), .Z(n798) );
  NAND U1195 ( .A(n800), .B(n801), .Z(z3[644]) );
  NANDN U1196 ( .A(N1030), .B(z2[644]), .Z(n801) );
  NANDN U1197 ( .A(n3), .B(N1676), .Z(n800) );
  NAND U1198 ( .A(n802), .B(n803), .Z(z3[643]) );
  NANDN U1199 ( .A(N1030), .B(z2[643]), .Z(n803) );
  NANDN U1200 ( .A(n3), .B(N1675), .Z(n802) );
  NAND U1201 ( .A(n804), .B(n805), .Z(z3[642]) );
  NANDN U1202 ( .A(N1030), .B(z2[642]), .Z(n805) );
  NANDN U1203 ( .A(n3), .B(N1674), .Z(n804) );
  NAND U1204 ( .A(n806), .B(n807), .Z(z3[641]) );
  NANDN U1205 ( .A(N1030), .B(z2[641]), .Z(n807) );
  NANDN U1206 ( .A(n3), .B(N1673), .Z(n806) );
  NAND U1207 ( .A(n808), .B(n809), .Z(z3[640]) );
  NANDN U1208 ( .A(N1030), .B(z2[640]), .Z(n809) );
  NANDN U1209 ( .A(n3), .B(N1672), .Z(n808) );
  NAND U1210 ( .A(n810), .B(n811), .Z(z3[63]) );
  NANDN U1211 ( .A(N1030), .B(z2[63]), .Z(n811) );
  NANDN U1212 ( .A(n3), .B(N1095), .Z(n810) );
  NAND U1213 ( .A(n812), .B(n813), .Z(z3[639]) );
  NANDN U1214 ( .A(N1030), .B(z2[639]), .Z(n813) );
  NANDN U1215 ( .A(n3), .B(N1671), .Z(n812) );
  NAND U1216 ( .A(n814), .B(n815), .Z(z3[638]) );
  NANDN U1217 ( .A(N1030), .B(z2[638]), .Z(n815) );
  NANDN U1218 ( .A(n3), .B(N1670), .Z(n814) );
  NAND U1219 ( .A(n816), .B(n817), .Z(z3[637]) );
  NANDN U1220 ( .A(N1030), .B(z2[637]), .Z(n817) );
  NANDN U1221 ( .A(n3), .B(N1669), .Z(n816) );
  NAND U1222 ( .A(n818), .B(n819), .Z(z3[636]) );
  NANDN U1223 ( .A(N1030), .B(z2[636]), .Z(n819) );
  NANDN U1224 ( .A(n3), .B(N1668), .Z(n818) );
  NAND U1225 ( .A(n820), .B(n821), .Z(z3[635]) );
  NANDN U1226 ( .A(N1030), .B(z2[635]), .Z(n821) );
  NANDN U1227 ( .A(n3), .B(N1667), .Z(n820) );
  NAND U1228 ( .A(n822), .B(n823), .Z(z3[634]) );
  NANDN U1229 ( .A(N1030), .B(z2[634]), .Z(n823) );
  NANDN U1230 ( .A(n3), .B(N1666), .Z(n822) );
  NAND U1231 ( .A(n824), .B(n825), .Z(z3[633]) );
  NANDN U1232 ( .A(N1030), .B(z2[633]), .Z(n825) );
  NANDN U1233 ( .A(n3), .B(N1665), .Z(n824) );
  NAND U1234 ( .A(n826), .B(n827), .Z(z3[632]) );
  NANDN U1235 ( .A(N1030), .B(z2[632]), .Z(n827) );
  NANDN U1236 ( .A(n3), .B(N1664), .Z(n826) );
  NAND U1237 ( .A(n828), .B(n829), .Z(z3[631]) );
  NANDN U1238 ( .A(N1030), .B(z2[631]), .Z(n829) );
  NANDN U1239 ( .A(n3), .B(N1663), .Z(n828) );
  NAND U1240 ( .A(n830), .B(n831), .Z(z3[630]) );
  NANDN U1241 ( .A(N1030), .B(z2[630]), .Z(n831) );
  NANDN U1242 ( .A(n3), .B(N1662), .Z(n830) );
  NAND U1243 ( .A(n832), .B(n833), .Z(z3[62]) );
  NANDN U1244 ( .A(N1030), .B(z2[62]), .Z(n833) );
  NANDN U1245 ( .A(n3), .B(N1094), .Z(n832) );
  NAND U1246 ( .A(n834), .B(n835), .Z(z3[629]) );
  NANDN U1247 ( .A(N1030), .B(z2[629]), .Z(n835) );
  NANDN U1248 ( .A(n3), .B(N1661), .Z(n834) );
  NAND U1249 ( .A(n836), .B(n837), .Z(z3[628]) );
  NANDN U1250 ( .A(N1030), .B(z2[628]), .Z(n837) );
  NANDN U1251 ( .A(n3), .B(N1660), .Z(n836) );
  NAND U1252 ( .A(n838), .B(n839), .Z(z3[627]) );
  NANDN U1253 ( .A(N1030), .B(z2[627]), .Z(n839) );
  NANDN U1254 ( .A(n3), .B(N1659), .Z(n838) );
  NAND U1255 ( .A(n840), .B(n841), .Z(z3[626]) );
  NANDN U1256 ( .A(N1030), .B(z2[626]), .Z(n841) );
  NANDN U1257 ( .A(n3), .B(N1658), .Z(n840) );
  NAND U1258 ( .A(n842), .B(n843), .Z(z3[625]) );
  NANDN U1259 ( .A(N1030), .B(z2[625]), .Z(n843) );
  NANDN U1260 ( .A(n3), .B(N1657), .Z(n842) );
  NAND U1261 ( .A(n844), .B(n845), .Z(z3[624]) );
  NANDN U1262 ( .A(N1030), .B(z2[624]), .Z(n845) );
  NANDN U1263 ( .A(n3), .B(N1656), .Z(n844) );
  NAND U1264 ( .A(n846), .B(n847), .Z(z3[623]) );
  NANDN U1265 ( .A(N1030), .B(z2[623]), .Z(n847) );
  NANDN U1266 ( .A(n3), .B(N1655), .Z(n846) );
  NAND U1267 ( .A(n848), .B(n849), .Z(z3[622]) );
  NANDN U1268 ( .A(N1030), .B(z2[622]), .Z(n849) );
  NANDN U1269 ( .A(n3), .B(N1654), .Z(n848) );
  NAND U1270 ( .A(n850), .B(n851), .Z(z3[621]) );
  NANDN U1271 ( .A(N1030), .B(z2[621]), .Z(n851) );
  NANDN U1272 ( .A(n3), .B(N1653), .Z(n850) );
  NAND U1273 ( .A(n852), .B(n853), .Z(z3[620]) );
  NANDN U1274 ( .A(N1030), .B(z2[620]), .Z(n853) );
  NANDN U1275 ( .A(n3), .B(N1652), .Z(n852) );
  NAND U1276 ( .A(n854), .B(n855), .Z(z3[61]) );
  NANDN U1277 ( .A(N1030), .B(z2[61]), .Z(n855) );
  NANDN U1278 ( .A(n3), .B(N1093), .Z(n854) );
  NAND U1279 ( .A(n856), .B(n857), .Z(z3[619]) );
  NANDN U1280 ( .A(N1030), .B(z2[619]), .Z(n857) );
  NANDN U1281 ( .A(n3), .B(N1651), .Z(n856) );
  NAND U1282 ( .A(n858), .B(n859), .Z(z3[618]) );
  NANDN U1283 ( .A(N1030), .B(z2[618]), .Z(n859) );
  NANDN U1284 ( .A(n3), .B(N1650), .Z(n858) );
  NAND U1285 ( .A(n860), .B(n861), .Z(z3[617]) );
  NANDN U1286 ( .A(N1030), .B(z2[617]), .Z(n861) );
  NANDN U1287 ( .A(n3), .B(N1649), .Z(n860) );
  NAND U1288 ( .A(n862), .B(n863), .Z(z3[616]) );
  NANDN U1289 ( .A(N1030), .B(z2[616]), .Z(n863) );
  NANDN U1290 ( .A(n3), .B(N1648), .Z(n862) );
  NAND U1291 ( .A(n864), .B(n865), .Z(z3[615]) );
  NANDN U1292 ( .A(N1030), .B(z2[615]), .Z(n865) );
  NANDN U1293 ( .A(n3), .B(N1647), .Z(n864) );
  NAND U1294 ( .A(n866), .B(n867), .Z(z3[614]) );
  NANDN U1295 ( .A(N1030), .B(z2[614]), .Z(n867) );
  NANDN U1296 ( .A(n3), .B(N1646), .Z(n866) );
  NAND U1297 ( .A(n868), .B(n869), .Z(z3[613]) );
  NANDN U1298 ( .A(N1030), .B(z2[613]), .Z(n869) );
  NANDN U1299 ( .A(n3), .B(N1645), .Z(n868) );
  NAND U1300 ( .A(n870), .B(n871), .Z(z3[612]) );
  NANDN U1301 ( .A(N1030), .B(z2[612]), .Z(n871) );
  NANDN U1302 ( .A(n3), .B(N1644), .Z(n870) );
  NAND U1303 ( .A(n872), .B(n873), .Z(z3[611]) );
  NANDN U1304 ( .A(N1030), .B(z2[611]), .Z(n873) );
  NANDN U1305 ( .A(n3), .B(N1643), .Z(n872) );
  NAND U1306 ( .A(n874), .B(n875), .Z(z3[610]) );
  NANDN U1307 ( .A(N1030), .B(z2[610]), .Z(n875) );
  NANDN U1308 ( .A(n3), .B(N1642), .Z(n874) );
  NAND U1309 ( .A(n876), .B(n877), .Z(z3[60]) );
  NANDN U1310 ( .A(N1030), .B(z2[60]), .Z(n877) );
  NANDN U1311 ( .A(n3), .B(N1092), .Z(n876) );
  NAND U1312 ( .A(n878), .B(n879), .Z(z3[609]) );
  NANDN U1313 ( .A(N1030), .B(z2[609]), .Z(n879) );
  NANDN U1314 ( .A(n3), .B(N1641), .Z(n878) );
  NAND U1315 ( .A(n880), .B(n881), .Z(z3[608]) );
  NANDN U1316 ( .A(N1030), .B(z2[608]), .Z(n881) );
  NANDN U1317 ( .A(n3), .B(N1640), .Z(n880) );
  NAND U1318 ( .A(n882), .B(n883), .Z(z3[607]) );
  NANDN U1319 ( .A(N1030), .B(z2[607]), .Z(n883) );
  NANDN U1320 ( .A(n3), .B(N1639), .Z(n882) );
  NAND U1321 ( .A(n884), .B(n885), .Z(z3[606]) );
  NANDN U1322 ( .A(N1030), .B(z2[606]), .Z(n885) );
  NANDN U1323 ( .A(n3), .B(N1638), .Z(n884) );
  NAND U1324 ( .A(n886), .B(n887), .Z(z3[605]) );
  NANDN U1325 ( .A(N1030), .B(z2[605]), .Z(n887) );
  NANDN U1326 ( .A(n3), .B(N1637), .Z(n886) );
  NAND U1327 ( .A(n888), .B(n889), .Z(z3[604]) );
  NANDN U1328 ( .A(N1030), .B(z2[604]), .Z(n889) );
  NANDN U1329 ( .A(n3), .B(N1636), .Z(n888) );
  NAND U1330 ( .A(n890), .B(n891), .Z(z3[603]) );
  NANDN U1331 ( .A(N1030), .B(z2[603]), .Z(n891) );
  NANDN U1332 ( .A(n3), .B(N1635), .Z(n890) );
  NAND U1333 ( .A(n892), .B(n893), .Z(z3[602]) );
  NANDN U1334 ( .A(N1030), .B(z2[602]), .Z(n893) );
  NANDN U1335 ( .A(n3), .B(N1634), .Z(n892) );
  NAND U1336 ( .A(n894), .B(n895), .Z(z3[601]) );
  NANDN U1337 ( .A(N1030), .B(z2[601]), .Z(n895) );
  NANDN U1338 ( .A(n3), .B(N1633), .Z(n894) );
  NAND U1339 ( .A(n896), .B(n897), .Z(z3[600]) );
  NANDN U1340 ( .A(N1030), .B(z2[600]), .Z(n897) );
  NANDN U1341 ( .A(n3), .B(N1632), .Z(n896) );
  NAND U1342 ( .A(n898), .B(n899), .Z(z3[5]) );
  NANDN U1343 ( .A(N1030), .B(z2[5]), .Z(n899) );
  NANDN U1344 ( .A(n3), .B(N1037), .Z(n898) );
  NAND U1345 ( .A(n900), .B(n901), .Z(z3[59]) );
  NANDN U1346 ( .A(N1030), .B(z2[59]), .Z(n901) );
  NANDN U1347 ( .A(n3), .B(N1091), .Z(n900) );
  NAND U1348 ( .A(n902), .B(n903), .Z(z3[599]) );
  NANDN U1349 ( .A(N1030), .B(z2[599]), .Z(n903) );
  NANDN U1350 ( .A(n3), .B(N1631), .Z(n902) );
  NAND U1351 ( .A(n904), .B(n905), .Z(z3[598]) );
  NANDN U1352 ( .A(N1030), .B(z2[598]), .Z(n905) );
  NANDN U1353 ( .A(n3), .B(N1630), .Z(n904) );
  NAND U1354 ( .A(n906), .B(n907), .Z(z3[597]) );
  NANDN U1355 ( .A(N1030), .B(z2[597]), .Z(n907) );
  NANDN U1356 ( .A(n3), .B(N1629), .Z(n906) );
  NAND U1357 ( .A(n908), .B(n909), .Z(z3[596]) );
  NANDN U1358 ( .A(N1030), .B(z2[596]), .Z(n909) );
  NANDN U1359 ( .A(n3), .B(N1628), .Z(n908) );
  NAND U1360 ( .A(n910), .B(n911), .Z(z3[595]) );
  NANDN U1361 ( .A(N1030), .B(z2[595]), .Z(n911) );
  NANDN U1362 ( .A(n3), .B(N1627), .Z(n910) );
  NAND U1363 ( .A(n912), .B(n913), .Z(z3[594]) );
  NANDN U1364 ( .A(N1030), .B(z2[594]), .Z(n913) );
  NANDN U1365 ( .A(n3), .B(N1626), .Z(n912) );
  NAND U1366 ( .A(n914), .B(n915), .Z(z3[593]) );
  NANDN U1367 ( .A(N1030), .B(z2[593]), .Z(n915) );
  NANDN U1368 ( .A(n3), .B(N1625), .Z(n914) );
  NAND U1369 ( .A(n916), .B(n917), .Z(z3[592]) );
  NANDN U1370 ( .A(N1030), .B(z2[592]), .Z(n917) );
  NANDN U1371 ( .A(n3), .B(N1624), .Z(n916) );
  NAND U1372 ( .A(n918), .B(n919), .Z(z3[591]) );
  NANDN U1373 ( .A(N1030), .B(z2[591]), .Z(n919) );
  NANDN U1374 ( .A(n3), .B(N1623), .Z(n918) );
  NAND U1375 ( .A(n920), .B(n921), .Z(z3[590]) );
  NANDN U1376 ( .A(N1030), .B(z2[590]), .Z(n921) );
  NANDN U1377 ( .A(n3), .B(N1622), .Z(n920) );
  NAND U1378 ( .A(n922), .B(n923), .Z(z3[58]) );
  NANDN U1379 ( .A(N1030), .B(z2[58]), .Z(n923) );
  NANDN U1380 ( .A(n3), .B(N1090), .Z(n922) );
  NAND U1381 ( .A(n924), .B(n925), .Z(z3[589]) );
  NANDN U1382 ( .A(N1030), .B(z2[589]), .Z(n925) );
  NANDN U1383 ( .A(n3), .B(N1621), .Z(n924) );
  NAND U1384 ( .A(n926), .B(n927), .Z(z3[588]) );
  NANDN U1385 ( .A(N1030), .B(z2[588]), .Z(n927) );
  NANDN U1386 ( .A(n3), .B(N1620), .Z(n926) );
  NAND U1387 ( .A(n928), .B(n929), .Z(z3[587]) );
  NANDN U1388 ( .A(N1030), .B(z2[587]), .Z(n929) );
  NANDN U1389 ( .A(n3), .B(N1619), .Z(n928) );
  NAND U1390 ( .A(n930), .B(n931), .Z(z3[586]) );
  NANDN U1391 ( .A(N1030), .B(z2[586]), .Z(n931) );
  NANDN U1392 ( .A(n3), .B(N1618), .Z(n930) );
  NAND U1393 ( .A(n932), .B(n933), .Z(z3[585]) );
  NANDN U1394 ( .A(N1030), .B(z2[585]), .Z(n933) );
  NANDN U1395 ( .A(n3), .B(N1617), .Z(n932) );
  NAND U1396 ( .A(n934), .B(n935), .Z(z3[584]) );
  NANDN U1397 ( .A(N1030), .B(z2[584]), .Z(n935) );
  NANDN U1398 ( .A(n3), .B(N1616), .Z(n934) );
  NAND U1399 ( .A(n936), .B(n937), .Z(z3[583]) );
  NANDN U1400 ( .A(N1030), .B(z2[583]), .Z(n937) );
  NANDN U1401 ( .A(n3), .B(N1615), .Z(n936) );
  NAND U1402 ( .A(n938), .B(n939), .Z(z3[582]) );
  NANDN U1403 ( .A(N1030), .B(z2[582]), .Z(n939) );
  NANDN U1404 ( .A(n3), .B(N1614), .Z(n938) );
  NAND U1405 ( .A(n940), .B(n941), .Z(z3[581]) );
  NANDN U1406 ( .A(N1030), .B(z2[581]), .Z(n941) );
  NANDN U1407 ( .A(n3), .B(N1613), .Z(n940) );
  NAND U1408 ( .A(n942), .B(n943), .Z(z3[580]) );
  NANDN U1409 ( .A(N1030), .B(z2[580]), .Z(n943) );
  NANDN U1410 ( .A(n3), .B(N1612), .Z(n942) );
  NAND U1411 ( .A(n944), .B(n945), .Z(z3[57]) );
  NANDN U1412 ( .A(N1030), .B(z2[57]), .Z(n945) );
  NANDN U1413 ( .A(n3), .B(N1089), .Z(n944) );
  NAND U1414 ( .A(n946), .B(n947), .Z(z3[579]) );
  NANDN U1415 ( .A(N1030), .B(z2[579]), .Z(n947) );
  NANDN U1416 ( .A(n3), .B(N1611), .Z(n946) );
  NAND U1417 ( .A(n948), .B(n949), .Z(z3[578]) );
  NANDN U1418 ( .A(N1030), .B(z2[578]), .Z(n949) );
  NANDN U1419 ( .A(n3), .B(N1610), .Z(n948) );
  NAND U1420 ( .A(n950), .B(n951), .Z(z3[577]) );
  NANDN U1421 ( .A(N1030), .B(z2[577]), .Z(n951) );
  NANDN U1422 ( .A(n3), .B(N1609), .Z(n950) );
  NAND U1423 ( .A(n952), .B(n953), .Z(z3[576]) );
  NANDN U1424 ( .A(N1030), .B(z2[576]), .Z(n953) );
  NANDN U1425 ( .A(n3), .B(N1608), .Z(n952) );
  NAND U1426 ( .A(n954), .B(n955), .Z(z3[575]) );
  NANDN U1427 ( .A(N1030), .B(z2[575]), .Z(n955) );
  NANDN U1428 ( .A(n3), .B(N1607), .Z(n954) );
  NAND U1429 ( .A(n956), .B(n957), .Z(z3[574]) );
  NANDN U1430 ( .A(N1030), .B(z2[574]), .Z(n957) );
  NANDN U1431 ( .A(n3), .B(N1606), .Z(n956) );
  NAND U1432 ( .A(n958), .B(n959), .Z(z3[573]) );
  NANDN U1433 ( .A(N1030), .B(z2[573]), .Z(n959) );
  NANDN U1434 ( .A(n3), .B(N1605), .Z(n958) );
  NAND U1435 ( .A(n960), .B(n961), .Z(z3[572]) );
  NANDN U1436 ( .A(N1030), .B(z2[572]), .Z(n961) );
  NANDN U1437 ( .A(n3), .B(N1604), .Z(n960) );
  NAND U1438 ( .A(n962), .B(n963), .Z(z3[571]) );
  NANDN U1439 ( .A(N1030), .B(z2[571]), .Z(n963) );
  NANDN U1440 ( .A(n3), .B(N1603), .Z(n962) );
  NAND U1441 ( .A(n964), .B(n965), .Z(z3[570]) );
  NANDN U1442 ( .A(N1030), .B(z2[570]), .Z(n965) );
  NANDN U1443 ( .A(n3), .B(N1602), .Z(n964) );
  NAND U1444 ( .A(n966), .B(n967), .Z(z3[56]) );
  NANDN U1445 ( .A(N1030), .B(z2[56]), .Z(n967) );
  NANDN U1446 ( .A(n3), .B(N1088), .Z(n966) );
  NAND U1447 ( .A(n968), .B(n969), .Z(z3[569]) );
  NANDN U1448 ( .A(N1030), .B(z2[569]), .Z(n969) );
  NANDN U1449 ( .A(n3), .B(N1601), .Z(n968) );
  NAND U1450 ( .A(n970), .B(n971), .Z(z3[568]) );
  NANDN U1451 ( .A(N1030), .B(z2[568]), .Z(n971) );
  NANDN U1452 ( .A(n3), .B(N1600), .Z(n970) );
  NAND U1453 ( .A(n972), .B(n973), .Z(z3[567]) );
  NANDN U1454 ( .A(N1030), .B(z2[567]), .Z(n973) );
  NANDN U1455 ( .A(n3), .B(N1599), .Z(n972) );
  NAND U1456 ( .A(n974), .B(n975), .Z(z3[566]) );
  NANDN U1457 ( .A(N1030), .B(z2[566]), .Z(n975) );
  NANDN U1458 ( .A(n3), .B(N1598), .Z(n974) );
  NAND U1459 ( .A(n976), .B(n977), .Z(z3[565]) );
  NANDN U1460 ( .A(N1030), .B(z2[565]), .Z(n977) );
  NANDN U1461 ( .A(n3), .B(N1597), .Z(n976) );
  NAND U1462 ( .A(n978), .B(n979), .Z(z3[564]) );
  NANDN U1463 ( .A(N1030), .B(z2[564]), .Z(n979) );
  NANDN U1464 ( .A(n3), .B(N1596), .Z(n978) );
  NAND U1465 ( .A(n980), .B(n981), .Z(z3[563]) );
  NANDN U1466 ( .A(N1030), .B(z2[563]), .Z(n981) );
  NANDN U1467 ( .A(n3), .B(N1595), .Z(n980) );
  NAND U1468 ( .A(n982), .B(n983), .Z(z3[562]) );
  NANDN U1469 ( .A(N1030), .B(z2[562]), .Z(n983) );
  NANDN U1470 ( .A(n3), .B(N1594), .Z(n982) );
  NAND U1471 ( .A(n984), .B(n985), .Z(z3[561]) );
  NANDN U1472 ( .A(N1030), .B(z2[561]), .Z(n985) );
  NANDN U1473 ( .A(n3), .B(N1593), .Z(n984) );
  NAND U1474 ( .A(n986), .B(n987), .Z(z3[560]) );
  NANDN U1475 ( .A(N1030), .B(z2[560]), .Z(n987) );
  NANDN U1476 ( .A(n3), .B(N1592), .Z(n986) );
  NAND U1477 ( .A(n988), .B(n989), .Z(z3[55]) );
  NANDN U1478 ( .A(N1030), .B(z2[55]), .Z(n989) );
  NANDN U1479 ( .A(n3), .B(N1087), .Z(n988) );
  NAND U1480 ( .A(n990), .B(n991), .Z(z3[559]) );
  NANDN U1481 ( .A(N1030), .B(z2[559]), .Z(n991) );
  NANDN U1482 ( .A(n3), .B(N1591), .Z(n990) );
  NAND U1483 ( .A(n992), .B(n993), .Z(z3[558]) );
  NANDN U1484 ( .A(N1030), .B(z2[558]), .Z(n993) );
  NANDN U1485 ( .A(n3), .B(N1590), .Z(n992) );
  NAND U1486 ( .A(n994), .B(n995), .Z(z3[557]) );
  NANDN U1487 ( .A(N1030), .B(z2[557]), .Z(n995) );
  NANDN U1488 ( .A(n3), .B(N1589), .Z(n994) );
  NAND U1489 ( .A(n996), .B(n997), .Z(z3[556]) );
  NANDN U1490 ( .A(N1030), .B(z2[556]), .Z(n997) );
  NANDN U1491 ( .A(n3), .B(N1588), .Z(n996) );
  NAND U1492 ( .A(n998), .B(n999), .Z(z3[555]) );
  NANDN U1493 ( .A(N1030), .B(z2[555]), .Z(n999) );
  NANDN U1494 ( .A(n3), .B(N1587), .Z(n998) );
  NAND U1495 ( .A(n1000), .B(n1001), .Z(z3[554]) );
  NANDN U1496 ( .A(N1030), .B(z2[554]), .Z(n1001) );
  NANDN U1497 ( .A(n3), .B(N1586), .Z(n1000) );
  NAND U1498 ( .A(n1002), .B(n1003), .Z(z3[553]) );
  NANDN U1499 ( .A(N1030), .B(z2[553]), .Z(n1003) );
  NANDN U1500 ( .A(n3), .B(N1585), .Z(n1002) );
  NAND U1501 ( .A(n1004), .B(n1005), .Z(z3[552]) );
  NANDN U1502 ( .A(N1030), .B(z2[552]), .Z(n1005) );
  NANDN U1503 ( .A(n3), .B(N1584), .Z(n1004) );
  NAND U1504 ( .A(n1006), .B(n1007), .Z(z3[551]) );
  NANDN U1505 ( .A(N1030), .B(z2[551]), .Z(n1007) );
  NANDN U1506 ( .A(n3), .B(N1583), .Z(n1006) );
  NAND U1507 ( .A(n1008), .B(n1009), .Z(z3[550]) );
  NANDN U1508 ( .A(N1030), .B(z2[550]), .Z(n1009) );
  NANDN U1509 ( .A(n3), .B(N1582), .Z(n1008) );
  NAND U1510 ( .A(n1010), .B(n1011), .Z(z3[54]) );
  NANDN U1511 ( .A(N1030), .B(z2[54]), .Z(n1011) );
  NANDN U1512 ( .A(n3), .B(N1086), .Z(n1010) );
  NAND U1513 ( .A(n1012), .B(n1013), .Z(z3[549]) );
  NANDN U1514 ( .A(N1030), .B(z2[549]), .Z(n1013) );
  NANDN U1515 ( .A(n3), .B(N1581), .Z(n1012) );
  NAND U1516 ( .A(n1014), .B(n1015), .Z(z3[548]) );
  NANDN U1517 ( .A(N1030), .B(z2[548]), .Z(n1015) );
  NANDN U1518 ( .A(n3), .B(N1580), .Z(n1014) );
  NAND U1519 ( .A(n1016), .B(n1017), .Z(z3[547]) );
  NANDN U1520 ( .A(N1030), .B(z2[547]), .Z(n1017) );
  NANDN U1521 ( .A(n3), .B(N1579), .Z(n1016) );
  NAND U1522 ( .A(n1018), .B(n1019), .Z(z3[546]) );
  NANDN U1523 ( .A(N1030), .B(z2[546]), .Z(n1019) );
  NANDN U1524 ( .A(n3), .B(N1578), .Z(n1018) );
  NAND U1525 ( .A(n1020), .B(n1021), .Z(z3[545]) );
  NANDN U1526 ( .A(N1030), .B(z2[545]), .Z(n1021) );
  NANDN U1527 ( .A(n3), .B(N1577), .Z(n1020) );
  NAND U1528 ( .A(n1022), .B(n1023), .Z(z3[544]) );
  NANDN U1529 ( .A(N1030), .B(z2[544]), .Z(n1023) );
  NANDN U1530 ( .A(n3), .B(N1576), .Z(n1022) );
  NAND U1531 ( .A(n1024), .B(n1025), .Z(z3[543]) );
  NANDN U1532 ( .A(N1030), .B(z2[543]), .Z(n1025) );
  NANDN U1533 ( .A(n3), .B(N1575), .Z(n1024) );
  NAND U1534 ( .A(n1026), .B(n1027), .Z(z3[542]) );
  NANDN U1535 ( .A(N1030), .B(z2[542]), .Z(n1027) );
  NANDN U1536 ( .A(n3), .B(N1574), .Z(n1026) );
  NAND U1537 ( .A(n1028), .B(n1029), .Z(z3[541]) );
  NANDN U1538 ( .A(N1030), .B(z2[541]), .Z(n1029) );
  NANDN U1539 ( .A(n3), .B(N1573), .Z(n1028) );
  NAND U1540 ( .A(n1030), .B(n1031), .Z(z3[540]) );
  NANDN U1541 ( .A(N1030), .B(z2[540]), .Z(n1031) );
  NANDN U1542 ( .A(n3), .B(N1572), .Z(n1030) );
  NAND U1543 ( .A(n1032), .B(n1033), .Z(z3[53]) );
  NANDN U1544 ( .A(N1030), .B(z2[53]), .Z(n1033) );
  NANDN U1545 ( .A(n3), .B(N1085), .Z(n1032) );
  NAND U1546 ( .A(n1034), .B(n1035), .Z(z3[539]) );
  NANDN U1547 ( .A(N1030), .B(z2[539]), .Z(n1035) );
  NANDN U1548 ( .A(n3), .B(N1571), .Z(n1034) );
  NAND U1549 ( .A(n1036), .B(n1037), .Z(z3[538]) );
  NANDN U1550 ( .A(N1030), .B(z2[538]), .Z(n1037) );
  NANDN U1551 ( .A(n3), .B(N1570), .Z(n1036) );
  NAND U1552 ( .A(n1038), .B(n1039), .Z(z3[537]) );
  NANDN U1553 ( .A(N1030), .B(z2[537]), .Z(n1039) );
  NANDN U1554 ( .A(n3), .B(N1569), .Z(n1038) );
  NAND U1555 ( .A(n1040), .B(n1041), .Z(z3[536]) );
  NANDN U1556 ( .A(N1030), .B(z2[536]), .Z(n1041) );
  NANDN U1557 ( .A(n3), .B(N1568), .Z(n1040) );
  NAND U1558 ( .A(n1042), .B(n1043), .Z(z3[535]) );
  NANDN U1559 ( .A(N1030), .B(z2[535]), .Z(n1043) );
  NANDN U1560 ( .A(n3), .B(N1567), .Z(n1042) );
  NAND U1561 ( .A(n1044), .B(n1045), .Z(z3[534]) );
  NANDN U1562 ( .A(N1030), .B(z2[534]), .Z(n1045) );
  NANDN U1563 ( .A(n3), .B(N1566), .Z(n1044) );
  NAND U1564 ( .A(n1046), .B(n1047), .Z(z3[533]) );
  NANDN U1565 ( .A(N1030), .B(z2[533]), .Z(n1047) );
  NANDN U1566 ( .A(n3), .B(N1565), .Z(n1046) );
  NAND U1567 ( .A(n1048), .B(n1049), .Z(z3[532]) );
  NANDN U1568 ( .A(N1030), .B(z2[532]), .Z(n1049) );
  NANDN U1569 ( .A(n3), .B(N1564), .Z(n1048) );
  NAND U1570 ( .A(n1050), .B(n1051), .Z(z3[531]) );
  NANDN U1571 ( .A(N1030), .B(z2[531]), .Z(n1051) );
  NANDN U1572 ( .A(n3), .B(N1563), .Z(n1050) );
  NAND U1573 ( .A(n1052), .B(n1053), .Z(z3[530]) );
  NANDN U1574 ( .A(N1030), .B(z2[530]), .Z(n1053) );
  NANDN U1575 ( .A(n3), .B(N1562), .Z(n1052) );
  NAND U1576 ( .A(n1054), .B(n1055), .Z(z3[52]) );
  NANDN U1577 ( .A(N1030), .B(z2[52]), .Z(n1055) );
  NANDN U1578 ( .A(n3), .B(N1084), .Z(n1054) );
  NAND U1579 ( .A(n1056), .B(n1057), .Z(z3[529]) );
  NANDN U1580 ( .A(N1030), .B(z2[529]), .Z(n1057) );
  NANDN U1581 ( .A(n3), .B(N1561), .Z(n1056) );
  NAND U1582 ( .A(n1058), .B(n1059), .Z(z3[528]) );
  NANDN U1583 ( .A(N1030), .B(z2[528]), .Z(n1059) );
  NANDN U1584 ( .A(n3), .B(N1560), .Z(n1058) );
  NAND U1585 ( .A(n1060), .B(n1061), .Z(z3[527]) );
  NANDN U1586 ( .A(N1030), .B(z2[527]), .Z(n1061) );
  NANDN U1587 ( .A(n3), .B(N1559), .Z(n1060) );
  NAND U1588 ( .A(n1062), .B(n1063), .Z(z3[526]) );
  NANDN U1589 ( .A(N1030), .B(z2[526]), .Z(n1063) );
  NANDN U1590 ( .A(n3), .B(N1558), .Z(n1062) );
  NAND U1591 ( .A(n1064), .B(n1065), .Z(z3[525]) );
  NANDN U1592 ( .A(N1030), .B(z2[525]), .Z(n1065) );
  NANDN U1593 ( .A(n3), .B(N1557), .Z(n1064) );
  NAND U1594 ( .A(n1066), .B(n1067), .Z(z3[524]) );
  NANDN U1595 ( .A(N1030), .B(z2[524]), .Z(n1067) );
  NANDN U1596 ( .A(n3), .B(N1556), .Z(n1066) );
  NAND U1597 ( .A(n1068), .B(n1069), .Z(z3[523]) );
  NANDN U1598 ( .A(N1030), .B(z2[523]), .Z(n1069) );
  NANDN U1599 ( .A(n3), .B(N1555), .Z(n1068) );
  NAND U1600 ( .A(n1070), .B(n1071), .Z(z3[522]) );
  NANDN U1601 ( .A(N1030), .B(z2[522]), .Z(n1071) );
  NANDN U1602 ( .A(n3), .B(N1554), .Z(n1070) );
  NAND U1603 ( .A(n1072), .B(n1073), .Z(z3[521]) );
  NANDN U1604 ( .A(N1030), .B(z2[521]), .Z(n1073) );
  NANDN U1605 ( .A(n3), .B(N1553), .Z(n1072) );
  NAND U1606 ( .A(n1074), .B(n1075), .Z(z3[520]) );
  NANDN U1607 ( .A(N1030), .B(z2[520]), .Z(n1075) );
  NANDN U1608 ( .A(n3), .B(N1552), .Z(n1074) );
  NAND U1609 ( .A(n1076), .B(n1077), .Z(z3[51]) );
  NANDN U1610 ( .A(N1030), .B(z2[51]), .Z(n1077) );
  NANDN U1611 ( .A(n3), .B(N1083), .Z(n1076) );
  NAND U1612 ( .A(n1078), .B(n1079), .Z(z3[519]) );
  NANDN U1613 ( .A(N1030), .B(z2[519]), .Z(n1079) );
  NANDN U1614 ( .A(n3), .B(N1551), .Z(n1078) );
  NAND U1615 ( .A(n1080), .B(n1081), .Z(z3[518]) );
  NANDN U1616 ( .A(N1030), .B(z2[518]), .Z(n1081) );
  NANDN U1617 ( .A(n3), .B(N1550), .Z(n1080) );
  NAND U1618 ( .A(n1082), .B(n1083), .Z(z3[517]) );
  NANDN U1619 ( .A(N1030), .B(z2[517]), .Z(n1083) );
  NANDN U1620 ( .A(n3), .B(N1549), .Z(n1082) );
  NAND U1621 ( .A(n1084), .B(n1085), .Z(z3[516]) );
  NANDN U1622 ( .A(N1030), .B(z2[516]), .Z(n1085) );
  NANDN U1623 ( .A(n3), .B(N1548), .Z(n1084) );
  NAND U1624 ( .A(n1086), .B(n1087), .Z(z3[515]) );
  NANDN U1625 ( .A(N1030), .B(z2[515]), .Z(n1087) );
  NANDN U1626 ( .A(n3), .B(N1547), .Z(n1086) );
  NAND U1627 ( .A(n1088), .B(n1089), .Z(z3[514]) );
  NANDN U1628 ( .A(N1030), .B(z2[514]), .Z(n1089) );
  NANDN U1629 ( .A(n3), .B(N1546), .Z(n1088) );
  NAND U1630 ( .A(n1090), .B(n1091), .Z(z3[513]) );
  NANDN U1631 ( .A(N1030), .B(z2[513]), .Z(n1091) );
  NANDN U1632 ( .A(n3), .B(N1545), .Z(n1090) );
  NAND U1633 ( .A(n1092), .B(n1093), .Z(z3[512]) );
  NANDN U1634 ( .A(N1030), .B(z2[512]), .Z(n1093) );
  NANDN U1635 ( .A(n3), .B(N1544), .Z(n1092) );
  NAND U1636 ( .A(n1094), .B(n1095), .Z(z3[511]) );
  NANDN U1637 ( .A(N1030), .B(z2[511]), .Z(n1095) );
  NANDN U1638 ( .A(n3), .B(N1543), .Z(n1094) );
  NAND U1639 ( .A(n1096), .B(n1097), .Z(z3[510]) );
  NANDN U1640 ( .A(N1030), .B(z2[510]), .Z(n1097) );
  NANDN U1641 ( .A(n3), .B(N1542), .Z(n1096) );
  NAND U1642 ( .A(n1098), .B(n1099), .Z(z3[50]) );
  NANDN U1643 ( .A(N1030), .B(z2[50]), .Z(n1099) );
  NANDN U1644 ( .A(n3), .B(N1082), .Z(n1098) );
  NAND U1645 ( .A(n1100), .B(n1101), .Z(z3[509]) );
  NANDN U1646 ( .A(N1030), .B(z2[509]), .Z(n1101) );
  NANDN U1647 ( .A(n3), .B(N1541), .Z(n1100) );
  NAND U1648 ( .A(n1102), .B(n1103), .Z(z3[508]) );
  NANDN U1649 ( .A(N1030), .B(z2[508]), .Z(n1103) );
  NANDN U1650 ( .A(n3), .B(N1540), .Z(n1102) );
  NAND U1651 ( .A(n1104), .B(n1105), .Z(z3[507]) );
  NANDN U1652 ( .A(N1030), .B(z2[507]), .Z(n1105) );
  NANDN U1653 ( .A(n3), .B(N1539), .Z(n1104) );
  NAND U1654 ( .A(n1106), .B(n1107), .Z(z3[506]) );
  NANDN U1655 ( .A(N1030), .B(z2[506]), .Z(n1107) );
  NANDN U1656 ( .A(n3), .B(N1538), .Z(n1106) );
  NAND U1657 ( .A(n1108), .B(n1109), .Z(z3[505]) );
  NANDN U1658 ( .A(N1030), .B(z2[505]), .Z(n1109) );
  NANDN U1659 ( .A(n3), .B(N1537), .Z(n1108) );
  NAND U1660 ( .A(n1110), .B(n1111), .Z(z3[504]) );
  NANDN U1661 ( .A(N1030), .B(z2[504]), .Z(n1111) );
  NANDN U1662 ( .A(n3), .B(N1536), .Z(n1110) );
  NAND U1663 ( .A(n1112), .B(n1113), .Z(z3[503]) );
  NANDN U1664 ( .A(N1030), .B(z2[503]), .Z(n1113) );
  NANDN U1665 ( .A(n3), .B(N1535), .Z(n1112) );
  NAND U1666 ( .A(n1114), .B(n1115), .Z(z3[502]) );
  NANDN U1667 ( .A(N1030), .B(z2[502]), .Z(n1115) );
  NANDN U1668 ( .A(n3), .B(N1534), .Z(n1114) );
  NAND U1669 ( .A(n1116), .B(n1117), .Z(z3[501]) );
  NANDN U1670 ( .A(N1030), .B(z2[501]), .Z(n1117) );
  NANDN U1671 ( .A(n3), .B(N1533), .Z(n1116) );
  NAND U1672 ( .A(n1118), .B(n1119), .Z(z3[500]) );
  NANDN U1673 ( .A(N1030), .B(z2[500]), .Z(n1119) );
  NANDN U1674 ( .A(n3), .B(N1532), .Z(n1118) );
  NAND U1675 ( .A(n1120), .B(n1121), .Z(z3[4]) );
  NANDN U1676 ( .A(N1030), .B(z2[4]), .Z(n1121) );
  NANDN U1677 ( .A(n3), .B(N1036), .Z(n1120) );
  NAND U1678 ( .A(n1122), .B(n1123), .Z(z3[49]) );
  NANDN U1679 ( .A(N1030), .B(z2[49]), .Z(n1123) );
  NANDN U1680 ( .A(n3), .B(N1081), .Z(n1122) );
  NAND U1681 ( .A(n1124), .B(n1125), .Z(z3[499]) );
  NANDN U1682 ( .A(N1030), .B(z2[499]), .Z(n1125) );
  NANDN U1683 ( .A(n3), .B(N1531), .Z(n1124) );
  NAND U1684 ( .A(n1126), .B(n1127), .Z(z3[498]) );
  NANDN U1685 ( .A(N1030), .B(z2[498]), .Z(n1127) );
  NANDN U1686 ( .A(n3), .B(N1530), .Z(n1126) );
  NAND U1687 ( .A(n1128), .B(n1129), .Z(z3[497]) );
  NANDN U1688 ( .A(N1030), .B(z2[497]), .Z(n1129) );
  NANDN U1689 ( .A(n3), .B(N1529), .Z(n1128) );
  NAND U1690 ( .A(n1130), .B(n1131), .Z(z3[496]) );
  NANDN U1691 ( .A(N1030), .B(z2[496]), .Z(n1131) );
  NANDN U1692 ( .A(n3), .B(N1528), .Z(n1130) );
  NAND U1693 ( .A(n1132), .B(n1133), .Z(z3[495]) );
  NANDN U1694 ( .A(N1030), .B(z2[495]), .Z(n1133) );
  NANDN U1695 ( .A(n3), .B(N1527), .Z(n1132) );
  NAND U1696 ( .A(n1134), .B(n1135), .Z(z3[494]) );
  NANDN U1697 ( .A(N1030), .B(z2[494]), .Z(n1135) );
  NANDN U1698 ( .A(n3), .B(N1526), .Z(n1134) );
  NAND U1699 ( .A(n1136), .B(n1137), .Z(z3[493]) );
  NANDN U1700 ( .A(N1030), .B(z2[493]), .Z(n1137) );
  NANDN U1701 ( .A(n3), .B(N1525), .Z(n1136) );
  NAND U1702 ( .A(n1138), .B(n1139), .Z(z3[492]) );
  NANDN U1703 ( .A(N1030), .B(z2[492]), .Z(n1139) );
  NANDN U1704 ( .A(n3), .B(N1524), .Z(n1138) );
  NAND U1705 ( .A(n1140), .B(n1141), .Z(z3[491]) );
  NANDN U1706 ( .A(N1030), .B(z2[491]), .Z(n1141) );
  NANDN U1707 ( .A(n3), .B(N1523), .Z(n1140) );
  NAND U1708 ( .A(n1142), .B(n1143), .Z(z3[490]) );
  NANDN U1709 ( .A(N1030), .B(z2[490]), .Z(n1143) );
  NANDN U1710 ( .A(n3), .B(N1522), .Z(n1142) );
  NAND U1711 ( .A(n1144), .B(n1145), .Z(z3[48]) );
  NANDN U1712 ( .A(N1030), .B(z2[48]), .Z(n1145) );
  NANDN U1713 ( .A(n3), .B(N1080), .Z(n1144) );
  NAND U1714 ( .A(n1146), .B(n1147), .Z(z3[489]) );
  NANDN U1715 ( .A(N1030), .B(z2[489]), .Z(n1147) );
  NANDN U1716 ( .A(n3), .B(N1521), .Z(n1146) );
  NAND U1717 ( .A(n1148), .B(n1149), .Z(z3[488]) );
  NANDN U1718 ( .A(N1030), .B(z2[488]), .Z(n1149) );
  NANDN U1719 ( .A(n3), .B(N1520), .Z(n1148) );
  NAND U1720 ( .A(n1150), .B(n1151), .Z(z3[487]) );
  NANDN U1721 ( .A(N1030), .B(z2[487]), .Z(n1151) );
  NANDN U1722 ( .A(n3), .B(N1519), .Z(n1150) );
  NAND U1723 ( .A(n1152), .B(n1153), .Z(z3[486]) );
  NANDN U1724 ( .A(N1030), .B(z2[486]), .Z(n1153) );
  NANDN U1725 ( .A(n3), .B(N1518), .Z(n1152) );
  NAND U1726 ( .A(n1154), .B(n1155), .Z(z3[485]) );
  NANDN U1727 ( .A(N1030), .B(z2[485]), .Z(n1155) );
  NANDN U1728 ( .A(n3), .B(N1517), .Z(n1154) );
  NAND U1729 ( .A(n1156), .B(n1157), .Z(z3[484]) );
  NANDN U1730 ( .A(N1030), .B(z2[484]), .Z(n1157) );
  NANDN U1731 ( .A(n3), .B(N1516), .Z(n1156) );
  NAND U1732 ( .A(n1158), .B(n1159), .Z(z3[483]) );
  NANDN U1733 ( .A(N1030), .B(z2[483]), .Z(n1159) );
  NANDN U1734 ( .A(n3), .B(N1515), .Z(n1158) );
  NAND U1735 ( .A(n1160), .B(n1161), .Z(z3[482]) );
  NANDN U1736 ( .A(N1030), .B(z2[482]), .Z(n1161) );
  NANDN U1737 ( .A(n3), .B(N1514), .Z(n1160) );
  NAND U1738 ( .A(n1162), .B(n1163), .Z(z3[481]) );
  NANDN U1739 ( .A(N1030), .B(z2[481]), .Z(n1163) );
  NANDN U1740 ( .A(n3), .B(N1513), .Z(n1162) );
  NAND U1741 ( .A(n1164), .B(n1165), .Z(z3[480]) );
  NANDN U1742 ( .A(N1030), .B(z2[480]), .Z(n1165) );
  NANDN U1743 ( .A(n3), .B(N1512), .Z(n1164) );
  NAND U1744 ( .A(n1166), .B(n1167), .Z(z3[47]) );
  NANDN U1745 ( .A(N1030), .B(z2[47]), .Z(n1167) );
  NANDN U1746 ( .A(n3), .B(N1079), .Z(n1166) );
  NAND U1747 ( .A(n1168), .B(n1169), .Z(z3[479]) );
  NANDN U1748 ( .A(N1030), .B(z2[479]), .Z(n1169) );
  NANDN U1749 ( .A(n3), .B(N1511), .Z(n1168) );
  NAND U1750 ( .A(n1170), .B(n1171), .Z(z3[478]) );
  NANDN U1751 ( .A(N1030), .B(z2[478]), .Z(n1171) );
  NANDN U1752 ( .A(n3), .B(N1510), .Z(n1170) );
  NAND U1753 ( .A(n1172), .B(n1173), .Z(z3[477]) );
  NANDN U1754 ( .A(N1030), .B(z2[477]), .Z(n1173) );
  NANDN U1755 ( .A(n3), .B(N1509), .Z(n1172) );
  NAND U1756 ( .A(n1174), .B(n1175), .Z(z3[476]) );
  NANDN U1757 ( .A(N1030), .B(z2[476]), .Z(n1175) );
  NANDN U1758 ( .A(n3), .B(N1508), .Z(n1174) );
  NAND U1759 ( .A(n1176), .B(n1177), .Z(z3[475]) );
  NANDN U1760 ( .A(N1030), .B(z2[475]), .Z(n1177) );
  NANDN U1761 ( .A(n3), .B(N1507), .Z(n1176) );
  NAND U1762 ( .A(n1178), .B(n1179), .Z(z3[474]) );
  NANDN U1763 ( .A(N1030), .B(z2[474]), .Z(n1179) );
  NANDN U1764 ( .A(n3), .B(N1506), .Z(n1178) );
  NAND U1765 ( .A(n1180), .B(n1181), .Z(z3[473]) );
  NANDN U1766 ( .A(N1030), .B(z2[473]), .Z(n1181) );
  NANDN U1767 ( .A(n3), .B(N1505), .Z(n1180) );
  NAND U1768 ( .A(n1182), .B(n1183), .Z(z3[472]) );
  NANDN U1769 ( .A(N1030), .B(z2[472]), .Z(n1183) );
  NANDN U1770 ( .A(n3), .B(N1504), .Z(n1182) );
  NAND U1771 ( .A(n1184), .B(n1185), .Z(z3[471]) );
  NANDN U1772 ( .A(N1030), .B(z2[471]), .Z(n1185) );
  NANDN U1773 ( .A(n3), .B(N1503), .Z(n1184) );
  NAND U1774 ( .A(n1186), .B(n1187), .Z(z3[470]) );
  NANDN U1775 ( .A(N1030), .B(z2[470]), .Z(n1187) );
  NANDN U1776 ( .A(n3), .B(N1502), .Z(n1186) );
  NAND U1777 ( .A(n1188), .B(n1189), .Z(z3[46]) );
  NANDN U1778 ( .A(N1030), .B(z2[46]), .Z(n1189) );
  NANDN U1779 ( .A(n3), .B(N1078), .Z(n1188) );
  NAND U1780 ( .A(n1190), .B(n1191), .Z(z3[469]) );
  NANDN U1781 ( .A(N1030), .B(z2[469]), .Z(n1191) );
  NANDN U1782 ( .A(n3), .B(N1501), .Z(n1190) );
  NAND U1783 ( .A(n1192), .B(n1193), .Z(z3[468]) );
  NANDN U1784 ( .A(N1030), .B(z2[468]), .Z(n1193) );
  NANDN U1785 ( .A(n3), .B(N1500), .Z(n1192) );
  NAND U1786 ( .A(n1194), .B(n1195), .Z(z3[467]) );
  NANDN U1787 ( .A(N1030), .B(z2[467]), .Z(n1195) );
  NANDN U1788 ( .A(n3), .B(N1499), .Z(n1194) );
  NAND U1789 ( .A(n1196), .B(n1197), .Z(z3[466]) );
  NANDN U1790 ( .A(N1030), .B(z2[466]), .Z(n1197) );
  NANDN U1791 ( .A(n3), .B(N1498), .Z(n1196) );
  NAND U1792 ( .A(n1198), .B(n1199), .Z(z3[465]) );
  NANDN U1793 ( .A(N1030), .B(z2[465]), .Z(n1199) );
  NANDN U1794 ( .A(n3), .B(N1497), .Z(n1198) );
  NAND U1795 ( .A(n1200), .B(n1201), .Z(z3[464]) );
  NANDN U1796 ( .A(N1030), .B(z2[464]), .Z(n1201) );
  NANDN U1797 ( .A(n3), .B(N1496), .Z(n1200) );
  NAND U1798 ( .A(n1202), .B(n1203), .Z(z3[463]) );
  NANDN U1799 ( .A(N1030), .B(z2[463]), .Z(n1203) );
  NANDN U1800 ( .A(n3), .B(N1495), .Z(n1202) );
  NAND U1801 ( .A(n1204), .B(n1205), .Z(z3[462]) );
  NANDN U1802 ( .A(N1030), .B(z2[462]), .Z(n1205) );
  NANDN U1803 ( .A(n3), .B(N1494), .Z(n1204) );
  NAND U1804 ( .A(n1206), .B(n1207), .Z(z3[461]) );
  NANDN U1805 ( .A(N1030), .B(z2[461]), .Z(n1207) );
  NANDN U1806 ( .A(n3), .B(N1493), .Z(n1206) );
  NAND U1807 ( .A(n1208), .B(n1209), .Z(z3[460]) );
  NANDN U1808 ( .A(N1030), .B(z2[460]), .Z(n1209) );
  NANDN U1809 ( .A(n3), .B(N1492), .Z(n1208) );
  NAND U1810 ( .A(n1210), .B(n1211), .Z(z3[45]) );
  NANDN U1811 ( .A(N1030), .B(z2[45]), .Z(n1211) );
  NANDN U1812 ( .A(n3), .B(N1077), .Z(n1210) );
  NAND U1813 ( .A(n1212), .B(n1213), .Z(z3[459]) );
  NANDN U1814 ( .A(N1030), .B(z2[459]), .Z(n1213) );
  NANDN U1815 ( .A(n3), .B(N1491), .Z(n1212) );
  NAND U1816 ( .A(n1214), .B(n1215), .Z(z3[458]) );
  NANDN U1817 ( .A(N1030), .B(z2[458]), .Z(n1215) );
  NANDN U1818 ( .A(n3), .B(N1490), .Z(n1214) );
  NAND U1819 ( .A(n1216), .B(n1217), .Z(z3[457]) );
  NANDN U1820 ( .A(N1030), .B(z2[457]), .Z(n1217) );
  NANDN U1821 ( .A(n3), .B(N1489), .Z(n1216) );
  NAND U1822 ( .A(n1218), .B(n1219), .Z(z3[456]) );
  NANDN U1823 ( .A(N1030), .B(z2[456]), .Z(n1219) );
  NANDN U1824 ( .A(n3), .B(N1488), .Z(n1218) );
  NAND U1825 ( .A(n1220), .B(n1221), .Z(z3[455]) );
  NANDN U1826 ( .A(N1030), .B(z2[455]), .Z(n1221) );
  NANDN U1827 ( .A(n3), .B(N1487), .Z(n1220) );
  NAND U1828 ( .A(n1222), .B(n1223), .Z(z3[454]) );
  NANDN U1829 ( .A(N1030), .B(z2[454]), .Z(n1223) );
  NANDN U1830 ( .A(n3), .B(N1486), .Z(n1222) );
  NAND U1831 ( .A(n1224), .B(n1225), .Z(z3[453]) );
  NANDN U1832 ( .A(N1030), .B(z2[453]), .Z(n1225) );
  NANDN U1833 ( .A(n3), .B(N1485), .Z(n1224) );
  NAND U1834 ( .A(n1226), .B(n1227), .Z(z3[452]) );
  NANDN U1835 ( .A(N1030), .B(z2[452]), .Z(n1227) );
  NANDN U1836 ( .A(n3), .B(N1484), .Z(n1226) );
  NAND U1837 ( .A(n1228), .B(n1229), .Z(z3[451]) );
  NANDN U1838 ( .A(N1030), .B(z2[451]), .Z(n1229) );
  NANDN U1839 ( .A(n3), .B(N1483), .Z(n1228) );
  NAND U1840 ( .A(n1230), .B(n1231), .Z(z3[450]) );
  NANDN U1841 ( .A(N1030), .B(z2[450]), .Z(n1231) );
  NANDN U1842 ( .A(n3), .B(N1482), .Z(n1230) );
  NAND U1843 ( .A(n1232), .B(n1233), .Z(z3[44]) );
  NANDN U1844 ( .A(N1030), .B(z2[44]), .Z(n1233) );
  NANDN U1845 ( .A(n3), .B(N1076), .Z(n1232) );
  NAND U1846 ( .A(n1234), .B(n1235), .Z(z3[449]) );
  NANDN U1847 ( .A(N1030), .B(z2[449]), .Z(n1235) );
  NANDN U1848 ( .A(n3), .B(N1481), .Z(n1234) );
  NAND U1849 ( .A(n1236), .B(n1237), .Z(z3[448]) );
  NANDN U1850 ( .A(N1030), .B(z2[448]), .Z(n1237) );
  NANDN U1851 ( .A(n3), .B(N1480), .Z(n1236) );
  NAND U1852 ( .A(n1238), .B(n1239), .Z(z3[447]) );
  NANDN U1853 ( .A(N1030), .B(z2[447]), .Z(n1239) );
  NANDN U1854 ( .A(n3), .B(N1479), .Z(n1238) );
  NAND U1855 ( .A(n1240), .B(n1241), .Z(z3[446]) );
  NANDN U1856 ( .A(N1030), .B(z2[446]), .Z(n1241) );
  NANDN U1857 ( .A(n3), .B(N1478), .Z(n1240) );
  NAND U1858 ( .A(n1242), .B(n1243), .Z(z3[445]) );
  NANDN U1859 ( .A(N1030), .B(z2[445]), .Z(n1243) );
  NANDN U1860 ( .A(n3), .B(N1477), .Z(n1242) );
  NAND U1861 ( .A(n1244), .B(n1245), .Z(z3[444]) );
  NANDN U1862 ( .A(N1030), .B(z2[444]), .Z(n1245) );
  NANDN U1863 ( .A(n3), .B(N1476), .Z(n1244) );
  NAND U1864 ( .A(n1246), .B(n1247), .Z(z3[443]) );
  NANDN U1865 ( .A(N1030), .B(z2[443]), .Z(n1247) );
  NANDN U1866 ( .A(n3), .B(N1475), .Z(n1246) );
  NAND U1867 ( .A(n1248), .B(n1249), .Z(z3[442]) );
  NANDN U1868 ( .A(N1030), .B(z2[442]), .Z(n1249) );
  NANDN U1869 ( .A(n3), .B(N1474), .Z(n1248) );
  NAND U1870 ( .A(n1250), .B(n1251), .Z(z3[441]) );
  NANDN U1871 ( .A(N1030), .B(z2[441]), .Z(n1251) );
  NANDN U1872 ( .A(n3), .B(N1473), .Z(n1250) );
  NAND U1873 ( .A(n1252), .B(n1253), .Z(z3[440]) );
  NANDN U1874 ( .A(N1030), .B(z2[440]), .Z(n1253) );
  NANDN U1875 ( .A(n3), .B(N1472), .Z(n1252) );
  NAND U1876 ( .A(n1254), .B(n1255), .Z(z3[43]) );
  NANDN U1877 ( .A(N1030), .B(z2[43]), .Z(n1255) );
  NANDN U1878 ( .A(n3), .B(N1075), .Z(n1254) );
  NAND U1879 ( .A(n1256), .B(n1257), .Z(z3[439]) );
  NANDN U1880 ( .A(N1030), .B(z2[439]), .Z(n1257) );
  NANDN U1881 ( .A(n3), .B(N1471), .Z(n1256) );
  NAND U1882 ( .A(n1258), .B(n1259), .Z(z3[438]) );
  NANDN U1883 ( .A(N1030), .B(z2[438]), .Z(n1259) );
  NANDN U1884 ( .A(n3), .B(N1470), .Z(n1258) );
  NAND U1885 ( .A(n1260), .B(n1261), .Z(z3[437]) );
  NANDN U1886 ( .A(N1030), .B(z2[437]), .Z(n1261) );
  NANDN U1887 ( .A(n3), .B(N1469), .Z(n1260) );
  NAND U1888 ( .A(n1262), .B(n1263), .Z(z3[436]) );
  NANDN U1889 ( .A(N1030), .B(z2[436]), .Z(n1263) );
  NANDN U1890 ( .A(n3), .B(N1468), .Z(n1262) );
  NAND U1891 ( .A(n1264), .B(n1265), .Z(z3[435]) );
  NANDN U1892 ( .A(N1030), .B(z2[435]), .Z(n1265) );
  NANDN U1893 ( .A(n3), .B(N1467), .Z(n1264) );
  NAND U1894 ( .A(n1266), .B(n1267), .Z(z3[434]) );
  NANDN U1895 ( .A(N1030), .B(z2[434]), .Z(n1267) );
  NANDN U1896 ( .A(n3), .B(N1466), .Z(n1266) );
  NAND U1897 ( .A(n1268), .B(n1269), .Z(z3[433]) );
  NANDN U1898 ( .A(N1030), .B(z2[433]), .Z(n1269) );
  NANDN U1899 ( .A(n3), .B(N1465), .Z(n1268) );
  NAND U1900 ( .A(n1270), .B(n1271), .Z(z3[432]) );
  NANDN U1901 ( .A(N1030), .B(z2[432]), .Z(n1271) );
  NANDN U1902 ( .A(n3), .B(N1464), .Z(n1270) );
  NAND U1903 ( .A(n1272), .B(n1273), .Z(z3[431]) );
  NANDN U1904 ( .A(N1030), .B(z2[431]), .Z(n1273) );
  NANDN U1905 ( .A(n3), .B(N1463), .Z(n1272) );
  NAND U1906 ( .A(n1274), .B(n1275), .Z(z3[430]) );
  NANDN U1907 ( .A(N1030), .B(z2[430]), .Z(n1275) );
  NANDN U1908 ( .A(n3), .B(N1462), .Z(n1274) );
  NAND U1909 ( .A(n1276), .B(n1277), .Z(z3[42]) );
  NANDN U1910 ( .A(N1030), .B(z2[42]), .Z(n1277) );
  NANDN U1911 ( .A(n3), .B(N1074), .Z(n1276) );
  NAND U1912 ( .A(n1278), .B(n1279), .Z(z3[429]) );
  NANDN U1913 ( .A(N1030), .B(z2[429]), .Z(n1279) );
  NANDN U1914 ( .A(n3), .B(N1461), .Z(n1278) );
  NAND U1915 ( .A(n1280), .B(n1281), .Z(z3[428]) );
  NANDN U1916 ( .A(N1030), .B(z2[428]), .Z(n1281) );
  NANDN U1917 ( .A(n3), .B(N1460), .Z(n1280) );
  NAND U1918 ( .A(n1282), .B(n1283), .Z(z3[427]) );
  NANDN U1919 ( .A(N1030), .B(z2[427]), .Z(n1283) );
  NANDN U1920 ( .A(n3), .B(N1459), .Z(n1282) );
  NAND U1921 ( .A(n1284), .B(n1285), .Z(z3[426]) );
  NANDN U1922 ( .A(N1030), .B(z2[426]), .Z(n1285) );
  NANDN U1923 ( .A(n3), .B(N1458), .Z(n1284) );
  NAND U1924 ( .A(n1286), .B(n1287), .Z(z3[425]) );
  NANDN U1925 ( .A(N1030), .B(z2[425]), .Z(n1287) );
  NANDN U1926 ( .A(n3), .B(N1457), .Z(n1286) );
  NAND U1927 ( .A(n1288), .B(n1289), .Z(z3[424]) );
  NANDN U1928 ( .A(N1030), .B(z2[424]), .Z(n1289) );
  NANDN U1929 ( .A(n3), .B(N1456), .Z(n1288) );
  NAND U1930 ( .A(n1290), .B(n1291), .Z(z3[423]) );
  NANDN U1931 ( .A(N1030), .B(z2[423]), .Z(n1291) );
  NANDN U1932 ( .A(n3), .B(N1455), .Z(n1290) );
  NAND U1933 ( .A(n1292), .B(n1293), .Z(z3[422]) );
  NANDN U1934 ( .A(N1030), .B(z2[422]), .Z(n1293) );
  NANDN U1935 ( .A(n3), .B(N1454), .Z(n1292) );
  NAND U1936 ( .A(n1294), .B(n1295), .Z(z3[421]) );
  NANDN U1937 ( .A(N1030), .B(z2[421]), .Z(n1295) );
  NANDN U1938 ( .A(n3), .B(N1453), .Z(n1294) );
  NAND U1939 ( .A(n1296), .B(n1297), .Z(z3[420]) );
  NANDN U1940 ( .A(N1030), .B(z2[420]), .Z(n1297) );
  NANDN U1941 ( .A(n3), .B(N1452), .Z(n1296) );
  NAND U1942 ( .A(n1298), .B(n1299), .Z(z3[41]) );
  NANDN U1943 ( .A(N1030), .B(z2[41]), .Z(n1299) );
  NANDN U1944 ( .A(n3), .B(N1073), .Z(n1298) );
  NAND U1945 ( .A(n1300), .B(n1301), .Z(z3[419]) );
  NANDN U1946 ( .A(N1030), .B(z2[419]), .Z(n1301) );
  NANDN U1947 ( .A(n3), .B(N1451), .Z(n1300) );
  NAND U1948 ( .A(n1302), .B(n1303), .Z(z3[418]) );
  NANDN U1949 ( .A(N1030), .B(z2[418]), .Z(n1303) );
  NANDN U1950 ( .A(n3), .B(N1450), .Z(n1302) );
  NAND U1951 ( .A(n1304), .B(n1305), .Z(z3[417]) );
  NANDN U1952 ( .A(N1030), .B(z2[417]), .Z(n1305) );
  NANDN U1953 ( .A(n3), .B(N1449), .Z(n1304) );
  NAND U1954 ( .A(n1306), .B(n1307), .Z(z3[416]) );
  NANDN U1955 ( .A(N1030), .B(z2[416]), .Z(n1307) );
  NANDN U1956 ( .A(n3), .B(N1448), .Z(n1306) );
  NAND U1957 ( .A(n1308), .B(n1309), .Z(z3[415]) );
  NANDN U1958 ( .A(N1030), .B(z2[415]), .Z(n1309) );
  NANDN U1959 ( .A(n3), .B(N1447), .Z(n1308) );
  NAND U1960 ( .A(n1310), .B(n1311), .Z(z3[414]) );
  NANDN U1961 ( .A(N1030), .B(z2[414]), .Z(n1311) );
  NANDN U1962 ( .A(n3), .B(N1446), .Z(n1310) );
  NAND U1963 ( .A(n1312), .B(n1313), .Z(z3[413]) );
  NANDN U1964 ( .A(N1030), .B(z2[413]), .Z(n1313) );
  NANDN U1965 ( .A(n3), .B(N1445), .Z(n1312) );
  NAND U1966 ( .A(n1314), .B(n1315), .Z(z3[412]) );
  NANDN U1967 ( .A(N1030), .B(z2[412]), .Z(n1315) );
  NANDN U1968 ( .A(n3), .B(N1444), .Z(n1314) );
  NAND U1969 ( .A(n1316), .B(n1317), .Z(z3[411]) );
  NANDN U1970 ( .A(N1030), .B(z2[411]), .Z(n1317) );
  NANDN U1971 ( .A(n3), .B(N1443), .Z(n1316) );
  NAND U1972 ( .A(n1318), .B(n1319), .Z(z3[410]) );
  NANDN U1973 ( .A(N1030), .B(z2[410]), .Z(n1319) );
  NANDN U1974 ( .A(n3), .B(N1442), .Z(n1318) );
  NAND U1975 ( .A(n1320), .B(n1321), .Z(z3[40]) );
  NANDN U1976 ( .A(N1030), .B(z2[40]), .Z(n1321) );
  NANDN U1977 ( .A(n3), .B(N1072), .Z(n1320) );
  NAND U1978 ( .A(n1322), .B(n1323), .Z(z3[409]) );
  NANDN U1979 ( .A(N1030), .B(z2[409]), .Z(n1323) );
  NANDN U1980 ( .A(n3), .B(N1441), .Z(n1322) );
  NAND U1981 ( .A(n1324), .B(n1325), .Z(z3[408]) );
  NANDN U1982 ( .A(N1030), .B(z2[408]), .Z(n1325) );
  NANDN U1983 ( .A(n3), .B(N1440), .Z(n1324) );
  NAND U1984 ( .A(n1326), .B(n1327), .Z(z3[407]) );
  NANDN U1985 ( .A(N1030), .B(z2[407]), .Z(n1327) );
  NANDN U1986 ( .A(n3), .B(N1439), .Z(n1326) );
  NAND U1987 ( .A(n1328), .B(n1329), .Z(z3[406]) );
  NANDN U1988 ( .A(N1030), .B(z2[406]), .Z(n1329) );
  NANDN U1989 ( .A(n3), .B(N1438), .Z(n1328) );
  NAND U1990 ( .A(n1330), .B(n1331), .Z(z3[405]) );
  NANDN U1991 ( .A(N1030), .B(z2[405]), .Z(n1331) );
  NANDN U1992 ( .A(n3), .B(N1437), .Z(n1330) );
  NAND U1993 ( .A(n1332), .B(n1333), .Z(z3[404]) );
  NANDN U1994 ( .A(N1030), .B(z2[404]), .Z(n1333) );
  NANDN U1995 ( .A(n3), .B(N1436), .Z(n1332) );
  NAND U1996 ( .A(n1334), .B(n1335), .Z(z3[403]) );
  NANDN U1997 ( .A(N1030), .B(z2[403]), .Z(n1335) );
  NANDN U1998 ( .A(n3), .B(N1435), .Z(n1334) );
  NAND U1999 ( .A(n1336), .B(n1337), .Z(z3[402]) );
  NANDN U2000 ( .A(N1030), .B(z2[402]), .Z(n1337) );
  NANDN U2001 ( .A(n3), .B(N1434), .Z(n1336) );
  NAND U2002 ( .A(n1338), .B(n1339), .Z(z3[401]) );
  NANDN U2003 ( .A(N1030), .B(z2[401]), .Z(n1339) );
  NANDN U2004 ( .A(n3), .B(N1433), .Z(n1338) );
  NAND U2005 ( .A(n1340), .B(n1341), .Z(z3[400]) );
  NANDN U2006 ( .A(N1030), .B(z2[400]), .Z(n1341) );
  NANDN U2007 ( .A(n3), .B(N1432), .Z(n1340) );
  NAND U2008 ( .A(n1342), .B(n1343), .Z(z3[3]) );
  NANDN U2009 ( .A(N1030), .B(z2[3]), .Z(n1343) );
  NANDN U2010 ( .A(n3), .B(N1035), .Z(n1342) );
  NAND U2011 ( .A(n1344), .B(n1345), .Z(z3[39]) );
  NANDN U2012 ( .A(N1030), .B(z2[39]), .Z(n1345) );
  NANDN U2013 ( .A(n3), .B(N1071), .Z(n1344) );
  NAND U2014 ( .A(n1346), .B(n1347), .Z(z3[399]) );
  NANDN U2015 ( .A(N1030), .B(z2[399]), .Z(n1347) );
  NANDN U2016 ( .A(n3), .B(N1431), .Z(n1346) );
  NAND U2017 ( .A(n1348), .B(n1349), .Z(z3[398]) );
  NANDN U2018 ( .A(N1030), .B(z2[398]), .Z(n1349) );
  NANDN U2019 ( .A(n3), .B(N1430), .Z(n1348) );
  NAND U2020 ( .A(n1350), .B(n1351), .Z(z3[397]) );
  NANDN U2021 ( .A(N1030), .B(z2[397]), .Z(n1351) );
  NANDN U2022 ( .A(n3), .B(N1429), .Z(n1350) );
  NAND U2023 ( .A(n1352), .B(n1353), .Z(z3[396]) );
  NANDN U2024 ( .A(N1030), .B(z2[396]), .Z(n1353) );
  NANDN U2025 ( .A(n3), .B(N1428), .Z(n1352) );
  NAND U2026 ( .A(n1354), .B(n1355), .Z(z3[395]) );
  NANDN U2027 ( .A(N1030), .B(z2[395]), .Z(n1355) );
  NANDN U2028 ( .A(n3), .B(N1427), .Z(n1354) );
  NAND U2029 ( .A(n1356), .B(n1357), .Z(z3[394]) );
  NANDN U2030 ( .A(N1030), .B(z2[394]), .Z(n1357) );
  NANDN U2031 ( .A(n3), .B(N1426), .Z(n1356) );
  NAND U2032 ( .A(n1358), .B(n1359), .Z(z3[393]) );
  NANDN U2033 ( .A(N1030), .B(z2[393]), .Z(n1359) );
  NANDN U2034 ( .A(n3), .B(N1425), .Z(n1358) );
  NAND U2035 ( .A(n1360), .B(n1361), .Z(z3[392]) );
  NANDN U2036 ( .A(N1030), .B(z2[392]), .Z(n1361) );
  NANDN U2037 ( .A(n3), .B(N1424), .Z(n1360) );
  NAND U2038 ( .A(n1362), .B(n1363), .Z(z3[391]) );
  NANDN U2039 ( .A(N1030), .B(z2[391]), .Z(n1363) );
  NANDN U2040 ( .A(n3), .B(N1423), .Z(n1362) );
  NAND U2041 ( .A(n1364), .B(n1365), .Z(z3[390]) );
  NANDN U2042 ( .A(N1030), .B(z2[390]), .Z(n1365) );
  NANDN U2043 ( .A(n3), .B(N1422), .Z(n1364) );
  NAND U2044 ( .A(n1366), .B(n1367), .Z(z3[38]) );
  NANDN U2045 ( .A(N1030), .B(z2[38]), .Z(n1367) );
  NANDN U2046 ( .A(n3), .B(N1070), .Z(n1366) );
  NAND U2047 ( .A(n1368), .B(n1369), .Z(z3[389]) );
  NANDN U2048 ( .A(N1030), .B(z2[389]), .Z(n1369) );
  NANDN U2049 ( .A(n3), .B(N1421), .Z(n1368) );
  NAND U2050 ( .A(n1370), .B(n1371), .Z(z3[388]) );
  NANDN U2051 ( .A(N1030), .B(z2[388]), .Z(n1371) );
  NANDN U2052 ( .A(n3), .B(N1420), .Z(n1370) );
  NAND U2053 ( .A(n1372), .B(n1373), .Z(z3[387]) );
  NANDN U2054 ( .A(N1030), .B(z2[387]), .Z(n1373) );
  NANDN U2055 ( .A(n3), .B(N1419), .Z(n1372) );
  NAND U2056 ( .A(n1374), .B(n1375), .Z(z3[386]) );
  NANDN U2057 ( .A(N1030), .B(z2[386]), .Z(n1375) );
  NANDN U2058 ( .A(n3), .B(N1418), .Z(n1374) );
  NAND U2059 ( .A(n1376), .B(n1377), .Z(z3[385]) );
  NANDN U2060 ( .A(N1030), .B(z2[385]), .Z(n1377) );
  NANDN U2061 ( .A(n3), .B(N1417), .Z(n1376) );
  NAND U2062 ( .A(n1378), .B(n1379), .Z(z3[384]) );
  NANDN U2063 ( .A(N1030), .B(z2[384]), .Z(n1379) );
  NANDN U2064 ( .A(n3), .B(N1416), .Z(n1378) );
  NAND U2065 ( .A(n1380), .B(n1381), .Z(z3[383]) );
  NANDN U2066 ( .A(N1030), .B(z2[383]), .Z(n1381) );
  NANDN U2067 ( .A(n3), .B(N1415), .Z(n1380) );
  NAND U2068 ( .A(n1382), .B(n1383), .Z(z3[382]) );
  NANDN U2069 ( .A(N1030), .B(z2[382]), .Z(n1383) );
  NANDN U2070 ( .A(n3), .B(N1414), .Z(n1382) );
  NAND U2071 ( .A(n1384), .B(n1385), .Z(z3[381]) );
  NANDN U2072 ( .A(N1030), .B(z2[381]), .Z(n1385) );
  NANDN U2073 ( .A(n3), .B(N1413), .Z(n1384) );
  NAND U2074 ( .A(n1386), .B(n1387), .Z(z3[380]) );
  NANDN U2075 ( .A(N1030), .B(z2[380]), .Z(n1387) );
  NANDN U2076 ( .A(n3), .B(N1412), .Z(n1386) );
  NAND U2077 ( .A(n1388), .B(n1389), .Z(z3[37]) );
  NANDN U2078 ( .A(N1030), .B(z2[37]), .Z(n1389) );
  NANDN U2079 ( .A(n3), .B(N1069), .Z(n1388) );
  NAND U2080 ( .A(n1390), .B(n1391), .Z(z3[379]) );
  NANDN U2081 ( .A(N1030), .B(z2[379]), .Z(n1391) );
  NANDN U2082 ( .A(n3), .B(N1411), .Z(n1390) );
  NAND U2083 ( .A(n1392), .B(n1393), .Z(z3[378]) );
  NANDN U2084 ( .A(N1030), .B(z2[378]), .Z(n1393) );
  NANDN U2085 ( .A(n3), .B(N1410), .Z(n1392) );
  NAND U2086 ( .A(n1394), .B(n1395), .Z(z3[377]) );
  NANDN U2087 ( .A(N1030), .B(z2[377]), .Z(n1395) );
  NANDN U2088 ( .A(n3), .B(N1409), .Z(n1394) );
  NAND U2089 ( .A(n1396), .B(n1397), .Z(z3[376]) );
  NANDN U2090 ( .A(N1030), .B(z2[376]), .Z(n1397) );
  NANDN U2091 ( .A(n3), .B(N1408), .Z(n1396) );
  NAND U2092 ( .A(n1398), .B(n1399), .Z(z3[375]) );
  NANDN U2093 ( .A(N1030), .B(z2[375]), .Z(n1399) );
  NANDN U2094 ( .A(n3), .B(N1407), .Z(n1398) );
  NAND U2095 ( .A(n1400), .B(n1401), .Z(z3[374]) );
  NANDN U2096 ( .A(N1030), .B(z2[374]), .Z(n1401) );
  NANDN U2097 ( .A(n3), .B(N1406), .Z(n1400) );
  NAND U2098 ( .A(n1402), .B(n1403), .Z(z3[373]) );
  NANDN U2099 ( .A(N1030), .B(z2[373]), .Z(n1403) );
  NANDN U2100 ( .A(n3), .B(N1405), .Z(n1402) );
  NAND U2101 ( .A(n1404), .B(n1405), .Z(z3[372]) );
  NANDN U2102 ( .A(N1030), .B(z2[372]), .Z(n1405) );
  NANDN U2103 ( .A(n3), .B(N1404), .Z(n1404) );
  NAND U2104 ( .A(n1406), .B(n1407), .Z(z3[371]) );
  NANDN U2105 ( .A(N1030), .B(z2[371]), .Z(n1407) );
  NANDN U2106 ( .A(n3), .B(N1403), .Z(n1406) );
  NAND U2107 ( .A(n1408), .B(n1409), .Z(z3[370]) );
  NANDN U2108 ( .A(N1030), .B(z2[370]), .Z(n1409) );
  NANDN U2109 ( .A(n3), .B(N1402), .Z(n1408) );
  NAND U2110 ( .A(n1410), .B(n1411), .Z(z3[36]) );
  NANDN U2111 ( .A(N1030), .B(z2[36]), .Z(n1411) );
  NANDN U2112 ( .A(n3), .B(N1068), .Z(n1410) );
  NAND U2113 ( .A(n1412), .B(n1413), .Z(z3[369]) );
  NANDN U2114 ( .A(N1030), .B(z2[369]), .Z(n1413) );
  NANDN U2115 ( .A(n3), .B(N1401), .Z(n1412) );
  NAND U2116 ( .A(n1414), .B(n1415), .Z(z3[368]) );
  NANDN U2117 ( .A(N1030), .B(z2[368]), .Z(n1415) );
  NANDN U2118 ( .A(n3), .B(N1400), .Z(n1414) );
  NAND U2119 ( .A(n1416), .B(n1417), .Z(z3[367]) );
  NANDN U2120 ( .A(N1030), .B(z2[367]), .Z(n1417) );
  NANDN U2121 ( .A(n3), .B(N1399), .Z(n1416) );
  NAND U2122 ( .A(n1418), .B(n1419), .Z(z3[366]) );
  NANDN U2123 ( .A(N1030), .B(z2[366]), .Z(n1419) );
  NANDN U2124 ( .A(n3), .B(N1398), .Z(n1418) );
  NAND U2125 ( .A(n1420), .B(n1421), .Z(z3[365]) );
  NANDN U2126 ( .A(N1030), .B(z2[365]), .Z(n1421) );
  NANDN U2127 ( .A(n3), .B(N1397), .Z(n1420) );
  NAND U2128 ( .A(n1422), .B(n1423), .Z(z3[364]) );
  NANDN U2129 ( .A(N1030), .B(z2[364]), .Z(n1423) );
  NANDN U2130 ( .A(n3), .B(N1396), .Z(n1422) );
  NAND U2131 ( .A(n1424), .B(n1425), .Z(z3[363]) );
  NANDN U2132 ( .A(N1030), .B(z2[363]), .Z(n1425) );
  NANDN U2133 ( .A(n3), .B(N1395), .Z(n1424) );
  NAND U2134 ( .A(n1426), .B(n1427), .Z(z3[362]) );
  NANDN U2135 ( .A(N1030), .B(z2[362]), .Z(n1427) );
  NANDN U2136 ( .A(n3), .B(N1394), .Z(n1426) );
  NAND U2137 ( .A(n1428), .B(n1429), .Z(z3[361]) );
  NANDN U2138 ( .A(N1030), .B(z2[361]), .Z(n1429) );
  NANDN U2139 ( .A(n3), .B(N1393), .Z(n1428) );
  NAND U2140 ( .A(n1430), .B(n1431), .Z(z3[360]) );
  NANDN U2141 ( .A(N1030), .B(z2[360]), .Z(n1431) );
  NANDN U2142 ( .A(n3), .B(N1392), .Z(n1430) );
  NAND U2143 ( .A(n1432), .B(n1433), .Z(z3[35]) );
  NANDN U2144 ( .A(N1030), .B(z2[35]), .Z(n1433) );
  NANDN U2145 ( .A(n3), .B(N1067), .Z(n1432) );
  NAND U2146 ( .A(n1434), .B(n1435), .Z(z3[359]) );
  NANDN U2147 ( .A(N1030), .B(z2[359]), .Z(n1435) );
  NANDN U2148 ( .A(n3), .B(N1391), .Z(n1434) );
  NAND U2149 ( .A(n1436), .B(n1437), .Z(z3[358]) );
  NANDN U2150 ( .A(N1030), .B(z2[358]), .Z(n1437) );
  NANDN U2151 ( .A(n3), .B(N1390), .Z(n1436) );
  NAND U2152 ( .A(n1438), .B(n1439), .Z(z3[357]) );
  NANDN U2153 ( .A(N1030), .B(z2[357]), .Z(n1439) );
  NANDN U2154 ( .A(n3), .B(N1389), .Z(n1438) );
  NAND U2155 ( .A(n1440), .B(n1441), .Z(z3[356]) );
  NANDN U2156 ( .A(N1030), .B(z2[356]), .Z(n1441) );
  NANDN U2157 ( .A(n3), .B(N1388), .Z(n1440) );
  NAND U2158 ( .A(n1442), .B(n1443), .Z(z3[355]) );
  NANDN U2159 ( .A(N1030), .B(z2[355]), .Z(n1443) );
  NANDN U2160 ( .A(n3), .B(N1387), .Z(n1442) );
  NAND U2161 ( .A(n1444), .B(n1445), .Z(z3[354]) );
  NANDN U2162 ( .A(N1030), .B(z2[354]), .Z(n1445) );
  NANDN U2163 ( .A(n3), .B(N1386), .Z(n1444) );
  NAND U2164 ( .A(n1446), .B(n1447), .Z(z3[353]) );
  NANDN U2165 ( .A(N1030), .B(z2[353]), .Z(n1447) );
  NANDN U2166 ( .A(n3), .B(N1385), .Z(n1446) );
  NAND U2167 ( .A(n1448), .B(n1449), .Z(z3[352]) );
  NANDN U2168 ( .A(N1030), .B(z2[352]), .Z(n1449) );
  NANDN U2169 ( .A(n3), .B(N1384), .Z(n1448) );
  NAND U2170 ( .A(n1450), .B(n1451), .Z(z3[351]) );
  NANDN U2171 ( .A(N1030), .B(z2[351]), .Z(n1451) );
  NANDN U2172 ( .A(n3), .B(N1383), .Z(n1450) );
  NAND U2173 ( .A(n1452), .B(n1453), .Z(z3[350]) );
  NANDN U2174 ( .A(N1030), .B(z2[350]), .Z(n1453) );
  NANDN U2175 ( .A(n3), .B(N1382), .Z(n1452) );
  NAND U2176 ( .A(n1454), .B(n1455), .Z(z3[34]) );
  NANDN U2177 ( .A(N1030), .B(z2[34]), .Z(n1455) );
  NANDN U2178 ( .A(n3), .B(N1066), .Z(n1454) );
  NAND U2179 ( .A(n1456), .B(n1457), .Z(z3[349]) );
  NANDN U2180 ( .A(N1030), .B(z2[349]), .Z(n1457) );
  NANDN U2181 ( .A(n3), .B(N1381), .Z(n1456) );
  NAND U2182 ( .A(n1458), .B(n1459), .Z(z3[348]) );
  NANDN U2183 ( .A(N1030), .B(z2[348]), .Z(n1459) );
  NANDN U2184 ( .A(n3), .B(N1380), .Z(n1458) );
  NAND U2185 ( .A(n1460), .B(n1461), .Z(z3[347]) );
  NANDN U2186 ( .A(N1030), .B(z2[347]), .Z(n1461) );
  NANDN U2187 ( .A(n3), .B(N1379), .Z(n1460) );
  NAND U2188 ( .A(n1462), .B(n1463), .Z(z3[346]) );
  NANDN U2189 ( .A(N1030), .B(z2[346]), .Z(n1463) );
  NANDN U2190 ( .A(n3), .B(N1378), .Z(n1462) );
  NAND U2191 ( .A(n1464), .B(n1465), .Z(z3[345]) );
  NANDN U2192 ( .A(N1030), .B(z2[345]), .Z(n1465) );
  NANDN U2193 ( .A(n3), .B(N1377), .Z(n1464) );
  NAND U2194 ( .A(n1466), .B(n1467), .Z(z3[344]) );
  NANDN U2195 ( .A(N1030), .B(z2[344]), .Z(n1467) );
  NANDN U2196 ( .A(n3), .B(N1376), .Z(n1466) );
  NAND U2197 ( .A(n1468), .B(n1469), .Z(z3[343]) );
  NANDN U2198 ( .A(N1030), .B(z2[343]), .Z(n1469) );
  NANDN U2199 ( .A(n3), .B(N1375), .Z(n1468) );
  NAND U2200 ( .A(n1470), .B(n1471), .Z(z3[342]) );
  NANDN U2201 ( .A(N1030), .B(z2[342]), .Z(n1471) );
  NANDN U2202 ( .A(n3), .B(N1374), .Z(n1470) );
  NAND U2203 ( .A(n1472), .B(n1473), .Z(z3[341]) );
  NANDN U2204 ( .A(N1030), .B(z2[341]), .Z(n1473) );
  NANDN U2205 ( .A(n3), .B(N1373), .Z(n1472) );
  NAND U2206 ( .A(n1474), .B(n1475), .Z(z3[340]) );
  NANDN U2207 ( .A(N1030), .B(z2[340]), .Z(n1475) );
  NANDN U2208 ( .A(n3), .B(N1372), .Z(n1474) );
  NAND U2209 ( .A(n1476), .B(n1477), .Z(z3[33]) );
  NANDN U2210 ( .A(N1030), .B(z2[33]), .Z(n1477) );
  NANDN U2211 ( .A(n3), .B(N1065), .Z(n1476) );
  NAND U2212 ( .A(n1478), .B(n1479), .Z(z3[339]) );
  NANDN U2213 ( .A(N1030), .B(z2[339]), .Z(n1479) );
  NANDN U2214 ( .A(n3), .B(N1371), .Z(n1478) );
  NAND U2215 ( .A(n1480), .B(n1481), .Z(z3[338]) );
  NANDN U2216 ( .A(N1030), .B(z2[338]), .Z(n1481) );
  NANDN U2217 ( .A(n3), .B(N1370), .Z(n1480) );
  NAND U2218 ( .A(n1482), .B(n1483), .Z(z3[337]) );
  NANDN U2219 ( .A(N1030), .B(z2[337]), .Z(n1483) );
  NANDN U2220 ( .A(n3), .B(N1369), .Z(n1482) );
  NAND U2221 ( .A(n1484), .B(n1485), .Z(z3[336]) );
  NANDN U2222 ( .A(N1030), .B(z2[336]), .Z(n1485) );
  NANDN U2223 ( .A(n3), .B(N1368), .Z(n1484) );
  NAND U2224 ( .A(n1486), .B(n1487), .Z(z3[335]) );
  NANDN U2225 ( .A(N1030), .B(z2[335]), .Z(n1487) );
  NANDN U2226 ( .A(n3), .B(N1367), .Z(n1486) );
  NAND U2227 ( .A(n1488), .B(n1489), .Z(z3[334]) );
  NANDN U2228 ( .A(N1030), .B(z2[334]), .Z(n1489) );
  NANDN U2229 ( .A(n3), .B(N1366), .Z(n1488) );
  NAND U2230 ( .A(n1490), .B(n1491), .Z(z3[333]) );
  NANDN U2231 ( .A(N1030), .B(z2[333]), .Z(n1491) );
  NANDN U2232 ( .A(n3), .B(N1365), .Z(n1490) );
  NAND U2233 ( .A(n1492), .B(n1493), .Z(z3[332]) );
  NANDN U2234 ( .A(N1030), .B(z2[332]), .Z(n1493) );
  NANDN U2235 ( .A(n3), .B(N1364), .Z(n1492) );
  NAND U2236 ( .A(n1494), .B(n1495), .Z(z3[331]) );
  NANDN U2237 ( .A(N1030), .B(z2[331]), .Z(n1495) );
  NANDN U2238 ( .A(n3), .B(N1363), .Z(n1494) );
  NAND U2239 ( .A(n1496), .B(n1497), .Z(z3[330]) );
  NANDN U2240 ( .A(N1030), .B(z2[330]), .Z(n1497) );
  NANDN U2241 ( .A(n3), .B(N1362), .Z(n1496) );
  NAND U2242 ( .A(n1498), .B(n1499), .Z(z3[32]) );
  NANDN U2243 ( .A(N1030), .B(z2[32]), .Z(n1499) );
  NANDN U2244 ( .A(n3), .B(N1064), .Z(n1498) );
  NAND U2245 ( .A(n1500), .B(n1501), .Z(z3[329]) );
  NANDN U2246 ( .A(N1030), .B(z2[329]), .Z(n1501) );
  NANDN U2247 ( .A(n3), .B(N1361), .Z(n1500) );
  NAND U2248 ( .A(n1502), .B(n1503), .Z(z3[328]) );
  NANDN U2249 ( .A(N1030), .B(z2[328]), .Z(n1503) );
  NANDN U2250 ( .A(n3), .B(N1360), .Z(n1502) );
  NAND U2251 ( .A(n1504), .B(n1505), .Z(z3[327]) );
  NANDN U2252 ( .A(N1030), .B(z2[327]), .Z(n1505) );
  NANDN U2253 ( .A(n3), .B(N1359), .Z(n1504) );
  NAND U2254 ( .A(n1506), .B(n1507), .Z(z3[326]) );
  NANDN U2255 ( .A(N1030), .B(z2[326]), .Z(n1507) );
  NANDN U2256 ( .A(n3), .B(N1358), .Z(n1506) );
  NAND U2257 ( .A(n1508), .B(n1509), .Z(z3[325]) );
  NANDN U2258 ( .A(N1030), .B(z2[325]), .Z(n1509) );
  NANDN U2259 ( .A(n3), .B(N1357), .Z(n1508) );
  NAND U2260 ( .A(n1510), .B(n1511), .Z(z3[324]) );
  NANDN U2261 ( .A(N1030), .B(z2[324]), .Z(n1511) );
  NANDN U2262 ( .A(n3), .B(N1356), .Z(n1510) );
  NAND U2263 ( .A(n1512), .B(n1513), .Z(z3[323]) );
  NANDN U2264 ( .A(N1030), .B(z2[323]), .Z(n1513) );
  NANDN U2265 ( .A(n3), .B(N1355), .Z(n1512) );
  NAND U2266 ( .A(n1514), .B(n1515), .Z(z3[322]) );
  NANDN U2267 ( .A(N1030), .B(z2[322]), .Z(n1515) );
  NANDN U2268 ( .A(n3), .B(N1354), .Z(n1514) );
  NAND U2269 ( .A(n1516), .B(n1517), .Z(z3[321]) );
  NANDN U2270 ( .A(N1030), .B(z2[321]), .Z(n1517) );
  NANDN U2271 ( .A(n3), .B(N1353), .Z(n1516) );
  NAND U2272 ( .A(n1518), .B(n1519), .Z(z3[320]) );
  NANDN U2273 ( .A(N1030), .B(z2[320]), .Z(n1519) );
  NANDN U2274 ( .A(n3), .B(N1352), .Z(n1518) );
  NAND U2275 ( .A(n1520), .B(n1521), .Z(z3[31]) );
  NANDN U2276 ( .A(N1030), .B(z2[31]), .Z(n1521) );
  NANDN U2277 ( .A(n3), .B(N1063), .Z(n1520) );
  NAND U2278 ( .A(n1522), .B(n1523), .Z(z3[319]) );
  NANDN U2279 ( .A(N1030), .B(z2[319]), .Z(n1523) );
  NANDN U2280 ( .A(n3), .B(N1351), .Z(n1522) );
  NAND U2281 ( .A(n1524), .B(n1525), .Z(z3[318]) );
  NANDN U2282 ( .A(N1030), .B(z2[318]), .Z(n1525) );
  NANDN U2283 ( .A(n3), .B(N1350), .Z(n1524) );
  NAND U2284 ( .A(n1526), .B(n1527), .Z(z3[317]) );
  NANDN U2285 ( .A(N1030), .B(z2[317]), .Z(n1527) );
  NANDN U2286 ( .A(n3), .B(N1349), .Z(n1526) );
  NAND U2287 ( .A(n1528), .B(n1529), .Z(z3[316]) );
  NANDN U2288 ( .A(N1030), .B(z2[316]), .Z(n1529) );
  NANDN U2289 ( .A(n3), .B(N1348), .Z(n1528) );
  NAND U2290 ( .A(n1530), .B(n1531), .Z(z3[315]) );
  NANDN U2291 ( .A(N1030), .B(z2[315]), .Z(n1531) );
  NANDN U2292 ( .A(n3), .B(N1347), .Z(n1530) );
  NAND U2293 ( .A(n1532), .B(n1533), .Z(z3[314]) );
  NANDN U2294 ( .A(N1030), .B(z2[314]), .Z(n1533) );
  NANDN U2295 ( .A(n3), .B(N1346), .Z(n1532) );
  NAND U2296 ( .A(n1534), .B(n1535), .Z(z3[313]) );
  NANDN U2297 ( .A(N1030), .B(z2[313]), .Z(n1535) );
  NANDN U2298 ( .A(n3), .B(N1345), .Z(n1534) );
  NAND U2299 ( .A(n1536), .B(n1537), .Z(z3[312]) );
  NANDN U2300 ( .A(N1030), .B(z2[312]), .Z(n1537) );
  NANDN U2301 ( .A(n3), .B(N1344), .Z(n1536) );
  NAND U2302 ( .A(n1538), .B(n1539), .Z(z3[311]) );
  NANDN U2303 ( .A(N1030), .B(z2[311]), .Z(n1539) );
  NANDN U2304 ( .A(n3), .B(N1343), .Z(n1538) );
  NAND U2305 ( .A(n1540), .B(n1541), .Z(z3[310]) );
  NANDN U2306 ( .A(N1030), .B(z2[310]), .Z(n1541) );
  NANDN U2307 ( .A(n3), .B(N1342), .Z(n1540) );
  NAND U2308 ( .A(n1542), .B(n1543), .Z(z3[30]) );
  NANDN U2309 ( .A(N1030), .B(z2[30]), .Z(n1543) );
  NANDN U2310 ( .A(n3), .B(N1062), .Z(n1542) );
  NAND U2311 ( .A(n1544), .B(n1545), .Z(z3[309]) );
  NANDN U2312 ( .A(N1030), .B(z2[309]), .Z(n1545) );
  NANDN U2313 ( .A(n3), .B(N1341), .Z(n1544) );
  NAND U2314 ( .A(n1546), .B(n1547), .Z(z3[308]) );
  NANDN U2315 ( .A(N1030), .B(z2[308]), .Z(n1547) );
  NANDN U2316 ( .A(n3), .B(N1340), .Z(n1546) );
  NAND U2317 ( .A(n1548), .B(n1549), .Z(z3[307]) );
  NANDN U2318 ( .A(N1030), .B(z2[307]), .Z(n1549) );
  NANDN U2319 ( .A(n3), .B(N1339), .Z(n1548) );
  NAND U2320 ( .A(n1550), .B(n1551), .Z(z3[306]) );
  NANDN U2321 ( .A(N1030), .B(z2[306]), .Z(n1551) );
  NANDN U2322 ( .A(n3), .B(N1338), .Z(n1550) );
  NAND U2323 ( .A(n1552), .B(n1553), .Z(z3[305]) );
  NANDN U2324 ( .A(N1030), .B(z2[305]), .Z(n1553) );
  NANDN U2325 ( .A(n3), .B(N1337), .Z(n1552) );
  NAND U2326 ( .A(n1554), .B(n1555), .Z(z3[304]) );
  NANDN U2327 ( .A(N1030), .B(z2[304]), .Z(n1555) );
  NANDN U2328 ( .A(n3), .B(N1336), .Z(n1554) );
  NAND U2329 ( .A(n1556), .B(n1557), .Z(z3[303]) );
  NANDN U2330 ( .A(N1030), .B(z2[303]), .Z(n1557) );
  NANDN U2331 ( .A(n3), .B(N1335), .Z(n1556) );
  NAND U2332 ( .A(n1558), .B(n1559), .Z(z3[302]) );
  NANDN U2333 ( .A(N1030), .B(z2[302]), .Z(n1559) );
  NANDN U2334 ( .A(n3), .B(N1334), .Z(n1558) );
  NAND U2335 ( .A(n1560), .B(n1561), .Z(z3[301]) );
  NANDN U2336 ( .A(N1030), .B(z2[301]), .Z(n1561) );
  NANDN U2337 ( .A(n3), .B(N1333), .Z(n1560) );
  NAND U2338 ( .A(n1562), .B(n1563), .Z(z3[300]) );
  NANDN U2339 ( .A(N1030), .B(z2[300]), .Z(n1563) );
  NANDN U2340 ( .A(n3), .B(N1332), .Z(n1562) );
  NAND U2341 ( .A(n1564), .B(n1565), .Z(z3[2]) );
  NANDN U2342 ( .A(N1030), .B(z2[2]), .Z(n1565) );
  NANDN U2343 ( .A(n3), .B(N1034), .Z(n1564) );
  NAND U2344 ( .A(n1566), .B(n1567), .Z(z3[29]) );
  NANDN U2345 ( .A(N1030), .B(z2[29]), .Z(n1567) );
  NANDN U2346 ( .A(n3), .B(N1061), .Z(n1566) );
  NAND U2347 ( .A(n1568), .B(n1569), .Z(z3[299]) );
  NANDN U2348 ( .A(N1030), .B(z2[299]), .Z(n1569) );
  NANDN U2349 ( .A(n3), .B(N1331), .Z(n1568) );
  NAND U2350 ( .A(n1570), .B(n1571), .Z(z3[298]) );
  NANDN U2351 ( .A(N1030), .B(z2[298]), .Z(n1571) );
  NANDN U2352 ( .A(n3), .B(N1330), .Z(n1570) );
  NAND U2353 ( .A(n1572), .B(n1573), .Z(z3[297]) );
  NANDN U2354 ( .A(N1030), .B(z2[297]), .Z(n1573) );
  NANDN U2355 ( .A(n3), .B(N1329), .Z(n1572) );
  NAND U2356 ( .A(n1574), .B(n1575), .Z(z3[296]) );
  NANDN U2357 ( .A(N1030), .B(z2[296]), .Z(n1575) );
  NANDN U2358 ( .A(n3), .B(N1328), .Z(n1574) );
  NAND U2359 ( .A(n1576), .B(n1577), .Z(z3[295]) );
  NANDN U2360 ( .A(N1030), .B(z2[295]), .Z(n1577) );
  NANDN U2361 ( .A(n3), .B(N1327), .Z(n1576) );
  NAND U2362 ( .A(n1578), .B(n1579), .Z(z3[294]) );
  NANDN U2363 ( .A(N1030), .B(z2[294]), .Z(n1579) );
  NANDN U2364 ( .A(n3), .B(N1326), .Z(n1578) );
  NAND U2365 ( .A(n1580), .B(n1581), .Z(z3[293]) );
  NANDN U2366 ( .A(N1030), .B(z2[293]), .Z(n1581) );
  NANDN U2367 ( .A(n3), .B(N1325), .Z(n1580) );
  NAND U2368 ( .A(n1582), .B(n1583), .Z(z3[292]) );
  NANDN U2369 ( .A(N1030), .B(z2[292]), .Z(n1583) );
  NANDN U2370 ( .A(n3), .B(N1324), .Z(n1582) );
  NAND U2371 ( .A(n1584), .B(n1585), .Z(z3[291]) );
  NANDN U2372 ( .A(N1030), .B(z2[291]), .Z(n1585) );
  NANDN U2373 ( .A(n3), .B(N1323), .Z(n1584) );
  NAND U2374 ( .A(n1586), .B(n1587), .Z(z3[290]) );
  NANDN U2375 ( .A(N1030), .B(z2[290]), .Z(n1587) );
  NANDN U2376 ( .A(n3), .B(N1322), .Z(n1586) );
  NAND U2377 ( .A(n1588), .B(n1589), .Z(z3[28]) );
  NANDN U2378 ( .A(N1030), .B(z2[28]), .Z(n1589) );
  NANDN U2379 ( .A(n3), .B(N1060), .Z(n1588) );
  NAND U2380 ( .A(n1590), .B(n1591), .Z(z3[289]) );
  NANDN U2381 ( .A(N1030), .B(z2[289]), .Z(n1591) );
  NANDN U2382 ( .A(n3), .B(N1321), .Z(n1590) );
  NAND U2383 ( .A(n1592), .B(n1593), .Z(z3[288]) );
  NANDN U2384 ( .A(N1030), .B(z2[288]), .Z(n1593) );
  NANDN U2385 ( .A(n3), .B(N1320), .Z(n1592) );
  NAND U2386 ( .A(n1594), .B(n1595), .Z(z3[287]) );
  NANDN U2387 ( .A(N1030), .B(z2[287]), .Z(n1595) );
  NANDN U2388 ( .A(n3), .B(N1319), .Z(n1594) );
  NAND U2389 ( .A(n1596), .B(n1597), .Z(z3[286]) );
  NANDN U2390 ( .A(N1030), .B(z2[286]), .Z(n1597) );
  NANDN U2391 ( .A(n3), .B(N1318), .Z(n1596) );
  NAND U2392 ( .A(n1598), .B(n1599), .Z(z3[285]) );
  NANDN U2393 ( .A(N1030), .B(z2[285]), .Z(n1599) );
  NANDN U2394 ( .A(n3), .B(N1317), .Z(n1598) );
  NAND U2395 ( .A(n1600), .B(n1601), .Z(z3[284]) );
  NANDN U2396 ( .A(N1030), .B(z2[284]), .Z(n1601) );
  NANDN U2397 ( .A(n3), .B(N1316), .Z(n1600) );
  NAND U2398 ( .A(n1602), .B(n1603), .Z(z3[283]) );
  NANDN U2399 ( .A(N1030), .B(z2[283]), .Z(n1603) );
  NANDN U2400 ( .A(n3), .B(N1315), .Z(n1602) );
  NAND U2401 ( .A(n1604), .B(n1605), .Z(z3[282]) );
  NANDN U2402 ( .A(N1030), .B(z2[282]), .Z(n1605) );
  NANDN U2403 ( .A(n3), .B(N1314), .Z(n1604) );
  NAND U2404 ( .A(n1606), .B(n1607), .Z(z3[281]) );
  NANDN U2405 ( .A(N1030), .B(z2[281]), .Z(n1607) );
  NANDN U2406 ( .A(n3), .B(N1313), .Z(n1606) );
  NAND U2407 ( .A(n1608), .B(n1609), .Z(z3[280]) );
  NANDN U2408 ( .A(N1030), .B(z2[280]), .Z(n1609) );
  NANDN U2409 ( .A(n3), .B(N1312), .Z(n1608) );
  NAND U2410 ( .A(n1610), .B(n1611), .Z(z3[27]) );
  NANDN U2411 ( .A(N1030), .B(z2[27]), .Z(n1611) );
  NANDN U2412 ( .A(n3), .B(N1059), .Z(n1610) );
  NAND U2413 ( .A(n1612), .B(n1613), .Z(z3[279]) );
  NANDN U2414 ( .A(N1030), .B(z2[279]), .Z(n1613) );
  NANDN U2415 ( .A(n3), .B(N1311), .Z(n1612) );
  NAND U2416 ( .A(n1614), .B(n1615), .Z(z3[278]) );
  NANDN U2417 ( .A(N1030), .B(z2[278]), .Z(n1615) );
  NANDN U2418 ( .A(n3), .B(N1310), .Z(n1614) );
  NAND U2419 ( .A(n1616), .B(n1617), .Z(z3[277]) );
  NANDN U2420 ( .A(N1030), .B(z2[277]), .Z(n1617) );
  NANDN U2421 ( .A(n3), .B(N1309), .Z(n1616) );
  NAND U2422 ( .A(n1618), .B(n1619), .Z(z3[276]) );
  NANDN U2423 ( .A(N1030), .B(z2[276]), .Z(n1619) );
  NANDN U2424 ( .A(n3), .B(N1308), .Z(n1618) );
  NAND U2425 ( .A(n1620), .B(n1621), .Z(z3[275]) );
  NANDN U2426 ( .A(N1030), .B(z2[275]), .Z(n1621) );
  NANDN U2427 ( .A(n3), .B(N1307), .Z(n1620) );
  NAND U2428 ( .A(n1622), .B(n1623), .Z(z3[274]) );
  NANDN U2429 ( .A(N1030), .B(z2[274]), .Z(n1623) );
  NANDN U2430 ( .A(n3), .B(N1306), .Z(n1622) );
  NAND U2431 ( .A(n1624), .B(n1625), .Z(z3[273]) );
  NANDN U2432 ( .A(N1030), .B(z2[273]), .Z(n1625) );
  NANDN U2433 ( .A(n3), .B(N1305), .Z(n1624) );
  NAND U2434 ( .A(n1626), .B(n1627), .Z(z3[272]) );
  NANDN U2435 ( .A(N1030), .B(z2[272]), .Z(n1627) );
  NANDN U2436 ( .A(n3), .B(N1304), .Z(n1626) );
  NAND U2437 ( .A(n1628), .B(n1629), .Z(z3[271]) );
  NANDN U2438 ( .A(N1030), .B(z2[271]), .Z(n1629) );
  NANDN U2439 ( .A(n3), .B(N1303), .Z(n1628) );
  NAND U2440 ( .A(n1630), .B(n1631), .Z(z3[270]) );
  NANDN U2441 ( .A(N1030), .B(z2[270]), .Z(n1631) );
  NANDN U2442 ( .A(n3), .B(N1302), .Z(n1630) );
  NAND U2443 ( .A(n1632), .B(n1633), .Z(z3[26]) );
  NANDN U2444 ( .A(N1030), .B(z2[26]), .Z(n1633) );
  NANDN U2445 ( .A(n3), .B(N1058), .Z(n1632) );
  NAND U2446 ( .A(n1634), .B(n1635), .Z(z3[269]) );
  NANDN U2447 ( .A(N1030), .B(z2[269]), .Z(n1635) );
  NANDN U2448 ( .A(n3), .B(N1301), .Z(n1634) );
  NAND U2449 ( .A(n1636), .B(n1637), .Z(z3[268]) );
  NANDN U2450 ( .A(N1030), .B(z2[268]), .Z(n1637) );
  NANDN U2451 ( .A(n3), .B(N1300), .Z(n1636) );
  NAND U2452 ( .A(n1638), .B(n1639), .Z(z3[267]) );
  NANDN U2453 ( .A(N1030), .B(z2[267]), .Z(n1639) );
  NANDN U2454 ( .A(n3), .B(N1299), .Z(n1638) );
  NAND U2455 ( .A(n1640), .B(n1641), .Z(z3[266]) );
  NANDN U2456 ( .A(N1030), .B(z2[266]), .Z(n1641) );
  NANDN U2457 ( .A(n3), .B(N1298), .Z(n1640) );
  NAND U2458 ( .A(n1642), .B(n1643), .Z(z3[265]) );
  NANDN U2459 ( .A(N1030), .B(z2[265]), .Z(n1643) );
  NANDN U2460 ( .A(n3), .B(N1297), .Z(n1642) );
  NAND U2461 ( .A(n1644), .B(n1645), .Z(z3[264]) );
  NANDN U2462 ( .A(N1030), .B(z2[264]), .Z(n1645) );
  NANDN U2463 ( .A(n3), .B(N1296), .Z(n1644) );
  NAND U2464 ( .A(n1646), .B(n1647), .Z(z3[263]) );
  NANDN U2465 ( .A(N1030), .B(z2[263]), .Z(n1647) );
  NANDN U2466 ( .A(n3), .B(N1295), .Z(n1646) );
  NAND U2467 ( .A(n1648), .B(n1649), .Z(z3[262]) );
  NANDN U2468 ( .A(N1030), .B(z2[262]), .Z(n1649) );
  NANDN U2469 ( .A(n3), .B(N1294), .Z(n1648) );
  NAND U2470 ( .A(n1650), .B(n1651), .Z(z3[261]) );
  NANDN U2471 ( .A(N1030), .B(z2[261]), .Z(n1651) );
  NANDN U2472 ( .A(n3), .B(N1293), .Z(n1650) );
  NAND U2473 ( .A(n1652), .B(n1653), .Z(z3[260]) );
  NANDN U2474 ( .A(N1030), .B(z2[260]), .Z(n1653) );
  NANDN U2475 ( .A(n3), .B(N1292), .Z(n1652) );
  NAND U2476 ( .A(n1654), .B(n1655), .Z(z3[25]) );
  NANDN U2477 ( .A(N1030), .B(z2[25]), .Z(n1655) );
  NANDN U2478 ( .A(n3), .B(N1057), .Z(n1654) );
  NAND U2479 ( .A(n1656), .B(n1657), .Z(z3[259]) );
  NANDN U2480 ( .A(N1030), .B(z2[259]), .Z(n1657) );
  NANDN U2481 ( .A(n3), .B(N1291), .Z(n1656) );
  NAND U2482 ( .A(n1658), .B(n1659), .Z(z3[258]) );
  NANDN U2483 ( .A(N1030), .B(z2[258]), .Z(n1659) );
  NANDN U2484 ( .A(n3), .B(N1290), .Z(n1658) );
  NAND U2485 ( .A(n1660), .B(n1661), .Z(z3[257]) );
  NANDN U2486 ( .A(N1030), .B(z2[257]), .Z(n1661) );
  NANDN U2487 ( .A(n3), .B(N1289), .Z(n1660) );
  NAND U2488 ( .A(n1662), .B(n1663), .Z(z3[256]) );
  NANDN U2489 ( .A(N1030), .B(z2[256]), .Z(n1663) );
  NANDN U2490 ( .A(n3), .B(N1288), .Z(n1662) );
  NAND U2491 ( .A(n1664), .B(n1665), .Z(z3[255]) );
  NANDN U2492 ( .A(N1030), .B(z2[255]), .Z(n1665) );
  NANDN U2493 ( .A(n3), .B(N1287), .Z(n1664) );
  NAND U2494 ( .A(n1666), .B(n1667), .Z(z3[254]) );
  NANDN U2495 ( .A(N1030), .B(z2[254]), .Z(n1667) );
  NANDN U2496 ( .A(n3), .B(N1286), .Z(n1666) );
  NAND U2497 ( .A(n1668), .B(n1669), .Z(z3[253]) );
  NANDN U2498 ( .A(N1030), .B(z2[253]), .Z(n1669) );
  NANDN U2499 ( .A(n3), .B(N1285), .Z(n1668) );
  NAND U2500 ( .A(n1670), .B(n1671), .Z(z3[252]) );
  NANDN U2501 ( .A(N1030), .B(z2[252]), .Z(n1671) );
  NANDN U2502 ( .A(n3), .B(N1284), .Z(n1670) );
  NAND U2503 ( .A(n1672), .B(n1673), .Z(z3[251]) );
  NANDN U2504 ( .A(N1030), .B(z2[251]), .Z(n1673) );
  NANDN U2505 ( .A(n3), .B(N1283), .Z(n1672) );
  NAND U2506 ( .A(n1674), .B(n1675), .Z(z3[250]) );
  NANDN U2507 ( .A(N1030), .B(z2[250]), .Z(n1675) );
  NANDN U2508 ( .A(n3), .B(N1282), .Z(n1674) );
  NAND U2509 ( .A(n1676), .B(n1677), .Z(z3[24]) );
  NANDN U2510 ( .A(N1030), .B(z2[24]), .Z(n1677) );
  NANDN U2511 ( .A(n3), .B(N1056), .Z(n1676) );
  NAND U2512 ( .A(n1678), .B(n1679), .Z(z3[249]) );
  NANDN U2513 ( .A(N1030), .B(z2[249]), .Z(n1679) );
  NANDN U2514 ( .A(n3), .B(N1281), .Z(n1678) );
  NAND U2515 ( .A(n1680), .B(n1681), .Z(z3[248]) );
  NANDN U2516 ( .A(N1030), .B(z2[248]), .Z(n1681) );
  NANDN U2517 ( .A(n3), .B(N1280), .Z(n1680) );
  NAND U2518 ( .A(n1682), .B(n1683), .Z(z3[247]) );
  NANDN U2519 ( .A(N1030), .B(z2[247]), .Z(n1683) );
  NANDN U2520 ( .A(n3), .B(N1279), .Z(n1682) );
  NAND U2521 ( .A(n1684), .B(n1685), .Z(z3[246]) );
  NANDN U2522 ( .A(N1030), .B(z2[246]), .Z(n1685) );
  NANDN U2523 ( .A(n3), .B(N1278), .Z(n1684) );
  NAND U2524 ( .A(n1686), .B(n1687), .Z(z3[245]) );
  NANDN U2525 ( .A(N1030), .B(z2[245]), .Z(n1687) );
  NANDN U2526 ( .A(n3), .B(N1277), .Z(n1686) );
  NAND U2527 ( .A(n1688), .B(n1689), .Z(z3[244]) );
  NANDN U2528 ( .A(N1030), .B(z2[244]), .Z(n1689) );
  NANDN U2529 ( .A(n3), .B(N1276), .Z(n1688) );
  NAND U2530 ( .A(n1690), .B(n1691), .Z(z3[243]) );
  NANDN U2531 ( .A(N1030), .B(z2[243]), .Z(n1691) );
  NANDN U2532 ( .A(n3), .B(N1275), .Z(n1690) );
  NAND U2533 ( .A(n1692), .B(n1693), .Z(z3[242]) );
  NANDN U2534 ( .A(N1030), .B(z2[242]), .Z(n1693) );
  NANDN U2535 ( .A(n3), .B(N1274), .Z(n1692) );
  NAND U2536 ( .A(n1694), .B(n1695), .Z(z3[241]) );
  NANDN U2537 ( .A(N1030), .B(z2[241]), .Z(n1695) );
  NANDN U2538 ( .A(n3), .B(N1273), .Z(n1694) );
  NAND U2539 ( .A(n1696), .B(n1697), .Z(z3[240]) );
  NANDN U2540 ( .A(N1030), .B(z2[240]), .Z(n1697) );
  NANDN U2541 ( .A(n3), .B(N1272), .Z(n1696) );
  NAND U2542 ( .A(n1698), .B(n1699), .Z(z3[23]) );
  NANDN U2543 ( .A(N1030), .B(z2[23]), .Z(n1699) );
  NANDN U2544 ( .A(n3), .B(N1055), .Z(n1698) );
  NAND U2545 ( .A(n1700), .B(n1701), .Z(z3[239]) );
  NANDN U2546 ( .A(N1030), .B(z2[239]), .Z(n1701) );
  NANDN U2547 ( .A(n3), .B(N1271), .Z(n1700) );
  NAND U2548 ( .A(n1702), .B(n1703), .Z(z3[238]) );
  NANDN U2549 ( .A(N1030), .B(z2[238]), .Z(n1703) );
  NANDN U2550 ( .A(n3), .B(N1270), .Z(n1702) );
  NAND U2551 ( .A(n1704), .B(n1705), .Z(z3[237]) );
  NANDN U2552 ( .A(N1030), .B(z2[237]), .Z(n1705) );
  NANDN U2553 ( .A(n3), .B(N1269), .Z(n1704) );
  NAND U2554 ( .A(n1706), .B(n1707), .Z(z3[236]) );
  NANDN U2555 ( .A(N1030), .B(z2[236]), .Z(n1707) );
  NANDN U2556 ( .A(n3), .B(N1268), .Z(n1706) );
  NAND U2557 ( .A(n1708), .B(n1709), .Z(z3[235]) );
  NANDN U2558 ( .A(N1030), .B(z2[235]), .Z(n1709) );
  NANDN U2559 ( .A(n3), .B(N1267), .Z(n1708) );
  NAND U2560 ( .A(n1710), .B(n1711), .Z(z3[234]) );
  NANDN U2561 ( .A(N1030), .B(z2[234]), .Z(n1711) );
  NANDN U2562 ( .A(n3), .B(N1266), .Z(n1710) );
  NAND U2563 ( .A(n1712), .B(n1713), .Z(z3[233]) );
  NANDN U2564 ( .A(N1030), .B(z2[233]), .Z(n1713) );
  NANDN U2565 ( .A(n3), .B(N1265), .Z(n1712) );
  NAND U2566 ( .A(n1714), .B(n1715), .Z(z3[232]) );
  NANDN U2567 ( .A(N1030), .B(z2[232]), .Z(n1715) );
  NANDN U2568 ( .A(n3), .B(N1264), .Z(n1714) );
  NAND U2569 ( .A(n1716), .B(n1717), .Z(z3[231]) );
  NANDN U2570 ( .A(N1030), .B(z2[231]), .Z(n1717) );
  NANDN U2571 ( .A(n3), .B(N1263), .Z(n1716) );
  NAND U2572 ( .A(n1718), .B(n1719), .Z(z3[230]) );
  NANDN U2573 ( .A(N1030), .B(z2[230]), .Z(n1719) );
  NANDN U2574 ( .A(n3), .B(N1262), .Z(n1718) );
  NAND U2575 ( .A(n1720), .B(n1721), .Z(z3[22]) );
  NANDN U2576 ( .A(N1030), .B(z2[22]), .Z(n1721) );
  NANDN U2577 ( .A(n3), .B(N1054), .Z(n1720) );
  NAND U2578 ( .A(n1722), .B(n1723), .Z(z3[229]) );
  NANDN U2579 ( .A(N1030), .B(z2[229]), .Z(n1723) );
  NANDN U2580 ( .A(n3), .B(N1261), .Z(n1722) );
  NAND U2581 ( .A(n1724), .B(n1725), .Z(z3[228]) );
  NANDN U2582 ( .A(N1030), .B(z2[228]), .Z(n1725) );
  NANDN U2583 ( .A(n3), .B(N1260), .Z(n1724) );
  NAND U2584 ( .A(n1726), .B(n1727), .Z(z3[227]) );
  NANDN U2585 ( .A(N1030), .B(z2[227]), .Z(n1727) );
  NANDN U2586 ( .A(n3), .B(N1259), .Z(n1726) );
  NAND U2587 ( .A(n1728), .B(n1729), .Z(z3[226]) );
  NANDN U2588 ( .A(N1030), .B(z2[226]), .Z(n1729) );
  NANDN U2589 ( .A(n3), .B(N1258), .Z(n1728) );
  NAND U2590 ( .A(n1730), .B(n1731), .Z(z3[225]) );
  NANDN U2591 ( .A(N1030), .B(z2[225]), .Z(n1731) );
  NANDN U2592 ( .A(n3), .B(N1257), .Z(n1730) );
  NAND U2593 ( .A(n1732), .B(n1733), .Z(z3[224]) );
  NANDN U2594 ( .A(N1030), .B(z2[224]), .Z(n1733) );
  NANDN U2595 ( .A(n3), .B(N1256), .Z(n1732) );
  NAND U2596 ( .A(n1734), .B(n1735), .Z(z3[223]) );
  NANDN U2597 ( .A(N1030), .B(z2[223]), .Z(n1735) );
  NANDN U2598 ( .A(n3), .B(N1255), .Z(n1734) );
  NAND U2599 ( .A(n1736), .B(n1737), .Z(z3[222]) );
  NANDN U2600 ( .A(N1030), .B(z2[222]), .Z(n1737) );
  NANDN U2601 ( .A(n3), .B(N1254), .Z(n1736) );
  NAND U2602 ( .A(n1738), .B(n1739), .Z(z3[221]) );
  NANDN U2603 ( .A(N1030), .B(z2[221]), .Z(n1739) );
  NANDN U2604 ( .A(n3), .B(N1253), .Z(n1738) );
  NAND U2605 ( .A(n1740), .B(n1741), .Z(z3[220]) );
  NANDN U2606 ( .A(N1030), .B(z2[220]), .Z(n1741) );
  NANDN U2607 ( .A(n3), .B(N1252), .Z(n1740) );
  NAND U2608 ( .A(n1742), .B(n1743), .Z(z3[21]) );
  NANDN U2609 ( .A(N1030), .B(z2[21]), .Z(n1743) );
  NANDN U2610 ( .A(n3), .B(N1053), .Z(n1742) );
  NAND U2611 ( .A(n1744), .B(n1745), .Z(z3[219]) );
  NANDN U2612 ( .A(N1030), .B(z2[219]), .Z(n1745) );
  NANDN U2613 ( .A(n3), .B(N1251), .Z(n1744) );
  NAND U2614 ( .A(n1746), .B(n1747), .Z(z3[218]) );
  NANDN U2615 ( .A(N1030), .B(z2[218]), .Z(n1747) );
  NANDN U2616 ( .A(n3), .B(N1250), .Z(n1746) );
  NAND U2617 ( .A(n1748), .B(n1749), .Z(z3[217]) );
  NANDN U2618 ( .A(N1030), .B(z2[217]), .Z(n1749) );
  NANDN U2619 ( .A(n3), .B(N1249), .Z(n1748) );
  NAND U2620 ( .A(n1750), .B(n1751), .Z(z3[216]) );
  NANDN U2621 ( .A(N1030), .B(z2[216]), .Z(n1751) );
  NANDN U2622 ( .A(n3), .B(N1248), .Z(n1750) );
  NAND U2623 ( .A(n1752), .B(n1753), .Z(z3[215]) );
  NANDN U2624 ( .A(N1030), .B(z2[215]), .Z(n1753) );
  NANDN U2625 ( .A(n3), .B(N1247), .Z(n1752) );
  NAND U2626 ( .A(n1754), .B(n1755), .Z(z3[214]) );
  NANDN U2627 ( .A(N1030), .B(z2[214]), .Z(n1755) );
  NANDN U2628 ( .A(n3), .B(N1246), .Z(n1754) );
  NAND U2629 ( .A(n1756), .B(n1757), .Z(z3[213]) );
  NANDN U2630 ( .A(N1030), .B(z2[213]), .Z(n1757) );
  NANDN U2631 ( .A(n3), .B(N1245), .Z(n1756) );
  NAND U2632 ( .A(n1758), .B(n1759), .Z(z3[212]) );
  NANDN U2633 ( .A(N1030), .B(z2[212]), .Z(n1759) );
  NANDN U2634 ( .A(n3), .B(N1244), .Z(n1758) );
  NAND U2635 ( .A(n1760), .B(n1761), .Z(z3[211]) );
  NANDN U2636 ( .A(N1030), .B(z2[211]), .Z(n1761) );
  NANDN U2637 ( .A(n3), .B(N1243), .Z(n1760) );
  NAND U2638 ( .A(n1762), .B(n1763), .Z(z3[210]) );
  NANDN U2639 ( .A(N1030), .B(z2[210]), .Z(n1763) );
  NANDN U2640 ( .A(n3), .B(N1242), .Z(n1762) );
  NAND U2641 ( .A(n1764), .B(n1765), .Z(z3[20]) );
  NANDN U2642 ( .A(N1030), .B(z2[20]), .Z(n1765) );
  NANDN U2643 ( .A(n3), .B(N1052), .Z(n1764) );
  NAND U2644 ( .A(n1766), .B(n1767), .Z(z3[209]) );
  NANDN U2645 ( .A(N1030), .B(z2[209]), .Z(n1767) );
  NANDN U2646 ( .A(n3), .B(N1241), .Z(n1766) );
  NAND U2647 ( .A(n1768), .B(n1769), .Z(z3[208]) );
  NANDN U2648 ( .A(N1030), .B(z2[208]), .Z(n1769) );
  NANDN U2649 ( .A(n3), .B(N1240), .Z(n1768) );
  NAND U2650 ( .A(n1770), .B(n1771), .Z(z3[207]) );
  NANDN U2651 ( .A(N1030), .B(z2[207]), .Z(n1771) );
  NANDN U2652 ( .A(n3), .B(N1239), .Z(n1770) );
  NAND U2653 ( .A(n1772), .B(n1773), .Z(z3[206]) );
  NANDN U2654 ( .A(N1030), .B(z2[206]), .Z(n1773) );
  NANDN U2655 ( .A(n3), .B(N1238), .Z(n1772) );
  NAND U2656 ( .A(n1774), .B(n1775), .Z(z3[205]) );
  NANDN U2657 ( .A(N1030), .B(z2[205]), .Z(n1775) );
  NANDN U2658 ( .A(n3), .B(N1237), .Z(n1774) );
  NAND U2659 ( .A(n1776), .B(n1777), .Z(z3[204]) );
  NANDN U2660 ( .A(N1030), .B(z2[204]), .Z(n1777) );
  NANDN U2661 ( .A(n3), .B(N1236), .Z(n1776) );
  NAND U2662 ( .A(n1778), .B(n1779), .Z(z3[203]) );
  NANDN U2663 ( .A(N1030), .B(z2[203]), .Z(n1779) );
  NANDN U2664 ( .A(n3), .B(N1235), .Z(n1778) );
  NAND U2665 ( .A(n1780), .B(n1781), .Z(z3[202]) );
  NANDN U2666 ( .A(N1030), .B(z2[202]), .Z(n1781) );
  NANDN U2667 ( .A(n3), .B(N1234), .Z(n1780) );
  NAND U2668 ( .A(n1782), .B(n1783), .Z(z3[201]) );
  NANDN U2669 ( .A(N1030), .B(z2[201]), .Z(n1783) );
  NANDN U2670 ( .A(n3), .B(N1233), .Z(n1782) );
  NAND U2671 ( .A(n1784), .B(n1785), .Z(z3[200]) );
  NANDN U2672 ( .A(N1030), .B(z2[200]), .Z(n1785) );
  NANDN U2673 ( .A(n3), .B(N1232), .Z(n1784) );
  NAND U2674 ( .A(n1786), .B(n1787), .Z(z3[1]) );
  NANDN U2675 ( .A(N1030), .B(z2[1]), .Z(n1787) );
  NANDN U2676 ( .A(n3), .B(N1033), .Z(n1786) );
  NAND U2677 ( .A(n1788), .B(n1789), .Z(z3[19]) );
  NANDN U2678 ( .A(N1030), .B(z2[19]), .Z(n1789) );
  NANDN U2679 ( .A(n3), .B(N1051), .Z(n1788) );
  NAND U2680 ( .A(n1790), .B(n1791), .Z(z3[199]) );
  NANDN U2681 ( .A(N1030), .B(z2[199]), .Z(n1791) );
  NANDN U2682 ( .A(n3), .B(N1231), .Z(n1790) );
  NAND U2683 ( .A(n1792), .B(n1793), .Z(z3[198]) );
  NANDN U2684 ( .A(N1030), .B(z2[198]), .Z(n1793) );
  NANDN U2685 ( .A(n3), .B(N1230), .Z(n1792) );
  NAND U2686 ( .A(n1794), .B(n1795), .Z(z3[197]) );
  NANDN U2687 ( .A(N1030), .B(z2[197]), .Z(n1795) );
  NANDN U2688 ( .A(n3), .B(N1229), .Z(n1794) );
  NAND U2689 ( .A(n1796), .B(n1797), .Z(z3[196]) );
  NANDN U2690 ( .A(N1030), .B(z2[196]), .Z(n1797) );
  NANDN U2691 ( .A(n3), .B(N1228), .Z(n1796) );
  NAND U2692 ( .A(n1798), .B(n1799), .Z(z3[195]) );
  NANDN U2693 ( .A(N1030), .B(z2[195]), .Z(n1799) );
  NANDN U2694 ( .A(n3), .B(N1227), .Z(n1798) );
  NAND U2695 ( .A(n1800), .B(n1801), .Z(z3[194]) );
  NANDN U2696 ( .A(N1030), .B(z2[194]), .Z(n1801) );
  NANDN U2697 ( .A(n3), .B(N1226), .Z(n1800) );
  NAND U2698 ( .A(n1802), .B(n1803), .Z(z3[193]) );
  NANDN U2699 ( .A(N1030), .B(z2[193]), .Z(n1803) );
  NANDN U2700 ( .A(n3), .B(N1225), .Z(n1802) );
  NAND U2701 ( .A(n1804), .B(n1805), .Z(z3[192]) );
  NANDN U2702 ( .A(N1030), .B(z2[192]), .Z(n1805) );
  NANDN U2703 ( .A(n3), .B(N1224), .Z(n1804) );
  NAND U2704 ( .A(n1806), .B(n1807), .Z(z3[191]) );
  NANDN U2705 ( .A(N1030), .B(z2[191]), .Z(n1807) );
  NANDN U2706 ( .A(n3), .B(N1223), .Z(n1806) );
  NAND U2707 ( .A(n1808), .B(n1809), .Z(z3[190]) );
  NANDN U2708 ( .A(N1030), .B(z2[190]), .Z(n1809) );
  NANDN U2709 ( .A(n3), .B(N1222), .Z(n1808) );
  NAND U2710 ( .A(n1810), .B(n1811), .Z(z3[18]) );
  NANDN U2711 ( .A(N1030), .B(z2[18]), .Z(n1811) );
  NANDN U2712 ( .A(n3), .B(N1050), .Z(n1810) );
  NAND U2713 ( .A(n1812), .B(n1813), .Z(z3[189]) );
  NANDN U2714 ( .A(N1030), .B(z2[189]), .Z(n1813) );
  NANDN U2715 ( .A(n3), .B(N1221), .Z(n1812) );
  NAND U2716 ( .A(n1814), .B(n1815), .Z(z3[188]) );
  NANDN U2717 ( .A(N1030), .B(z2[188]), .Z(n1815) );
  NANDN U2718 ( .A(n3), .B(N1220), .Z(n1814) );
  NAND U2719 ( .A(n1816), .B(n1817), .Z(z3[187]) );
  NANDN U2720 ( .A(N1030), .B(z2[187]), .Z(n1817) );
  NANDN U2721 ( .A(n3), .B(N1219), .Z(n1816) );
  NAND U2722 ( .A(n1818), .B(n1819), .Z(z3[186]) );
  NANDN U2723 ( .A(N1030), .B(z2[186]), .Z(n1819) );
  NANDN U2724 ( .A(n3), .B(N1218), .Z(n1818) );
  NAND U2725 ( .A(n1820), .B(n1821), .Z(z3[185]) );
  NANDN U2726 ( .A(N1030), .B(z2[185]), .Z(n1821) );
  NANDN U2727 ( .A(n3), .B(N1217), .Z(n1820) );
  NAND U2728 ( .A(n1822), .B(n1823), .Z(z3[184]) );
  NANDN U2729 ( .A(N1030), .B(z2[184]), .Z(n1823) );
  NANDN U2730 ( .A(n3), .B(N1216), .Z(n1822) );
  NAND U2731 ( .A(n1824), .B(n1825), .Z(z3[183]) );
  NANDN U2732 ( .A(N1030), .B(z2[183]), .Z(n1825) );
  NANDN U2733 ( .A(n3), .B(N1215), .Z(n1824) );
  NAND U2734 ( .A(n1826), .B(n1827), .Z(z3[182]) );
  NANDN U2735 ( .A(N1030), .B(z2[182]), .Z(n1827) );
  NANDN U2736 ( .A(n3), .B(N1214), .Z(n1826) );
  NAND U2737 ( .A(n1828), .B(n1829), .Z(z3[181]) );
  NANDN U2738 ( .A(N1030), .B(z2[181]), .Z(n1829) );
  NANDN U2739 ( .A(n3), .B(N1213), .Z(n1828) );
  NAND U2740 ( .A(n1830), .B(n1831), .Z(z3[180]) );
  NANDN U2741 ( .A(N1030), .B(z2[180]), .Z(n1831) );
  NANDN U2742 ( .A(n3), .B(N1212), .Z(n1830) );
  NAND U2743 ( .A(n1832), .B(n1833), .Z(z3[17]) );
  NANDN U2744 ( .A(N1030), .B(z2[17]), .Z(n1833) );
  NANDN U2745 ( .A(n3), .B(N1049), .Z(n1832) );
  NAND U2746 ( .A(n1834), .B(n1835), .Z(z3[179]) );
  NANDN U2747 ( .A(N1030), .B(z2[179]), .Z(n1835) );
  NANDN U2748 ( .A(n3), .B(N1211), .Z(n1834) );
  NAND U2749 ( .A(n1836), .B(n1837), .Z(z3[178]) );
  NANDN U2750 ( .A(N1030), .B(z2[178]), .Z(n1837) );
  NANDN U2751 ( .A(n3), .B(N1210), .Z(n1836) );
  NAND U2752 ( .A(n1838), .B(n1839), .Z(z3[177]) );
  NANDN U2753 ( .A(N1030), .B(z2[177]), .Z(n1839) );
  NANDN U2754 ( .A(n3), .B(N1209), .Z(n1838) );
  NAND U2755 ( .A(n1840), .B(n1841), .Z(z3[176]) );
  NANDN U2756 ( .A(N1030), .B(z2[176]), .Z(n1841) );
  NANDN U2757 ( .A(n3), .B(N1208), .Z(n1840) );
  NAND U2758 ( .A(n1842), .B(n1843), .Z(z3[175]) );
  NANDN U2759 ( .A(N1030), .B(z2[175]), .Z(n1843) );
  NANDN U2760 ( .A(n3), .B(N1207), .Z(n1842) );
  NAND U2761 ( .A(n1844), .B(n1845), .Z(z3[174]) );
  NANDN U2762 ( .A(N1030), .B(z2[174]), .Z(n1845) );
  NANDN U2763 ( .A(n3), .B(N1206), .Z(n1844) );
  NAND U2764 ( .A(n1846), .B(n1847), .Z(z3[173]) );
  NANDN U2765 ( .A(N1030), .B(z2[173]), .Z(n1847) );
  NANDN U2766 ( .A(n3), .B(N1205), .Z(n1846) );
  NAND U2767 ( .A(n1848), .B(n1849), .Z(z3[172]) );
  NANDN U2768 ( .A(N1030), .B(z2[172]), .Z(n1849) );
  NANDN U2769 ( .A(n3), .B(N1204), .Z(n1848) );
  NAND U2770 ( .A(n1850), .B(n1851), .Z(z3[171]) );
  NANDN U2771 ( .A(N1030), .B(z2[171]), .Z(n1851) );
  NANDN U2772 ( .A(n3), .B(N1203), .Z(n1850) );
  NAND U2773 ( .A(n1852), .B(n1853), .Z(z3[170]) );
  NANDN U2774 ( .A(N1030), .B(z2[170]), .Z(n1853) );
  NANDN U2775 ( .A(n3), .B(N1202), .Z(n1852) );
  NAND U2776 ( .A(n1854), .B(n1855), .Z(z3[16]) );
  NANDN U2777 ( .A(N1030), .B(z2[16]), .Z(n1855) );
  NANDN U2778 ( .A(n3), .B(N1048), .Z(n1854) );
  NAND U2779 ( .A(n1856), .B(n1857), .Z(z3[169]) );
  NANDN U2780 ( .A(N1030), .B(z2[169]), .Z(n1857) );
  NANDN U2781 ( .A(n3), .B(N1201), .Z(n1856) );
  NAND U2782 ( .A(n1858), .B(n1859), .Z(z3[168]) );
  NANDN U2783 ( .A(N1030), .B(z2[168]), .Z(n1859) );
  NANDN U2784 ( .A(n3), .B(N1200), .Z(n1858) );
  NAND U2785 ( .A(n1860), .B(n1861), .Z(z3[167]) );
  NANDN U2786 ( .A(N1030), .B(z2[167]), .Z(n1861) );
  NANDN U2787 ( .A(n3), .B(N1199), .Z(n1860) );
  NAND U2788 ( .A(n1862), .B(n1863), .Z(z3[166]) );
  NANDN U2789 ( .A(N1030), .B(z2[166]), .Z(n1863) );
  NANDN U2790 ( .A(n3), .B(N1198), .Z(n1862) );
  NAND U2791 ( .A(n1864), .B(n1865), .Z(z3[165]) );
  NANDN U2792 ( .A(N1030), .B(z2[165]), .Z(n1865) );
  NANDN U2793 ( .A(n3), .B(N1197), .Z(n1864) );
  NAND U2794 ( .A(n1866), .B(n1867), .Z(z3[164]) );
  NANDN U2795 ( .A(N1030), .B(z2[164]), .Z(n1867) );
  NANDN U2796 ( .A(n3), .B(N1196), .Z(n1866) );
  NAND U2797 ( .A(n1868), .B(n1869), .Z(z3[163]) );
  NANDN U2798 ( .A(N1030), .B(z2[163]), .Z(n1869) );
  NANDN U2799 ( .A(n3), .B(N1195), .Z(n1868) );
  NAND U2800 ( .A(n1870), .B(n1871), .Z(z3[162]) );
  NANDN U2801 ( .A(N1030), .B(z2[162]), .Z(n1871) );
  NANDN U2802 ( .A(n3), .B(N1194), .Z(n1870) );
  NAND U2803 ( .A(n1872), .B(n1873), .Z(z3[161]) );
  NANDN U2804 ( .A(N1030), .B(z2[161]), .Z(n1873) );
  NANDN U2805 ( .A(n3), .B(N1193), .Z(n1872) );
  NAND U2806 ( .A(n1874), .B(n1875), .Z(z3[160]) );
  NANDN U2807 ( .A(N1030), .B(z2[160]), .Z(n1875) );
  NANDN U2808 ( .A(n3), .B(N1192), .Z(n1874) );
  NAND U2809 ( .A(n1876), .B(n1877), .Z(z3[15]) );
  NANDN U2810 ( .A(N1030), .B(z2[15]), .Z(n1877) );
  NANDN U2811 ( .A(n3), .B(N1047), .Z(n1876) );
  NAND U2812 ( .A(n1878), .B(n1879), .Z(z3[159]) );
  NANDN U2813 ( .A(N1030), .B(z2[159]), .Z(n1879) );
  NANDN U2814 ( .A(n3), .B(N1191), .Z(n1878) );
  NAND U2815 ( .A(n1880), .B(n1881), .Z(z3[158]) );
  NANDN U2816 ( .A(N1030), .B(z2[158]), .Z(n1881) );
  NANDN U2817 ( .A(n3), .B(N1190), .Z(n1880) );
  NAND U2818 ( .A(n1882), .B(n1883), .Z(z3[157]) );
  NANDN U2819 ( .A(N1030), .B(z2[157]), .Z(n1883) );
  NANDN U2820 ( .A(n3), .B(N1189), .Z(n1882) );
  NAND U2821 ( .A(n1884), .B(n1885), .Z(z3[156]) );
  NANDN U2822 ( .A(N1030), .B(z2[156]), .Z(n1885) );
  NANDN U2823 ( .A(n3), .B(N1188), .Z(n1884) );
  NAND U2824 ( .A(n1886), .B(n1887), .Z(z3[155]) );
  NANDN U2825 ( .A(N1030), .B(z2[155]), .Z(n1887) );
  NANDN U2826 ( .A(n3), .B(N1187), .Z(n1886) );
  NAND U2827 ( .A(n1888), .B(n1889), .Z(z3[154]) );
  NANDN U2828 ( .A(N1030), .B(z2[154]), .Z(n1889) );
  NANDN U2829 ( .A(n3), .B(N1186), .Z(n1888) );
  NAND U2830 ( .A(n1890), .B(n1891), .Z(z3[153]) );
  NANDN U2831 ( .A(N1030), .B(z2[153]), .Z(n1891) );
  NANDN U2832 ( .A(n3), .B(N1185), .Z(n1890) );
  NAND U2833 ( .A(n1892), .B(n1893), .Z(z3[152]) );
  NANDN U2834 ( .A(N1030), .B(z2[152]), .Z(n1893) );
  NANDN U2835 ( .A(n3), .B(N1184), .Z(n1892) );
  NAND U2836 ( .A(n1894), .B(n1895), .Z(z3[151]) );
  NANDN U2837 ( .A(N1030), .B(z2[151]), .Z(n1895) );
  NANDN U2838 ( .A(n3), .B(N1183), .Z(n1894) );
  NAND U2839 ( .A(n1896), .B(n1897), .Z(z3[150]) );
  NANDN U2840 ( .A(N1030), .B(z2[150]), .Z(n1897) );
  NANDN U2841 ( .A(n3), .B(N1182), .Z(n1896) );
  NAND U2842 ( .A(n1898), .B(n1899), .Z(z3[14]) );
  NANDN U2843 ( .A(N1030), .B(z2[14]), .Z(n1899) );
  NANDN U2844 ( .A(n3), .B(N1046), .Z(n1898) );
  NAND U2845 ( .A(n1900), .B(n1901), .Z(z3[149]) );
  NANDN U2846 ( .A(N1030), .B(z2[149]), .Z(n1901) );
  NANDN U2847 ( .A(n3), .B(N1181), .Z(n1900) );
  NAND U2848 ( .A(n1902), .B(n1903), .Z(z3[148]) );
  NANDN U2849 ( .A(N1030), .B(z2[148]), .Z(n1903) );
  NANDN U2850 ( .A(n3), .B(N1180), .Z(n1902) );
  NAND U2851 ( .A(n1904), .B(n1905), .Z(z3[147]) );
  NANDN U2852 ( .A(N1030), .B(z2[147]), .Z(n1905) );
  NANDN U2853 ( .A(n3), .B(N1179), .Z(n1904) );
  NAND U2854 ( .A(n1906), .B(n1907), .Z(z3[146]) );
  NANDN U2855 ( .A(N1030), .B(z2[146]), .Z(n1907) );
  NANDN U2856 ( .A(n3), .B(N1178), .Z(n1906) );
  NAND U2857 ( .A(n1908), .B(n1909), .Z(z3[145]) );
  NANDN U2858 ( .A(N1030), .B(z2[145]), .Z(n1909) );
  NANDN U2859 ( .A(n3), .B(N1177), .Z(n1908) );
  NAND U2860 ( .A(n1910), .B(n1911), .Z(z3[144]) );
  NANDN U2861 ( .A(N1030), .B(z2[144]), .Z(n1911) );
  NANDN U2862 ( .A(n3), .B(N1176), .Z(n1910) );
  NAND U2863 ( .A(n1912), .B(n1913), .Z(z3[143]) );
  NANDN U2864 ( .A(N1030), .B(z2[143]), .Z(n1913) );
  NANDN U2865 ( .A(n3), .B(N1175), .Z(n1912) );
  NAND U2866 ( .A(n1914), .B(n1915), .Z(z3[142]) );
  NANDN U2867 ( .A(N1030), .B(z2[142]), .Z(n1915) );
  NANDN U2868 ( .A(n3), .B(N1174), .Z(n1914) );
  NAND U2869 ( .A(n1916), .B(n1917), .Z(z3[141]) );
  NANDN U2870 ( .A(N1030), .B(z2[141]), .Z(n1917) );
  NANDN U2871 ( .A(n3), .B(N1173), .Z(n1916) );
  NAND U2872 ( .A(n1918), .B(n1919), .Z(z3[140]) );
  NANDN U2873 ( .A(N1030), .B(z2[140]), .Z(n1919) );
  NANDN U2874 ( .A(n3), .B(N1172), .Z(n1918) );
  NAND U2875 ( .A(n1920), .B(n1921), .Z(z3[13]) );
  NANDN U2876 ( .A(N1030), .B(z2[13]), .Z(n1921) );
  NANDN U2877 ( .A(n3), .B(N1045), .Z(n1920) );
  NAND U2878 ( .A(n1922), .B(n1923), .Z(z3[139]) );
  NANDN U2879 ( .A(N1030), .B(z2[139]), .Z(n1923) );
  NANDN U2880 ( .A(n3), .B(N1171), .Z(n1922) );
  NAND U2881 ( .A(n1924), .B(n1925), .Z(z3[138]) );
  NANDN U2882 ( .A(N1030), .B(z2[138]), .Z(n1925) );
  NANDN U2883 ( .A(n3), .B(N1170), .Z(n1924) );
  NAND U2884 ( .A(n1926), .B(n1927), .Z(z3[137]) );
  NANDN U2885 ( .A(N1030), .B(z2[137]), .Z(n1927) );
  NANDN U2886 ( .A(n3), .B(N1169), .Z(n1926) );
  NAND U2887 ( .A(n1928), .B(n1929), .Z(z3[136]) );
  NANDN U2888 ( .A(N1030), .B(z2[136]), .Z(n1929) );
  NANDN U2889 ( .A(n3), .B(N1168), .Z(n1928) );
  NAND U2890 ( .A(n1930), .B(n1931), .Z(z3[135]) );
  NANDN U2891 ( .A(N1030), .B(z2[135]), .Z(n1931) );
  NANDN U2892 ( .A(n3), .B(N1167), .Z(n1930) );
  NAND U2893 ( .A(n1932), .B(n1933), .Z(z3[134]) );
  NANDN U2894 ( .A(N1030), .B(z2[134]), .Z(n1933) );
  NANDN U2895 ( .A(n3), .B(N1166), .Z(n1932) );
  NAND U2896 ( .A(n1934), .B(n1935), .Z(z3[133]) );
  NANDN U2897 ( .A(N1030), .B(z2[133]), .Z(n1935) );
  NANDN U2898 ( .A(n3), .B(N1165), .Z(n1934) );
  NAND U2899 ( .A(n1936), .B(n1937), .Z(z3[132]) );
  NANDN U2900 ( .A(N1030), .B(z2[132]), .Z(n1937) );
  NANDN U2901 ( .A(n3), .B(N1164), .Z(n1936) );
  NAND U2902 ( .A(n1938), .B(n1939), .Z(z3[131]) );
  NANDN U2903 ( .A(N1030), .B(z2[131]), .Z(n1939) );
  NANDN U2904 ( .A(n3), .B(N1163), .Z(n1938) );
  NAND U2905 ( .A(n1940), .B(n1941), .Z(z3[130]) );
  NANDN U2906 ( .A(N1030), .B(z2[130]), .Z(n1941) );
  NANDN U2907 ( .A(n3), .B(N1162), .Z(n1940) );
  NAND U2908 ( .A(n1942), .B(n1943), .Z(z3[12]) );
  NANDN U2909 ( .A(N1030), .B(z2[12]), .Z(n1943) );
  NANDN U2910 ( .A(n3), .B(N1044), .Z(n1942) );
  NAND U2911 ( .A(n1944), .B(n1945), .Z(z3[129]) );
  NANDN U2912 ( .A(N1030), .B(z2[129]), .Z(n1945) );
  NANDN U2913 ( .A(n3), .B(N1161), .Z(n1944) );
  NAND U2914 ( .A(n1946), .B(n1947), .Z(z3[128]) );
  NANDN U2915 ( .A(N1030), .B(z2[128]), .Z(n1947) );
  NANDN U2916 ( .A(n3), .B(N1160), .Z(n1946) );
  NAND U2917 ( .A(n1948), .B(n1949), .Z(z3[127]) );
  NANDN U2918 ( .A(N1030), .B(z2[127]), .Z(n1949) );
  NANDN U2919 ( .A(n3), .B(N1159), .Z(n1948) );
  NAND U2920 ( .A(n1950), .B(n1951), .Z(z3[126]) );
  NANDN U2921 ( .A(N1030), .B(z2[126]), .Z(n1951) );
  NANDN U2922 ( .A(n3), .B(N1158), .Z(n1950) );
  NAND U2923 ( .A(n1952), .B(n1953), .Z(z3[125]) );
  NANDN U2924 ( .A(N1030), .B(z2[125]), .Z(n1953) );
  NANDN U2925 ( .A(n3), .B(N1157), .Z(n1952) );
  NAND U2926 ( .A(n1954), .B(n1955), .Z(z3[124]) );
  NANDN U2927 ( .A(N1030), .B(z2[124]), .Z(n1955) );
  NANDN U2928 ( .A(n3), .B(N1156), .Z(n1954) );
  NAND U2929 ( .A(n1956), .B(n1957), .Z(z3[123]) );
  NANDN U2930 ( .A(N1030), .B(z2[123]), .Z(n1957) );
  NANDN U2931 ( .A(n3), .B(N1155), .Z(n1956) );
  NAND U2932 ( .A(n1958), .B(n1959), .Z(z3[122]) );
  NANDN U2933 ( .A(N1030), .B(z2[122]), .Z(n1959) );
  NANDN U2934 ( .A(n3), .B(N1154), .Z(n1958) );
  NAND U2935 ( .A(n1960), .B(n1961), .Z(z3[121]) );
  NANDN U2936 ( .A(N1030), .B(z2[121]), .Z(n1961) );
  NANDN U2937 ( .A(n3), .B(N1153), .Z(n1960) );
  NAND U2938 ( .A(n1962), .B(n1963), .Z(z3[120]) );
  NANDN U2939 ( .A(N1030), .B(z2[120]), .Z(n1963) );
  NANDN U2940 ( .A(n3), .B(N1152), .Z(n1962) );
  NAND U2941 ( .A(n1964), .B(n1965), .Z(z3[11]) );
  NANDN U2942 ( .A(N1030), .B(z2[11]), .Z(n1965) );
  NANDN U2943 ( .A(n3), .B(N1043), .Z(n1964) );
  NAND U2944 ( .A(n1966), .B(n1967), .Z(z3[119]) );
  NANDN U2945 ( .A(N1030), .B(z2[119]), .Z(n1967) );
  NANDN U2946 ( .A(n3), .B(N1151), .Z(n1966) );
  NAND U2947 ( .A(n1968), .B(n1969), .Z(z3[118]) );
  NANDN U2948 ( .A(N1030), .B(z2[118]), .Z(n1969) );
  NANDN U2949 ( .A(n3), .B(N1150), .Z(n1968) );
  NAND U2950 ( .A(n1970), .B(n1971), .Z(z3[117]) );
  NANDN U2951 ( .A(N1030), .B(z2[117]), .Z(n1971) );
  NANDN U2952 ( .A(n3), .B(N1149), .Z(n1970) );
  NAND U2953 ( .A(n1972), .B(n1973), .Z(z3[116]) );
  NANDN U2954 ( .A(N1030), .B(z2[116]), .Z(n1973) );
  NANDN U2955 ( .A(n3), .B(N1148), .Z(n1972) );
  NAND U2956 ( .A(n1974), .B(n1975), .Z(z3[115]) );
  NANDN U2957 ( .A(N1030), .B(z2[115]), .Z(n1975) );
  NANDN U2958 ( .A(n3), .B(N1147), .Z(n1974) );
  NAND U2959 ( .A(n1976), .B(n1977), .Z(z3[114]) );
  NANDN U2960 ( .A(N1030), .B(z2[114]), .Z(n1977) );
  NANDN U2961 ( .A(n3), .B(N1146), .Z(n1976) );
  NAND U2962 ( .A(n1978), .B(n1979), .Z(z3[113]) );
  NANDN U2963 ( .A(N1030), .B(z2[113]), .Z(n1979) );
  NANDN U2964 ( .A(n3), .B(N1145), .Z(n1978) );
  NAND U2965 ( .A(n1980), .B(n1981), .Z(z3[112]) );
  NANDN U2966 ( .A(N1030), .B(z2[112]), .Z(n1981) );
  NANDN U2967 ( .A(n3), .B(N1144), .Z(n1980) );
  NAND U2968 ( .A(n1982), .B(n1983), .Z(z3[111]) );
  NANDN U2969 ( .A(N1030), .B(z2[111]), .Z(n1983) );
  NANDN U2970 ( .A(n3), .B(N1143), .Z(n1982) );
  NAND U2971 ( .A(n1984), .B(n1985), .Z(z3[110]) );
  NANDN U2972 ( .A(N1030), .B(z2[110]), .Z(n1985) );
  NANDN U2973 ( .A(n3), .B(N1142), .Z(n1984) );
  NAND U2974 ( .A(n1986), .B(n1987), .Z(z3[10]) );
  NANDN U2975 ( .A(N1030), .B(z2[10]), .Z(n1987) );
  NANDN U2976 ( .A(n3), .B(N1042), .Z(n1986) );
  NAND U2977 ( .A(n1988), .B(n1989), .Z(z3[109]) );
  NANDN U2978 ( .A(N1030), .B(z2[109]), .Z(n1989) );
  NANDN U2979 ( .A(n3), .B(N1141), .Z(n1988) );
  NAND U2980 ( .A(n1990), .B(n1991), .Z(z3[108]) );
  NANDN U2981 ( .A(N1030), .B(z2[108]), .Z(n1991) );
  NANDN U2982 ( .A(n3), .B(N1140), .Z(n1990) );
  NAND U2983 ( .A(n1992), .B(n1993), .Z(z3[107]) );
  NANDN U2984 ( .A(N1030), .B(z2[107]), .Z(n1993) );
  NANDN U2985 ( .A(n3), .B(N1139), .Z(n1992) );
  NAND U2986 ( .A(n1994), .B(n1995), .Z(z3[106]) );
  NANDN U2987 ( .A(N1030), .B(z2[106]), .Z(n1995) );
  NANDN U2988 ( .A(n3), .B(N1138), .Z(n1994) );
  NAND U2989 ( .A(n1996), .B(n1997), .Z(z3[105]) );
  NANDN U2990 ( .A(N1030), .B(z2[105]), .Z(n1997) );
  NANDN U2991 ( .A(n3), .B(N1137), .Z(n1996) );
  NAND U2992 ( .A(n1998), .B(n1999), .Z(z3[104]) );
  NANDN U2993 ( .A(N1030), .B(z2[104]), .Z(n1999) );
  NANDN U2994 ( .A(n3), .B(N1136), .Z(n1998) );
  NAND U2995 ( .A(n2000), .B(n2001), .Z(z3[103]) );
  NANDN U2996 ( .A(N1030), .B(z2[103]), .Z(n2001) );
  NANDN U2997 ( .A(n3), .B(N1135), .Z(n2000) );
  NAND U2998 ( .A(n2002), .B(n2003), .Z(z3[102]) );
  NANDN U2999 ( .A(N1030), .B(z2[102]), .Z(n2003) );
  NANDN U3000 ( .A(n3), .B(N1134), .Z(n2002) );
  NAND U3001 ( .A(n2004), .B(n2005), .Z(z3[1025]) );
  NANDN U3002 ( .A(N1030), .B(z2[1025]), .Z(n2005) );
  NANDN U3003 ( .A(n3), .B(N2057), .Z(n2004) );
  NAND U3004 ( .A(n2006), .B(n2007), .Z(z3[1024]) );
  NANDN U3005 ( .A(N1030), .B(z2[1024]), .Z(n2007) );
  NANDN U3006 ( .A(n3), .B(N2056), .Z(n2006) );
  NAND U3007 ( .A(n2008), .B(n2009), .Z(z3[1023]) );
  NANDN U3008 ( .A(N1030), .B(z2[1023]), .Z(n2009) );
  NANDN U3009 ( .A(n3), .B(N2055), .Z(n2008) );
  NAND U3010 ( .A(n2010), .B(n2011), .Z(z3[1022]) );
  NANDN U3011 ( .A(N1030), .B(z2[1022]), .Z(n2011) );
  NANDN U3012 ( .A(n3), .B(N2054), .Z(n2010) );
  NAND U3013 ( .A(n2012), .B(n2013), .Z(z3[1021]) );
  NANDN U3014 ( .A(N1030), .B(z2[1021]), .Z(n2013) );
  NANDN U3015 ( .A(n3), .B(N2053), .Z(n2012) );
  NAND U3016 ( .A(n2014), .B(n2015), .Z(z3[1020]) );
  NANDN U3017 ( .A(N1030), .B(z2[1020]), .Z(n2015) );
  NANDN U3018 ( .A(n3), .B(N2052), .Z(n2014) );
  NAND U3019 ( .A(n2016), .B(n2017), .Z(z3[101]) );
  NANDN U3020 ( .A(N1030), .B(z2[101]), .Z(n2017) );
  NANDN U3021 ( .A(n3), .B(N1133), .Z(n2016) );
  NAND U3022 ( .A(n2018), .B(n2019), .Z(z3[1019]) );
  NANDN U3023 ( .A(N1030), .B(z2[1019]), .Z(n2019) );
  NANDN U3024 ( .A(n3), .B(N2051), .Z(n2018) );
  NAND U3025 ( .A(n2020), .B(n2021), .Z(z3[1018]) );
  NANDN U3026 ( .A(N1030), .B(z2[1018]), .Z(n2021) );
  NANDN U3027 ( .A(n3), .B(N2050), .Z(n2020) );
  NAND U3028 ( .A(n2022), .B(n2023), .Z(z3[1017]) );
  NANDN U3029 ( .A(N1030), .B(z2[1017]), .Z(n2023) );
  NANDN U3030 ( .A(n3), .B(N2049), .Z(n2022) );
  NAND U3031 ( .A(n2024), .B(n2025), .Z(z3[1016]) );
  NANDN U3032 ( .A(N1030), .B(z2[1016]), .Z(n2025) );
  NANDN U3033 ( .A(n3), .B(N2048), .Z(n2024) );
  NAND U3034 ( .A(n2026), .B(n2027), .Z(z3[1015]) );
  NANDN U3035 ( .A(N1030), .B(z2[1015]), .Z(n2027) );
  NANDN U3036 ( .A(n3), .B(N2047), .Z(n2026) );
  NAND U3037 ( .A(n2028), .B(n2029), .Z(z3[1014]) );
  NANDN U3038 ( .A(N1030), .B(z2[1014]), .Z(n2029) );
  NANDN U3039 ( .A(n3), .B(N2046), .Z(n2028) );
  NAND U3040 ( .A(n2030), .B(n2031), .Z(z3[1013]) );
  NANDN U3041 ( .A(N1030), .B(z2[1013]), .Z(n2031) );
  NANDN U3042 ( .A(n3), .B(N2045), .Z(n2030) );
  NAND U3043 ( .A(n2032), .B(n2033), .Z(z3[1012]) );
  NANDN U3044 ( .A(N1030), .B(z2[1012]), .Z(n2033) );
  NANDN U3045 ( .A(n3), .B(N2044), .Z(n2032) );
  NAND U3046 ( .A(n2034), .B(n2035), .Z(z3[1011]) );
  NANDN U3047 ( .A(N1030), .B(z2[1011]), .Z(n2035) );
  NANDN U3048 ( .A(n3), .B(N2043), .Z(n2034) );
  NAND U3049 ( .A(n2036), .B(n2037), .Z(z3[1010]) );
  NANDN U3050 ( .A(N1030), .B(z2[1010]), .Z(n2037) );
  NANDN U3051 ( .A(n3), .B(N2042), .Z(n2036) );
  NAND U3052 ( .A(n2038), .B(n2039), .Z(z3[100]) );
  NANDN U3053 ( .A(N1030), .B(z2[100]), .Z(n2039) );
  NANDN U3054 ( .A(n3), .B(N1132), .Z(n2038) );
  NAND U3055 ( .A(n2040), .B(n2041), .Z(z3[1009]) );
  NANDN U3056 ( .A(N1030), .B(z2[1009]), .Z(n2041) );
  NANDN U3057 ( .A(n3), .B(N2041), .Z(n2040) );
  NAND U3058 ( .A(n2042), .B(n2043), .Z(z3[1008]) );
  NANDN U3059 ( .A(N1030), .B(z2[1008]), .Z(n2043) );
  NANDN U3060 ( .A(n3), .B(N2040), .Z(n2042) );
  NAND U3061 ( .A(n2044), .B(n2045), .Z(z3[1007]) );
  NANDN U3062 ( .A(N1030), .B(z2[1007]), .Z(n2045) );
  NANDN U3063 ( .A(n3), .B(N2039), .Z(n2044) );
  NAND U3064 ( .A(n2046), .B(n2047), .Z(z3[1006]) );
  NANDN U3065 ( .A(N1030), .B(z2[1006]), .Z(n2047) );
  NANDN U3066 ( .A(n3), .B(N2038), .Z(n2046) );
  NAND U3067 ( .A(n2048), .B(n2049), .Z(z3[1005]) );
  NANDN U3068 ( .A(N1030), .B(z2[1005]), .Z(n2049) );
  NANDN U3069 ( .A(n3), .B(N2037), .Z(n2048) );
  NAND U3070 ( .A(n2050), .B(n2051), .Z(z3[1004]) );
  NANDN U3071 ( .A(N1030), .B(z2[1004]), .Z(n2051) );
  NANDN U3072 ( .A(n3), .B(N2036), .Z(n2050) );
  NAND U3073 ( .A(n2052), .B(n2053), .Z(z3[1003]) );
  NANDN U3074 ( .A(N1030), .B(z2[1003]), .Z(n2053) );
  NANDN U3075 ( .A(n3), .B(N2035), .Z(n2052) );
  NAND U3076 ( .A(n2054), .B(n2055), .Z(z3[1002]) );
  NANDN U3077 ( .A(N1030), .B(z2[1002]), .Z(n2055) );
  NANDN U3078 ( .A(n3), .B(N2034), .Z(n2054) );
  NAND U3079 ( .A(n2056), .B(n2057), .Z(z3[1001]) );
  NANDN U3080 ( .A(N1030), .B(z2[1001]), .Z(n2057) );
  NANDN U3081 ( .A(n3), .B(N2033), .Z(n2056) );
  NAND U3082 ( .A(n2058), .B(n2059), .Z(z3[1000]) );
  NANDN U3083 ( .A(N1030), .B(z2[1000]), .Z(n2059) );
  NANDN U3084 ( .A(n3), .B(N2032), .Z(n2058) );
  NAND U3085 ( .A(n2060), .B(n2061), .Z(z3[0]) );
  NANDN U3086 ( .A(N1030), .B(z2[0]), .Z(n2061) );
  NANDN U3087 ( .A(n3), .B(N1032), .Z(n2060) );
  IV U3088 ( .A(N1030), .Z(n3) );
  NAND U3089 ( .A(n2062), .B(n2063), .Z(z2[9]) );
  NANDN U3090 ( .A(xregN_1), .B(zin[8]), .Z(n2063) );
  NAND U3091 ( .A(N13), .B(xregN_1), .Z(n2062) );
  NAND U3092 ( .A(n2064), .B(n2065), .Z(z2[99]) );
  NANDN U3093 ( .A(xregN_1), .B(zin[98]), .Z(n2065) );
  NAND U3094 ( .A(N103), .B(xregN_1), .Z(n2064) );
  NAND U3095 ( .A(n2066), .B(n2067), .Z(z2[999]) );
  NANDN U3096 ( .A(xregN_1), .B(zin[998]), .Z(n2067) );
  NAND U3097 ( .A(N1003), .B(xregN_1), .Z(n2066) );
  NAND U3098 ( .A(n2068), .B(n2069), .Z(z2[998]) );
  NANDN U3099 ( .A(xregN_1), .B(zin[997]), .Z(n2069) );
  NAND U3100 ( .A(N1002), .B(xregN_1), .Z(n2068) );
  NAND U3101 ( .A(n2070), .B(n2071), .Z(z2[997]) );
  NANDN U3102 ( .A(xregN_1), .B(zin[996]), .Z(n2071) );
  NAND U3103 ( .A(N1001), .B(xregN_1), .Z(n2070) );
  NAND U3104 ( .A(n2072), .B(n2073), .Z(z2[996]) );
  NANDN U3105 ( .A(xregN_1), .B(zin[995]), .Z(n2073) );
  NAND U3106 ( .A(N1000), .B(xregN_1), .Z(n2072) );
  NAND U3107 ( .A(n2074), .B(n2075), .Z(z2[995]) );
  NANDN U3108 ( .A(xregN_1), .B(zin[994]), .Z(n2075) );
  NAND U3109 ( .A(N999), .B(xregN_1), .Z(n2074) );
  NAND U3110 ( .A(n2076), .B(n2077), .Z(z2[994]) );
  NANDN U3111 ( .A(xregN_1), .B(zin[993]), .Z(n2077) );
  NAND U3112 ( .A(N998), .B(xregN_1), .Z(n2076) );
  NAND U3113 ( .A(n2078), .B(n2079), .Z(z2[993]) );
  NANDN U3114 ( .A(xregN_1), .B(zin[992]), .Z(n2079) );
  NAND U3115 ( .A(N997), .B(xregN_1), .Z(n2078) );
  NAND U3116 ( .A(n2080), .B(n2081), .Z(z2[992]) );
  NANDN U3117 ( .A(xregN_1), .B(zin[991]), .Z(n2081) );
  NAND U3118 ( .A(N996), .B(xregN_1), .Z(n2080) );
  NAND U3119 ( .A(n2082), .B(n2083), .Z(z2[991]) );
  NANDN U3120 ( .A(xregN_1), .B(zin[990]), .Z(n2083) );
  NAND U3121 ( .A(N995), .B(xregN_1), .Z(n2082) );
  NAND U3122 ( .A(n2084), .B(n2085), .Z(z2[990]) );
  NANDN U3123 ( .A(xregN_1), .B(zin[989]), .Z(n2085) );
  NAND U3124 ( .A(N994), .B(xregN_1), .Z(n2084) );
  NAND U3125 ( .A(n2086), .B(n2087), .Z(z2[98]) );
  NANDN U3126 ( .A(xregN_1), .B(zin[97]), .Z(n2087) );
  NAND U3127 ( .A(N102), .B(xregN_1), .Z(n2086) );
  NAND U3128 ( .A(n2088), .B(n2089), .Z(z2[989]) );
  NANDN U3129 ( .A(xregN_1), .B(zin[988]), .Z(n2089) );
  NAND U3130 ( .A(N993), .B(xregN_1), .Z(n2088) );
  NAND U3131 ( .A(n2090), .B(n2091), .Z(z2[988]) );
  NANDN U3132 ( .A(xregN_1), .B(zin[987]), .Z(n2091) );
  NAND U3133 ( .A(N992), .B(xregN_1), .Z(n2090) );
  NAND U3134 ( .A(n2092), .B(n2093), .Z(z2[987]) );
  NANDN U3135 ( .A(xregN_1), .B(zin[986]), .Z(n2093) );
  NAND U3136 ( .A(N991), .B(xregN_1), .Z(n2092) );
  NAND U3137 ( .A(n2094), .B(n2095), .Z(z2[986]) );
  NANDN U3138 ( .A(xregN_1), .B(zin[985]), .Z(n2095) );
  NAND U3139 ( .A(N990), .B(xregN_1), .Z(n2094) );
  NAND U3140 ( .A(n2096), .B(n2097), .Z(z2[985]) );
  NANDN U3141 ( .A(xregN_1), .B(zin[984]), .Z(n2097) );
  NAND U3142 ( .A(N989), .B(xregN_1), .Z(n2096) );
  NAND U3143 ( .A(n2098), .B(n2099), .Z(z2[984]) );
  NANDN U3144 ( .A(xregN_1), .B(zin[983]), .Z(n2099) );
  NAND U3145 ( .A(N988), .B(xregN_1), .Z(n2098) );
  NAND U3146 ( .A(n2100), .B(n2101), .Z(z2[983]) );
  NANDN U3147 ( .A(xregN_1), .B(zin[982]), .Z(n2101) );
  NAND U3148 ( .A(N987), .B(xregN_1), .Z(n2100) );
  NAND U3149 ( .A(n2102), .B(n2103), .Z(z2[982]) );
  NANDN U3150 ( .A(xregN_1), .B(zin[981]), .Z(n2103) );
  NAND U3151 ( .A(N986), .B(xregN_1), .Z(n2102) );
  NAND U3152 ( .A(n2104), .B(n2105), .Z(z2[981]) );
  NANDN U3153 ( .A(xregN_1), .B(zin[980]), .Z(n2105) );
  NAND U3154 ( .A(N985), .B(xregN_1), .Z(n2104) );
  NAND U3155 ( .A(n2106), .B(n2107), .Z(z2[980]) );
  NANDN U3156 ( .A(xregN_1), .B(zin[979]), .Z(n2107) );
  NAND U3157 ( .A(N984), .B(xregN_1), .Z(n2106) );
  NAND U3158 ( .A(n2108), .B(n2109), .Z(z2[97]) );
  NANDN U3159 ( .A(xregN_1), .B(zin[96]), .Z(n2109) );
  NAND U3160 ( .A(N101), .B(xregN_1), .Z(n2108) );
  NAND U3161 ( .A(n2110), .B(n2111), .Z(z2[979]) );
  NANDN U3162 ( .A(xregN_1), .B(zin[978]), .Z(n2111) );
  NAND U3163 ( .A(N983), .B(xregN_1), .Z(n2110) );
  NAND U3164 ( .A(n2112), .B(n2113), .Z(z2[978]) );
  NANDN U3165 ( .A(xregN_1), .B(zin[977]), .Z(n2113) );
  NAND U3166 ( .A(N982), .B(xregN_1), .Z(n2112) );
  NAND U3167 ( .A(n2114), .B(n2115), .Z(z2[977]) );
  NANDN U3168 ( .A(xregN_1), .B(zin[976]), .Z(n2115) );
  NAND U3169 ( .A(N981), .B(xregN_1), .Z(n2114) );
  NAND U3170 ( .A(n2116), .B(n2117), .Z(z2[976]) );
  NANDN U3171 ( .A(xregN_1), .B(zin[975]), .Z(n2117) );
  NAND U3172 ( .A(N980), .B(xregN_1), .Z(n2116) );
  NAND U3173 ( .A(n2118), .B(n2119), .Z(z2[975]) );
  NANDN U3174 ( .A(xregN_1), .B(zin[974]), .Z(n2119) );
  NAND U3175 ( .A(N979), .B(xregN_1), .Z(n2118) );
  NAND U3176 ( .A(n2120), .B(n2121), .Z(z2[974]) );
  NANDN U3177 ( .A(xregN_1), .B(zin[973]), .Z(n2121) );
  NAND U3178 ( .A(N978), .B(xregN_1), .Z(n2120) );
  NAND U3179 ( .A(n2122), .B(n2123), .Z(z2[973]) );
  NANDN U3180 ( .A(xregN_1), .B(zin[972]), .Z(n2123) );
  NAND U3181 ( .A(N977), .B(xregN_1), .Z(n2122) );
  NAND U3182 ( .A(n2124), .B(n2125), .Z(z2[972]) );
  NANDN U3183 ( .A(xregN_1), .B(zin[971]), .Z(n2125) );
  NAND U3184 ( .A(N976), .B(xregN_1), .Z(n2124) );
  NAND U3185 ( .A(n2126), .B(n2127), .Z(z2[971]) );
  NANDN U3186 ( .A(xregN_1), .B(zin[970]), .Z(n2127) );
  NAND U3187 ( .A(N975), .B(xregN_1), .Z(n2126) );
  NAND U3188 ( .A(n2128), .B(n2129), .Z(z2[970]) );
  NANDN U3189 ( .A(xregN_1), .B(zin[969]), .Z(n2129) );
  NAND U3190 ( .A(N974), .B(xregN_1), .Z(n2128) );
  NAND U3191 ( .A(n2130), .B(n2131), .Z(z2[96]) );
  NANDN U3192 ( .A(xregN_1), .B(zin[95]), .Z(n2131) );
  NAND U3193 ( .A(N100), .B(xregN_1), .Z(n2130) );
  NAND U3194 ( .A(n2132), .B(n2133), .Z(z2[969]) );
  NANDN U3195 ( .A(xregN_1), .B(zin[968]), .Z(n2133) );
  NAND U3196 ( .A(N973), .B(xregN_1), .Z(n2132) );
  NAND U3197 ( .A(n2134), .B(n2135), .Z(z2[968]) );
  NANDN U3198 ( .A(xregN_1), .B(zin[967]), .Z(n2135) );
  NAND U3199 ( .A(N972), .B(xregN_1), .Z(n2134) );
  NAND U3200 ( .A(n2136), .B(n2137), .Z(z2[967]) );
  NANDN U3201 ( .A(xregN_1), .B(zin[966]), .Z(n2137) );
  NAND U3202 ( .A(N971), .B(xregN_1), .Z(n2136) );
  NAND U3203 ( .A(n2138), .B(n2139), .Z(z2[966]) );
  NANDN U3204 ( .A(xregN_1), .B(zin[965]), .Z(n2139) );
  NAND U3205 ( .A(N970), .B(xregN_1), .Z(n2138) );
  NAND U3206 ( .A(n2140), .B(n2141), .Z(z2[965]) );
  NANDN U3207 ( .A(xregN_1), .B(zin[964]), .Z(n2141) );
  NAND U3208 ( .A(N969), .B(xregN_1), .Z(n2140) );
  NAND U3209 ( .A(n2142), .B(n2143), .Z(z2[964]) );
  NANDN U3210 ( .A(xregN_1), .B(zin[963]), .Z(n2143) );
  NAND U3211 ( .A(N968), .B(xregN_1), .Z(n2142) );
  NAND U3212 ( .A(n2144), .B(n2145), .Z(z2[963]) );
  NANDN U3213 ( .A(xregN_1), .B(zin[962]), .Z(n2145) );
  NAND U3214 ( .A(N967), .B(xregN_1), .Z(n2144) );
  NAND U3215 ( .A(n2146), .B(n2147), .Z(z2[962]) );
  NANDN U3216 ( .A(xregN_1), .B(zin[961]), .Z(n2147) );
  NAND U3217 ( .A(N966), .B(xregN_1), .Z(n2146) );
  NAND U3218 ( .A(n2148), .B(n2149), .Z(z2[961]) );
  NANDN U3219 ( .A(xregN_1), .B(zin[960]), .Z(n2149) );
  NAND U3220 ( .A(N965), .B(xregN_1), .Z(n2148) );
  NAND U3221 ( .A(n2150), .B(n2151), .Z(z2[960]) );
  NANDN U3222 ( .A(xregN_1), .B(zin[959]), .Z(n2151) );
  NAND U3223 ( .A(N964), .B(xregN_1), .Z(n2150) );
  NAND U3224 ( .A(n2152), .B(n2153), .Z(z2[95]) );
  NANDN U3225 ( .A(xregN_1), .B(zin[94]), .Z(n2153) );
  NAND U3226 ( .A(N99), .B(xregN_1), .Z(n2152) );
  NAND U3227 ( .A(n2154), .B(n2155), .Z(z2[959]) );
  NANDN U3228 ( .A(xregN_1), .B(zin[958]), .Z(n2155) );
  NAND U3229 ( .A(N963), .B(xregN_1), .Z(n2154) );
  NAND U3230 ( .A(n2156), .B(n2157), .Z(z2[958]) );
  NANDN U3231 ( .A(xregN_1), .B(zin[957]), .Z(n2157) );
  NAND U3232 ( .A(N962), .B(xregN_1), .Z(n2156) );
  NAND U3233 ( .A(n2158), .B(n2159), .Z(z2[957]) );
  NANDN U3234 ( .A(xregN_1), .B(zin[956]), .Z(n2159) );
  NAND U3235 ( .A(N961), .B(xregN_1), .Z(n2158) );
  NAND U3236 ( .A(n2160), .B(n2161), .Z(z2[956]) );
  NANDN U3237 ( .A(xregN_1), .B(zin[955]), .Z(n2161) );
  NAND U3238 ( .A(N960), .B(xregN_1), .Z(n2160) );
  NAND U3239 ( .A(n2162), .B(n2163), .Z(z2[955]) );
  NANDN U3240 ( .A(xregN_1), .B(zin[954]), .Z(n2163) );
  NAND U3241 ( .A(N959), .B(xregN_1), .Z(n2162) );
  NAND U3242 ( .A(n2164), .B(n2165), .Z(z2[954]) );
  NANDN U3243 ( .A(xregN_1), .B(zin[953]), .Z(n2165) );
  NAND U3244 ( .A(N958), .B(xregN_1), .Z(n2164) );
  NAND U3245 ( .A(n2166), .B(n2167), .Z(z2[953]) );
  NANDN U3246 ( .A(xregN_1), .B(zin[952]), .Z(n2167) );
  NAND U3247 ( .A(N957), .B(xregN_1), .Z(n2166) );
  NAND U3248 ( .A(n2168), .B(n2169), .Z(z2[952]) );
  NANDN U3249 ( .A(xregN_1), .B(zin[951]), .Z(n2169) );
  NAND U3250 ( .A(N956), .B(xregN_1), .Z(n2168) );
  NAND U3251 ( .A(n2170), .B(n2171), .Z(z2[951]) );
  NANDN U3252 ( .A(xregN_1), .B(zin[950]), .Z(n2171) );
  NAND U3253 ( .A(N955), .B(xregN_1), .Z(n2170) );
  NAND U3254 ( .A(n2172), .B(n2173), .Z(z2[950]) );
  NANDN U3255 ( .A(xregN_1), .B(zin[949]), .Z(n2173) );
  NAND U3256 ( .A(N954), .B(xregN_1), .Z(n2172) );
  NAND U3257 ( .A(n2174), .B(n2175), .Z(z2[94]) );
  NANDN U3258 ( .A(xregN_1), .B(zin[93]), .Z(n2175) );
  NAND U3259 ( .A(N98), .B(xregN_1), .Z(n2174) );
  NAND U3260 ( .A(n2176), .B(n2177), .Z(z2[949]) );
  NANDN U3261 ( .A(xregN_1), .B(zin[948]), .Z(n2177) );
  NAND U3262 ( .A(N953), .B(xregN_1), .Z(n2176) );
  NAND U3263 ( .A(n2178), .B(n2179), .Z(z2[948]) );
  NANDN U3264 ( .A(xregN_1), .B(zin[947]), .Z(n2179) );
  NAND U3265 ( .A(N952), .B(xregN_1), .Z(n2178) );
  NAND U3266 ( .A(n2180), .B(n2181), .Z(z2[947]) );
  NANDN U3267 ( .A(xregN_1), .B(zin[946]), .Z(n2181) );
  NAND U3268 ( .A(N951), .B(xregN_1), .Z(n2180) );
  NAND U3269 ( .A(n2182), .B(n2183), .Z(z2[946]) );
  NANDN U3270 ( .A(xregN_1), .B(zin[945]), .Z(n2183) );
  NAND U3271 ( .A(N950), .B(xregN_1), .Z(n2182) );
  NAND U3272 ( .A(n2184), .B(n2185), .Z(z2[945]) );
  NANDN U3273 ( .A(xregN_1), .B(zin[944]), .Z(n2185) );
  NAND U3274 ( .A(N949), .B(xregN_1), .Z(n2184) );
  NAND U3275 ( .A(n2186), .B(n2187), .Z(z2[944]) );
  NANDN U3276 ( .A(xregN_1), .B(zin[943]), .Z(n2187) );
  NAND U3277 ( .A(N948), .B(xregN_1), .Z(n2186) );
  NAND U3278 ( .A(n2188), .B(n2189), .Z(z2[943]) );
  NANDN U3279 ( .A(xregN_1), .B(zin[942]), .Z(n2189) );
  NAND U3280 ( .A(N947), .B(xregN_1), .Z(n2188) );
  NAND U3281 ( .A(n2190), .B(n2191), .Z(z2[942]) );
  NANDN U3282 ( .A(xregN_1), .B(zin[941]), .Z(n2191) );
  NAND U3283 ( .A(N946), .B(xregN_1), .Z(n2190) );
  NAND U3284 ( .A(n2192), .B(n2193), .Z(z2[941]) );
  NANDN U3285 ( .A(xregN_1), .B(zin[940]), .Z(n2193) );
  NAND U3286 ( .A(N945), .B(xregN_1), .Z(n2192) );
  NAND U3287 ( .A(n2194), .B(n2195), .Z(z2[940]) );
  NANDN U3288 ( .A(xregN_1), .B(zin[939]), .Z(n2195) );
  NAND U3289 ( .A(N944), .B(xregN_1), .Z(n2194) );
  NAND U3290 ( .A(n2196), .B(n2197), .Z(z2[93]) );
  NANDN U3291 ( .A(xregN_1), .B(zin[92]), .Z(n2197) );
  NAND U3292 ( .A(N97), .B(xregN_1), .Z(n2196) );
  NAND U3293 ( .A(n2198), .B(n2199), .Z(z2[939]) );
  NANDN U3294 ( .A(xregN_1), .B(zin[938]), .Z(n2199) );
  NAND U3295 ( .A(N943), .B(xregN_1), .Z(n2198) );
  NAND U3296 ( .A(n2200), .B(n2201), .Z(z2[938]) );
  NANDN U3297 ( .A(xregN_1), .B(zin[937]), .Z(n2201) );
  NAND U3298 ( .A(N942), .B(xregN_1), .Z(n2200) );
  NAND U3299 ( .A(n2202), .B(n2203), .Z(z2[937]) );
  NANDN U3300 ( .A(xregN_1), .B(zin[936]), .Z(n2203) );
  NAND U3301 ( .A(N941), .B(xregN_1), .Z(n2202) );
  NAND U3302 ( .A(n2204), .B(n2205), .Z(z2[936]) );
  NANDN U3303 ( .A(xregN_1), .B(zin[935]), .Z(n2205) );
  NAND U3304 ( .A(N940), .B(xregN_1), .Z(n2204) );
  NAND U3305 ( .A(n2206), .B(n2207), .Z(z2[935]) );
  NANDN U3306 ( .A(xregN_1), .B(zin[934]), .Z(n2207) );
  NAND U3307 ( .A(N939), .B(xregN_1), .Z(n2206) );
  NAND U3308 ( .A(n2208), .B(n2209), .Z(z2[934]) );
  NANDN U3309 ( .A(xregN_1), .B(zin[933]), .Z(n2209) );
  NAND U3310 ( .A(N938), .B(xregN_1), .Z(n2208) );
  NAND U3311 ( .A(n2210), .B(n2211), .Z(z2[933]) );
  NANDN U3312 ( .A(xregN_1), .B(zin[932]), .Z(n2211) );
  NAND U3313 ( .A(N937), .B(xregN_1), .Z(n2210) );
  NAND U3314 ( .A(n2212), .B(n2213), .Z(z2[932]) );
  NANDN U3315 ( .A(xregN_1), .B(zin[931]), .Z(n2213) );
  NAND U3316 ( .A(N936), .B(xregN_1), .Z(n2212) );
  NAND U3317 ( .A(n2214), .B(n2215), .Z(z2[931]) );
  NANDN U3318 ( .A(xregN_1), .B(zin[930]), .Z(n2215) );
  NAND U3319 ( .A(N935), .B(xregN_1), .Z(n2214) );
  NAND U3320 ( .A(n2216), .B(n2217), .Z(z2[930]) );
  NANDN U3321 ( .A(xregN_1), .B(zin[929]), .Z(n2217) );
  NAND U3322 ( .A(N934), .B(xregN_1), .Z(n2216) );
  NAND U3323 ( .A(n2218), .B(n2219), .Z(z2[92]) );
  NANDN U3324 ( .A(xregN_1), .B(zin[91]), .Z(n2219) );
  NAND U3325 ( .A(N96), .B(xregN_1), .Z(n2218) );
  NAND U3326 ( .A(n2220), .B(n2221), .Z(z2[929]) );
  NANDN U3327 ( .A(xregN_1), .B(zin[928]), .Z(n2221) );
  NAND U3328 ( .A(N933), .B(xregN_1), .Z(n2220) );
  NAND U3329 ( .A(n2222), .B(n2223), .Z(z2[928]) );
  NANDN U3330 ( .A(xregN_1), .B(zin[927]), .Z(n2223) );
  NAND U3331 ( .A(N932), .B(xregN_1), .Z(n2222) );
  NAND U3332 ( .A(n2224), .B(n2225), .Z(z2[927]) );
  NANDN U3333 ( .A(xregN_1), .B(zin[926]), .Z(n2225) );
  NAND U3334 ( .A(N931), .B(xregN_1), .Z(n2224) );
  NAND U3335 ( .A(n2226), .B(n2227), .Z(z2[926]) );
  NANDN U3336 ( .A(xregN_1), .B(zin[925]), .Z(n2227) );
  NAND U3337 ( .A(N930), .B(xregN_1), .Z(n2226) );
  NAND U3338 ( .A(n2228), .B(n2229), .Z(z2[925]) );
  NANDN U3339 ( .A(xregN_1), .B(zin[924]), .Z(n2229) );
  NAND U3340 ( .A(N929), .B(xregN_1), .Z(n2228) );
  NAND U3341 ( .A(n2230), .B(n2231), .Z(z2[924]) );
  NANDN U3342 ( .A(xregN_1), .B(zin[923]), .Z(n2231) );
  NAND U3343 ( .A(N928), .B(xregN_1), .Z(n2230) );
  NAND U3344 ( .A(n2232), .B(n2233), .Z(z2[923]) );
  NANDN U3345 ( .A(xregN_1), .B(zin[922]), .Z(n2233) );
  NAND U3346 ( .A(N927), .B(xregN_1), .Z(n2232) );
  NAND U3347 ( .A(n2234), .B(n2235), .Z(z2[922]) );
  NANDN U3348 ( .A(xregN_1), .B(zin[921]), .Z(n2235) );
  NAND U3349 ( .A(N926), .B(xregN_1), .Z(n2234) );
  NAND U3350 ( .A(n2236), .B(n2237), .Z(z2[921]) );
  NANDN U3351 ( .A(xregN_1), .B(zin[920]), .Z(n2237) );
  NAND U3352 ( .A(N925), .B(xregN_1), .Z(n2236) );
  NAND U3353 ( .A(n2238), .B(n2239), .Z(z2[920]) );
  NANDN U3354 ( .A(xregN_1), .B(zin[919]), .Z(n2239) );
  NAND U3355 ( .A(N924), .B(xregN_1), .Z(n2238) );
  NAND U3356 ( .A(n2240), .B(n2241), .Z(z2[91]) );
  NANDN U3357 ( .A(xregN_1), .B(zin[90]), .Z(n2241) );
  NAND U3358 ( .A(N95), .B(xregN_1), .Z(n2240) );
  NAND U3359 ( .A(n2242), .B(n2243), .Z(z2[919]) );
  NANDN U3360 ( .A(xregN_1), .B(zin[918]), .Z(n2243) );
  NAND U3361 ( .A(N923), .B(xregN_1), .Z(n2242) );
  NAND U3362 ( .A(n2244), .B(n2245), .Z(z2[918]) );
  NANDN U3363 ( .A(xregN_1), .B(zin[917]), .Z(n2245) );
  NAND U3364 ( .A(N922), .B(xregN_1), .Z(n2244) );
  NAND U3365 ( .A(n2246), .B(n2247), .Z(z2[917]) );
  NANDN U3366 ( .A(xregN_1), .B(zin[916]), .Z(n2247) );
  NAND U3367 ( .A(N921), .B(xregN_1), .Z(n2246) );
  NAND U3368 ( .A(n2248), .B(n2249), .Z(z2[916]) );
  NANDN U3369 ( .A(xregN_1), .B(zin[915]), .Z(n2249) );
  NAND U3370 ( .A(N920), .B(xregN_1), .Z(n2248) );
  NAND U3371 ( .A(n2250), .B(n2251), .Z(z2[915]) );
  NANDN U3372 ( .A(xregN_1), .B(zin[914]), .Z(n2251) );
  NAND U3373 ( .A(N919), .B(xregN_1), .Z(n2250) );
  NAND U3374 ( .A(n2252), .B(n2253), .Z(z2[914]) );
  NANDN U3375 ( .A(xregN_1), .B(zin[913]), .Z(n2253) );
  NAND U3376 ( .A(N918), .B(xregN_1), .Z(n2252) );
  NAND U3377 ( .A(n2254), .B(n2255), .Z(z2[913]) );
  NANDN U3378 ( .A(xregN_1), .B(zin[912]), .Z(n2255) );
  NAND U3379 ( .A(N917), .B(xregN_1), .Z(n2254) );
  NAND U3380 ( .A(n2256), .B(n2257), .Z(z2[912]) );
  NANDN U3381 ( .A(xregN_1), .B(zin[911]), .Z(n2257) );
  NAND U3382 ( .A(N916), .B(xregN_1), .Z(n2256) );
  NAND U3383 ( .A(n2258), .B(n2259), .Z(z2[911]) );
  NANDN U3384 ( .A(xregN_1), .B(zin[910]), .Z(n2259) );
  NAND U3385 ( .A(N915), .B(xregN_1), .Z(n2258) );
  NAND U3386 ( .A(n2260), .B(n2261), .Z(z2[910]) );
  NANDN U3387 ( .A(xregN_1), .B(zin[909]), .Z(n2261) );
  NAND U3388 ( .A(N914), .B(xregN_1), .Z(n2260) );
  NAND U3389 ( .A(n2262), .B(n2263), .Z(z2[90]) );
  NANDN U3390 ( .A(xregN_1), .B(zin[89]), .Z(n2263) );
  NAND U3391 ( .A(N94), .B(xregN_1), .Z(n2262) );
  NAND U3392 ( .A(n2264), .B(n2265), .Z(z2[909]) );
  NANDN U3393 ( .A(xregN_1), .B(zin[908]), .Z(n2265) );
  NAND U3394 ( .A(N913), .B(xregN_1), .Z(n2264) );
  NAND U3395 ( .A(n2266), .B(n2267), .Z(z2[908]) );
  NANDN U3396 ( .A(xregN_1), .B(zin[907]), .Z(n2267) );
  NAND U3397 ( .A(N912), .B(xregN_1), .Z(n2266) );
  NAND U3398 ( .A(n2268), .B(n2269), .Z(z2[907]) );
  NANDN U3399 ( .A(xregN_1), .B(zin[906]), .Z(n2269) );
  NAND U3400 ( .A(N911), .B(xregN_1), .Z(n2268) );
  NAND U3401 ( .A(n2270), .B(n2271), .Z(z2[906]) );
  NANDN U3402 ( .A(xregN_1), .B(zin[905]), .Z(n2271) );
  NAND U3403 ( .A(N910), .B(xregN_1), .Z(n2270) );
  NAND U3404 ( .A(n2272), .B(n2273), .Z(z2[905]) );
  NANDN U3405 ( .A(xregN_1), .B(zin[904]), .Z(n2273) );
  NAND U3406 ( .A(N909), .B(xregN_1), .Z(n2272) );
  NAND U3407 ( .A(n2274), .B(n2275), .Z(z2[904]) );
  NANDN U3408 ( .A(xregN_1), .B(zin[903]), .Z(n2275) );
  NAND U3409 ( .A(N908), .B(xregN_1), .Z(n2274) );
  NAND U3410 ( .A(n2276), .B(n2277), .Z(z2[903]) );
  NANDN U3411 ( .A(xregN_1), .B(zin[902]), .Z(n2277) );
  NAND U3412 ( .A(N907), .B(xregN_1), .Z(n2276) );
  NAND U3413 ( .A(n2278), .B(n2279), .Z(z2[902]) );
  NANDN U3414 ( .A(xregN_1), .B(zin[901]), .Z(n2279) );
  NAND U3415 ( .A(N906), .B(xregN_1), .Z(n2278) );
  NAND U3416 ( .A(n2280), .B(n2281), .Z(z2[901]) );
  NANDN U3417 ( .A(xregN_1), .B(zin[900]), .Z(n2281) );
  NAND U3418 ( .A(N905), .B(xregN_1), .Z(n2280) );
  NAND U3419 ( .A(n2282), .B(n2283), .Z(z2[900]) );
  NANDN U3420 ( .A(xregN_1), .B(zin[899]), .Z(n2283) );
  NAND U3421 ( .A(N904), .B(xregN_1), .Z(n2282) );
  NAND U3422 ( .A(n2284), .B(n2285), .Z(z2[8]) );
  NANDN U3423 ( .A(xregN_1), .B(zin[7]), .Z(n2285) );
  NAND U3424 ( .A(N12), .B(xregN_1), .Z(n2284) );
  NAND U3425 ( .A(n2286), .B(n2287), .Z(z2[89]) );
  NANDN U3426 ( .A(xregN_1), .B(zin[88]), .Z(n2287) );
  NAND U3427 ( .A(N93), .B(xregN_1), .Z(n2286) );
  NAND U3428 ( .A(n2288), .B(n2289), .Z(z2[899]) );
  NANDN U3429 ( .A(xregN_1), .B(zin[898]), .Z(n2289) );
  NAND U3430 ( .A(N903), .B(xregN_1), .Z(n2288) );
  NAND U3431 ( .A(n2290), .B(n2291), .Z(z2[898]) );
  NANDN U3432 ( .A(xregN_1), .B(zin[897]), .Z(n2291) );
  NAND U3433 ( .A(N902), .B(xregN_1), .Z(n2290) );
  NAND U3434 ( .A(n2292), .B(n2293), .Z(z2[897]) );
  NANDN U3435 ( .A(xregN_1), .B(zin[896]), .Z(n2293) );
  NAND U3436 ( .A(N901), .B(xregN_1), .Z(n2292) );
  NAND U3437 ( .A(n2294), .B(n2295), .Z(z2[896]) );
  NANDN U3438 ( .A(xregN_1), .B(zin[895]), .Z(n2295) );
  NAND U3439 ( .A(N900), .B(xregN_1), .Z(n2294) );
  NAND U3440 ( .A(n2296), .B(n2297), .Z(z2[895]) );
  NANDN U3441 ( .A(xregN_1), .B(zin[894]), .Z(n2297) );
  NAND U3442 ( .A(N899), .B(xregN_1), .Z(n2296) );
  NAND U3443 ( .A(n2298), .B(n2299), .Z(z2[894]) );
  NANDN U3444 ( .A(xregN_1), .B(zin[893]), .Z(n2299) );
  NAND U3445 ( .A(N898), .B(xregN_1), .Z(n2298) );
  NAND U3446 ( .A(n2300), .B(n2301), .Z(z2[893]) );
  NANDN U3447 ( .A(xregN_1), .B(zin[892]), .Z(n2301) );
  NAND U3448 ( .A(N897), .B(xregN_1), .Z(n2300) );
  NAND U3449 ( .A(n2302), .B(n2303), .Z(z2[892]) );
  NANDN U3450 ( .A(xregN_1), .B(zin[891]), .Z(n2303) );
  NAND U3451 ( .A(N896), .B(xregN_1), .Z(n2302) );
  NAND U3452 ( .A(n2304), .B(n2305), .Z(z2[891]) );
  NANDN U3453 ( .A(xregN_1), .B(zin[890]), .Z(n2305) );
  NAND U3454 ( .A(N895), .B(xregN_1), .Z(n2304) );
  NAND U3455 ( .A(n2306), .B(n2307), .Z(z2[890]) );
  NANDN U3456 ( .A(xregN_1), .B(zin[889]), .Z(n2307) );
  NAND U3457 ( .A(N894), .B(xregN_1), .Z(n2306) );
  NAND U3458 ( .A(n2308), .B(n2309), .Z(z2[88]) );
  NANDN U3459 ( .A(xregN_1), .B(zin[87]), .Z(n2309) );
  NAND U3460 ( .A(N92), .B(xregN_1), .Z(n2308) );
  NAND U3461 ( .A(n2310), .B(n2311), .Z(z2[889]) );
  NANDN U3462 ( .A(xregN_1), .B(zin[888]), .Z(n2311) );
  NAND U3463 ( .A(N893), .B(xregN_1), .Z(n2310) );
  NAND U3464 ( .A(n2312), .B(n2313), .Z(z2[888]) );
  NANDN U3465 ( .A(xregN_1), .B(zin[887]), .Z(n2313) );
  NAND U3466 ( .A(N892), .B(xregN_1), .Z(n2312) );
  NAND U3467 ( .A(n2314), .B(n2315), .Z(z2[887]) );
  NANDN U3468 ( .A(xregN_1), .B(zin[886]), .Z(n2315) );
  NAND U3469 ( .A(N891), .B(xregN_1), .Z(n2314) );
  NAND U3470 ( .A(n2316), .B(n2317), .Z(z2[886]) );
  NANDN U3471 ( .A(xregN_1), .B(zin[885]), .Z(n2317) );
  NAND U3472 ( .A(N890), .B(xregN_1), .Z(n2316) );
  NAND U3473 ( .A(n2318), .B(n2319), .Z(z2[885]) );
  NANDN U3474 ( .A(xregN_1), .B(zin[884]), .Z(n2319) );
  NAND U3475 ( .A(N889), .B(xregN_1), .Z(n2318) );
  NAND U3476 ( .A(n2320), .B(n2321), .Z(z2[884]) );
  NANDN U3477 ( .A(xregN_1), .B(zin[883]), .Z(n2321) );
  NAND U3478 ( .A(N888), .B(xregN_1), .Z(n2320) );
  NAND U3479 ( .A(n2322), .B(n2323), .Z(z2[883]) );
  NANDN U3480 ( .A(xregN_1), .B(zin[882]), .Z(n2323) );
  NAND U3481 ( .A(N887), .B(xregN_1), .Z(n2322) );
  NAND U3482 ( .A(n2324), .B(n2325), .Z(z2[882]) );
  NANDN U3483 ( .A(xregN_1), .B(zin[881]), .Z(n2325) );
  NAND U3484 ( .A(N886), .B(xregN_1), .Z(n2324) );
  NAND U3485 ( .A(n2326), .B(n2327), .Z(z2[881]) );
  NANDN U3486 ( .A(xregN_1), .B(zin[880]), .Z(n2327) );
  NAND U3487 ( .A(N885), .B(xregN_1), .Z(n2326) );
  NAND U3488 ( .A(n2328), .B(n2329), .Z(z2[880]) );
  NANDN U3489 ( .A(xregN_1), .B(zin[879]), .Z(n2329) );
  NAND U3490 ( .A(N884), .B(xregN_1), .Z(n2328) );
  NAND U3491 ( .A(n2330), .B(n2331), .Z(z2[87]) );
  NANDN U3492 ( .A(xregN_1), .B(zin[86]), .Z(n2331) );
  NAND U3493 ( .A(N91), .B(xregN_1), .Z(n2330) );
  NAND U3494 ( .A(n2332), .B(n2333), .Z(z2[879]) );
  NANDN U3495 ( .A(xregN_1), .B(zin[878]), .Z(n2333) );
  NAND U3496 ( .A(N883), .B(xregN_1), .Z(n2332) );
  NAND U3497 ( .A(n2334), .B(n2335), .Z(z2[878]) );
  NANDN U3498 ( .A(xregN_1), .B(zin[877]), .Z(n2335) );
  NAND U3499 ( .A(N882), .B(xregN_1), .Z(n2334) );
  NAND U3500 ( .A(n2336), .B(n2337), .Z(z2[877]) );
  NANDN U3501 ( .A(xregN_1), .B(zin[876]), .Z(n2337) );
  NAND U3502 ( .A(N881), .B(xregN_1), .Z(n2336) );
  NAND U3503 ( .A(n2338), .B(n2339), .Z(z2[876]) );
  NANDN U3504 ( .A(xregN_1), .B(zin[875]), .Z(n2339) );
  NAND U3505 ( .A(N880), .B(xregN_1), .Z(n2338) );
  NAND U3506 ( .A(n2340), .B(n2341), .Z(z2[875]) );
  NANDN U3507 ( .A(xregN_1), .B(zin[874]), .Z(n2341) );
  NAND U3508 ( .A(N879), .B(xregN_1), .Z(n2340) );
  NAND U3509 ( .A(n2342), .B(n2343), .Z(z2[874]) );
  NANDN U3510 ( .A(xregN_1), .B(zin[873]), .Z(n2343) );
  NAND U3511 ( .A(N878), .B(xregN_1), .Z(n2342) );
  NAND U3512 ( .A(n2344), .B(n2345), .Z(z2[873]) );
  NANDN U3513 ( .A(xregN_1), .B(zin[872]), .Z(n2345) );
  NAND U3514 ( .A(N877), .B(xregN_1), .Z(n2344) );
  NAND U3515 ( .A(n2346), .B(n2347), .Z(z2[872]) );
  NANDN U3516 ( .A(xregN_1), .B(zin[871]), .Z(n2347) );
  NAND U3517 ( .A(N876), .B(xregN_1), .Z(n2346) );
  NAND U3518 ( .A(n2348), .B(n2349), .Z(z2[871]) );
  NANDN U3519 ( .A(xregN_1), .B(zin[870]), .Z(n2349) );
  NAND U3520 ( .A(N875), .B(xregN_1), .Z(n2348) );
  NAND U3521 ( .A(n2350), .B(n2351), .Z(z2[870]) );
  NANDN U3522 ( .A(xregN_1), .B(zin[869]), .Z(n2351) );
  NAND U3523 ( .A(N874), .B(xregN_1), .Z(n2350) );
  NAND U3524 ( .A(n2352), .B(n2353), .Z(z2[86]) );
  NANDN U3525 ( .A(xregN_1), .B(zin[85]), .Z(n2353) );
  NAND U3526 ( .A(N90), .B(xregN_1), .Z(n2352) );
  NAND U3527 ( .A(n2354), .B(n2355), .Z(z2[869]) );
  NANDN U3528 ( .A(xregN_1), .B(zin[868]), .Z(n2355) );
  NAND U3529 ( .A(N873), .B(xregN_1), .Z(n2354) );
  NAND U3530 ( .A(n2356), .B(n2357), .Z(z2[868]) );
  NANDN U3531 ( .A(xregN_1), .B(zin[867]), .Z(n2357) );
  NAND U3532 ( .A(N872), .B(xregN_1), .Z(n2356) );
  NAND U3533 ( .A(n2358), .B(n2359), .Z(z2[867]) );
  NANDN U3534 ( .A(xregN_1), .B(zin[866]), .Z(n2359) );
  NAND U3535 ( .A(N871), .B(xregN_1), .Z(n2358) );
  NAND U3536 ( .A(n2360), .B(n2361), .Z(z2[866]) );
  NANDN U3537 ( .A(xregN_1), .B(zin[865]), .Z(n2361) );
  NAND U3538 ( .A(N870), .B(xregN_1), .Z(n2360) );
  NAND U3539 ( .A(n2362), .B(n2363), .Z(z2[865]) );
  NANDN U3540 ( .A(xregN_1), .B(zin[864]), .Z(n2363) );
  NAND U3541 ( .A(N869), .B(xregN_1), .Z(n2362) );
  NAND U3542 ( .A(n2364), .B(n2365), .Z(z2[864]) );
  NANDN U3543 ( .A(xregN_1), .B(zin[863]), .Z(n2365) );
  NAND U3544 ( .A(N868), .B(xregN_1), .Z(n2364) );
  NAND U3545 ( .A(n2366), .B(n2367), .Z(z2[863]) );
  NANDN U3546 ( .A(xregN_1), .B(zin[862]), .Z(n2367) );
  NAND U3547 ( .A(N867), .B(xregN_1), .Z(n2366) );
  NAND U3548 ( .A(n2368), .B(n2369), .Z(z2[862]) );
  NANDN U3549 ( .A(xregN_1), .B(zin[861]), .Z(n2369) );
  NAND U3550 ( .A(N866), .B(xregN_1), .Z(n2368) );
  NAND U3551 ( .A(n2370), .B(n2371), .Z(z2[861]) );
  NANDN U3552 ( .A(xregN_1), .B(zin[860]), .Z(n2371) );
  NAND U3553 ( .A(N865), .B(xregN_1), .Z(n2370) );
  NAND U3554 ( .A(n2372), .B(n2373), .Z(z2[860]) );
  NANDN U3555 ( .A(xregN_1), .B(zin[859]), .Z(n2373) );
  NAND U3556 ( .A(N864), .B(xregN_1), .Z(n2372) );
  NAND U3557 ( .A(n2374), .B(n2375), .Z(z2[85]) );
  NANDN U3558 ( .A(xregN_1), .B(zin[84]), .Z(n2375) );
  NAND U3559 ( .A(N89), .B(xregN_1), .Z(n2374) );
  NAND U3560 ( .A(n2376), .B(n2377), .Z(z2[859]) );
  NANDN U3561 ( .A(xregN_1), .B(zin[858]), .Z(n2377) );
  NAND U3562 ( .A(N863), .B(xregN_1), .Z(n2376) );
  NAND U3563 ( .A(n2378), .B(n2379), .Z(z2[858]) );
  NANDN U3564 ( .A(xregN_1), .B(zin[857]), .Z(n2379) );
  NAND U3565 ( .A(N862), .B(xregN_1), .Z(n2378) );
  NAND U3566 ( .A(n2380), .B(n2381), .Z(z2[857]) );
  NANDN U3567 ( .A(xregN_1), .B(zin[856]), .Z(n2381) );
  NAND U3568 ( .A(N861), .B(xregN_1), .Z(n2380) );
  NAND U3569 ( .A(n2382), .B(n2383), .Z(z2[856]) );
  NANDN U3570 ( .A(xregN_1), .B(zin[855]), .Z(n2383) );
  NAND U3571 ( .A(N860), .B(xregN_1), .Z(n2382) );
  NAND U3572 ( .A(n2384), .B(n2385), .Z(z2[855]) );
  NANDN U3573 ( .A(xregN_1), .B(zin[854]), .Z(n2385) );
  NAND U3574 ( .A(N859), .B(xregN_1), .Z(n2384) );
  NAND U3575 ( .A(n2386), .B(n2387), .Z(z2[854]) );
  NANDN U3576 ( .A(xregN_1), .B(zin[853]), .Z(n2387) );
  NAND U3577 ( .A(N858), .B(xregN_1), .Z(n2386) );
  NAND U3578 ( .A(n2388), .B(n2389), .Z(z2[853]) );
  NANDN U3579 ( .A(xregN_1), .B(zin[852]), .Z(n2389) );
  NAND U3580 ( .A(N857), .B(xregN_1), .Z(n2388) );
  NAND U3581 ( .A(n2390), .B(n2391), .Z(z2[852]) );
  NANDN U3582 ( .A(xregN_1), .B(zin[851]), .Z(n2391) );
  NAND U3583 ( .A(N856), .B(xregN_1), .Z(n2390) );
  NAND U3584 ( .A(n2392), .B(n2393), .Z(z2[851]) );
  NANDN U3585 ( .A(xregN_1), .B(zin[850]), .Z(n2393) );
  NAND U3586 ( .A(N855), .B(xregN_1), .Z(n2392) );
  NAND U3587 ( .A(n2394), .B(n2395), .Z(z2[850]) );
  NANDN U3588 ( .A(xregN_1), .B(zin[849]), .Z(n2395) );
  NAND U3589 ( .A(N854), .B(xregN_1), .Z(n2394) );
  NAND U3590 ( .A(n2396), .B(n2397), .Z(z2[84]) );
  NANDN U3591 ( .A(xregN_1), .B(zin[83]), .Z(n2397) );
  NAND U3592 ( .A(N88), .B(xregN_1), .Z(n2396) );
  NAND U3593 ( .A(n2398), .B(n2399), .Z(z2[849]) );
  NANDN U3594 ( .A(xregN_1), .B(zin[848]), .Z(n2399) );
  NAND U3595 ( .A(N853), .B(xregN_1), .Z(n2398) );
  NAND U3596 ( .A(n2400), .B(n2401), .Z(z2[848]) );
  NANDN U3597 ( .A(xregN_1), .B(zin[847]), .Z(n2401) );
  NAND U3598 ( .A(N852), .B(xregN_1), .Z(n2400) );
  NAND U3599 ( .A(n2402), .B(n2403), .Z(z2[847]) );
  NANDN U3600 ( .A(xregN_1), .B(zin[846]), .Z(n2403) );
  NAND U3601 ( .A(N851), .B(xregN_1), .Z(n2402) );
  NAND U3602 ( .A(n2404), .B(n2405), .Z(z2[846]) );
  NANDN U3603 ( .A(xregN_1), .B(zin[845]), .Z(n2405) );
  NAND U3604 ( .A(N850), .B(xregN_1), .Z(n2404) );
  NAND U3605 ( .A(n2406), .B(n2407), .Z(z2[845]) );
  NANDN U3606 ( .A(xregN_1), .B(zin[844]), .Z(n2407) );
  NAND U3607 ( .A(N849), .B(xregN_1), .Z(n2406) );
  NAND U3608 ( .A(n2408), .B(n2409), .Z(z2[844]) );
  NANDN U3609 ( .A(xregN_1), .B(zin[843]), .Z(n2409) );
  NAND U3610 ( .A(N848), .B(xregN_1), .Z(n2408) );
  NAND U3611 ( .A(n2410), .B(n2411), .Z(z2[843]) );
  NANDN U3612 ( .A(xregN_1), .B(zin[842]), .Z(n2411) );
  NAND U3613 ( .A(N847), .B(xregN_1), .Z(n2410) );
  NAND U3614 ( .A(n2412), .B(n2413), .Z(z2[842]) );
  NANDN U3615 ( .A(xregN_1), .B(zin[841]), .Z(n2413) );
  NAND U3616 ( .A(N846), .B(xregN_1), .Z(n2412) );
  NAND U3617 ( .A(n2414), .B(n2415), .Z(z2[841]) );
  NANDN U3618 ( .A(xregN_1), .B(zin[840]), .Z(n2415) );
  NAND U3619 ( .A(N845), .B(xregN_1), .Z(n2414) );
  NAND U3620 ( .A(n2416), .B(n2417), .Z(z2[840]) );
  NANDN U3621 ( .A(xregN_1), .B(zin[839]), .Z(n2417) );
  NAND U3622 ( .A(N844), .B(xregN_1), .Z(n2416) );
  NAND U3623 ( .A(n2418), .B(n2419), .Z(z2[83]) );
  NANDN U3624 ( .A(xregN_1), .B(zin[82]), .Z(n2419) );
  NAND U3625 ( .A(N87), .B(xregN_1), .Z(n2418) );
  NAND U3626 ( .A(n2420), .B(n2421), .Z(z2[839]) );
  NANDN U3627 ( .A(xregN_1), .B(zin[838]), .Z(n2421) );
  NAND U3628 ( .A(N843), .B(xregN_1), .Z(n2420) );
  NAND U3629 ( .A(n2422), .B(n2423), .Z(z2[838]) );
  NANDN U3630 ( .A(xregN_1), .B(zin[837]), .Z(n2423) );
  NAND U3631 ( .A(N842), .B(xregN_1), .Z(n2422) );
  NAND U3632 ( .A(n2424), .B(n2425), .Z(z2[837]) );
  NANDN U3633 ( .A(xregN_1), .B(zin[836]), .Z(n2425) );
  NAND U3634 ( .A(N841), .B(xregN_1), .Z(n2424) );
  NAND U3635 ( .A(n2426), .B(n2427), .Z(z2[836]) );
  NANDN U3636 ( .A(xregN_1), .B(zin[835]), .Z(n2427) );
  NAND U3637 ( .A(N840), .B(xregN_1), .Z(n2426) );
  NAND U3638 ( .A(n2428), .B(n2429), .Z(z2[835]) );
  NANDN U3639 ( .A(xregN_1), .B(zin[834]), .Z(n2429) );
  NAND U3640 ( .A(N839), .B(xregN_1), .Z(n2428) );
  NAND U3641 ( .A(n2430), .B(n2431), .Z(z2[834]) );
  NANDN U3642 ( .A(xregN_1), .B(zin[833]), .Z(n2431) );
  NAND U3643 ( .A(N838), .B(xregN_1), .Z(n2430) );
  NAND U3644 ( .A(n2432), .B(n2433), .Z(z2[833]) );
  NANDN U3645 ( .A(xregN_1), .B(zin[832]), .Z(n2433) );
  NAND U3646 ( .A(N837), .B(xregN_1), .Z(n2432) );
  NAND U3647 ( .A(n2434), .B(n2435), .Z(z2[832]) );
  NANDN U3648 ( .A(xregN_1), .B(zin[831]), .Z(n2435) );
  NAND U3649 ( .A(N836), .B(xregN_1), .Z(n2434) );
  NAND U3650 ( .A(n2436), .B(n2437), .Z(z2[831]) );
  NANDN U3651 ( .A(xregN_1), .B(zin[830]), .Z(n2437) );
  NAND U3652 ( .A(N835), .B(xregN_1), .Z(n2436) );
  NAND U3653 ( .A(n2438), .B(n2439), .Z(z2[830]) );
  NANDN U3654 ( .A(xregN_1), .B(zin[829]), .Z(n2439) );
  NAND U3655 ( .A(N834), .B(xregN_1), .Z(n2438) );
  NAND U3656 ( .A(n2440), .B(n2441), .Z(z2[82]) );
  NANDN U3657 ( .A(xregN_1), .B(zin[81]), .Z(n2441) );
  NAND U3658 ( .A(N86), .B(xregN_1), .Z(n2440) );
  NAND U3659 ( .A(n2442), .B(n2443), .Z(z2[829]) );
  NANDN U3660 ( .A(xregN_1), .B(zin[828]), .Z(n2443) );
  NAND U3661 ( .A(N833), .B(xregN_1), .Z(n2442) );
  NAND U3662 ( .A(n2444), .B(n2445), .Z(z2[828]) );
  NANDN U3663 ( .A(xregN_1), .B(zin[827]), .Z(n2445) );
  NAND U3664 ( .A(N832), .B(xregN_1), .Z(n2444) );
  NAND U3665 ( .A(n2446), .B(n2447), .Z(z2[827]) );
  NANDN U3666 ( .A(xregN_1), .B(zin[826]), .Z(n2447) );
  NAND U3667 ( .A(N831), .B(xregN_1), .Z(n2446) );
  NAND U3668 ( .A(n2448), .B(n2449), .Z(z2[826]) );
  NANDN U3669 ( .A(xregN_1), .B(zin[825]), .Z(n2449) );
  NAND U3670 ( .A(N830), .B(xregN_1), .Z(n2448) );
  NAND U3671 ( .A(n2450), .B(n2451), .Z(z2[825]) );
  NANDN U3672 ( .A(xregN_1), .B(zin[824]), .Z(n2451) );
  NAND U3673 ( .A(N829), .B(xregN_1), .Z(n2450) );
  NAND U3674 ( .A(n2452), .B(n2453), .Z(z2[824]) );
  NANDN U3675 ( .A(xregN_1), .B(zin[823]), .Z(n2453) );
  NAND U3676 ( .A(N828), .B(xregN_1), .Z(n2452) );
  NAND U3677 ( .A(n2454), .B(n2455), .Z(z2[823]) );
  NANDN U3678 ( .A(xregN_1), .B(zin[822]), .Z(n2455) );
  NAND U3679 ( .A(N827), .B(xregN_1), .Z(n2454) );
  NAND U3680 ( .A(n2456), .B(n2457), .Z(z2[822]) );
  NANDN U3681 ( .A(xregN_1), .B(zin[821]), .Z(n2457) );
  NAND U3682 ( .A(N826), .B(xregN_1), .Z(n2456) );
  NAND U3683 ( .A(n2458), .B(n2459), .Z(z2[821]) );
  NANDN U3684 ( .A(xregN_1), .B(zin[820]), .Z(n2459) );
  NAND U3685 ( .A(N825), .B(xregN_1), .Z(n2458) );
  NAND U3686 ( .A(n2460), .B(n2461), .Z(z2[820]) );
  NANDN U3687 ( .A(xregN_1), .B(zin[819]), .Z(n2461) );
  NAND U3688 ( .A(N824), .B(xregN_1), .Z(n2460) );
  NAND U3689 ( .A(n2462), .B(n2463), .Z(z2[81]) );
  NANDN U3690 ( .A(xregN_1), .B(zin[80]), .Z(n2463) );
  NAND U3691 ( .A(N85), .B(xregN_1), .Z(n2462) );
  NAND U3692 ( .A(n2464), .B(n2465), .Z(z2[819]) );
  NANDN U3693 ( .A(xregN_1), .B(zin[818]), .Z(n2465) );
  NAND U3694 ( .A(N823), .B(xregN_1), .Z(n2464) );
  NAND U3695 ( .A(n2466), .B(n2467), .Z(z2[818]) );
  NANDN U3696 ( .A(xregN_1), .B(zin[817]), .Z(n2467) );
  NAND U3697 ( .A(N822), .B(xregN_1), .Z(n2466) );
  NAND U3698 ( .A(n2468), .B(n2469), .Z(z2[817]) );
  NANDN U3699 ( .A(xregN_1), .B(zin[816]), .Z(n2469) );
  NAND U3700 ( .A(N821), .B(xregN_1), .Z(n2468) );
  NAND U3701 ( .A(n2470), .B(n2471), .Z(z2[816]) );
  NANDN U3702 ( .A(xregN_1), .B(zin[815]), .Z(n2471) );
  NAND U3703 ( .A(N820), .B(xregN_1), .Z(n2470) );
  NAND U3704 ( .A(n2472), .B(n2473), .Z(z2[815]) );
  NANDN U3705 ( .A(xregN_1), .B(zin[814]), .Z(n2473) );
  NAND U3706 ( .A(N819), .B(xregN_1), .Z(n2472) );
  NAND U3707 ( .A(n2474), .B(n2475), .Z(z2[814]) );
  NANDN U3708 ( .A(xregN_1), .B(zin[813]), .Z(n2475) );
  NAND U3709 ( .A(N818), .B(xregN_1), .Z(n2474) );
  NAND U3710 ( .A(n2476), .B(n2477), .Z(z2[813]) );
  NANDN U3711 ( .A(xregN_1), .B(zin[812]), .Z(n2477) );
  NAND U3712 ( .A(N817), .B(xregN_1), .Z(n2476) );
  NAND U3713 ( .A(n2478), .B(n2479), .Z(z2[812]) );
  NANDN U3714 ( .A(xregN_1), .B(zin[811]), .Z(n2479) );
  NAND U3715 ( .A(N816), .B(xregN_1), .Z(n2478) );
  NAND U3716 ( .A(n2480), .B(n2481), .Z(z2[811]) );
  NANDN U3717 ( .A(xregN_1), .B(zin[810]), .Z(n2481) );
  NAND U3718 ( .A(N815), .B(xregN_1), .Z(n2480) );
  NAND U3719 ( .A(n2482), .B(n2483), .Z(z2[810]) );
  NANDN U3720 ( .A(xregN_1), .B(zin[809]), .Z(n2483) );
  NAND U3721 ( .A(N814), .B(xregN_1), .Z(n2482) );
  NAND U3722 ( .A(n2484), .B(n2485), .Z(z2[80]) );
  NANDN U3723 ( .A(xregN_1), .B(zin[79]), .Z(n2485) );
  NAND U3724 ( .A(N84), .B(xregN_1), .Z(n2484) );
  NAND U3725 ( .A(n2486), .B(n2487), .Z(z2[809]) );
  NANDN U3726 ( .A(xregN_1), .B(zin[808]), .Z(n2487) );
  NAND U3727 ( .A(N813), .B(xregN_1), .Z(n2486) );
  NAND U3728 ( .A(n2488), .B(n2489), .Z(z2[808]) );
  NANDN U3729 ( .A(xregN_1), .B(zin[807]), .Z(n2489) );
  NAND U3730 ( .A(N812), .B(xregN_1), .Z(n2488) );
  NAND U3731 ( .A(n2490), .B(n2491), .Z(z2[807]) );
  NANDN U3732 ( .A(xregN_1), .B(zin[806]), .Z(n2491) );
  NAND U3733 ( .A(N811), .B(xregN_1), .Z(n2490) );
  NAND U3734 ( .A(n2492), .B(n2493), .Z(z2[806]) );
  NANDN U3735 ( .A(xregN_1), .B(zin[805]), .Z(n2493) );
  NAND U3736 ( .A(N810), .B(xregN_1), .Z(n2492) );
  NAND U3737 ( .A(n2494), .B(n2495), .Z(z2[805]) );
  NANDN U3738 ( .A(xregN_1), .B(zin[804]), .Z(n2495) );
  NAND U3739 ( .A(N809), .B(xregN_1), .Z(n2494) );
  NAND U3740 ( .A(n2496), .B(n2497), .Z(z2[804]) );
  NANDN U3741 ( .A(xregN_1), .B(zin[803]), .Z(n2497) );
  NAND U3742 ( .A(N808), .B(xregN_1), .Z(n2496) );
  NAND U3743 ( .A(n2498), .B(n2499), .Z(z2[803]) );
  NANDN U3744 ( .A(xregN_1), .B(zin[802]), .Z(n2499) );
  NAND U3745 ( .A(N807), .B(xregN_1), .Z(n2498) );
  NAND U3746 ( .A(n2500), .B(n2501), .Z(z2[802]) );
  NANDN U3747 ( .A(xregN_1), .B(zin[801]), .Z(n2501) );
  NAND U3748 ( .A(N806), .B(xregN_1), .Z(n2500) );
  NAND U3749 ( .A(n2502), .B(n2503), .Z(z2[801]) );
  NANDN U3750 ( .A(xregN_1), .B(zin[800]), .Z(n2503) );
  NAND U3751 ( .A(N805), .B(xregN_1), .Z(n2502) );
  NAND U3752 ( .A(n2504), .B(n2505), .Z(z2[800]) );
  NANDN U3753 ( .A(xregN_1), .B(zin[799]), .Z(n2505) );
  NAND U3754 ( .A(N804), .B(xregN_1), .Z(n2504) );
  NAND U3755 ( .A(n2506), .B(n2507), .Z(z2[7]) );
  NANDN U3756 ( .A(xregN_1), .B(zin[6]), .Z(n2507) );
  NAND U3757 ( .A(N11), .B(xregN_1), .Z(n2506) );
  NAND U3758 ( .A(n2508), .B(n2509), .Z(z2[79]) );
  NANDN U3759 ( .A(xregN_1), .B(zin[78]), .Z(n2509) );
  NAND U3760 ( .A(N83), .B(xregN_1), .Z(n2508) );
  NAND U3761 ( .A(n2510), .B(n2511), .Z(z2[799]) );
  NANDN U3762 ( .A(xregN_1), .B(zin[798]), .Z(n2511) );
  NAND U3763 ( .A(N803), .B(xregN_1), .Z(n2510) );
  NAND U3764 ( .A(n2512), .B(n2513), .Z(z2[798]) );
  NANDN U3765 ( .A(xregN_1), .B(zin[797]), .Z(n2513) );
  NAND U3766 ( .A(N802), .B(xregN_1), .Z(n2512) );
  NAND U3767 ( .A(n2514), .B(n2515), .Z(z2[797]) );
  NANDN U3768 ( .A(xregN_1), .B(zin[796]), .Z(n2515) );
  NAND U3769 ( .A(N801), .B(xregN_1), .Z(n2514) );
  NAND U3770 ( .A(n2516), .B(n2517), .Z(z2[796]) );
  NANDN U3771 ( .A(xregN_1), .B(zin[795]), .Z(n2517) );
  NAND U3772 ( .A(N800), .B(xregN_1), .Z(n2516) );
  NAND U3773 ( .A(n2518), .B(n2519), .Z(z2[795]) );
  NANDN U3774 ( .A(xregN_1), .B(zin[794]), .Z(n2519) );
  NAND U3775 ( .A(N799), .B(xregN_1), .Z(n2518) );
  NAND U3776 ( .A(n2520), .B(n2521), .Z(z2[794]) );
  NANDN U3777 ( .A(xregN_1), .B(zin[793]), .Z(n2521) );
  NAND U3778 ( .A(N798), .B(xregN_1), .Z(n2520) );
  NAND U3779 ( .A(n2522), .B(n2523), .Z(z2[793]) );
  NANDN U3780 ( .A(xregN_1), .B(zin[792]), .Z(n2523) );
  NAND U3781 ( .A(N797), .B(xregN_1), .Z(n2522) );
  NAND U3782 ( .A(n2524), .B(n2525), .Z(z2[792]) );
  NANDN U3783 ( .A(xregN_1), .B(zin[791]), .Z(n2525) );
  NAND U3784 ( .A(N796), .B(xregN_1), .Z(n2524) );
  NAND U3785 ( .A(n2526), .B(n2527), .Z(z2[791]) );
  NANDN U3786 ( .A(xregN_1), .B(zin[790]), .Z(n2527) );
  NAND U3787 ( .A(N795), .B(xregN_1), .Z(n2526) );
  NAND U3788 ( .A(n2528), .B(n2529), .Z(z2[790]) );
  NANDN U3789 ( .A(xregN_1), .B(zin[789]), .Z(n2529) );
  NAND U3790 ( .A(N794), .B(xregN_1), .Z(n2528) );
  NAND U3791 ( .A(n2530), .B(n2531), .Z(z2[78]) );
  NANDN U3792 ( .A(xregN_1), .B(zin[77]), .Z(n2531) );
  NAND U3793 ( .A(N82), .B(xregN_1), .Z(n2530) );
  NAND U3794 ( .A(n2532), .B(n2533), .Z(z2[789]) );
  NANDN U3795 ( .A(xregN_1), .B(zin[788]), .Z(n2533) );
  NAND U3796 ( .A(N793), .B(xregN_1), .Z(n2532) );
  NAND U3797 ( .A(n2534), .B(n2535), .Z(z2[788]) );
  NANDN U3798 ( .A(xregN_1), .B(zin[787]), .Z(n2535) );
  NAND U3799 ( .A(N792), .B(xregN_1), .Z(n2534) );
  NAND U3800 ( .A(n2536), .B(n2537), .Z(z2[787]) );
  NANDN U3801 ( .A(xregN_1), .B(zin[786]), .Z(n2537) );
  NAND U3802 ( .A(N791), .B(xregN_1), .Z(n2536) );
  NAND U3803 ( .A(n2538), .B(n2539), .Z(z2[786]) );
  NANDN U3804 ( .A(xregN_1), .B(zin[785]), .Z(n2539) );
  NAND U3805 ( .A(N790), .B(xregN_1), .Z(n2538) );
  NAND U3806 ( .A(n2540), .B(n2541), .Z(z2[785]) );
  NANDN U3807 ( .A(xregN_1), .B(zin[784]), .Z(n2541) );
  NAND U3808 ( .A(N789), .B(xregN_1), .Z(n2540) );
  NAND U3809 ( .A(n2542), .B(n2543), .Z(z2[784]) );
  NANDN U3810 ( .A(xregN_1), .B(zin[783]), .Z(n2543) );
  NAND U3811 ( .A(N788), .B(xregN_1), .Z(n2542) );
  NAND U3812 ( .A(n2544), .B(n2545), .Z(z2[783]) );
  NANDN U3813 ( .A(xregN_1), .B(zin[782]), .Z(n2545) );
  NAND U3814 ( .A(N787), .B(xregN_1), .Z(n2544) );
  NAND U3815 ( .A(n2546), .B(n2547), .Z(z2[782]) );
  NANDN U3816 ( .A(xregN_1), .B(zin[781]), .Z(n2547) );
  NAND U3817 ( .A(N786), .B(xregN_1), .Z(n2546) );
  NAND U3818 ( .A(n2548), .B(n2549), .Z(z2[781]) );
  NANDN U3819 ( .A(xregN_1), .B(zin[780]), .Z(n2549) );
  NAND U3820 ( .A(N785), .B(xregN_1), .Z(n2548) );
  NAND U3821 ( .A(n2550), .B(n2551), .Z(z2[780]) );
  NANDN U3822 ( .A(xregN_1), .B(zin[779]), .Z(n2551) );
  NAND U3823 ( .A(N784), .B(xregN_1), .Z(n2550) );
  NAND U3824 ( .A(n2552), .B(n2553), .Z(z2[77]) );
  NANDN U3825 ( .A(xregN_1), .B(zin[76]), .Z(n2553) );
  NAND U3826 ( .A(N81), .B(xregN_1), .Z(n2552) );
  NAND U3827 ( .A(n2554), .B(n2555), .Z(z2[779]) );
  NANDN U3828 ( .A(xregN_1), .B(zin[778]), .Z(n2555) );
  NAND U3829 ( .A(N783), .B(xregN_1), .Z(n2554) );
  NAND U3830 ( .A(n2556), .B(n2557), .Z(z2[778]) );
  NANDN U3831 ( .A(xregN_1), .B(zin[777]), .Z(n2557) );
  NAND U3832 ( .A(N782), .B(xregN_1), .Z(n2556) );
  NAND U3833 ( .A(n2558), .B(n2559), .Z(z2[777]) );
  NANDN U3834 ( .A(xregN_1), .B(zin[776]), .Z(n2559) );
  NAND U3835 ( .A(N781), .B(xregN_1), .Z(n2558) );
  NAND U3836 ( .A(n2560), .B(n2561), .Z(z2[776]) );
  NANDN U3837 ( .A(xregN_1), .B(zin[775]), .Z(n2561) );
  NAND U3838 ( .A(N780), .B(xregN_1), .Z(n2560) );
  NAND U3839 ( .A(n2562), .B(n2563), .Z(z2[775]) );
  NANDN U3840 ( .A(xregN_1), .B(zin[774]), .Z(n2563) );
  NAND U3841 ( .A(N779), .B(xregN_1), .Z(n2562) );
  NAND U3842 ( .A(n2564), .B(n2565), .Z(z2[774]) );
  NANDN U3843 ( .A(xregN_1), .B(zin[773]), .Z(n2565) );
  NAND U3844 ( .A(N778), .B(xregN_1), .Z(n2564) );
  NAND U3845 ( .A(n2566), .B(n2567), .Z(z2[773]) );
  NANDN U3846 ( .A(xregN_1), .B(zin[772]), .Z(n2567) );
  NAND U3847 ( .A(N777), .B(xregN_1), .Z(n2566) );
  NAND U3848 ( .A(n2568), .B(n2569), .Z(z2[772]) );
  NANDN U3849 ( .A(xregN_1), .B(zin[771]), .Z(n2569) );
  NAND U3850 ( .A(N776), .B(xregN_1), .Z(n2568) );
  NAND U3851 ( .A(n2570), .B(n2571), .Z(z2[771]) );
  NANDN U3852 ( .A(xregN_1), .B(zin[770]), .Z(n2571) );
  NAND U3853 ( .A(N775), .B(xregN_1), .Z(n2570) );
  NAND U3854 ( .A(n2572), .B(n2573), .Z(z2[770]) );
  NANDN U3855 ( .A(xregN_1), .B(zin[769]), .Z(n2573) );
  NAND U3856 ( .A(N774), .B(xregN_1), .Z(n2572) );
  NAND U3857 ( .A(n2574), .B(n2575), .Z(z2[76]) );
  NANDN U3858 ( .A(xregN_1), .B(zin[75]), .Z(n2575) );
  NAND U3859 ( .A(N80), .B(xregN_1), .Z(n2574) );
  NAND U3860 ( .A(n2576), .B(n2577), .Z(z2[769]) );
  NANDN U3861 ( .A(xregN_1), .B(zin[768]), .Z(n2577) );
  NAND U3862 ( .A(N773), .B(xregN_1), .Z(n2576) );
  NAND U3863 ( .A(n2578), .B(n2579), .Z(z2[768]) );
  NANDN U3864 ( .A(xregN_1), .B(zin[767]), .Z(n2579) );
  NAND U3865 ( .A(N772), .B(xregN_1), .Z(n2578) );
  NAND U3866 ( .A(n2580), .B(n2581), .Z(z2[767]) );
  NANDN U3867 ( .A(xregN_1), .B(zin[766]), .Z(n2581) );
  NAND U3868 ( .A(N771), .B(xregN_1), .Z(n2580) );
  NAND U3869 ( .A(n2582), .B(n2583), .Z(z2[766]) );
  NANDN U3870 ( .A(xregN_1), .B(zin[765]), .Z(n2583) );
  NAND U3871 ( .A(N770), .B(xregN_1), .Z(n2582) );
  NAND U3872 ( .A(n2584), .B(n2585), .Z(z2[765]) );
  NANDN U3873 ( .A(xregN_1), .B(zin[764]), .Z(n2585) );
  NAND U3874 ( .A(N769), .B(xregN_1), .Z(n2584) );
  NAND U3875 ( .A(n2586), .B(n2587), .Z(z2[764]) );
  NANDN U3876 ( .A(xregN_1), .B(zin[763]), .Z(n2587) );
  NAND U3877 ( .A(N768), .B(xregN_1), .Z(n2586) );
  NAND U3878 ( .A(n2588), .B(n2589), .Z(z2[763]) );
  NANDN U3879 ( .A(xregN_1), .B(zin[762]), .Z(n2589) );
  NAND U3880 ( .A(N767), .B(xregN_1), .Z(n2588) );
  NAND U3881 ( .A(n2590), .B(n2591), .Z(z2[762]) );
  NANDN U3882 ( .A(xregN_1), .B(zin[761]), .Z(n2591) );
  NAND U3883 ( .A(N766), .B(xregN_1), .Z(n2590) );
  NAND U3884 ( .A(n2592), .B(n2593), .Z(z2[761]) );
  NANDN U3885 ( .A(xregN_1), .B(zin[760]), .Z(n2593) );
  NAND U3886 ( .A(N765), .B(xregN_1), .Z(n2592) );
  NAND U3887 ( .A(n2594), .B(n2595), .Z(z2[760]) );
  NANDN U3888 ( .A(xregN_1), .B(zin[759]), .Z(n2595) );
  NAND U3889 ( .A(N764), .B(xregN_1), .Z(n2594) );
  NAND U3890 ( .A(n2596), .B(n2597), .Z(z2[75]) );
  NANDN U3891 ( .A(xregN_1), .B(zin[74]), .Z(n2597) );
  NAND U3892 ( .A(N79), .B(xregN_1), .Z(n2596) );
  NAND U3893 ( .A(n2598), .B(n2599), .Z(z2[759]) );
  NANDN U3894 ( .A(xregN_1), .B(zin[758]), .Z(n2599) );
  NAND U3895 ( .A(N763), .B(xregN_1), .Z(n2598) );
  NAND U3896 ( .A(n2600), .B(n2601), .Z(z2[758]) );
  NANDN U3897 ( .A(xregN_1), .B(zin[757]), .Z(n2601) );
  NAND U3898 ( .A(N762), .B(xregN_1), .Z(n2600) );
  NAND U3899 ( .A(n2602), .B(n2603), .Z(z2[757]) );
  NANDN U3900 ( .A(xregN_1), .B(zin[756]), .Z(n2603) );
  NAND U3901 ( .A(N761), .B(xregN_1), .Z(n2602) );
  NAND U3902 ( .A(n2604), .B(n2605), .Z(z2[756]) );
  NANDN U3903 ( .A(xregN_1), .B(zin[755]), .Z(n2605) );
  NAND U3904 ( .A(N760), .B(xregN_1), .Z(n2604) );
  NAND U3905 ( .A(n2606), .B(n2607), .Z(z2[755]) );
  NANDN U3906 ( .A(xregN_1), .B(zin[754]), .Z(n2607) );
  NAND U3907 ( .A(N759), .B(xregN_1), .Z(n2606) );
  NAND U3908 ( .A(n2608), .B(n2609), .Z(z2[754]) );
  NANDN U3909 ( .A(xregN_1), .B(zin[753]), .Z(n2609) );
  NAND U3910 ( .A(N758), .B(xregN_1), .Z(n2608) );
  NAND U3911 ( .A(n2610), .B(n2611), .Z(z2[753]) );
  NANDN U3912 ( .A(xregN_1), .B(zin[752]), .Z(n2611) );
  NAND U3913 ( .A(N757), .B(xregN_1), .Z(n2610) );
  NAND U3914 ( .A(n2612), .B(n2613), .Z(z2[752]) );
  NANDN U3915 ( .A(xregN_1), .B(zin[751]), .Z(n2613) );
  NAND U3916 ( .A(N756), .B(xregN_1), .Z(n2612) );
  NAND U3917 ( .A(n2614), .B(n2615), .Z(z2[751]) );
  NANDN U3918 ( .A(xregN_1), .B(zin[750]), .Z(n2615) );
  NAND U3919 ( .A(N755), .B(xregN_1), .Z(n2614) );
  NAND U3920 ( .A(n2616), .B(n2617), .Z(z2[750]) );
  NANDN U3921 ( .A(xregN_1), .B(zin[749]), .Z(n2617) );
  NAND U3922 ( .A(N754), .B(xregN_1), .Z(n2616) );
  NAND U3923 ( .A(n2618), .B(n2619), .Z(z2[74]) );
  NANDN U3924 ( .A(xregN_1), .B(zin[73]), .Z(n2619) );
  NAND U3925 ( .A(N78), .B(xregN_1), .Z(n2618) );
  NAND U3926 ( .A(n2620), .B(n2621), .Z(z2[749]) );
  NANDN U3927 ( .A(xregN_1), .B(zin[748]), .Z(n2621) );
  NAND U3928 ( .A(N753), .B(xregN_1), .Z(n2620) );
  NAND U3929 ( .A(n2622), .B(n2623), .Z(z2[748]) );
  NANDN U3930 ( .A(xregN_1), .B(zin[747]), .Z(n2623) );
  NAND U3931 ( .A(N752), .B(xregN_1), .Z(n2622) );
  NAND U3932 ( .A(n2624), .B(n2625), .Z(z2[747]) );
  NANDN U3933 ( .A(xregN_1), .B(zin[746]), .Z(n2625) );
  NAND U3934 ( .A(N751), .B(xregN_1), .Z(n2624) );
  NAND U3935 ( .A(n2626), .B(n2627), .Z(z2[746]) );
  NANDN U3936 ( .A(xregN_1), .B(zin[745]), .Z(n2627) );
  NAND U3937 ( .A(N750), .B(xregN_1), .Z(n2626) );
  NAND U3938 ( .A(n2628), .B(n2629), .Z(z2[745]) );
  NANDN U3939 ( .A(xregN_1), .B(zin[744]), .Z(n2629) );
  NAND U3940 ( .A(N749), .B(xregN_1), .Z(n2628) );
  NAND U3941 ( .A(n2630), .B(n2631), .Z(z2[744]) );
  NANDN U3942 ( .A(xregN_1), .B(zin[743]), .Z(n2631) );
  NAND U3943 ( .A(N748), .B(xregN_1), .Z(n2630) );
  NAND U3944 ( .A(n2632), .B(n2633), .Z(z2[743]) );
  NANDN U3945 ( .A(xregN_1), .B(zin[742]), .Z(n2633) );
  NAND U3946 ( .A(N747), .B(xregN_1), .Z(n2632) );
  NAND U3947 ( .A(n2634), .B(n2635), .Z(z2[742]) );
  NANDN U3948 ( .A(xregN_1), .B(zin[741]), .Z(n2635) );
  NAND U3949 ( .A(N746), .B(xregN_1), .Z(n2634) );
  NAND U3950 ( .A(n2636), .B(n2637), .Z(z2[741]) );
  NANDN U3951 ( .A(xregN_1), .B(zin[740]), .Z(n2637) );
  NAND U3952 ( .A(N745), .B(xregN_1), .Z(n2636) );
  NAND U3953 ( .A(n2638), .B(n2639), .Z(z2[740]) );
  NANDN U3954 ( .A(xregN_1), .B(zin[739]), .Z(n2639) );
  NAND U3955 ( .A(N744), .B(xregN_1), .Z(n2638) );
  NAND U3956 ( .A(n2640), .B(n2641), .Z(z2[73]) );
  NANDN U3957 ( .A(xregN_1), .B(zin[72]), .Z(n2641) );
  NAND U3958 ( .A(N77), .B(xregN_1), .Z(n2640) );
  NAND U3959 ( .A(n2642), .B(n2643), .Z(z2[739]) );
  NANDN U3960 ( .A(xregN_1), .B(zin[738]), .Z(n2643) );
  NAND U3961 ( .A(N743), .B(xregN_1), .Z(n2642) );
  NAND U3962 ( .A(n2644), .B(n2645), .Z(z2[738]) );
  NANDN U3963 ( .A(xregN_1), .B(zin[737]), .Z(n2645) );
  NAND U3964 ( .A(N742), .B(xregN_1), .Z(n2644) );
  NAND U3965 ( .A(n2646), .B(n2647), .Z(z2[737]) );
  NANDN U3966 ( .A(xregN_1), .B(zin[736]), .Z(n2647) );
  NAND U3967 ( .A(N741), .B(xregN_1), .Z(n2646) );
  NAND U3968 ( .A(n2648), .B(n2649), .Z(z2[736]) );
  NANDN U3969 ( .A(xregN_1), .B(zin[735]), .Z(n2649) );
  NAND U3970 ( .A(N740), .B(xregN_1), .Z(n2648) );
  NAND U3971 ( .A(n2650), .B(n2651), .Z(z2[735]) );
  NANDN U3972 ( .A(xregN_1), .B(zin[734]), .Z(n2651) );
  NAND U3973 ( .A(N739), .B(xregN_1), .Z(n2650) );
  NAND U3974 ( .A(n2652), .B(n2653), .Z(z2[734]) );
  NANDN U3975 ( .A(xregN_1), .B(zin[733]), .Z(n2653) );
  NAND U3976 ( .A(N738), .B(xregN_1), .Z(n2652) );
  NAND U3977 ( .A(n2654), .B(n2655), .Z(z2[733]) );
  NANDN U3978 ( .A(xregN_1), .B(zin[732]), .Z(n2655) );
  NAND U3979 ( .A(N737), .B(xregN_1), .Z(n2654) );
  NAND U3980 ( .A(n2656), .B(n2657), .Z(z2[732]) );
  NANDN U3981 ( .A(xregN_1), .B(zin[731]), .Z(n2657) );
  NAND U3982 ( .A(N736), .B(xregN_1), .Z(n2656) );
  NAND U3983 ( .A(n2658), .B(n2659), .Z(z2[731]) );
  NANDN U3984 ( .A(xregN_1), .B(zin[730]), .Z(n2659) );
  NAND U3985 ( .A(N735), .B(xregN_1), .Z(n2658) );
  NAND U3986 ( .A(n2660), .B(n2661), .Z(z2[730]) );
  NANDN U3987 ( .A(xregN_1), .B(zin[729]), .Z(n2661) );
  NAND U3988 ( .A(N734), .B(xregN_1), .Z(n2660) );
  NAND U3989 ( .A(n2662), .B(n2663), .Z(z2[72]) );
  NANDN U3990 ( .A(xregN_1), .B(zin[71]), .Z(n2663) );
  NAND U3991 ( .A(N76), .B(xregN_1), .Z(n2662) );
  NAND U3992 ( .A(n2664), .B(n2665), .Z(z2[729]) );
  NANDN U3993 ( .A(xregN_1), .B(zin[728]), .Z(n2665) );
  NAND U3994 ( .A(N733), .B(xregN_1), .Z(n2664) );
  NAND U3995 ( .A(n2666), .B(n2667), .Z(z2[728]) );
  NANDN U3996 ( .A(xregN_1), .B(zin[727]), .Z(n2667) );
  NAND U3997 ( .A(N732), .B(xregN_1), .Z(n2666) );
  NAND U3998 ( .A(n2668), .B(n2669), .Z(z2[727]) );
  NANDN U3999 ( .A(xregN_1), .B(zin[726]), .Z(n2669) );
  NAND U4000 ( .A(N731), .B(xregN_1), .Z(n2668) );
  NAND U4001 ( .A(n2670), .B(n2671), .Z(z2[726]) );
  NANDN U4002 ( .A(xregN_1), .B(zin[725]), .Z(n2671) );
  NAND U4003 ( .A(N730), .B(xregN_1), .Z(n2670) );
  NAND U4004 ( .A(n2672), .B(n2673), .Z(z2[725]) );
  NANDN U4005 ( .A(xregN_1), .B(zin[724]), .Z(n2673) );
  NAND U4006 ( .A(N729), .B(xregN_1), .Z(n2672) );
  NAND U4007 ( .A(n2674), .B(n2675), .Z(z2[724]) );
  NANDN U4008 ( .A(xregN_1), .B(zin[723]), .Z(n2675) );
  NAND U4009 ( .A(N728), .B(xregN_1), .Z(n2674) );
  NAND U4010 ( .A(n2676), .B(n2677), .Z(z2[723]) );
  NANDN U4011 ( .A(xregN_1), .B(zin[722]), .Z(n2677) );
  NAND U4012 ( .A(N727), .B(xregN_1), .Z(n2676) );
  NAND U4013 ( .A(n2678), .B(n2679), .Z(z2[722]) );
  NANDN U4014 ( .A(xregN_1), .B(zin[721]), .Z(n2679) );
  NAND U4015 ( .A(N726), .B(xregN_1), .Z(n2678) );
  NAND U4016 ( .A(n2680), .B(n2681), .Z(z2[721]) );
  NANDN U4017 ( .A(xregN_1), .B(zin[720]), .Z(n2681) );
  NAND U4018 ( .A(N725), .B(xregN_1), .Z(n2680) );
  NAND U4019 ( .A(n2682), .B(n2683), .Z(z2[720]) );
  NANDN U4020 ( .A(xregN_1), .B(zin[719]), .Z(n2683) );
  NAND U4021 ( .A(N724), .B(xregN_1), .Z(n2682) );
  NAND U4022 ( .A(n2684), .B(n2685), .Z(z2[71]) );
  NANDN U4023 ( .A(xregN_1), .B(zin[70]), .Z(n2685) );
  NAND U4024 ( .A(N75), .B(xregN_1), .Z(n2684) );
  NAND U4025 ( .A(n2686), .B(n2687), .Z(z2[719]) );
  NANDN U4026 ( .A(xregN_1), .B(zin[718]), .Z(n2687) );
  NAND U4027 ( .A(N723), .B(xregN_1), .Z(n2686) );
  NAND U4028 ( .A(n2688), .B(n2689), .Z(z2[718]) );
  NANDN U4029 ( .A(xregN_1), .B(zin[717]), .Z(n2689) );
  NAND U4030 ( .A(N722), .B(xregN_1), .Z(n2688) );
  NAND U4031 ( .A(n2690), .B(n2691), .Z(z2[717]) );
  NANDN U4032 ( .A(xregN_1), .B(zin[716]), .Z(n2691) );
  NAND U4033 ( .A(N721), .B(xregN_1), .Z(n2690) );
  NAND U4034 ( .A(n2692), .B(n2693), .Z(z2[716]) );
  NANDN U4035 ( .A(xregN_1), .B(zin[715]), .Z(n2693) );
  NAND U4036 ( .A(N720), .B(xregN_1), .Z(n2692) );
  NAND U4037 ( .A(n2694), .B(n2695), .Z(z2[715]) );
  NANDN U4038 ( .A(xregN_1), .B(zin[714]), .Z(n2695) );
  NAND U4039 ( .A(N719), .B(xregN_1), .Z(n2694) );
  NAND U4040 ( .A(n2696), .B(n2697), .Z(z2[714]) );
  NANDN U4041 ( .A(xregN_1), .B(zin[713]), .Z(n2697) );
  NAND U4042 ( .A(N718), .B(xregN_1), .Z(n2696) );
  NAND U4043 ( .A(n2698), .B(n2699), .Z(z2[713]) );
  NANDN U4044 ( .A(xregN_1), .B(zin[712]), .Z(n2699) );
  NAND U4045 ( .A(N717), .B(xregN_1), .Z(n2698) );
  NAND U4046 ( .A(n2700), .B(n2701), .Z(z2[712]) );
  NANDN U4047 ( .A(xregN_1), .B(zin[711]), .Z(n2701) );
  NAND U4048 ( .A(N716), .B(xregN_1), .Z(n2700) );
  NAND U4049 ( .A(n2702), .B(n2703), .Z(z2[711]) );
  NANDN U4050 ( .A(xregN_1), .B(zin[710]), .Z(n2703) );
  NAND U4051 ( .A(N715), .B(xregN_1), .Z(n2702) );
  NAND U4052 ( .A(n2704), .B(n2705), .Z(z2[710]) );
  NANDN U4053 ( .A(xregN_1), .B(zin[709]), .Z(n2705) );
  NAND U4054 ( .A(N714), .B(xregN_1), .Z(n2704) );
  NAND U4055 ( .A(n2706), .B(n2707), .Z(z2[70]) );
  NANDN U4056 ( .A(xregN_1), .B(zin[69]), .Z(n2707) );
  NAND U4057 ( .A(N74), .B(xregN_1), .Z(n2706) );
  NAND U4058 ( .A(n2708), .B(n2709), .Z(z2[709]) );
  NANDN U4059 ( .A(xregN_1), .B(zin[708]), .Z(n2709) );
  NAND U4060 ( .A(N713), .B(xregN_1), .Z(n2708) );
  NAND U4061 ( .A(n2710), .B(n2711), .Z(z2[708]) );
  NANDN U4062 ( .A(xregN_1), .B(zin[707]), .Z(n2711) );
  NAND U4063 ( .A(N712), .B(xregN_1), .Z(n2710) );
  NAND U4064 ( .A(n2712), .B(n2713), .Z(z2[707]) );
  NANDN U4065 ( .A(xregN_1), .B(zin[706]), .Z(n2713) );
  NAND U4066 ( .A(N711), .B(xregN_1), .Z(n2712) );
  NAND U4067 ( .A(n2714), .B(n2715), .Z(z2[706]) );
  NANDN U4068 ( .A(xregN_1), .B(zin[705]), .Z(n2715) );
  NAND U4069 ( .A(N710), .B(xregN_1), .Z(n2714) );
  NAND U4070 ( .A(n2716), .B(n2717), .Z(z2[705]) );
  NANDN U4071 ( .A(xregN_1), .B(zin[704]), .Z(n2717) );
  NAND U4072 ( .A(N709), .B(xregN_1), .Z(n2716) );
  NAND U4073 ( .A(n2718), .B(n2719), .Z(z2[704]) );
  NANDN U4074 ( .A(xregN_1), .B(zin[703]), .Z(n2719) );
  NAND U4075 ( .A(N708), .B(xregN_1), .Z(n2718) );
  NAND U4076 ( .A(n2720), .B(n2721), .Z(z2[703]) );
  NANDN U4077 ( .A(xregN_1), .B(zin[702]), .Z(n2721) );
  NAND U4078 ( .A(N707), .B(xregN_1), .Z(n2720) );
  NAND U4079 ( .A(n2722), .B(n2723), .Z(z2[702]) );
  NANDN U4080 ( .A(xregN_1), .B(zin[701]), .Z(n2723) );
  NAND U4081 ( .A(N706), .B(xregN_1), .Z(n2722) );
  NAND U4082 ( .A(n2724), .B(n2725), .Z(z2[701]) );
  NANDN U4083 ( .A(xregN_1), .B(zin[700]), .Z(n2725) );
  NAND U4084 ( .A(N705), .B(xregN_1), .Z(n2724) );
  NAND U4085 ( .A(n2726), .B(n2727), .Z(z2[700]) );
  NANDN U4086 ( .A(xregN_1), .B(zin[699]), .Z(n2727) );
  NAND U4087 ( .A(N704), .B(xregN_1), .Z(n2726) );
  NAND U4088 ( .A(n2728), .B(n2729), .Z(z2[6]) );
  NANDN U4089 ( .A(xregN_1), .B(zin[5]), .Z(n2729) );
  NAND U4090 ( .A(N10), .B(xregN_1), .Z(n2728) );
  NAND U4091 ( .A(n2730), .B(n2731), .Z(z2[69]) );
  NANDN U4092 ( .A(xregN_1), .B(zin[68]), .Z(n2731) );
  NAND U4093 ( .A(N73), .B(xregN_1), .Z(n2730) );
  NAND U4094 ( .A(n2732), .B(n2733), .Z(z2[699]) );
  NANDN U4095 ( .A(xregN_1), .B(zin[698]), .Z(n2733) );
  NAND U4096 ( .A(N703), .B(xregN_1), .Z(n2732) );
  NAND U4097 ( .A(n2734), .B(n2735), .Z(z2[698]) );
  NANDN U4098 ( .A(xregN_1), .B(zin[697]), .Z(n2735) );
  NAND U4099 ( .A(N702), .B(xregN_1), .Z(n2734) );
  NAND U4100 ( .A(n2736), .B(n2737), .Z(z2[697]) );
  NANDN U4101 ( .A(xregN_1), .B(zin[696]), .Z(n2737) );
  NAND U4102 ( .A(N701), .B(xregN_1), .Z(n2736) );
  NAND U4103 ( .A(n2738), .B(n2739), .Z(z2[696]) );
  NANDN U4104 ( .A(xregN_1), .B(zin[695]), .Z(n2739) );
  NAND U4105 ( .A(N700), .B(xregN_1), .Z(n2738) );
  NAND U4106 ( .A(n2740), .B(n2741), .Z(z2[695]) );
  NANDN U4107 ( .A(xregN_1), .B(zin[694]), .Z(n2741) );
  NAND U4108 ( .A(N699), .B(xregN_1), .Z(n2740) );
  NAND U4109 ( .A(n2742), .B(n2743), .Z(z2[694]) );
  NANDN U4110 ( .A(xregN_1), .B(zin[693]), .Z(n2743) );
  NAND U4111 ( .A(N698), .B(xregN_1), .Z(n2742) );
  NAND U4112 ( .A(n2744), .B(n2745), .Z(z2[693]) );
  NANDN U4113 ( .A(xregN_1), .B(zin[692]), .Z(n2745) );
  NAND U4114 ( .A(N697), .B(xregN_1), .Z(n2744) );
  NAND U4115 ( .A(n2746), .B(n2747), .Z(z2[692]) );
  NANDN U4116 ( .A(xregN_1), .B(zin[691]), .Z(n2747) );
  NAND U4117 ( .A(N696), .B(xregN_1), .Z(n2746) );
  NAND U4118 ( .A(n2748), .B(n2749), .Z(z2[691]) );
  NANDN U4119 ( .A(xregN_1), .B(zin[690]), .Z(n2749) );
  NAND U4120 ( .A(N695), .B(xregN_1), .Z(n2748) );
  NAND U4121 ( .A(n2750), .B(n2751), .Z(z2[690]) );
  NANDN U4122 ( .A(xregN_1), .B(zin[689]), .Z(n2751) );
  NAND U4123 ( .A(N694), .B(xregN_1), .Z(n2750) );
  NAND U4124 ( .A(n2752), .B(n2753), .Z(z2[68]) );
  NANDN U4125 ( .A(xregN_1), .B(zin[67]), .Z(n2753) );
  NAND U4126 ( .A(N72), .B(xregN_1), .Z(n2752) );
  NAND U4127 ( .A(n2754), .B(n2755), .Z(z2[689]) );
  NANDN U4128 ( .A(xregN_1), .B(zin[688]), .Z(n2755) );
  NAND U4129 ( .A(N693), .B(xregN_1), .Z(n2754) );
  NAND U4130 ( .A(n2756), .B(n2757), .Z(z2[688]) );
  NANDN U4131 ( .A(xregN_1), .B(zin[687]), .Z(n2757) );
  NAND U4132 ( .A(N692), .B(xregN_1), .Z(n2756) );
  NAND U4133 ( .A(n2758), .B(n2759), .Z(z2[687]) );
  NANDN U4134 ( .A(xregN_1), .B(zin[686]), .Z(n2759) );
  NAND U4135 ( .A(N691), .B(xregN_1), .Z(n2758) );
  NAND U4136 ( .A(n2760), .B(n2761), .Z(z2[686]) );
  NANDN U4137 ( .A(xregN_1), .B(zin[685]), .Z(n2761) );
  NAND U4138 ( .A(N690), .B(xregN_1), .Z(n2760) );
  NAND U4139 ( .A(n2762), .B(n2763), .Z(z2[685]) );
  NANDN U4140 ( .A(xregN_1), .B(zin[684]), .Z(n2763) );
  NAND U4141 ( .A(N689), .B(xregN_1), .Z(n2762) );
  NAND U4142 ( .A(n2764), .B(n2765), .Z(z2[684]) );
  NANDN U4143 ( .A(xregN_1), .B(zin[683]), .Z(n2765) );
  NAND U4144 ( .A(N688), .B(xregN_1), .Z(n2764) );
  NAND U4145 ( .A(n2766), .B(n2767), .Z(z2[683]) );
  NANDN U4146 ( .A(xregN_1), .B(zin[682]), .Z(n2767) );
  NAND U4147 ( .A(N687), .B(xregN_1), .Z(n2766) );
  NAND U4148 ( .A(n2768), .B(n2769), .Z(z2[682]) );
  NANDN U4149 ( .A(xregN_1), .B(zin[681]), .Z(n2769) );
  NAND U4150 ( .A(N686), .B(xregN_1), .Z(n2768) );
  NAND U4151 ( .A(n2770), .B(n2771), .Z(z2[681]) );
  NANDN U4152 ( .A(xregN_1), .B(zin[680]), .Z(n2771) );
  NAND U4153 ( .A(N685), .B(xregN_1), .Z(n2770) );
  NAND U4154 ( .A(n2772), .B(n2773), .Z(z2[680]) );
  NANDN U4155 ( .A(xregN_1), .B(zin[679]), .Z(n2773) );
  NAND U4156 ( .A(N684), .B(xregN_1), .Z(n2772) );
  NAND U4157 ( .A(n2774), .B(n2775), .Z(z2[67]) );
  NANDN U4158 ( .A(xregN_1), .B(zin[66]), .Z(n2775) );
  NAND U4159 ( .A(N71), .B(xregN_1), .Z(n2774) );
  NAND U4160 ( .A(n2776), .B(n2777), .Z(z2[679]) );
  NANDN U4161 ( .A(xregN_1), .B(zin[678]), .Z(n2777) );
  NAND U4162 ( .A(N683), .B(xregN_1), .Z(n2776) );
  NAND U4163 ( .A(n2778), .B(n2779), .Z(z2[678]) );
  NANDN U4164 ( .A(xregN_1), .B(zin[677]), .Z(n2779) );
  NAND U4165 ( .A(N682), .B(xregN_1), .Z(n2778) );
  NAND U4166 ( .A(n2780), .B(n2781), .Z(z2[677]) );
  NANDN U4167 ( .A(xregN_1), .B(zin[676]), .Z(n2781) );
  NAND U4168 ( .A(N681), .B(xregN_1), .Z(n2780) );
  NAND U4169 ( .A(n2782), .B(n2783), .Z(z2[676]) );
  NANDN U4170 ( .A(xregN_1), .B(zin[675]), .Z(n2783) );
  NAND U4171 ( .A(N680), .B(xregN_1), .Z(n2782) );
  NAND U4172 ( .A(n2784), .B(n2785), .Z(z2[675]) );
  NANDN U4173 ( .A(xregN_1), .B(zin[674]), .Z(n2785) );
  NAND U4174 ( .A(N679), .B(xregN_1), .Z(n2784) );
  NAND U4175 ( .A(n2786), .B(n2787), .Z(z2[674]) );
  NANDN U4176 ( .A(xregN_1), .B(zin[673]), .Z(n2787) );
  NAND U4177 ( .A(N678), .B(xregN_1), .Z(n2786) );
  NAND U4178 ( .A(n2788), .B(n2789), .Z(z2[673]) );
  NANDN U4179 ( .A(xregN_1), .B(zin[672]), .Z(n2789) );
  NAND U4180 ( .A(N677), .B(xregN_1), .Z(n2788) );
  NAND U4181 ( .A(n2790), .B(n2791), .Z(z2[672]) );
  NANDN U4182 ( .A(xregN_1), .B(zin[671]), .Z(n2791) );
  NAND U4183 ( .A(N676), .B(xregN_1), .Z(n2790) );
  NAND U4184 ( .A(n2792), .B(n2793), .Z(z2[671]) );
  NANDN U4185 ( .A(xregN_1), .B(zin[670]), .Z(n2793) );
  NAND U4186 ( .A(N675), .B(xregN_1), .Z(n2792) );
  NAND U4187 ( .A(n2794), .B(n2795), .Z(z2[670]) );
  NANDN U4188 ( .A(xregN_1), .B(zin[669]), .Z(n2795) );
  NAND U4189 ( .A(N674), .B(xregN_1), .Z(n2794) );
  NAND U4190 ( .A(n2796), .B(n2797), .Z(z2[66]) );
  NANDN U4191 ( .A(xregN_1), .B(zin[65]), .Z(n2797) );
  NAND U4192 ( .A(N70), .B(xregN_1), .Z(n2796) );
  NAND U4193 ( .A(n2798), .B(n2799), .Z(z2[669]) );
  NANDN U4194 ( .A(xregN_1), .B(zin[668]), .Z(n2799) );
  NAND U4195 ( .A(N673), .B(xregN_1), .Z(n2798) );
  NAND U4196 ( .A(n2800), .B(n2801), .Z(z2[668]) );
  NANDN U4197 ( .A(xregN_1), .B(zin[667]), .Z(n2801) );
  NAND U4198 ( .A(N672), .B(xregN_1), .Z(n2800) );
  NAND U4199 ( .A(n2802), .B(n2803), .Z(z2[667]) );
  NANDN U4200 ( .A(xregN_1), .B(zin[666]), .Z(n2803) );
  NAND U4201 ( .A(N671), .B(xregN_1), .Z(n2802) );
  NAND U4202 ( .A(n2804), .B(n2805), .Z(z2[666]) );
  NANDN U4203 ( .A(xregN_1), .B(zin[665]), .Z(n2805) );
  NAND U4204 ( .A(N670), .B(xregN_1), .Z(n2804) );
  NAND U4205 ( .A(n2806), .B(n2807), .Z(z2[665]) );
  NANDN U4206 ( .A(xregN_1), .B(zin[664]), .Z(n2807) );
  NAND U4207 ( .A(N669), .B(xregN_1), .Z(n2806) );
  NAND U4208 ( .A(n2808), .B(n2809), .Z(z2[664]) );
  NANDN U4209 ( .A(xregN_1), .B(zin[663]), .Z(n2809) );
  NAND U4210 ( .A(N668), .B(xregN_1), .Z(n2808) );
  NAND U4211 ( .A(n2810), .B(n2811), .Z(z2[663]) );
  NANDN U4212 ( .A(xregN_1), .B(zin[662]), .Z(n2811) );
  NAND U4213 ( .A(N667), .B(xregN_1), .Z(n2810) );
  NAND U4214 ( .A(n2812), .B(n2813), .Z(z2[662]) );
  NANDN U4215 ( .A(xregN_1), .B(zin[661]), .Z(n2813) );
  NAND U4216 ( .A(N666), .B(xregN_1), .Z(n2812) );
  NAND U4217 ( .A(n2814), .B(n2815), .Z(z2[661]) );
  NANDN U4218 ( .A(xregN_1), .B(zin[660]), .Z(n2815) );
  NAND U4219 ( .A(N665), .B(xregN_1), .Z(n2814) );
  NAND U4220 ( .A(n2816), .B(n2817), .Z(z2[660]) );
  NANDN U4221 ( .A(xregN_1), .B(zin[659]), .Z(n2817) );
  NAND U4222 ( .A(N664), .B(xregN_1), .Z(n2816) );
  NAND U4223 ( .A(n2818), .B(n2819), .Z(z2[65]) );
  NANDN U4224 ( .A(xregN_1), .B(zin[64]), .Z(n2819) );
  NAND U4225 ( .A(N69), .B(xregN_1), .Z(n2818) );
  NAND U4226 ( .A(n2820), .B(n2821), .Z(z2[659]) );
  NANDN U4227 ( .A(xregN_1), .B(zin[658]), .Z(n2821) );
  NAND U4228 ( .A(N663), .B(xregN_1), .Z(n2820) );
  NAND U4229 ( .A(n2822), .B(n2823), .Z(z2[658]) );
  NANDN U4230 ( .A(xregN_1), .B(zin[657]), .Z(n2823) );
  NAND U4231 ( .A(N662), .B(xregN_1), .Z(n2822) );
  NAND U4232 ( .A(n2824), .B(n2825), .Z(z2[657]) );
  NANDN U4233 ( .A(xregN_1), .B(zin[656]), .Z(n2825) );
  NAND U4234 ( .A(N661), .B(xregN_1), .Z(n2824) );
  NAND U4235 ( .A(n2826), .B(n2827), .Z(z2[656]) );
  NANDN U4236 ( .A(xregN_1), .B(zin[655]), .Z(n2827) );
  NAND U4237 ( .A(N660), .B(xregN_1), .Z(n2826) );
  NAND U4238 ( .A(n2828), .B(n2829), .Z(z2[655]) );
  NANDN U4239 ( .A(xregN_1), .B(zin[654]), .Z(n2829) );
  NAND U4240 ( .A(N659), .B(xregN_1), .Z(n2828) );
  NAND U4241 ( .A(n2830), .B(n2831), .Z(z2[654]) );
  NANDN U4242 ( .A(xregN_1), .B(zin[653]), .Z(n2831) );
  NAND U4243 ( .A(N658), .B(xregN_1), .Z(n2830) );
  NAND U4244 ( .A(n2832), .B(n2833), .Z(z2[653]) );
  NANDN U4245 ( .A(xregN_1), .B(zin[652]), .Z(n2833) );
  NAND U4246 ( .A(N657), .B(xregN_1), .Z(n2832) );
  NAND U4247 ( .A(n2834), .B(n2835), .Z(z2[652]) );
  NANDN U4248 ( .A(xregN_1), .B(zin[651]), .Z(n2835) );
  NAND U4249 ( .A(N656), .B(xregN_1), .Z(n2834) );
  NAND U4250 ( .A(n2836), .B(n2837), .Z(z2[651]) );
  NANDN U4251 ( .A(xregN_1), .B(zin[650]), .Z(n2837) );
  NAND U4252 ( .A(N655), .B(xregN_1), .Z(n2836) );
  NAND U4253 ( .A(n2838), .B(n2839), .Z(z2[650]) );
  NANDN U4254 ( .A(xregN_1), .B(zin[649]), .Z(n2839) );
  NAND U4255 ( .A(N654), .B(xregN_1), .Z(n2838) );
  NAND U4256 ( .A(n2840), .B(n2841), .Z(z2[64]) );
  NANDN U4257 ( .A(xregN_1), .B(zin[63]), .Z(n2841) );
  NAND U4258 ( .A(N68), .B(xregN_1), .Z(n2840) );
  NAND U4259 ( .A(n2842), .B(n2843), .Z(z2[649]) );
  NANDN U4260 ( .A(xregN_1), .B(zin[648]), .Z(n2843) );
  NAND U4261 ( .A(N653), .B(xregN_1), .Z(n2842) );
  NAND U4262 ( .A(n2844), .B(n2845), .Z(z2[648]) );
  NANDN U4263 ( .A(xregN_1), .B(zin[647]), .Z(n2845) );
  NAND U4264 ( .A(N652), .B(xregN_1), .Z(n2844) );
  NAND U4265 ( .A(n2846), .B(n2847), .Z(z2[647]) );
  NANDN U4266 ( .A(xregN_1), .B(zin[646]), .Z(n2847) );
  NAND U4267 ( .A(N651), .B(xregN_1), .Z(n2846) );
  NAND U4268 ( .A(n2848), .B(n2849), .Z(z2[646]) );
  NANDN U4269 ( .A(xregN_1), .B(zin[645]), .Z(n2849) );
  NAND U4270 ( .A(N650), .B(xregN_1), .Z(n2848) );
  NAND U4271 ( .A(n2850), .B(n2851), .Z(z2[645]) );
  NANDN U4272 ( .A(xregN_1), .B(zin[644]), .Z(n2851) );
  NAND U4273 ( .A(N649), .B(xregN_1), .Z(n2850) );
  NAND U4274 ( .A(n2852), .B(n2853), .Z(z2[644]) );
  NANDN U4275 ( .A(xregN_1), .B(zin[643]), .Z(n2853) );
  NAND U4276 ( .A(N648), .B(xregN_1), .Z(n2852) );
  NAND U4277 ( .A(n2854), .B(n2855), .Z(z2[643]) );
  NANDN U4278 ( .A(xregN_1), .B(zin[642]), .Z(n2855) );
  NAND U4279 ( .A(N647), .B(xregN_1), .Z(n2854) );
  NAND U4280 ( .A(n2856), .B(n2857), .Z(z2[642]) );
  NANDN U4281 ( .A(xregN_1), .B(zin[641]), .Z(n2857) );
  NAND U4282 ( .A(N646), .B(xregN_1), .Z(n2856) );
  NAND U4283 ( .A(n2858), .B(n2859), .Z(z2[641]) );
  NANDN U4284 ( .A(xregN_1), .B(zin[640]), .Z(n2859) );
  NAND U4285 ( .A(N645), .B(xregN_1), .Z(n2858) );
  NAND U4286 ( .A(n2860), .B(n2861), .Z(z2[640]) );
  NANDN U4287 ( .A(xregN_1), .B(zin[639]), .Z(n2861) );
  NAND U4288 ( .A(N644), .B(xregN_1), .Z(n2860) );
  NAND U4289 ( .A(n2862), .B(n2863), .Z(z2[63]) );
  NANDN U4290 ( .A(xregN_1), .B(zin[62]), .Z(n2863) );
  NAND U4291 ( .A(N67), .B(xregN_1), .Z(n2862) );
  NAND U4292 ( .A(n2864), .B(n2865), .Z(z2[639]) );
  NANDN U4293 ( .A(xregN_1), .B(zin[638]), .Z(n2865) );
  NAND U4294 ( .A(N643), .B(xregN_1), .Z(n2864) );
  NAND U4295 ( .A(n2866), .B(n2867), .Z(z2[638]) );
  NANDN U4296 ( .A(xregN_1), .B(zin[637]), .Z(n2867) );
  NAND U4297 ( .A(N642), .B(xregN_1), .Z(n2866) );
  NAND U4298 ( .A(n2868), .B(n2869), .Z(z2[637]) );
  NANDN U4299 ( .A(xregN_1), .B(zin[636]), .Z(n2869) );
  NAND U4300 ( .A(N641), .B(xregN_1), .Z(n2868) );
  NAND U4301 ( .A(n2870), .B(n2871), .Z(z2[636]) );
  NANDN U4302 ( .A(xregN_1), .B(zin[635]), .Z(n2871) );
  NAND U4303 ( .A(N640), .B(xregN_1), .Z(n2870) );
  NAND U4304 ( .A(n2872), .B(n2873), .Z(z2[635]) );
  NANDN U4305 ( .A(xregN_1), .B(zin[634]), .Z(n2873) );
  NAND U4306 ( .A(N639), .B(xregN_1), .Z(n2872) );
  NAND U4307 ( .A(n2874), .B(n2875), .Z(z2[634]) );
  NANDN U4308 ( .A(xregN_1), .B(zin[633]), .Z(n2875) );
  NAND U4309 ( .A(N638), .B(xregN_1), .Z(n2874) );
  NAND U4310 ( .A(n2876), .B(n2877), .Z(z2[633]) );
  NANDN U4311 ( .A(xregN_1), .B(zin[632]), .Z(n2877) );
  NAND U4312 ( .A(N637), .B(xregN_1), .Z(n2876) );
  NAND U4313 ( .A(n2878), .B(n2879), .Z(z2[632]) );
  NANDN U4314 ( .A(xregN_1), .B(zin[631]), .Z(n2879) );
  NAND U4315 ( .A(N636), .B(xregN_1), .Z(n2878) );
  NAND U4316 ( .A(n2880), .B(n2881), .Z(z2[631]) );
  NANDN U4317 ( .A(xregN_1), .B(zin[630]), .Z(n2881) );
  NAND U4318 ( .A(N635), .B(xregN_1), .Z(n2880) );
  NAND U4319 ( .A(n2882), .B(n2883), .Z(z2[630]) );
  NANDN U4320 ( .A(xregN_1), .B(zin[629]), .Z(n2883) );
  NAND U4321 ( .A(N634), .B(xregN_1), .Z(n2882) );
  NAND U4322 ( .A(n2884), .B(n2885), .Z(z2[62]) );
  NANDN U4323 ( .A(xregN_1), .B(zin[61]), .Z(n2885) );
  NAND U4324 ( .A(N66), .B(xregN_1), .Z(n2884) );
  NAND U4325 ( .A(n2886), .B(n2887), .Z(z2[629]) );
  NANDN U4326 ( .A(xregN_1), .B(zin[628]), .Z(n2887) );
  NAND U4327 ( .A(N633), .B(xregN_1), .Z(n2886) );
  NAND U4328 ( .A(n2888), .B(n2889), .Z(z2[628]) );
  NANDN U4329 ( .A(xregN_1), .B(zin[627]), .Z(n2889) );
  NAND U4330 ( .A(N632), .B(xregN_1), .Z(n2888) );
  NAND U4331 ( .A(n2890), .B(n2891), .Z(z2[627]) );
  NANDN U4332 ( .A(xregN_1), .B(zin[626]), .Z(n2891) );
  NAND U4333 ( .A(N631), .B(xregN_1), .Z(n2890) );
  NAND U4334 ( .A(n2892), .B(n2893), .Z(z2[626]) );
  NANDN U4335 ( .A(xregN_1), .B(zin[625]), .Z(n2893) );
  NAND U4336 ( .A(N630), .B(xregN_1), .Z(n2892) );
  NAND U4337 ( .A(n2894), .B(n2895), .Z(z2[625]) );
  NANDN U4338 ( .A(xregN_1), .B(zin[624]), .Z(n2895) );
  NAND U4339 ( .A(N629), .B(xregN_1), .Z(n2894) );
  NAND U4340 ( .A(n2896), .B(n2897), .Z(z2[624]) );
  NANDN U4341 ( .A(xregN_1), .B(zin[623]), .Z(n2897) );
  NAND U4342 ( .A(N628), .B(xregN_1), .Z(n2896) );
  NAND U4343 ( .A(n2898), .B(n2899), .Z(z2[623]) );
  NANDN U4344 ( .A(xregN_1), .B(zin[622]), .Z(n2899) );
  NAND U4345 ( .A(N627), .B(xregN_1), .Z(n2898) );
  NAND U4346 ( .A(n2900), .B(n2901), .Z(z2[622]) );
  NANDN U4347 ( .A(xregN_1), .B(zin[621]), .Z(n2901) );
  NAND U4348 ( .A(N626), .B(xregN_1), .Z(n2900) );
  NAND U4349 ( .A(n2902), .B(n2903), .Z(z2[621]) );
  NANDN U4350 ( .A(xregN_1), .B(zin[620]), .Z(n2903) );
  NAND U4351 ( .A(N625), .B(xregN_1), .Z(n2902) );
  NAND U4352 ( .A(n2904), .B(n2905), .Z(z2[620]) );
  NANDN U4353 ( .A(xregN_1), .B(zin[619]), .Z(n2905) );
  NAND U4354 ( .A(N624), .B(xregN_1), .Z(n2904) );
  NAND U4355 ( .A(n2906), .B(n2907), .Z(z2[61]) );
  NANDN U4356 ( .A(xregN_1), .B(zin[60]), .Z(n2907) );
  NAND U4357 ( .A(N65), .B(xregN_1), .Z(n2906) );
  NAND U4358 ( .A(n2908), .B(n2909), .Z(z2[619]) );
  NANDN U4359 ( .A(xregN_1), .B(zin[618]), .Z(n2909) );
  NAND U4360 ( .A(N623), .B(xregN_1), .Z(n2908) );
  NAND U4361 ( .A(n2910), .B(n2911), .Z(z2[618]) );
  NANDN U4362 ( .A(xregN_1), .B(zin[617]), .Z(n2911) );
  NAND U4363 ( .A(N622), .B(xregN_1), .Z(n2910) );
  NAND U4364 ( .A(n2912), .B(n2913), .Z(z2[617]) );
  NANDN U4365 ( .A(xregN_1), .B(zin[616]), .Z(n2913) );
  NAND U4366 ( .A(N621), .B(xregN_1), .Z(n2912) );
  NAND U4367 ( .A(n2914), .B(n2915), .Z(z2[616]) );
  NANDN U4368 ( .A(xregN_1), .B(zin[615]), .Z(n2915) );
  NAND U4369 ( .A(N620), .B(xregN_1), .Z(n2914) );
  NAND U4370 ( .A(n2916), .B(n2917), .Z(z2[615]) );
  NANDN U4371 ( .A(xregN_1), .B(zin[614]), .Z(n2917) );
  NAND U4372 ( .A(N619), .B(xregN_1), .Z(n2916) );
  NAND U4373 ( .A(n2918), .B(n2919), .Z(z2[614]) );
  NANDN U4374 ( .A(xregN_1), .B(zin[613]), .Z(n2919) );
  NAND U4375 ( .A(N618), .B(xregN_1), .Z(n2918) );
  NAND U4376 ( .A(n2920), .B(n2921), .Z(z2[613]) );
  NANDN U4377 ( .A(xregN_1), .B(zin[612]), .Z(n2921) );
  NAND U4378 ( .A(N617), .B(xregN_1), .Z(n2920) );
  NAND U4379 ( .A(n2922), .B(n2923), .Z(z2[612]) );
  NANDN U4380 ( .A(xregN_1), .B(zin[611]), .Z(n2923) );
  NAND U4381 ( .A(N616), .B(xregN_1), .Z(n2922) );
  NAND U4382 ( .A(n2924), .B(n2925), .Z(z2[611]) );
  NANDN U4383 ( .A(xregN_1), .B(zin[610]), .Z(n2925) );
  NAND U4384 ( .A(N615), .B(xregN_1), .Z(n2924) );
  NAND U4385 ( .A(n2926), .B(n2927), .Z(z2[610]) );
  NANDN U4386 ( .A(xregN_1), .B(zin[609]), .Z(n2927) );
  NAND U4387 ( .A(N614), .B(xregN_1), .Z(n2926) );
  NAND U4388 ( .A(n2928), .B(n2929), .Z(z2[60]) );
  NANDN U4389 ( .A(xregN_1), .B(zin[59]), .Z(n2929) );
  NAND U4390 ( .A(N64), .B(xregN_1), .Z(n2928) );
  NAND U4391 ( .A(n2930), .B(n2931), .Z(z2[609]) );
  NANDN U4392 ( .A(xregN_1), .B(zin[608]), .Z(n2931) );
  NAND U4393 ( .A(N613), .B(xregN_1), .Z(n2930) );
  NAND U4394 ( .A(n2932), .B(n2933), .Z(z2[608]) );
  NANDN U4395 ( .A(xregN_1), .B(zin[607]), .Z(n2933) );
  NAND U4396 ( .A(N612), .B(xregN_1), .Z(n2932) );
  NAND U4397 ( .A(n2934), .B(n2935), .Z(z2[607]) );
  NANDN U4398 ( .A(xregN_1), .B(zin[606]), .Z(n2935) );
  NAND U4399 ( .A(N611), .B(xregN_1), .Z(n2934) );
  NAND U4400 ( .A(n2936), .B(n2937), .Z(z2[606]) );
  NANDN U4401 ( .A(xregN_1), .B(zin[605]), .Z(n2937) );
  NAND U4402 ( .A(N610), .B(xregN_1), .Z(n2936) );
  NAND U4403 ( .A(n2938), .B(n2939), .Z(z2[605]) );
  NANDN U4404 ( .A(xregN_1), .B(zin[604]), .Z(n2939) );
  NAND U4405 ( .A(N609), .B(xregN_1), .Z(n2938) );
  NAND U4406 ( .A(n2940), .B(n2941), .Z(z2[604]) );
  NANDN U4407 ( .A(xregN_1), .B(zin[603]), .Z(n2941) );
  NAND U4408 ( .A(N608), .B(xregN_1), .Z(n2940) );
  NAND U4409 ( .A(n2942), .B(n2943), .Z(z2[603]) );
  NANDN U4410 ( .A(xregN_1), .B(zin[602]), .Z(n2943) );
  NAND U4411 ( .A(N607), .B(xregN_1), .Z(n2942) );
  NAND U4412 ( .A(n2944), .B(n2945), .Z(z2[602]) );
  NANDN U4413 ( .A(xregN_1), .B(zin[601]), .Z(n2945) );
  NAND U4414 ( .A(N606), .B(xregN_1), .Z(n2944) );
  NAND U4415 ( .A(n2946), .B(n2947), .Z(z2[601]) );
  NANDN U4416 ( .A(xregN_1), .B(zin[600]), .Z(n2947) );
  NAND U4417 ( .A(N605), .B(xregN_1), .Z(n2946) );
  NAND U4418 ( .A(n2948), .B(n2949), .Z(z2[600]) );
  NANDN U4419 ( .A(xregN_1), .B(zin[599]), .Z(n2949) );
  NAND U4420 ( .A(N604), .B(xregN_1), .Z(n2948) );
  NAND U4421 ( .A(n2950), .B(n2951), .Z(z2[5]) );
  NANDN U4422 ( .A(xregN_1), .B(zin[4]), .Z(n2951) );
  NAND U4423 ( .A(N9), .B(xregN_1), .Z(n2950) );
  NAND U4424 ( .A(n2952), .B(n2953), .Z(z2[59]) );
  NANDN U4425 ( .A(xregN_1), .B(zin[58]), .Z(n2953) );
  NAND U4426 ( .A(N63), .B(xregN_1), .Z(n2952) );
  NAND U4427 ( .A(n2954), .B(n2955), .Z(z2[599]) );
  NANDN U4428 ( .A(xregN_1), .B(zin[598]), .Z(n2955) );
  NAND U4429 ( .A(N603), .B(xregN_1), .Z(n2954) );
  NAND U4430 ( .A(n2956), .B(n2957), .Z(z2[598]) );
  NANDN U4431 ( .A(xregN_1), .B(zin[597]), .Z(n2957) );
  NAND U4432 ( .A(N602), .B(xregN_1), .Z(n2956) );
  NAND U4433 ( .A(n2958), .B(n2959), .Z(z2[597]) );
  NANDN U4434 ( .A(xregN_1), .B(zin[596]), .Z(n2959) );
  NAND U4435 ( .A(N601), .B(xregN_1), .Z(n2958) );
  NAND U4436 ( .A(n2960), .B(n2961), .Z(z2[596]) );
  NANDN U4437 ( .A(xregN_1), .B(zin[595]), .Z(n2961) );
  NAND U4438 ( .A(N600), .B(xregN_1), .Z(n2960) );
  NAND U4439 ( .A(n2962), .B(n2963), .Z(z2[595]) );
  NANDN U4440 ( .A(xregN_1), .B(zin[594]), .Z(n2963) );
  NAND U4441 ( .A(N599), .B(xregN_1), .Z(n2962) );
  NAND U4442 ( .A(n2964), .B(n2965), .Z(z2[594]) );
  NANDN U4443 ( .A(xregN_1), .B(zin[593]), .Z(n2965) );
  NAND U4444 ( .A(N598), .B(xregN_1), .Z(n2964) );
  NAND U4445 ( .A(n2966), .B(n2967), .Z(z2[593]) );
  NANDN U4446 ( .A(xregN_1), .B(zin[592]), .Z(n2967) );
  NAND U4447 ( .A(N597), .B(xregN_1), .Z(n2966) );
  NAND U4448 ( .A(n2968), .B(n2969), .Z(z2[592]) );
  NANDN U4449 ( .A(xregN_1), .B(zin[591]), .Z(n2969) );
  NAND U4450 ( .A(N596), .B(xregN_1), .Z(n2968) );
  NAND U4451 ( .A(n2970), .B(n2971), .Z(z2[591]) );
  NANDN U4452 ( .A(xregN_1), .B(zin[590]), .Z(n2971) );
  NAND U4453 ( .A(N595), .B(xregN_1), .Z(n2970) );
  NAND U4454 ( .A(n2972), .B(n2973), .Z(z2[590]) );
  NANDN U4455 ( .A(xregN_1), .B(zin[589]), .Z(n2973) );
  NAND U4456 ( .A(N594), .B(xregN_1), .Z(n2972) );
  NAND U4457 ( .A(n2974), .B(n2975), .Z(z2[58]) );
  NANDN U4458 ( .A(xregN_1), .B(zin[57]), .Z(n2975) );
  NAND U4459 ( .A(N62), .B(xregN_1), .Z(n2974) );
  NAND U4460 ( .A(n2976), .B(n2977), .Z(z2[589]) );
  NANDN U4461 ( .A(xregN_1), .B(zin[588]), .Z(n2977) );
  NAND U4462 ( .A(N593), .B(xregN_1), .Z(n2976) );
  NAND U4463 ( .A(n2978), .B(n2979), .Z(z2[588]) );
  NANDN U4464 ( .A(xregN_1), .B(zin[587]), .Z(n2979) );
  NAND U4465 ( .A(N592), .B(xregN_1), .Z(n2978) );
  NAND U4466 ( .A(n2980), .B(n2981), .Z(z2[587]) );
  NANDN U4467 ( .A(xregN_1), .B(zin[586]), .Z(n2981) );
  NAND U4468 ( .A(N591), .B(xregN_1), .Z(n2980) );
  NAND U4469 ( .A(n2982), .B(n2983), .Z(z2[586]) );
  NANDN U4470 ( .A(xregN_1), .B(zin[585]), .Z(n2983) );
  NAND U4471 ( .A(N590), .B(xregN_1), .Z(n2982) );
  NAND U4472 ( .A(n2984), .B(n2985), .Z(z2[585]) );
  NANDN U4473 ( .A(xregN_1), .B(zin[584]), .Z(n2985) );
  NAND U4474 ( .A(N589), .B(xregN_1), .Z(n2984) );
  NAND U4475 ( .A(n2986), .B(n2987), .Z(z2[584]) );
  NANDN U4476 ( .A(xregN_1), .B(zin[583]), .Z(n2987) );
  NAND U4477 ( .A(N588), .B(xregN_1), .Z(n2986) );
  NAND U4478 ( .A(n2988), .B(n2989), .Z(z2[583]) );
  NANDN U4479 ( .A(xregN_1), .B(zin[582]), .Z(n2989) );
  NAND U4480 ( .A(N587), .B(xregN_1), .Z(n2988) );
  NAND U4481 ( .A(n2990), .B(n2991), .Z(z2[582]) );
  NANDN U4482 ( .A(xregN_1), .B(zin[581]), .Z(n2991) );
  NAND U4483 ( .A(N586), .B(xregN_1), .Z(n2990) );
  NAND U4484 ( .A(n2992), .B(n2993), .Z(z2[581]) );
  NANDN U4485 ( .A(xregN_1), .B(zin[580]), .Z(n2993) );
  NAND U4486 ( .A(N585), .B(xregN_1), .Z(n2992) );
  NAND U4487 ( .A(n2994), .B(n2995), .Z(z2[580]) );
  NANDN U4488 ( .A(xregN_1), .B(zin[579]), .Z(n2995) );
  NAND U4489 ( .A(N584), .B(xregN_1), .Z(n2994) );
  NAND U4490 ( .A(n2996), .B(n2997), .Z(z2[57]) );
  NANDN U4491 ( .A(xregN_1), .B(zin[56]), .Z(n2997) );
  NAND U4492 ( .A(N61), .B(xregN_1), .Z(n2996) );
  NAND U4493 ( .A(n2998), .B(n2999), .Z(z2[579]) );
  NANDN U4494 ( .A(xregN_1), .B(zin[578]), .Z(n2999) );
  NAND U4495 ( .A(N583), .B(xregN_1), .Z(n2998) );
  NAND U4496 ( .A(n3000), .B(n3001), .Z(z2[578]) );
  NANDN U4497 ( .A(xregN_1), .B(zin[577]), .Z(n3001) );
  NAND U4498 ( .A(N582), .B(xregN_1), .Z(n3000) );
  NAND U4499 ( .A(n3002), .B(n3003), .Z(z2[577]) );
  NANDN U4500 ( .A(xregN_1), .B(zin[576]), .Z(n3003) );
  NAND U4501 ( .A(N581), .B(xregN_1), .Z(n3002) );
  NAND U4502 ( .A(n3004), .B(n3005), .Z(z2[576]) );
  NANDN U4503 ( .A(xregN_1), .B(zin[575]), .Z(n3005) );
  NAND U4504 ( .A(N580), .B(xregN_1), .Z(n3004) );
  NAND U4505 ( .A(n3006), .B(n3007), .Z(z2[575]) );
  NANDN U4506 ( .A(xregN_1), .B(zin[574]), .Z(n3007) );
  NAND U4507 ( .A(N579), .B(xregN_1), .Z(n3006) );
  NAND U4508 ( .A(n3008), .B(n3009), .Z(z2[574]) );
  NANDN U4509 ( .A(xregN_1), .B(zin[573]), .Z(n3009) );
  NAND U4510 ( .A(N578), .B(xregN_1), .Z(n3008) );
  NAND U4511 ( .A(n3010), .B(n3011), .Z(z2[573]) );
  NANDN U4512 ( .A(xregN_1), .B(zin[572]), .Z(n3011) );
  NAND U4513 ( .A(N577), .B(xregN_1), .Z(n3010) );
  NAND U4514 ( .A(n3012), .B(n3013), .Z(z2[572]) );
  NANDN U4515 ( .A(xregN_1), .B(zin[571]), .Z(n3013) );
  NAND U4516 ( .A(N576), .B(xregN_1), .Z(n3012) );
  NAND U4517 ( .A(n3014), .B(n3015), .Z(z2[571]) );
  NANDN U4518 ( .A(xregN_1), .B(zin[570]), .Z(n3015) );
  NAND U4519 ( .A(N575), .B(xregN_1), .Z(n3014) );
  NAND U4520 ( .A(n3016), .B(n3017), .Z(z2[570]) );
  NANDN U4521 ( .A(xregN_1), .B(zin[569]), .Z(n3017) );
  NAND U4522 ( .A(N574), .B(xregN_1), .Z(n3016) );
  NAND U4523 ( .A(n3018), .B(n3019), .Z(z2[56]) );
  NANDN U4524 ( .A(xregN_1), .B(zin[55]), .Z(n3019) );
  NAND U4525 ( .A(N60), .B(xregN_1), .Z(n3018) );
  NAND U4526 ( .A(n3020), .B(n3021), .Z(z2[569]) );
  NANDN U4527 ( .A(xregN_1), .B(zin[568]), .Z(n3021) );
  NAND U4528 ( .A(N573), .B(xregN_1), .Z(n3020) );
  NAND U4529 ( .A(n3022), .B(n3023), .Z(z2[568]) );
  NANDN U4530 ( .A(xregN_1), .B(zin[567]), .Z(n3023) );
  NAND U4531 ( .A(N572), .B(xregN_1), .Z(n3022) );
  NAND U4532 ( .A(n3024), .B(n3025), .Z(z2[567]) );
  NANDN U4533 ( .A(xregN_1), .B(zin[566]), .Z(n3025) );
  NAND U4534 ( .A(N571), .B(xregN_1), .Z(n3024) );
  NAND U4535 ( .A(n3026), .B(n3027), .Z(z2[566]) );
  NANDN U4536 ( .A(xregN_1), .B(zin[565]), .Z(n3027) );
  NAND U4537 ( .A(N570), .B(xregN_1), .Z(n3026) );
  NAND U4538 ( .A(n3028), .B(n3029), .Z(z2[565]) );
  NANDN U4539 ( .A(xregN_1), .B(zin[564]), .Z(n3029) );
  NAND U4540 ( .A(N569), .B(xregN_1), .Z(n3028) );
  NAND U4541 ( .A(n3030), .B(n3031), .Z(z2[564]) );
  NANDN U4542 ( .A(xregN_1), .B(zin[563]), .Z(n3031) );
  NAND U4543 ( .A(N568), .B(xregN_1), .Z(n3030) );
  NAND U4544 ( .A(n3032), .B(n3033), .Z(z2[563]) );
  NANDN U4545 ( .A(xregN_1), .B(zin[562]), .Z(n3033) );
  NAND U4546 ( .A(N567), .B(xregN_1), .Z(n3032) );
  NAND U4547 ( .A(n3034), .B(n3035), .Z(z2[562]) );
  NANDN U4548 ( .A(xregN_1), .B(zin[561]), .Z(n3035) );
  NAND U4549 ( .A(N566), .B(xregN_1), .Z(n3034) );
  NAND U4550 ( .A(n3036), .B(n3037), .Z(z2[561]) );
  NANDN U4551 ( .A(xregN_1), .B(zin[560]), .Z(n3037) );
  NAND U4552 ( .A(N565), .B(xregN_1), .Z(n3036) );
  NAND U4553 ( .A(n3038), .B(n3039), .Z(z2[560]) );
  NANDN U4554 ( .A(xregN_1), .B(zin[559]), .Z(n3039) );
  NAND U4555 ( .A(N564), .B(xregN_1), .Z(n3038) );
  NAND U4556 ( .A(n3040), .B(n3041), .Z(z2[55]) );
  NANDN U4557 ( .A(xregN_1), .B(zin[54]), .Z(n3041) );
  NAND U4558 ( .A(N59), .B(xregN_1), .Z(n3040) );
  NAND U4559 ( .A(n3042), .B(n3043), .Z(z2[559]) );
  NANDN U4560 ( .A(xregN_1), .B(zin[558]), .Z(n3043) );
  NAND U4561 ( .A(N563), .B(xregN_1), .Z(n3042) );
  NAND U4562 ( .A(n3044), .B(n3045), .Z(z2[558]) );
  NANDN U4563 ( .A(xregN_1), .B(zin[557]), .Z(n3045) );
  NAND U4564 ( .A(N562), .B(xregN_1), .Z(n3044) );
  NAND U4565 ( .A(n3046), .B(n3047), .Z(z2[557]) );
  NANDN U4566 ( .A(xregN_1), .B(zin[556]), .Z(n3047) );
  NAND U4567 ( .A(N561), .B(xregN_1), .Z(n3046) );
  NAND U4568 ( .A(n3048), .B(n3049), .Z(z2[556]) );
  NANDN U4569 ( .A(xregN_1), .B(zin[555]), .Z(n3049) );
  NAND U4570 ( .A(N560), .B(xregN_1), .Z(n3048) );
  NAND U4571 ( .A(n3050), .B(n3051), .Z(z2[555]) );
  NANDN U4572 ( .A(xregN_1), .B(zin[554]), .Z(n3051) );
  NAND U4573 ( .A(N559), .B(xregN_1), .Z(n3050) );
  NAND U4574 ( .A(n3052), .B(n3053), .Z(z2[554]) );
  NANDN U4575 ( .A(xregN_1), .B(zin[553]), .Z(n3053) );
  NAND U4576 ( .A(N558), .B(xregN_1), .Z(n3052) );
  NAND U4577 ( .A(n3054), .B(n3055), .Z(z2[553]) );
  NANDN U4578 ( .A(xregN_1), .B(zin[552]), .Z(n3055) );
  NAND U4579 ( .A(N557), .B(xregN_1), .Z(n3054) );
  NAND U4580 ( .A(n3056), .B(n3057), .Z(z2[552]) );
  NANDN U4581 ( .A(xregN_1), .B(zin[551]), .Z(n3057) );
  NAND U4582 ( .A(N556), .B(xregN_1), .Z(n3056) );
  NAND U4583 ( .A(n3058), .B(n3059), .Z(z2[551]) );
  NANDN U4584 ( .A(xregN_1), .B(zin[550]), .Z(n3059) );
  NAND U4585 ( .A(N555), .B(xregN_1), .Z(n3058) );
  NAND U4586 ( .A(n3060), .B(n3061), .Z(z2[550]) );
  NANDN U4587 ( .A(xregN_1), .B(zin[549]), .Z(n3061) );
  NAND U4588 ( .A(N554), .B(xregN_1), .Z(n3060) );
  NAND U4589 ( .A(n3062), .B(n3063), .Z(z2[54]) );
  NANDN U4590 ( .A(xregN_1), .B(zin[53]), .Z(n3063) );
  NAND U4591 ( .A(N58), .B(xregN_1), .Z(n3062) );
  NAND U4592 ( .A(n3064), .B(n3065), .Z(z2[549]) );
  NANDN U4593 ( .A(xregN_1), .B(zin[548]), .Z(n3065) );
  NAND U4594 ( .A(N553), .B(xregN_1), .Z(n3064) );
  NAND U4595 ( .A(n3066), .B(n3067), .Z(z2[548]) );
  NANDN U4596 ( .A(xregN_1), .B(zin[547]), .Z(n3067) );
  NAND U4597 ( .A(N552), .B(xregN_1), .Z(n3066) );
  NAND U4598 ( .A(n3068), .B(n3069), .Z(z2[547]) );
  NANDN U4599 ( .A(xregN_1), .B(zin[546]), .Z(n3069) );
  NAND U4600 ( .A(N551), .B(xregN_1), .Z(n3068) );
  NAND U4601 ( .A(n3070), .B(n3071), .Z(z2[546]) );
  NANDN U4602 ( .A(xregN_1), .B(zin[545]), .Z(n3071) );
  NAND U4603 ( .A(N550), .B(xregN_1), .Z(n3070) );
  NAND U4604 ( .A(n3072), .B(n3073), .Z(z2[545]) );
  NANDN U4605 ( .A(xregN_1), .B(zin[544]), .Z(n3073) );
  NAND U4606 ( .A(N549), .B(xregN_1), .Z(n3072) );
  NAND U4607 ( .A(n3074), .B(n3075), .Z(z2[544]) );
  NANDN U4608 ( .A(xregN_1), .B(zin[543]), .Z(n3075) );
  NAND U4609 ( .A(N548), .B(xregN_1), .Z(n3074) );
  NAND U4610 ( .A(n3076), .B(n3077), .Z(z2[543]) );
  NANDN U4611 ( .A(xregN_1), .B(zin[542]), .Z(n3077) );
  NAND U4612 ( .A(N547), .B(xregN_1), .Z(n3076) );
  NAND U4613 ( .A(n3078), .B(n3079), .Z(z2[542]) );
  NANDN U4614 ( .A(xregN_1), .B(zin[541]), .Z(n3079) );
  NAND U4615 ( .A(N546), .B(xregN_1), .Z(n3078) );
  NAND U4616 ( .A(n3080), .B(n3081), .Z(z2[541]) );
  NANDN U4617 ( .A(xregN_1), .B(zin[540]), .Z(n3081) );
  NAND U4618 ( .A(N545), .B(xregN_1), .Z(n3080) );
  NAND U4619 ( .A(n3082), .B(n3083), .Z(z2[540]) );
  NANDN U4620 ( .A(xregN_1), .B(zin[539]), .Z(n3083) );
  NAND U4621 ( .A(N544), .B(xregN_1), .Z(n3082) );
  NAND U4622 ( .A(n3084), .B(n3085), .Z(z2[53]) );
  NANDN U4623 ( .A(xregN_1), .B(zin[52]), .Z(n3085) );
  NAND U4624 ( .A(N57), .B(xregN_1), .Z(n3084) );
  NAND U4625 ( .A(n3086), .B(n3087), .Z(z2[539]) );
  NANDN U4626 ( .A(xregN_1), .B(zin[538]), .Z(n3087) );
  NAND U4627 ( .A(N543), .B(xregN_1), .Z(n3086) );
  NAND U4628 ( .A(n3088), .B(n3089), .Z(z2[538]) );
  NANDN U4629 ( .A(xregN_1), .B(zin[537]), .Z(n3089) );
  NAND U4630 ( .A(N542), .B(xregN_1), .Z(n3088) );
  NAND U4631 ( .A(n3090), .B(n3091), .Z(z2[537]) );
  NANDN U4632 ( .A(xregN_1), .B(zin[536]), .Z(n3091) );
  NAND U4633 ( .A(N541), .B(xregN_1), .Z(n3090) );
  NAND U4634 ( .A(n3092), .B(n3093), .Z(z2[536]) );
  NANDN U4635 ( .A(xregN_1), .B(zin[535]), .Z(n3093) );
  NAND U4636 ( .A(N540), .B(xregN_1), .Z(n3092) );
  NAND U4637 ( .A(n3094), .B(n3095), .Z(z2[535]) );
  NANDN U4638 ( .A(xregN_1), .B(zin[534]), .Z(n3095) );
  NAND U4639 ( .A(N539), .B(xregN_1), .Z(n3094) );
  NAND U4640 ( .A(n3096), .B(n3097), .Z(z2[534]) );
  NANDN U4641 ( .A(xregN_1), .B(zin[533]), .Z(n3097) );
  NAND U4642 ( .A(N538), .B(xregN_1), .Z(n3096) );
  NAND U4643 ( .A(n3098), .B(n3099), .Z(z2[533]) );
  NANDN U4644 ( .A(xregN_1), .B(zin[532]), .Z(n3099) );
  NAND U4645 ( .A(N537), .B(xregN_1), .Z(n3098) );
  NAND U4646 ( .A(n3100), .B(n3101), .Z(z2[532]) );
  NANDN U4647 ( .A(xregN_1), .B(zin[531]), .Z(n3101) );
  NAND U4648 ( .A(N536), .B(xregN_1), .Z(n3100) );
  NAND U4649 ( .A(n3102), .B(n3103), .Z(z2[531]) );
  NANDN U4650 ( .A(xregN_1), .B(zin[530]), .Z(n3103) );
  NAND U4651 ( .A(N535), .B(xregN_1), .Z(n3102) );
  NAND U4652 ( .A(n3104), .B(n3105), .Z(z2[530]) );
  NANDN U4653 ( .A(xregN_1), .B(zin[529]), .Z(n3105) );
  NAND U4654 ( .A(N534), .B(xregN_1), .Z(n3104) );
  NAND U4655 ( .A(n3106), .B(n3107), .Z(z2[52]) );
  NANDN U4656 ( .A(xregN_1), .B(zin[51]), .Z(n3107) );
  NAND U4657 ( .A(N56), .B(xregN_1), .Z(n3106) );
  NAND U4658 ( .A(n3108), .B(n3109), .Z(z2[529]) );
  NANDN U4659 ( .A(xregN_1), .B(zin[528]), .Z(n3109) );
  NAND U4660 ( .A(N533), .B(xregN_1), .Z(n3108) );
  NAND U4661 ( .A(n3110), .B(n3111), .Z(z2[528]) );
  NANDN U4662 ( .A(xregN_1), .B(zin[527]), .Z(n3111) );
  NAND U4663 ( .A(N532), .B(xregN_1), .Z(n3110) );
  NAND U4664 ( .A(n3112), .B(n3113), .Z(z2[527]) );
  NANDN U4665 ( .A(xregN_1), .B(zin[526]), .Z(n3113) );
  NAND U4666 ( .A(N531), .B(xregN_1), .Z(n3112) );
  NAND U4667 ( .A(n3114), .B(n3115), .Z(z2[526]) );
  NANDN U4668 ( .A(xregN_1), .B(zin[525]), .Z(n3115) );
  NAND U4669 ( .A(N530), .B(xregN_1), .Z(n3114) );
  NAND U4670 ( .A(n3116), .B(n3117), .Z(z2[525]) );
  NANDN U4671 ( .A(xregN_1), .B(zin[524]), .Z(n3117) );
  NAND U4672 ( .A(N529), .B(xregN_1), .Z(n3116) );
  NAND U4673 ( .A(n3118), .B(n3119), .Z(z2[524]) );
  NANDN U4674 ( .A(xregN_1), .B(zin[523]), .Z(n3119) );
  NAND U4675 ( .A(N528), .B(xregN_1), .Z(n3118) );
  NAND U4676 ( .A(n3120), .B(n3121), .Z(z2[523]) );
  NANDN U4677 ( .A(xregN_1), .B(zin[522]), .Z(n3121) );
  NAND U4678 ( .A(N527), .B(xregN_1), .Z(n3120) );
  NAND U4679 ( .A(n3122), .B(n3123), .Z(z2[522]) );
  NANDN U4680 ( .A(xregN_1), .B(zin[521]), .Z(n3123) );
  NAND U4681 ( .A(N526), .B(xregN_1), .Z(n3122) );
  NAND U4682 ( .A(n3124), .B(n3125), .Z(z2[521]) );
  NANDN U4683 ( .A(xregN_1), .B(zin[520]), .Z(n3125) );
  NAND U4684 ( .A(N525), .B(xregN_1), .Z(n3124) );
  NAND U4685 ( .A(n3126), .B(n3127), .Z(z2[520]) );
  NANDN U4686 ( .A(xregN_1), .B(zin[519]), .Z(n3127) );
  NAND U4687 ( .A(N524), .B(xregN_1), .Z(n3126) );
  NAND U4688 ( .A(n3128), .B(n3129), .Z(z2[51]) );
  NANDN U4689 ( .A(xregN_1), .B(zin[50]), .Z(n3129) );
  NAND U4690 ( .A(N55), .B(xregN_1), .Z(n3128) );
  NAND U4691 ( .A(n3130), .B(n3131), .Z(z2[519]) );
  NANDN U4692 ( .A(xregN_1), .B(zin[518]), .Z(n3131) );
  NAND U4693 ( .A(N523), .B(xregN_1), .Z(n3130) );
  NAND U4694 ( .A(n3132), .B(n3133), .Z(z2[518]) );
  NANDN U4695 ( .A(xregN_1), .B(zin[517]), .Z(n3133) );
  NAND U4696 ( .A(N522), .B(xregN_1), .Z(n3132) );
  NAND U4697 ( .A(n3134), .B(n3135), .Z(z2[517]) );
  NANDN U4698 ( .A(xregN_1), .B(zin[516]), .Z(n3135) );
  NAND U4699 ( .A(N521), .B(xregN_1), .Z(n3134) );
  NAND U4700 ( .A(n3136), .B(n3137), .Z(z2[516]) );
  NANDN U4701 ( .A(xregN_1), .B(zin[515]), .Z(n3137) );
  NAND U4702 ( .A(N520), .B(xregN_1), .Z(n3136) );
  NAND U4703 ( .A(n3138), .B(n3139), .Z(z2[515]) );
  NANDN U4704 ( .A(xregN_1), .B(zin[514]), .Z(n3139) );
  NAND U4705 ( .A(N519), .B(xregN_1), .Z(n3138) );
  NAND U4706 ( .A(n3140), .B(n3141), .Z(z2[514]) );
  NANDN U4707 ( .A(xregN_1), .B(zin[513]), .Z(n3141) );
  NAND U4708 ( .A(N518), .B(xregN_1), .Z(n3140) );
  NAND U4709 ( .A(n3142), .B(n3143), .Z(z2[513]) );
  NANDN U4710 ( .A(xregN_1), .B(zin[512]), .Z(n3143) );
  NAND U4711 ( .A(N517), .B(xregN_1), .Z(n3142) );
  NAND U4712 ( .A(n3144), .B(n3145), .Z(z2[512]) );
  NANDN U4713 ( .A(xregN_1), .B(zin[511]), .Z(n3145) );
  NAND U4714 ( .A(N516), .B(xregN_1), .Z(n3144) );
  NAND U4715 ( .A(n3146), .B(n3147), .Z(z2[511]) );
  NANDN U4716 ( .A(xregN_1), .B(zin[510]), .Z(n3147) );
  NAND U4717 ( .A(N515), .B(xregN_1), .Z(n3146) );
  NAND U4718 ( .A(n3148), .B(n3149), .Z(z2[510]) );
  NANDN U4719 ( .A(xregN_1), .B(zin[509]), .Z(n3149) );
  NAND U4720 ( .A(N514), .B(xregN_1), .Z(n3148) );
  NAND U4721 ( .A(n3150), .B(n3151), .Z(z2[50]) );
  NANDN U4722 ( .A(xregN_1), .B(zin[49]), .Z(n3151) );
  NAND U4723 ( .A(N54), .B(xregN_1), .Z(n3150) );
  NAND U4724 ( .A(n3152), .B(n3153), .Z(z2[509]) );
  NANDN U4725 ( .A(xregN_1), .B(zin[508]), .Z(n3153) );
  NAND U4726 ( .A(N513), .B(xregN_1), .Z(n3152) );
  NAND U4727 ( .A(n3154), .B(n3155), .Z(z2[508]) );
  NANDN U4728 ( .A(xregN_1), .B(zin[507]), .Z(n3155) );
  NAND U4729 ( .A(N512), .B(xregN_1), .Z(n3154) );
  NAND U4730 ( .A(n3156), .B(n3157), .Z(z2[507]) );
  NANDN U4731 ( .A(xregN_1), .B(zin[506]), .Z(n3157) );
  NAND U4732 ( .A(N511), .B(xregN_1), .Z(n3156) );
  NAND U4733 ( .A(n3158), .B(n3159), .Z(z2[506]) );
  NANDN U4734 ( .A(xregN_1), .B(zin[505]), .Z(n3159) );
  NAND U4735 ( .A(N510), .B(xregN_1), .Z(n3158) );
  NAND U4736 ( .A(n3160), .B(n3161), .Z(z2[505]) );
  NANDN U4737 ( .A(xregN_1), .B(zin[504]), .Z(n3161) );
  NAND U4738 ( .A(N509), .B(xregN_1), .Z(n3160) );
  NAND U4739 ( .A(n3162), .B(n3163), .Z(z2[504]) );
  NANDN U4740 ( .A(xregN_1), .B(zin[503]), .Z(n3163) );
  NAND U4741 ( .A(N508), .B(xregN_1), .Z(n3162) );
  NAND U4742 ( .A(n3164), .B(n3165), .Z(z2[503]) );
  NANDN U4743 ( .A(xregN_1), .B(zin[502]), .Z(n3165) );
  NAND U4744 ( .A(N507), .B(xregN_1), .Z(n3164) );
  NAND U4745 ( .A(n3166), .B(n3167), .Z(z2[502]) );
  NANDN U4746 ( .A(xregN_1), .B(zin[501]), .Z(n3167) );
  NAND U4747 ( .A(N506), .B(xregN_1), .Z(n3166) );
  NAND U4748 ( .A(n3168), .B(n3169), .Z(z2[501]) );
  NANDN U4749 ( .A(xregN_1), .B(zin[500]), .Z(n3169) );
  NAND U4750 ( .A(N505), .B(xregN_1), .Z(n3168) );
  NAND U4751 ( .A(n3170), .B(n3171), .Z(z2[500]) );
  NANDN U4752 ( .A(xregN_1), .B(zin[499]), .Z(n3171) );
  NAND U4753 ( .A(N504), .B(xregN_1), .Z(n3170) );
  NAND U4754 ( .A(n3172), .B(n3173), .Z(z2[4]) );
  NANDN U4755 ( .A(xregN_1), .B(zin[3]), .Z(n3173) );
  NAND U4756 ( .A(N8), .B(xregN_1), .Z(n3172) );
  NAND U4757 ( .A(n3174), .B(n3175), .Z(z2[49]) );
  NANDN U4758 ( .A(xregN_1), .B(zin[48]), .Z(n3175) );
  NAND U4759 ( .A(N53), .B(xregN_1), .Z(n3174) );
  NAND U4760 ( .A(n3176), .B(n3177), .Z(z2[499]) );
  NANDN U4761 ( .A(xregN_1), .B(zin[498]), .Z(n3177) );
  NAND U4762 ( .A(N503), .B(xregN_1), .Z(n3176) );
  NAND U4763 ( .A(n3178), .B(n3179), .Z(z2[498]) );
  NANDN U4764 ( .A(xregN_1), .B(zin[497]), .Z(n3179) );
  NAND U4765 ( .A(N502), .B(xregN_1), .Z(n3178) );
  NAND U4766 ( .A(n3180), .B(n3181), .Z(z2[497]) );
  NANDN U4767 ( .A(xregN_1), .B(zin[496]), .Z(n3181) );
  NAND U4768 ( .A(N501), .B(xregN_1), .Z(n3180) );
  NAND U4769 ( .A(n3182), .B(n3183), .Z(z2[496]) );
  NANDN U4770 ( .A(xregN_1), .B(zin[495]), .Z(n3183) );
  NAND U4771 ( .A(N500), .B(xregN_1), .Z(n3182) );
  NAND U4772 ( .A(n3184), .B(n3185), .Z(z2[495]) );
  NANDN U4773 ( .A(xregN_1), .B(zin[494]), .Z(n3185) );
  NAND U4774 ( .A(N499), .B(xregN_1), .Z(n3184) );
  NAND U4775 ( .A(n3186), .B(n3187), .Z(z2[494]) );
  NANDN U4776 ( .A(xregN_1), .B(zin[493]), .Z(n3187) );
  NAND U4777 ( .A(N498), .B(xregN_1), .Z(n3186) );
  NAND U4778 ( .A(n3188), .B(n3189), .Z(z2[493]) );
  NANDN U4779 ( .A(xregN_1), .B(zin[492]), .Z(n3189) );
  NAND U4780 ( .A(N497), .B(xregN_1), .Z(n3188) );
  NAND U4781 ( .A(n3190), .B(n3191), .Z(z2[492]) );
  NANDN U4782 ( .A(xregN_1), .B(zin[491]), .Z(n3191) );
  NAND U4783 ( .A(N496), .B(xregN_1), .Z(n3190) );
  NAND U4784 ( .A(n3192), .B(n3193), .Z(z2[491]) );
  NANDN U4785 ( .A(xregN_1), .B(zin[490]), .Z(n3193) );
  NAND U4786 ( .A(N495), .B(xregN_1), .Z(n3192) );
  NAND U4787 ( .A(n3194), .B(n3195), .Z(z2[490]) );
  NANDN U4788 ( .A(xregN_1), .B(zin[489]), .Z(n3195) );
  NAND U4789 ( .A(N494), .B(xregN_1), .Z(n3194) );
  NAND U4790 ( .A(n3196), .B(n3197), .Z(z2[48]) );
  NANDN U4791 ( .A(xregN_1), .B(zin[47]), .Z(n3197) );
  NAND U4792 ( .A(N52), .B(xregN_1), .Z(n3196) );
  NAND U4793 ( .A(n3198), .B(n3199), .Z(z2[489]) );
  NANDN U4794 ( .A(xregN_1), .B(zin[488]), .Z(n3199) );
  NAND U4795 ( .A(N493), .B(xregN_1), .Z(n3198) );
  NAND U4796 ( .A(n3200), .B(n3201), .Z(z2[488]) );
  NANDN U4797 ( .A(xregN_1), .B(zin[487]), .Z(n3201) );
  NAND U4798 ( .A(N492), .B(xregN_1), .Z(n3200) );
  NAND U4799 ( .A(n3202), .B(n3203), .Z(z2[487]) );
  NANDN U4800 ( .A(xregN_1), .B(zin[486]), .Z(n3203) );
  NAND U4801 ( .A(N491), .B(xregN_1), .Z(n3202) );
  NAND U4802 ( .A(n3204), .B(n3205), .Z(z2[486]) );
  NANDN U4803 ( .A(xregN_1), .B(zin[485]), .Z(n3205) );
  NAND U4804 ( .A(N490), .B(xregN_1), .Z(n3204) );
  NAND U4805 ( .A(n3206), .B(n3207), .Z(z2[485]) );
  NANDN U4806 ( .A(xregN_1), .B(zin[484]), .Z(n3207) );
  NAND U4807 ( .A(N489), .B(xregN_1), .Z(n3206) );
  NAND U4808 ( .A(n3208), .B(n3209), .Z(z2[484]) );
  NANDN U4809 ( .A(xregN_1), .B(zin[483]), .Z(n3209) );
  NAND U4810 ( .A(N488), .B(xregN_1), .Z(n3208) );
  NAND U4811 ( .A(n3210), .B(n3211), .Z(z2[483]) );
  NANDN U4812 ( .A(xregN_1), .B(zin[482]), .Z(n3211) );
  NAND U4813 ( .A(N487), .B(xregN_1), .Z(n3210) );
  NAND U4814 ( .A(n3212), .B(n3213), .Z(z2[482]) );
  NANDN U4815 ( .A(xregN_1), .B(zin[481]), .Z(n3213) );
  NAND U4816 ( .A(N486), .B(xregN_1), .Z(n3212) );
  NAND U4817 ( .A(n3214), .B(n3215), .Z(z2[481]) );
  NANDN U4818 ( .A(xregN_1), .B(zin[480]), .Z(n3215) );
  NAND U4819 ( .A(N485), .B(xregN_1), .Z(n3214) );
  NAND U4820 ( .A(n3216), .B(n3217), .Z(z2[480]) );
  NANDN U4821 ( .A(xregN_1), .B(zin[479]), .Z(n3217) );
  NAND U4822 ( .A(N484), .B(xregN_1), .Z(n3216) );
  NAND U4823 ( .A(n3218), .B(n3219), .Z(z2[47]) );
  NANDN U4824 ( .A(xregN_1), .B(zin[46]), .Z(n3219) );
  NAND U4825 ( .A(N51), .B(xregN_1), .Z(n3218) );
  NAND U4826 ( .A(n3220), .B(n3221), .Z(z2[479]) );
  NANDN U4827 ( .A(xregN_1), .B(zin[478]), .Z(n3221) );
  NAND U4828 ( .A(N483), .B(xregN_1), .Z(n3220) );
  NAND U4829 ( .A(n3222), .B(n3223), .Z(z2[478]) );
  NANDN U4830 ( .A(xregN_1), .B(zin[477]), .Z(n3223) );
  NAND U4831 ( .A(N482), .B(xregN_1), .Z(n3222) );
  NAND U4832 ( .A(n3224), .B(n3225), .Z(z2[477]) );
  NANDN U4833 ( .A(xregN_1), .B(zin[476]), .Z(n3225) );
  NAND U4834 ( .A(N481), .B(xregN_1), .Z(n3224) );
  NAND U4835 ( .A(n3226), .B(n3227), .Z(z2[476]) );
  NANDN U4836 ( .A(xregN_1), .B(zin[475]), .Z(n3227) );
  NAND U4837 ( .A(N480), .B(xregN_1), .Z(n3226) );
  NAND U4838 ( .A(n3228), .B(n3229), .Z(z2[475]) );
  NANDN U4839 ( .A(xregN_1), .B(zin[474]), .Z(n3229) );
  NAND U4840 ( .A(N479), .B(xregN_1), .Z(n3228) );
  NAND U4841 ( .A(n3230), .B(n3231), .Z(z2[474]) );
  NANDN U4842 ( .A(xregN_1), .B(zin[473]), .Z(n3231) );
  NAND U4843 ( .A(N478), .B(xregN_1), .Z(n3230) );
  NAND U4844 ( .A(n3232), .B(n3233), .Z(z2[473]) );
  NANDN U4845 ( .A(xregN_1), .B(zin[472]), .Z(n3233) );
  NAND U4846 ( .A(N477), .B(xregN_1), .Z(n3232) );
  NAND U4847 ( .A(n3234), .B(n3235), .Z(z2[472]) );
  NANDN U4848 ( .A(xregN_1), .B(zin[471]), .Z(n3235) );
  NAND U4849 ( .A(N476), .B(xregN_1), .Z(n3234) );
  NAND U4850 ( .A(n3236), .B(n3237), .Z(z2[471]) );
  NANDN U4851 ( .A(xregN_1), .B(zin[470]), .Z(n3237) );
  NAND U4852 ( .A(N475), .B(xregN_1), .Z(n3236) );
  NAND U4853 ( .A(n3238), .B(n3239), .Z(z2[470]) );
  NANDN U4854 ( .A(xregN_1), .B(zin[469]), .Z(n3239) );
  NAND U4855 ( .A(N474), .B(xregN_1), .Z(n3238) );
  NAND U4856 ( .A(n3240), .B(n3241), .Z(z2[46]) );
  NANDN U4857 ( .A(xregN_1), .B(zin[45]), .Z(n3241) );
  NAND U4858 ( .A(N50), .B(xregN_1), .Z(n3240) );
  NAND U4859 ( .A(n3242), .B(n3243), .Z(z2[469]) );
  NANDN U4860 ( .A(xregN_1), .B(zin[468]), .Z(n3243) );
  NAND U4861 ( .A(N473), .B(xregN_1), .Z(n3242) );
  NAND U4862 ( .A(n3244), .B(n3245), .Z(z2[468]) );
  NANDN U4863 ( .A(xregN_1), .B(zin[467]), .Z(n3245) );
  NAND U4864 ( .A(N472), .B(xregN_1), .Z(n3244) );
  NAND U4865 ( .A(n3246), .B(n3247), .Z(z2[467]) );
  NANDN U4866 ( .A(xregN_1), .B(zin[466]), .Z(n3247) );
  NAND U4867 ( .A(N471), .B(xregN_1), .Z(n3246) );
  NAND U4868 ( .A(n3248), .B(n3249), .Z(z2[466]) );
  NANDN U4869 ( .A(xregN_1), .B(zin[465]), .Z(n3249) );
  NAND U4870 ( .A(N470), .B(xregN_1), .Z(n3248) );
  NAND U4871 ( .A(n3250), .B(n3251), .Z(z2[465]) );
  NANDN U4872 ( .A(xregN_1), .B(zin[464]), .Z(n3251) );
  NAND U4873 ( .A(N469), .B(xregN_1), .Z(n3250) );
  NAND U4874 ( .A(n3252), .B(n3253), .Z(z2[464]) );
  NANDN U4875 ( .A(xregN_1), .B(zin[463]), .Z(n3253) );
  NAND U4876 ( .A(N468), .B(xregN_1), .Z(n3252) );
  NAND U4877 ( .A(n3254), .B(n3255), .Z(z2[463]) );
  NANDN U4878 ( .A(xregN_1), .B(zin[462]), .Z(n3255) );
  NAND U4879 ( .A(N467), .B(xregN_1), .Z(n3254) );
  NAND U4880 ( .A(n3256), .B(n3257), .Z(z2[462]) );
  NANDN U4881 ( .A(xregN_1), .B(zin[461]), .Z(n3257) );
  NAND U4882 ( .A(N466), .B(xregN_1), .Z(n3256) );
  NAND U4883 ( .A(n3258), .B(n3259), .Z(z2[461]) );
  NANDN U4884 ( .A(xregN_1), .B(zin[460]), .Z(n3259) );
  NAND U4885 ( .A(N465), .B(xregN_1), .Z(n3258) );
  NAND U4886 ( .A(n3260), .B(n3261), .Z(z2[460]) );
  NANDN U4887 ( .A(xregN_1), .B(zin[459]), .Z(n3261) );
  NAND U4888 ( .A(N464), .B(xregN_1), .Z(n3260) );
  NAND U4889 ( .A(n3262), .B(n3263), .Z(z2[45]) );
  NANDN U4890 ( .A(xregN_1), .B(zin[44]), .Z(n3263) );
  NAND U4891 ( .A(N49), .B(xregN_1), .Z(n3262) );
  NAND U4892 ( .A(n3264), .B(n3265), .Z(z2[459]) );
  NANDN U4893 ( .A(xregN_1), .B(zin[458]), .Z(n3265) );
  NAND U4894 ( .A(N463), .B(xregN_1), .Z(n3264) );
  NAND U4895 ( .A(n3266), .B(n3267), .Z(z2[458]) );
  NANDN U4896 ( .A(xregN_1), .B(zin[457]), .Z(n3267) );
  NAND U4897 ( .A(N462), .B(xregN_1), .Z(n3266) );
  NAND U4898 ( .A(n3268), .B(n3269), .Z(z2[457]) );
  NANDN U4899 ( .A(xregN_1), .B(zin[456]), .Z(n3269) );
  NAND U4900 ( .A(N461), .B(xregN_1), .Z(n3268) );
  NAND U4901 ( .A(n3270), .B(n3271), .Z(z2[456]) );
  NANDN U4902 ( .A(xregN_1), .B(zin[455]), .Z(n3271) );
  NAND U4903 ( .A(N460), .B(xregN_1), .Z(n3270) );
  NAND U4904 ( .A(n3272), .B(n3273), .Z(z2[455]) );
  NANDN U4905 ( .A(xregN_1), .B(zin[454]), .Z(n3273) );
  NAND U4906 ( .A(N459), .B(xregN_1), .Z(n3272) );
  NAND U4907 ( .A(n3274), .B(n3275), .Z(z2[454]) );
  NANDN U4908 ( .A(xregN_1), .B(zin[453]), .Z(n3275) );
  NAND U4909 ( .A(N458), .B(xregN_1), .Z(n3274) );
  NAND U4910 ( .A(n3276), .B(n3277), .Z(z2[453]) );
  NANDN U4911 ( .A(xregN_1), .B(zin[452]), .Z(n3277) );
  NAND U4912 ( .A(N457), .B(xregN_1), .Z(n3276) );
  NAND U4913 ( .A(n3278), .B(n3279), .Z(z2[452]) );
  NANDN U4914 ( .A(xregN_1), .B(zin[451]), .Z(n3279) );
  NAND U4915 ( .A(N456), .B(xregN_1), .Z(n3278) );
  NAND U4916 ( .A(n3280), .B(n3281), .Z(z2[451]) );
  NANDN U4917 ( .A(xregN_1), .B(zin[450]), .Z(n3281) );
  NAND U4918 ( .A(N455), .B(xregN_1), .Z(n3280) );
  NAND U4919 ( .A(n3282), .B(n3283), .Z(z2[450]) );
  NANDN U4920 ( .A(xregN_1), .B(zin[449]), .Z(n3283) );
  NAND U4921 ( .A(N454), .B(xregN_1), .Z(n3282) );
  NAND U4922 ( .A(n3284), .B(n3285), .Z(z2[44]) );
  NANDN U4923 ( .A(xregN_1), .B(zin[43]), .Z(n3285) );
  NAND U4924 ( .A(N48), .B(xregN_1), .Z(n3284) );
  NAND U4925 ( .A(n3286), .B(n3287), .Z(z2[449]) );
  NANDN U4926 ( .A(xregN_1), .B(zin[448]), .Z(n3287) );
  NAND U4927 ( .A(N453), .B(xregN_1), .Z(n3286) );
  NAND U4928 ( .A(n3288), .B(n3289), .Z(z2[448]) );
  NANDN U4929 ( .A(xregN_1), .B(zin[447]), .Z(n3289) );
  NAND U4930 ( .A(N452), .B(xregN_1), .Z(n3288) );
  NAND U4931 ( .A(n3290), .B(n3291), .Z(z2[447]) );
  NANDN U4932 ( .A(xregN_1), .B(zin[446]), .Z(n3291) );
  NAND U4933 ( .A(N451), .B(xregN_1), .Z(n3290) );
  NAND U4934 ( .A(n3292), .B(n3293), .Z(z2[446]) );
  NANDN U4935 ( .A(xregN_1), .B(zin[445]), .Z(n3293) );
  NAND U4936 ( .A(N450), .B(xregN_1), .Z(n3292) );
  NAND U4937 ( .A(n3294), .B(n3295), .Z(z2[445]) );
  NANDN U4938 ( .A(xregN_1), .B(zin[444]), .Z(n3295) );
  NAND U4939 ( .A(N449), .B(xregN_1), .Z(n3294) );
  NAND U4940 ( .A(n3296), .B(n3297), .Z(z2[444]) );
  NANDN U4941 ( .A(xregN_1), .B(zin[443]), .Z(n3297) );
  NAND U4942 ( .A(N448), .B(xregN_1), .Z(n3296) );
  NAND U4943 ( .A(n3298), .B(n3299), .Z(z2[443]) );
  NANDN U4944 ( .A(xregN_1), .B(zin[442]), .Z(n3299) );
  NAND U4945 ( .A(N447), .B(xregN_1), .Z(n3298) );
  NAND U4946 ( .A(n3300), .B(n3301), .Z(z2[442]) );
  NANDN U4947 ( .A(xregN_1), .B(zin[441]), .Z(n3301) );
  NAND U4948 ( .A(N446), .B(xregN_1), .Z(n3300) );
  NAND U4949 ( .A(n3302), .B(n3303), .Z(z2[441]) );
  NANDN U4950 ( .A(xregN_1), .B(zin[440]), .Z(n3303) );
  NAND U4951 ( .A(N445), .B(xregN_1), .Z(n3302) );
  NAND U4952 ( .A(n3304), .B(n3305), .Z(z2[440]) );
  NANDN U4953 ( .A(xregN_1), .B(zin[439]), .Z(n3305) );
  NAND U4954 ( .A(N444), .B(xregN_1), .Z(n3304) );
  NAND U4955 ( .A(n3306), .B(n3307), .Z(z2[43]) );
  NANDN U4956 ( .A(xregN_1), .B(zin[42]), .Z(n3307) );
  NAND U4957 ( .A(N47), .B(xregN_1), .Z(n3306) );
  NAND U4958 ( .A(n3308), .B(n3309), .Z(z2[439]) );
  NANDN U4959 ( .A(xregN_1), .B(zin[438]), .Z(n3309) );
  NAND U4960 ( .A(N443), .B(xregN_1), .Z(n3308) );
  NAND U4961 ( .A(n3310), .B(n3311), .Z(z2[438]) );
  NANDN U4962 ( .A(xregN_1), .B(zin[437]), .Z(n3311) );
  NAND U4963 ( .A(N442), .B(xregN_1), .Z(n3310) );
  NAND U4964 ( .A(n3312), .B(n3313), .Z(z2[437]) );
  NANDN U4965 ( .A(xregN_1), .B(zin[436]), .Z(n3313) );
  NAND U4966 ( .A(N441), .B(xregN_1), .Z(n3312) );
  NAND U4967 ( .A(n3314), .B(n3315), .Z(z2[436]) );
  NANDN U4968 ( .A(xregN_1), .B(zin[435]), .Z(n3315) );
  NAND U4969 ( .A(N440), .B(xregN_1), .Z(n3314) );
  NAND U4970 ( .A(n3316), .B(n3317), .Z(z2[435]) );
  NANDN U4971 ( .A(xregN_1), .B(zin[434]), .Z(n3317) );
  NAND U4972 ( .A(N439), .B(xregN_1), .Z(n3316) );
  NAND U4973 ( .A(n3318), .B(n3319), .Z(z2[434]) );
  NANDN U4974 ( .A(xregN_1), .B(zin[433]), .Z(n3319) );
  NAND U4975 ( .A(N438), .B(xregN_1), .Z(n3318) );
  NAND U4976 ( .A(n3320), .B(n3321), .Z(z2[433]) );
  NANDN U4977 ( .A(xregN_1), .B(zin[432]), .Z(n3321) );
  NAND U4978 ( .A(N437), .B(xregN_1), .Z(n3320) );
  NAND U4979 ( .A(n3322), .B(n3323), .Z(z2[432]) );
  NANDN U4980 ( .A(xregN_1), .B(zin[431]), .Z(n3323) );
  NAND U4981 ( .A(N436), .B(xregN_1), .Z(n3322) );
  NAND U4982 ( .A(n3324), .B(n3325), .Z(z2[431]) );
  NANDN U4983 ( .A(xregN_1), .B(zin[430]), .Z(n3325) );
  NAND U4984 ( .A(N435), .B(xregN_1), .Z(n3324) );
  NAND U4985 ( .A(n3326), .B(n3327), .Z(z2[430]) );
  NANDN U4986 ( .A(xregN_1), .B(zin[429]), .Z(n3327) );
  NAND U4987 ( .A(N434), .B(xregN_1), .Z(n3326) );
  NAND U4988 ( .A(n3328), .B(n3329), .Z(z2[42]) );
  NANDN U4989 ( .A(xregN_1), .B(zin[41]), .Z(n3329) );
  NAND U4990 ( .A(N46), .B(xregN_1), .Z(n3328) );
  NAND U4991 ( .A(n3330), .B(n3331), .Z(z2[429]) );
  NANDN U4992 ( .A(xregN_1), .B(zin[428]), .Z(n3331) );
  NAND U4993 ( .A(N433), .B(xregN_1), .Z(n3330) );
  NAND U4994 ( .A(n3332), .B(n3333), .Z(z2[428]) );
  NANDN U4995 ( .A(xregN_1), .B(zin[427]), .Z(n3333) );
  NAND U4996 ( .A(N432), .B(xregN_1), .Z(n3332) );
  NAND U4997 ( .A(n3334), .B(n3335), .Z(z2[427]) );
  NANDN U4998 ( .A(xregN_1), .B(zin[426]), .Z(n3335) );
  NAND U4999 ( .A(N431), .B(xregN_1), .Z(n3334) );
  NAND U5000 ( .A(n3336), .B(n3337), .Z(z2[426]) );
  NANDN U5001 ( .A(xregN_1), .B(zin[425]), .Z(n3337) );
  NAND U5002 ( .A(N430), .B(xregN_1), .Z(n3336) );
  NAND U5003 ( .A(n3338), .B(n3339), .Z(z2[425]) );
  NANDN U5004 ( .A(xregN_1), .B(zin[424]), .Z(n3339) );
  NAND U5005 ( .A(N429), .B(xregN_1), .Z(n3338) );
  NAND U5006 ( .A(n3340), .B(n3341), .Z(z2[424]) );
  NANDN U5007 ( .A(xregN_1), .B(zin[423]), .Z(n3341) );
  NAND U5008 ( .A(N428), .B(xregN_1), .Z(n3340) );
  NAND U5009 ( .A(n3342), .B(n3343), .Z(z2[423]) );
  NANDN U5010 ( .A(xregN_1), .B(zin[422]), .Z(n3343) );
  NAND U5011 ( .A(N427), .B(xregN_1), .Z(n3342) );
  NAND U5012 ( .A(n3344), .B(n3345), .Z(z2[422]) );
  NANDN U5013 ( .A(xregN_1), .B(zin[421]), .Z(n3345) );
  NAND U5014 ( .A(N426), .B(xregN_1), .Z(n3344) );
  NAND U5015 ( .A(n3346), .B(n3347), .Z(z2[421]) );
  NANDN U5016 ( .A(xregN_1), .B(zin[420]), .Z(n3347) );
  NAND U5017 ( .A(N425), .B(xregN_1), .Z(n3346) );
  NAND U5018 ( .A(n3348), .B(n3349), .Z(z2[420]) );
  NANDN U5019 ( .A(xregN_1), .B(zin[419]), .Z(n3349) );
  NAND U5020 ( .A(N424), .B(xregN_1), .Z(n3348) );
  NAND U5021 ( .A(n3350), .B(n3351), .Z(z2[41]) );
  NANDN U5022 ( .A(xregN_1), .B(zin[40]), .Z(n3351) );
  NAND U5023 ( .A(N45), .B(xregN_1), .Z(n3350) );
  NAND U5024 ( .A(n3352), .B(n3353), .Z(z2[419]) );
  NANDN U5025 ( .A(xregN_1), .B(zin[418]), .Z(n3353) );
  NAND U5026 ( .A(N423), .B(xregN_1), .Z(n3352) );
  NAND U5027 ( .A(n3354), .B(n3355), .Z(z2[418]) );
  NANDN U5028 ( .A(xregN_1), .B(zin[417]), .Z(n3355) );
  NAND U5029 ( .A(N422), .B(xregN_1), .Z(n3354) );
  NAND U5030 ( .A(n3356), .B(n3357), .Z(z2[417]) );
  NANDN U5031 ( .A(xregN_1), .B(zin[416]), .Z(n3357) );
  NAND U5032 ( .A(N421), .B(xregN_1), .Z(n3356) );
  NAND U5033 ( .A(n3358), .B(n3359), .Z(z2[416]) );
  NANDN U5034 ( .A(xregN_1), .B(zin[415]), .Z(n3359) );
  NAND U5035 ( .A(N420), .B(xregN_1), .Z(n3358) );
  NAND U5036 ( .A(n3360), .B(n3361), .Z(z2[415]) );
  NANDN U5037 ( .A(xregN_1), .B(zin[414]), .Z(n3361) );
  NAND U5038 ( .A(N419), .B(xregN_1), .Z(n3360) );
  NAND U5039 ( .A(n3362), .B(n3363), .Z(z2[414]) );
  NANDN U5040 ( .A(xregN_1), .B(zin[413]), .Z(n3363) );
  NAND U5041 ( .A(N418), .B(xregN_1), .Z(n3362) );
  NAND U5042 ( .A(n3364), .B(n3365), .Z(z2[413]) );
  NANDN U5043 ( .A(xregN_1), .B(zin[412]), .Z(n3365) );
  NAND U5044 ( .A(N417), .B(xregN_1), .Z(n3364) );
  NAND U5045 ( .A(n3366), .B(n3367), .Z(z2[412]) );
  NANDN U5046 ( .A(xregN_1), .B(zin[411]), .Z(n3367) );
  NAND U5047 ( .A(N416), .B(xregN_1), .Z(n3366) );
  NAND U5048 ( .A(n3368), .B(n3369), .Z(z2[411]) );
  NANDN U5049 ( .A(xregN_1), .B(zin[410]), .Z(n3369) );
  NAND U5050 ( .A(N415), .B(xregN_1), .Z(n3368) );
  NAND U5051 ( .A(n3370), .B(n3371), .Z(z2[410]) );
  NANDN U5052 ( .A(xregN_1), .B(zin[409]), .Z(n3371) );
  NAND U5053 ( .A(N414), .B(xregN_1), .Z(n3370) );
  NAND U5054 ( .A(n3372), .B(n3373), .Z(z2[40]) );
  NANDN U5055 ( .A(xregN_1), .B(zin[39]), .Z(n3373) );
  NAND U5056 ( .A(N44), .B(xregN_1), .Z(n3372) );
  NAND U5057 ( .A(n3374), .B(n3375), .Z(z2[409]) );
  NANDN U5058 ( .A(xregN_1), .B(zin[408]), .Z(n3375) );
  NAND U5059 ( .A(N413), .B(xregN_1), .Z(n3374) );
  NAND U5060 ( .A(n3376), .B(n3377), .Z(z2[408]) );
  NANDN U5061 ( .A(xregN_1), .B(zin[407]), .Z(n3377) );
  NAND U5062 ( .A(N412), .B(xregN_1), .Z(n3376) );
  NAND U5063 ( .A(n3378), .B(n3379), .Z(z2[407]) );
  NANDN U5064 ( .A(xregN_1), .B(zin[406]), .Z(n3379) );
  NAND U5065 ( .A(N411), .B(xregN_1), .Z(n3378) );
  NAND U5066 ( .A(n3380), .B(n3381), .Z(z2[406]) );
  NANDN U5067 ( .A(xregN_1), .B(zin[405]), .Z(n3381) );
  NAND U5068 ( .A(N410), .B(xregN_1), .Z(n3380) );
  NAND U5069 ( .A(n3382), .B(n3383), .Z(z2[405]) );
  NANDN U5070 ( .A(xregN_1), .B(zin[404]), .Z(n3383) );
  NAND U5071 ( .A(N409), .B(xregN_1), .Z(n3382) );
  NAND U5072 ( .A(n3384), .B(n3385), .Z(z2[404]) );
  NANDN U5073 ( .A(xregN_1), .B(zin[403]), .Z(n3385) );
  NAND U5074 ( .A(N408), .B(xregN_1), .Z(n3384) );
  NAND U5075 ( .A(n3386), .B(n3387), .Z(z2[403]) );
  NANDN U5076 ( .A(xregN_1), .B(zin[402]), .Z(n3387) );
  NAND U5077 ( .A(N407), .B(xregN_1), .Z(n3386) );
  NAND U5078 ( .A(n3388), .B(n3389), .Z(z2[402]) );
  NANDN U5079 ( .A(xregN_1), .B(zin[401]), .Z(n3389) );
  NAND U5080 ( .A(N406), .B(xregN_1), .Z(n3388) );
  NAND U5081 ( .A(n3390), .B(n3391), .Z(z2[401]) );
  NANDN U5082 ( .A(xregN_1), .B(zin[400]), .Z(n3391) );
  NAND U5083 ( .A(N405), .B(xregN_1), .Z(n3390) );
  NAND U5084 ( .A(n3392), .B(n3393), .Z(z2[400]) );
  NANDN U5085 ( .A(xregN_1), .B(zin[399]), .Z(n3393) );
  NAND U5086 ( .A(N404), .B(xregN_1), .Z(n3392) );
  NAND U5087 ( .A(n3394), .B(n3395), .Z(z2[3]) );
  NANDN U5088 ( .A(xregN_1), .B(zin[2]), .Z(n3395) );
  NAND U5089 ( .A(N7), .B(xregN_1), .Z(n3394) );
  NAND U5090 ( .A(n3396), .B(n3397), .Z(z2[39]) );
  NANDN U5091 ( .A(xregN_1), .B(zin[38]), .Z(n3397) );
  NAND U5092 ( .A(N43), .B(xregN_1), .Z(n3396) );
  NAND U5093 ( .A(n3398), .B(n3399), .Z(z2[399]) );
  NANDN U5094 ( .A(xregN_1), .B(zin[398]), .Z(n3399) );
  NAND U5095 ( .A(N403), .B(xregN_1), .Z(n3398) );
  NAND U5096 ( .A(n3400), .B(n3401), .Z(z2[398]) );
  NANDN U5097 ( .A(xregN_1), .B(zin[397]), .Z(n3401) );
  NAND U5098 ( .A(N402), .B(xregN_1), .Z(n3400) );
  NAND U5099 ( .A(n3402), .B(n3403), .Z(z2[397]) );
  NANDN U5100 ( .A(xregN_1), .B(zin[396]), .Z(n3403) );
  NAND U5101 ( .A(N401), .B(xregN_1), .Z(n3402) );
  NAND U5102 ( .A(n3404), .B(n3405), .Z(z2[396]) );
  NANDN U5103 ( .A(xregN_1), .B(zin[395]), .Z(n3405) );
  NAND U5104 ( .A(N400), .B(xregN_1), .Z(n3404) );
  NAND U5105 ( .A(n3406), .B(n3407), .Z(z2[395]) );
  NANDN U5106 ( .A(xregN_1), .B(zin[394]), .Z(n3407) );
  NAND U5107 ( .A(N399), .B(xregN_1), .Z(n3406) );
  NAND U5108 ( .A(n3408), .B(n3409), .Z(z2[394]) );
  NANDN U5109 ( .A(xregN_1), .B(zin[393]), .Z(n3409) );
  NAND U5110 ( .A(N398), .B(xregN_1), .Z(n3408) );
  NAND U5111 ( .A(n3410), .B(n3411), .Z(z2[393]) );
  NANDN U5112 ( .A(xregN_1), .B(zin[392]), .Z(n3411) );
  NAND U5113 ( .A(N397), .B(xregN_1), .Z(n3410) );
  NAND U5114 ( .A(n3412), .B(n3413), .Z(z2[392]) );
  NANDN U5115 ( .A(xregN_1), .B(zin[391]), .Z(n3413) );
  NAND U5116 ( .A(N396), .B(xregN_1), .Z(n3412) );
  NAND U5117 ( .A(n3414), .B(n3415), .Z(z2[391]) );
  NANDN U5118 ( .A(xregN_1), .B(zin[390]), .Z(n3415) );
  NAND U5119 ( .A(N395), .B(xregN_1), .Z(n3414) );
  NAND U5120 ( .A(n3416), .B(n3417), .Z(z2[390]) );
  NANDN U5121 ( .A(xregN_1), .B(zin[389]), .Z(n3417) );
  NAND U5122 ( .A(N394), .B(xregN_1), .Z(n3416) );
  NAND U5123 ( .A(n3418), .B(n3419), .Z(z2[38]) );
  NANDN U5124 ( .A(xregN_1), .B(zin[37]), .Z(n3419) );
  NAND U5125 ( .A(N42), .B(xregN_1), .Z(n3418) );
  NAND U5126 ( .A(n3420), .B(n3421), .Z(z2[389]) );
  NANDN U5127 ( .A(xregN_1), .B(zin[388]), .Z(n3421) );
  NAND U5128 ( .A(N393), .B(xregN_1), .Z(n3420) );
  NAND U5129 ( .A(n3422), .B(n3423), .Z(z2[388]) );
  NANDN U5130 ( .A(xregN_1), .B(zin[387]), .Z(n3423) );
  NAND U5131 ( .A(N392), .B(xregN_1), .Z(n3422) );
  NAND U5132 ( .A(n3424), .B(n3425), .Z(z2[387]) );
  NANDN U5133 ( .A(xregN_1), .B(zin[386]), .Z(n3425) );
  NAND U5134 ( .A(N391), .B(xregN_1), .Z(n3424) );
  NAND U5135 ( .A(n3426), .B(n3427), .Z(z2[386]) );
  NANDN U5136 ( .A(xregN_1), .B(zin[385]), .Z(n3427) );
  NAND U5137 ( .A(N390), .B(xregN_1), .Z(n3426) );
  NAND U5138 ( .A(n3428), .B(n3429), .Z(z2[385]) );
  NANDN U5139 ( .A(xregN_1), .B(zin[384]), .Z(n3429) );
  NAND U5140 ( .A(N389), .B(xregN_1), .Z(n3428) );
  NAND U5141 ( .A(n3430), .B(n3431), .Z(z2[384]) );
  NANDN U5142 ( .A(xregN_1), .B(zin[383]), .Z(n3431) );
  NAND U5143 ( .A(N388), .B(xregN_1), .Z(n3430) );
  NAND U5144 ( .A(n3432), .B(n3433), .Z(z2[383]) );
  NANDN U5145 ( .A(xregN_1), .B(zin[382]), .Z(n3433) );
  NAND U5146 ( .A(N387), .B(xregN_1), .Z(n3432) );
  NAND U5147 ( .A(n3434), .B(n3435), .Z(z2[382]) );
  NANDN U5148 ( .A(xregN_1), .B(zin[381]), .Z(n3435) );
  NAND U5149 ( .A(N386), .B(xregN_1), .Z(n3434) );
  NAND U5150 ( .A(n3436), .B(n3437), .Z(z2[381]) );
  NANDN U5151 ( .A(xregN_1), .B(zin[380]), .Z(n3437) );
  NAND U5152 ( .A(N385), .B(xregN_1), .Z(n3436) );
  NAND U5153 ( .A(n3438), .B(n3439), .Z(z2[380]) );
  NANDN U5154 ( .A(xregN_1), .B(zin[379]), .Z(n3439) );
  NAND U5155 ( .A(N384), .B(xregN_1), .Z(n3438) );
  NAND U5156 ( .A(n3440), .B(n3441), .Z(z2[37]) );
  NANDN U5157 ( .A(xregN_1), .B(zin[36]), .Z(n3441) );
  NAND U5158 ( .A(N41), .B(xregN_1), .Z(n3440) );
  NAND U5159 ( .A(n3442), .B(n3443), .Z(z2[379]) );
  NANDN U5160 ( .A(xregN_1), .B(zin[378]), .Z(n3443) );
  NAND U5161 ( .A(N383), .B(xregN_1), .Z(n3442) );
  NAND U5162 ( .A(n3444), .B(n3445), .Z(z2[378]) );
  NANDN U5163 ( .A(xregN_1), .B(zin[377]), .Z(n3445) );
  NAND U5164 ( .A(N382), .B(xregN_1), .Z(n3444) );
  NAND U5165 ( .A(n3446), .B(n3447), .Z(z2[377]) );
  NANDN U5166 ( .A(xregN_1), .B(zin[376]), .Z(n3447) );
  NAND U5167 ( .A(N381), .B(xregN_1), .Z(n3446) );
  NAND U5168 ( .A(n3448), .B(n3449), .Z(z2[376]) );
  NANDN U5169 ( .A(xregN_1), .B(zin[375]), .Z(n3449) );
  NAND U5170 ( .A(N380), .B(xregN_1), .Z(n3448) );
  NAND U5171 ( .A(n3450), .B(n3451), .Z(z2[375]) );
  NANDN U5172 ( .A(xregN_1), .B(zin[374]), .Z(n3451) );
  NAND U5173 ( .A(N379), .B(xregN_1), .Z(n3450) );
  NAND U5174 ( .A(n3452), .B(n3453), .Z(z2[374]) );
  NANDN U5175 ( .A(xregN_1), .B(zin[373]), .Z(n3453) );
  NAND U5176 ( .A(N378), .B(xregN_1), .Z(n3452) );
  NAND U5177 ( .A(n3454), .B(n3455), .Z(z2[373]) );
  NANDN U5178 ( .A(xregN_1), .B(zin[372]), .Z(n3455) );
  NAND U5179 ( .A(N377), .B(xregN_1), .Z(n3454) );
  NAND U5180 ( .A(n3456), .B(n3457), .Z(z2[372]) );
  NANDN U5181 ( .A(xregN_1), .B(zin[371]), .Z(n3457) );
  NAND U5182 ( .A(N376), .B(xregN_1), .Z(n3456) );
  NAND U5183 ( .A(n3458), .B(n3459), .Z(z2[371]) );
  NANDN U5184 ( .A(xregN_1), .B(zin[370]), .Z(n3459) );
  NAND U5185 ( .A(N375), .B(xregN_1), .Z(n3458) );
  NAND U5186 ( .A(n3460), .B(n3461), .Z(z2[370]) );
  NANDN U5187 ( .A(xregN_1), .B(zin[369]), .Z(n3461) );
  NAND U5188 ( .A(N374), .B(xregN_1), .Z(n3460) );
  NAND U5189 ( .A(n3462), .B(n3463), .Z(z2[36]) );
  NANDN U5190 ( .A(xregN_1), .B(zin[35]), .Z(n3463) );
  NAND U5191 ( .A(N40), .B(xregN_1), .Z(n3462) );
  NAND U5192 ( .A(n3464), .B(n3465), .Z(z2[369]) );
  NANDN U5193 ( .A(xregN_1), .B(zin[368]), .Z(n3465) );
  NAND U5194 ( .A(N373), .B(xregN_1), .Z(n3464) );
  NAND U5195 ( .A(n3466), .B(n3467), .Z(z2[368]) );
  NANDN U5196 ( .A(xregN_1), .B(zin[367]), .Z(n3467) );
  NAND U5197 ( .A(N372), .B(xregN_1), .Z(n3466) );
  NAND U5198 ( .A(n3468), .B(n3469), .Z(z2[367]) );
  NANDN U5199 ( .A(xregN_1), .B(zin[366]), .Z(n3469) );
  NAND U5200 ( .A(N371), .B(xregN_1), .Z(n3468) );
  NAND U5201 ( .A(n3470), .B(n3471), .Z(z2[366]) );
  NANDN U5202 ( .A(xregN_1), .B(zin[365]), .Z(n3471) );
  NAND U5203 ( .A(N370), .B(xregN_1), .Z(n3470) );
  NAND U5204 ( .A(n3472), .B(n3473), .Z(z2[365]) );
  NANDN U5205 ( .A(xregN_1), .B(zin[364]), .Z(n3473) );
  NAND U5206 ( .A(N369), .B(xregN_1), .Z(n3472) );
  NAND U5207 ( .A(n3474), .B(n3475), .Z(z2[364]) );
  NANDN U5208 ( .A(xregN_1), .B(zin[363]), .Z(n3475) );
  NAND U5209 ( .A(N368), .B(xregN_1), .Z(n3474) );
  NAND U5210 ( .A(n3476), .B(n3477), .Z(z2[363]) );
  NANDN U5211 ( .A(xregN_1), .B(zin[362]), .Z(n3477) );
  NAND U5212 ( .A(N367), .B(xregN_1), .Z(n3476) );
  NAND U5213 ( .A(n3478), .B(n3479), .Z(z2[362]) );
  NANDN U5214 ( .A(xregN_1), .B(zin[361]), .Z(n3479) );
  NAND U5215 ( .A(N366), .B(xregN_1), .Z(n3478) );
  NAND U5216 ( .A(n3480), .B(n3481), .Z(z2[361]) );
  NANDN U5217 ( .A(xregN_1), .B(zin[360]), .Z(n3481) );
  NAND U5218 ( .A(N365), .B(xregN_1), .Z(n3480) );
  NAND U5219 ( .A(n3482), .B(n3483), .Z(z2[360]) );
  NANDN U5220 ( .A(xregN_1), .B(zin[359]), .Z(n3483) );
  NAND U5221 ( .A(N364), .B(xregN_1), .Z(n3482) );
  NAND U5222 ( .A(n3484), .B(n3485), .Z(z2[35]) );
  NANDN U5223 ( .A(xregN_1), .B(zin[34]), .Z(n3485) );
  NAND U5224 ( .A(N39), .B(xregN_1), .Z(n3484) );
  NAND U5225 ( .A(n3486), .B(n3487), .Z(z2[359]) );
  NANDN U5226 ( .A(xregN_1), .B(zin[358]), .Z(n3487) );
  NAND U5227 ( .A(N363), .B(xregN_1), .Z(n3486) );
  NAND U5228 ( .A(n3488), .B(n3489), .Z(z2[358]) );
  NANDN U5229 ( .A(xregN_1), .B(zin[357]), .Z(n3489) );
  NAND U5230 ( .A(N362), .B(xregN_1), .Z(n3488) );
  NAND U5231 ( .A(n3490), .B(n3491), .Z(z2[357]) );
  NANDN U5232 ( .A(xregN_1), .B(zin[356]), .Z(n3491) );
  NAND U5233 ( .A(N361), .B(xregN_1), .Z(n3490) );
  NAND U5234 ( .A(n3492), .B(n3493), .Z(z2[356]) );
  NANDN U5235 ( .A(xregN_1), .B(zin[355]), .Z(n3493) );
  NAND U5236 ( .A(N360), .B(xregN_1), .Z(n3492) );
  NAND U5237 ( .A(n3494), .B(n3495), .Z(z2[355]) );
  NANDN U5238 ( .A(xregN_1), .B(zin[354]), .Z(n3495) );
  NAND U5239 ( .A(N359), .B(xregN_1), .Z(n3494) );
  NAND U5240 ( .A(n3496), .B(n3497), .Z(z2[354]) );
  NANDN U5241 ( .A(xregN_1), .B(zin[353]), .Z(n3497) );
  NAND U5242 ( .A(N358), .B(xregN_1), .Z(n3496) );
  NAND U5243 ( .A(n3498), .B(n3499), .Z(z2[353]) );
  NANDN U5244 ( .A(xregN_1), .B(zin[352]), .Z(n3499) );
  NAND U5245 ( .A(N357), .B(xregN_1), .Z(n3498) );
  NAND U5246 ( .A(n3500), .B(n3501), .Z(z2[352]) );
  NANDN U5247 ( .A(xregN_1), .B(zin[351]), .Z(n3501) );
  NAND U5248 ( .A(N356), .B(xregN_1), .Z(n3500) );
  NAND U5249 ( .A(n3502), .B(n3503), .Z(z2[351]) );
  NANDN U5250 ( .A(xregN_1), .B(zin[350]), .Z(n3503) );
  NAND U5251 ( .A(N355), .B(xregN_1), .Z(n3502) );
  NAND U5252 ( .A(n3504), .B(n3505), .Z(z2[350]) );
  NANDN U5253 ( .A(xregN_1), .B(zin[349]), .Z(n3505) );
  NAND U5254 ( .A(N354), .B(xregN_1), .Z(n3504) );
  NAND U5255 ( .A(n3506), .B(n3507), .Z(z2[34]) );
  NANDN U5256 ( .A(xregN_1), .B(zin[33]), .Z(n3507) );
  NAND U5257 ( .A(N38), .B(xregN_1), .Z(n3506) );
  NAND U5258 ( .A(n3508), .B(n3509), .Z(z2[349]) );
  NANDN U5259 ( .A(xregN_1), .B(zin[348]), .Z(n3509) );
  NAND U5260 ( .A(N353), .B(xregN_1), .Z(n3508) );
  NAND U5261 ( .A(n3510), .B(n3511), .Z(z2[348]) );
  NANDN U5262 ( .A(xregN_1), .B(zin[347]), .Z(n3511) );
  NAND U5263 ( .A(N352), .B(xregN_1), .Z(n3510) );
  NAND U5264 ( .A(n3512), .B(n3513), .Z(z2[347]) );
  NANDN U5265 ( .A(xregN_1), .B(zin[346]), .Z(n3513) );
  NAND U5266 ( .A(N351), .B(xregN_1), .Z(n3512) );
  NAND U5267 ( .A(n3514), .B(n3515), .Z(z2[346]) );
  NANDN U5268 ( .A(xregN_1), .B(zin[345]), .Z(n3515) );
  NAND U5269 ( .A(N350), .B(xregN_1), .Z(n3514) );
  NAND U5270 ( .A(n3516), .B(n3517), .Z(z2[345]) );
  NANDN U5271 ( .A(xregN_1), .B(zin[344]), .Z(n3517) );
  NAND U5272 ( .A(N349), .B(xregN_1), .Z(n3516) );
  NAND U5273 ( .A(n3518), .B(n3519), .Z(z2[344]) );
  NANDN U5274 ( .A(xregN_1), .B(zin[343]), .Z(n3519) );
  NAND U5275 ( .A(N348), .B(xregN_1), .Z(n3518) );
  NAND U5276 ( .A(n3520), .B(n3521), .Z(z2[343]) );
  NANDN U5277 ( .A(xregN_1), .B(zin[342]), .Z(n3521) );
  NAND U5278 ( .A(N347), .B(xregN_1), .Z(n3520) );
  NAND U5279 ( .A(n3522), .B(n3523), .Z(z2[342]) );
  NANDN U5280 ( .A(xregN_1), .B(zin[341]), .Z(n3523) );
  NAND U5281 ( .A(N346), .B(xregN_1), .Z(n3522) );
  NAND U5282 ( .A(n3524), .B(n3525), .Z(z2[341]) );
  NANDN U5283 ( .A(xregN_1), .B(zin[340]), .Z(n3525) );
  NAND U5284 ( .A(N345), .B(xregN_1), .Z(n3524) );
  NAND U5285 ( .A(n3526), .B(n3527), .Z(z2[340]) );
  NANDN U5286 ( .A(xregN_1), .B(zin[339]), .Z(n3527) );
  NAND U5287 ( .A(N344), .B(xregN_1), .Z(n3526) );
  NAND U5288 ( .A(n3528), .B(n3529), .Z(z2[33]) );
  NANDN U5289 ( .A(xregN_1), .B(zin[32]), .Z(n3529) );
  NAND U5290 ( .A(N37), .B(xregN_1), .Z(n3528) );
  NAND U5291 ( .A(n3530), .B(n3531), .Z(z2[339]) );
  NANDN U5292 ( .A(xregN_1), .B(zin[338]), .Z(n3531) );
  NAND U5293 ( .A(N343), .B(xregN_1), .Z(n3530) );
  NAND U5294 ( .A(n3532), .B(n3533), .Z(z2[338]) );
  NANDN U5295 ( .A(xregN_1), .B(zin[337]), .Z(n3533) );
  NAND U5296 ( .A(N342), .B(xregN_1), .Z(n3532) );
  NAND U5297 ( .A(n3534), .B(n3535), .Z(z2[337]) );
  NANDN U5298 ( .A(xregN_1), .B(zin[336]), .Z(n3535) );
  NAND U5299 ( .A(N341), .B(xregN_1), .Z(n3534) );
  NAND U5300 ( .A(n3536), .B(n3537), .Z(z2[336]) );
  NANDN U5301 ( .A(xregN_1), .B(zin[335]), .Z(n3537) );
  NAND U5302 ( .A(N340), .B(xregN_1), .Z(n3536) );
  NAND U5303 ( .A(n3538), .B(n3539), .Z(z2[335]) );
  NANDN U5304 ( .A(xregN_1), .B(zin[334]), .Z(n3539) );
  NAND U5305 ( .A(N339), .B(xregN_1), .Z(n3538) );
  NAND U5306 ( .A(n3540), .B(n3541), .Z(z2[334]) );
  NANDN U5307 ( .A(xregN_1), .B(zin[333]), .Z(n3541) );
  NAND U5308 ( .A(N338), .B(xregN_1), .Z(n3540) );
  NAND U5309 ( .A(n3542), .B(n3543), .Z(z2[333]) );
  NANDN U5310 ( .A(xregN_1), .B(zin[332]), .Z(n3543) );
  NAND U5311 ( .A(N337), .B(xregN_1), .Z(n3542) );
  NAND U5312 ( .A(n3544), .B(n3545), .Z(z2[332]) );
  NANDN U5313 ( .A(xregN_1), .B(zin[331]), .Z(n3545) );
  NAND U5314 ( .A(N336), .B(xregN_1), .Z(n3544) );
  NAND U5315 ( .A(n3546), .B(n3547), .Z(z2[331]) );
  NANDN U5316 ( .A(xregN_1), .B(zin[330]), .Z(n3547) );
  NAND U5317 ( .A(N335), .B(xregN_1), .Z(n3546) );
  NAND U5318 ( .A(n3548), .B(n3549), .Z(z2[330]) );
  NANDN U5319 ( .A(xregN_1), .B(zin[329]), .Z(n3549) );
  NAND U5320 ( .A(N334), .B(xregN_1), .Z(n3548) );
  NAND U5321 ( .A(n3550), .B(n3551), .Z(z2[32]) );
  NANDN U5322 ( .A(xregN_1), .B(zin[31]), .Z(n3551) );
  NAND U5323 ( .A(N36), .B(xregN_1), .Z(n3550) );
  NAND U5324 ( .A(n3552), .B(n3553), .Z(z2[329]) );
  NANDN U5325 ( .A(xregN_1), .B(zin[328]), .Z(n3553) );
  NAND U5326 ( .A(N333), .B(xregN_1), .Z(n3552) );
  NAND U5327 ( .A(n3554), .B(n3555), .Z(z2[328]) );
  NANDN U5328 ( .A(xregN_1), .B(zin[327]), .Z(n3555) );
  NAND U5329 ( .A(N332), .B(xregN_1), .Z(n3554) );
  NAND U5330 ( .A(n3556), .B(n3557), .Z(z2[327]) );
  NANDN U5331 ( .A(xregN_1), .B(zin[326]), .Z(n3557) );
  NAND U5332 ( .A(N331), .B(xregN_1), .Z(n3556) );
  NAND U5333 ( .A(n3558), .B(n3559), .Z(z2[326]) );
  NANDN U5334 ( .A(xregN_1), .B(zin[325]), .Z(n3559) );
  NAND U5335 ( .A(N330), .B(xregN_1), .Z(n3558) );
  NAND U5336 ( .A(n3560), .B(n3561), .Z(z2[325]) );
  NANDN U5337 ( .A(xregN_1), .B(zin[324]), .Z(n3561) );
  NAND U5338 ( .A(N329), .B(xregN_1), .Z(n3560) );
  NAND U5339 ( .A(n3562), .B(n3563), .Z(z2[324]) );
  NANDN U5340 ( .A(xregN_1), .B(zin[323]), .Z(n3563) );
  NAND U5341 ( .A(N328), .B(xregN_1), .Z(n3562) );
  NAND U5342 ( .A(n3564), .B(n3565), .Z(z2[323]) );
  NANDN U5343 ( .A(xregN_1), .B(zin[322]), .Z(n3565) );
  NAND U5344 ( .A(N327), .B(xregN_1), .Z(n3564) );
  NAND U5345 ( .A(n3566), .B(n3567), .Z(z2[322]) );
  NANDN U5346 ( .A(xregN_1), .B(zin[321]), .Z(n3567) );
  NAND U5347 ( .A(N326), .B(xregN_1), .Z(n3566) );
  NAND U5348 ( .A(n3568), .B(n3569), .Z(z2[321]) );
  NANDN U5349 ( .A(xregN_1), .B(zin[320]), .Z(n3569) );
  NAND U5350 ( .A(N325), .B(xregN_1), .Z(n3568) );
  NAND U5351 ( .A(n3570), .B(n3571), .Z(z2[320]) );
  NANDN U5352 ( .A(xregN_1), .B(zin[319]), .Z(n3571) );
  NAND U5353 ( .A(N324), .B(xregN_1), .Z(n3570) );
  NAND U5354 ( .A(n3572), .B(n3573), .Z(z2[31]) );
  NANDN U5355 ( .A(xregN_1), .B(zin[30]), .Z(n3573) );
  NAND U5356 ( .A(N35), .B(xregN_1), .Z(n3572) );
  NAND U5357 ( .A(n3574), .B(n3575), .Z(z2[319]) );
  NANDN U5358 ( .A(xregN_1), .B(zin[318]), .Z(n3575) );
  NAND U5359 ( .A(N323), .B(xregN_1), .Z(n3574) );
  NAND U5360 ( .A(n3576), .B(n3577), .Z(z2[318]) );
  NANDN U5361 ( .A(xregN_1), .B(zin[317]), .Z(n3577) );
  NAND U5362 ( .A(N322), .B(xregN_1), .Z(n3576) );
  NAND U5363 ( .A(n3578), .B(n3579), .Z(z2[317]) );
  NANDN U5364 ( .A(xregN_1), .B(zin[316]), .Z(n3579) );
  NAND U5365 ( .A(N321), .B(xregN_1), .Z(n3578) );
  NAND U5366 ( .A(n3580), .B(n3581), .Z(z2[316]) );
  NANDN U5367 ( .A(xregN_1), .B(zin[315]), .Z(n3581) );
  NAND U5368 ( .A(N320), .B(xregN_1), .Z(n3580) );
  NAND U5369 ( .A(n3582), .B(n3583), .Z(z2[315]) );
  NANDN U5370 ( .A(xregN_1), .B(zin[314]), .Z(n3583) );
  NAND U5371 ( .A(N319), .B(xregN_1), .Z(n3582) );
  NAND U5372 ( .A(n3584), .B(n3585), .Z(z2[314]) );
  NANDN U5373 ( .A(xregN_1), .B(zin[313]), .Z(n3585) );
  NAND U5374 ( .A(N318), .B(xregN_1), .Z(n3584) );
  NAND U5375 ( .A(n3586), .B(n3587), .Z(z2[313]) );
  NANDN U5376 ( .A(xregN_1), .B(zin[312]), .Z(n3587) );
  NAND U5377 ( .A(N317), .B(xregN_1), .Z(n3586) );
  NAND U5378 ( .A(n3588), .B(n3589), .Z(z2[312]) );
  NANDN U5379 ( .A(xregN_1), .B(zin[311]), .Z(n3589) );
  NAND U5380 ( .A(N316), .B(xregN_1), .Z(n3588) );
  NAND U5381 ( .A(n3590), .B(n3591), .Z(z2[311]) );
  NANDN U5382 ( .A(xregN_1), .B(zin[310]), .Z(n3591) );
  NAND U5383 ( .A(N315), .B(xregN_1), .Z(n3590) );
  NAND U5384 ( .A(n3592), .B(n3593), .Z(z2[310]) );
  NANDN U5385 ( .A(xregN_1), .B(zin[309]), .Z(n3593) );
  NAND U5386 ( .A(N314), .B(xregN_1), .Z(n3592) );
  NAND U5387 ( .A(n3594), .B(n3595), .Z(z2[30]) );
  NANDN U5388 ( .A(xregN_1), .B(zin[29]), .Z(n3595) );
  NAND U5389 ( .A(N34), .B(xregN_1), .Z(n3594) );
  NAND U5390 ( .A(n3596), .B(n3597), .Z(z2[309]) );
  NANDN U5391 ( .A(xregN_1), .B(zin[308]), .Z(n3597) );
  NAND U5392 ( .A(N313), .B(xregN_1), .Z(n3596) );
  NAND U5393 ( .A(n3598), .B(n3599), .Z(z2[308]) );
  NANDN U5394 ( .A(xregN_1), .B(zin[307]), .Z(n3599) );
  NAND U5395 ( .A(N312), .B(xregN_1), .Z(n3598) );
  NAND U5396 ( .A(n3600), .B(n3601), .Z(z2[307]) );
  NANDN U5397 ( .A(xregN_1), .B(zin[306]), .Z(n3601) );
  NAND U5398 ( .A(N311), .B(xregN_1), .Z(n3600) );
  NAND U5399 ( .A(n3602), .B(n3603), .Z(z2[306]) );
  NANDN U5400 ( .A(xregN_1), .B(zin[305]), .Z(n3603) );
  NAND U5401 ( .A(N310), .B(xregN_1), .Z(n3602) );
  NAND U5402 ( .A(n3604), .B(n3605), .Z(z2[305]) );
  NANDN U5403 ( .A(xregN_1), .B(zin[304]), .Z(n3605) );
  NAND U5404 ( .A(N309), .B(xregN_1), .Z(n3604) );
  NAND U5405 ( .A(n3606), .B(n3607), .Z(z2[304]) );
  NANDN U5406 ( .A(xregN_1), .B(zin[303]), .Z(n3607) );
  NAND U5407 ( .A(N308), .B(xregN_1), .Z(n3606) );
  NAND U5408 ( .A(n3608), .B(n3609), .Z(z2[303]) );
  NANDN U5409 ( .A(xregN_1), .B(zin[302]), .Z(n3609) );
  NAND U5410 ( .A(N307), .B(xregN_1), .Z(n3608) );
  NAND U5411 ( .A(n3610), .B(n3611), .Z(z2[302]) );
  NANDN U5412 ( .A(xregN_1), .B(zin[301]), .Z(n3611) );
  NAND U5413 ( .A(N306), .B(xregN_1), .Z(n3610) );
  NAND U5414 ( .A(n3612), .B(n3613), .Z(z2[301]) );
  NANDN U5415 ( .A(xregN_1), .B(zin[300]), .Z(n3613) );
  NAND U5416 ( .A(N305), .B(xregN_1), .Z(n3612) );
  NAND U5417 ( .A(n3614), .B(n3615), .Z(z2[300]) );
  NANDN U5418 ( .A(xregN_1), .B(zin[299]), .Z(n3615) );
  NAND U5419 ( .A(N304), .B(xregN_1), .Z(n3614) );
  NAND U5420 ( .A(n3616), .B(n3617), .Z(z2[2]) );
  NANDN U5421 ( .A(xregN_1), .B(zin[1]), .Z(n3617) );
  NAND U5422 ( .A(N6), .B(xregN_1), .Z(n3616) );
  NAND U5423 ( .A(n3618), .B(n3619), .Z(z2[29]) );
  NANDN U5424 ( .A(xregN_1), .B(zin[28]), .Z(n3619) );
  NAND U5425 ( .A(N33), .B(xregN_1), .Z(n3618) );
  NAND U5426 ( .A(n3620), .B(n3621), .Z(z2[299]) );
  NANDN U5427 ( .A(xregN_1), .B(zin[298]), .Z(n3621) );
  NAND U5428 ( .A(N303), .B(xregN_1), .Z(n3620) );
  NAND U5429 ( .A(n3622), .B(n3623), .Z(z2[298]) );
  NANDN U5430 ( .A(xregN_1), .B(zin[297]), .Z(n3623) );
  NAND U5431 ( .A(N302), .B(xregN_1), .Z(n3622) );
  NAND U5432 ( .A(n3624), .B(n3625), .Z(z2[297]) );
  NANDN U5433 ( .A(xregN_1), .B(zin[296]), .Z(n3625) );
  NAND U5434 ( .A(N301), .B(xregN_1), .Z(n3624) );
  NAND U5435 ( .A(n3626), .B(n3627), .Z(z2[296]) );
  NANDN U5436 ( .A(xregN_1), .B(zin[295]), .Z(n3627) );
  NAND U5437 ( .A(N300), .B(xregN_1), .Z(n3626) );
  NAND U5438 ( .A(n3628), .B(n3629), .Z(z2[295]) );
  NANDN U5439 ( .A(xregN_1), .B(zin[294]), .Z(n3629) );
  NAND U5440 ( .A(N299), .B(xregN_1), .Z(n3628) );
  NAND U5441 ( .A(n3630), .B(n3631), .Z(z2[294]) );
  NANDN U5442 ( .A(xregN_1), .B(zin[293]), .Z(n3631) );
  NAND U5443 ( .A(N298), .B(xregN_1), .Z(n3630) );
  NAND U5444 ( .A(n3632), .B(n3633), .Z(z2[293]) );
  NANDN U5445 ( .A(xregN_1), .B(zin[292]), .Z(n3633) );
  NAND U5446 ( .A(N297), .B(xregN_1), .Z(n3632) );
  NAND U5447 ( .A(n3634), .B(n3635), .Z(z2[292]) );
  NANDN U5448 ( .A(xregN_1), .B(zin[291]), .Z(n3635) );
  NAND U5449 ( .A(N296), .B(xregN_1), .Z(n3634) );
  NAND U5450 ( .A(n3636), .B(n3637), .Z(z2[291]) );
  NANDN U5451 ( .A(xregN_1), .B(zin[290]), .Z(n3637) );
  NAND U5452 ( .A(N295), .B(xregN_1), .Z(n3636) );
  NAND U5453 ( .A(n3638), .B(n3639), .Z(z2[290]) );
  NANDN U5454 ( .A(xregN_1), .B(zin[289]), .Z(n3639) );
  NAND U5455 ( .A(N294), .B(xregN_1), .Z(n3638) );
  NAND U5456 ( .A(n3640), .B(n3641), .Z(z2[28]) );
  NANDN U5457 ( .A(xregN_1), .B(zin[27]), .Z(n3641) );
  NAND U5458 ( .A(N32), .B(xregN_1), .Z(n3640) );
  NAND U5459 ( .A(n3642), .B(n3643), .Z(z2[289]) );
  NANDN U5460 ( .A(xregN_1), .B(zin[288]), .Z(n3643) );
  NAND U5461 ( .A(N293), .B(xregN_1), .Z(n3642) );
  NAND U5462 ( .A(n3644), .B(n3645), .Z(z2[288]) );
  NANDN U5463 ( .A(xregN_1), .B(zin[287]), .Z(n3645) );
  NAND U5464 ( .A(N292), .B(xregN_1), .Z(n3644) );
  NAND U5465 ( .A(n3646), .B(n3647), .Z(z2[287]) );
  NANDN U5466 ( .A(xregN_1), .B(zin[286]), .Z(n3647) );
  NAND U5467 ( .A(N291), .B(xregN_1), .Z(n3646) );
  NAND U5468 ( .A(n3648), .B(n3649), .Z(z2[286]) );
  NANDN U5469 ( .A(xregN_1), .B(zin[285]), .Z(n3649) );
  NAND U5470 ( .A(N290), .B(xregN_1), .Z(n3648) );
  NAND U5471 ( .A(n3650), .B(n3651), .Z(z2[285]) );
  NANDN U5472 ( .A(xregN_1), .B(zin[284]), .Z(n3651) );
  NAND U5473 ( .A(N289), .B(xregN_1), .Z(n3650) );
  NAND U5474 ( .A(n3652), .B(n3653), .Z(z2[284]) );
  NANDN U5475 ( .A(xregN_1), .B(zin[283]), .Z(n3653) );
  NAND U5476 ( .A(N288), .B(xregN_1), .Z(n3652) );
  NAND U5477 ( .A(n3654), .B(n3655), .Z(z2[283]) );
  NANDN U5478 ( .A(xregN_1), .B(zin[282]), .Z(n3655) );
  NAND U5479 ( .A(N287), .B(xregN_1), .Z(n3654) );
  NAND U5480 ( .A(n3656), .B(n3657), .Z(z2[282]) );
  NANDN U5481 ( .A(xregN_1), .B(zin[281]), .Z(n3657) );
  NAND U5482 ( .A(N286), .B(xregN_1), .Z(n3656) );
  NAND U5483 ( .A(n3658), .B(n3659), .Z(z2[281]) );
  NANDN U5484 ( .A(xregN_1), .B(zin[280]), .Z(n3659) );
  NAND U5485 ( .A(N285), .B(xregN_1), .Z(n3658) );
  NAND U5486 ( .A(n3660), .B(n3661), .Z(z2[280]) );
  NANDN U5487 ( .A(xregN_1), .B(zin[279]), .Z(n3661) );
  NAND U5488 ( .A(N284), .B(xregN_1), .Z(n3660) );
  NAND U5489 ( .A(n3662), .B(n3663), .Z(z2[27]) );
  NANDN U5490 ( .A(xregN_1), .B(zin[26]), .Z(n3663) );
  NAND U5491 ( .A(N31), .B(xregN_1), .Z(n3662) );
  NAND U5492 ( .A(n3664), .B(n3665), .Z(z2[279]) );
  NANDN U5493 ( .A(xregN_1), .B(zin[278]), .Z(n3665) );
  NAND U5494 ( .A(N283), .B(xregN_1), .Z(n3664) );
  NAND U5495 ( .A(n3666), .B(n3667), .Z(z2[278]) );
  NANDN U5496 ( .A(xregN_1), .B(zin[277]), .Z(n3667) );
  NAND U5497 ( .A(N282), .B(xregN_1), .Z(n3666) );
  NAND U5498 ( .A(n3668), .B(n3669), .Z(z2[277]) );
  NANDN U5499 ( .A(xregN_1), .B(zin[276]), .Z(n3669) );
  NAND U5500 ( .A(N281), .B(xregN_1), .Z(n3668) );
  NAND U5501 ( .A(n3670), .B(n3671), .Z(z2[276]) );
  NANDN U5502 ( .A(xregN_1), .B(zin[275]), .Z(n3671) );
  NAND U5503 ( .A(N280), .B(xregN_1), .Z(n3670) );
  NAND U5504 ( .A(n3672), .B(n3673), .Z(z2[275]) );
  NANDN U5505 ( .A(xregN_1), .B(zin[274]), .Z(n3673) );
  NAND U5506 ( .A(N279), .B(xregN_1), .Z(n3672) );
  NAND U5507 ( .A(n3674), .B(n3675), .Z(z2[274]) );
  NANDN U5508 ( .A(xregN_1), .B(zin[273]), .Z(n3675) );
  NAND U5509 ( .A(N278), .B(xregN_1), .Z(n3674) );
  NAND U5510 ( .A(n3676), .B(n3677), .Z(z2[273]) );
  NANDN U5511 ( .A(xregN_1), .B(zin[272]), .Z(n3677) );
  NAND U5512 ( .A(N277), .B(xregN_1), .Z(n3676) );
  NAND U5513 ( .A(n3678), .B(n3679), .Z(z2[272]) );
  NANDN U5514 ( .A(xregN_1), .B(zin[271]), .Z(n3679) );
  NAND U5515 ( .A(N276), .B(xregN_1), .Z(n3678) );
  NAND U5516 ( .A(n3680), .B(n3681), .Z(z2[271]) );
  NANDN U5517 ( .A(xregN_1), .B(zin[270]), .Z(n3681) );
  NAND U5518 ( .A(N275), .B(xregN_1), .Z(n3680) );
  NAND U5519 ( .A(n3682), .B(n3683), .Z(z2[270]) );
  NANDN U5520 ( .A(xregN_1), .B(zin[269]), .Z(n3683) );
  NAND U5521 ( .A(N274), .B(xregN_1), .Z(n3682) );
  NAND U5522 ( .A(n3684), .B(n3685), .Z(z2[26]) );
  NANDN U5523 ( .A(xregN_1), .B(zin[25]), .Z(n3685) );
  NAND U5524 ( .A(N30), .B(xregN_1), .Z(n3684) );
  NAND U5525 ( .A(n3686), .B(n3687), .Z(z2[269]) );
  NANDN U5526 ( .A(xregN_1), .B(zin[268]), .Z(n3687) );
  NAND U5527 ( .A(N273), .B(xregN_1), .Z(n3686) );
  NAND U5528 ( .A(n3688), .B(n3689), .Z(z2[268]) );
  NANDN U5529 ( .A(xregN_1), .B(zin[267]), .Z(n3689) );
  NAND U5530 ( .A(N272), .B(xregN_1), .Z(n3688) );
  NAND U5531 ( .A(n3690), .B(n3691), .Z(z2[267]) );
  NANDN U5532 ( .A(xregN_1), .B(zin[266]), .Z(n3691) );
  NAND U5533 ( .A(N271), .B(xregN_1), .Z(n3690) );
  NAND U5534 ( .A(n3692), .B(n3693), .Z(z2[266]) );
  NANDN U5535 ( .A(xregN_1), .B(zin[265]), .Z(n3693) );
  NAND U5536 ( .A(N270), .B(xregN_1), .Z(n3692) );
  NAND U5537 ( .A(n3694), .B(n3695), .Z(z2[265]) );
  NANDN U5538 ( .A(xregN_1), .B(zin[264]), .Z(n3695) );
  NAND U5539 ( .A(N269), .B(xregN_1), .Z(n3694) );
  NAND U5540 ( .A(n3696), .B(n3697), .Z(z2[264]) );
  NANDN U5541 ( .A(xregN_1), .B(zin[263]), .Z(n3697) );
  NAND U5542 ( .A(N268), .B(xregN_1), .Z(n3696) );
  NAND U5543 ( .A(n3698), .B(n3699), .Z(z2[263]) );
  NANDN U5544 ( .A(xregN_1), .B(zin[262]), .Z(n3699) );
  NAND U5545 ( .A(N267), .B(xregN_1), .Z(n3698) );
  NAND U5546 ( .A(n3700), .B(n3701), .Z(z2[262]) );
  NANDN U5547 ( .A(xregN_1), .B(zin[261]), .Z(n3701) );
  NAND U5548 ( .A(N266), .B(xregN_1), .Z(n3700) );
  NAND U5549 ( .A(n3702), .B(n3703), .Z(z2[261]) );
  NANDN U5550 ( .A(xregN_1), .B(zin[260]), .Z(n3703) );
  NAND U5551 ( .A(N265), .B(xregN_1), .Z(n3702) );
  NAND U5552 ( .A(n3704), .B(n3705), .Z(z2[260]) );
  NANDN U5553 ( .A(xregN_1), .B(zin[259]), .Z(n3705) );
  NAND U5554 ( .A(N264), .B(xregN_1), .Z(n3704) );
  NAND U5555 ( .A(n3706), .B(n3707), .Z(z2[25]) );
  NANDN U5556 ( .A(xregN_1), .B(zin[24]), .Z(n3707) );
  NAND U5557 ( .A(N29), .B(xregN_1), .Z(n3706) );
  NAND U5558 ( .A(n3708), .B(n3709), .Z(z2[259]) );
  NANDN U5559 ( .A(xregN_1), .B(zin[258]), .Z(n3709) );
  NAND U5560 ( .A(N263), .B(xregN_1), .Z(n3708) );
  NAND U5561 ( .A(n3710), .B(n3711), .Z(z2[258]) );
  NANDN U5562 ( .A(xregN_1), .B(zin[257]), .Z(n3711) );
  NAND U5563 ( .A(N262), .B(xregN_1), .Z(n3710) );
  NAND U5564 ( .A(n3712), .B(n3713), .Z(z2[257]) );
  NANDN U5565 ( .A(xregN_1), .B(zin[256]), .Z(n3713) );
  NAND U5566 ( .A(N261), .B(xregN_1), .Z(n3712) );
  NAND U5567 ( .A(n3714), .B(n3715), .Z(z2[256]) );
  NANDN U5568 ( .A(xregN_1), .B(zin[255]), .Z(n3715) );
  NAND U5569 ( .A(N260), .B(xregN_1), .Z(n3714) );
  NAND U5570 ( .A(n3716), .B(n3717), .Z(z2[255]) );
  NANDN U5571 ( .A(xregN_1), .B(zin[254]), .Z(n3717) );
  NAND U5572 ( .A(N259), .B(xregN_1), .Z(n3716) );
  NAND U5573 ( .A(n3718), .B(n3719), .Z(z2[254]) );
  NANDN U5574 ( .A(xregN_1), .B(zin[253]), .Z(n3719) );
  NAND U5575 ( .A(N258), .B(xregN_1), .Z(n3718) );
  NAND U5576 ( .A(n3720), .B(n3721), .Z(z2[253]) );
  NANDN U5577 ( .A(xregN_1), .B(zin[252]), .Z(n3721) );
  NAND U5578 ( .A(N257), .B(xregN_1), .Z(n3720) );
  NAND U5579 ( .A(n3722), .B(n3723), .Z(z2[252]) );
  NANDN U5580 ( .A(xregN_1), .B(zin[251]), .Z(n3723) );
  NAND U5581 ( .A(N256), .B(xregN_1), .Z(n3722) );
  NAND U5582 ( .A(n3724), .B(n3725), .Z(z2[251]) );
  NANDN U5583 ( .A(xregN_1), .B(zin[250]), .Z(n3725) );
  NAND U5584 ( .A(N255), .B(xregN_1), .Z(n3724) );
  NAND U5585 ( .A(n3726), .B(n3727), .Z(z2[250]) );
  NANDN U5586 ( .A(xregN_1), .B(zin[249]), .Z(n3727) );
  NAND U5587 ( .A(N254), .B(xregN_1), .Z(n3726) );
  NAND U5588 ( .A(n3728), .B(n3729), .Z(z2[24]) );
  NANDN U5589 ( .A(xregN_1), .B(zin[23]), .Z(n3729) );
  NAND U5590 ( .A(N28), .B(xregN_1), .Z(n3728) );
  NAND U5591 ( .A(n3730), .B(n3731), .Z(z2[249]) );
  NANDN U5592 ( .A(xregN_1), .B(zin[248]), .Z(n3731) );
  NAND U5593 ( .A(N253), .B(xregN_1), .Z(n3730) );
  NAND U5594 ( .A(n3732), .B(n3733), .Z(z2[248]) );
  NANDN U5595 ( .A(xregN_1), .B(zin[247]), .Z(n3733) );
  NAND U5596 ( .A(N252), .B(xregN_1), .Z(n3732) );
  NAND U5597 ( .A(n3734), .B(n3735), .Z(z2[247]) );
  NANDN U5598 ( .A(xregN_1), .B(zin[246]), .Z(n3735) );
  NAND U5599 ( .A(N251), .B(xregN_1), .Z(n3734) );
  NAND U5600 ( .A(n3736), .B(n3737), .Z(z2[246]) );
  NANDN U5601 ( .A(xregN_1), .B(zin[245]), .Z(n3737) );
  NAND U5602 ( .A(N250), .B(xregN_1), .Z(n3736) );
  NAND U5603 ( .A(n3738), .B(n3739), .Z(z2[245]) );
  NANDN U5604 ( .A(xregN_1), .B(zin[244]), .Z(n3739) );
  NAND U5605 ( .A(N249), .B(xregN_1), .Z(n3738) );
  NAND U5606 ( .A(n3740), .B(n3741), .Z(z2[244]) );
  NANDN U5607 ( .A(xregN_1), .B(zin[243]), .Z(n3741) );
  NAND U5608 ( .A(N248), .B(xregN_1), .Z(n3740) );
  NAND U5609 ( .A(n3742), .B(n3743), .Z(z2[243]) );
  NANDN U5610 ( .A(xregN_1), .B(zin[242]), .Z(n3743) );
  NAND U5611 ( .A(N247), .B(xregN_1), .Z(n3742) );
  NAND U5612 ( .A(n3744), .B(n3745), .Z(z2[242]) );
  NANDN U5613 ( .A(xregN_1), .B(zin[241]), .Z(n3745) );
  NAND U5614 ( .A(N246), .B(xregN_1), .Z(n3744) );
  NAND U5615 ( .A(n3746), .B(n3747), .Z(z2[241]) );
  NANDN U5616 ( .A(xregN_1), .B(zin[240]), .Z(n3747) );
  NAND U5617 ( .A(N245), .B(xregN_1), .Z(n3746) );
  NAND U5618 ( .A(n3748), .B(n3749), .Z(z2[240]) );
  NANDN U5619 ( .A(xregN_1), .B(zin[239]), .Z(n3749) );
  NAND U5620 ( .A(N244), .B(xregN_1), .Z(n3748) );
  NAND U5621 ( .A(n3750), .B(n3751), .Z(z2[23]) );
  NANDN U5622 ( .A(xregN_1), .B(zin[22]), .Z(n3751) );
  NAND U5623 ( .A(N27), .B(xregN_1), .Z(n3750) );
  NAND U5624 ( .A(n3752), .B(n3753), .Z(z2[239]) );
  NANDN U5625 ( .A(xregN_1), .B(zin[238]), .Z(n3753) );
  NAND U5626 ( .A(N243), .B(xregN_1), .Z(n3752) );
  NAND U5627 ( .A(n3754), .B(n3755), .Z(z2[238]) );
  NANDN U5628 ( .A(xregN_1), .B(zin[237]), .Z(n3755) );
  NAND U5629 ( .A(N242), .B(xregN_1), .Z(n3754) );
  NAND U5630 ( .A(n3756), .B(n3757), .Z(z2[237]) );
  NANDN U5631 ( .A(xregN_1), .B(zin[236]), .Z(n3757) );
  NAND U5632 ( .A(N241), .B(xregN_1), .Z(n3756) );
  NAND U5633 ( .A(n3758), .B(n3759), .Z(z2[236]) );
  NANDN U5634 ( .A(xregN_1), .B(zin[235]), .Z(n3759) );
  NAND U5635 ( .A(N240), .B(xregN_1), .Z(n3758) );
  NAND U5636 ( .A(n3760), .B(n3761), .Z(z2[235]) );
  NANDN U5637 ( .A(xregN_1), .B(zin[234]), .Z(n3761) );
  NAND U5638 ( .A(N239), .B(xregN_1), .Z(n3760) );
  NAND U5639 ( .A(n3762), .B(n3763), .Z(z2[234]) );
  NANDN U5640 ( .A(xregN_1), .B(zin[233]), .Z(n3763) );
  NAND U5641 ( .A(N238), .B(xregN_1), .Z(n3762) );
  NAND U5642 ( .A(n3764), .B(n3765), .Z(z2[233]) );
  NANDN U5643 ( .A(xregN_1), .B(zin[232]), .Z(n3765) );
  NAND U5644 ( .A(N237), .B(xregN_1), .Z(n3764) );
  NAND U5645 ( .A(n3766), .B(n3767), .Z(z2[232]) );
  NANDN U5646 ( .A(xregN_1), .B(zin[231]), .Z(n3767) );
  NAND U5647 ( .A(N236), .B(xregN_1), .Z(n3766) );
  NAND U5648 ( .A(n3768), .B(n3769), .Z(z2[231]) );
  NANDN U5649 ( .A(xregN_1), .B(zin[230]), .Z(n3769) );
  NAND U5650 ( .A(N235), .B(xregN_1), .Z(n3768) );
  NAND U5651 ( .A(n3770), .B(n3771), .Z(z2[230]) );
  NANDN U5652 ( .A(xregN_1), .B(zin[229]), .Z(n3771) );
  NAND U5653 ( .A(N234), .B(xregN_1), .Z(n3770) );
  NAND U5654 ( .A(n3772), .B(n3773), .Z(z2[22]) );
  NANDN U5655 ( .A(xregN_1), .B(zin[21]), .Z(n3773) );
  NAND U5656 ( .A(N26), .B(xregN_1), .Z(n3772) );
  NAND U5657 ( .A(n3774), .B(n3775), .Z(z2[229]) );
  NANDN U5658 ( .A(xregN_1), .B(zin[228]), .Z(n3775) );
  NAND U5659 ( .A(N233), .B(xregN_1), .Z(n3774) );
  NAND U5660 ( .A(n3776), .B(n3777), .Z(z2[228]) );
  NANDN U5661 ( .A(xregN_1), .B(zin[227]), .Z(n3777) );
  NAND U5662 ( .A(N232), .B(xregN_1), .Z(n3776) );
  NAND U5663 ( .A(n3778), .B(n3779), .Z(z2[227]) );
  NANDN U5664 ( .A(xregN_1), .B(zin[226]), .Z(n3779) );
  NAND U5665 ( .A(N231), .B(xregN_1), .Z(n3778) );
  NAND U5666 ( .A(n3780), .B(n3781), .Z(z2[226]) );
  NANDN U5667 ( .A(xregN_1), .B(zin[225]), .Z(n3781) );
  NAND U5668 ( .A(N230), .B(xregN_1), .Z(n3780) );
  NAND U5669 ( .A(n3782), .B(n3783), .Z(z2[225]) );
  NANDN U5670 ( .A(xregN_1), .B(zin[224]), .Z(n3783) );
  NAND U5671 ( .A(N229), .B(xregN_1), .Z(n3782) );
  NAND U5672 ( .A(n3784), .B(n3785), .Z(z2[224]) );
  NANDN U5673 ( .A(xregN_1), .B(zin[223]), .Z(n3785) );
  NAND U5674 ( .A(N228), .B(xregN_1), .Z(n3784) );
  NAND U5675 ( .A(n3786), .B(n3787), .Z(z2[223]) );
  NANDN U5676 ( .A(xregN_1), .B(zin[222]), .Z(n3787) );
  NAND U5677 ( .A(N227), .B(xregN_1), .Z(n3786) );
  NAND U5678 ( .A(n3788), .B(n3789), .Z(z2[222]) );
  NANDN U5679 ( .A(xregN_1), .B(zin[221]), .Z(n3789) );
  NAND U5680 ( .A(N226), .B(xregN_1), .Z(n3788) );
  NAND U5681 ( .A(n3790), .B(n3791), .Z(z2[221]) );
  NANDN U5682 ( .A(xregN_1), .B(zin[220]), .Z(n3791) );
  NAND U5683 ( .A(N225), .B(xregN_1), .Z(n3790) );
  NAND U5684 ( .A(n3792), .B(n3793), .Z(z2[220]) );
  NANDN U5685 ( .A(xregN_1), .B(zin[219]), .Z(n3793) );
  NAND U5686 ( .A(N224), .B(xregN_1), .Z(n3792) );
  NAND U5687 ( .A(n3794), .B(n3795), .Z(z2[21]) );
  NANDN U5688 ( .A(xregN_1), .B(zin[20]), .Z(n3795) );
  NAND U5689 ( .A(N25), .B(xregN_1), .Z(n3794) );
  NAND U5690 ( .A(n3796), .B(n3797), .Z(z2[219]) );
  NANDN U5691 ( .A(xregN_1), .B(zin[218]), .Z(n3797) );
  NAND U5692 ( .A(N223), .B(xregN_1), .Z(n3796) );
  NAND U5693 ( .A(n3798), .B(n3799), .Z(z2[218]) );
  NANDN U5694 ( .A(xregN_1), .B(zin[217]), .Z(n3799) );
  NAND U5695 ( .A(N222), .B(xregN_1), .Z(n3798) );
  NAND U5696 ( .A(n3800), .B(n3801), .Z(z2[217]) );
  NANDN U5697 ( .A(xregN_1), .B(zin[216]), .Z(n3801) );
  NAND U5698 ( .A(N221), .B(xregN_1), .Z(n3800) );
  NAND U5699 ( .A(n3802), .B(n3803), .Z(z2[216]) );
  NANDN U5700 ( .A(xregN_1), .B(zin[215]), .Z(n3803) );
  NAND U5701 ( .A(N220), .B(xregN_1), .Z(n3802) );
  NAND U5702 ( .A(n3804), .B(n3805), .Z(z2[215]) );
  NANDN U5703 ( .A(xregN_1), .B(zin[214]), .Z(n3805) );
  NAND U5704 ( .A(N219), .B(xregN_1), .Z(n3804) );
  NAND U5705 ( .A(n3806), .B(n3807), .Z(z2[214]) );
  NANDN U5706 ( .A(xregN_1), .B(zin[213]), .Z(n3807) );
  NAND U5707 ( .A(N218), .B(xregN_1), .Z(n3806) );
  NAND U5708 ( .A(n3808), .B(n3809), .Z(z2[213]) );
  NANDN U5709 ( .A(xregN_1), .B(zin[212]), .Z(n3809) );
  NAND U5710 ( .A(N217), .B(xregN_1), .Z(n3808) );
  NAND U5711 ( .A(n3810), .B(n3811), .Z(z2[212]) );
  NANDN U5712 ( .A(xregN_1), .B(zin[211]), .Z(n3811) );
  NAND U5713 ( .A(N216), .B(xregN_1), .Z(n3810) );
  NAND U5714 ( .A(n3812), .B(n3813), .Z(z2[211]) );
  NANDN U5715 ( .A(xregN_1), .B(zin[210]), .Z(n3813) );
  NAND U5716 ( .A(N215), .B(xregN_1), .Z(n3812) );
  NAND U5717 ( .A(n3814), .B(n3815), .Z(z2[210]) );
  NANDN U5718 ( .A(xregN_1), .B(zin[209]), .Z(n3815) );
  NAND U5719 ( .A(N214), .B(xregN_1), .Z(n3814) );
  NAND U5720 ( .A(n3816), .B(n3817), .Z(z2[20]) );
  NANDN U5721 ( .A(xregN_1), .B(zin[19]), .Z(n3817) );
  NAND U5722 ( .A(N24), .B(xregN_1), .Z(n3816) );
  NAND U5723 ( .A(n3818), .B(n3819), .Z(z2[209]) );
  NANDN U5724 ( .A(xregN_1), .B(zin[208]), .Z(n3819) );
  NAND U5725 ( .A(N213), .B(xregN_1), .Z(n3818) );
  NAND U5726 ( .A(n3820), .B(n3821), .Z(z2[208]) );
  NANDN U5727 ( .A(xregN_1), .B(zin[207]), .Z(n3821) );
  NAND U5728 ( .A(N212), .B(xregN_1), .Z(n3820) );
  NAND U5729 ( .A(n3822), .B(n3823), .Z(z2[207]) );
  NANDN U5730 ( .A(xregN_1), .B(zin[206]), .Z(n3823) );
  NAND U5731 ( .A(N211), .B(xregN_1), .Z(n3822) );
  NAND U5732 ( .A(n3824), .B(n3825), .Z(z2[206]) );
  NANDN U5733 ( .A(xregN_1), .B(zin[205]), .Z(n3825) );
  NAND U5734 ( .A(N210), .B(xregN_1), .Z(n3824) );
  NAND U5735 ( .A(n3826), .B(n3827), .Z(z2[205]) );
  NANDN U5736 ( .A(xregN_1), .B(zin[204]), .Z(n3827) );
  NAND U5737 ( .A(N209), .B(xregN_1), .Z(n3826) );
  NAND U5738 ( .A(n3828), .B(n3829), .Z(z2[204]) );
  NANDN U5739 ( .A(xregN_1), .B(zin[203]), .Z(n3829) );
  NAND U5740 ( .A(N208), .B(xregN_1), .Z(n3828) );
  NAND U5741 ( .A(n3830), .B(n3831), .Z(z2[203]) );
  NANDN U5742 ( .A(xregN_1), .B(zin[202]), .Z(n3831) );
  NAND U5743 ( .A(N207), .B(xregN_1), .Z(n3830) );
  NAND U5744 ( .A(n3832), .B(n3833), .Z(z2[202]) );
  NANDN U5745 ( .A(xregN_1), .B(zin[201]), .Z(n3833) );
  NAND U5746 ( .A(N206), .B(xregN_1), .Z(n3832) );
  NAND U5747 ( .A(n3834), .B(n3835), .Z(z2[201]) );
  NANDN U5748 ( .A(xregN_1), .B(zin[200]), .Z(n3835) );
  NAND U5749 ( .A(N205), .B(xregN_1), .Z(n3834) );
  NAND U5750 ( .A(n3836), .B(n3837), .Z(z2[200]) );
  NANDN U5751 ( .A(xregN_1), .B(zin[199]), .Z(n3837) );
  NAND U5752 ( .A(N204), .B(xregN_1), .Z(n3836) );
  NAND U5753 ( .A(n3838), .B(n3839), .Z(z2[1]) );
  NANDN U5754 ( .A(xregN_1), .B(zin[0]), .Z(n3839) );
  NAND U5755 ( .A(N5), .B(xregN_1), .Z(n3838) );
  NAND U5756 ( .A(n3840), .B(n3841), .Z(z2[19]) );
  NANDN U5757 ( .A(xregN_1), .B(zin[18]), .Z(n3841) );
  NAND U5758 ( .A(N23), .B(xregN_1), .Z(n3840) );
  NAND U5759 ( .A(n3842), .B(n3843), .Z(z2[199]) );
  NANDN U5760 ( .A(xregN_1), .B(zin[198]), .Z(n3843) );
  NAND U5761 ( .A(N203), .B(xregN_1), .Z(n3842) );
  NAND U5762 ( .A(n3844), .B(n3845), .Z(z2[198]) );
  NANDN U5763 ( .A(xregN_1), .B(zin[197]), .Z(n3845) );
  NAND U5764 ( .A(N202), .B(xregN_1), .Z(n3844) );
  NAND U5765 ( .A(n3846), .B(n3847), .Z(z2[197]) );
  NANDN U5766 ( .A(xregN_1), .B(zin[196]), .Z(n3847) );
  NAND U5767 ( .A(N201), .B(xregN_1), .Z(n3846) );
  NAND U5768 ( .A(n3848), .B(n3849), .Z(z2[196]) );
  NANDN U5769 ( .A(xregN_1), .B(zin[195]), .Z(n3849) );
  NAND U5770 ( .A(N200), .B(xregN_1), .Z(n3848) );
  NAND U5771 ( .A(n3850), .B(n3851), .Z(z2[195]) );
  NANDN U5772 ( .A(xregN_1), .B(zin[194]), .Z(n3851) );
  NAND U5773 ( .A(N199), .B(xregN_1), .Z(n3850) );
  NAND U5774 ( .A(n3852), .B(n3853), .Z(z2[194]) );
  NANDN U5775 ( .A(xregN_1), .B(zin[193]), .Z(n3853) );
  NAND U5776 ( .A(N198), .B(xregN_1), .Z(n3852) );
  NAND U5777 ( .A(n3854), .B(n3855), .Z(z2[193]) );
  NANDN U5778 ( .A(xregN_1), .B(zin[192]), .Z(n3855) );
  NAND U5779 ( .A(N197), .B(xregN_1), .Z(n3854) );
  NAND U5780 ( .A(n3856), .B(n3857), .Z(z2[192]) );
  NANDN U5781 ( .A(xregN_1), .B(zin[191]), .Z(n3857) );
  NAND U5782 ( .A(N196), .B(xregN_1), .Z(n3856) );
  NAND U5783 ( .A(n3858), .B(n3859), .Z(z2[191]) );
  NANDN U5784 ( .A(xregN_1), .B(zin[190]), .Z(n3859) );
  NAND U5785 ( .A(N195), .B(xregN_1), .Z(n3858) );
  NAND U5786 ( .A(n3860), .B(n3861), .Z(z2[190]) );
  NANDN U5787 ( .A(xregN_1), .B(zin[189]), .Z(n3861) );
  NAND U5788 ( .A(N194), .B(xregN_1), .Z(n3860) );
  NAND U5789 ( .A(n3862), .B(n3863), .Z(z2[18]) );
  NANDN U5790 ( .A(xregN_1), .B(zin[17]), .Z(n3863) );
  NAND U5791 ( .A(N22), .B(xregN_1), .Z(n3862) );
  NAND U5792 ( .A(n3864), .B(n3865), .Z(z2[189]) );
  NANDN U5793 ( .A(xregN_1), .B(zin[188]), .Z(n3865) );
  NAND U5794 ( .A(N193), .B(xregN_1), .Z(n3864) );
  NAND U5795 ( .A(n3866), .B(n3867), .Z(z2[188]) );
  NANDN U5796 ( .A(xregN_1), .B(zin[187]), .Z(n3867) );
  NAND U5797 ( .A(N192), .B(xregN_1), .Z(n3866) );
  NAND U5798 ( .A(n3868), .B(n3869), .Z(z2[187]) );
  NANDN U5799 ( .A(xregN_1), .B(zin[186]), .Z(n3869) );
  NAND U5800 ( .A(N191), .B(xregN_1), .Z(n3868) );
  NAND U5801 ( .A(n3870), .B(n3871), .Z(z2[186]) );
  NANDN U5802 ( .A(xregN_1), .B(zin[185]), .Z(n3871) );
  NAND U5803 ( .A(N190), .B(xregN_1), .Z(n3870) );
  NAND U5804 ( .A(n3872), .B(n3873), .Z(z2[185]) );
  NANDN U5805 ( .A(xregN_1), .B(zin[184]), .Z(n3873) );
  NAND U5806 ( .A(N189), .B(xregN_1), .Z(n3872) );
  NAND U5807 ( .A(n3874), .B(n3875), .Z(z2[184]) );
  NANDN U5808 ( .A(xregN_1), .B(zin[183]), .Z(n3875) );
  NAND U5809 ( .A(N188), .B(xregN_1), .Z(n3874) );
  NAND U5810 ( .A(n3876), .B(n3877), .Z(z2[183]) );
  NANDN U5811 ( .A(xregN_1), .B(zin[182]), .Z(n3877) );
  NAND U5812 ( .A(N187), .B(xregN_1), .Z(n3876) );
  NAND U5813 ( .A(n3878), .B(n3879), .Z(z2[182]) );
  NANDN U5814 ( .A(xregN_1), .B(zin[181]), .Z(n3879) );
  NAND U5815 ( .A(N186), .B(xregN_1), .Z(n3878) );
  NAND U5816 ( .A(n3880), .B(n3881), .Z(z2[181]) );
  NANDN U5817 ( .A(xregN_1), .B(zin[180]), .Z(n3881) );
  NAND U5818 ( .A(N185), .B(xregN_1), .Z(n3880) );
  NAND U5819 ( .A(n3882), .B(n3883), .Z(z2[180]) );
  NANDN U5820 ( .A(xregN_1), .B(zin[179]), .Z(n3883) );
  NAND U5821 ( .A(N184), .B(xregN_1), .Z(n3882) );
  NAND U5822 ( .A(n3884), .B(n3885), .Z(z2[17]) );
  NANDN U5823 ( .A(xregN_1), .B(zin[16]), .Z(n3885) );
  NAND U5824 ( .A(N21), .B(xregN_1), .Z(n3884) );
  NAND U5825 ( .A(n3886), .B(n3887), .Z(z2[179]) );
  NANDN U5826 ( .A(xregN_1), .B(zin[178]), .Z(n3887) );
  NAND U5827 ( .A(N183), .B(xregN_1), .Z(n3886) );
  NAND U5828 ( .A(n3888), .B(n3889), .Z(z2[178]) );
  NANDN U5829 ( .A(xregN_1), .B(zin[177]), .Z(n3889) );
  NAND U5830 ( .A(N182), .B(xregN_1), .Z(n3888) );
  NAND U5831 ( .A(n3890), .B(n3891), .Z(z2[177]) );
  NANDN U5832 ( .A(xregN_1), .B(zin[176]), .Z(n3891) );
  NAND U5833 ( .A(N181), .B(xregN_1), .Z(n3890) );
  NAND U5834 ( .A(n3892), .B(n3893), .Z(z2[176]) );
  NANDN U5835 ( .A(xregN_1), .B(zin[175]), .Z(n3893) );
  NAND U5836 ( .A(N180), .B(xregN_1), .Z(n3892) );
  NAND U5837 ( .A(n3894), .B(n3895), .Z(z2[175]) );
  NANDN U5838 ( .A(xregN_1), .B(zin[174]), .Z(n3895) );
  NAND U5839 ( .A(N179), .B(xregN_1), .Z(n3894) );
  NAND U5840 ( .A(n3896), .B(n3897), .Z(z2[174]) );
  NANDN U5841 ( .A(xregN_1), .B(zin[173]), .Z(n3897) );
  NAND U5842 ( .A(N178), .B(xregN_1), .Z(n3896) );
  NAND U5843 ( .A(n3898), .B(n3899), .Z(z2[173]) );
  NANDN U5844 ( .A(xregN_1), .B(zin[172]), .Z(n3899) );
  NAND U5845 ( .A(N177), .B(xregN_1), .Z(n3898) );
  NAND U5846 ( .A(n3900), .B(n3901), .Z(z2[172]) );
  NANDN U5847 ( .A(xregN_1), .B(zin[171]), .Z(n3901) );
  NAND U5848 ( .A(N176), .B(xregN_1), .Z(n3900) );
  NAND U5849 ( .A(n3902), .B(n3903), .Z(z2[171]) );
  NANDN U5850 ( .A(xregN_1), .B(zin[170]), .Z(n3903) );
  NAND U5851 ( .A(N175), .B(xregN_1), .Z(n3902) );
  NAND U5852 ( .A(n3904), .B(n3905), .Z(z2[170]) );
  NANDN U5853 ( .A(xregN_1), .B(zin[169]), .Z(n3905) );
  NAND U5854 ( .A(N174), .B(xregN_1), .Z(n3904) );
  NAND U5855 ( .A(n3906), .B(n3907), .Z(z2[16]) );
  NANDN U5856 ( .A(xregN_1), .B(zin[15]), .Z(n3907) );
  NAND U5857 ( .A(N20), .B(xregN_1), .Z(n3906) );
  NAND U5858 ( .A(n3908), .B(n3909), .Z(z2[169]) );
  NANDN U5859 ( .A(xregN_1), .B(zin[168]), .Z(n3909) );
  NAND U5860 ( .A(N173), .B(xregN_1), .Z(n3908) );
  NAND U5861 ( .A(n3910), .B(n3911), .Z(z2[168]) );
  NANDN U5862 ( .A(xregN_1), .B(zin[167]), .Z(n3911) );
  NAND U5863 ( .A(N172), .B(xregN_1), .Z(n3910) );
  NAND U5864 ( .A(n3912), .B(n3913), .Z(z2[167]) );
  NANDN U5865 ( .A(xregN_1), .B(zin[166]), .Z(n3913) );
  NAND U5866 ( .A(N171), .B(xregN_1), .Z(n3912) );
  NAND U5867 ( .A(n3914), .B(n3915), .Z(z2[166]) );
  NANDN U5868 ( .A(xregN_1), .B(zin[165]), .Z(n3915) );
  NAND U5869 ( .A(N170), .B(xregN_1), .Z(n3914) );
  NAND U5870 ( .A(n3916), .B(n3917), .Z(z2[165]) );
  NANDN U5871 ( .A(xregN_1), .B(zin[164]), .Z(n3917) );
  NAND U5872 ( .A(N169), .B(xregN_1), .Z(n3916) );
  NAND U5873 ( .A(n3918), .B(n3919), .Z(z2[164]) );
  NANDN U5874 ( .A(xregN_1), .B(zin[163]), .Z(n3919) );
  NAND U5875 ( .A(N168), .B(xregN_1), .Z(n3918) );
  NAND U5876 ( .A(n3920), .B(n3921), .Z(z2[163]) );
  NANDN U5877 ( .A(xregN_1), .B(zin[162]), .Z(n3921) );
  NAND U5878 ( .A(N167), .B(xregN_1), .Z(n3920) );
  NAND U5879 ( .A(n3922), .B(n3923), .Z(z2[162]) );
  NANDN U5880 ( .A(xregN_1), .B(zin[161]), .Z(n3923) );
  NAND U5881 ( .A(N166), .B(xregN_1), .Z(n3922) );
  NAND U5882 ( .A(n3924), .B(n3925), .Z(z2[161]) );
  NANDN U5883 ( .A(xregN_1), .B(zin[160]), .Z(n3925) );
  NAND U5884 ( .A(N165), .B(xregN_1), .Z(n3924) );
  NAND U5885 ( .A(n3926), .B(n3927), .Z(z2[160]) );
  NANDN U5886 ( .A(xregN_1), .B(zin[159]), .Z(n3927) );
  NAND U5887 ( .A(N164), .B(xregN_1), .Z(n3926) );
  NAND U5888 ( .A(n3928), .B(n3929), .Z(z2[15]) );
  NANDN U5889 ( .A(xregN_1), .B(zin[14]), .Z(n3929) );
  NAND U5890 ( .A(N19), .B(xregN_1), .Z(n3928) );
  NAND U5891 ( .A(n3930), .B(n3931), .Z(z2[159]) );
  NANDN U5892 ( .A(xregN_1), .B(zin[158]), .Z(n3931) );
  NAND U5893 ( .A(N163), .B(xregN_1), .Z(n3930) );
  NAND U5894 ( .A(n3932), .B(n3933), .Z(z2[158]) );
  NANDN U5895 ( .A(xregN_1), .B(zin[157]), .Z(n3933) );
  NAND U5896 ( .A(N162), .B(xregN_1), .Z(n3932) );
  NAND U5897 ( .A(n3934), .B(n3935), .Z(z2[157]) );
  NANDN U5898 ( .A(xregN_1), .B(zin[156]), .Z(n3935) );
  NAND U5899 ( .A(N161), .B(xregN_1), .Z(n3934) );
  NAND U5900 ( .A(n3936), .B(n3937), .Z(z2[156]) );
  NANDN U5901 ( .A(xregN_1), .B(zin[155]), .Z(n3937) );
  NAND U5902 ( .A(N160), .B(xregN_1), .Z(n3936) );
  NAND U5903 ( .A(n3938), .B(n3939), .Z(z2[155]) );
  NANDN U5904 ( .A(xregN_1), .B(zin[154]), .Z(n3939) );
  NAND U5905 ( .A(N159), .B(xregN_1), .Z(n3938) );
  NAND U5906 ( .A(n3940), .B(n3941), .Z(z2[154]) );
  NANDN U5907 ( .A(xregN_1), .B(zin[153]), .Z(n3941) );
  NAND U5908 ( .A(N158), .B(xregN_1), .Z(n3940) );
  NAND U5909 ( .A(n3942), .B(n3943), .Z(z2[153]) );
  NANDN U5910 ( .A(xregN_1), .B(zin[152]), .Z(n3943) );
  NAND U5911 ( .A(N157), .B(xregN_1), .Z(n3942) );
  NAND U5912 ( .A(n3944), .B(n3945), .Z(z2[152]) );
  NANDN U5913 ( .A(xregN_1), .B(zin[151]), .Z(n3945) );
  NAND U5914 ( .A(N156), .B(xregN_1), .Z(n3944) );
  NAND U5915 ( .A(n3946), .B(n3947), .Z(z2[151]) );
  NANDN U5916 ( .A(xregN_1), .B(zin[150]), .Z(n3947) );
  NAND U5917 ( .A(N155), .B(xregN_1), .Z(n3946) );
  NAND U5918 ( .A(n3948), .B(n3949), .Z(z2[150]) );
  NANDN U5919 ( .A(xregN_1), .B(zin[149]), .Z(n3949) );
  NAND U5920 ( .A(N154), .B(xregN_1), .Z(n3948) );
  NAND U5921 ( .A(n3950), .B(n3951), .Z(z2[14]) );
  NANDN U5922 ( .A(xregN_1), .B(zin[13]), .Z(n3951) );
  NAND U5923 ( .A(N18), .B(xregN_1), .Z(n3950) );
  NAND U5924 ( .A(n3952), .B(n3953), .Z(z2[149]) );
  NANDN U5925 ( .A(xregN_1), .B(zin[148]), .Z(n3953) );
  NAND U5926 ( .A(N153), .B(xregN_1), .Z(n3952) );
  NAND U5927 ( .A(n3954), .B(n3955), .Z(z2[148]) );
  NANDN U5928 ( .A(xregN_1), .B(zin[147]), .Z(n3955) );
  NAND U5929 ( .A(N152), .B(xregN_1), .Z(n3954) );
  NAND U5930 ( .A(n3956), .B(n3957), .Z(z2[147]) );
  NANDN U5931 ( .A(xregN_1), .B(zin[146]), .Z(n3957) );
  NAND U5932 ( .A(N151), .B(xregN_1), .Z(n3956) );
  NAND U5933 ( .A(n3958), .B(n3959), .Z(z2[146]) );
  NANDN U5934 ( .A(xregN_1), .B(zin[145]), .Z(n3959) );
  NAND U5935 ( .A(N150), .B(xregN_1), .Z(n3958) );
  NAND U5936 ( .A(n3960), .B(n3961), .Z(z2[145]) );
  NANDN U5937 ( .A(xregN_1), .B(zin[144]), .Z(n3961) );
  NAND U5938 ( .A(N149), .B(xregN_1), .Z(n3960) );
  NAND U5939 ( .A(n3962), .B(n3963), .Z(z2[144]) );
  NANDN U5940 ( .A(xregN_1), .B(zin[143]), .Z(n3963) );
  NAND U5941 ( .A(N148), .B(xregN_1), .Z(n3962) );
  NAND U5942 ( .A(n3964), .B(n3965), .Z(z2[143]) );
  NANDN U5943 ( .A(xregN_1), .B(zin[142]), .Z(n3965) );
  NAND U5944 ( .A(N147), .B(xregN_1), .Z(n3964) );
  NAND U5945 ( .A(n3966), .B(n3967), .Z(z2[142]) );
  NANDN U5946 ( .A(xregN_1), .B(zin[141]), .Z(n3967) );
  NAND U5947 ( .A(N146), .B(xregN_1), .Z(n3966) );
  NAND U5948 ( .A(n3968), .B(n3969), .Z(z2[141]) );
  NANDN U5949 ( .A(xregN_1), .B(zin[140]), .Z(n3969) );
  NAND U5950 ( .A(N145), .B(xregN_1), .Z(n3968) );
  NAND U5951 ( .A(n3970), .B(n3971), .Z(z2[140]) );
  NANDN U5952 ( .A(xregN_1), .B(zin[139]), .Z(n3971) );
  NAND U5953 ( .A(N144), .B(xregN_1), .Z(n3970) );
  NAND U5954 ( .A(n3972), .B(n3973), .Z(z2[13]) );
  NANDN U5955 ( .A(xregN_1), .B(zin[12]), .Z(n3973) );
  NAND U5956 ( .A(N17), .B(xregN_1), .Z(n3972) );
  NAND U5957 ( .A(n3974), .B(n3975), .Z(z2[139]) );
  NANDN U5958 ( .A(xregN_1), .B(zin[138]), .Z(n3975) );
  NAND U5959 ( .A(N143), .B(xregN_1), .Z(n3974) );
  NAND U5960 ( .A(n3976), .B(n3977), .Z(z2[138]) );
  NANDN U5961 ( .A(xregN_1), .B(zin[137]), .Z(n3977) );
  NAND U5962 ( .A(N142), .B(xregN_1), .Z(n3976) );
  NAND U5963 ( .A(n3978), .B(n3979), .Z(z2[137]) );
  NANDN U5964 ( .A(xregN_1), .B(zin[136]), .Z(n3979) );
  NAND U5965 ( .A(N141), .B(xregN_1), .Z(n3978) );
  NAND U5966 ( .A(n3980), .B(n3981), .Z(z2[136]) );
  NANDN U5967 ( .A(xregN_1), .B(zin[135]), .Z(n3981) );
  NAND U5968 ( .A(N140), .B(xregN_1), .Z(n3980) );
  NAND U5969 ( .A(n3982), .B(n3983), .Z(z2[135]) );
  NANDN U5970 ( .A(xregN_1), .B(zin[134]), .Z(n3983) );
  NAND U5971 ( .A(N139), .B(xregN_1), .Z(n3982) );
  NAND U5972 ( .A(n3984), .B(n3985), .Z(z2[134]) );
  NANDN U5973 ( .A(xregN_1), .B(zin[133]), .Z(n3985) );
  NAND U5974 ( .A(N138), .B(xregN_1), .Z(n3984) );
  NAND U5975 ( .A(n3986), .B(n3987), .Z(z2[133]) );
  NANDN U5976 ( .A(xregN_1), .B(zin[132]), .Z(n3987) );
  NAND U5977 ( .A(N137), .B(xregN_1), .Z(n3986) );
  NAND U5978 ( .A(n3988), .B(n3989), .Z(z2[132]) );
  NANDN U5979 ( .A(xregN_1), .B(zin[131]), .Z(n3989) );
  NAND U5980 ( .A(N136), .B(xregN_1), .Z(n3988) );
  NAND U5981 ( .A(n3990), .B(n3991), .Z(z2[131]) );
  NANDN U5982 ( .A(xregN_1), .B(zin[130]), .Z(n3991) );
  NAND U5983 ( .A(N135), .B(xregN_1), .Z(n3990) );
  NAND U5984 ( .A(n3992), .B(n3993), .Z(z2[130]) );
  NANDN U5985 ( .A(xregN_1), .B(zin[129]), .Z(n3993) );
  NAND U5986 ( .A(N134), .B(xregN_1), .Z(n3992) );
  NAND U5987 ( .A(n3994), .B(n3995), .Z(z2[12]) );
  NANDN U5988 ( .A(xregN_1), .B(zin[11]), .Z(n3995) );
  NAND U5989 ( .A(N16), .B(xregN_1), .Z(n3994) );
  NAND U5990 ( .A(n3996), .B(n3997), .Z(z2[129]) );
  NANDN U5991 ( .A(xregN_1), .B(zin[128]), .Z(n3997) );
  NAND U5992 ( .A(N133), .B(xregN_1), .Z(n3996) );
  NAND U5993 ( .A(n3998), .B(n3999), .Z(z2[128]) );
  NANDN U5994 ( .A(xregN_1), .B(zin[127]), .Z(n3999) );
  NAND U5995 ( .A(N132), .B(xregN_1), .Z(n3998) );
  NAND U5996 ( .A(n4000), .B(n4001), .Z(z2[127]) );
  NANDN U5997 ( .A(xregN_1), .B(zin[126]), .Z(n4001) );
  NAND U5998 ( .A(N131), .B(xregN_1), .Z(n4000) );
  NAND U5999 ( .A(n4002), .B(n4003), .Z(z2[126]) );
  NANDN U6000 ( .A(xregN_1), .B(zin[125]), .Z(n4003) );
  NAND U6001 ( .A(N130), .B(xregN_1), .Z(n4002) );
  NAND U6002 ( .A(n4004), .B(n4005), .Z(z2[125]) );
  NANDN U6003 ( .A(xregN_1), .B(zin[124]), .Z(n4005) );
  NAND U6004 ( .A(N129), .B(xregN_1), .Z(n4004) );
  NAND U6005 ( .A(n4006), .B(n4007), .Z(z2[124]) );
  NANDN U6006 ( .A(xregN_1), .B(zin[123]), .Z(n4007) );
  NAND U6007 ( .A(N128), .B(xregN_1), .Z(n4006) );
  NAND U6008 ( .A(n4008), .B(n4009), .Z(z2[123]) );
  NANDN U6009 ( .A(xregN_1), .B(zin[122]), .Z(n4009) );
  NAND U6010 ( .A(N127), .B(xregN_1), .Z(n4008) );
  NAND U6011 ( .A(n4010), .B(n4011), .Z(z2[122]) );
  NANDN U6012 ( .A(xregN_1), .B(zin[121]), .Z(n4011) );
  NAND U6013 ( .A(N126), .B(xregN_1), .Z(n4010) );
  NAND U6014 ( .A(n4012), .B(n4013), .Z(z2[121]) );
  NANDN U6015 ( .A(xregN_1), .B(zin[120]), .Z(n4013) );
  NAND U6016 ( .A(N125), .B(xregN_1), .Z(n4012) );
  NAND U6017 ( .A(n4014), .B(n4015), .Z(z2[120]) );
  NANDN U6018 ( .A(xregN_1), .B(zin[119]), .Z(n4015) );
  NAND U6019 ( .A(N124), .B(xregN_1), .Z(n4014) );
  NAND U6020 ( .A(n4016), .B(n4017), .Z(z2[11]) );
  NANDN U6021 ( .A(xregN_1), .B(zin[10]), .Z(n4017) );
  NAND U6022 ( .A(N15), .B(xregN_1), .Z(n4016) );
  NAND U6023 ( .A(n4018), .B(n4019), .Z(z2[119]) );
  NANDN U6024 ( .A(xregN_1), .B(zin[118]), .Z(n4019) );
  NAND U6025 ( .A(N123), .B(xregN_1), .Z(n4018) );
  NAND U6026 ( .A(n4020), .B(n4021), .Z(z2[118]) );
  NANDN U6027 ( .A(xregN_1), .B(zin[117]), .Z(n4021) );
  NAND U6028 ( .A(N122), .B(xregN_1), .Z(n4020) );
  NAND U6029 ( .A(n4022), .B(n4023), .Z(z2[117]) );
  NANDN U6030 ( .A(xregN_1), .B(zin[116]), .Z(n4023) );
  NAND U6031 ( .A(N121), .B(xregN_1), .Z(n4022) );
  NAND U6032 ( .A(n4024), .B(n4025), .Z(z2[116]) );
  NANDN U6033 ( .A(xregN_1), .B(zin[115]), .Z(n4025) );
  NAND U6034 ( .A(N120), .B(xregN_1), .Z(n4024) );
  NAND U6035 ( .A(n4026), .B(n4027), .Z(z2[115]) );
  NANDN U6036 ( .A(xregN_1), .B(zin[114]), .Z(n4027) );
  NAND U6037 ( .A(N119), .B(xregN_1), .Z(n4026) );
  NAND U6038 ( .A(n4028), .B(n4029), .Z(z2[114]) );
  NANDN U6039 ( .A(xregN_1), .B(zin[113]), .Z(n4029) );
  NAND U6040 ( .A(N118), .B(xregN_1), .Z(n4028) );
  NAND U6041 ( .A(n4030), .B(n4031), .Z(z2[113]) );
  NANDN U6042 ( .A(xregN_1), .B(zin[112]), .Z(n4031) );
  NAND U6043 ( .A(N117), .B(xregN_1), .Z(n4030) );
  NAND U6044 ( .A(n4032), .B(n4033), .Z(z2[112]) );
  NANDN U6045 ( .A(xregN_1), .B(zin[111]), .Z(n4033) );
  NAND U6046 ( .A(N116), .B(xregN_1), .Z(n4032) );
  NAND U6047 ( .A(n4034), .B(n4035), .Z(z2[111]) );
  NANDN U6048 ( .A(xregN_1), .B(zin[110]), .Z(n4035) );
  NAND U6049 ( .A(N115), .B(xregN_1), .Z(n4034) );
  NAND U6050 ( .A(n4036), .B(n4037), .Z(z2[110]) );
  NANDN U6051 ( .A(xregN_1), .B(zin[109]), .Z(n4037) );
  NAND U6052 ( .A(N114), .B(xregN_1), .Z(n4036) );
  NAND U6053 ( .A(n4038), .B(n4039), .Z(z2[10]) );
  NANDN U6054 ( .A(xregN_1), .B(zin[9]), .Z(n4039) );
  NAND U6055 ( .A(N14), .B(xregN_1), .Z(n4038) );
  NAND U6056 ( .A(n4040), .B(n4041), .Z(z2[109]) );
  NANDN U6057 ( .A(xregN_1), .B(zin[108]), .Z(n4041) );
  NAND U6058 ( .A(N113), .B(xregN_1), .Z(n4040) );
  NAND U6059 ( .A(n4042), .B(n4043), .Z(z2[108]) );
  NANDN U6060 ( .A(xregN_1), .B(zin[107]), .Z(n4043) );
  NAND U6061 ( .A(N112), .B(xregN_1), .Z(n4042) );
  NAND U6062 ( .A(n4044), .B(n4045), .Z(z2[107]) );
  NANDN U6063 ( .A(xregN_1), .B(zin[106]), .Z(n4045) );
  NAND U6064 ( .A(N111), .B(xregN_1), .Z(n4044) );
  NAND U6065 ( .A(n4046), .B(n4047), .Z(z2[106]) );
  NANDN U6066 ( .A(xregN_1), .B(zin[105]), .Z(n4047) );
  NAND U6067 ( .A(N110), .B(xregN_1), .Z(n4046) );
  NAND U6068 ( .A(n4048), .B(n4049), .Z(z2[105]) );
  NANDN U6069 ( .A(xregN_1), .B(zin[104]), .Z(n4049) );
  NAND U6070 ( .A(N109), .B(xregN_1), .Z(n4048) );
  NAND U6071 ( .A(n4050), .B(n4051), .Z(z2[104]) );
  NANDN U6072 ( .A(xregN_1), .B(zin[103]), .Z(n4051) );
  NAND U6073 ( .A(N108), .B(xregN_1), .Z(n4050) );
  NAND U6074 ( .A(n4052), .B(n4053), .Z(z2[103]) );
  NANDN U6075 ( .A(xregN_1), .B(zin[102]), .Z(n4053) );
  NAND U6076 ( .A(N107), .B(xregN_1), .Z(n4052) );
  NAND U6077 ( .A(n4054), .B(n4055), .Z(z2[102]) );
  NANDN U6078 ( .A(xregN_1), .B(zin[101]), .Z(n4055) );
  NAND U6079 ( .A(N106), .B(xregN_1), .Z(n4054) );
  NAND U6080 ( .A(n4056), .B(n4057), .Z(z2[1025]) );
  NANDN U6081 ( .A(xregN_1), .B(zin[1024]), .Z(n4057) );
  NAND U6082 ( .A(N1029), .B(xregN_1), .Z(n4056) );
  NAND U6083 ( .A(n4058), .B(n4059), .Z(z2[1024]) );
  NANDN U6084 ( .A(xregN_1), .B(zin[1023]), .Z(n4059) );
  NAND U6085 ( .A(N1028), .B(xregN_1), .Z(n4058) );
  NAND U6086 ( .A(n4060), .B(n4061), .Z(z2[1023]) );
  NANDN U6087 ( .A(xregN_1), .B(zin[1022]), .Z(n4061) );
  NAND U6088 ( .A(N1027), .B(xregN_1), .Z(n4060) );
  NAND U6089 ( .A(n4062), .B(n4063), .Z(z2[1022]) );
  NANDN U6090 ( .A(xregN_1), .B(zin[1021]), .Z(n4063) );
  NAND U6091 ( .A(N1026), .B(xregN_1), .Z(n4062) );
  NAND U6092 ( .A(n4064), .B(n4065), .Z(z2[1021]) );
  NANDN U6093 ( .A(xregN_1), .B(zin[1020]), .Z(n4065) );
  NAND U6094 ( .A(N1025), .B(xregN_1), .Z(n4064) );
  NAND U6095 ( .A(n4066), .B(n4067), .Z(z2[1020]) );
  NANDN U6096 ( .A(xregN_1), .B(zin[1019]), .Z(n4067) );
  NAND U6097 ( .A(N1024), .B(xregN_1), .Z(n4066) );
  NAND U6098 ( .A(n4068), .B(n4069), .Z(z2[101]) );
  NANDN U6099 ( .A(xregN_1), .B(zin[100]), .Z(n4069) );
  NAND U6100 ( .A(N105), .B(xregN_1), .Z(n4068) );
  NAND U6101 ( .A(n4070), .B(n4071), .Z(z2[1019]) );
  NANDN U6102 ( .A(xregN_1), .B(zin[1018]), .Z(n4071) );
  NAND U6103 ( .A(N1023), .B(xregN_1), .Z(n4070) );
  NAND U6104 ( .A(n4072), .B(n4073), .Z(z2[1018]) );
  NANDN U6105 ( .A(xregN_1), .B(zin[1017]), .Z(n4073) );
  NAND U6106 ( .A(N1022), .B(xregN_1), .Z(n4072) );
  NAND U6107 ( .A(n4074), .B(n4075), .Z(z2[1017]) );
  NANDN U6108 ( .A(xregN_1), .B(zin[1016]), .Z(n4075) );
  NAND U6109 ( .A(N1021), .B(xregN_1), .Z(n4074) );
  NAND U6110 ( .A(n4076), .B(n4077), .Z(z2[1016]) );
  NANDN U6111 ( .A(xregN_1), .B(zin[1015]), .Z(n4077) );
  NAND U6112 ( .A(N1020), .B(xregN_1), .Z(n4076) );
  NAND U6113 ( .A(n4078), .B(n4079), .Z(z2[1015]) );
  NANDN U6114 ( .A(xregN_1), .B(zin[1014]), .Z(n4079) );
  NAND U6115 ( .A(N1019), .B(xregN_1), .Z(n4078) );
  NAND U6116 ( .A(n4080), .B(n4081), .Z(z2[1014]) );
  NANDN U6117 ( .A(xregN_1), .B(zin[1013]), .Z(n4081) );
  NAND U6118 ( .A(N1018), .B(xregN_1), .Z(n4080) );
  NAND U6119 ( .A(n4082), .B(n4083), .Z(z2[1013]) );
  NANDN U6120 ( .A(xregN_1), .B(zin[1012]), .Z(n4083) );
  NAND U6121 ( .A(N1017), .B(xregN_1), .Z(n4082) );
  NAND U6122 ( .A(n4084), .B(n4085), .Z(z2[1012]) );
  NANDN U6123 ( .A(xregN_1), .B(zin[1011]), .Z(n4085) );
  NAND U6124 ( .A(N1016), .B(xregN_1), .Z(n4084) );
  NAND U6125 ( .A(n4086), .B(n4087), .Z(z2[1011]) );
  NANDN U6126 ( .A(xregN_1), .B(zin[1010]), .Z(n4087) );
  NAND U6127 ( .A(N1015), .B(xregN_1), .Z(n4086) );
  NAND U6128 ( .A(n4088), .B(n4089), .Z(z2[1010]) );
  NANDN U6129 ( .A(xregN_1), .B(zin[1009]), .Z(n4089) );
  NAND U6130 ( .A(N1014), .B(xregN_1), .Z(n4088) );
  NAND U6131 ( .A(n4090), .B(n4091), .Z(z2[100]) );
  NANDN U6132 ( .A(xregN_1), .B(zin[99]), .Z(n4091) );
  NAND U6133 ( .A(N104), .B(xregN_1), .Z(n4090) );
  NAND U6134 ( .A(n4092), .B(n4093), .Z(z2[1009]) );
  NANDN U6135 ( .A(xregN_1), .B(zin[1008]), .Z(n4093) );
  NAND U6136 ( .A(N1013), .B(xregN_1), .Z(n4092) );
  NAND U6137 ( .A(n4094), .B(n4095), .Z(z2[1008]) );
  NANDN U6138 ( .A(xregN_1), .B(zin[1007]), .Z(n4095) );
  NAND U6139 ( .A(N1012), .B(xregN_1), .Z(n4094) );
  NAND U6140 ( .A(n4096), .B(n4097), .Z(z2[1007]) );
  NANDN U6141 ( .A(xregN_1), .B(zin[1006]), .Z(n4097) );
  NAND U6142 ( .A(N1011), .B(xregN_1), .Z(n4096) );
  NAND U6143 ( .A(n4098), .B(n4099), .Z(z2[1006]) );
  NANDN U6144 ( .A(xregN_1), .B(zin[1005]), .Z(n4099) );
  NAND U6145 ( .A(N1010), .B(xregN_1), .Z(n4098) );
  NAND U6146 ( .A(n4100), .B(n4101), .Z(z2[1005]) );
  NANDN U6147 ( .A(xregN_1), .B(zin[1004]), .Z(n4101) );
  NAND U6148 ( .A(N1009), .B(xregN_1), .Z(n4100) );
  NAND U6149 ( .A(n4102), .B(n4103), .Z(z2[1004]) );
  NANDN U6150 ( .A(xregN_1), .B(zin[1003]), .Z(n4103) );
  NAND U6151 ( .A(N1008), .B(xregN_1), .Z(n4102) );
  NAND U6152 ( .A(n4104), .B(n4105), .Z(z2[1003]) );
  NANDN U6153 ( .A(xregN_1), .B(zin[1002]), .Z(n4105) );
  NAND U6154 ( .A(N1007), .B(xregN_1), .Z(n4104) );
  NAND U6155 ( .A(n4106), .B(n4107), .Z(z2[1002]) );
  NANDN U6156 ( .A(xregN_1), .B(zin[1001]), .Z(n4107) );
  NAND U6157 ( .A(N1006), .B(xregN_1), .Z(n4106) );
  NAND U6158 ( .A(n4108), .B(n4109), .Z(z2[1001]) );
  NANDN U6159 ( .A(xregN_1), .B(zin[1000]), .Z(n4109) );
  NAND U6160 ( .A(N1005), .B(xregN_1), .Z(n4108) );
  NAND U6161 ( .A(n4110), .B(n4111), .Z(z2[1000]) );
  NANDN U6162 ( .A(xregN_1), .B(zin[999]), .Z(n4111) );
  NAND U6163 ( .A(N1004), .B(xregN_1), .Z(n4110) );
  AND U6164 ( .A(N4), .B(xregN_1), .Z(z2[0]) );
endmodule


module modmult_N1024_CC1024 ( clk, rst, start, x, y, n, o );
  input [1023:0] x;
  input [1023:0] y;
  input [1023:0] n;
  output [1023:0] o;
  input clk, rst, start;
  wire   \zout[0][1025] , \zout[0][1024] , \zin[0][1025] , \zin[0][1024] ,
         \zin[0][1023] , \zin[0][1022] , \zin[0][1021] , \zin[0][1020] ,
         \zin[0][1019] , \zin[0][1018] , \zin[0][1017] , \zin[0][1016] ,
         \zin[0][1015] , \zin[0][1014] , \zin[0][1013] , \zin[0][1012] ,
         \zin[0][1011] , \zin[0][1010] , \zin[0][1009] , \zin[0][1008] ,
         \zin[0][1007] , \zin[0][1006] , \zin[0][1005] , \zin[0][1004] ,
         \zin[0][1003] , \zin[0][1002] , \zin[0][1001] , \zin[0][1000] ,
         \zin[0][999] , \zin[0][998] , \zin[0][997] , \zin[0][996] ,
         \zin[0][995] , \zin[0][994] , \zin[0][993] , \zin[0][992] ,
         \zin[0][991] , \zin[0][990] , \zin[0][989] , \zin[0][988] ,
         \zin[0][987] , \zin[0][986] , \zin[0][985] , \zin[0][984] ,
         \zin[0][983] , \zin[0][982] , \zin[0][981] , \zin[0][980] ,
         \zin[0][979] , \zin[0][978] , \zin[0][977] , \zin[0][976] ,
         \zin[0][975] , \zin[0][974] , \zin[0][973] , \zin[0][972] ,
         \zin[0][971] , \zin[0][970] , \zin[0][969] , \zin[0][968] ,
         \zin[0][967] , \zin[0][966] , \zin[0][965] , \zin[0][964] ,
         \zin[0][963] , \zin[0][962] , \zin[0][961] , \zin[0][960] ,
         \zin[0][959] , \zin[0][958] , \zin[0][957] , \zin[0][956] ,
         \zin[0][955] , \zin[0][954] , \zin[0][953] , \zin[0][952] ,
         \zin[0][951] , \zin[0][950] , \zin[0][949] , \zin[0][948] ,
         \zin[0][947] , \zin[0][946] , \zin[0][945] , \zin[0][944] ,
         \zin[0][943] , \zin[0][942] , \zin[0][941] , \zin[0][940] ,
         \zin[0][939] , \zin[0][938] , \zin[0][937] , \zin[0][936] ,
         \zin[0][935] , \zin[0][934] , \zin[0][933] , \zin[0][932] ,
         \zin[0][931] , \zin[0][930] , \zin[0][929] , \zin[0][928] ,
         \zin[0][927] , \zin[0][926] , \zin[0][925] , \zin[0][924] ,
         \zin[0][923] , \zin[0][922] , \zin[0][921] , \zin[0][920] ,
         \zin[0][919] , \zin[0][918] , \zin[0][917] , \zin[0][916] ,
         \zin[0][915] , \zin[0][914] , \zin[0][913] , \zin[0][912] ,
         \zin[0][911] , \zin[0][910] , \zin[0][909] , \zin[0][908] ,
         \zin[0][907] , \zin[0][906] , \zin[0][905] , \zin[0][904] ,
         \zin[0][903] , \zin[0][902] , \zin[0][901] , \zin[0][900] ,
         \zin[0][899] , \zin[0][898] , \zin[0][897] , \zin[0][896] ,
         \zin[0][895] , \zin[0][894] , \zin[0][893] , \zin[0][892] ,
         \zin[0][891] , \zin[0][890] , \zin[0][889] , \zin[0][888] ,
         \zin[0][887] , \zin[0][886] , \zin[0][885] , \zin[0][884] ,
         \zin[0][883] , \zin[0][882] , \zin[0][881] , \zin[0][880] ,
         \zin[0][879] , \zin[0][878] , \zin[0][877] , \zin[0][876] ,
         \zin[0][875] , \zin[0][874] , \zin[0][873] , \zin[0][872] ,
         \zin[0][871] , \zin[0][870] , \zin[0][869] , \zin[0][868] ,
         \zin[0][867] , \zin[0][866] , \zin[0][865] , \zin[0][864] ,
         \zin[0][863] , \zin[0][862] , \zin[0][861] , \zin[0][860] ,
         \zin[0][859] , \zin[0][858] , \zin[0][857] , \zin[0][856] ,
         \zin[0][855] , \zin[0][854] , \zin[0][853] , \zin[0][852] ,
         \zin[0][851] , \zin[0][850] , \zin[0][849] , \zin[0][848] ,
         \zin[0][847] , \zin[0][846] , \zin[0][845] , \zin[0][844] ,
         \zin[0][843] , \zin[0][842] , \zin[0][841] , \zin[0][840] ,
         \zin[0][839] , \zin[0][838] , \zin[0][837] , \zin[0][836] ,
         \zin[0][835] , \zin[0][834] , \zin[0][833] , \zin[0][832] ,
         \zin[0][831] , \zin[0][830] , \zin[0][829] , \zin[0][828] ,
         \zin[0][827] , \zin[0][826] , \zin[0][825] , \zin[0][824] ,
         \zin[0][823] , \zin[0][822] , \zin[0][821] , \zin[0][820] ,
         \zin[0][819] , \zin[0][818] , \zin[0][817] , \zin[0][816] ,
         \zin[0][815] , \zin[0][814] , \zin[0][813] , \zin[0][812] ,
         \zin[0][811] , \zin[0][810] , \zin[0][809] , \zin[0][808] ,
         \zin[0][807] , \zin[0][806] , \zin[0][805] , \zin[0][804] ,
         \zin[0][803] , \zin[0][802] , \zin[0][801] , \zin[0][800] ,
         \zin[0][799] , \zin[0][798] , \zin[0][797] , \zin[0][796] ,
         \zin[0][795] , \zin[0][794] , \zin[0][793] , \zin[0][792] ,
         \zin[0][791] , \zin[0][790] , \zin[0][789] , \zin[0][788] ,
         \zin[0][787] , \zin[0][786] , \zin[0][785] , \zin[0][784] ,
         \zin[0][783] , \zin[0][782] , \zin[0][781] , \zin[0][780] ,
         \zin[0][779] , \zin[0][778] , \zin[0][777] , \zin[0][776] ,
         \zin[0][775] , \zin[0][774] , \zin[0][773] , \zin[0][772] ,
         \zin[0][771] , \zin[0][770] , \zin[0][769] , \zin[0][768] ,
         \zin[0][767] , \zin[0][766] , \zin[0][765] , \zin[0][764] ,
         \zin[0][763] , \zin[0][762] , \zin[0][761] , \zin[0][760] ,
         \zin[0][759] , \zin[0][758] , \zin[0][757] , \zin[0][756] ,
         \zin[0][755] , \zin[0][754] , \zin[0][753] , \zin[0][752] ,
         \zin[0][751] , \zin[0][750] , \zin[0][749] , \zin[0][748] ,
         \zin[0][747] , \zin[0][746] , \zin[0][745] , \zin[0][744] ,
         \zin[0][743] , \zin[0][742] , \zin[0][741] , \zin[0][740] ,
         \zin[0][739] , \zin[0][738] , \zin[0][737] , \zin[0][736] ,
         \zin[0][735] , \zin[0][734] , \zin[0][733] , \zin[0][732] ,
         \zin[0][731] , \zin[0][730] , \zin[0][729] , \zin[0][728] ,
         \zin[0][727] , \zin[0][726] , \zin[0][725] , \zin[0][724] ,
         \zin[0][723] , \zin[0][722] , \zin[0][721] , \zin[0][720] ,
         \zin[0][719] , \zin[0][718] , \zin[0][717] , \zin[0][716] ,
         \zin[0][715] , \zin[0][714] , \zin[0][713] , \zin[0][712] ,
         \zin[0][711] , \zin[0][710] , \zin[0][709] , \zin[0][708] ,
         \zin[0][707] , \zin[0][706] , \zin[0][705] , \zin[0][704] ,
         \zin[0][703] , \zin[0][702] , \zin[0][701] , \zin[0][700] ,
         \zin[0][699] , \zin[0][698] , \zin[0][697] , \zin[0][696] ,
         \zin[0][695] , \zin[0][694] , \zin[0][693] , \zin[0][692] ,
         \zin[0][691] , \zin[0][690] , \zin[0][689] , \zin[0][688] ,
         \zin[0][687] , \zin[0][686] , \zin[0][685] , \zin[0][684] ,
         \zin[0][683] , \zin[0][682] , \zin[0][681] , \zin[0][680] ,
         \zin[0][679] , \zin[0][678] , \zin[0][677] , \zin[0][676] ,
         \zin[0][675] , \zin[0][674] , \zin[0][673] , \zin[0][672] ,
         \zin[0][671] , \zin[0][670] , \zin[0][669] , \zin[0][668] ,
         \zin[0][667] , \zin[0][666] , \zin[0][665] , \zin[0][664] ,
         \zin[0][663] , \zin[0][662] , \zin[0][661] , \zin[0][660] ,
         \zin[0][659] , \zin[0][658] , \zin[0][657] , \zin[0][656] ,
         \zin[0][655] , \zin[0][654] , \zin[0][653] , \zin[0][652] ,
         \zin[0][651] , \zin[0][650] , \zin[0][649] , \zin[0][648] ,
         \zin[0][647] , \zin[0][646] , \zin[0][645] , \zin[0][644] ,
         \zin[0][643] , \zin[0][642] , \zin[0][641] , \zin[0][640] ,
         \zin[0][639] , \zin[0][638] , \zin[0][637] , \zin[0][636] ,
         \zin[0][635] , \zin[0][634] , \zin[0][633] , \zin[0][632] ,
         \zin[0][631] , \zin[0][630] , \zin[0][629] , \zin[0][628] ,
         \zin[0][627] , \zin[0][626] , \zin[0][625] , \zin[0][624] ,
         \zin[0][623] , \zin[0][622] , \zin[0][621] , \zin[0][620] ,
         \zin[0][619] , \zin[0][618] , \zin[0][617] , \zin[0][616] ,
         \zin[0][615] , \zin[0][614] , \zin[0][613] , \zin[0][612] ,
         \zin[0][611] , \zin[0][610] , \zin[0][609] , \zin[0][608] ,
         \zin[0][607] , \zin[0][606] , \zin[0][605] , \zin[0][604] ,
         \zin[0][603] , \zin[0][602] , \zin[0][601] , \zin[0][600] ,
         \zin[0][599] , \zin[0][598] , \zin[0][597] , \zin[0][596] ,
         \zin[0][595] , \zin[0][594] , \zin[0][593] , \zin[0][592] ,
         \zin[0][591] , \zin[0][590] , \zin[0][589] , \zin[0][588] ,
         \zin[0][587] , \zin[0][586] , \zin[0][585] , \zin[0][584] ,
         \zin[0][583] , \zin[0][582] , \zin[0][581] , \zin[0][580] ,
         \zin[0][579] , \zin[0][578] , \zin[0][577] , \zin[0][576] ,
         \zin[0][575] , \zin[0][574] , \zin[0][573] , \zin[0][572] ,
         \zin[0][571] , \zin[0][570] , \zin[0][569] , \zin[0][568] ,
         \zin[0][567] , \zin[0][566] , \zin[0][565] , \zin[0][564] ,
         \zin[0][563] , \zin[0][562] , \zin[0][561] , \zin[0][560] ,
         \zin[0][559] , \zin[0][558] , \zin[0][557] , \zin[0][556] ,
         \zin[0][555] , \zin[0][554] , \zin[0][553] , \zin[0][552] ,
         \zin[0][551] , \zin[0][550] , \zin[0][549] , \zin[0][548] ,
         \zin[0][547] , \zin[0][546] , \zin[0][545] , \zin[0][544] ,
         \zin[0][543] , \zin[0][542] , \zin[0][541] , \zin[0][540] ,
         \zin[0][539] , \zin[0][538] , \zin[0][537] , \zin[0][536] ,
         \zin[0][535] , \zin[0][534] , \zin[0][533] , \zin[0][532] ,
         \zin[0][531] , \zin[0][530] , \zin[0][529] , \zin[0][528] ,
         \zin[0][527] , \zin[0][526] , \zin[0][525] , \zin[0][524] ,
         \zin[0][523] , \zin[0][522] , \zin[0][521] , \zin[0][520] ,
         \zin[0][519] , \zin[0][518] , \zin[0][517] , \zin[0][516] ,
         \zin[0][515] , \zin[0][514] , \zin[0][513] , \zin[0][512] ,
         \zin[0][511] , \zin[0][510] , \zin[0][509] , \zin[0][508] ,
         \zin[0][507] , \zin[0][506] , \zin[0][505] , \zin[0][504] ,
         \zin[0][503] , \zin[0][502] , \zin[0][501] , \zin[0][500] ,
         \zin[0][499] , \zin[0][498] , \zin[0][497] , \zin[0][496] ,
         \zin[0][495] , \zin[0][494] , \zin[0][493] , \zin[0][492] ,
         \zin[0][491] , \zin[0][490] , \zin[0][489] , \zin[0][488] ,
         \zin[0][487] , \zin[0][486] , \zin[0][485] , \zin[0][484] ,
         \zin[0][483] , \zin[0][482] , \zin[0][481] , \zin[0][480] ,
         \zin[0][479] , \zin[0][478] , \zin[0][477] , \zin[0][476] ,
         \zin[0][475] , \zin[0][474] , \zin[0][473] , \zin[0][472] ,
         \zin[0][471] , \zin[0][470] , \zin[0][469] , \zin[0][468] ,
         \zin[0][467] , \zin[0][466] , \zin[0][465] , \zin[0][464] ,
         \zin[0][463] , \zin[0][462] , \zin[0][461] , \zin[0][460] ,
         \zin[0][459] , \zin[0][458] , \zin[0][457] , \zin[0][456] ,
         \zin[0][455] , \zin[0][454] , \zin[0][453] , \zin[0][452] ,
         \zin[0][451] , \zin[0][450] , \zin[0][449] , \zin[0][448] ,
         \zin[0][447] , \zin[0][446] , \zin[0][445] , \zin[0][444] ,
         \zin[0][443] , \zin[0][442] , \zin[0][441] , \zin[0][440] ,
         \zin[0][439] , \zin[0][438] , \zin[0][437] , \zin[0][436] ,
         \zin[0][435] , \zin[0][434] , \zin[0][433] , \zin[0][432] ,
         \zin[0][431] , \zin[0][430] , \zin[0][429] , \zin[0][428] ,
         \zin[0][427] , \zin[0][426] , \zin[0][425] , \zin[0][424] ,
         \zin[0][423] , \zin[0][422] , \zin[0][421] , \zin[0][420] ,
         \zin[0][419] , \zin[0][418] , \zin[0][417] , \zin[0][416] ,
         \zin[0][415] , \zin[0][414] , \zin[0][413] , \zin[0][412] ,
         \zin[0][411] , \zin[0][410] , \zin[0][409] , \zin[0][408] ,
         \zin[0][407] , \zin[0][406] , \zin[0][405] , \zin[0][404] ,
         \zin[0][403] , \zin[0][402] , \zin[0][401] , \zin[0][400] ,
         \zin[0][399] , \zin[0][398] , \zin[0][397] , \zin[0][396] ,
         \zin[0][395] , \zin[0][394] , \zin[0][393] , \zin[0][392] ,
         \zin[0][391] , \zin[0][390] , \zin[0][389] , \zin[0][388] ,
         \zin[0][387] , \zin[0][386] , \zin[0][385] , \zin[0][384] ,
         \zin[0][383] , \zin[0][382] , \zin[0][381] , \zin[0][380] ,
         \zin[0][379] , \zin[0][378] , \zin[0][377] , \zin[0][376] ,
         \zin[0][375] , \zin[0][374] , \zin[0][373] , \zin[0][372] ,
         \zin[0][371] , \zin[0][370] , \zin[0][369] , \zin[0][368] ,
         \zin[0][367] , \zin[0][366] , \zin[0][365] , \zin[0][364] ,
         \zin[0][363] , \zin[0][362] , \zin[0][361] , \zin[0][360] ,
         \zin[0][359] , \zin[0][358] , \zin[0][357] , \zin[0][356] ,
         \zin[0][355] , \zin[0][354] , \zin[0][353] , \zin[0][352] ,
         \zin[0][351] , \zin[0][350] , \zin[0][349] , \zin[0][348] ,
         \zin[0][347] , \zin[0][346] , \zin[0][345] , \zin[0][344] ,
         \zin[0][343] , \zin[0][342] , \zin[0][341] , \zin[0][340] ,
         \zin[0][339] , \zin[0][338] , \zin[0][337] , \zin[0][336] ,
         \zin[0][335] , \zin[0][334] , \zin[0][333] , \zin[0][332] ,
         \zin[0][331] , \zin[0][330] , \zin[0][329] , \zin[0][328] ,
         \zin[0][327] , \zin[0][326] , \zin[0][325] , \zin[0][324] ,
         \zin[0][323] , \zin[0][322] , \zin[0][321] , \zin[0][320] ,
         \zin[0][319] , \zin[0][318] , \zin[0][317] , \zin[0][316] ,
         \zin[0][315] , \zin[0][314] , \zin[0][313] , \zin[0][312] ,
         \zin[0][311] , \zin[0][310] , \zin[0][309] , \zin[0][308] ,
         \zin[0][307] , \zin[0][306] , \zin[0][305] , \zin[0][304] ,
         \zin[0][303] , \zin[0][302] , \zin[0][301] , \zin[0][300] ,
         \zin[0][299] , \zin[0][298] , \zin[0][297] , \zin[0][296] ,
         \zin[0][295] , \zin[0][294] , \zin[0][293] , \zin[0][292] ,
         \zin[0][291] , \zin[0][290] , \zin[0][289] , \zin[0][288] ,
         \zin[0][287] , \zin[0][286] , \zin[0][285] , \zin[0][284] ,
         \zin[0][283] , \zin[0][282] , \zin[0][281] , \zin[0][280] ,
         \zin[0][279] , \zin[0][278] , \zin[0][277] , \zin[0][276] ,
         \zin[0][275] , \zin[0][274] , \zin[0][273] , \zin[0][272] ,
         \zin[0][271] , \zin[0][270] , \zin[0][269] , \zin[0][268] ,
         \zin[0][267] , \zin[0][266] , \zin[0][265] , \zin[0][264] ,
         \zin[0][263] , \zin[0][262] , \zin[0][261] , \zin[0][260] ,
         \zin[0][259] , \zin[0][258] , \zin[0][257] , \zin[0][256] ,
         \zin[0][255] , \zin[0][254] , \zin[0][253] , \zin[0][252] ,
         \zin[0][251] , \zin[0][250] , \zin[0][249] , \zin[0][248] ,
         \zin[0][247] , \zin[0][246] , \zin[0][245] , \zin[0][244] ,
         \zin[0][243] , \zin[0][242] , \zin[0][241] , \zin[0][240] ,
         \zin[0][239] , \zin[0][238] , \zin[0][237] , \zin[0][236] ,
         \zin[0][235] , \zin[0][234] , \zin[0][233] , \zin[0][232] ,
         \zin[0][231] , \zin[0][230] , \zin[0][229] , \zin[0][228] ,
         \zin[0][227] , \zin[0][226] , \zin[0][225] , \zin[0][224] ,
         \zin[0][223] , \zin[0][222] , \zin[0][221] , \zin[0][220] ,
         \zin[0][219] , \zin[0][218] , \zin[0][217] , \zin[0][216] ,
         \zin[0][215] , \zin[0][214] , \zin[0][213] , \zin[0][212] ,
         \zin[0][211] , \zin[0][210] , \zin[0][209] , \zin[0][208] ,
         \zin[0][207] , \zin[0][206] , \zin[0][205] , \zin[0][204] ,
         \zin[0][203] , \zin[0][202] , \zin[0][201] , \zin[0][200] ,
         \zin[0][199] , \zin[0][198] , \zin[0][197] , \zin[0][196] ,
         \zin[0][195] , \zin[0][194] , \zin[0][193] , \zin[0][192] ,
         \zin[0][191] , \zin[0][190] , \zin[0][189] , \zin[0][188] ,
         \zin[0][187] , \zin[0][186] , \zin[0][185] , \zin[0][184] ,
         \zin[0][183] , \zin[0][182] , \zin[0][181] , \zin[0][180] ,
         \zin[0][179] , \zin[0][178] , \zin[0][177] , \zin[0][176] ,
         \zin[0][175] , \zin[0][174] , \zin[0][173] , \zin[0][172] ,
         \zin[0][171] , \zin[0][170] , \zin[0][169] , \zin[0][168] ,
         \zin[0][167] , \zin[0][166] , \zin[0][165] , \zin[0][164] ,
         \zin[0][163] , \zin[0][162] , \zin[0][161] , \zin[0][160] ,
         \zin[0][159] , \zin[0][158] , \zin[0][157] , \zin[0][156] ,
         \zin[0][155] , \zin[0][154] , \zin[0][153] , \zin[0][152] ,
         \zin[0][151] , \zin[0][150] , \zin[0][149] , \zin[0][148] ,
         \zin[0][147] , \zin[0][146] , \zin[0][145] , \zin[0][144] ,
         \zin[0][143] , \zin[0][142] , \zin[0][141] , \zin[0][140] ,
         \zin[0][139] , \zin[0][138] , \zin[0][137] , \zin[0][136] ,
         \zin[0][135] , \zin[0][134] , \zin[0][133] , \zin[0][132] ,
         \zin[0][131] , \zin[0][130] , \zin[0][129] , \zin[0][128] ,
         \zin[0][127] , \zin[0][126] , \zin[0][125] , \zin[0][124] ,
         \zin[0][123] , \zin[0][122] , \zin[0][121] , \zin[0][120] ,
         \zin[0][119] , \zin[0][118] , \zin[0][117] , \zin[0][116] ,
         \zin[0][115] , \zin[0][114] , \zin[0][113] , \zin[0][112] ,
         \zin[0][111] , \zin[0][110] , \zin[0][109] , \zin[0][108] ,
         \zin[0][107] , \zin[0][106] , \zin[0][105] , \zin[0][104] ,
         \zin[0][103] , \zin[0][102] , \zin[0][101] , \zin[0][100] ,
         \zin[0][99] , \zin[0][98] , \zin[0][97] , \zin[0][96] , \zin[0][95] ,
         \zin[0][94] , \zin[0][93] , \zin[0][92] , \zin[0][91] , \zin[0][90] ,
         \zin[0][89] , \zin[0][88] , \zin[0][87] , \zin[0][86] , \zin[0][85] ,
         \zin[0][84] , \zin[0][83] , \zin[0][82] , \zin[0][81] , \zin[0][80] ,
         \zin[0][79] , \zin[0][78] , \zin[0][77] , \zin[0][76] , \zin[0][75] ,
         \zin[0][74] , \zin[0][73] , \zin[0][72] , \zin[0][71] , \zin[0][70] ,
         \zin[0][69] , \zin[0][68] , \zin[0][67] , \zin[0][66] , \zin[0][65] ,
         \zin[0][64] , \zin[0][63] , \zin[0][62] , \zin[0][61] , \zin[0][60] ,
         \zin[0][59] , \zin[0][58] , \zin[0][57] , \zin[0][56] , \zin[0][55] ,
         \zin[0][54] , \zin[0][53] , \zin[0][52] , \zin[0][51] , \zin[0][50] ,
         \zin[0][49] , \zin[0][48] , \zin[0][47] , \zin[0][46] , \zin[0][45] ,
         \zin[0][44] , \zin[0][43] , \zin[0][42] , \zin[0][41] , \zin[0][40] ,
         \zin[0][39] , \zin[0][38] , \zin[0][37] , \zin[0][36] , \zin[0][35] ,
         \zin[0][34] , \zin[0][33] , \zin[0][32] , \zin[0][31] , \zin[0][30] ,
         \zin[0][29] , \zin[0][28] , \zin[0][27] , \zin[0][26] , \zin[0][25] ,
         \zin[0][24] , \zin[0][23] , \zin[0][22] , \zin[0][21] , \zin[0][20] ,
         \zin[0][19] , \zin[0][18] , \zin[0][17] , \zin[0][16] , \zin[0][15] ,
         \zin[0][14] , \zin[0][13] , \zin[0][12] , \zin[0][11] , \zin[0][10] ,
         \zin[0][9] , \zin[0][8] , \zin[0][7] , \zin[0][6] , \zin[0][5] ,
         \zin[0][4] , \zin[0][3] , \zin[0][2] , \zin[0][1] , \zin[0][0] , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047;
  wire   [1025:0] zreg;
  wire   [1023:0] xin;
  wire   [1023:0] xreg;

  DFF \xreg_reg[1]  ( .D(n2047), .CLK(clk), .RST(rst), .Q(xreg[1]) );
  DFF \xreg_reg[2]  ( .D(xin[1]), .CLK(clk), .RST(rst), .Q(xreg[2]) );
  DFF \xreg_reg[3]  ( .D(xin[2]), .CLK(clk), .RST(rst), .Q(xreg[3]) );
  DFF \xreg_reg[4]  ( .D(xin[3]), .CLK(clk), .RST(rst), .Q(xreg[4]) );
  DFF \xreg_reg[5]  ( .D(xin[4]), .CLK(clk), .RST(rst), .Q(xreg[5]) );
  DFF \xreg_reg[6]  ( .D(xin[5]), .CLK(clk), .RST(rst), .Q(xreg[6]) );
  DFF \xreg_reg[7]  ( .D(xin[6]), .CLK(clk), .RST(rst), .Q(xreg[7]) );
  DFF \xreg_reg[8]  ( .D(xin[7]), .CLK(clk), .RST(rst), .Q(xreg[8]) );
  DFF \xreg_reg[9]  ( .D(xin[8]), .CLK(clk), .RST(rst), .Q(xreg[9]) );
  DFF \xreg_reg[10]  ( .D(xin[9]), .CLK(clk), .RST(rst), .Q(xreg[10]) );
  DFF \xreg_reg[11]  ( .D(xin[10]), .CLK(clk), .RST(rst), .Q(xreg[11]) );
  DFF \xreg_reg[12]  ( .D(xin[11]), .CLK(clk), .RST(rst), .Q(xreg[12]) );
  DFF \xreg_reg[13]  ( .D(xin[12]), .CLK(clk), .RST(rst), .Q(xreg[13]) );
  DFF \xreg_reg[14]  ( .D(xin[13]), .CLK(clk), .RST(rst), .Q(xreg[14]) );
  DFF \xreg_reg[15]  ( .D(xin[14]), .CLK(clk), .RST(rst), .Q(xreg[15]) );
  DFF \xreg_reg[16]  ( .D(xin[15]), .CLK(clk), .RST(rst), .Q(xreg[16]) );
  DFF \xreg_reg[17]  ( .D(xin[16]), .CLK(clk), .RST(rst), .Q(xreg[17]) );
  DFF \xreg_reg[18]  ( .D(xin[17]), .CLK(clk), .RST(rst), .Q(xreg[18]) );
  DFF \xreg_reg[19]  ( .D(xin[18]), .CLK(clk), .RST(rst), .Q(xreg[19]) );
  DFF \xreg_reg[20]  ( .D(xin[19]), .CLK(clk), .RST(rst), .Q(xreg[20]) );
  DFF \xreg_reg[21]  ( .D(xin[20]), .CLK(clk), .RST(rst), .Q(xreg[21]) );
  DFF \xreg_reg[22]  ( .D(xin[21]), .CLK(clk), .RST(rst), .Q(xreg[22]) );
  DFF \xreg_reg[23]  ( .D(xin[22]), .CLK(clk), .RST(rst), .Q(xreg[23]) );
  DFF \xreg_reg[24]  ( .D(xin[23]), .CLK(clk), .RST(rst), .Q(xreg[24]) );
  DFF \xreg_reg[25]  ( .D(xin[24]), .CLK(clk), .RST(rst), .Q(xreg[25]) );
  DFF \xreg_reg[26]  ( .D(xin[25]), .CLK(clk), .RST(rst), .Q(xreg[26]) );
  DFF \xreg_reg[27]  ( .D(xin[26]), .CLK(clk), .RST(rst), .Q(xreg[27]) );
  DFF \xreg_reg[28]  ( .D(xin[27]), .CLK(clk), .RST(rst), .Q(xreg[28]) );
  DFF \xreg_reg[29]  ( .D(xin[28]), .CLK(clk), .RST(rst), .Q(xreg[29]) );
  DFF \xreg_reg[30]  ( .D(xin[29]), .CLK(clk), .RST(rst), .Q(xreg[30]) );
  DFF \xreg_reg[31]  ( .D(xin[30]), .CLK(clk), .RST(rst), .Q(xreg[31]) );
  DFF \xreg_reg[32]  ( .D(xin[31]), .CLK(clk), .RST(rst), .Q(xreg[32]) );
  DFF \xreg_reg[33]  ( .D(xin[32]), .CLK(clk), .RST(rst), .Q(xreg[33]) );
  DFF \xreg_reg[34]  ( .D(xin[33]), .CLK(clk), .RST(rst), .Q(xreg[34]) );
  DFF \xreg_reg[35]  ( .D(xin[34]), .CLK(clk), .RST(rst), .Q(xreg[35]) );
  DFF \xreg_reg[36]  ( .D(xin[35]), .CLK(clk), .RST(rst), .Q(xreg[36]) );
  DFF \xreg_reg[37]  ( .D(xin[36]), .CLK(clk), .RST(rst), .Q(xreg[37]) );
  DFF \xreg_reg[38]  ( .D(xin[37]), .CLK(clk), .RST(rst), .Q(xreg[38]) );
  DFF \xreg_reg[39]  ( .D(xin[38]), .CLK(clk), .RST(rst), .Q(xreg[39]) );
  DFF \xreg_reg[40]  ( .D(xin[39]), .CLK(clk), .RST(rst), .Q(xreg[40]) );
  DFF \xreg_reg[41]  ( .D(xin[40]), .CLK(clk), .RST(rst), .Q(xreg[41]) );
  DFF \xreg_reg[42]  ( .D(xin[41]), .CLK(clk), .RST(rst), .Q(xreg[42]) );
  DFF \xreg_reg[43]  ( .D(xin[42]), .CLK(clk), .RST(rst), .Q(xreg[43]) );
  DFF \xreg_reg[44]  ( .D(xin[43]), .CLK(clk), .RST(rst), .Q(xreg[44]) );
  DFF \xreg_reg[45]  ( .D(xin[44]), .CLK(clk), .RST(rst), .Q(xreg[45]) );
  DFF \xreg_reg[46]  ( .D(xin[45]), .CLK(clk), .RST(rst), .Q(xreg[46]) );
  DFF \xreg_reg[47]  ( .D(xin[46]), .CLK(clk), .RST(rst), .Q(xreg[47]) );
  DFF \xreg_reg[48]  ( .D(xin[47]), .CLK(clk), .RST(rst), .Q(xreg[48]) );
  DFF \xreg_reg[49]  ( .D(xin[48]), .CLK(clk), .RST(rst), .Q(xreg[49]) );
  DFF \xreg_reg[50]  ( .D(xin[49]), .CLK(clk), .RST(rst), .Q(xreg[50]) );
  DFF \xreg_reg[51]  ( .D(xin[50]), .CLK(clk), .RST(rst), .Q(xreg[51]) );
  DFF \xreg_reg[52]  ( .D(xin[51]), .CLK(clk), .RST(rst), .Q(xreg[52]) );
  DFF \xreg_reg[53]  ( .D(xin[52]), .CLK(clk), .RST(rst), .Q(xreg[53]) );
  DFF \xreg_reg[54]  ( .D(xin[53]), .CLK(clk), .RST(rst), .Q(xreg[54]) );
  DFF \xreg_reg[55]  ( .D(xin[54]), .CLK(clk), .RST(rst), .Q(xreg[55]) );
  DFF \xreg_reg[56]  ( .D(xin[55]), .CLK(clk), .RST(rst), .Q(xreg[56]) );
  DFF \xreg_reg[57]  ( .D(xin[56]), .CLK(clk), .RST(rst), .Q(xreg[57]) );
  DFF \xreg_reg[58]  ( .D(xin[57]), .CLK(clk), .RST(rst), .Q(xreg[58]) );
  DFF \xreg_reg[59]  ( .D(xin[58]), .CLK(clk), .RST(rst), .Q(xreg[59]) );
  DFF \xreg_reg[60]  ( .D(xin[59]), .CLK(clk), .RST(rst), .Q(xreg[60]) );
  DFF \xreg_reg[61]  ( .D(xin[60]), .CLK(clk), .RST(rst), .Q(xreg[61]) );
  DFF \xreg_reg[62]  ( .D(xin[61]), .CLK(clk), .RST(rst), .Q(xreg[62]) );
  DFF \xreg_reg[63]  ( .D(xin[62]), .CLK(clk), .RST(rst), .Q(xreg[63]) );
  DFF \xreg_reg[64]  ( .D(xin[63]), .CLK(clk), .RST(rst), .Q(xreg[64]) );
  DFF \xreg_reg[65]  ( .D(xin[64]), .CLK(clk), .RST(rst), .Q(xreg[65]) );
  DFF \xreg_reg[66]  ( .D(xin[65]), .CLK(clk), .RST(rst), .Q(xreg[66]) );
  DFF \xreg_reg[67]  ( .D(xin[66]), .CLK(clk), .RST(rst), .Q(xreg[67]) );
  DFF \xreg_reg[68]  ( .D(xin[67]), .CLK(clk), .RST(rst), .Q(xreg[68]) );
  DFF \xreg_reg[69]  ( .D(xin[68]), .CLK(clk), .RST(rst), .Q(xreg[69]) );
  DFF \xreg_reg[70]  ( .D(xin[69]), .CLK(clk), .RST(rst), .Q(xreg[70]) );
  DFF \xreg_reg[71]  ( .D(xin[70]), .CLK(clk), .RST(rst), .Q(xreg[71]) );
  DFF \xreg_reg[72]  ( .D(xin[71]), .CLK(clk), .RST(rst), .Q(xreg[72]) );
  DFF \xreg_reg[73]  ( .D(xin[72]), .CLK(clk), .RST(rst), .Q(xreg[73]) );
  DFF \xreg_reg[74]  ( .D(xin[73]), .CLK(clk), .RST(rst), .Q(xreg[74]) );
  DFF \xreg_reg[75]  ( .D(xin[74]), .CLK(clk), .RST(rst), .Q(xreg[75]) );
  DFF \xreg_reg[76]  ( .D(xin[75]), .CLK(clk), .RST(rst), .Q(xreg[76]) );
  DFF \xreg_reg[77]  ( .D(xin[76]), .CLK(clk), .RST(rst), .Q(xreg[77]) );
  DFF \xreg_reg[78]  ( .D(xin[77]), .CLK(clk), .RST(rst), .Q(xreg[78]) );
  DFF \xreg_reg[79]  ( .D(xin[78]), .CLK(clk), .RST(rst), .Q(xreg[79]) );
  DFF \xreg_reg[80]  ( .D(xin[79]), .CLK(clk), .RST(rst), .Q(xreg[80]) );
  DFF \xreg_reg[81]  ( .D(xin[80]), .CLK(clk), .RST(rst), .Q(xreg[81]) );
  DFF \xreg_reg[82]  ( .D(xin[81]), .CLK(clk), .RST(rst), .Q(xreg[82]) );
  DFF \xreg_reg[83]  ( .D(xin[82]), .CLK(clk), .RST(rst), .Q(xreg[83]) );
  DFF \xreg_reg[84]  ( .D(xin[83]), .CLK(clk), .RST(rst), .Q(xreg[84]) );
  DFF \xreg_reg[85]  ( .D(xin[84]), .CLK(clk), .RST(rst), .Q(xreg[85]) );
  DFF \xreg_reg[86]  ( .D(xin[85]), .CLK(clk), .RST(rst), .Q(xreg[86]) );
  DFF \xreg_reg[87]  ( .D(xin[86]), .CLK(clk), .RST(rst), .Q(xreg[87]) );
  DFF \xreg_reg[88]  ( .D(xin[87]), .CLK(clk), .RST(rst), .Q(xreg[88]) );
  DFF \xreg_reg[89]  ( .D(xin[88]), .CLK(clk), .RST(rst), .Q(xreg[89]) );
  DFF \xreg_reg[90]  ( .D(xin[89]), .CLK(clk), .RST(rst), .Q(xreg[90]) );
  DFF \xreg_reg[91]  ( .D(xin[90]), .CLK(clk), .RST(rst), .Q(xreg[91]) );
  DFF \xreg_reg[92]  ( .D(xin[91]), .CLK(clk), .RST(rst), .Q(xreg[92]) );
  DFF \xreg_reg[93]  ( .D(xin[92]), .CLK(clk), .RST(rst), .Q(xreg[93]) );
  DFF \xreg_reg[94]  ( .D(xin[93]), .CLK(clk), .RST(rst), .Q(xreg[94]) );
  DFF \xreg_reg[95]  ( .D(xin[94]), .CLK(clk), .RST(rst), .Q(xreg[95]) );
  DFF \xreg_reg[96]  ( .D(xin[95]), .CLK(clk), .RST(rst), .Q(xreg[96]) );
  DFF \xreg_reg[97]  ( .D(xin[96]), .CLK(clk), .RST(rst), .Q(xreg[97]) );
  DFF \xreg_reg[98]  ( .D(xin[97]), .CLK(clk), .RST(rst), .Q(xreg[98]) );
  DFF \xreg_reg[99]  ( .D(xin[98]), .CLK(clk), .RST(rst), .Q(xreg[99]) );
  DFF \xreg_reg[100]  ( .D(xin[99]), .CLK(clk), .RST(rst), .Q(xreg[100]) );
  DFF \xreg_reg[101]  ( .D(xin[100]), .CLK(clk), .RST(rst), .Q(xreg[101]) );
  DFF \xreg_reg[102]  ( .D(xin[101]), .CLK(clk), .RST(rst), .Q(xreg[102]) );
  DFF \xreg_reg[103]  ( .D(xin[102]), .CLK(clk), .RST(rst), .Q(xreg[103]) );
  DFF \xreg_reg[104]  ( .D(xin[103]), .CLK(clk), .RST(rst), .Q(xreg[104]) );
  DFF \xreg_reg[105]  ( .D(xin[104]), .CLK(clk), .RST(rst), .Q(xreg[105]) );
  DFF \xreg_reg[106]  ( .D(xin[105]), .CLK(clk), .RST(rst), .Q(xreg[106]) );
  DFF \xreg_reg[107]  ( .D(xin[106]), .CLK(clk), .RST(rst), .Q(xreg[107]) );
  DFF \xreg_reg[108]  ( .D(xin[107]), .CLK(clk), .RST(rst), .Q(xreg[108]) );
  DFF \xreg_reg[109]  ( .D(xin[108]), .CLK(clk), .RST(rst), .Q(xreg[109]) );
  DFF \xreg_reg[110]  ( .D(xin[109]), .CLK(clk), .RST(rst), .Q(xreg[110]) );
  DFF \xreg_reg[111]  ( .D(xin[110]), .CLK(clk), .RST(rst), .Q(xreg[111]) );
  DFF \xreg_reg[112]  ( .D(xin[111]), .CLK(clk), .RST(rst), .Q(xreg[112]) );
  DFF \xreg_reg[113]  ( .D(xin[112]), .CLK(clk), .RST(rst), .Q(xreg[113]) );
  DFF \xreg_reg[114]  ( .D(xin[113]), .CLK(clk), .RST(rst), .Q(xreg[114]) );
  DFF \xreg_reg[115]  ( .D(xin[114]), .CLK(clk), .RST(rst), .Q(xreg[115]) );
  DFF \xreg_reg[116]  ( .D(xin[115]), .CLK(clk), .RST(rst), .Q(xreg[116]) );
  DFF \xreg_reg[117]  ( .D(xin[116]), .CLK(clk), .RST(rst), .Q(xreg[117]) );
  DFF \xreg_reg[118]  ( .D(xin[117]), .CLK(clk), .RST(rst), .Q(xreg[118]) );
  DFF \xreg_reg[119]  ( .D(xin[118]), .CLK(clk), .RST(rst), .Q(xreg[119]) );
  DFF \xreg_reg[120]  ( .D(xin[119]), .CLK(clk), .RST(rst), .Q(xreg[120]) );
  DFF \xreg_reg[121]  ( .D(xin[120]), .CLK(clk), .RST(rst), .Q(xreg[121]) );
  DFF \xreg_reg[122]  ( .D(xin[121]), .CLK(clk), .RST(rst), .Q(xreg[122]) );
  DFF \xreg_reg[123]  ( .D(xin[122]), .CLK(clk), .RST(rst), .Q(xreg[123]) );
  DFF \xreg_reg[124]  ( .D(xin[123]), .CLK(clk), .RST(rst), .Q(xreg[124]) );
  DFF \xreg_reg[125]  ( .D(xin[124]), .CLK(clk), .RST(rst), .Q(xreg[125]) );
  DFF \xreg_reg[126]  ( .D(xin[125]), .CLK(clk), .RST(rst), .Q(xreg[126]) );
  DFF \xreg_reg[127]  ( .D(xin[126]), .CLK(clk), .RST(rst), .Q(xreg[127]) );
  DFF \xreg_reg[128]  ( .D(xin[127]), .CLK(clk), .RST(rst), .Q(xreg[128]) );
  DFF \xreg_reg[129]  ( .D(xin[128]), .CLK(clk), .RST(rst), .Q(xreg[129]) );
  DFF \xreg_reg[130]  ( .D(xin[129]), .CLK(clk), .RST(rst), .Q(xreg[130]) );
  DFF \xreg_reg[131]  ( .D(xin[130]), .CLK(clk), .RST(rst), .Q(xreg[131]) );
  DFF \xreg_reg[132]  ( .D(xin[131]), .CLK(clk), .RST(rst), .Q(xreg[132]) );
  DFF \xreg_reg[133]  ( .D(xin[132]), .CLK(clk), .RST(rst), .Q(xreg[133]) );
  DFF \xreg_reg[134]  ( .D(xin[133]), .CLK(clk), .RST(rst), .Q(xreg[134]) );
  DFF \xreg_reg[135]  ( .D(xin[134]), .CLK(clk), .RST(rst), .Q(xreg[135]) );
  DFF \xreg_reg[136]  ( .D(xin[135]), .CLK(clk), .RST(rst), .Q(xreg[136]) );
  DFF \xreg_reg[137]  ( .D(xin[136]), .CLK(clk), .RST(rst), .Q(xreg[137]) );
  DFF \xreg_reg[138]  ( .D(xin[137]), .CLK(clk), .RST(rst), .Q(xreg[138]) );
  DFF \xreg_reg[139]  ( .D(xin[138]), .CLK(clk), .RST(rst), .Q(xreg[139]) );
  DFF \xreg_reg[140]  ( .D(xin[139]), .CLK(clk), .RST(rst), .Q(xreg[140]) );
  DFF \xreg_reg[141]  ( .D(xin[140]), .CLK(clk), .RST(rst), .Q(xreg[141]) );
  DFF \xreg_reg[142]  ( .D(xin[141]), .CLK(clk), .RST(rst), .Q(xreg[142]) );
  DFF \xreg_reg[143]  ( .D(xin[142]), .CLK(clk), .RST(rst), .Q(xreg[143]) );
  DFF \xreg_reg[144]  ( .D(xin[143]), .CLK(clk), .RST(rst), .Q(xreg[144]) );
  DFF \xreg_reg[145]  ( .D(xin[144]), .CLK(clk), .RST(rst), .Q(xreg[145]) );
  DFF \xreg_reg[146]  ( .D(xin[145]), .CLK(clk), .RST(rst), .Q(xreg[146]) );
  DFF \xreg_reg[147]  ( .D(xin[146]), .CLK(clk), .RST(rst), .Q(xreg[147]) );
  DFF \xreg_reg[148]  ( .D(xin[147]), .CLK(clk), .RST(rst), .Q(xreg[148]) );
  DFF \xreg_reg[149]  ( .D(xin[148]), .CLK(clk), .RST(rst), .Q(xreg[149]) );
  DFF \xreg_reg[150]  ( .D(xin[149]), .CLK(clk), .RST(rst), .Q(xreg[150]) );
  DFF \xreg_reg[151]  ( .D(xin[150]), .CLK(clk), .RST(rst), .Q(xreg[151]) );
  DFF \xreg_reg[152]  ( .D(xin[151]), .CLK(clk), .RST(rst), .Q(xreg[152]) );
  DFF \xreg_reg[153]  ( .D(xin[152]), .CLK(clk), .RST(rst), .Q(xreg[153]) );
  DFF \xreg_reg[154]  ( .D(xin[153]), .CLK(clk), .RST(rst), .Q(xreg[154]) );
  DFF \xreg_reg[155]  ( .D(xin[154]), .CLK(clk), .RST(rst), .Q(xreg[155]) );
  DFF \xreg_reg[156]  ( .D(xin[155]), .CLK(clk), .RST(rst), .Q(xreg[156]) );
  DFF \xreg_reg[157]  ( .D(xin[156]), .CLK(clk), .RST(rst), .Q(xreg[157]) );
  DFF \xreg_reg[158]  ( .D(xin[157]), .CLK(clk), .RST(rst), .Q(xreg[158]) );
  DFF \xreg_reg[159]  ( .D(xin[158]), .CLK(clk), .RST(rst), .Q(xreg[159]) );
  DFF \xreg_reg[160]  ( .D(xin[159]), .CLK(clk), .RST(rst), .Q(xreg[160]) );
  DFF \xreg_reg[161]  ( .D(xin[160]), .CLK(clk), .RST(rst), .Q(xreg[161]) );
  DFF \xreg_reg[162]  ( .D(xin[161]), .CLK(clk), .RST(rst), .Q(xreg[162]) );
  DFF \xreg_reg[163]  ( .D(xin[162]), .CLK(clk), .RST(rst), .Q(xreg[163]) );
  DFF \xreg_reg[164]  ( .D(xin[163]), .CLK(clk), .RST(rst), .Q(xreg[164]) );
  DFF \xreg_reg[165]  ( .D(xin[164]), .CLK(clk), .RST(rst), .Q(xreg[165]) );
  DFF \xreg_reg[166]  ( .D(xin[165]), .CLK(clk), .RST(rst), .Q(xreg[166]) );
  DFF \xreg_reg[167]  ( .D(xin[166]), .CLK(clk), .RST(rst), .Q(xreg[167]) );
  DFF \xreg_reg[168]  ( .D(xin[167]), .CLK(clk), .RST(rst), .Q(xreg[168]) );
  DFF \xreg_reg[169]  ( .D(xin[168]), .CLK(clk), .RST(rst), .Q(xreg[169]) );
  DFF \xreg_reg[170]  ( .D(xin[169]), .CLK(clk), .RST(rst), .Q(xreg[170]) );
  DFF \xreg_reg[171]  ( .D(xin[170]), .CLK(clk), .RST(rst), .Q(xreg[171]) );
  DFF \xreg_reg[172]  ( .D(xin[171]), .CLK(clk), .RST(rst), .Q(xreg[172]) );
  DFF \xreg_reg[173]  ( .D(xin[172]), .CLK(clk), .RST(rst), .Q(xreg[173]) );
  DFF \xreg_reg[174]  ( .D(xin[173]), .CLK(clk), .RST(rst), .Q(xreg[174]) );
  DFF \xreg_reg[175]  ( .D(xin[174]), .CLK(clk), .RST(rst), .Q(xreg[175]) );
  DFF \xreg_reg[176]  ( .D(xin[175]), .CLK(clk), .RST(rst), .Q(xreg[176]) );
  DFF \xreg_reg[177]  ( .D(xin[176]), .CLK(clk), .RST(rst), .Q(xreg[177]) );
  DFF \xreg_reg[178]  ( .D(xin[177]), .CLK(clk), .RST(rst), .Q(xreg[178]) );
  DFF \xreg_reg[179]  ( .D(xin[178]), .CLK(clk), .RST(rst), .Q(xreg[179]) );
  DFF \xreg_reg[180]  ( .D(xin[179]), .CLK(clk), .RST(rst), .Q(xreg[180]) );
  DFF \xreg_reg[181]  ( .D(xin[180]), .CLK(clk), .RST(rst), .Q(xreg[181]) );
  DFF \xreg_reg[182]  ( .D(xin[181]), .CLK(clk), .RST(rst), .Q(xreg[182]) );
  DFF \xreg_reg[183]  ( .D(xin[182]), .CLK(clk), .RST(rst), .Q(xreg[183]) );
  DFF \xreg_reg[184]  ( .D(xin[183]), .CLK(clk), .RST(rst), .Q(xreg[184]) );
  DFF \xreg_reg[185]  ( .D(xin[184]), .CLK(clk), .RST(rst), .Q(xreg[185]) );
  DFF \xreg_reg[186]  ( .D(xin[185]), .CLK(clk), .RST(rst), .Q(xreg[186]) );
  DFF \xreg_reg[187]  ( .D(xin[186]), .CLK(clk), .RST(rst), .Q(xreg[187]) );
  DFF \xreg_reg[188]  ( .D(xin[187]), .CLK(clk), .RST(rst), .Q(xreg[188]) );
  DFF \xreg_reg[189]  ( .D(xin[188]), .CLK(clk), .RST(rst), .Q(xreg[189]) );
  DFF \xreg_reg[190]  ( .D(xin[189]), .CLK(clk), .RST(rst), .Q(xreg[190]) );
  DFF \xreg_reg[191]  ( .D(xin[190]), .CLK(clk), .RST(rst), .Q(xreg[191]) );
  DFF \xreg_reg[192]  ( .D(xin[191]), .CLK(clk), .RST(rst), .Q(xreg[192]) );
  DFF \xreg_reg[193]  ( .D(xin[192]), .CLK(clk), .RST(rst), .Q(xreg[193]) );
  DFF \xreg_reg[194]  ( .D(xin[193]), .CLK(clk), .RST(rst), .Q(xreg[194]) );
  DFF \xreg_reg[195]  ( .D(xin[194]), .CLK(clk), .RST(rst), .Q(xreg[195]) );
  DFF \xreg_reg[196]  ( .D(xin[195]), .CLK(clk), .RST(rst), .Q(xreg[196]) );
  DFF \xreg_reg[197]  ( .D(xin[196]), .CLK(clk), .RST(rst), .Q(xreg[197]) );
  DFF \xreg_reg[198]  ( .D(xin[197]), .CLK(clk), .RST(rst), .Q(xreg[198]) );
  DFF \xreg_reg[199]  ( .D(xin[198]), .CLK(clk), .RST(rst), .Q(xreg[199]) );
  DFF \xreg_reg[200]  ( .D(xin[199]), .CLK(clk), .RST(rst), .Q(xreg[200]) );
  DFF \xreg_reg[201]  ( .D(xin[200]), .CLK(clk), .RST(rst), .Q(xreg[201]) );
  DFF \xreg_reg[202]  ( .D(xin[201]), .CLK(clk), .RST(rst), .Q(xreg[202]) );
  DFF \xreg_reg[203]  ( .D(xin[202]), .CLK(clk), .RST(rst), .Q(xreg[203]) );
  DFF \xreg_reg[204]  ( .D(xin[203]), .CLK(clk), .RST(rst), .Q(xreg[204]) );
  DFF \xreg_reg[205]  ( .D(xin[204]), .CLK(clk), .RST(rst), .Q(xreg[205]) );
  DFF \xreg_reg[206]  ( .D(xin[205]), .CLK(clk), .RST(rst), .Q(xreg[206]) );
  DFF \xreg_reg[207]  ( .D(xin[206]), .CLK(clk), .RST(rst), .Q(xreg[207]) );
  DFF \xreg_reg[208]  ( .D(xin[207]), .CLK(clk), .RST(rst), .Q(xreg[208]) );
  DFF \xreg_reg[209]  ( .D(xin[208]), .CLK(clk), .RST(rst), .Q(xreg[209]) );
  DFF \xreg_reg[210]  ( .D(xin[209]), .CLK(clk), .RST(rst), .Q(xreg[210]) );
  DFF \xreg_reg[211]  ( .D(xin[210]), .CLK(clk), .RST(rst), .Q(xreg[211]) );
  DFF \xreg_reg[212]  ( .D(xin[211]), .CLK(clk), .RST(rst), .Q(xreg[212]) );
  DFF \xreg_reg[213]  ( .D(xin[212]), .CLK(clk), .RST(rst), .Q(xreg[213]) );
  DFF \xreg_reg[214]  ( .D(xin[213]), .CLK(clk), .RST(rst), .Q(xreg[214]) );
  DFF \xreg_reg[215]  ( .D(xin[214]), .CLK(clk), .RST(rst), .Q(xreg[215]) );
  DFF \xreg_reg[216]  ( .D(xin[215]), .CLK(clk), .RST(rst), .Q(xreg[216]) );
  DFF \xreg_reg[217]  ( .D(xin[216]), .CLK(clk), .RST(rst), .Q(xreg[217]) );
  DFF \xreg_reg[218]  ( .D(xin[217]), .CLK(clk), .RST(rst), .Q(xreg[218]) );
  DFF \xreg_reg[219]  ( .D(xin[218]), .CLK(clk), .RST(rst), .Q(xreg[219]) );
  DFF \xreg_reg[220]  ( .D(xin[219]), .CLK(clk), .RST(rst), .Q(xreg[220]) );
  DFF \xreg_reg[221]  ( .D(xin[220]), .CLK(clk), .RST(rst), .Q(xreg[221]) );
  DFF \xreg_reg[222]  ( .D(xin[221]), .CLK(clk), .RST(rst), .Q(xreg[222]) );
  DFF \xreg_reg[223]  ( .D(xin[222]), .CLK(clk), .RST(rst), .Q(xreg[223]) );
  DFF \xreg_reg[224]  ( .D(xin[223]), .CLK(clk), .RST(rst), .Q(xreg[224]) );
  DFF \xreg_reg[225]  ( .D(xin[224]), .CLK(clk), .RST(rst), .Q(xreg[225]) );
  DFF \xreg_reg[226]  ( .D(xin[225]), .CLK(clk), .RST(rst), .Q(xreg[226]) );
  DFF \xreg_reg[227]  ( .D(xin[226]), .CLK(clk), .RST(rst), .Q(xreg[227]) );
  DFF \xreg_reg[228]  ( .D(xin[227]), .CLK(clk), .RST(rst), .Q(xreg[228]) );
  DFF \xreg_reg[229]  ( .D(xin[228]), .CLK(clk), .RST(rst), .Q(xreg[229]) );
  DFF \xreg_reg[230]  ( .D(xin[229]), .CLK(clk), .RST(rst), .Q(xreg[230]) );
  DFF \xreg_reg[231]  ( .D(xin[230]), .CLK(clk), .RST(rst), .Q(xreg[231]) );
  DFF \xreg_reg[232]  ( .D(xin[231]), .CLK(clk), .RST(rst), .Q(xreg[232]) );
  DFF \xreg_reg[233]  ( .D(xin[232]), .CLK(clk), .RST(rst), .Q(xreg[233]) );
  DFF \xreg_reg[234]  ( .D(xin[233]), .CLK(clk), .RST(rst), .Q(xreg[234]) );
  DFF \xreg_reg[235]  ( .D(xin[234]), .CLK(clk), .RST(rst), .Q(xreg[235]) );
  DFF \xreg_reg[236]  ( .D(xin[235]), .CLK(clk), .RST(rst), .Q(xreg[236]) );
  DFF \xreg_reg[237]  ( .D(xin[236]), .CLK(clk), .RST(rst), .Q(xreg[237]) );
  DFF \xreg_reg[238]  ( .D(xin[237]), .CLK(clk), .RST(rst), .Q(xreg[238]) );
  DFF \xreg_reg[239]  ( .D(xin[238]), .CLK(clk), .RST(rst), .Q(xreg[239]) );
  DFF \xreg_reg[240]  ( .D(xin[239]), .CLK(clk), .RST(rst), .Q(xreg[240]) );
  DFF \xreg_reg[241]  ( .D(xin[240]), .CLK(clk), .RST(rst), .Q(xreg[241]) );
  DFF \xreg_reg[242]  ( .D(xin[241]), .CLK(clk), .RST(rst), .Q(xreg[242]) );
  DFF \xreg_reg[243]  ( .D(xin[242]), .CLK(clk), .RST(rst), .Q(xreg[243]) );
  DFF \xreg_reg[244]  ( .D(xin[243]), .CLK(clk), .RST(rst), .Q(xreg[244]) );
  DFF \xreg_reg[245]  ( .D(xin[244]), .CLK(clk), .RST(rst), .Q(xreg[245]) );
  DFF \xreg_reg[246]  ( .D(xin[245]), .CLK(clk), .RST(rst), .Q(xreg[246]) );
  DFF \xreg_reg[247]  ( .D(xin[246]), .CLK(clk), .RST(rst), .Q(xreg[247]) );
  DFF \xreg_reg[248]  ( .D(xin[247]), .CLK(clk), .RST(rst), .Q(xreg[248]) );
  DFF \xreg_reg[249]  ( .D(xin[248]), .CLK(clk), .RST(rst), .Q(xreg[249]) );
  DFF \xreg_reg[250]  ( .D(xin[249]), .CLK(clk), .RST(rst), .Q(xreg[250]) );
  DFF \xreg_reg[251]  ( .D(xin[250]), .CLK(clk), .RST(rst), .Q(xreg[251]) );
  DFF \xreg_reg[252]  ( .D(xin[251]), .CLK(clk), .RST(rst), .Q(xreg[252]) );
  DFF \xreg_reg[253]  ( .D(xin[252]), .CLK(clk), .RST(rst), .Q(xreg[253]) );
  DFF \xreg_reg[254]  ( .D(xin[253]), .CLK(clk), .RST(rst), .Q(xreg[254]) );
  DFF \xreg_reg[255]  ( .D(xin[254]), .CLK(clk), .RST(rst), .Q(xreg[255]) );
  DFF \xreg_reg[256]  ( .D(xin[255]), .CLK(clk), .RST(rst), .Q(xreg[256]) );
  DFF \xreg_reg[257]  ( .D(xin[256]), .CLK(clk), .RST(rst), .Q(xreg[257]) );
  DFF \xreg_reg[258]  ( .D(xin[257]), .CLK(clk), .RST(rst), .Q(xreg[258]) );
  DFF \xreg_reg[259]  ( .D(xin[258]), .CLK(clk), .RST(rst), .Q(xreg[259]) );
  DFF \xreg_reg[260]  ( .D(xin[259]), .CLK(clk), .RST(rst), .Q(xreg[260]) );
  DFF \xreg_reg[261]  ( .D(xin[260]), .CLK(clk), .RST(rst), .Q(xreg[261]) );
  DFF \xreg_reg[262]  ( .D(xin[261]), .CLK(clk), .RST(rst), .Q(xreg[262]) );
  DFF \xreg_reg[263]  ( .D(xin[262]), .CLK(clk), .RST(rst), .Q(xreg[263]) );
  DFF \xreg_reg[264]  ( .D(xin[263]), .CLK(clk), .RST(rst), .Q(xreg[264]) );
  DFF \xreg_reg[265]  ( .D(xin[264]), .CLK(clk), .RST(rst), .Q(xreg[265]) );
  DFF \xreg_reg[266]  ( .D(xin[265]), .CLK(clk), .RST(rst), .Q(xreg[266]) );
  DFF \xreg_reg[267]  ( .D(xin[266]), .CLK(clk), .RST(rst), .Q(xreg[267]) );
  DFF \xreg_reg[268]  ( .D(xin[267]), .CLK(clk), .RST(rst), .Q(xreg[268]) );
  DFF \xreg_reg[269]  ( .D(xin[268]), .CLK(clk), .RST(rst), .Q(xreg[269]) );
  DFF \xreg_reg[270]  ( .D(xin[269]), .CLK(clk), .RST(rst), .Q(xreg[270]) );
  DFF \xreg_reg[271]  ( .D(xin[270]), .CLK(clk), .RST(rst), .Q(xreg[271]) );
  DFF \xreg_reg[272]  ( .D(xin[271]), .CLK(clk), .RST(rst), .Q(xreg[272]) );
  DFF \xreg_reg[273]  ( .D(xin[272]), .CLK(clk), .RST(rst), .Q(xreg[273]) );
  DFF \xreg_reg[274]  ( .D(xin[273]), .CLK(clk), .RST(rst), .Q(xreg[274]) );
  DFF \xreg_reg[275]  ( .D(xin[274]), .CLK(clk), .RST(rst), .Q(xreg[275]) );
  DFF \xreg_reg[276]  ( .D(xin[275]), .CLK(clk), .RST(rst), .Q(xreg[276]) );
  DFF \xreg_reg[277]  ( .D(xin[276]), .CLK(clk), .RST(rst), .Q(xreg[277]) );
  DFF \xreg_reg[278]  ( .D(xin[277]), .CLK(clk), .RST(rst), .Q(xreg[278]) );
  DFF \xreg_reg[279]  ( .D(xin[278]), .CLK(clk), .RST(rst), .Q(xreg[279]) );
  DFF \xreg_reg[280]  ( .D(xin[279]), .CLK(clk), .RST(rst), .Q(xreg[280]) );
  DFF \xreg_reg[281]  ( .D(xin[280]), .CLK(clk), .RST(rst), .Q(xreg[281]) );
  DFF \xreg_reg[282]  ( .D(xin[281]), .CLK(clk), .RST(rst), .Q(xreg[282]) );
  DFF \xreg_reg[283]  ( .D(xin[282]), .CLK(clk), .RST(rst), .Q(xreg[283]) );
  DFF \xreg_reg[284]  ( .D(xin[283]), .CLK(clk), .RST(rst), .Q(xreg[284]) );
  DFF \xreg_reg[285]  ( .D(xin[284]), .CLK(clk), .RST(rst), .Q(xreg[285]) );
  DFF \xreg_reg[286]  ( .D(xin[285]), .CLK(clk), .RST(rst), .Q(xreg[286]) );
  DFF \xreg_reg[287]  ( .D(xin[286]), .CLK(clk), .RST(rst), .Q(xreg[287]) );
  DFF \xreg_reg[288]  ( .D(xin[287]), .CLK(clk), .RST(rst), .Q(xreg[288]) );
  DFF \xreg_reg[289]  ( .D(xin[288]), .CLK(clk), .RST(rst), .Q(xreg[289]) );
  DFF \xreg_reg[290]  ( .D(xin[289]), .CLK(clk), .RST(rst), .Q(xreg[290]) );
  DFF \xreg_reg[291]  ( .D(xin[290]), .CLK(clk), .RST(rst), .Q(xreg[291]) );
  DFF \xreg_reg[292]  ( .D(xin[291]), .CLK(clk), .RST(rst), .Q(xreg[292]) );
  DFF \xreg_reg[293]  ( .D(xin[292]), .CLK(clk), .RST(rst), .Q(xreg[293]) );
  DFF \xreg_reg[294]  ( .D(xin[293]), .CLK(clk), .RST(rst), .Q(xreg[294]) );
  DFF \xreg_reg[295]  ( .D(xin[294]), .CLK(clk), .RST(rst), .Q(xreg[295]) );
  DFF \xreg_reg[296]  ( .D(xin[295]), .CLK(clk), .RST(rst), .Q(xreg[296]) );
  DFF \xreg_reg[297]  ( .D(xin[296]), .CLK(clk), .RST(rst), .Q(xreg[297]) );
  DFF \xreg_reg[298]  ( .D(xin[297]), .CLK(clk), .RST(rst), .Q(xreg[298]) );
  DFF \xreg_reg[299]  ( .D(xin[298]), .CLK(clk), .RST(rst), .Q(xreg[299]) );
  DFF \xreg_reg[300]  ( .D(xin[299]), .CLK(clk), .RST(rst), .Q(xreg[300]) );
  DFF \xreg_reg[301]  ( .D(xin[300]), .CLK(clk), .RST(rst), .Q(xreg[301]) );
  DFF \xreg_reg[302]  ( .D(xin[301]), .CLK(clk), .RST(rst), .Q(xreg[302]) );
  DFF \xreg_reg[303]  ( .D(xin[302]), .CLK(clk), .RST(rst), .Q(xreg[303]) );
  DFF \xreg_reg[304]  ( .D(xin[303]), .CLK(clk), .RST(rst), .Q(xreg[304]) );
  DFF \xreg_reg[305]  ( .D(xin[304]), .CLK(clk), .RST(rst), .Q(xreg[305]) );
  DFF \xreg_reg[306]  ( .D(xin[305]), .CLK(clk), .RST(rst), .Q(xreg[306]) );
  DFF \xreg_reg[307]  ( .D(xin[306]), .CLK(clk), .RST(rst), .Q(xreg[307]) );
  DFF \xreg_reg[308]  ( .D(xin[307]), .CLK(clk), .RST(rst), .Q(xreg[308]) );
  DFF \xreg_reg[309]  ( .D(xin[308]), .CLK(clk), .RST(rst), .Q(xreg[309]) );
  DFF \xreg_reg[310]  ( .D(xin[309]), .CLK(clk), .RST(rst), .Q(xreg[310]) );
  DFF \xreg_reg[311]  ( .D(xin[310]), .CLK(clk), .RST(rst), .Q(xreg[311]) );
  DFF \xreg_reg[312]  ( .D(xin[311]), .CLK(clk), .RST(rst), .Q(xreg[312]) );
  DFF \xreg_reg[313]  ( .D(xin[312]), .CLK(clk), .RST(rst), .Q(xreg[313]) );
  DFF \xreg_reg[314]  ( .D(xin[313]), .CLK(clk), .RST(rst), .Q(xreg[314]) );
  DFF \xreg_reg[315]  ( .D(xin[314]), .CLK(clk), .RST(rst), .Q(xreg[315]) );
  DFF \xreg_reg[316]  ( .D(xin[315]), .CLK(clk), .RST(rst), .Q(xreg[316]) );
  DFF \xreg_reg[317]  ( .D(xin[316]), .CLK(clk), .RST(rst), .Q(xreg[317]) );
  DFF \xreg_reg[318]  ( .D(xin[317]), .CLK(clk), .RST(rst), .Q(xreg[318]) );
  DFF \xreg_reg[319]  ( .D(xin[318]), .CLK(clk), .RST(rst), .Q(xreg[319]) );
  DFF \xreg_reg[320]  ( .D(xin[319]), .CLK(clk), .RST(rst), .Q(xreg[320]) );
  DFF \xreg_reg[321]  ( .D(xin[320]), .CLK(clk), .RST(rst), .Q(xreg[321]) );
  DFF \xreg_reg[322]  ( .D(xin[321]), .CLK(clk), .RST(rst), .Q(xreg[322]) );
  DFF \xreg_reg[323]  ( .D(xin[322]), .CLK(clk), .RST(rst), .Q(xreg[323]) );
  DFF \xreg_reg[324]  ( .D(xin[323]), .CLK(clk), .RST(rst), .Q(xreg[324]) );
  DFF \xreg_reg[325]  ( .D(xin[324]), .CLK(clk), .RST(rst), .Q(xreg[325]) );
  DFF \xreg_reg[326]  ( .D(xin[325]), .CLK(clk), .RST(rst), .Q(xreg[326]) );
  DFF \xreg_reg[327]  ( .D(xin[326]), .CLK(clk), .RST(rst), .Q(xreg[327]) );
  DFF \xreg_reg[328]  ( .D(xin[327]), .CLK(clk), .RST(rst), .Q(xreg[328]) );
  DFF \xreg_reg[329]  ( .D(xin[328]), .CLK(clk), .RST(rst), .Q(xreg[329]) );
  DFF \xreg_reg[330]  ( .D(xin[329]), .CLK(clk), .RST(rst), .Q(xreg[330]) );
  DFF \xreg_reg[331]  ( .D(xin[330]), .CLK(clk), .RST(rst), .Q(xreg[331]) );
  DFF \xreg_reg[332]  ( .D(xin[331]), .CLK(clk), .RST(rst), .Q(xreg[332]) );
  DFF \xreg_reg[333]  ( .D(xin[332]), .CLK(clk), .RST(rst), .Q(xreg[333]) );
  DFF \xreg_reg[334]  ( .D(xin[333]), .CLK(clk), .RST(rst), .Q(xreg[334]) );
  DFF \xreg_reg[335]  ( .D(xin[334]), .CLK(clk), .RST(rst), .Q(xreg[335]) );
  DFF \xreg_reg[336]  ( .D(xin[335]), .CLK(clk), .RST(rst), .Q(xreg[336]) );
  DFF \xreg_reg[337]  ( .D(xin[336]), .CLK(clk), .RST(rst), .Q(xreg[337]) );
  DFF \xreg_reg[338]  ( .D(xin[337]), .CLK(clk), .RST(rst), .Q(xreg[338]) );
  DFF \xreg_reg[339]  ( .D(xin[338]), .CLK(clk), .RST(rst), .Q(xreg[339]) );
  DFF \xreg_reg[340]  ( .D(xin[339]), .CLK(clk), .RST(rst), .Q(xreg[340]) );
  DFF \xreg_reg[341]  ( .D(xin[340]), .CLK(clk), .RST(rst), .Q(xreg[341]) );
  DFF \xreg_reg[342]  ( .D(xin[341]), .CLK(clk), .RST(rst), .Q(xreg[342]) );
  DFF \xreg_reg[343]  ( .D(xin[342]), .CLK(clk), .RST(rst), .Q(xreg[343]) );
  DFF \xreg_reg[344]  ( .D(xin[343]), .CLK(clk), .RST(rst), .Q(xreg[344]) );
  DFF \xreg_reg[345]  ( .D(xin[344]), .CLK(clk), .RST(rst), .Q(xreg[345]) );
  DFF \xreg_reg[346]  ( .D(xin[345]), .CLK(clk), .RST(rst), .Q(xreg[346]) );
  DFF \xreg_reg[347]  ( .D(xin[346]), .CLK(clk), .RST(rst), .Q(xreg[347]) );
  DFF \xreg_reg[348]  ( .D(xin[347]), .CLK(clk), .RST(rst), .Q(xreg[348]) );
  DFF \xreg_reg[349]  ( .D(xin[348]), .CLK(clk), .RST(rst), .Q(xreg[349]) );
  DFF \xreg_reg[350]  ( .D(xin[349]), .CLK(clk), .RST(rst), .Q(xreg[350]) );
  DFF \xreg_reg[351]  ( .D(xin[350]), .CLK(clk), .RST(rst), .Q(xreg[351]) );
  DFF \xreg_reg[352]  ( .D(xin[351]), .CLK(clk), .RST(rst), .Q(xreg[352]) );
  DFF \xreg_reg[353]  ( .D(xin[352]), .CLK(clk), .RST(rst), .Q(xreg[353]) );
  DFF \xreg_reg[354]  ( .D(xin[353]), .CLK(clk), .RST(rst), .Q(xreg[354]) );
  DFF \xreg_reg[355]  ( .D(xin[354]), .CLK(clk), .RST(rst), .Q(xreg[355]) );
  DFF \xreg_reg[356]  ( .D(xin[355]), .CLK(clk), .RST(rst), .Q(xreg[356]) );
  DFF \xreg_reg[357]  ( .D(xin[356]), .CLK(clk), .RST(rst), .Q(xreg[357]) );
  DFF \xreg_reg[358]  ( .D(xin[357]), .CLK(clk), .RST(rst), .Q(xreg[358]) );
  DFF \xreg_reg[359]  ( .D(xin[358]), .CLK(clk), .RST(rst), .Q(xreg[359]) );
  DFF \xreg_reg[360]  ( .D(xin[359]), .CLK(clk), .RST(rst), .Q(xreg[360]) );
  DFF \xreg_reg[361]  ( .D(xin[360]), .CLK(clk), .RST(rst), .Q(xreg[361]) );
  DFF \xreg_reg[362]  ( .D(xin[361]), .CLK(clk), .RST(rst), .Q(xreg[362]) );
  DFF \xreg_reg[363]  ( .D(xin[362]), .CLK(clk), .RST(rst), .Q(xreg[363]) );
  DFF \xreg_reg[364]  ( .D(xin[363]), .CLK(clk), .RST(rst), .Q(xreg[364]) );
  DFF \xreg_reg[365]  ( .D(xin[364]), .CLK(clk), .RST(rst), .Q(xreg[365]) );
  DFF \xreg_reg[366]  ( .D(xin[365]), .CLK(clk), .RST(rst), .Q(xreg[366]) );
  DFF \xreg_reg[367]  ( .D(xin[366]), .CLK(clk), .RST(rst), .Q(xreg[367]) );
  DFF \xreg_reg[368]  ( .D(xin[367]), .CLK(clk), .RST(rst), .Q(xreg[368]) );
  DFF \xreg_reg[369]  ( .D(xin[368]), .CLK(clk), .RST(rst), .Q(xreg[369]) );
  DFF \xreg_reg[370]  ( .D(xin[369]), .CLK(clk), .RST(rst), .Q(xreg[370]) );
  DFF \xreg_reg[371]  ( .D(xin[370]), .CLK(clk), .RST(rst), .Q(xreg[371]) );
  DFF \xreg_reg[372]  ( .D(xin[371]), .CLK(clk), .RST(rst), .Q(xreg[372]) );
  DFF \xreg_reg[373]  ( .D(xin[372]), .CLK(clk), .RST(rst), .Q(xreg[373]) );
  DFF \xreg_reg[374]  ( .D(xin[373]), .CLK(clk), .RST(rst), .Q(xreg[374]) );
  DFF \xreg_reg[375]  ( .D(xin[374]), .CLK(clk), .RST(rst), .Q(xreg[375]) );
  DFF \xreg_reg[376]  ( .D(xin[375]), .CLK(clk), .RST(rst), .Q(xreg[376]) );
  DFF \xreg_reg[377]  ( .D(xin[376]), .CLK(clk), .RST(rst), .Q(xreg[377]) );
  DFF \xreg_reg[378]  ( .D(xin[377]), .CLK(clk), .RST(rst), .Q(xreg[378]) );
  DFF \xreg_reg[379]  ( .D(xin[378]), .CLK(clk), .RST(rst), .Q(xreg[379]) );
  DFF \xreg_reg[380]  ( .D(xin[379]), .CLK(clk), .RST(rst), .Q(xreg[380]) );
  DFF \xreg_reg[381]  ( .D(xin[380]), .CLK(clk), .RST(rst), .Q(xreg[381]) );
  DFF \xreg_reg[382]  ( .D(xin[381]), .CLK(clk), .RST(rst), .Q(xreg[382]) );
  DFF \xreg_reg[383]  ( .D(xin[382]), .CLK(clk), .RST(rst), .Q(xreg[383]) );
  DFF \xreg_reg[384]  ( .D(xin[383]), .CLK(clk), .RST(rst), .Q(xreg[384]) );
  DFF \xreg_reg[385]  ( .D(xin[384]), .CLK(clk), .RST(rst), .Q(xreg[385]) );
  DFF \xreg_reg[386]  ( .D(xin[385]), .CLK(clk), .RST(rst), .Q(xreg[386]) );
  DFF \xreg_reg[387]  ( .D(xin[386]), .CLK(clk), .RST(rst), .Q(xreg[387]) );
  DFF \xreg_reg[388]  ( .D(xin[387]), .CLK(clk), .RST(rst), .Q(xreg[388]) );
  DFF \xreg_reg[389]  ( .D(xin[388]), .CLK(clk), .RST(rst), .Q(xreg[389]) );
  DFF \xreg_reg[390]  ( .D(xin[389]), .CLK(clk), .RST(rst), .Q(xreg[390]) );
  DFF \xreg_reg[391]  ( .D(xin[390]), .CLK(clk), .RST(rst), .Q(xreg[391]) );
  DFF \xreg_reg[392]  ( .D(xin[391]), .CLK(clk), .RST(rst), .Q(xreg[392]) );
  DFF \xreg_reg[393]  ( .D(xin[392]), .CLK(clk), .RST(rst), .Q(xreg[393]) );
  DFF \xreg_reg[394]  ( .D(xin[393]), .CLK(clk), .RST(rst), .Q(xreg[394]) );
  DFF \xreg_reg[395]  ( .D(xin[394]), .CLK(clk), .RST(rst), .Q(xreg[395]) );
  DFF \xreg_reg[396]  ( .D(xin[395]), .CLK(clk), .RST(rst), .Q(xreg[396]) );
  DFF \xreg_reg[397]  ( .D(xin[396]), .CLK(clk), .RST(rst), .Q(xreg[397]) );
  DFF \xreg_reg[398]  ( .D(xin[397]), .CLK(clk), .RST(rst), .Q(xreg[398]) );
  DFF \xreg_reg[399]  ( .D(xin[398]), .CLK(clk), .RST(rst), .Q(xreg[399]) );
  DFF \xreg_reg[400]  ( .D(xin[399]), .CLK(clk), .RST(rst), .Q(xreg[400]) );
  DFF \xreg_reg[401]  ( .D(xin[400]), .CLK(clk), .RST(rst), .Q(xreg[401]) );
  DFF \xreg_reg[402]  ( .D(xin[401]), .CLK(clk), .RST(rst), .Q(xreg[402]) );
  DFF \xreg_reg[403]  ( .D(xin[402]), .CLK(clk), .RST(rst), .Q(xreg[403]) );
  DFF \xreg_reg[404]  ( .D(xin[403]), .CLK(clk), .RST(rst), .Q(xreg[404]) );
  DFF \xreg_reg[405]  ( .D(xin[404]), .CLK(clk), .RST(rst), .Q(xreg[405]) );
  DFF \xreg_reg[406]  ( .D(xin[405]), .CLK(clk), .RST(rst), .Q(xreg[406]) );
  DFF \xreg_reg[407]  ( .D(xin[406]), .CLK(clk), .RST(rst), .Q(xreg[407]) );
  DFF \xreg_reg[408]  ( .D(xin[407]), .CLK(clk), .RST(rst), .Q(xreg[408]) );
  DFF \xreg_reg[409]  ( .D(xin[408]), .CLK(clk), .RST(rst), .Q(xreg[409]) );
  DFF \xreg_reg[410]  ( .D(xin[409]), .CLK(clk), .RST(rst), .Q(xreg[410]) );
  DFF \xreg_reg[411]  ( .D(xin[410]), .CLK(clk), .RST(rst), .Q(xreg[411]) );
  DFF \xreg_reg[412]  ( .D(xin[411]), .CLK(clk), .RST(rst), .Q(xreg[412]) );
  DFF \xreg_reg[413]  ( .D(xin[412]), .CLK(clk), .RST(rst), .Q(xreg[413]) );
  DFF \xreg_reg[414]  ( .D(xin[413]), .CLK(clk), .RST(rst), .Q(xreg[414]) );
  DFF \xreg_reg[415]  ( .D(xin[414]), .CLK(clk), .RST(rst), .Q(xreg[415]) );
  DFF \xreg_reg[416]  ( .D(xin[415]), .CLK(clk), .RST(rst), .Q(xreg[416]) );
  DFF \xreg_reg[417]  ( .D(xin[416]), .CLK(clk), .RST(rst), .Q(xreg[417]) );
  DFF \xreg_reg[418]  ( .D(xin[417]), .CLK(clk), .RST(rst), .Q(xreg[418]) );
  DFF \xreg_reg[419]  ( .D(xin[418]), .CLK(clk), .RST(rst), .Q(xreg[419]) );
  DFF \xreg_reg[420]  ( .D(xin[419]), .CLK(clk), .RST(rst), .Q(xreg[420]) );
  DFF \xreg_reg[421]  ( .D(xin[420]), .CLK(clk), .RST(rst), .Q(xreg[421]) );
  DFF \xreg_reg[422]  ( .D(xin[421]), .CLK(clk), .RST(rst), .Q(xreg[422]) );
  DFF \xreg_reg[423]  ( .D(xin[422]), .CLK(clk), .RST(rst), .Q(xreg[423]) );
  DFF \xreg_reg[424]  ( .D(xin[423]), .CLK(clk), .RST(rst), .Q(xreg[424]) );
  DFF \xreg_reg[425]  ( .D(xin[424]), .CLK(clk), .RST(rst), .Q(xreg[425]) );
  DFF \xreg_reg[426]  ( .D(xin[425]), .CLK(clk), .RST(rst), .Q(xreg[426]) );
  DFF \xreg_reg[427]  ( .D(xin[426]), .CLK(clk), .RST(rst), .Q(xreg[427]) );
  DFF \xreg_reg[428]  ( .D(xin[427]), .CLK(clk), .RST(rst), .Q(xreg[428]) );
  DFF \xreg_reg[429]  ( .D(xin[428]), .CLK(clk), .RST(rst), .Q(xreg[429]) );
  DFF \xreg_reg[430]  ( .D(xin[429]), .CLK(clk), .RST(rst), .Q(xreg[430]) );
  DFF \xreg_reg[431]  ( .D(xin[430]), .CLK(clk), .RST(rst), .Q(xreg[431]) );
  DFF \xreg_reg[432]  ( .D(xin[431]), .CLK(clk), .RST(rst), .Q(xreg[432]) );
  DFF \xreg_reg[433]  ( .D(xin[432]), .CLK(clk), .RST(rst), .Q(xreg[433]) );
  DFF \xreg_reg[434]  ( .D(xin[433]), .CLK(clk), .RST(rst), .Q(xreg[434]) );
  DFF \xreg_reg[435]  ( .D(xin[434]), .CLK(clk), .RST(rst), .Q(xreg[435]) );
  DFF \xreg_reg[436]  ( .D(xin[435]), .CLK(clk), .RST(rst), .Q(xreg[436]) );
  DFF \xreg_reg[437]  ( .D(xin[436]), .CLK(clk), .RST(rst), .Q(xreg[437]) );
  DFF \xreg_reg[438]  ( .D(xin[437]), .CLK(clk), .RST(rst), .Q(xreg[438]) );
  DFF \xreg_reg[439]  ( .D(xin[438]), .CLK(clk), .RST(rst), .Q(xreg[439]) );
  DFF \xreg_reg[440]  ( .D(xin[439]), .CLK(clk), .RST(rst), .Q(xreg[440]) );
  DFF \xreg_reg[441]  ( .D(xin[440]), .CLK(clk), .RST(rst), .Q(xreg[441]) );
  DFF \xreg_reg[442]  ( .D(xin[441]), .CLK(clk), .RST(rst), .Q(xreg[442]) );
  DFF \xreg_reg[443]  ( .D(xin[442]), .CLK(clk), .RST(rst), .Q(xreg[443]) );
  DFF \xreg_reg[444]  ( .D(xin[443]), .CLK(clk), .RST(rst), .Q(xreg[444]) );
  DFF \xreg_reg[445]  ( .D(xin[444]), .CLK(clk), .RST(rst), .Q(xreg[445]) );
  DFF \xreg_reg[446]  ( .D(xin[445]), .CLK(clk), .RST(rst), .Q(xreg[446]) );
  DFF \xreg_reg[447]  ( .D(xin[446]), .CLK(clk), .RST(rst), .Q(xreg[447]) );
  DFF \xreg_reg[448]  ( .D(xin[447]), .CLK(clk), .RST(rst), .Q(xreg[448]) );
  DFF \xreg_reg[449]  ( .D(xin[448]), .CLK(clk), .RST(rst), .Q(xreg[449]) );
  DFF \xreg_reg[450]  ( .D(xin[449]), .CLK(clk), .RST(rst), .Q(xreg[450]) );
  DFF \xreg_reg[451]  ( .D(xin[450]), .CLK(clk), .RST(rst), .Q(xreg[451]) );
  DFF \xreg_reg[452]  ( .D(xin[451]), .CLK(clk), .RST(rst), .Q(xreg[452]) );
  DFF \xreg_reg[453]  ( .D(xin[452]), .CLK(clk), .RST(rst), .Q(xreg[453]) );
  DFF \xreg_reg[454]  ( .D(xin[453]), .CLK(clk), .RST(rst), .Q(xreg[454]) );
  DFF \xreg_reg[455]  ( .D(xin[454]), .CLK(clk), .RST(rst), .Q(xreg[455]) );
  DFF \xreg_reg[456]  ( .D(xin[455]), .CLK(clk), .RST(rst), .Q(xreg[456]) );
  DFF \xreg_reg[457]  ( .D(xin[456]), .CLK(clk), .RST(rst), .Q(xreg[457]) );
  DFF \xreg_reg[458]  ( .D(xin[457]), .CLK(clk), .RST(rst), .Q(xreg[458]) );
  DFF \xreg_reg[459]  ( .D(xin[458]), .CLK(clk), .RST(rst), .Q(xreg[459]) );
  DFF \xreg_reg[460]  ( .D(xin[459]), .CLK(clk), .RST(rst), .Q(xreg[460]) );
  DFF \xreg_reg[461]  ( .D(xin[460]), .CLK(clk), .RST(rst), .Q(xreg[461]) );
  DFF \xreg_reg[462]  ( .D(xin[461]), .CLK(clk), .RST(rst), .Q(xreg[462]) );
  DFF \xreg_reg[463]  ( .D(xin[462]), .CLK(clk), .RST(rst), .Q(xreg[463]) );
  DFF \xreg_reg[464]  ( .D(xin[463]), .CLK(clk), .RST(rst), .Q(xreg[464]) );
  DFF \xreg_reg[465]  ( .D(xin[464]), .CLK(clk), .RST(rst), .Q(xreg[465]) );
  DFF \xreg_reg[466]  ( .D(xin[465]), .CLK(clk), .RST(rst), .Q(xreg[466]) );
  DFF \xreg_reg[467]  ( .D(xin[466]), .CLK(clk), .RST(rst), .Q(xreg[467]) );
  DFF \xreg_reg[468]  ( .D(xin[467]), .CLK(clk), .RST(rst), .Q(xreg[468]) );
  DFF \xreg_reg[469]  ( .D(xin[468]), .CLK(clk), .RST(rst), .Q(xreg[469]) );
  DFF \xreg_reg[470]  ( .D(xin[469]), .CLK(clk), .RST(rst), .Q(xreg[470]) );
  DFF \xreg_reg[471]  ( .D(xin[470]), .CLK(clk), .RST(rst), .Q(xreg[471]) );
  DFF \xreg_reg[472]  ( .D(xin[471]), .CLK(clk), .RST(rst), .Q(xreg[472]) );
  DFF \xreg_reg[473]  ( .D(xin[472]), .CLK(clk), .RST(rst), .Q(xreg[473]) );
  DFF \xreg_reg[474]  ( .D(xin[473]), .CLK(clk), .RST(rst), .Q(xreg[474]) );
  DFF \xreg_reg[475]  ( .D(xin[474]), .CLK(clk), .RST(rst), .Q(xreg[475]) );
  DFF \xreg_reg[476]  ( .D(xin[475]), .CLK(clk), .RST(rst), .Q(xreg[476]) );
  DFF \xreg_reg[477]  ( .D(xin[476]), .CLK(clk), .RST(rst), .Q(xreg[477]) );
  DFF \xreg_reg[478]  ( .D(xin[477]), .CLK(clk), .RST(rst), .Q(xreg[478]) );
  DFF \xreg_reg[479]  ( .D(xin[478]), .CLK(clk), .RST(rst), .Q(xreg[479]) );
  DFF \xreg_reg[480]  ( .D(xin[479]), .CLK(clk), .RST(rst), .Q(xreg[480]) );
  DFF \xreg_reg[481]  ( .D(xin[480]), .CLK(clk), .RST(rst), .Q(xreg[481]) );
  DFF \xreg_reg[482]  ( .D(xin[481]), .CLK(clk), .RST(rst), .Q(xreg[482]) );
  DFF \xreg_reg[483]  ( .D(xin[482]), .CLK(clk), .RST(rst), .Q(xreg[483]) );
  DFF \xreg_reg[484]  ( .D(xin[483]), .CLK(clk), .RST(rst), .Q(xreg[484]) );
  DFF \xreg_reg[485]  ( .D(xin[484]), .CLK(clk), .RST(rst), .Q(xreg[485]) );
  DFF \xreg_reg[486]  ( .D(xin[485]), .CLK(clk), .RST(rst), .Q(xreg[486]) );
  DFF \xreg_reg[487]  ( .D(xin[486]), .CLK(clk), .RST(rst), .Q(xreg[487]) );
  DFF \xreg_reg[488]  ( .D(xin[487]), .CLK(clk), .RST(rst), .Q(xreg[488]) );
  DFF \xreg_reg[489]  ( .D(xin[488]), .CLK(clk), .RST(rst), .Q(xreg[489]) );
  DFF \xreg_reg[490]  ( .D(xin[489]), .CLK(clk), .RST(rst), .Q(xreg[490]) );
  DFF \xreg_reg[491]  ( .D(xin[490]), .CLK(clk), .RST(rst), .Q(xreg[491]) );
  DFF \xreg_reg[492]  ( .D(xin[491]), .CLK(clk), .RST(rst), .Q(xreg[492]) );
  DFF \xreg_reg[493]  ( .D(xin[492]), .CLK(clk), .RST(rst), .Q(xreg[493]) );
  DFF \xreg_reg[494]  ( .D(xin[493]), .CLK(clk), .RST(rst), .Q(xreg[494]) );
  DFF \xreg_reg[495]  ( .D(xin[494]), .CLK(clk), .RST(rst), .Q(xreg[495]) );
  DFF \xreg_reg[496]  ( .D(xin[495]), .CLK(clk), .RST(rst), .Q(xreg[496]) );
  DFF \xreg_reg[497]  ( .D(xin[496]), .CLK(clk), .RST(rst), .Q(xreg[497]) );
  DFF \xreg_reg[498]  ( .D(xin[497]), .CLK(clk), .RST(rst), .Q(xreg[498]) );
  DFF \xreg_reg[499]  ( .D(xin[498]), .CLK(clk), .RST(rst), .Q(xreg[499]) );
  DFF \xreg_reg[500]  ( .D(xin[499]), .CLK(clk), .RST(rst), .Q(xreg[500]) );
  DFF \xreg_reg[501]  ( .D(xin[500]), .CLK(clk), .RST(rst), .Q(xreg[501]) );
  DFF \xreg_reg[502]  ( .D(xin[501]), .CLK(clk), .RST(rst), .Q(xreg[502]) );
  DFF \xreg_reg[503]  ( .D(xin[502]), .CLK(clk), .RST(rst), .Q(xreg[503]) );
  DFF \xreg_reg[504]  ( .D(xin[503]), .CLK(clk), .RST(rst), .Q(xreg[504]) );
  DFF \xreg_reg[505]  ( .D(xin[504]), .CLK(clk), .RST(rst), .Q(xreg[505]) );
  DFF \xreg_reg[506]  ( .D(xin[505]), .CLK(clk), .RST(rst), .Q(xreg[506]) );
  DFF \xreg_reg[507]  ( .D(xin[506]), .CLK(clk), .RST(rst), .Q(xreg[507]) );
  DFF \xreg_reg[508]  ( .D(xin[507]), .CLK(clk), .RST(rst), .Q(xreg[508]) );
  DFF \xreg_reg[509]  ( .D(xin[508]), .CLK(clk), .RST(rst), .Q(xreg[509]) );
  DFF \xreg_reg[510]  ( .D(xin[509]), .CLK(clk), .RST(rst), .Q(xreg[510]) );
  DFF \xreg_reg[511]  ( .D(xin[510]), .CLK(clk), .RST(rst), .Q(xreg[511]) );
  DFF \xreg_reg[512]  ( .D(xin[511]), .CLK(clk), .RST(rst), .Q(xreg[512]) );
  DFF \xreg_reg[513]  ( .D(xin[512]), .CLK(clk), .RST(rst), .Q(xreg[513]) );
  DFF \xreg_reg[514]  ( .D(xin[513]), .CLK(clk), .RST(rst), .Q(xreg[514]) );
  DFF \xreg_reg[515]  ( .D(xin[514]), .CLK(clk), .RST(rst), .Q(xreg[515]) );
  DFF \xreg_reg[516]  ( .D(xin[515]), .CLK(clk), .RST(rst), .Q(xreg[516]) );
  DFF \xreg_reg[517]  ( .D(xin[516]), .CLK(clk), .RST(rst), .Q(xreg[517]) );
  DFF \xreg_reg[518]  ( .D(xin[517]), .CLK(clk), .RST(rst), .Q(xreg[518]) );
  DFF \xreg_reg[519]  ( .D(xin[518]), .CLK(clk), .RST(rst), .Q(xreg[519]) );
  DFF \xreg_reg[520]  ( .D(xin[519]), .CLK(clk), .RST(rst), .Q(xreg[520]) );
  DFF \xreg_reg[521]  ( .D(xin[520]), .CLK(clk), .RST(rst), .Q(xreg[521]) );
  DFF \xreg_reg[522]  ( .D(xin[521]), .CLK(clk), .RST(rst), .Q(xreg[522]) );
  DFF \xreg_reg[523]  ( .D(xin[522]), .CLK(clk), .RST(rst), .Q(xreg[523]) );
  DFF \xreg_reg[524]  ( .D(xin[523]), .CLK(clk), .RST(rst), .Q(xreg[524]) );
  DFF \xreg_reg[525]  ( .D(xin[524]), .CLK(clk), .RST(rst), .Q(xreg[525]) );
  DFF \xreg_reg[526]  ( .D(xin[525]), .CLK(clk), .RST(rst), .Q(xreg[526]) );
  DFF \xreg_reg[527]  ( .D(xin[526]), .CLK(clk), .RST(rst), .Q(xreg[527]) );
  DFF \xreg_reg[528]  ( .D(xin[527]), .CLK(clk), .RST(rst), .Q(xreg[528]) );
  DFF \xreg_reg[529]  ( .D(xin[528]), .CLK(clk), .RST(rst), .Q(xreg[529]) );
  DFF \xreg_reg[530]  ( .D(xin[529]), .CLK(clk), .RST(rst), .Q(xreg[530]) );
  DFF \xreg_reg[531]  ( .D(xin[530]), .CLK(clk), .RST(rst), .Q(xreg[531]) );
  DFF \xreg_reg[532]  ( .D(xin[531]), .CLK(clk), .RST(rst), .Q(xreg[532]) );
  DFF \xreg_reg[533]  ( .D(xin[532]), .CLK(clk), .RST(rst), .Q(xreg[533]) );
  DFF \xreg_reg[534]  ( .D(xin[533]), .CLK(clk), .RST(rst), .Q(xreg[534]) );
  DFF \xreg_reg[535]  ( .D(xin[534]), .CLK(clk), .RST(rst), .Q(xreg[535]) );
  DFF \xreg_reg[536]  ( .D(xin[535]), .CLK(clk), .RST(rst), .Q(xreg[536]) );
  DFF \xreg_reg[537]  ( .D(xin[536]), .CLK(clk), .RST(rst), .Q(xreg[537]) );
  DFF \xreg_reg[538]  ( .D(xin[537]), .CLK(clk), .RST(rst), .Q(xreg[538]) );
  DFF \xreg_reg[539]  ( .D(xin[538]), .CLK(clk), .RST(rst), .Q(xreg[539]) );
  DFF \xreg_reg[540]  ( .D(xin[539]), .CLK(clk), .RST(rst), .Q(xreg[540]) );
  DFF \xreg_reg[541]  ( .D(xin[540]), .CLK(clk), .RST(rst), .Q(xreg[541]) );
  DFF \xreg_reg[542]  ( .D(xin[541]), .CLK(clk), .RST(rst), .Q(xreg[542]) );
  DFF \xreg_reg[543]  ( .D(xin[542]), .CLK(clk), .RST(rst), .Q(xreg[543]) );
  DFF \xreg_reg[544]  ( .D(xin[543]), .CLK(clk), .RST(rst), .Q(xreg[544]) );
  DFF \xreg_reg[545]  ( .D(xin[544]), .CLK(clk), .RST(rst), .Q(xreg[545]) );
  DFF \xreg_reg[546]  ( .D(xin[545]), .CLK(clk), .RST(rst), .Q(xreg[546]) );
  DFF \xreg_reg[547]  ( .D(xin[546]), .CLK(clk), .RST(rst), .Q(xreg[547]) );
  DFF \xreg_reg[548]  ( .D(xin[547]), .CLK(clk), .RST(rst), .Q(xreg[548]) );
  DFF \xreg_reg[549]  ( .D(xin[548]), .CLK(clk), .RST(rst), .Q(xreg[549]) );
  DFF \xreg_reg[550]  ( .D(xin[549]), .CLK(clk), .RST(rst), .Q(xreg[550]) );
  DFF \xreg_reg[551]  ( .D(xin[550]), .CLK(clk), .RST(rst), .Q(xreg[551]) );
  DFF \xreg_reg[552]  ( .D(xin[551]), .CLK(clk), .RST(rst), .Q(xreg[552]) );
  DFF \xreg_reg[553]  ( .D(xin[552]), .CLK(clk), .RST(rst), .Q(xreg[553]) );
  DFF \xreg_reg[554]  ( .D(xin[553]), .CLK(clk), .RST(rst), .Q(xreg[554]) );
  DFF \xreg_reg[555]  ( .D(xin[554]), .CLK(clk), .RST(rst), .Q(xreg[555]) );
  DFF \xreg_reg[556]  ( .D(xin[555]), .CLK(clk), .RST(rst), .Q(xreg[556]) );
  DFF \xreg_reg[557]  ( .D(xin[556]), .CLK(clk), .RST(rst), .Q(xreg[557]) );
  DFF \xreg_reg[558]  ( .D(xin[557]), .CLK(clk), .RST(rst), .Q(xreg[558]) );
  DFF \xreg_reg[559]  ( .D(xin[558]), .CLK(clk), .RST(rst), .Q(xreg[559]) );
  DFF \xreg_reg[560]  ( .D(xin[559]), .CLK(clk), .RST(rst), .Q(xreg[560]) );
  DFF \xreg_reg[561]  ( .D(xin[560]), .CLK(clk), .RST(rst), .Q(xreg[561]) );
  DFF \xreg_reg[562]  ( .D(xin[561]), .CLK(clk), .RST(rst), .Q(xreg[562]) );
  DFF \xreg_reg[563]  ( .D(xin[562]), .CLK(clk), .RST(rst), .Q(xreg[563]) );
  DFF \xreg_reg[564]  ( .D(xin[563]), .CLK(clk), .RST(rst), .Q(xreg[564]) );
  DFF \xreg_reg[565]  ( .D(xin[564]), .CLK(clk), .RST(rst), .Q(xreg[565]) );
  DFF \xreg_reg[566]  ( .D(xin[565]), .CLK(clk), .RST(rst), .Q(xreg[566]) );
  DFF \xreg_reg[567]  ( .D(xin[566]), .CLK(clk), .RST(rst), .Q(xreg[567]) );
  DFF \xreg_reg[568]  ( .D(xin[567]), .CLK(clk), .RST(rst), .Q(xreg[568]) );
  DFF \xreg_reg[569]  ( .D(xin[568]), .CLK(clk), .RST(rst), .Q(xreg[569]) );
  DFF \xreg_reg[570]  ( .D(xin[569]), .CLK(clk), .RST(rst), .Q(xreg[570]) );
  DFF \xreg_reg[571]  ( .D(xin[570]), .CLK(clk), .RST(rst), .Q(xreg[571]) );
  DFF \xreg_reg[572]  ( .D(xin[571]), .CLK(clk), .RST(rst), .Q(xreg[572]) );
  DFF \xreg_reg[573]  ( .D(xin[572]), .CLK(clk), .RST(rst), .Q(xreg[573]) );
  DFF \xreg_reg[574]  ( .D(xin[573]), .CLK(clk), .RST(rst), .Q(xreg[574]) );
  DFF \xreg_reg[575]  ( .D(xin[574]), .CLK(clk), .RST(rst), .Q(xreg[575]) );
  DFF \xreg_reg[576]  ( .D(xin[575]), .CLK(clk), .RST(rst), .Q(xreg[576]) );
  DFF \xreg_reg[577]  ( .D(xin[576]), .CLK(clk), .RST(rst), .Q(xreg[577]) );
  DFF \xreg_reg[578]  ( .D(xin[577]), .CLK(clk), .RST(rst), .Q(xreg[578]) );
  DFF \xreg_reg[579]  ( .D(xin[578]), .CLK(clk), .RST(rst), .Q(xreg[579]) );
  DFF \xreg_reg[580]  ( .D(xin[579]), .CLK(clk), .RST(rst), .Q(xreg[580]) );
  DFF \xreg_reg[581]  ( .D(xin[580]), .CLK(clk), .RST(rst), .Q(xreg[581]) );
  DFF \xreg_reg[582]  ( .D(xin[581]), .CLK(clk), .RST(rst), .Q(xreg[582]) );
  DFF \xreg_reg[583]  ( .D(xin[582]), .CLK(clk), .RST(rst), .Q(xreg[583]) );
  DFF \xreg_reg[584]  ( .D(xin[583]), .CLK(clk), .RST(rst), .Q(xreg[584]) );
  DFF \xreg_reg[585]  ( .D(xin[584]), .CLK(clk), .RST(rst), .Q(xreg[585]) );
  DFF \xreg_reg[586]  ( .D(xin[585]), .CLK(clk), .RST(rst), .Q(xreg[586]) );
  DFF \xreg_reg[587]  ( .D(xin[586]), .CLK(clk), .RST(rst), .Q(xreg[587]) );
  DFF \xreg_reg[588]  ( .D(xin[587]), .CLK(clk), .RST(rst), .Q(xreg[588]) );
  DFF \xreg_reg[589]  ( .D(xin[588]), .CLK(clk), .RST(rst), .Q(xreg[589]) );
  DFF \xreg_reg[590]  ( .D(xin[589]), .CLK(clk), .RST(rst), .Q(xreg[590]) );
  DFF \xreg_reg[591]  ( .D(xin[590]), .CLK(clk), .RST(rst), .Q(xreg[591]) );
  DFF \xreg_reg[592]  ( .D(xin[591]), .CLK(clk), .RST(rst), .Q(xreg[592]) );
  DFF \xreg_reg[593]  ( .D(xin[592]), .CLK(clk), .RST(rst), .Q(xreg[593]) );
  DFF \xreg_reg[594]  ( .D(xin[593]), .CLK(clk), .RST(rst), .Q(xreg[594]) );
  DFF \xreg_reg[595]  ( .D(xin[594]), .CLK(clk), .RST(rst), .Q(xreg[595]) );
  DFF \xreg_reg[596]  ( .D(xin[595]), .CLK(clk), .RST(rst), .Q(xreg[596]) );
  DFF \xreg_reg[597]  ( .D(xin[596]), .CLK(clk), .RST(rst), .Q(xreg[597]) );
  DFF \xreg_reg[598]  ( .D(xin[597]), .CLK(clk), .RST(rst), .Q(xreg[598]) );
  DFF \xreg_reg[599]  ( .D(xin[598]), .CLK(clk), .RST(rst), .Q(xreg[599]) );
  DFF \xreg_reg[600]  ( .D(xin[599]), .CLK(clk), .RST(rst), .Q(xreg[600]) );
  DFF \xreg_reg[601]  ( .D(xin[600]), .CLK(clk), .RST(rst), .Q(xreg[601]) );
  DFF \xreg_reg[602]  ( .D(xin[601]), .CLK(clk), .RST(rst), .Q(xreg[602]) );
  DFF \xreg_reg[603]  ( .D(xin[602]), .CLK(clk), .RST(rst), .Q(xreg[603]) );
  DFF \xreg_reg[604]  ( .D(xin[603]), .CLK(clk), .RST(rst), .Q(xreg[604]) );
  DFF \xreg_reg[605]  ( .D(xin[604]), .CLK(clk), .RST(rst), .Q(xreg[605]) );
  DFF \xreg_reg[606]  ( .D(xin[605]), .CLK(clk), .RST(rst), .Q(xreg[606]) );
  DFF \xreg_reg[607]  ( .D(xin[606]), .CLK(clk), .RST(rst), .Q(xreg[607]) );
  DFF \xreg_reg[608]  ( .D(xin[607]), .CLK(clk), .RST(rst), .Q(xreg[608]) );
  DFF \xreg_reg[609]  ( .D(xin[608]), .CLK(clk), .RST(rst), .Q(xreg[609]) );
  DFF \xreg_reg[610]  ( .D(xin[609]), .CLK(clk), .RST(rst), .Q(xreg[610]) );
  DFF \xreg_reg[611]  ( .D(xin[610]), .CLK(clk), .RST(rst), .Q(xreg[611]) );
  DFF \xreg_reg[612]  ( .D(xin[611]), .CLK(clk), .RST(rst), .Q(xreg[612]) );
  DFF \xreg_reg[613]  ( .D(xin[612]), .CLK(clk), .RST(rst), .Q(xreg[613]) );
  DFF \xreg_reg[614]  ( .D(xin[613]), .CLK(clk), .RST(rst), .Q(xreg[614]) );
  DFF \xreg_reg[615]  ( .D(xin[614]), .CLK(clk), .RST(rst), .Q(xreg[615]) );
  DFF \xreg_reg[616]  ( .D(xin[615]), .CLK(clk), .RST(rst), .Q(xreg[616]) );
  DFF \xreg_reg[617]  ( .D(xin[616]), .CLK(clk), .RST(rst), .Q(xreg[617]) );
  DFF \xreg_reg[618]  ( .D(xin[617]), .CLK(clk), .RST(rst), .Q(xreg[618]) );
  DFF \xreg_reg[619]  ( .D(xin[618]), .CLK(clk), .RST(rst), .Q(xreg[619]) );
  DFF \xreg_reg[620]  ( .D(xin[619]), .CLK(clk), .RST(rst), .Q(xreg[620]) );
  DFF \xreg_reg[621]  ( .D(xin[620]), .CLK(clk), .RST(rst), .Q(xreg[621]) );
  DFF \xreg_reg[622]  ( .D(xin[621]), .CLK(clk), .RST(rst), .Q(xreg[622]) );
  DFF \xreg_reg[623]  ( .D(xin[622]), .CLK(clk), .RST(rst), .Q(xreg[623]) );
  DFF \xreg_reg[624]  ( .D(xin[623]), .CLK(clk), .RST(rst), .Q(xreg[624]) );
  DFF \xreg_reg[625]  ( .D(xin[624]), .CLK(clk), .RST(rst), .Q(xreg[625]) );
  DFF \xreg_reg[626]  ( .D(xin[625]), .CLK(clk), .RST(rst), .Q(xreg[626]) );
  DFF \xreg_reg[627]  ( .D(xin[626]), .CLK(clk), .RST(rst), .Q(xreg[627]) );
  DFF \xreg_reg[628]  ( .D(xin[627]), .CLK(clk), .RST(rst), .Q(xreg[628]) );
  DFF \xreg_reg[629]  ( .D(xin[628]), .CLK(clk), .RST(rst), .Q(xreg[629]) );
  DFF \xreg_reg[630]  ( .D(xin[629]), .CLK(clk), .RST(rst), .Q(xreg[630]) );
  DFF \xreg_reg[631]  ( .D(xin[630]), .CLK(clk), .RST(rst), .Q(xreg[631]) );
  DFF \xreg_reg[632]  ( .D(xin[631]), .CLK(clk), .RST(rst), .Q(xreg[632]) );
  DFF \xreg_reg[633]  ( .D(xin[632]), .CLK(clk), .RST(rst), .Q(xreg[633]) );
  DFF \xreg_reg[634]  ( .D(xin[633]), .CLK(clk), .RST(rst), .Q(xreg[634]) );
  DFF \xreg_reg[635]  ( .D(xin[634]), .CLK(clk), .RST(rst), .Q(xreg[635]) );
  DFF \xreg_reg[636]  ( .D(xin[635]), .CLK(clk), .RST(rst), .Q(xreg[636]) );
  DFF \xreg_reg[637]  ( .D(xin[636]), .CLK(clk), .RST(rst), .Q(xreg[637]) );
  DFF \xreg_reg[638]  ( .D(xin[637]), .CLK(clk), .RST(rst), .Q(xreg[638]) );
  DFF \xreg_reg[639]  ( .D(xin[638]), .CLK(clk), .RST(rst), .Q(xreg[639]) );
  DFF \xreg_reg[640]  ( .D(xin[639]), .CLK(clk), .RST(rst), .Q(xreg[640]) );
  DFF \xreg_reg[641]  ( .D(xin[640]), .CLK(clk), .RST(rst), .Q(xreg[641]) );
  DFF \xreg_reg[642]  ( .D(xin[641]), .CLK(clk), .RST(rst), .Q(xreg[642]) );
  DFF \xreg_reg[643]  ( .D(xin[642]), .CLK(clk), .RST(rst), .Q(xreg[643]) );
  DFF \xreg_reg[644]  ( .D(xin[643]), .CLK(clk), .RST(rst), .Q(xreg[644]) );
  DFF \xreg_reg[645]  ( .D(xin[644]), .CLK(clk), .RST(rst), .Q(xreg[645]) );
  DFF \xreg_reg[646]  ( .D(xin[645]), .CLK(clk), .RST(rst), .Q(xreg[646]) );
  DFF \xreg_reg[647]  ( .D(xin[646]), .CLK(clk), .RST(rst), .Q(xreg[647]) );
  DFF \xreg_reg[648]  ( .D(xin[647]), .CLK(clk), .RST(rst), .Q(xreg[648]) );
  DFF \xreg_reg[649]  ( .D(xin[648]), .CLK(clk), .RST(rst), .Q(xreg[649]) );
  DFF \xreg_reg[650]  ( .D(xin[649]), .CLK(clk), .RST(rst), .Q(xreg[650]) );
  DFF \xreg_reg[651]  ( .D(xin[650]), .CLK(clk), .RST(rst), .Q(xreg[651]) );
  DFF \xreg_reg[652]  ( .D(xin[651]), .CLK(clk), .RST(rst), .Q(xreg[652]) );
  DFF \xreg_reg[653]  ( .D(xin[652]), .CLK(clk), .RST(rst), .Q(xreg[653]) );
  DFF \xreg_reg[654]  ( .D(xin[653]), .CLK(clk), .RST(rst), .Q(xreg[654]) );
  DFF \xreg_reg[655]  ( .D(xin[654]), .CLK(clk), .RST(rst), .Q(xreg[655]) );
  DFF \xreg_reg[656]  ( .D(xin[655]), .CLK(clk), .RST(rst), .Q(xreg[656]) );
  DFF \xreg_reg[657]  ( .D(xin[656]), .CLK(clk), .RST(rst), .Q(xreg[657]) );
  DFF \xreg_reg[658]  ( .D(xin[657]), .CLK(clk), .RST(rst), .Q(xreg[658]) );
  DFF \xreg_reg[659]  ( .D(xin[658]), .CLK(clk), .RST(rst), .Q(xreg[659]) );
  DFF \xreg_reg[660]  ( .D(xin[659]), .CLK(clk), .RST(rst), .Q(xreg[660]) );
  DFF \xreg_reg[661]  ( .D(xin[660]), .CLK(clk), .RST(rst), .Q(xreg[661]) );
  DFF \xreg_reg[662]  ( .D(xin[661]), .CLK(clk), .RST(rst), .Q(xreg[662]) );
  DFF \xreg_reg[663]  ( .D(xin[662]), .CLK(clk), .RST(rst), .Q(xreg[663]) );
  DFF \xreg_reg[664]  ( .D(xin[663]), .CLK(clk), .RST(rst), .Q(xreg[664]) );
  DFF \xreg_reg[665]  ( .D(xin[664]), .CLK(clk), .RST(rst), .Q(xreg[665]) );
  DFF \xreg_reg[666]  ( .D(xin[665]), .CLK(clk), .RST(rst), .Q(xreg[666]) );
  DFF \xreg_reg[667]  ( .D(xin[666]), .CLK(clk), .RST(rst), .Q(xreg[667]) );
  DFF \xreg_reg[668]  ( .D(xin[667]), .CLK(clk), .RST(rst), .Q(xreg[668]) );
  DFF \xreg_reg[669]  ( .D(xin[668]), .CLK(clk), .RST(rst), .Q(xreg[669]) );
  DFF \xreg_reg[670]  ( .D(xin[669]), .CLK(clk), .RST(rst), .Q(xreg[670]) );
  DFF \xreg_reg[671]  ( .D(xin[670]), .CLK(clk), .RST(rst), .Q(xreg[671]) );
  DFF \xreg_reg[672]  ( .D(xin[671]), .CLK(clk), .RST(rst), .Q(xreg[672]) );
  DFF \xreg_reg[673]  ( .D(xin[672]), .CLK(clk), .RST(rst), .Q(xreg[673]) );
  DFF \xreg_reg[674]  ( .D(xin[673]), .CLK(clk), .RST(rst), .Q(xreg[674]) );
  DFF \xreg_reg[675]  ( .D(xin[674]), .CLK(clk), .RST(rst), .Q(xreg[675]) );
  DFF \xreg_reg[676]  ( .D(xin[675]), .CLK(clk), .RST(rst), .Q(xreg[676]) );
  DFF \xreg_reg[677]  ( .D(xin[676]), .CLK(clk), .RST(rst), .Q(xreg[677]) );
  DFF \xreg_reg[678]  ( .D(xin[677]), .CLK(clk), .RST(rst), .Q(xreg[678]) );
  DFF \xreg_reg[679]  ( .D(xin[678]), .CLK(clk), .RST(rst), .Q(xreg[679]) );
  DFF \xreg_reg[680]  ( .D(xin[679]), .CLK(clk), .RST(rst), .Q(xreg[680]) );
  DFF \xreg_reg[681]  ( .D(xin[680]), .CLK(clk), .RST(rst), .Q(xreg[681]) );
  DFF \xreg_reg[682]  ( .D(xin[681]), .CLK(clk), .RST(rst), .Q(xreg[682]) );
  DFF \xreg_reg[683]  ( .D(xin[682]), .CLK(clk), .RST(rst), .Q(xreg[683]) );
  DFF \xreg_reg[684]  ( .D(xin[683]), .CLK(clk), .RST(rst), .Q(xreg[684]) );
  DFF \xreg_reg[685]  ( .D(xin[684]), .CLK(clk), .RST(rst), .Q(xreg[685]) );
  DFF \xreg_reg[686]  ( .D(xin[685]), .CLK(clk), .RST(rst), .Q(xreg[686]) );
  DFF \xreg_reg[687]  ( .D(xin[686]), .CLK(clk), .RST(rst), .Q(xreg[687]) );
  DFF \xreg_reg[688]  ( .D(xin[687]), .CLK(clk), .RST(rst), .Q(xreg[688]) );
  DFF \xreg_reg[689]  ( .D(xin[688]), .CLK(clk), .RST(rst), .Q(xreg[689]) );
  DFF \xreg_reg[690]  ( .D(xin[689]), .CLK(clk), .RST(rst), .Q(xreg[690]) );
  DFF \xreg_reg[691]  ( .D(xin[690]), .CLK(clk), .RST(rst), .Q(xreg[691]) );
  DFF \xreg_reg[692]  ( .D(xin[691]), .CLK(clk), .RST(rst), .Q(xreg[692]) );
  DFF \xreg_reg[693]  ( .D(xin[692]), .CLK(clk), .RST(rst), .Q(xreg[693]) );
  DFF \xreg_reg[694]  ( .D(xin[693]), .CLK(clk), .RST(rst), .Q(xreg[694]) );
  DFF \xreg_reg[695]  ( .D(xin[694]), .CLK(clk), .RST(rst), .Q(xreg[695]) );
  DFF \xreg_reg[696]  ( .D(xin[695]), .CLK(clk), .RST(rst), .Q(xreg[696]) );
  DFF \xreg_reg[697]  ( .D(xin[696]), .CLK(clk), .RST(rst), .Q(xreg[697]) );
  DFF \xreg_reg[698]  ( .D(xin[697]), .CLK(clk), .RST(rst), .Q(xreg[698]) );
  DFF \xreg_reg[699]  ( .D(xin[698]), .CLK(clk), .RST(rst), .Q(xreg[699]) );
  DFF \xreg_reg[700]  ( .D(xin[699]), .CLK(clk), .RST(rst), .Q(xreg[700]) );
  DFF \xreg_reg[701]  ( .D(xin[700]), .CLK(clk), .RST(rst), .Q(xreg[701]) );
  DFF \xreg_reg[702]  ( .D(xin[701]), .CLK(clk), .RST(rst), .Q(xreg[702]) );
  DFF \xreg_reg[703]  ( .D(xin[702]), .CLK(clk), .RST(rst), .Q(xreg[703]) );
  DFF \xreg_reg[704]  ( .D(xin[703]), .CLK(clk), .RST(rst), .Q(xreg[704]) );
  DFF \xreg_reg[705]  ( .D(xin[704]), .CLK(clk), .RST(rst), .Q(xreg[705]) );
  DFF \xreg_reg[706]  ( .D(xin[705]), .CLK(clk), .RST(rst), .Q(xreg[706]) );
  DFF \xreg_reg[707]  ( .D(xin[706]), .CLK(clk), .RST(rst), .Q(xreg[707]) );
  DFF \xreg_reg[708]  ( .D(xin[707]), .CLK(clk), .RST(rst), .Q(xreg[708]) );
  DFF \xreg_reg[709]  ( .D(xin[708]), .CLK(clk), .RST(rst), .Q(xreg[709]) );
  DFF \xreg_reg[710]  ( .D(xin[709]), .CLK(clk), .RST(rst), .Q(xreg[710]) );
  DFF \xreg_reg[711]  ( .D(xin[710]), .CLK(clk), .RST(rst), .Q(xreg[711]) );
  DFF \xreg_reg[712]  ( .D(xin[711]), .CLK(clk), .RST(rst), .Q(xreg[712]) );
  DFF \xreg_reg[713]  ( .D(xin[712]), .CLK(clk), .RST(rst), .Q(xreg[713]) );
  DFF \xreg_reg[714]  ( .D(xin[713]), .CLK(clk), .RST(rst), .Q(xreg[714]) );
  DFF \xreg_reg[715]  ( .D(xin[714]), .CLK(clk), .RST(rst), .Q(xreg[715]) );
  DFF \xreg_reg[716]  ( .D(xin[715]), .CLK(clk), .RST(rst), .Q(xreg[716]) );
  DFF \xreg_reg[717]  ( .D(xin[716]), .CLK(clk), .RST(rst), .Q(xreg[717]) );
  DFF \xreg_reg[718]  ( .D(xin[717]), .CLK(clk), .RST(rst), .Q(xreg[718]) );
  DFF \xreg_reg[719]  ( .D(xin[718]), .CLK(clk), .RST(rst), .Q(xreg[719]) );
  DFF \xreg_reg[720]  ( .D(xin[719]), .CLK(clk), .RST(rst), .Q(xreg[720]) );
  DFF \xreg_reg[721]  ( .D(xin[720]), .CLK(clk), .RST(rst), .Q(xreg[721]) );
  DFF \xreg_reg[722]  ( .D(xin[721]), .CLK(clk), .RST(rst), .Q(xreg[722]) );
  DFF \xreg_reg[723]  ( .D(xin[722]), .CLK(clk), .RST(rst), .Q(xreg[723]) );
  DFF \xreg_reg[724]  ( .D(xin[723]), .CLK(clk), .RST(rst), .Q(xreg[724]) );
  DFF \xreg_reg[725]  ( .D(xin[724]), .CLK(clk), .RST(rst), .Q(xreg[725]) );
  DFF \xreg_reg[726]  ( .D(xin[725]), .CLK(clk), .RST(rst), .Q(xreg[726]) );
  DFF \xreg_reg[727]  ( .D(xin[726]), .CLK(clk), .RST(rst), .Q(xreg[727]) );
  DFF \xreg_reg[728]  ( .D(xin[727]), .CLK(clk), .RST(rst), .Q(xreg[728]) );
  DFF \xreg_reg[729]  ( .D(xin[728]), .CLK(clk), .RST(rst), .Q(xreg[729]) );
  DFF \xreg_reg[730]  ( .D(xin[729]), .CLK(clk), .RST(rst), .Q(xreg[730]) );
  DFF \xreg_reg[731]  ( .D(xin[730]), .CLK(clk), .RST(rst), .Q(xreg[731]) );
  DFF \xreg_reg[732]  ( .D(xin[731]), .CLK(clk), .RST(rst), .Q(xreg[732]) );
  DFF \xreg_reg[733]  ( .D(xin[732]), .CLK(clk), .RST(rst), .Q(xreg[733]) );
  DFF \xreg_reg[734]  ( .D(xin[733]), .CLK(clk), .RST(rst), .Q(xreg[734]) );
  DFF \xreg_reg[735]  ( .D(xin[734]), .CLK(clk), .RST(rst), .Q(xreg[735]) );
  DFF \xreg_reg[736]  ( .D(xin[735]), .CLK(clk), .RST(rst), .Q(xreg[736]) );
  DFF \xreg_reg[737]  ( .D(xin[736]), .CLK(clk), .RST(rst), .Q(xreg[737]) );
  DFF \xreg_reg[738]  ( .D(xin[737]), .CLK(clk), .RST(rst), .Q(xreg[738]) );
  DFF \xreg_reg[739]  ( .D(xin[738]), .CLK(clk), .RST(rst), .Q(xreg[739]) );
  DFF \xreg_reg[740]  ( .D(xin[739]), .CLK(clk), .RST(rst), .Q(xreg[740]) );
  DFF \xreg_reg[741]  ( .D(xin[740]), .CLK(clk), .RST(rst), .Q(xreg[741]) );
  DFF \xreg_reg[742]  ( .D(xin[741]), .CLK(clk), .RST(rst), .Q(xreg[742]) );
  DFF \xreg_reg[743]  ( .D(xin[742]), .CLK(clk), .RST(rst), .Q(xreg[743]) );
  DFF \xreg_reg[744]  ( .D(xin[743]), .CLK(clk), .RST(rst), .Q(xreg[744]) );
  DFF \xreg_reg[745]  ( .D(xin[744]), .CLK(clk), .RST(rst), .Q(xreg[745]) );
  DFF \xreg_reg[746]  ( .D(xin[745]), .CLK(clk), .RST(rst), .Q(xreg[746]) );
  DFF \xreg_reg[747]  ( .D(xin[746]), .CLK(clk), .RST(rst), .Q(xreg[747]) );
  DFF \xreg_reg[748]  ( .D(xin[747]), .CLK(clk), .RST(rst), .Q(xreg[748]) );
  DFF \xreg_reg[749]  ( .D(xin[748]), .CLK(clk), .RST(rst), .Q(xreg[749]) );
  DFF \xreg_reg[750]  ( .D(xin[749]), .CLK(clk), .RST(rst), .Q(xreg[750]) );
  DFF \xreg_reg[751]  ( .D(xin[750]), .CLK(clk), .RST(rst), .Q(xreg[751]) );
  DFF \xreg_reg[752]  ( .D(xin[751]), .CLK(clk), .RST(rst), .Q(xreg[752]) );
  DFF \xreg_reg[753]  ( .D(xin[752]), .CLK(clk), .RST(rst), .Q(xreg[753]) );
  DFF \xreg_reg[754]  ( .D(xin[753]), .CLK(clk), .RST(rst), .Q(xreg[754]) );
  DFF \xreg_reg[755]  ( .D(xin[754]), .CLK(clk), .RST(rst), .Q(xreg[755]) );
  DFF \xreg_reg[756]  ( .D(xin[755]), .CLK(clk), .RST(rst), .Q(xreg[756]) );
  DFF \xreg_reg[757]  ( .D(xin[756]), .CLK(clk), .RST(rst), .Q(xreg[757]) );
  DFF \xreg_reg[758]  ( .D(xin[757]), .CLK(clk), .RST(rst), .Q(xreg[758]) );
  DFF \xreg_reg[759]  ( .D(xin[758]), .CLK(clk), .RST(rst), .Q(xreg[759]) );
  DFF \xreg_reg[760]  ( .D(xin[759]), .CLK(clk), .RST(rst), .Q(xreg[760]) );
  DFF \xreg_reg[761]  ( .D(xin[760]), .CLK(clk), .RST(rst), .Q(xreg[761]) );
  DFF \xreg_reg[762]  ( .D(xin[761]), .CLK(clk), .RST(rst), .Q(xreg[762]) );
  DFF \xreg_reg[763]  ( .D(xin[762]), .CLK(clk), .RST(rst), .Q(xreg[763]) );
  DFF \xreg_reg[764]  ( .D(xin[763]), .CLK(clk), .RST(rst), .Q(xreg[764]) );
  DFF \xreg_reg[765]  ( .D(xin[764]), .CLK(clk), .RST(rst), .Q(xreg[765]) );
  DFF \xreg_reg[766]  ( .D(xin[765]), .CLK(clk), .RST(rst), .Q(xreg[766]) );
  DFF \xreg_reg[767]  ( .D(xin[766]), .CLK(clk), .RST(rst), .Q(xreg[767]) );
  DFF \xreg_reg[768]  ( .D(xin[767]), .CLK(clk), .RST(rst), .Q(xreg[768]) );
  DFF \xreg_reg[769]  ( .D(xin[768]), .CLK(clk), .RST(rst), .Q(xreg[769]) );
  DFF \xreg_reg[770]  ( .D(xin[769]), .CLK(clk), .RST(rst), .Q(xreg[770]) );
  DFF \xreg_reg[771]  ( .D(xin[770]), .CLK(clk), .RST(rst), .Q(xreg[771]) );
  DFF \xreg_reg[772]  ( .D(xin[771]), .CLK(clk), .RST(rst), .Q(xreg[772]) );
  DFF \xreg_reg[773]  ( .D(xin[772]), .CLK(clk), .RST(rst), .Q(xreg[773]) );
  DFF \xreg_reg[774]  ( .D(xin[773]), .CLK(clk), .RST(rst), .Q(xreg[774]) );
  DFF \xreg_reg[775]  ( .D(xin[774]), .CLK(clk), .RST(rst), .Q(xreg[775]) );
  DFF \xreg_reg[776]  ( .D(xin[775]), .CLK(clk), .RST(rst), .Q(xreg[776]) );
  DFF \xreg_reg[777]  ( .D(xin[776]), .CLK(clk), .RST(rst), .Q(xreg[777]) );
  DFF \xreg_reg[778]  ( .D(xin[777]), .CLK(clk), .RST(rst), .Q(xreg[778]) );
  DFF \xreg_reg[779]  ( .D(xin[778]), .CLK(clk), .RST(rst), .Q(xreg[779]) );
  DFF \xreg_reg[780]  ( .D(xin[779]), .CLK(clk), .RST(rst), .Q(xreg[780]) );
  DFF \xreg_reg[781]  ( .D(xin[780]), .CLK(clk), .RST(rst), .Q(xreg[781]) );
  DFF \xreg_reg[782]  ( .D(xin[781]), .CLK(clk), .RST(rst), .Q(xreg[782]) );
  DFF \xreg_reg[783]  ( .D(xin[782]), .CLK(clk), .RST(rst), .Q(xreg[783]) );
  DFF \xreg_reg[784]  ( .D(xin[783]), .CLK(clk), .RST(rst), .Q(xreg[784]) );
  DFF \xreg_reg[785]  ( .D(xin[784]), .CLK(clk), .RST(rst), .Q(xreg[785]) );
  DFF \xreg_reg[786]  ( .D(xin[785]), .CLK(clk), .RST(rst), .Q(xreg[786]) );
  DFF \xreg_reg[787]  ( .D(xin[786]), .CLK(clk), .RST(rst), .Q(xreg[787]) );
  DFF \xreg_reg[788]  ( .D(xin[787]), .CLK(clk), .RST(rst), .Q(xreg[788]) );
  DFF \xreg_reg[789]  ( .D(xin[788]), .CLK(clk), .RST(rst), .Q(xreg[789]) );
  DFF \xreg_reg[790]  ( .D(xin[789]), .CLK(clk), .RST(rst), .Q(xreg[790]) );
  DFF \xreg_reg[791]  ( .D(xin[790]), .CLK(clk), .RST(rst), .Q(xreg[791]) );
  DFF \xreg_reg[792]  ( .D(xin[791]), .CLK(clk), .RST(rst), .Q(xreg[792]) );
  DFF \xreg_reg[793]  ( .D(xin[792]), .CLK(clk), .RST(rst), .Q(xreg[793]) );
  DFF \xreg_reg[794]  ( .D(xin[793]), .CLK(clk), .RST(rst), .Q(xreg[794]) );
  DFF \xreg_reg[795]  ( .D(xin[794]), .CLK(clk), .RST(rst), .Q(xreg[795]) );
  DFF \xreg_reg[796]  ( .D(xin[795]), .CLK(clk), .RST(rst), .Q(xreg[796]) );
  DFF \xreg_reg[797]  ( .D(xin[796]), .CLK(clk), .RST(rst), .Q(xreg[797]) );
  DFF \xreg_reg[798]  ( .D(xin[797]), .CLK(clk), .RST(rst), .Q(xreg[798]) );
  DFF \xreg_reg[799]  ( .D(xin[798]), .CLK(clk), .RST(rst), .Q(xreg[799]) );
  DFF \xreg_reg[800]  ( .D(xin[799]), .CLK(clk), .RST(rst), .Q(xreg[800]) );
  DFF \xreg_reg[801]  ( .D(xin[800]), .CLK(clk), .RST(rst), .Q(xreg[801]) );
  DFF \xreg_reg[802]  ( .D(xin[801]), .CLK(clk), .RST(rst), .Q(xreg[802]) );
  DFF \xreg_reg[803]  ( .D(xin[802]), .CLK(clk), .RST(rst), .Q(xreg[803]) );
  DFF \xreg_reg[804]  ( .D(xin[803]), .CLK(clk), .RST(rst), .Q(xreg[804]) );
  DFF \xreg_reg[805]  ( .D(xin[804]), .CLK(clk), .RST(rst), .Q(xreg[805]) );
  DFF \xreg_reg[806]  ( .D(xin[805]), .CLK(clk), .RST(rst), .Q(xreg[806]) );
  DFF \xreg_reg[807]  ( .D(xin[806]), .CLK(clk), .RST(rst), .Q(xreg[807]) );
  DFF \xreg_reg[808]  ( .D(xin[807]), .CLK(clk), .RST(rst), .Q(xreg[808]) );
  DFF \xreg_reg[809]  ( .D(xin[808]), .CLK(clk), .RST(rst), .Q(xreg[809]) );
  DFF \xreg_reg[810]  ( .D(xin[809]), .CLK(clk), .RST(rst), .Q(xreg[810]) );
  DFF \xreg_reg[811]  ( .D(xin[810]), .CLK(clk), .RST(rst), .Q(xreg[811]) );
  DFF \xreg_reg[812]  ( .D(xin[811]), .CLK(clk), .RST(rst), .Q(xreg[812]) );
  DFF \xreg_reg[813]  ( .D(xin[812]), .CLK(clk), .RST(rst), .Q(xreg[813]) );
  DFF \xreg_reg[814]  ( .D(xin[813]), .CLK(clk), .RST(rst), .Q(xreg[814]) );
  DFF \xreg_reg[815]  ( .D(xin[814]), .CLK(clk), .RST(rst), .Q(xreg[815]) );
  DFF \xreg_reg[816]  ( .D(xin[815]), .CLK(clk), .RST(rst), .Q(xreg[816]) );
  DFF \xreg_reg[817]  ( .D(xin[816]), .CLK(clk), .RST(rst), .Q(xreg[817]) );
  DFF \xreg_reg[818]  ( .D(xin[817]), .CLK(clk), .RST(rst), .Q(xreg[818]) );
  DFF \xreg_reg[819]  ( .D(xin[818]), .CLK(clk), .RST(rst), .Q(xreg[819]) );
  DFF \xreg_reg[820]  ( .D(xin[819]), .CLK(clk), .RST(rst), .Q(xreg[820]) );
  DFF \xreg_reg[821]  ( .D(xin[820]), .CLK(clk), .RST(rst), .Q(xreg[821]) );
  DFF \xreg_reg[822]  ( .D(xin[821]), .CLK(clk), .RST(rst), .Q(xreg[822]) );
  DFF \xreg_reg[823]  ( .D(xin[822]), .CLK(clk), .RST(rst), .Q(xreg[823]) );
  DFF \xreg_reg[824]  ( .D(xin[823]), .CLK(clk), .RST(rst), .Q(xreg[824]) );
  DFF \xreg_reg[825]  ( .D(xin[824]), .CLK(clk), .RST(rst), .Q(xreg[825]) );
  DFF \xreg_reg[826]  ( .D(xin[825]), .CLK(clk), .RST(rst), .Q(xreg[826]) );
  DFF \xreg_reg[827]  ( .D(xin[826]), .CLK(clk), .RST(rst), .Q(xreg[827]) );
  DFF \xreg_reg[828]  ( .D(xin[827]), .CLK(clk), .RST(rst), .Q(xreg[828]) );
  DFF \xreg_reg[829]  ( .D(xin[828]), .CLK(clk), .RST(rst), .Q(xreg[829]) );
  DFF \xreg_reg[830]  ( .D(xin[829]), .CLK(clk), .RST(rst), .Q(xreg[830]) );
  DFF \xreg_reg[831]  ( .D(xin[830]), .CLK(clk), .RST(rst), .Q(xreg[831]) );
  DFF \xreg_reg[832]  ( .D(xin[831]), .CLK(clk), .RST(rst), .Q(xreg[832]) );
  DFF \xreg_reg[833]  ( .D(xin[832]), .CLK(clk), .RST(rst), .Q(xreg[833]) );
  DFF \xreg_reg[834]  ( .D(xin[833]), .CLK(clk), .RST(rst), .Q(xreg[834]) );
  DFF \xreg_reg[835]  ( .D(xin[834]), .CLK(clk), .RST(rst), .Q(xreg[835]) );
  DFF \xreg_reg[836]  ( .D(xin[835]), .CLK(clk), .RST(rst), .Q(xreg[836]) );
  DFF \xreg_reg[837]  ( .D(xin[836]), .CLK(clk), .RST(rst), .Q(xreg[837]) );
  DFF \xreg_reg[838]  ( .D(xin[837]), .CLK(clk), .RST(rst), .Q(xreg[838]) );
  DFF \xreg_reg[839]  ( .D(xin[838]), .CLK(clk), .RST(rst), .Q(xreg[839]) );
  DFF \xreg_reg[840]  ( .D(xin[839]), .CLK(clk), .RST(rst), .Q(xreg[840]) );
  DFF \xreg_reg[841]  ( .D(xin[840]), .CLK(clk), .RST(rst), .Q(xreg[841]) );
  DFF \xreg_reg[842]  ( .D(xin[841]), .CLK(clk), .RST(rst), .Q(xreg[842]) );
  DFF \xreg_reg[843]  ( .D(xin[842]), .CLK(clk), .RST(rst), .Q(xreg[843]) );
  DFF \xreg_reg[844]  ( .D(xin[843]), .CLK(clk), .RST(rst), .Q(xreg[844]) );
  DFF \xreg_reg[845]  ( .D(xin[844]), .CLK(clk), .RST(rst), .Q(xreg[845]) );
  DFF \xreg_reg[846]  ( .D(xin[845]), .CLK(clk), .RST(rst), .Q(xreg[846]) );
  DFF \xreg_reg[847]  ( .D(xin[846]), .CLK(clk), .RST(rst), .Q(xreg[847]) );
  DFF \xreg_reg[848]  ( .D(xin[847]), .CLK(clk), .RST(rst), .Q(xreg[848]) );
  DFF \xreg_reg[849]  ( .D(xin[848]), .CLK(clk), .RST(rst), .Q(xreg[849]) );
  DFF \xreg_reg[850]  ( .D(xin[849]), .CLK(clk), .RST(rst), .Q(xreg[850]) );
  DFF \xreg_reg[851]  ( .D(xin[850]), .CLK(clk), .RST(rst), .Q(xreg[851]) );
  DFF \xreg_reg[852]  ( .D(xin[851]), .CLK(clk), .RST(rst), .Q(xreg[852]) );
  DFF \xreg_reg[853]  ( .D(xin[852]), .CLK(clk), .RST(rst), .Q(xreg[853]) );
  DFF \xreg_reg[854]  ( .D(xin[853]), .CLK(clk), .RST(rst), .Q(xreg[854]) );
  DFF \xreg_reg[855]  ( .D(xin[854]), .CLK(clk), .RST(rst), .Q(xreg[855]) );
  DFF \xreg_reg[856]  ( .D(xin[855]), .CLK(clk), .RST(rst), .Q(xreg[856]) );
  DFF \xreg_reg[857]  ( .D(xin[856]), .CLK(clk), .RST(rst), .Q(xreg[857]) );
  DFF \xreg_reg[858]  ( .D(xin[857]), .CLK(clk), .RST(rst), .Q(xreg[858]) );
  DFF \xreg_reg[859]  ( .D(xin[858]), .CLK(clk), .RST(rst), .Q(xreg[859]) );
  DFF \xreg_reg[860]  ( .D(xin[859]), .CLK(clk), .RST(rst), .Q(xreg[860]) );
  DFF \xreg_reg[861]  ( .D(xin[860]), .CLK(clk), .RST(rst), .Q(xreg[861]) );
  DFF \xreg_reg[862]  ( .D(xin[861]), .CLK(clk), .RST(rst), .Q(xreg[862]) );
  DFF \xreg_reg[863]  ( .D(xin[862]), .CLK(clk), .RST(rst), .Q(xreg[863]) );
  DFF \xreg_reg[864]  ( .D(xin[863]), .CLK(clk), .RST(rst), .Q(xreg[864]) );
  DFF \xreg_reg[865]  ( .D(xin[864]), .CLK(clk), .RST(rst), .Q(xreg[865]) );
  DFF \xreg_reg[866]  ( .D(xin[865]), .CLK(clk), .RST(rst), .Q(xreg[866]) );
  DFF \xreg_reg[867]  ( .D(xin[866]), .CLK(clk), .RST(rst), .Q(xreg[867]) );
  DFF \xreg_reg[868]  ( .D(xin[867]), .CLK(clk), .RST(rst), .Q(xreg[868]) );
  DFF \xreg_reg[869]  ( .D(xin[868]), .CLK(clk), .RST(rst), .Q(xreg[869]) );
  DFF \xreg_reg[870]  ( .D(xin[869]), .CLK(clk), .RST(rst), .Q(xreg[870]) );
  DFF \xreg_reg[871]  ( .D(xin[870]), .CLK(clk), .RST(rst), .Q(xreg[871]) );
  DFF \xreg_reg[872]  ( .D(xin[871]), .CLK(clk), .RST(rst), .Q(xreg[872]) );
  DFF \xreg_reg[873]  ( .D(xin[872]), .CLK(clk), .RST(rst), .Q(xreg[873]) );
  DFF \xreg_reg[874]  ( .D(xin[873]), .CLK(clk), .RST(rst), .Q(xreg[874]) );
  DFF \xreg_reg[875]  ( .D(xin[874]), .CLK(clk), .RST(rst), .Q(xreg[875]) );
  DFF \xreg_reg[876]  ( .D(xin[875]), .CLK(clk), .RST(rst), .Q(xreg[876]) );
  DFF \xreg_reg[877]  ( .D(xin[876]), .CLK(clk), .RST(rst), .Q(xreg[877]) );
  DFF \xreg_reg[878]  ( .D(xin[877]), .CLK(clk), .RST(rst), .Q(xreg[878]) );
  DFF \xreg_reg[879]  ( .D(xin[878]), .CLK(clk), .RST(rst), .Q(xreg[879]) );
  DFF \xreg_reg[880]  ( .D(xin[879]), .CLK(clk), .RST(rst), .Q(xreg[880]) );
  DFF \xreg_reg[881]  ( .D(xin[880]), .CLK(clk), .RST(rst), .Q(xreg[881]) );
  DFF \xreg_reg[882]  ( .D(xin[881]), .CLK(clk), .RST(rst), .Q(xreg[882]) );
  DFF \xreg_reg[883]  ( .D(xin[882]), .CLK(clk), .RST(rst), .Q(xreg[883]) );
  DFF \xreg_reg[884]  ( .D(xin[883]), .CLK(clk), .RST(rst), .Q(xreg[884]) );
  DFF \xreg_reg[885]  ( .D(xin[884]), .CLK(clk), .RST(rst), .Q(xreg[885]) );
  DFF \xreg_reg[886]  ( .D(xin[885]), .CLK(clk), .RST(rst), .Q(xreg[886]) );
  DFF \xreg_reg[887]  ( .D(xin[886]), .CLK(clk), .RST(rst), .Q(xreg[887]) );
  DFF \xreg_reg[888]  ( .D(xin[887]), .CLK(clk), .RST(rst), .Q(xreg[888]) );
  DFF \xreg_reg[889]  ( .D(xin[888]), .CLK(clk), .RST(rst), .Q(xreg[889]) );
  DFF \xreg_reg[890]  ( .D(xin[889]), .CLK(clk), .RST(rst), .Q(xreg[890]) );
  DFF \xreg_reg[891]  ( .D(xin[890]), .CLK(clk), .RST(rst), .Q(xreg[891]) );
  DFF \xreg_reg[892]  ( .D(xin[891]), .CLK(clk), .RST(rst), .Q(xreg[892]) );
  DFF \xreg_reg[893]  ( .D(xin[892]), .CLK(clk), .RST(rst), .Q(xreg[893]) );
  DFF \xreg_reg[894]  ( .D(xin[893]), .CLK(clk), .RST(rst), .Q(xreg[894]) );
  DFF \xreg_reg[895]  ( .D(xin[894]), .CLK(clk), .RST(rst), .Q(xreg[895]) );
  DFF \xreg_reg[896]  ( .D(xin[895]), .CLK(clk), .RST(rst), .Q(xreg[896]) );
  DFF \xreg_reg[897]  ( .D(xin[896]), .CLK(clk), .RST(rst), .Q(xreg[897]) );
  DFF \xreg_reg[898]  ( .D(xin[897]), .CLK(clk), .RST(rst), .Q(xreg[898]) );
  DFF \xreg_reg[899]  ( .D(xin[898]), .CLK(clk), .RST(rst), .Q(xreg[899]) );
  DFF \xreg_reg[900]  ( .D(xin[899]), .CLK(clk), .RST(rst), .Q(xreg[900]) );
  DFF \xreg_reg[901]  ( .D(xin[900]), .CLK(clk), .RST(rst), .Q(xreg[901]) );
  DFF \xreg_reg[902]  ( .D(xin[901]), .CLK(clk), .RST(rst), .Q(xreg[902]) );
  DFF \xreg_reg[903]  ( .D(xin[902]), .CLK(clk), .RST(rst), .Q(xreg[903]) );
  DFF \xreg_reg[904]  ( .D(xin[903]), .CLK(clk), .RST(rst), .Q(xreg[904]) );
  DFF \xreg_reg[905]  ( .D(xin[904]), .CLK(clk), .RST(rst), .Q(xreg[905]) );
  DFF \xreg_reg[906]  ( .D(xin[905]), .CLK(clk), .RST(rst), .Q(xreg[906]) );
  DFF \xreg_reg[907]  ( .D(xin[906]), .CLK(clk), .RST(rst), .Q(xreg[907]) );
  DFF \xreg_reg[908]  ( .D(xin[907]), .CLK(clk), .RST(rst), .Q(xreg[908]) );
  DFF \xreg_reg[909]  ( .D(xin[908]), .CLK(clk), .RST(rst), .Q(xreg[909]) );
  DFF \xreg_reg[910]  ( .D(xin[909]), .CLK(clk), .RST(rst), .Q(xreg[910]) );
  DFF \xreg_reg[911]  ( .D(xin[910]), .CLK(clk), .RST(rst), .Q(xreg[911]) );
  DFF \xreg_reg[912]  ( .D(xin[911]), .CLK(clk), .RST(rst), .Q(xreg[912]) );
  DFF \xreg_reg[913]  ( .D(xin[912]), .CLK(clk), .RST(rst), .Q(xreg[913]) );
  DFF \xreg_reg[914]  ( .D(xin[913]), .CLK(clk), .RST(rst), .Q(xreg[914]) );
  DFF \xreg_reg[915]  ( .D(xin[914]), .CLK(clk), .RST(rst), .Q(xreg[915]) );
  DFF \xreg_reg[916]  ( .D(xin[915]), .CLK(clk), .RST(rst), .Q(xreg[916]) );
  DFF \xreg_reg[917]  ( .D(xin[916]), .CLK(clk), .RST(rst), .Q(xreg[917]) );
  DFF \xreg_reg[918]  ( .D(xin[917]), .CLK(clk), .RST(rst), .Q(xreg[918]) );
  DFF \xreg_reg[919]  ( .D(xin[918]), .CLK(clk), .RST(rst), .Q(xreg[919]) );
  DFF \xreg_reg[920]  ( .D(xin[919]), .CLK(clk), .RST(rst), .Q(xreg[920]) );
  DFF \xreg_reg[921]  ( .D(xin[920]), .CLK(clk), .RST(rst), .Q(xreg[921]) );
  DFF \xreg_reg[922]  ( .D(xin[921]), .CLK(clk), .RST(rst), .Q(xreg[922]) );
  DFF \xreg_reg[923]  ( .D(xin[922]), .CLK(clk), .RST(rst), .Q(xreg[923]) );
  DFF \xreg_reg[924]  ( .D(xin[923]), .CLK(clk), .RST(rst), .Q(xreg[924]) );
  DFF \xreg_reg[925]  ( .D(xin[924]), .CLK(clk), .RST(rst), .Q(xreg[925]) );
  DFF \xreg_reg[926]  ( .D(xin[925]), .CLK(clk), .RST(rst), .Q(xreg[926]) );
  DFF \xreg_reg[927]  ( .D(xin[926]), .CLK(clk), .RST(rst), .Q(xreg[927]) );
  DFF \xreg_reg[928]  ( .D(xin[927]), .CLK(clk), .RST(rst), .Q(xreg[928]) );
  DFF \xreg_reg[929]  ( .D(xin[928]), .CLK(clk), .RST(rst), .Q(xreg[929]) );
  DFF \xreg_reg[930]  ( .D(xin[929]), .CLK(clk), .RST(rst), .Q(xreg[930]) );
  DFF \xreg_reg[931]  ( .D(xin[930]), .CLK(clk), .RST(rst), .Q(xreg[931]) );
  DFF \xreg_reg[932]  ( .D(xin[931]), .CLK(clk), .RST(rst), .Q(xreg[932]) );
  DFF \xreg_reg[933]  ( .D(xin[932]), .CLK(clk), .RST(rst), .Q(xreg[933]) );
  DFF \xreg_reg[934]  ( .D(xin[933]), .CLK(clk), .RST(rst), .Q(xreg[934]) );
  DFF \xreg_reg[935]  ( .D(xin[934]), .CLK(clk), .RST(rst), .Q(xreg[935]) );
  DFF \xreg_reg[936]  ( .D(xin[935]), .CLK(clk), .RST(rst), .Q(xreg[936]) );
  DFF \xreg_reg[937]  ( .D(xin[936]), .CLK(clk), .RST(rst), .Q(xreg[937]) );
  DFF \xreg_reg[938]  ( .D(xin[937]), .CLK(clk), .RST(rst), .Q(xreg[938]) );
  DFF \xreg_reg[939]  ( .D(xin[938]), .CLK(clk), .RST(rst), .Q(xreg[939]) );
  DFF \xreg_reg[940]  ( .D(xin[939]), .CLK(clk), .RST(rst), .Q(xreg[940]) );
  DFF \xreg_reg[941]  ( .D(xin[940]), .CLK(clk), .RST(rst), .Q(xreg[941]) );
  DFF \xreg_reg[942]  ( .D(xin[941]), .CLK(clk), .RST(rst), .Q(xreg[942]) );
  DFF \xreg_reg[943]  ( .D(xin[942]), .CLK(clk), .RST(rst), .Q(xreg[943]) );
  DFF \xreg_reg[944]  ( .D(xin[943]), .CLK(clk), .RST(rst), .Q(xreg[944]) );
  DFF \xreg_reg[945]  ( .D(xin[944]), .CLK(clk), .RST(rst), .Q(xreg[945]) );
  DFF \xreg_reg[946]  ( .D(xin[945]), .CLK(clk), .RST(rst), .Q(xreg[946]) );
  DFF \xreg_reg[947]  ( .D(xin[946]), .CLK(clk), .RST(rst), .Q(xreg[947]) );
  DFF \xreg_reg[948]  ( .D(xin[947]), .CLK(clk), .RST(rst), .Q(xreg[948]) );
  DFF \xreg_reg[949]  ( .D(xin[948]), .CLK(clk), .RST(rst), .Q(xreg[949]) );
  DFF \xreg_reg[950]  ( .D(xin[949]), .CLK(clk), .RST(rst), .Q(xreg[950]) );
  DFF \xreg_reg[951]  ( .D(xin[950]), .CLK(clk), .RST(rst), .Q(xreg[951]) );
  DFF \xreg_reg[952]  ( .D(xin[951]), .CLK(clk), .RST(rst), .Q(xreg[952]) );
  DFF \xreg_reg[953]  ( .D(xin[952]), .CLK(clk), .RST(rst), .Q(xreg[953]) );
  DFF \xreg_reg[954]  ( .D(xin[953]), .CLK(clk), .RST(rst), .Q(xreg[954]) );
  DFF \xreg_reg[955]  ( .D(xin[954]), .CLK(clk), .RST(rst), .Q(xreg[955]) );
  DFF \xreg_reg[956]  ( .D(xin[955]), .CLK(clk), .RST(rst), .Q(xreg[956]) );
  DFF \xreg_reg[957]  ( .D(xin[956]), .CLK(clk), .RST(rst), .Q(xreg[957]) );
  DFF \xreg_reg[958]  ( .D(xin[957]), .CLK(clk), .RST(rst), .Q(xreg[958]) );
  DFF \xreg_reg[959]  ( .D(xin[958]), .CLK(clk), .RST(rst), .Q(xreg[959]) );
  DFF \xreg_reg[960]  ( .D(xin[959]), .CLK(clk), .RST(rst), .Q(xreg[960]) );
  DFF \xreg_reg[961]  ( .D(xin[960]), .CLK(clk), .RST(rst), .Q(xreg[961]) );
  DFF \xreg_reg[962]  ( .D(xin[961]), .CLK(clk), .RST(rst), .Q(xreg[962]) );
  DFF \xreg_reg[963]  ( .D(xin[962]), .CLK(clk), .RST(rst), .Q(xreg[963]) );
  DFF \xreg_reg[964]  ( .D(xin[963]), .CLK(clk), .RST(rst), .Q(xreg[964]) );
  DFF \xreg_reg[965]  ( .D(xin[964]), .CLK(clk), .RST(rst), .Q(xreg[965]) );
  DFF \xreg_reg[966]  ( .D(xin[965]), .CLK(clk), .RST(rst), .Q(xreg[966]) );
  DFF \xreg_reg[967]  ( .D(xin[966]), .CLK(clk), .RST(rst), .Q(xreg[967]) );
  DFF \xreg_reg[968]  ( .D(xin[967]), .CLK(clk), .RST(rst), .Q(xreg[968]) );
  DFF \xreg_reg[969]  ( .D(xin[968]), .CLK(clk), .RST(rst), .Q(xreg[969]) );
  DFF \xreg_reg[970]  ( .D(xin[969]), .CLK(clk), .RST(rst), .Q(xreg[970]) );
  DFF \xreg_reg[971]  ( .D(xin[970]), .CLK(clk), .RST(rst), .Q(xreg[971]) );
  DFF \xreg_reg[972]  ( .D(xin[971]), .CLK(clk), .RST(rst), .Q(xreg[972]) );
  DFF \xreg_reg[973]  ( .D(xin[972]), .CLK(clk), .RST(rst), .Q(xreg[973]) );
  DFF \xreg_reg[974]  ( .D(xin[973]), .CLK(clk), .RST(rst), .Q(xreg[974]) );
  DFF \xreg_reg[975]  ( .D(xin[974]), .CLK(clk), .RST(rst), .Q(xreg[975]) );
  DFF \xreg_reg[976]  ( .D(xin[975]), .CLK(clk), .RST(rst), .Q(xreg[976]) );
  DFF \xreg_reg[977]  ( .D(xin[976]), .CLK(clk), .RST(rst), .Q(xreg[977]) );
  DFF \xreg_reg[978]  ( .D(xin[977]), .CLK(clk), .RST(rst), .Q(xreg[978]) );
  DFF \xreg_reg[979]  ( .D(xin[978]), .CLK(clk), .RST(rst), .Q(xreg[979]) );
  DFF \xreg_reg[980]  ( .D(xin[979]), .CLK(clk), .RST(rst), .Q(xreg[980]) );
  DFF \xreg_reg[981]  ( .D(xin[980]), .CLK(clk), .RST(rst), .Q(xreg[981]) );
  DFF \xreg_reg[982]  ( .D(xin[981]), .CLK(clk), .RST(rst), .Q(xreg[982]) );
  DFF \xreg_reg[983]  ( .D(xin[982]), .CLK(clk), .RST(rst), .Q(xreg[983]) );
  DFF \xreg_reg[984]  ( .D(xin[983]), .CLK(clk), .RST(rst), .Q(xreg[984]) );
  DFF \xreg_reg[985]  ( .D(xin[984]), .CLK(clk), .RST(rst), .Q(xreg[985]) );
  DFF \xreg_reg[986]  ( .D(xin[985]), .CLK(clk), .RST(rst), .Q(xreg[986]) );
  DFF \xreg_reg[987]  ( .D(xin[986]), .CLK(clk), .RST(rst), .Q(xreg[987]) );
  DFF \xreg_reg[988]  ( .D(xin[987]), .CLK(clk), .RST(rst), .Q(xreg[988]) );
  DFF \xreg_reg[989]  ( .D(xin[988]), .CLK(clk), .RST(rst), .Q(xreg[989]) );
  DFF \xreg_reg[990]  ( .D(xin[989]), .CLK(clk), .RST(rst), .Q(xreg[990]) );
  DFF \xreg_reg[991]  ( .D(xin[990]), .CLK(clk), .RST(rst), .Q(xreg[991]) );
  DFF \xreg_reg[992]  ( .D(xin[991]), .CLK(clk), .RST(rst), .Q(xreg[992]) );
  DFF \xreg_reg[993]  ( .D(xin[992]), .CLK(clk), .RST(rst), .Q(xreg[993]) );
  DFF \xreg_reg[994]  ( .D(xin[993]), .CLK(clk), .RST(rst), .Q(xreg[994]) );
  DFF \xreg_reg[995]  ( .D(xin[994]), .CLK(clk), .RST(rst), .Q(xreg[995]) );
  DFF \xreg_reg[996]  ( .D(xin[995]), .CLK(clk), .RST(rst), .Q(xreg[996]) );
  DFF \xreg_reg[997]  ( .D(xin[996]), .CLK(clk), .RST(rst), .Q(xreg[997]) );
  DFF \xreg_reg[998]  ( .D(xin[997]), .CLK(clk), .RST(rst), .Q(xreg[998]) );
  DFF \xreg_reg[999]  ( .D(xin[998]), .CLK(clk), .RST(rst), .Q(xreg[999]) );
  DFF \xreg_reg[1000]  ( .D(xin[999]), .CLK(clk), .RST(rst), .Q(xreg[1000]) );
  DFF \xreg_reg[1001]  ( .D(xin[1000]), .CLK(clk), .RST(rst), .Q(xreg[1001])
         );
  DFF \xreg_reg[1002]  ( .D(xin[1001]), .CLK(clk), .RST(rst), .Q(xreg[1002])
         );
  DFF \xreg_reg[1003]  ( .D(xin[1002]), .CLK(clk), .RST(rst), .Q(xreg[1003])
         );
  DFF \xreg_reg[1004]  ( .D(xin[1003]), .CLK(clk), .RST(rst), .Q(xreg[1004])
         );
  DFF \xreg_reg[1005]  ( .D(xin[1004]), .CLK(clk), .RST(rst), .Q(xreg[1005])
         );
  DFF \xreg_reg[1006]  ( .D(xin[1005]), .CLK(clk), .RST(rst), .Q(xreg[1006])
         );
  DFF \xreg_reg[1007]  ( .D(xin[1006]), .CLK(clk), .RST(rst), .Q(xreg[1007])
         );
  DFF \xreg_reg[1008]  ( .D(xin[1007]), .CLK(clk), .RST(rst), .Q(xreg[1008])
         );
  DFF \xreg_reg[1009]  ( .D(xin[1008]), .CLK(clk), .RST(rst), .Q(xreg[1009])
         );
  DFF \xreg_reg[1010]  ( .D(xin[1009]), .CLK(clk), .RST(rst), .Q(xreg[1010])
         );
  DFF \xreg_reg[1011]  ( .D(xin[1010]), .CLK(clk), .RST(rst), .Q(xreg[1011])
         );
  DFF \xreg_reg[1012]  ( .D(xin[1011]), .CLK(clk), .RST(rst), .Q(xreg[1012])
         );
  DFF \xreg_reg[1013]  ( .D(xin[1012]), .CLK(clk), .RST(rst), .Q(xreg[1013])
         );
  DFF \xreg_reg[1014]  ( .D(xin[1013]), .CLK(clk), .RST(rst), .Q(xreg[1014])
         );
  DFF \xreg_reg[1015]  ( .D(xin[1014]), .CLK(clk), .RST(rst), .Q(xreg[1015])
         );
  DFF \xreg_reg[1016]  ( .D(xin[1015]), .CLK(clk), .RST(rst), .Q(xreg[1016])
         );
  DFF \xreg_reg[1017]  ( .D(xin[1016]), .CLK(clk), .RST(rst), .Q(xreg[1017])
         );
  DFF \xreg_reg[1018]  ( .D(xin[1017]), .CLK(clk), .RST(rst), .Q(xreg[1018])
         );
  DFF \xreg_reg[1019]  ( .D(xin[1018]), .CLK(clk), .RST(rst), .Q(xreg[1019])
         );
  DFF \xreg_reg[1020]  ( .D(xin[1019]), .CLK(clk), .RST(rst), .Q(xreg[1020])
         );
  DFF \xreg_reg[1021]  ( .D(xin[1020]), .CLK(clk), .RST(rst), .Q(xreg[1021])
         );
  DFF \xreg_reg[1022]  ( .D(xin[1021]), .CLK(clk), .RST(rst), .Q(xreg[1022])
         );
  DFF \xreg_reg[1023]  ( .D(xin[1022]), .CLK(clk), .RST(rst), .Q(xreg[1023])
         );
  DFF \zreg_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .Q(zreg[0]) );
  DFF \zreg_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .Q(zreg[1]) );
  DFF \zreg_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .Q(zreg[2]) );
  DFF \zreg_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .Q(zreg[3]) );
  DFF \zreg_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .Q(zreg[4]) );
  DFF \zreg_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .Q(zreg[5]) );
  DFF \zreg_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .Q(zreg[6]) );
  DFF \zreg_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .Q(zreg[7]) );
  DFF \zreg_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .Q(zreg[8]) );
  DFF \zreg_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .Q(zreg[9]) );
  DFF \zreg_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .Q(zreg[10]) );
  DFF \zreg_reg[11]  ( .D(o[11]), .CLK(clk), .RST(rst), .Q(zreg[11]) );
  DFF \zreg_reg[12]  ( .D(o[12]), .CLK(clk), .RST(rst), .Q(zreg[12]) );
  DFF \zreg_reg[13]  ( .D(o[13]), .CLK(clk), .RST(rst), .Q(zreg[13]) );
  DFF \zreg_reg[14]  ( .D(o[14]), .CLK(clk), .RST(rst), .Q(zreg[14]) );
  DFF \zreg_reg[15]  ( .D(o[15]), .CLK(clk), .RST(rst), .Q(zreg[15]) );
  DFF \zreg_reg[16]  ( .D(o[16]), .CLK(clk), .RST(rst), .Q(zreg[16]) );
  DFF \zreg_reg[17]  ( .D(o[17]), .CLK(clk), .RST(rst), .Q(zreg[17]) );
  DFF \zreg_reg[18]  ( .D(o[18]), .CLK(clk), .RST(rst), .Q(zreg[18]) );
  DFF \zreg_reg[19]  ( .D(o[19]), .CLK(clk), .RST(rst), .Q(zreg[19]) );
  DFF \zreg_reg[20]  ( .D(o[20]), .CLK(clk), .RST(rst), .Q(zreg[20]) );
  DFF \zreg_reg[21]  ( .D(o[21]), .CLK(clk), .RST(rst), .Q(zreg[21]) );
  DFF \zreg_reg[22]  ( .D(o[22]), .CLK(clk), .RST(rst), .Q(zreg[22]) );
  DFF \zreg_reg[23]  ( .D(o[23]), .CLK(clk), .RST(rst), .Q(zreg[23]) );
  DFF \zreg_reg[24]  ( .D(o[24]), .CLK(clk), .RST(rst), .Q(zreg[24]) );
  DFF \zreg_reg[25]  ( .D(o[25]), .CLK(clk), .RST(rst), .Q(zreg[25]) );
  DFF \zreg_reg[26]  ( .D(o[26]), .CLK(clk), .RST(rst), .Q(zreg[26]) );
  DFF \zreg_reg[27]  ( .D(o[27]), .CLK(clk), .RST(rst), .Q(zreg[27]) );
  DFF \zreg_reg[28]  ( .D(o[28]), .CLK(clk), .RST(rst), .Q(zreg[28]) );
  DFF \zreg_reg[29]  ( .D(o[29]), .CLK(clk), .RST(rst), .Q(zreg[29]) );
  DFF \zreg_reg[30]  ( .D(o[30]), .CLK(clk), .RST(rst), .Q(zreg[30]) );
  DFF \zreg_reg[31]  ( .D(o[31]), .CLK(clk), .RST(rst), .Q(zreg[31]) );
  DFF \zreg_reg[32]  ( .D(o[32]), .CLK(clk), .RST(rst), .Q(zreg[32]) );
  DFF \zreg_reg[33]  ( .D(o[33]), .CLK(clk), .RST(rst), .Q(zreg[33]) );
  DFF \zreg_reg[34]  ( .D(o[34]), .CLK(clk), .RST(rst), .Q(zreg[34]) );
  DFF \zreg_reg[35]  ( .D(o[35]), .CLK(clk), .RST(rst), .Q(zreg[35]) );
  DFF \zreg_reg[36]  ( .D(o[36]), .CLK(clk), .RST(rst), .Q(zreg[36]) );
  DFF \zreg_reg[37]  ( .D(o[37]), .CLK(clk), .RST(rst), .Q(zreg[37]) );
  DFF \zreg_reg[38]  ( .D(o[38]), .CLK(clk), .RST(rst), .Q(zreg[38]) );
  DFF \zreg_reg[39]  ( .D(o[39]), .CLK(clk), .RST(rst), .Q(zreg[39]) );
  DFF \zreg_reg[40]  ( .D(o[40]), .CLK(clk), .RST(rst), .Q(zreg[40]) );
  DFF \zreg_reg[41]  ( .D(o[41]), .CLK(clk), .RST(rst), .Q(zreg[41]) );
  DFF \zreg_reg[42]  ( .D(o[42]), .CLK(clk), .RST(rst), .Q(zreg[42]) );
  DFF \zreg_reg[43]  ( .D(o[43]), .CLK(clk), .RST(rst), .Q(zreg[43]) );
  DFF \zreg_reg[44]  ( .D(o[44]), .CLK(clk), .RST(rst), .Q(zreg[44]) );
  DFF \zreg_reg[45]  ( .D(o[45]), .CLK(clk), .RST(rst), .Q(zreg[45]) );
  DFF \zreg_reg[46]  ( .D(o[46]), .CLK(clk), .RST(rst), .Q(zreg[46]) );
  DFF \zreg_reg[47]  ( .D(o[47]), .CLK(clk), .RST(rst), .Q(zreg[47]) );
  DFF \zreg_reg[48]  ( .D(o[48]), .CLK(clk), .RST(rst), .Q(zreg[48]) );
  DFF \zreg_reg[49]  ( .D(o[49]), .CLK(clk), .RST(rst), .Q(zreg[49]) );
  DFF \zreg_reg[50]  ( .D(o[50]), .CLK(clk), .RST(rst), .Q(zreg[50]) );
  DFF \zreg_reg[51]  ( .D(o[51]), .CLK(clk), .RST(rst), .Q(zreg[51]) );
  DFF \zreg_reg[52]  ( .D(o[52]), .CLK(clk), .RST(rst), .Q(zreg[52]) );
  DFF \zreg_reg[53]  ( .D(o[53]), .CLK(clk), .RST(rst), .Q(zreg[53]) );
  DFF \zreg_reg[54]  ( .D(o[54]), .CLK(clk), .RST(rst), .Q(zreg[54]) );
  DFF \zreg_reg[55]  ( .D(o[55]), .CLK(clk), .RST(rst), .Q(zreg[55]) );
  DFF \zreg_reg[56]  ( .D(o[56]), .CLK(clk), .RST(rst), .Q(zreg[56]) );
  DFF \zreg_reg[57]  ( .D(o[57]), .CLK(clk), .RST(rst), .Q(zreg[57]) );
  DFF \zreg_reg[58]  ( .D(o[58]), .CLK(clk), .RST(rst), .Q(zreg[58]) );
  DFF \zreg_reg[59]  ( .D(o[59]), .CLK(clk), .RST(rst), .Q(zreg[59]) );
  DFF \zreg_reg[60]  ( .D(o[60]), .CLK(clk), .RST(rst), .Q(zreg[60]) );
  DFF \zreg_reg[61]  ( .D(o[61]), .CLK(clk), .RST(rst), .Q(zreg[61]) );
  DFF \zreg_reg[62]  ( .D(o[62]), .CLK(clk), .RST(rst), .Q(zreg[62]) );
  DFF \zreg_reg[63]  ( .D(o[63]), .CLK(clk), .RST(rst), .Q(zreg[63]) );
  DFF \zreg_reg[64]  ( .D(o[64]), .CLK(clk), .RST(rst), .Q(zreg[64]) );
  DFF \zreg_reg[65]  ( .D(o[65]), .CLK(clk), .RST(rst), .Q(zreg[65]) );
  DFF \zreg_reg[66]  ( .D(o[66]), .CLK(clk), .RST(rst), .Q(zreg[66]) );
  DFF \zreg_reg[67]  ( .D(o[67]), .CLK(clk), .RST(rst), .Q(zreg[67]) );
  DFF \zreg_reg[68]  ( .D(o[68]), .CLK(clk), .RST(rst), .Q(zreg[68]) );
  DFF \zreg_reg[69]  ( .D(o[69]), .CLK(clk), .RST(rst), .Q(zreg[69]) );
  DFF \zreg_reg[70]  ( .D(o[70]), .CLK(clk), .RST(rst), .Q(zreg[70]) );
  DFF \zreg_reg[71]  ( .D(o[71]), .CLK(clk), .RST(rst), .Q(zreg[71]) );
  DFF \zreg_reg[72]  ( .D(o[72]), .CLK(clk), .RST(rst), .Q(zreg[72]) );
  DFF \zreg_reg[73]  ( .D(o[73]), .CLK(clk), .RST(rst), .Q(zreg[73]) );
  DFF \zreg_reg[74]  ( .D(o[74]), .CLK(clk), .RST(rst), .Q(zreg[74]) );
  DFF \zreg_reg[75]  ( .D(o[75]), .CLK(clk), .RST(rst), .Q(zreg[75]) );
  DFF \zreg_reg[76]  ( .D(o[76]), .CLK(clk), .RST(rst), .Q(zreg[76]) );
  DFF \zreg_reg[77]  ( .D(o[77]), .CLK(clk), .RST(rst), .Q(zreg[77]) );
  DFF \zreg_reg[78]  ( .D(o[78]), .CLK(clk), .RST(rst), .Q(zreg[78]) );
  DFF \zreg_reg[79]  ( .D(o[79]), .CLK(clk), .RST(rst), .Q(zreg[79]) );
  DFF \zreg_reg[80]  ( .D(o[80]), .CLK(clk), .RST(rst), .Q(zreg[80]) );
  DFF \zreg_reg[81]  ( .D(o[81]), .CLK(clk), .RST(rst), .Q(zreg[81]) );
  DFF \zreg_reg[82]  ( .D(o[82]), .CLK(clk), .RST(rst), .Q(zreg[82]) );
  DFF \zreg_reg[83]  ( .D(o[83]), .CLK(clk), .RST(rst), .Q(zreg[83]) );
  DFF \zreg_reg[84]  ( .D(o[84]), .CLK(clk), .RST(rst), .Q(zreg[84]) );
  DFF \zreg_reg[85]  ( .D(o[85]), .CLK(clk), .RST(rst), .Q(zreg[85]) );
  DFF \zreg_reg[86]  ( .D(o[86]), .CLK(clk), .RST(rst), .Q(zreg[86]) );
  DFF \zreg_reg[87]  ( .D(o[87]), .CLK(clk), .RST(rst), .Q(zreg[87]) );
  DFF \zreg_reg[88]  ( .D(o[88]), .CLK(clk), .RST(rst), .Q(zreg[88]) );
  DFF \zreg_reg[89]  ( .D(o[89]), .CLK(clk), .RST(rst), .Q(zreg[89]) );
  DFF \zreg_reg[90]  ( .D(o[90]), .CLK(clk), .RST(rst), .Q(zreg[90]) );
  DFF \zreg_reg[91]  ( .D(o[91]), .CLK(clk), .RST(rst), .Q(zreg[91]) );
  DFF \zreg_reg[92]  ( .D(o[92]), .CLK(clk), .RST(rst), .Q(zreg[92]) );
  DFF \zreg_reg[93]  ( .D(o[93]), .CLK(clk), .RST(rst), .Q(zreg[93]) );
  DFF \zreg_reg[94]  ( .D(o[94]), .CLK(clk), .RST(rst), .Q(zreg[94]) );
  DFF \zreg_reg[95]  ( .D(o[95]), .CLK(clk), .RST(rst), .Q(zreg[95]) );
  DFF \zreg_reg[96]  ( .D(o[96]), .CLK(clk), .RST(rst), .Q(zreg[96]) );
  DFF \zreg_reg[97]  ( .D(o[97]), .CLK(clk), .RST(rst), .Q(zreg[97]) );
  DFF \zreg_reg[98]  ( .D(o[98]), .CLK(clk), .RST(rst), .Q(zreg[98]) );
  DFF \zreg_reg[99]  ( .D(o[99]), .CLK(clk), .RST(rst), .Q(zreg[99]) );
  DFF \zreg_reg[100]  ( .D(o[100]), .CLK(clk), .RST(rst), .Q(zreg[100]) );
  DFF \zreg_reg[101]  ( .D(o[101]), .CLK(clk), .RST(rst), .Q(zreg[101]) );
  DFF \zreg_reg[102]  ( .D(o[102]), .CLK(clk), .RST(rst), .Q(zreg[102]) );
  DFF \zreg_reg[103]  ( .D(o[103]), .CLK(clk), .RST(rst), .Q(zreg[103]) );
  DFF \zreg_reg[104]  ( .D(o[104]), .CLK(clk), .RST(rst), .Q(zreg[104]) );
  DFF \zreg_reg[105]  ( .D(o[105]), .CLK(clk), .RST(rst), .Q(zreg[105]) );
  DFF \zreg_reg[106]  ( .D(o[106]), .CLK(clk), .RST(rst), .Q(zreg[106]) );
  DFF \zreg_reg[107]  ( .D(o[107]), .CLK(clk), .RST(rst), .Q(zreg[107]) );
  DFF \zreg_reg[108]  ( .D(o[108]), .CLK(clk), .RST(rst), .Q(zreg[108]) );
  DFF \zreg_reg[109]  ( .D(o[109]), .CLK(clk), .RST(rst), .Q(zreg[109]) );
  DFF \zreg_reg[110]  ( .D(o[110]), .CLK(clk), .RST(rst), .Q(zreg[110]) );
  DFF \zreg_reg[111]  ( .D(o[111]), .CLK(clk), .RST(rst), .Q(zreg[111]) );
  DFF \zreg_reg[112]  ( .D(o[112]), .CLK(clk), .RST(rst), .Q(zreg[112]) );
  DFF \zreg_reg[113]  ( .D(o[113]), .CLK(clk), .RST(rst), .Q(zreg[113]) );
  DFF \zreg_reg[114]  ( .D(o[114]), .CLK(clk), .RST(rst), .Q(zreg[114]) );
  DFF \zreg_reg[115]  ( .D(o[115]), .CLK(clk), .RST(rst), .Q(zreg[115]) );
  DFF \zreg_reg[116]  ( .D(o[116]), .CLK(clk), .RST(rst), .Q(zreg[116]) );
  DFF \zreg_reg[117]  ( .D(o[117]), .CLK(clk), .RST(rst), .Q(zreg[117]) );
  DFF \zreg_reg[118]  ( .D(o[118]), .CLK(clk), .RST(rst), .Q(zreg[118]) );
  DFF \zreg_reg[119]  ( .D(o[119]), .CLK(clk), .RST(rst), .Q(zreg[119]) );
  DFF \zreg_reg[120]  ( .D(o[120]), .CLK(clk), .RST(rst), .Q(zreg[120]) );
  DFF \zreg_reg[121]  ( .D(o[121]), .CLK(clk), .RST(rst), .Q(zreg[121]) );
  DFF \zreg_reg[122]  ( .D(o[122]), .CLK(clk), .RST(rst), .Q(zreg[122]) );
  DFF \zreg_reg[123]  ( .D(o[123]), .CLK(clk), .RST(rst), .Q(zreg[123]) );
  DFF \zreg_reg[124]  ( .D(o[124]), .CLK(clk), .RST(rst), .Q(zreg[124]) );
  DFF \zreg_reg[125]  ( .D(o[125]), .CLK(clk), .RST(rst), .Q(zreg[125]) );
  DFF \zreg_reg[126]  ( .D(o[126]), .CLK(clk), .RST(rst), .Q(zreg[126]) );
  DFF \zreg_reg[127]  ( .D(o[127]), .CLK(clk), .RST(rst), .Q(zreg[127]) );
  DFF \zreg_reg[128]  ( .D(o[128]), .CLK(clk), .RST(rst), .Q(zreg[128]) );
  DFF \zreg_reg[129]  ( .D(o[129]), .CLK(clk), .RST(rst), .Q(zreg[129]) );
  DFF \zreg_reg[130]  ( .D(o[130]), .CLK(clk), .RST(rst), .Q(zreg[130]) );
  DFF \zreg_reg[131]  ( .D(o[131]), .CLK(clk), .RST(rst), .Q(zreg[131]) );
  DFF \zreg_reg[132]  ( .D(o[132]), .CLK(clk), .RST(rst), .Q(zreg[132]) );
  DFF \zreg_reg[133]  ( .D(o[133]), .CLK(clk), .RST(rst), .Q(zreg[133]) );
  DFF \zreg_reg[134]  ( .D(o[134]), .CLK(clk), .RST(rst), .Q(zreg[134]) );
  DFF \zreg_reg[135]  ( .D(o[135]), .CLK(clk), .RST(rst), .Q(zreg[135]) );
  DFF \zreg_reg[136]  ( .D(o[136]), .CLK(clk), .RST(rst), .Q(zreg[136]) );
  DFF \zreg_reg[137]  ( .D(o[137]), .CLK(clk), .RST(rst), .Q(zreg[137]) );
  DFF \zreg_reg[138]  ( .D(o[138]), .CLK(clk), .RST(rst), .Q(zreg[138]) );
  DFF \zreg_reg[139]  ( .D(o[139]), .CLK(clk), .RST(rst), .Q(zreg[139]) );
  DFF \zreg_reg[140]  ( .D(o[140]), .CLK(clk), .RST(rst), .Q(zreg[140]) );
  DFF \zreg_reg[141]  ( .D(o[141]), .CLK(clk), .RST(rst), .Q(zreg[141]) );
  DFF \zreg_reg[142]  ( .D(o[142]), .CLK(clk), .RST(rst), .Q(zreg[142]) );
  DFF \zreg_reg[143]  ( .D(o[143]), .CLK(clk), .RST(rst), .Q(zreg[143]) );
  DFF \zreg_reg[144]  ( .D(o[144]), .CLK(clk), .RST(rst), .Q(zreg[144]) );
  DFF \zreg_reg[145]  ( .D(o[145]), .CLK(clk), .RST(rst), .Q(zreg[145]) );
  DFF \zreg_reg[146]  ( .D(o[146]), .CLK(clk), .RST(rst), .Q(zreg[146]) );
  DFF \zreg_reg[147]  ( .D(o[147]), .CLK(clk), .RST(rst), .Q(zreg[147]) );
  DFF \zreg_reg[148]  ( .D(o[148]), .CLK(clk), .RST(rst), .Q(zreg[148]) );
  DFF \zreg_reg[149]  ( .D(o[149]), .CLK(clk), .RST(rst), .Q(zreg[149]) );
  DFF \zreg_reg[150]  ( .D(o[150]), .CLK(clk), .RST(rst), .Q(zreg[150]) );
  DFF \zreg_reg[151]  ( .D(o[151]), .CLK(clk), .RST(rst), .Q(zreg[151]) );
  DFF \zreg_reg[152]  ( .D(o[152]), .CLK(clk), .RST(rst), .Q(zreg[152]) );
  DFF \zreg_reg[153]  ( .D(o[153]), .CLK(clk), .RST(rst), .Q(zreg[153]) );
  DFF \zreg_reg[154]  ( .D(o[154]), .CLK(clk), .RST(rst), .Q(zreg[154]) );
  DFF \zreg_reg[155]  ( .D(o[155]), .CLK(clk), .RST(rst), .Q(zreg[155]) );
  DFF \zreg_reg[156]  ( .D(o[156]), .CLK(clk), .RST(rst), .Q(zreg[156]) );
  DFF \zreg_reg[157]  ( .D(o[157]), .CLK(clk), .RST(rst), .Q(zreg[157]) );
  DFF \zreg_reg[158]  ( .D(o[158]), .CLK(clk), .RST(rst), .Q(zreg[158]) );
  DFF \zreg_reg[159]  ( .D(o[159]), .CLK(clk), .RST(rst), .Q(zreg[159]) );
  DFF \zreg_reg[160]  ( .D(o[160]), .CLK(clk), .RST(rst), .Q(zreg[160]) );
  DFF \zreg_reg[161]  ( .D(o[161]), .CLK(clk), .RST(rst), .Q(zreg[161]) );
  DFF \zreg_reg[162]  ( .D(o[162]), .CLK(clk), .RST(rst), .Q(zreg[162]) );
  DFF \zreg_reg[163]  ( .D(o[163]), .CLK(clk), .RST(rst), .Q(zreg[163]) );
  DFF \zreg_reg[164]  ( .D(o[164]), .CLK(clk), .RST(rst), .Q(zreg[164]) );
  DFF \zreg_reg[165]  ( .D(o[165]), .CLK(clk), .RST(rst), .Q(zreg[165]) );
  DFF \zreg_reg[166]  ( .D(o[166]), .CLK(clk), .RST(rst), .Q(zreg[166]) );
  DFF \zreg_reg[167]  ( .D(o[167]), .CLK(clk), .RST(rst), .Q(zreg[167]) );
  DFF \zreg_reg[168]  ( .D(o[168]), .CLK(clk), .RST(rst), .Q(zreg[168]) );
  DFF \zreg_reg[169]  ( .D(o[169]), .CLK(clk), .RST(rst), .Q(zreg[169]) );
  DFF \zreg_reg[170]  ( .D(o[170]), .CLK(clk), .RST(rst), .Q(zreg[170]) );
  DFF \zreg_reg[171]  ( .D(o[171]), .CLK(clk), .RST(rst), .Q(zreg[171]) );
  DFF \zreg_reg[172]  ( .D(o[172]), .CLK(clk), .RST(rst), .Q(zreg[172]) );
  DFF \zreg_reg[173]  ( .D(o[173]), .CLK(clk), .RST(rst), .Q(zreg[173]) );
  DFF \zreg_reg[174]  ( .D(o[174]), .CLK(clk), .RST(rst), .Q(zreg[174]) );
  DFF \zreg_reg[175]  ( .D(o[175]), .CLK(clk), .RST(rst), .Q(zreg[175]) );
  DFF \zreg_reg[176]  ( .D(o[176]), .CLK(clk), .RST(rst), .Q(zreg[176]) );
  DFF \zreg_reg[177]  ( .D(o[177]), .CLK(clk), .RST(rst), .Q(zreg[177]) );
  DFF \zreg_reg[178]  ( .D(o[178]), .CLK(clk), .RST(rst), .Q(zreg[178]) );
  DFF \zreg_reg[179]  ( .D(o[179]), .CLK(clk), .RST(rst), .Q(zreg[179]) );
  DFF \zreg_reg[180]  ( .D(o[180]), .CLK(clk), .RST(rst), .Q(zreg[180]) );
  DFF \zreg_reg[181]  ( .D(o[181]), .CLK(clk), .RST(rst), .Q(zreg[181]) );
  DFF \zreg_reg[182]  ( .D(o[182]), .CLK(clk), .RST(rst), .Q(zreg[182]) );
  DFF \zreg_reg[183]  ( .D(o[183]), .CLK(clk), .RST(rst), .Q(zreg[183]) );
  DFF \zreg_reg[184]  ( .D(o[184]), .CLK(clk), .RST(rst), .Q(zreg[184]) );
  DFF \zreg_reg[185]  ( .D(o[185]), .CLK(clk), .RST(rst), .Q(zreg[185]) );
  DFF \zreg_reg[186]  ( .D(o[186]), .CLK(clk), .RST(rst), .Q(zreg[186]) );
  DFF \zreg_reg[187]  ( .D(o[187]), .CLK(clk), .RST(rst), .Q(zreg[187]) );
  DFF \zreg_reg[188]  ( .D(o[188]), .CLK(clk), .RST(rst), .Q(zreg[188]) );
  DFF \zreg_reg[189]  ( .D(o[189]), .CLK(clk), .RST(rst), .Q(zreg[189]) );
  DFF \zreg_reg[190]  ( .D(o[190]), .CLK(clk), .RST(rst), .Q(zreg[190]) );
  DFF \zreg_reg[191]  ( .D(o[191]), .CLK(clk), .RST(rst), .Q(zreg[191]) );
  DFF \zreg_reg[192]  ( .D(o[192]), .CLK(clk), .RST(rst), .Q(zreg[192]) );
  DFF \zreg_reg[193]  ( .D(o[193]), .CLK(clk), .RST(rst), .Q(zreg[193]) );
  DFF \zreg_reg[194]  ( .D(o[194]), .CLK(clk), .RST(rst), .Q(zreg[194]) );
  DFF \zreg_reg[195]  ( .D(o[195]), .CLK(clk), .RST(rst), .Q(zreg[195]) );
  DFF \zreg_reg[196]  ( .D(o[196]), .CLK(clk), .RST(rst), .Q(zreg[196]) );
  DFF \zreg_reg[197]  ( .D(o[197]), .CLK(clk), .RST(rst), .Q(zreg[197]) );
  DFF \zreg_reg[198]  ( .D(o[198]), .CLK(clk), .RST(rst), .Q(zreg[198]) );
  DFF \zreg_reg[199]  ( .D(o[199]), .CLK(clk), .RST(rst), .Q(zreg[199]) );
  DFF \zreg_reg[200]  ( .D(o[200]), .CLK(clk), .RST(rst), .Q(zreg[200]) );
  DFF \zreg_reg[201]  ( .D(o[201]), .CLK(clk), .RST(rst), .Q(zreg[201]) );
  DFF \zreg_reg[202]  ( .D(o[202]), .CLK(clk), .RST(rst), .Q(zreg[202]) );
  DFF \zreg_reg[203]  ( .D(o[203]), .CLK(clk), .RST(rst), .Q(zreg[203]) );
  DFF \zreg_reg[204]  ( .D(o[204]), .CLK(clk), .RST(rst), .Q(zreg[204]) );
  DFF \zreg_reg[205]  ( .D(o[205]), .CLK(clk), .RST(rst), .Q(zreg[205]) );
  DFF \zreg_reg[206]  ( .D(o[206]), .CLK(clk), .RST(rst), .Q(zreg[206]) );
  DFF \zreg_reg[207]  ( .D(o[207]), .CLK(clk), .RST(rst), .Q(zreg[207]) );
  DFF \zreg_reg[208]  ( .D(o[208]), .CLK(clk), .RST(rst), .Q(zreg[208]) );
  DFF \zreg_reg[209]  ( .D(o[209]), .CLK(clk), .RST(rst), .Q(zreg[209]) );
  DFF \zreg_reg[210]  ( .D(o[210]), .CLK(clk), .RST(rst), .Q(zreg[210]) );
  DFF \zreg_reg[211]  ( .D(o[211]), .CLK(clk), .RST(rst), .Q(zreg[211]) );
  DFF \zreg_reg[212]  ( .D(o[212]), .CLK(clk), .RST(rst), .Q(zreg[212]) );
  DFF \zreg_reg[213]  ( .D(o[213]), .CLK(clk), .RST(rst), .Q(zreg[213]) );
  DFF \zreg_reg[214]  ( .D(o[214]), .CLK(clk), .RST(rst), .Q(zreg[214]) );
  DFF \zreg_reg[215]  ( .D(o[215]), .CLK(clk), .RST(rst), .Q(zreg[215]) );
  DFF \zreg_reg[216]  ( .D(o[216]), .CLK(clk), .RST(rst), .Q(zreg[216]) );
  DFF \zreg_reg[217]  ( .D(o[217]), .CLK(clk), .RST(rst), .Q(zreg[217]) );
  DFF \zreg_reg[218]  ( .D(o[218]), .CLK(clk), .RST(rst), .Q(zreg[218]) );
  DFF \zreg_reg[219]  ( .D(o[219]), .CLK(clk), .RST(rst), .Q(zreg[219]) );
  DFF \zreg_reg[220]  ( .D(o[220]), .CLK(clk), .RST(rst), .Q(zreg[220]) );
  DFF \zreg_reg[221]  ( .D(o[221]), .CLK(clk), .RST(rst), .Q(zreg[221]) );
  DFF \zreg_reg[222]  ( .D(o[222]), .CLK(clk), .RST(rst), .Q(zreg[222]) );
  DFF \zreg_reg[223]  ( .D(o[223]), .CLK(clk), .RST(rst), .Q(zreg[223]) );
  DFF \zreg_reg[224]  ( .D(o[224]), .CLK(clk), .RST(rst), .Q(zreg[224]) );
  DFF \zreg_reg[225]  ( .D(o[225]), .CLK(clk), .RST(rst), .Q(zreg[225]) );
  DFF \zreg_reg[226]  ( .D(o[226]), .CLK(clk), .RST(rst), .Q(zreg[226]) );
  DFF \zreg_reg[227]  ( .D(o[227]), .CLK(clk), .RST(rst), .Q(zreg[227]) );
  DFF \zreg_reg[228]  ( .D(o[228]), .CLK(clk), .RST(rst), .Q(zreg[228]) );
  DFF \zreg_reg[229]  ( .D(o[229]), .CLK(clk), .RST(rst), .Q(zreg[229]) );
  DFF \zreg_reg[230]  ( .D(o[230]), .CLK(clk), .RST(rst), .Q(zreg[230]) );
  DFF \zreg_reg[231]  ( .D(o[231]), .CLK(clk), .RST(rst), .Q(zreg[231]) );
  DFF \zreg_reg[232]  ( .D(o[232]), .CLK(clk), .RST(rst), .Q(zreg[232]) );
  DFF \zreg_reg[233]  ( .D(o[233]), .CLK(clk), .RST(rst), .Q(zreg[233]) );
  DFF \zreg_reg[234]  ( .D(o[234]), .CLK(clk), .RST(rst), .Q(zreg[234]) );
  DFF \zreg_reg[235]  ( .D(o[235]), .CLK(clk), .RST(rst), .Q(zreg[235]) );
  DFF \zreg_reg[236]  ( .D(o[236]), .CLK(clk), .RST(rst), .Q(zreg[236]) );
  DFF \zreg_reg[237]  ( .D(o[237]), .CLK(clk), .RST(rst), .Q(zreg[237]) );
  DFF \zreg_reg[238]  ( .D(o[238]), .CLK(clk), .RST(rst), .Q(zreg[238]) );
  DFF \zreg_reg[239]  ( .D(o[239]), .CLK(clk), .RST(rst), .Q(zreg[239]) );
  DFF \zreg_reg[240]  ( .D(o[240]), .CLK(clk), .RST(rst), .Q(zreg[240]) );
  DFF \zreg_reg[241]  ( .D(o[241]), .CLK(clk), .RST(rst), .Q(zreg[241]) );
  DFF \zreg_reg[242]  ( .D(o[242]), .CLK(clk), .RST(rst), .Q(zreg[242]) );
  DFF \zreg_reg[243]  ( .D(o[243]), .CLK(clk), .RST(rst), .Q(zreg[243]) );
  DFF \zreg_reg[244]  ( .D(o[244]), .CLK(clk), .RST(rst), .Q(zreg[244]) );
  DFF \zreg_reg[245]  ( .D(o[245]), .CLK(clk), .RST(rst), .Q(zreg[245]) );
  DFF \zreg_reg[246]  ( .D(o[246]), .CLK(clk), .RST(rst), .Q(zreg[246]) );
  DFF \zreg_reg[247]  ( .D(o[247]), .CLK(clk), .RST(rst), .Q(zreg[247]) );
  DFF \zreg_reg[248]  ( .D(o[248]), .CLK(clk), .RST(rst), .Q(zreg[248]) );
  DFF \zreg_reg[249]  ( .D(o[249]), .CLK(clk), .RST(rst), .Q(zreg[249]) );
  DFF \zreg_reg[250]  ( .D(o[250]), .CLK(clk), .RST(rst), .Q(zreg[250]) );
  DFF \zreg_reg[251]  ( .D(o[251]), .CLK(clk), .RST(rst), .Q(zreg[251]) );
  DFF \zreg_reg[252]  ( .D(o[252]), .CLK(clk), .RST(rst), .Q(zreg[252]) );
  DFF \zreg_reg[253]  ( .D(o[253]), .CLK(clk), .RST(rst), .Q(zreg[253]) );
  DFF \zreg_reg[254]  ( .D(o[254]), .CLK(clk), .RST(rst), .Q(zreg[254]) );
  DFF \zreg_reg[255]  ( .D(o[255]), .CLK(clk), .RST(rst), .Q(zreg[255]) );
  DFF \zreg_reg[256]  ( .D(o[256]), .CLK(clk), .RST(rst), .Q(zreg[256]) );
  DFF \zreg_reg[257]  ( .D(o[257]), .CLK(clk), .RST(rst), .Q(zreg[257]) );
  DFF \zreg_reg[258]  ( .D(o[258]), .CLK(clk), .RST(rst), .Q(zreg[258]) );
  DFF \zreg_reg[259]  ( .D(o[259]), .CLK(clk), .RST(rst), .Q(zreg[259]) );
  DFF \zreg_reg[260]  ( .D(o[260]), .CLK(clk), .RST(rst), .Q(zreg[260]) );
  DFF \zreg_reg[261]  ( .D(o[261]), .CLK(clk), .RST(rst), .Q(zreg[261]) );
  DFF \zreg_reg[262]  ( .D(o[262]), .CLK(clk), .RST(rst), .Q(zreg[262]) );
  DFF \zreg_reg[263]  ( .D(o[263]), .CLK(clk), .RST(rst), .Q(zreg[263]) );
  DFF \zreg_reg[264]  ( .D(o[264]), .CLK(clk), .RST(rst), .Q(zreg[264]) );
  DFF \zreg_reg[265]  ( .D(o[265]), .CLK(clk), .RST(rst), .Q(zreg[265]) );
  DFF \zreg_reg[266]  ( .D(o[266]), .CLK(clk), .RST(rst), .Q(zreg[266]) );
  DFF \zreg_reg[267]  ( .D(o[267]), .CLK(clk), .RST(rst), .Q(zreg[267]) );
  DFF \zreg_reg[268]  ( .D(o[268]), .CLK(clk), .RST(rst), .Q(zreg[268]) );
  DFF \zreg_reg[269]  ( .D(o[269]), .CLK(clk), .RST(rst), .Q(zreg[269]) );
  DFF \zreg_reg[270]  ( .D(o[270]), .CLK(clk), .RST(rst), .Q(zreg[270]) );
  DFF \zreg_reg[271]  ( .D(o[271]), .CLK(clk), .RST(rst), .Q(zreg[271]) );
  DFF \zreg_reg[272]  ( .D(o[272]), .CLK(clk), .RST(rst), .Q(zreg[272]) );
  DFF \zreg_reg[273]  ( .D(o[273]), .CLK(clk), .RST(rst), .Q(zreg[273]) );
  DFF \zreg_reg[274]  ( .D(o[274]), .CLK(clk), .RST(rst), .Q(zreg[274]) );
  DFF \zreg_reg[275]  ( .D(o[275]), .CLK(clk), .RST(rst), .Q(zreg[275]) );
  DFF \zreg_reg[276]  ( .D(o[276]), .CLK(clk), .RST(rst), .Q(zreg[276]) );
  DFF \zreg_reg[277]  ( .D(o[277]), .CLK(clk), .RST(rst), .Q(zreg[277]) );
  DFF \zreg_reg[278]  ( .D(o[278]), .CLK(clk), .RST(rst), .Q(zreg[278]) );
  DFF \zreg_reg[279]  ( .D(o[279]), .CLK(clk), .RST(rst), .Q(zreg[279]) );
  DFF \zreg_reg[280]  ( .D(o[280]), .CLK(clk), .RST(rst), .Q(zreg[280]) );
  DFF \zreg_reg[281]  ( .D(o[281]), .CLK(clk), .RST(rst), .Q(zreg[281]) );
  DFF \zreg_reg[282]  ( .D(o[282]), .CLK(clk), .RST(rst), .Q(zreg[282]) );
  DFF \zreg_reg[283]  ( .D(o[283]), .CLK(clk), .RST(rst), .Q(zreg[283]) );
  DFF \zreg_reg[284]  ( .D(o[284]), .CLK(clk), .RST(rst), .Q(zreg[284]) );
  DFF \zreg_reg[285]  ( .D(o[285]), .CLK(clk), .RST(rst), .Q(zreg[285]) );
  DFF \zreg_reg[286]  ( .D(o[286]), .CLK(clk), .RST(rst), .Q(zreg[286]) );
  DFF \zreg_reg[287]  ( .D(o[287]), .CLK(clk), .RST(rst), .Q(zreg[287]) );
  DFF \zreg_reg[288]  ( .D(o[288]), .CLK(clk), .RST(rst), .Q(zreg[288]) );
  DFF \zreg_reg[289]  ( .D(o[289]), .CLK(clk), .RST(rst), .Q(zreg[289]) );
  DFF \zreg_reg[290]  ( .D(o[290]), .CLK(clk), .RST(rst), .Q(zreg[290]) );
  DFF \zreg_reg[291]  ( .D(o[291]), .CLK(clk), .RST(rst), .Q(zreg[291]) );
  DFF \zreg_reg[292]  ( .D(o[292]), .CLK(clk), .RST(rst), .Q(zreg[292]) );
  DFF \zreg_reg[293]  ( .D(o[293]), .CLK(clk), .RST(rst), .Q(zreg[293]) );
  DFF \zreg_reg[294]  ( .D(o[294]), .CLK(clk), .RST(rst), .Q(zreg[294]) );
  DFF \zreg_reg[295]  ( .D(o[295]), .CLK(clk), .RST(rst), .Q(zreg[295]) );
  DFF \zreg_reg[296]  ( .D(o[296]), .CLK(clk), .RST(rst), .Q(zreg[296]) );
  DFF \zreg_reg[297]  ( .D(o[297]), .CLK(clk), .RST(rst), .Q(zreg[297]) );
  DFF \zreg_reg[298]  ( .D(o[298]), .CLK(clk), .RST(rst), .Q(zreg[298]) );
  DFF \zreg_reg[299]  ( .D(o[299]), .CLK(clk), .RST(rst), .Q(zreg[299]) );
  DFF \zreg_reg[300]  ( .D(o[300]), .CLK(clk), .RST(rst), .Q(zreg[300]) );
  DFF \zreg_reg[301]  ( .D(o[301]), .CLK(clk), .RST(rst), .Q(zreg[301]) );
  DFF \zreg_reg[302]  ( .D(o[302]), .CLK(clk), .RST(rst), .Q(zreg[302]) );
  DFF \zreg_reg[303]  ( .D(o[303]), .CLK(clk), .RST(rst), .Q(zreg[303]) );
  DFF \zreg_reg[304]  ( .D(o[304]), .CLK(clk), .RST(rst), .Q(zreg[304]) );
  DFF \zreg_reg[305]  ( .D(o[305]), .CLK(clk), .RST(rst), .Q(zreg[305]) );
  DFF \zreg_reg[306]  ( .D(o[306]), .CLK(clk), .RST(rst), .Q(zreg[306]) );
  DFF \zreg_reg[307]  ( .D(o[307]), .CLK(clk), .RST(rst), .Q(zreg[307]) );
  DFF \zreg_reg[308]  ( .D(o[308]), .CLK(clk), .RST(rst), .Q(zreg[308]) );
  DFF \zreg_reg[309]  ( .D(o[309]), .CLK(clk), .RST(rst), .Q(zreg[309]) );
  DFF \zreg_reg[310]  ( .D(o[310]), .CLK(clk), .RST(rst), .Q(zreg[310]) );
  DFF \zreg_reg[311]  ( .D(o[311]), .CLK(clk), .RST(rst), .Q(zreg[311]) );
  DFF \zreg_reg[312]  ( .D(o[312]), .CLK(clk), .RST(rst), .Q(zreg[312]) );
  DFF \zreg_reg[313]  ( .D(o[313]), .CLK(clk), .RST(rst), .Q(zreg[313]) );
  DFF \zreg_reg[314]  ( .D(o[314]), .CLK(clk), .RST(rst), .Q(zreg[314]) );
  DFF \zreg_reg[315]  ( .D(o[315]), .CLK(clk), .RST(rst), .Q(zreg[315]) );
  DFF \zreg_reg[316]  ( .D(o[316]), .CLK(clk), .RST(rst), .Q(zreg[316]) );
  DFF \zreg_reg[317]  ( .D(o[317]), .CLK(clk), .RST(rst), .Q(zreg[317]) );
  DFF \zreg_reg[318]  ( .D(o[318]), .CLK(clk), .RST(rst), .Q(zreg[318]) );
  DFF \zreg_reg[319]  ( .D(o[319]), .CLK(clk), .RST(rst), .Q(zreg[319]) );
  DFF \zreg_reg[320]  ( .D(o[320]), .CLK(clk), .RST(rst), .Q(zreg[320]) );
  DFF \zreg_reg[321]  ( .D(o[321]), .CLK(clk), .RST(rst), .Q(zreg[321]) );
  DFF \zreg_reg[322]  ( .D(o[322]), .CLK(clk), .RST(rst), .Q(zreg[322]) );
  DFF \zreg_reg[323]  ( .D(o[323]), .CLK(clk), .RST(rst), .Q(zreg[323]) );
  DFF \zreg_reg[324]  ( .D(o[324]), .CLK(clk), .RST(rst), .Q(zreg[324]) );
  DFF \zreg_reg[325]  ( .D(o[325]), .CLK(clk), .RST(rst), .Q(zreg[325]) );
  DFF \zreg_reg[326]  ( .D(o[326]), .CLK(clk), .RST(rst), .Q(zreg[326]) );
  DFF \zreg_reg[327]  ( .D(o[327]), .CLK(clk), .RST(rst), .Q(zreg[327]) );
  DFF \zreg_reg[328]  ( .D(o[328]), .CLK(clk), .RST(rst), .Q(zreg[328]) );
  DFF \zreg_reg[329]  ( .D(o[329]), .CLK(clk), .RST(rst), .Q(zreg[329]) );
  DFF \zreg_reg[330]  ( .D(o[330]), .CLK(clk), .RST(rst), .Q(zreg[330]) );
  DFF \zreg_reg[331]  ( .D(o[331]), .CLK(clk), .RST(rst), .Q(zreg[331]) );
  DFF \zreg_reg[332]  ( .D(o[332]), .CLK(clk), .RST(rst), .Q(zreg[332]) );
  DFF \zreg_reg[333]  ( .D(o[333]), .CLK(clk), .RST(rst), .Q(zreg[333]) );
  DFF \zreg_reg[334]  ( .D(o[334]), .CLK(clk), .RST(rst), .Q(zreg[334]) );
  DFF \zreg_reg[335]  ( .D(o[335]), .CLK(clk), .RST(rst), .Q(zreg[335]) );
  DFF \zreg_reg[336]  ( .D(o[336]), .CLK(clk), .RST(rst), .Q(zreg[336]) );
  DFF \zreg_reg[337]  ( .D(o[337]), .CLK(clk), .RST(rst), .Q(zreg[337]) );
  DFF \zreg_reg[338]  ( .D(o[338]), .CLK(clk), .RST(rst), .Q(zreg[338]) );
  DFF \zreg_reg[339]  ( .D(o[339]), .CLK(clk), .RST(rst), .Q(zreg[339]) );
  DFF \zreg_reg[340]  ( .D(o[340]), .CLK(clk), .RST(rst), .Q(zreg[340]) );
  DFF \zreg_reg[341]  ( .D(o[341]), .CLK(clk), .RST(rst), .Q(zreg[341]) );
  DFF \zreg_reg[342]  ( .D(o[342]), .CLK(clk), .RST(rst), .Q(zreg[342]) );
  DFF \zreg_reg[343]  ( .D(o[343]), .CLK(clk), .RST(rst), .Q(zreg[343]) );
  DFF \zreg_reg[344]  ( .D(o[344]), .CLK(clk), .RST(rst), .Q(zreg[344]) );
  DFF \zreg_reg[345]  ( .D(o[345]), .CLK(clk), .RST(rst), .Q(zreg[345]) );
  DFF \zreg_reg[346]  ( .D(o[346]), .CLK(clk), .RST(rst), .Q(zreg[346]) );
  DFF \zreg_reg[347]  ( .D(o[347]), .CLK(clk), .RST(rst), .Q(zreg[347]) );
  DFF \zreg_reg[348]  ( .D(o[348]), .CLK(clk), .RST(rst), .Q(zreg[348]) );
  DFF \zreg_reg[349]  ( .D(o[349]), .CLK(clk), .RST(rst), .Q(zreg[349]) );
  DFF \zreg_reg[350]  ( .D(o[350]), .CLK(clk), .RST(rst), .Q(zreg[350]) );
  DFF \zreg_reg[351]  ( .D(o[351]), .CLK(clk), .RST(rst), .Q(zreg[351]) );
  DFF \zreg_reg[352]  ( .D(o[352]), .CLK(clk), .RST(rst), .Q(zreg[352]) );
  DFF \zreg_reg[353]  ( .D(o[353]), .CLK(clk), .RST(rst), .Q(zreg[353]) );
  DFF \zreg_reg[354]  ( .D(o[354]), .CLK(clk), .RST(rst), .Q(zreg[354]) );
  DFF \zreg_reg[355]  ( .D(o[355]), .CLK(clk), .RST(rst), .Q(zreg[355]) );
  DFF \zreg_reg[356]  ( .D(o[356]), .CLK(clk), .RST(rst), .Q(zreg[356]) );
  DFF \zreg_reg[357]  ( .D(o[357]), .CLK(clk), .RST(rst), .Q(zreg[357]) );
  DFF \zreg_reg[358]  ( .D(o[358]), .CLK(clk), .RST(rst), .Q(zreg[358]) );
  DFF \zreg_reg[359]  ( .D(o[359]), .CLK(clk), .RST(rst), .Q(zreg[359]) );
  DFF \zreg_reg[360]  ( .D(o[360]), .CLK(clk), .RST(rst), .Q(zreg[360]) );
  DFF \zreg_reg[361]  ( .D(o[361]), .CLK(clk), .RST(rst), .Q(zreg[361]) );
  DFF \zreg_reg[362]  ( .D(o[362]), .CLK(clk), .RST(rst), .Q(zreg[362]) );
  DFF \zreg_reg[363]  ( .D(o[363]), .CLK(clk), .RST(rst), .Q(zreg[363]) );
  DFF \zreg_reg[364]  ( .D(o[364]), .CLK(clk), .RST(rst), .Q(zreg[364]) );
  DFF \zreg_reg[365]  ( .D(o[365]), .CLK(clk), .RST(rst), .Q(zreg[365]) );
  DFF \zreg_reg[366]  ( .D(o[366]), .CLK(clk), .RST(rst), .Q(zreg[366]) );
  DFF \zreg_reg[367]  ( .D(o[367]), .CLK(clk), .RST(rst), .Q(zreg[367]) );
  DFF \zreg_reg[368]  ( .D(o[368]), .CLK(clk), .RST(rst), .Q(zreg[368]) );
  DFF \zreg_reg[369]  ( .D(o[369]), .CLK(clk), .RST(rst), .Q(zreg[369]) );
  DFF \zreg_reg[370]  ( .D(o[370]), .CLK(clk), .RST(rst), .Q(zreg[370]) );
  DFF \zreg_reg[371]  ( .D(o[371]), .CLK(clk), .RST(rst), .Q(zreg[371]) );
  DFF \zreg_reg[372]  ( .D(o[372]), .CLK(clk), .RST(rst), .Q(zreg[372]) );
  DFF \zreg_reg[373]  ( .D(o[373]), .CLK(clk), .RST(rst), .Q(zreg[373]) );
  DFF \zreg_reg[374]  ( .D(o[374]), .CLK(clk), .RST(rst), .Q(zreg[374]) );
  DFF \zreg_reg[375]  ( .D(o[375]), .CLK(clk), .RST(rst), .Q(zreg[375]) );
  DFF \zreg_reg[376]  ( .D(o[376]), .CLK(clk), .RST(rst), .Q(zreg[376]) );
  DFF \zreg_reg[377]  ( .D(o[377]), .CLK(clk), .RST(rst), .Q(zreg[377]) );
  DFF \zreg_reg[378]  ( .D(o[378]), .CLK(clk), .RST(rst), .Q(zreg[378]) );
  DFF \zreg_reg[379]  ( .D(o[379]), .CLK(clk), .RST(rst), .Q(zreg[379]) );
  DFF \zreg_reg[380]  ( .D(o[380]), .CLK(clk), .RST(rst), .Q(zreg[380]) );
  DFF \zreg_reg[381]  ( .D(o[381]), .CLK(clk), .RST(rst), .Q(zreg[381]) );
  DFF \zreg_reg[382]  ( .D(o[382]), .CLK(clk), .RST(rst), .Q(zreg[382]) );
  DFF \zreg_reg[383]  ( .D(o[383]), .CLK(clk), .RST(rst), .Q(zreg[383]) );
  DFF \zreg_reg[384]  ( .D(o[384]), .CLK(clk), .RST(rst), .Q(zreg[384]) );
  DFF \zreg_reg[385]  ( .D(o[385]), .CLK(clk), .RST(rst), .Q(zreg[385]) );
  DFF \zreg_reg[386]  ( .D(o[386]), .CLK(clk), .RST(rst), .Q(zreg[386]) );
  DFF \zreg_reg[387]  ( .D(o[387]), .CLK(clk), .RST(rst), .Q(zreg[387]) );
  DFF \zreg_reg[388]  ( .D(o[388]), .CLK(clk), .RST(rst), .Q(zreg[388]) );
  DFF \zreg_reg[389]  ( .D(o[389]), .CLK(clk), .RST(rst), .Q(zreg[389]) );
  DFF \zreg_reg[390]  ( .D(o[390]), .CLK(clk), .RST(rst), .Q(zreg[390]) );
  DFF \zreg_reg[391]  ( .D(o[391]), .CLK(clk), .RST(rst), .Q(zreg[391]) );
  DFF \zreg_reg[392]  ( .D(o[392]), .CLK(clk), .RST(rst), .Q(zreg[392]) );
  DFF \zreg_reg[393]  ( .D(o[393]), .CLK(clk), .RST(rst), .Q(zreg[393]) );
  DFF \zreg_reg[394]  ( .D(o[394]), .CLK(clk), .RST(rst), .Q(zreg[394]) );
  DFF \zreg_reg[395]  ( .D(o[395]), .CLK(clk), .RST(rst), .Q(zreg[395]) );
  DFF \zreg_reg[396]  ( .D(o[396]), .CLK(clk), .RST(rst), .Q(zreg[396]) );
  DFF \zreg_reg[397]  ( .D(o[397]), .CLK(clk), .RST(rst), .Q(zreg[397]) );
  DFF \zreg_reg[398]  ( .D(o[398]), .CLK(clk), .RST(rst), .Q(zreg[398]) );
  DFF \zreg_reg[399]  ( .D(o[399]), .CLK(clk), .RST(rst), .Q(zreg[399]) );
  DFF \zreg_reg[400]  ( .D(o[400]), .CLK(clk), .RST(rst), .Q(zreg[400]) );
  DFF \zreg_reg[401]  ( .D(o[401]), .CLK(clk), .RST(rst), .Q(zreg[401]) );
  DFF \zreg_reg[402]  ( .D(o[402]), .CLK(clk), .RST(rst), .Q(zreg[402]) );
  DFF \zreg_reg[403]  ( .D(o[403]), .CLK(clk), .RST(rst), .Q(zreg[403]) );
  DFF \zreg_reg[404]  ( .D(o[404]), .CLK(clk), .RST(rst), .Q(zreg[404]) );
  DFF \zreg_reg[405]  ( .D(o[405]), .CLK(clk), .RST(rst), .Q(zreg[405]) );
  DFF \zreg_reg[406]  ( .D(o[406]), .CLK(clk), .RST(rst), .Q(zreg[406]) );
  DFF \zreg_reg[407]  ( .D(o[407]), .CLK(clk), .RST(rst), .Q(zreg[407]) );
  DFF \zreg_reg[408]  ( .D(o[408]), .CLK(clk), .RST(rst), .Q(zreg[408]) );
  DFF \zreg_reg[409]  ( .D(o[409]), .CLK(clk), .RST(rst), .Q(zreg[409]) );
  DFF \zreg_reg[410]  ( .D(o[410]), .CLK(clk), .RST(rst), .Q(zreg[410]) );
  DFF \zreg_reg[411]  ( .D(o[411]), .CLK(clk), .RST(rst), .Q(zreg[411]) );
  DFF \zreg_reg[412]  ( .D(o[412]), .CLK(clk), .RST(rst), .Q(zreg[412]) );
  DFF \zreg_reg[413]  ( .D(o[413]), .CLK(clk), .RST(rst), .Q(zreg[413]) );
  DFF \zreg_reg[414]  ( .D(o[414]), .CLK(clk), .RST(rst), .Q(zreg[414]) );
  DFF \zreg_reg[415]  ( .D(o[415]), .CLK(clk), .RST(rst), .Q(zreg[415]) );
  DFF \zreg_reg[416]  ( .D(o[416]), .CLK(clk), .RST(rst), .Q(zreg[416]) );
  DFF \zreg_reg[417]  ( .D(o[417]), .CLK(clk), .RST(rst), .Q(zreg[417]) );
  DFF \zreg_reg[418]  ( .D(o[418]), .CLK(clk), .RST(rst), .Q(zreg[418]) );
  DFF \zreg_reg[419]  ( .D(o[419]), .CLK(clk), .RST(rst), .Q(zreg[419]) );
  DFF \zreg_reg[420]  ( .D(o[420]), .CLK(clk), .RST(rst), .Q(zreg[420]) );
  DFF \zreg_reg[421]  ( .D(o[421]), .CLK(clk), .RST(rst), .Q(zreg[421]) );
  DFF \zreg_reg[422]  ( .D(o[422]), .CLK(clk), .RST(rst), .Q(zreg[422]) );
  DFF \zreg_reg[423]  ( .D(o[423]), .CLK(clk), .RST(rst), .Q(zreg[423]) );
  DFF \zreg_reg[424]  ( .D(o[424]), .CLK(clk), .RST(rst), .Q(zreg[424]) );
  DFF \zreg_reg[425]  ( .D(o[425]), .CLK(clk), .RST(rst), .Q(zreg[425]) );
  DFF \zreg_reg[426]  ( .D(o[426]), .CLK(clk), .RST(rst), .Q(zreg[426]) );
  DFF \zreg_reg[427]  ( .D(o[427]), .CLK(clk), .RST(rst), .Q(zreg[427]) );
  DFF \zreg_reg[428]  ( .D(o[428]), .CLK(clk), .RST(rst), .Q(zreg[428]) );
  DFF \zreg_reg[429]  ( .D(o[429]), .CLK(clk), .RST(rst), .Q(zreg[429]) );
  DFF \zreg_reg[430]  ( .D(o[430]), .CLK(clk), .RST(rst), .Q(zreg[430]) );
  DFF \zreg_reg[431]  ( .D(o[431]), .CLK(clk), .RST(rst), .Q(zreg[431]) );
  DFF \zreg_reg[432]  ( .D(o[432]), .CLK(clk), .RST(rst), .Q(zreg[432]) );
  DFF \zreg_reg[433]  ( .D(o[433]), .CLK(clk), .RST(rst), .Q(zreg[433]) );
  DFF \zreg_reg[434]  ( .D(o[434]), .CLK(clk), .RST(rst), .Q(zreg[434]) );
  DFF \zreg_reg[435]  ( .D(o[435]), .CLK(clk), .RST(rst), .Q(zreg[435]) );
  DFF \zreg_reg[436]  ( .D(o[436]), .CLK(clk), .RST(rst), .Q(zreg[436]) );
  DFF \zreg_reg[437]  ( .D(o[437]), .CLK(clk), .RST(rst), .Q(zreg[437]) );
  DFF \zreg_reg[438]  ( .D(o[438]), .CLK(clk), .RST(rst), .Q(zreg[438]) );
  DFF \zreg_reg[439]  ( .D(o[439]), .CLK(clk), .RST(rst), .Q(zreg[439]) );
  DFF \zreg_reg[440]  ( .D(o[440]), .CLK(clk), .RST(rst), .Q(zreg[440]) );
  DFF \zreg_reg[441]  ( .D(o[441]), .CLK(clk), .RST(rst), .Q(zreg[441]) );
  DFF \zreg_reg[442]  ( .D(o[442]), .CLK(clk), .RST(rst), .Q(zreg[442]) );
  DFF \zreg_reg[443]  ( .D(o[443]), .CLK(clk), .RST(rst), .Q(zreg[443]) );
  DFF \zreg_reg[444]  ( .D(o[444]), .CLK(clk), .RST(rst), .Q(zreg[444]) );
  DFF \zreg_reg[445]  ( .D(o[445]), .CLK(clk), .RST(rst), .Q(zreg[445]) );
  DFF \zreg_reg[446]  ( .D(o[446]), .CLK(clk), .RST(rst), .Q(zreg[446]) );
  DFF \zreg_reg[447]  ( .D(o[447]), .CLK(clk), .RST(rst), .Q(zreg[447]) );
  DFF \zreg_reg[448]  ( .D(o[448]), .CLK(clk), .RST(rst), .Q(zreg[448]) );
  DFF \zreg_reg[449]  ( .D(o[449]), .CLK(clk), .RST(rst), .Q(zreg[449]) );
  DFF \zreg_reg[450]  ( .D(o[450]), .CLK(clk), .RST(rst), .Q(zreg[450]) );
  DFF \zreg_reg[451]  ( .D(o[451]), .CLK(clk), .RST(rst), .Q(zreg[451]) );
  DFF \zreg_reg[452]  ( .D(o[452]), .CLK(clk), .RST(rst), .Q(zreg[452]) );
  DFF \zreg_reg[453]  ( .D(o[453]), .CLK(clk), .RST(rst), .Q(zreg[453]) );
  DFF \zreg_reg[454]  ( .D(o[454]), .CLK(clk), .RST(rst), .Q(zreg[454]) );
  DFF \zreg_reg[455]  ( .D(o[455]), .CLK(clk), .RST(rst), .Q(zreg[455]) );
  DFF \zreg_reg[456]  ( .D(o[456]), .CLK(clk), .RST(rst), .Q(zreg[456]) );
  DFF \zreg_reg[457]  ( .D(o[457]), .CLK(clk), .RST(rst), .Q(zreg[457]) );
  DFF \zreg_reg[458]  ( .D(o[458]), .CLK(clk), .RST(rst), .Q(zreg[458]) );
  DFF \zreg_reg[459]  ( .D(o[459]), .CLK(clk), .RST(rst), .Q(zreg[459]) );
  DFF \zreg_reg[460]  ( .D(o[460]), .CLK(clk), .RST(rst), .Q(zreg[460]) );
  DFF \zreg_reg[461]  ( .D(o[461]), .CLK(clk), .RST(rst), .Q(zreg[461]) );
  DFF \zreg_reg[462]  ( .D(o[462]), .CLK(clk), .RST(rst), .Q(zreg[462]) );
  DFF \zreg_reg[463]  ( .D(o[463]), .CLK(clk), .RST(rst), .Q(zreg[463]) );
  DFF \zreg_reg[464]  ( .D(o[464]), .CLK(clk), .RST(rst), .Q(zreg[464]) );
  DFF \zreg_reg[465]  ( .D(o[465]), .CLK(clk), .RST(rst), .Q(zreg[465]) );
  DFF \zreg_reg[466]  ( .D(o[466]), .CLK(clk), .RST(rst), .Q(zreg[466]) );
  DFF \zreg_reg[467]  ( .D(o[467]), .CLK(clk), .RST(rst), .Q(zreg[467]) );
  DFF \zreg_reg[468]  ( .D(o[468]), .CLK(clk), .RST(rst), .Q(zreg[468]) );
  DFF \zreg_reg[469]  ( .D(o[469]), .CLK(clk), .RST(rst), .Q(zreg[469]) );
  DFF \zreg_reg[470]  ( .D(o[470]), .CLK(clk), .RST(rst), .Q(zreg[470]) );
  DFF \zreg_reg[471]  ( .D(o[471]), .CLK(clk), .RST(rst), .Q(zreg[471]) );
  DFF \zreg_reg[472]  ( .D(o[472]), .CLK(clk), .RST(rst), .Q(zreg[472]) );
  DFF \zreg_reg[473]  ( .D(o[473]), .CLK(clk), .RST(rst), .Q(zreg[473]) );
  DFF \zreg_reg[474]  ( .D(o[474]), .CLK(clk), .RST(rst), .Q(zreg[474]) );
  DFF \zreg_reg[475]  ( .D(o[475]), .CLK(clk), .RST(rst), .Q(zreg[475]) );
  DFF \zreg_reg[476]  ( .D(o[476]), .CLK(clk), .RST(rst), .Q(zreg[476]) );
  DFF \zreg_reg[477]  ( .D(o[477]), .CLK(clk), .RST(rst), .Q(zreg[477]) );
  DFF \zreg_reg[478]  ( .D(o[478]), .CLK(clk), .RST(rst), .Q(zreg[478]) );
  DFF \zreg_reg[479]  ( .D(o[479]), .CLK(clk), .RST(rst), .Q(zreg[479]) );
  DFF \zreg_reg[480]  ( .D(o[480]), .CLK(clk), .RST(rst), .Q(zreg[480]) );
  DFF \zreg_reg[481]  ( .D(o[481]), .CLK(clk), .RST(rst), .Q(zreg[481]) );
  DFF \zreg_reg[482]  ( .D(o[482]), .CLK(clk), .RST(rst), .Q(zreg[482]) );
  DFF \zreg_reg[483]  ( .D(o[483]), .CLK(clk), .RST(rst), .Q(zreg[483]) );
  DFF \zreg_reg[484]  ( .D(o[484]), .CLK(clk), .RST(rst), .Q(zreg[484]) );
  DFF \zreg_reg[485]  ( .D(o[485]), .CLK(clk), .RST(rst), .Q(zreg[485]) );
  DFF \zreg_reg[486]  ( .D(o[486]), .CLK(clk), .RST(rst), .Q(zreg[486]) );
  DFF \zreg_reg[487]  ( .D(o[487]), .CLK(clk), .RST(rst), .Q(zreg[487]) );
  DFF \zreg_reg[488]  ( .D(o[488]), .CLK(clk), .RST(rst), .Q(zreg[488]) );
  DFF \zreg_reg[489]  ( .D(o[489]), .CLK(clk), .RST(rst), .Q(zreg[489]) );
  DFF \zreg_reg[490]  ( .D(o[490]), .CLK(clk), .RST(rst), .Q(zreg[490]) );
  DFF \zreg_reg[491]  ( .D(o[491]), .CLK(clk), .RST(rst), .Q(zreg[491]) );
  DFF \zreg_reg[492]  ( .D(o[492]), .CLK(clk), .RST(rst), .Q(zreg[492]) );
  DFF \zreg_reg[493]  ( .D(o[493]), .CLK(clk), .RST(rst), .Q(zreg[493]) );
  DFF \zreg_reg[494]  ( .D(o[494]), .CLK(clk), .RST(rst), .Q(zreg[494]) );
  DFF \zreg_reg[495]  ( .D(o[495]), .CLK(clk), .RST(rst), .Q(zreg[495]) );
  DFF \zreg_reg[496]  ( .D(o[496]), .CLK(clk), .RST(rst), .Q(zreg[496]) );
  DFF \zreg_reg[497]  ( .D(o[497]), .CLK(clk), .RST(rst), .Q(zreg[497]) );
  DFF \zreg_reg[498]  ( .D(o[498]), .CLK(clk), .RST(rst), .Q(zreg[498]) );
  DFF \zreg_reg[499]  ( .D(o[499]), .CLK(clk), .RST(rst), .Q(zreg[499]) );
  DFF \zreg_reg[500]  ( .D(o[500]), .CLK(clk), .RST(rst), .Q(zreg[500]) );
  DFF \zreg_reg[501]  ( .D(o[501]), .CLK(clk), .RST(rst), .Q(zreg[501]) );
  DFF \zreg_reg[502]  ( .D(o[502]), .CLK(clk), .RST(rst), .Q(zreg[502]) );
  DFF \zreg_reg[503]  ( .D(o[503]), .CLK(clk), .RST(rst), .Q(zreg[503]) );
  DFF \zreg_reg[504]  ( .D(o[504]), .CLK(clk), .RST(rst), .Q(zreg[504]) );
  DFF \zreg_reg[505]  ( .D(o[505]), .CLK(clk), .RST(rst), .Q(zreg[505]) );
  DFF \zreg_reg[506]  ( .D(o[506]), .CLK(clk), .RST(rst), .Q(zreg[506]) );
  DFF \zreg_reg[507]  ( .D(o[507]), .CLK(clk), .RST(rst), .Q(zreg[507]) );
  DFF \zreg_reg[508]  ( .D(o[508]), .CLK(clk), .RST(rst), .Q(zreg[508]) );
  DFF \zreg_reg[509]  ( .D(o[509]), .CLK(clk), .RST(rst), .Q(zreg[509]) );
  DFF \zreg_reg[510]  ( .D(o[510]), .CLK(clk), .RST(rst), .Q(zreg[510]) );
  DFF \zreg_reg[511]  ( .D(o[511]), .CLK(clk), .RST(rst), .Q(zreg[511]) );
  DFF \zreg_reg[512]  ( .D(o[512]), .CLK(clk), .RST(rst), .Q(zreg[512]) );
  DFF \zreg_reg[513]  ( .D(o[513]), .CLK(clk), .RST(rst), .Q(zreg[513]) );
  DFF \zreg_reg[514]  ( .D(o[514]), .CLK(clk), .RST(rst), .Q(zreg[514]) );
  DFF \zreg_reg[515]  ( .D(o[515]), .CLK(clk), .RST(rst), .Q(zreg[515]) );
  DFF \zreg_reg[516]  ( .D(o[516]), .CLK(clk), .RST(rst), .Q(zreg[516]) );
  DFF \zreg_reg[517]  ( .D(o[517]), .CLK(clk), .RST(rst), .Q(zreg[517]) );
  DFF \zreg_reg[518]  ( .D(o[518]), .CLK(clk), .RST(rst), .Q(zreg[518]) );
  DFF \zreg_reg[519]  ( .D(o[519]), .CLK(clk), .RST(rst), .Q(zreg[519]) );
  DFF \zreg_reg[520]  ( .D(o[520]), .CLK(clk), .RST(rst), .Q(zreg[520]) );
  DFF \zreg_reg[521]  ( .D(o[521]), .CLK(clk), .RST(rst), .Q(zreg[521]) );
  DFF \zreg_reg[522]  ( .D(o[522]), .CLK(clk), .RST(rst), .Q(zreg[522]) );
  DFF \zreg_reg[523]  ( .D(o[523]), .CLK(clk), .RST(rst), .Q(zreg[523]) );
  DFF \zreg_reg[524]  ( .D(o[524]), .CLK(clk), .RST(rst), .Q(zreg[524]) );
  DFF \zreg_reg[525]  ( .D(o[525]), .CLK(clk), .RST(rst), .Q(zreg[525]) );
  DFF \zreg_reg[526]  ( .D(o[526]), .CLK(clk), .RST(rst), .Q(zreg[526]) );
  DFF \zreg_reg[527]  ( .D(o[527]), .CLK(clk), .RST(rst), .Q(zreg[527]) );
  DFF \zreg_reg[528]  ( .D(o[528]), .CLK(clk), .RST(rst), .Q(zreg[528]) );
  DFF \zreg_reg[529]  ( .D(o[529]), .CLK(clk), .RST(rst), .Q(zreg[529]) );
  DFF \zreg_reg[530]  ( .D(o[530]), .CLK(clk), .RST(rst), .Q(zreg[530]) );
  DFF \zreg_reg[531]  ( .D(o[531]), .CLK(clk), .RST(rst), .Q(zreg[531]) );
  DFF \zreg_reg[532]  ( .D(o[532]), .CLK(clk), .RST(rst), .Q(zreg[532]) );
  DFF \zreg_reg[533]  ( .D(o[533]), .CLK(clk), .RST(rst), .Q(zreg[533]) );
  DFF \zreg_reg[534]  ( .D(o[534]), .CLK(clk), .RST(rst), .Q(zreg[534]) );
  DFF \zreg_reg[535]  ( .D(o[535]), .CLK(clk), .RST(rst), .Q(zreg[535]) );
  DFF \zreg_reg[536]  ( .D(o[536]), .CLK(clk), .RST(rst), .Q(zreg[536]) );
  DFF \zreg_reg[537]  ( .D(o[537]), .CLK(clk), .RST(rst), .Q(zreg[537]) );
  DFF \zreg_reg[538]  ( .D(o[538]), .CLK(clk), .RST(rst), .Q(zreg[538]) );
  DFF \zreg_reg[539]  ( .D(o[539]), .CLK(clk), .RST(rst), .Q(zreg[539]) );
  DFF \zreg_reg[540]  ( .D(o[540]), .CLK(clk), .RST(rst), .Q(zreg[540]) );
  DFF \zreg_reg[541]  ( .D(o[541]), .CLK(clk), .RST(rst), .Q(zreg[541]) );
  DFF \zreg_reg[542]  ( .D(o[542]), .CLK(clk), .RST(rst), .Q(zreg[542]) );
  DFF \zreg_reg[543]  ( .D(o[543]), .CLK(clk), .RST(rst), .Q(zreg[543]) );
  DFF \zreg_reg[544]  ( .D(o[544]), .CLK(clk), .RST(rst), .Q(zreg[544]) );
  DFF \zreg_reg[545]  ( .D(o[545]), .CLK(clk), .RST(rst), .Q(zreg[545]) );
  DFF \zreg_reg[546]  ( .D(o[546]), .CLK(clk), .RST(rst), .Q(zreg[546]) );
  DFF \zreg_reg[547]  ( .D(o[547]), .CLK(clk), .RST(rst), .Q(zreg[547]) );
  DFF \zreg_reg[548]  ( .D(o[548]), .CLK(clk), .RST(rst), .Q(zreg[548]) );
  DFF \zreg_reg[549]  ( .D(o[549]), .CLK(clk), .RST(rst), .Q(zreg[549]) );
  DFF \zreg_reg[550]  ( .D(o[550]), .CLK(clk), .RST(rst), .Q(zreg[550]) );
  DFF \zreg_reg[551]  ( .D(o[551]), .CLK(clk), .RST(rst), .Q(zreg[551]) );
  DFF \zreg_reg[552]  ( .D(o[552]), .CLK(clk), .RST(rst), .Q(zreg[552]) );
  DFF \zreg_reg[553]  ( .D(o[553]), .CLK(clk), .RST(rst), .Q(zreg[553]) );
  DFF \zreg_reg[554]  ( .D(o[554]), .CLK(clk), .RST(rst), .Q(zreg[554]) );
  DFF \zreg_reg[555]  ( .D(o[555]), .CLK(clk), .RST(rst), .Q(zreg[555]) );
  DFF \zreg_reg[556]  ( .D(o[556]), .CLK(clk), .RST(rst), .Q(zreg[556]) );
  DFF \zreg_reg[557]  ( .D(o[557]), .CLK(clk), .RST(rst), .Q(zreg[557]) );
  DFF \zreg_reg[558]  ( .D(o[558]), .CLK(clk), .RST(rst), .Q(zreg[558]) );
  DFF \zreg_reg[559]  ( .D(o[559]), .CLK(clk), .RST(rst), .Q(zreg[559]) );
  DFF \zreg_reg[560]  ( .D(o[560]), .CLK(clk), .RST(rst), .Q(zreg[560]) );
  DFF \zreg_reg[561]  ( .D(o[561]), .CLK(clk), .RST(rst), .Q(zreg[561]) );
  DFF \zreg_reg[562]  ( .D(o[562]), .CLK(clk), .RST(rst), .Q(zreg[562]) );
  DFF \zreg_reg[563]  ( .D(o[563]), .CLK(clk), .RST(rst), .Q(zreg[563]) );
  DFF \zreg_reg[564]  ( .D(o[564]), .CLK(clk), .RST(rst), .Q(zreg[564]) );
  DFF \zreg_reg[565]  ( .D(o[565]), .CLK(clk), .RST(rst), .Q(zreg[565]) );
  DFF \zreg_reg[566]  ( .D(o[566]), .CLK(clk), .RST(rst), .Q(zreg[566]) );
  DFF \zreg_reg[567]  ( .D(o[567]), .CLK(clk), .RST(rst), .Q(zreg[567]) );
  DFF \zreg_reg[568]  ( .D(o[568]), .CLK(clk), .RST(rst), .Q(zreg[568]) );
  DFF \zreg_reg[569]  ( .D(o[569]), .CLK(clk), .RST(rst), .Q(zreg[569]) );
  DFF \zreg_reg[570]  ( .D(o[570]), .CLK(clk), .RST(rst), .Q(zreg[570]) );
  DFF \zreg_reg[571]  ( .D(o[571]), .CLK(clk), .RST(rst), .Q(zreg[571]) );
  DFF \zreg_reg[572]  ( .D(o[572]), .CLK(clk), .RST(rst), .Q(zreg[572]) );
  DFF \zreg_reg[573]  ( .D(o[573]), .CLK(clk), .RST(rst), .Q(zreg[573]) );
  DFF \zreg_reg[574]  ( .D(o[574]), .CLK(clk), .RST(rst), .Q(zreg[574]) );
  DFF \zreg_reg[575]  ( .D(o[575]), .CLK(clk), .RST(rst), .Q(zreg[575]) );
  DFF \zreg_reg[576]  ( .D(o[576]), .CLK(clk), .RST(rst), .Q(zreg[576]) );
  DFF \zreg_reg[577]  ( .D(o[577]), .CLK(clk), .RST(rst), .Q(zreg[577]) );
  DFF \zreg_reg[578]  ( .D(o[578]), .CLK(clk), .RST(rst), .Q(zreg[578]) );
  DFF \zreg_reg[579]  ( .D(o[579]), .CLK(clk), .RST(rst), .Q(zreg[579]) );
  DFF \zreg_reg[580]  ( .D(o[580]), .CLK(clk), .RST(rst), .Q(zreg[580]) );
  DFF \zreg_reg[581]  ( .D(o[581]), .CLK(clk), .RST(rst), .Q(zreg[581]) );
  DFF \zreg_reg[582]  ( .D(o[582]), .CLK(clk), .RST(rst), .Q(zreg[582]) );
  DFF \zreg_reg[583]  ( .D(o[583]), .CLK(clk), .RST(rst), .Q(zreg[583]) );
  DFF \zreg_reg[584]  ( .D(o[584]), .CLK(clk), .RST(rst), .Q(zreg[584]) );
  DFF \zreg_reg[585]  ( .D(o[585]), .CLK(clk), .RST(rst), .Q(zreg[585]) );
  DFF \zreg_reg[586]  ( .D(o[586]), .CLK(clk), .RST(rst), .Q(zreg[586]) );
  DFF \zreg_reg[587]  ( .D(o[587]), .CLK(clk), .RST(rst), .Q(zreg[587]) );
  DFF \zreg_reg[588]  ( .D(o[588]), .CLK(clk), .RST(rst), .Q(zreg[588]) );
  DFF \zreg_reg[589]  ( .D(o[589]), .CLK(clk), .RST(rst), .Q(zreg[589]) );
  DFF \zreg_reg[590]  ( .D(o[590]), .CLK(clk), .RST(rst), .Q(zreg[590]) );
  DFF \zreg_reg[591]  ( .D(o[591]), .CLK(clk), .RST(rst), .Q(zreg[591]) );
  DFF \zreg_reg[592]  ( .D(o[592]), .CLK(clk), .RST(rst), .Q(zreg[592]) );
  DFF \zreg_reg[593]  ( .D(o[593]), .CLK(clk), .RST(rst), .Q(zreg[593]) );
  DFF \zreg_reg[594]  ( .D(o[594]), .CLK(clk), .RST(rst), .Q(zreg[594]) );
  DFF \zreg_reg[595]  ( .D(o[595]), .CLK(clk), .RST(rst), .Q(zreg[595]) );
  DFF \zreg_reg[596]  ( .D(o[596]), .CLK(clk), .RST(rst), .Q(zreg[596]) );
  DFF \zreg_reg[597]  ( .D(o[597]), .CLK(clk), .RST(rst), .Q(zreg[597]) );
  DFF \zreg_reg[598]  ( .D(o[598]), .CLK(clk), .RST(rst), .Q(zreg[598]) );
  DFF \zreg_reg[599]  ( .D(o[599]), .CLK(clk), .RST(rst), .Q(zreg[599]) );
  DFF \zreg_reg[600]  ( .D(o[600]), .CLK(clk), .RST(rst), .Q(zreg[600]) );
  DFF \zreg_reg[601]  ( .D(o[601]), .CLK(clk), .RST(rst), .Q(zreg[601]) );
  DFF \zreg_reg[602]  ( .D(o[602]), .CLK(clk), .RST(rst), .Q(zreg[602]) );
  DFF \zreg_reg[603]  ( .D(o[603]), .CLK(clk), .RST(rst), .Q(zreg[603]) );
  DFF \zreg_reg[604]  ( .D(o[604]), .CLK(clk), .RST(rst), .Q(zreg[604]) );
  DFF \zreg_reg[605]  ( .D(o[605]), .CLK(clk), .RST(rst), .Q(zreg[605]) );
  DFF \zreg_reg[606]  ( .D(o[606]), .CLK(clk), .RST(rst), .Q(zreg[606]) );
  DFF \zreg_reg[607]  ( .D(o[607]), .CLK(clk), .RST(rst), .Q(zreg[607]) );
  DFF \zreg_reg[608]  ( .D(o[608]), .CLK(clk), .RST(rst), .Q(zreg[608]) );
  DFF \zreg_reg[609]  ( .D(o[609]), .CLK(clk), .RST(rst), .Q(zreg[609]) );
  DFF \zreg_reg[610]  ( .D(o[610]), .CLK(clk), .RST(rst), .Q(zreg[610]) );
  DFF \zreg_reg[611]  ( .D(o[611]), .CLK(clk), .RST(rst), .Q(zreg[611]) );
  DFF \zreg_reg[612]  ( .D(o[612]), .CLK(clk), .RST(rst), .Q(zreg[612]) );
  DFF \zreg_reg[613]  ( .D(o[613]), .CLK(clk), .RST(rst), .Q(zreg[613]) );
  DFF \zreg_reg[614]  ( .D(o[614]), .CLK(clk), .RST(rst), .Q(zreg[614]) );
  DFF \zreg_reg[615]  ( .D(o[615]), .CLK(clk), .RST(rst), .Q(zreg[615]) );
  DFF \zreg_reg[616]  ( .D(o[616]), .CLK(clk), .RST(rst), .Q(zreg[616]) );
  DFF \zreg_reg[617]  ( .D(o[617]), .CLK(clk), .RST(rst), .Q(zreg[617]) );
  DFF \zreg_reg[618]  ( .D(o[618]), .CLK(clk), .RST(rst), .Q(zreg[618]) );
  DFF \zreg_reg[619]  ( .D(o[619]), .CLK(clk), .RST(rst), .Q(zreg[619]) );
  DFF \zreg_reg[620]  ( .D(o[620]), .CLK(clk), .RST(rst), .Q(zreg[620]) );
  DFF \zreg_reg[621]  ( .D(o[621]), .CLK(clk), .RST(rst), .Q(zreg[621]) );
  DFF \zreg_reg[622]  ( .D(o[622]), .CLK(clk), .RST(rst), .Q(zreg[622]) );
  DFF \zreg_reg[623]  ( .D(o[623]), .CLK(clk), .RST(rst), .Q(zreg[623]) );
  DFF \zreg_reg[624]  ( .D(o[624]), .CLK(clk), .RST(rst), .Q(zreg[624]) );
  DFF \zreg_reg[625]  ( .D(o[625]), .CLK(clk), .RST(rst), .Q(zreg[625]) );
  DFF \zreg_reg[626]  ( .D(o[626]), .CLK(clk), .RST(rst), .Q(zreg[626]) );
  DFF \zreg_reg[627]  ( .D(o[627]), .CLK(clk), .RST(rst), .Q(zreg[627]) );
  DFF \zreg_reg[628]  ( .D(o[628]), .CLK(clk), .RST(rst), .Q(zreg[628]) );
  DFF \zreg_reg[629]  ( .D(o[629]), .CLK(clk), .RST(rst), .Q(zreg[629]) );
  DFF \zreg_reg[630]  ( .D(o[630]), .CLK(clk), .RST(rst), .Q(zreg[630]) );
  DFF \zreg_reg[631]  ( .D(o[631]), .CLK(clk), .RST(rst), .Q(zreg[631]) );
  DFF \zreg_reg[632]  ( .D(o[632]), .CLK(clk), .RST(rst), .Q(zreg[632]) );
  DFF \zreg_reg[633]  ( .D(o[633]), .CLK(clk), .RST(rst), .Q(zreg[633]) );
  DFF \zreg_reg[634]  ( .D(o[634]), .CLK(clk), .RST(rst), .Q(zreg[634]) );
  DFF \zreg_reg[635]  ( .D(o[635]), .CLK(clk), .RST(rst), .Q(zreg[635]) );
  DFF \zreg_reg[636]  ( .D(o[636]), .CLK(clk), .RST(rst), .Q(zreg[636]) );
  DFF \zreg_reg[637]  ( .D(o[637]), .CLK(clk), .RST(rst), .Q(zreg[637]) );
  DFF \zreg_reg[638]  ( .D(o[638]), .CLK(clk), .RST(rst), .Q(zreg[638]) );
  DFF \zreg_reg[639]  ( .D(o[639]), .CLK(clk), .RST(rst), .Q(zreg[639]) );
  DFF \zreg_reg[640]  ( .D(o[640]), .CLK(clk), .RST(rst), .Q(zreg[640]) );
  DFF \zreg_reg[641]  ( .D(o[641]), .CLK(clk), .RST(rst), .Q(zreg[641]) );
  DFF \zreg_reg[642]  ( .D(o[642]), .CLK(clk), .RST(rst), .Q(zreg[642]) );
  DFF \zreg_reg[643]  ( .D(o[643]), .CLK(clk), .RST(rst), .Q(zreg[643]) );
  DFF \zreg_reg[644]  ( .D(o[644]), .CLK(clk), .RST(rst), .Q(zreg[644]) );
  DFF \zreg_reg[645]  ( .D(o[645]), .CLK(clk), .RST(rst), .Q(zreg[645]) );
  DFF \zreg_reg[646]  ( .D(o[646]), .CLK(clk), .RST(rst), .Q(zreg[646]) );
  DFF \zreg_reg[647]  ( .D(o[647]), .CLK(clk), .RST(rst), .Q(zreg[647]) );
  DFF \zreg_reg[648]  ( .D(o[648]), .CLK(clk), .RST(rst), .Q(zreg[648]) );
  DFF \zreg_reg[649]  ( .D(o[649]), .CLK(clk), .RST(rst), .Q(zreg[649]) );
  DFF \zreg_reg[650]  ( .D(o[650]), .CLK(clk), .RST(rst), .Q(zreg[650]) );
  DFF \zreg_reg[651]  ( .D(o[651]), .CLK(clk), .RST(rst), .Q(zreg[651]) );
  DFF \zreg_reg[652]  ( .D(o[652]), .CLK(clk), .RST(rst), .Q(zreg[652]) );
  DFF \zreg_reg[653]  ( .D(o[653]), .CLK(clk), .RST(rst), .Q(zreg[653]) );
  DFF \zreg_reg[654]  ( .D(o[654]), .CLK(clk), .RST(rst), .Q(zreg[654]) );
  DFF \zreg_reg[655]  ( .D(o[655]), .CLK(clk), .RST(rst), .Q(zreg[655]) );
  DFF \zreg_reg[656]  ( .D(o[656]), .CLK(clk), .RST(rst), .Q(zreg[656]) );
  DFF \zreg_reg[657]  ( .D(o[657]), .CLK(clk), .RST(rst), .Q(zreg[657]) );
  DFF \zreg_reg[658]  ( .D(o[658]), .CLK(clk), .RST(rst), .Q(zreg[658]) );
  DFF \zreg_reg[659]  ( .D(o[659]), .CLK(clk), .RST(rst), .Q(zreg[659]) );
  DFF \zreg_reg[660]  ( .D(o[660]), .CLK(clk), .RST(rst), .Q(zreg[660]) );
  DFF \zreg_reg[661]  ( .D(o[661]), .CLK(clk), .RST(rst), .Q(zreg[661]) );
  DFF \zreg_reg[662]  ( .D(o[662]), .CLK(clk), .RST(rst), .Q(zreg[662]) );
  DFF \zreg_reg[663]  ( .D(o[663]), .CLK(clk), .RST(rst), .Q(zreg[663]) );
  DFF \zreg_reg[664]  ( .D(o[664]), .CLK(clk), .RST(rst), .Q(zreg[664]) );
  DFF \zreg_reg[665]  ( .D(o[665]), .CLK(clk), .RST(rst), .Q(zreg[665]) );
  DFF \zreg_reg[666]  ( .D(o[666]), .CLK(clk), .RST(rst), .Q(zreg[666]) );
  DFF \zreg_reg[667]  ( .D(o[667]), .CLK(clk), .RST(rst), .Q(zreg[667]) );
  DFF \zreg_reg[668]  ( .D(o[668]), .CLK(clk), .RST(rst), .Q(zreg[668]) );
  DFF \zreg_reg[669]  ( .D(o[669]), .CLK(clk), .RST(rst), .Q(zreg[669]) );
  DFF \zreg_reg[670]  ( .D(o[670]), .CLK(clk), .RST(rst), .Q(zreg[670]) );
  DFF \zreg_reg[671]  ( .D(o[671]), .CLK(clk), .RST(rst), .Q(zreg[671]) );
  DFF \zreg_reg[672]  ( .D(o[672]), .CLK(clk), .RST(rst), .Q(zreg[672]) );
  DFF \zreg_reg[673]  ( .D(o[673]), .CLK(clk), .RST(rst), .Q(zreg[673]) );
  DFF \zreg_reg[674]  ( .D(o[674]), .CLK(clk), .RST(rst), .Q(zreg[674]) );
  DFF \zreg_reg[675]  ( .D(o[675]), .CLK(clk), .RST(rst), .Q(zreg[675]) );
  DFF \zreg_reg[676]  ( .D(o[676]), .CLK(clk), .RST(rst), .Q(zreg[676]) );
  DFF \zreg_reg[677]  ( .D(o[677]), .CLK(clk), .RST(rst), .Q(zreg[677]) );
  DFF \zreg_reg[678]  ( .D(o[678]), .CLK(clk), .RST(rst), .Q(zreg[678]) );
  DFF \zreg_reg[679]  ( .D(o[679]), .CLK(clk), .RST(rst), .Q(zreg[679]) );
  DFF \zreg_reg[680]  ( .D(o[680]), .CLK(clk), .RST(rst), .Q(zreg[680]) );
  DFF \zreg_reg[681]  ( .D(o[681]), .CLK(clk), .RST(rst), .Q(zreg[681]) );
  DFF \zreg_reg[682]  ( .D(o[682]), .CLK(clk), .RST(rst), .Q(zreg[682]) );
  DFF \zreg_reg[683]  ( .D(o[683]), .CLK(clk), .RST(rst), .Q(zreg[683]) );
  DFF \zreg_reg[684]  ( .D(o[684]), .CLK(clk), .RST(rst), .Q(zreg[684]) );
  DFF \zreg_reg[685]  ( .D(o[685]), .CLK(clk), .RST(rst), .Q(zreg[685]) );
  DFF \zreg_reg[686]  ( .D(o[686]), .CLK(clk), .RST(rst), .Q(zreg[686]) );
  DFF \zreg_reg[687]  ( .D(o[687]), .CLK(clk), .RST(rst), .Q(zreg[687]) );
  DFF \zreg_reg[688]  ( .D(o[688]), .CLK(clk), .RST(rst), .Q(zreg[688]) );
  DFF \zreg_reg[689]  ( .D(o[689]), .CLK(clk), .RST(rst), .Q(zreg[689]) );
  DFF \zreg_reg[690]  ( .D(o[690]), .CLK(clk), .RST(rst), .Q(zreg[690]) );
  DFF \zreg_reg[691]  ( .D(o[691]), .CLK(clk), .RST(rst), .Q(zreg[691]) );
  DFF \zreg_reg[692]  ( .D(o[692]), .CLK(clk), .RST(rst), .Q(zreg[692]) );
  DFF \zreg_reg[693]  ( .D(o[693]), .CLK(clk), .RST(rst), .Q(zreg[693]) );
  DFF \zreg_reg[694]  ( .D(o[694]), .CLK(clk), .RST(rst), .Q(zreg[694]) );
  DFF \zreg_reg[695]  ( .D(o[695]), .CLK(clk), .RST(rst), .Q(zreg[695]) );
  DFF \zreg_reg[696]  ( .D(o[696]), .CLK(clk), .RST(rst), .Q(zreg[696]) );
  DFF \zreg_reg[697]  ( .D(o[697]), .CLK(clk), .RST(rst), .Q(zreg[697]) );
  DFF \zreg_reg[698]  ( .D(o[698]), .CLK(clk), .RST(rst), .Q(zreg[698]) );
  DFF \zreg_reg[699]  ( .D(o[699]), .CLK(clk), .RST(rst), .Q(zreg[699]) );
  DFF \zreg_reg[700]  ( .D(o[700]), .CLK(clk), .RST(rst), .Q(zreg[700]) );
  DFF \zreg_reg[701]  ( .D(o[701]), .CLK(clk), .RST(rst), .Q(zreg[701]) );
  DFF \zreg_reg[702]  ( .D(o[702]), .CLK(clk), .RST(rst), .Q(zreg[702]) );
  DFF \zreg_reg[703]  ( .D(o[703]), .CLK(clk), .RST(rst), .Q(zreg[703]) );
  DFF \zreg_reg[704]  ( .D(o[704]), .CLK(clk), .RST(rst), .Q(zreg[704]) );
  DFF \zreg_reg[705]  ( .D(o[705]), .CLK(clk), .RST(rst), .Q(zreg[705]) );
  DFF \zreg_reg[706]  ( .D(o[706]), .CLK(clk), .RST(rst), .Q(zreg[706]) );
  DFF \zreg_reg[707]  ( .D(o[707]), .CLK(clk), .RST(rst), .Q(zreg[707]) );
  DFF \zreg_reg[708]  ( .D(o[708]), .CLK(clk), .RST(rst), .Q(zreg[708]) );
  DFF \zreg_reg[709]  ( .D(o[709]), .CLK(clk), .RST(rst), .Q(zreg[709]) );
  DFF \zreg_reg[710]  ( .D(o[710]), .CLK(clk), .RST(rst), .Q(zreg[710]) );
  DFF \zreg_reg[711]  ( .D(o[711]), .CLK(clk), .RST(rst), .Q(zreg[711]) );
  DFF \zreg_reg[712]  ( .D(o[712]), .CLK(clk), .RST(rst), .Q(zreg[712]) );
  DFF \zreg_reg[713]  ( .D(o[713]), .CLK(clk), .RST(rst), .Q(zreg[713]) );
  DFF \zreg_reg[714]  ( .D(o[714]), .CLK(clk), .RST(rst), .Q(zreg[714]) );
  DFF \zreg_reg[715]  ( .D(o[715]), .CLK(clk), .RST(rst), .Q(zreg[715]) );
  DFF \zreg_reg[716]  ( .D(o[716]), .CLK(clk), .RST(rst), .Q(zreg[716]) );
  DFF \zreg_reg[717]  ( .D(o[717]), .CLK(clk), .RST(rst), .Q(zreg[717]) );
  DFF \zreg_reg[718]  ( .D(o[718]), .CLK(clk), .RST(rst), .Q(zreg[718]) );
  DFF \zreg_reg[719]  ( .D(o[719]), .CLK(clk), .RST(rst), .Q(zreg[719]) );
  DFF \zreg_reg[720]  ( .D(o[720]), .CLK(clk), .RST(rst), .Q(zreg[720]) );
  DFF \zreg_reg[721]  ( .D(o[721]), .CLK(clk), .RST(rst), .Q(zreg[721]) );
  DFF \zreg_reg[722]  ( .D(o[722]), .CLK(clk), .RST(rst), .Q(zreg[722]) );
  DFF \zreg_reg[723]  ( .D(o[723]), .CLK(clk), .RST(rst), .Q(zreg[723]) );
  DFF \zreg_reg[724]  ( .D(o[724]), .CLK(clk), .RST(rst), .Q(zreg[724]) );
  DFF \zreg_reg[725]  ( .D(o[725]), .CLK(clk), .RST(rst), .Q(zreg[725]) );
  DFF \zreg_reg[726]  ( .D(o[726]), .CLK(clk), .RST(rst), .Q(zreg[726]) );
  DFF \zreg_reg[727]  ( .D(o[727]), .CLK(clk), .RST(rst), .Q(zreg[727]) );
  DFF \zreg_reg[728]  ( .D(o[728]), .CLK(clk), .RST(rst), .Q(zreg[728]) );
  DFF \zreg_reg[729]  ( .D(o[729]), .CLK(clk), .RST(rst), .Q(zreg[729]) );
  DFF \zreg_reg[730]  ( .D(o[730]), .CLK(clk), .RST(rst), .Q(zreg[730]) );
  DFF \zreg_reg[731]  ( .D(o[731]), .CLK(clk), .RST(rst), .Q(zreg[731]) );
  DFF \zreg_reg[732]  ( .D(o[732]), .CLK(clk), .RST(rst), .Q(zreg[732]) );
  DFF \zreg_reg[733]  ( .D(o[733]), .CLK(clk), .RST(rst), .Q(zreg[733]) );
  DFF \zreg_reg[734]  ( .D(o[734]), .CLK(clk), .RST(rst), .Q(zreg[734]) );
  DFF \zreg_reg[735]  ( .D(o[735]), .CLK(clk), .RST(rst), .Q(zreg[735]) );
  DFF \zreg_reg[736]  ( .D(o[736]), .CLK(clk), .RST(rst), .Q(zreg[736]) );
  DFF \zreg_reg[737]  ( .D(o[737]), .CLK(clk), .RST(rst), .Q(zreg[737]) );
  DFF \zreg_reg[738]  ( .D(o[738]), .CLK(clk), .RST(rst), .Q(zreg[738]) );
  DFF \zreg_reg[739]  ( .D(o[739]), .CLK(clk), .RST(rst), .Q(zreg[739]) );
  DFF \zreg_reg[740]  ( .D(o[740]), .CLK(clk), .RST(rst), .Q(zreg[740]) );
  DFF \zreg_reg[741]  ( .D(o[741]), .CLK(clk), .RST(rst), .Q(zreg[741]) );
  DFF \zreg_reg[742]  ( .D(o[742]), .CLK(clk), .RST(rst), .Q(zreg[742]) );
  DFF \zreg_reg[743]  ( .D(o[743]), .CLK(clk), .RST(rst), .Q(zreg[743]) );
  DFF \zreg_reg[744]  ( .D(o[744]), .CLK(clk), .RST(rst), .Q(zreg[744]) );
  DFF \zreg_reg[745]  ( .D(o[745]), .CLK(clk), .RST(rst), .Q(zreg[745]) );
  DFF \zreg_reg[746]  ( .D(o[746]), .CLK(clk), .RST(rst), .Q(zreg[746]) );
  DFF \zreg_reg[747]  ( .D(o[747]), .CLK(clk), .RST(rst), .Q(zreg[747]) );
  DFF \zreg_reg[748]  ( .D(o[748]), .CLK(clk), .RST(rst), .Q(zreg[748]) );
  DFF \zreg_reg[749]  ( .D(o[749]), .CLK(clk), .RST(rst), .Q(zreg[749]) );
  DFF \zreg_reg[750]  ( .D(o[750]), .CLK(clk), .RST(rst), .Q(zreg[750]) );
  DFF \zreg_reg[751]  ( .D(o[751]), .CLK(clk), .RST(rst), .Q(zreg[751]) );
  DFF \zreg_reg[752]  ( .D(o[752]), .CLK(clk), .RST(rst), .Q(zreg[752]) );
  DFF \zreg_reg[753]  ( .D(o[753]), .CLK(clk), .RST(rst), .Q(zreg[753]) );
  DFF \zreg_reg[754]  ( .D(o[754]), .CLK(clk), .RST(rst), .Q(zreg[754]) );
  DFF \zreg_reg[755]  ( .D(o[755]), .CLK(clk), .RST(rst), .Q(zreg[755]) );
  DFF \zreg_reg[756]  ( .D(o[756]), .CLK(clk), .RST(rst), .Q(zreg[756]) );
  DFF \zreg_reg[757]  ( .D(o[757]), .CLK(clk), .RST(rst), .Q(zreg[757]) );
  DFF \zreg_reg[758]  ( .D(o[758]), .CLK(clk), .RST(rst), .Q(zreg[758]) );
  DFF \zreg_reg[759]  ( .D(o[759]), .CLK(clk), .RST(rst), .Q(zreg[759]) );
  DFF \zreg_reg[760]  ( .D(o[760]), .CLK(clk), .RST(rst), .Q(zreg[760]) );
  DFF \zreg_reg[761]  ( .D(o[761]), .CLK(clk), .RST(rst), .Q(zreg[761]) );
  DFF \zreg_reg[762]  ( .D(o[762]), .CLK(clk), .RST(rst), .Q(zreg[762]) );
  DFF \zreg_reg[763]  ( .D(o[763]), .CLK(clk), .RST(rst), .Q(zreg[763]) );
  DFF \zreg_reg[764]  ( .D(o[764]), .CLK(clk), .RST(rst), .Q(zreg[764]) );
  DFF \zreg_reg[765]  ( .D(o[765]), .CLK(clk), .RST(rst), .Q(zreg[765]) );
  DFF \zreg_reg[766]  ( .D(o[766]), .CLK(clk), .RST(rst), .Q(zreg[766]) );
  DFF \zreg_reg[767]  ( .D(o[767]), .CLK(clk), .RST(rst), .Q(zreg[767]) );
  DFF \zreg_reg[768]  ( .D(o[768]), .CLK(clk), .RST(rst), .Q(zreg[768]) );
  DFF \zreg_reg[769]  ( .D(o[769]), .CLK(clk), .RST(rst), .Q(zreg[769]) );
  DFF \zreg_reg[770]  ( .D(o[770]), .CLK(clk), .RST(rst), .Q(zreg[770]) );
  DFF \zreg_reg[771]  ( .D(o[771]), .CLK(clk), .RST(rst), .Q(zreg[771]) );
  DFF \zreg_reg[772]  ( .D(o[772]), .CLK(clk), .RST(rst), .Q(zreg[772]) );
  DFF \zreg_reg[773]  ( .D(o[773]), .CLK(clk), .RST(rst), .Q(zreg[773]) );
  DFF \zreg_reg[774]  ( .D(o[774]), .CLK(clk), .RST(rst), .Q(zreg[774]) );
  DFF \zreg_reg[775]  ( .D(o[775]), .CLK(clk), .RST(rst), .Q(zreg[775]) );
  DFF \zreg_reg[776]  ( .D(o[776]), .CLK(clk), .RST(rst), .Q(zreg[776]) );
  DFF \zreg_reg[777]  ( .D(o[777]), .CLK(clk), .RST(rst), .Q(zreg[777]) );
  DFF \zreg_reg[778]  ( .D(o[778]), .CLK(clk), .RST(rst), .Q(zreg[778]) );
  DFF \zreg_reg[779]  ( .D(o[779]), .CLK(clk), .RST(rst), .Q(zreg[779]) );
  DFF \zreg_reg[780]  ( .D(o[780]), .CLK(clk), .RST(rst), .Q(zreg[780]) );
  DFF \zreg_reg[781]  ( .D(o[781]), .CLK(clk), .RST(rst), .Q(zreg[781]) );
  DFF \zreg_reg[782]  ( .D(o[782]), .CLK(clk), .RST(rst), .Q(zreg[782]) );
  DFF \zreg_reg[783]  ( .D(o[783]), .CLK(clk), .RST(rst), .Q(zreg[783]) );
  DFF \zreg_reg[784]  ( .D(o[784]), .CLK(clk), .RST(rst), .Q(zreg[784]) );
  DFF \zreg_reg[785]  ( .D(o[785]), .CLK(clk), .RST(rst), .Q(zreg[785]) );
  DFF \zreg_reg[786]  ( .D(o[786]), .CLK(clk), .RST(rst), .Q(zreg[786]) );
  DFF \zreg_reg[787]  ( .D(o[787]), .CLK(clk), .RST(rst), .Q(zreg[787]) );
  DFF \zreg_reg[788]  ( .D(o[788]), .CLK(clk), .RST(rst), .Q(zreg[788]) );
  DFF \zreg_reg[789]  ( .D(o[789]), .CLK(clk), .RST(rst), .Q(zreg[789]) );
  DFF \zreg_reg[790]  ( .D(o[790]), .CLK(clk), .RST(rst), .Q(zreg[790]) );
  DFF \zreg_reg[791]  ( .D(o[791]), .CLK(clk), .RST(rst), .Q(zreg[791]) );
  DFF \zreg_reg[792]  ( .D(o[792]), .CLK(clk), .RST(rst), .Q(zreg[792]) );
  DFF \zreg_reg[793]  ( .D(o[793]), .CLK(clk), .RST(rst), .Q(zreg[793]) );
  DFF \zreg_reg[794]  ( .D(o[794]), .CLK(clk), .RST(rst), .Q(zreg[794]) );
  DFF \zreg_reg[795]  ( .D(o[795]), .CLK(clk), .RST(rst), .Q(zreg[795]) );
  DFF \zreg_reg[796]  ( .D(o[796]), .CLK(clk), .RST(rst), .Q(zreg[796]) );
  DFF \zreg_reg[797]  ( .D(o[797]), .CLK(clk), .RST(rst), .Q(zreg[797]) );
  DFF \zreg_reg[798]  ( .D(o[798]), .CLK(clk), .RST(rst), .Q(zreg[798]) );
  DFF \zreg_reg[799]  ( .D(o[799]), .CLK(clk), .RST(rst), .Q(zreg[799]) );
  DFF \zreg_reg[800]  ( .D(o[800]), .CLK(clk), .RST(rst), .Q(zreg[800]) );
  DFF \zreg_reg[801]  ( .D(o[801]), .CLK(clk), .RST(rst), .Q(zreg[801]) );
  DFF \zreg_reg[802]  ( .D(o[802]), .CLK(clk), .RST(rst), .Q(zreg[802]) );
  DFF \zreg_reg[803]  ( .D(o[803]), .CLK(clk), .RST(rst), .Q(zreg[803]) );
  DFF \zreg_reg[804]  ( .D(o[804]), .CLK(clk), .RST(rst), .Q(zreg[804]) );
  DFF \zreg_reg[805]  ( .D(o[805]), .CLK(clk), .RST(rst), .Q(zreg[805]) );
  DFF \zreg_reg[806]  ( .D(o[806]), .CLK(clk), .RST(rst), .Q(zreg[806]) );
  DFF \zreg_reg[807]  ( .D(o[807]), .CLK(clk), .RST(rst), .Q(zreg[807]) );
  DFF \zreg_reg[808]  ( .D(o[808]), .CLK(clk), .RST(rst), .Q(zreg[808]) );
  DFF \zreg_reg[809]  ( .D(o[809]), .CLK(clk), .RST(rst), .Q(zreg[809]) );
  DFF \zreg_reg[810]  ( .D(o[810]), .CLK(clk), .RST(rst), .Q(zreg[810]) );
  DFF \zreg_reg[811]  ( .D(o[811]), .CLK(clk), .RST(rst), .Q(zreg[811]) );
  DFF \zreg_reg[812]  ( .D(o[812]), .CLK(clk), .RST(rst), .Q(zreg[812]) );
  DFF \zreg_reg[813]  ( .D(o[813]), .CLK(clk), .RST(rst), .Q(zreg[813]) );
  DFF \zreg_reg[814]  ( .D(o[814]), .CLK(clk), .RST(rst), .Q(zreg[814]) );
  DFF \zreg_reg[815]  ( .D(o[815]), .CLK(clk), .RST(rst), .Q(zreg[815]) );
  DFF \zreg_reg[816]  ( .D(o[816]), .CLK(clk), .RST(rst), .Q(zreg[816]) );
  DFF \zreg_reg[817]  ( .D(o[817]), .CLK(clk), .RST(rst), .Q(zreg[817]) );
  DFF \zreg_reg[818]  ( .D(o[818]), .CLK(clk), .RST(rst), .Q(zreg[818]) );
  DFF \zreg_reg[819]  ( .D(o[819]), .CLK(clk), .RST(rst), .Q(zreg[819]) );
  DFF \zreg_reg[820]  ( .D(o[820]), .CLK(clk), .RST(rst), .Q(zreg[820]) );
  DFF \zreg_reg[821]  ( .D(o[821]), .CLK(clk), .RST(rst), .Q(zreg[821]) );
  DFF \zreg_reg[822]  ( .D(o[822]), .CLK(clk), .RST(rst), .Q(zreg[822]) );
  DFF \zreg_reg[823]  ( .D(o[823]), .CLK(clk), .RST(rst), .Q(zreg[823]) );
  DFF \zreg_reg[824]  ( .D(o[824]), .CLK(clk), .RST(rst), .Q(zreg[824]) );
  DFF \zreg_reg[825]  ( .D(o[825]), .CLK(clk), .RST(rst), .Q(zreg[825]) );
  DFF \zreg_reg[826]  ( .D(o[826]), .CLK(clk), .RST(rst), .Q(zreg[826]) );
  DFF \zreg_reg[827]  ( .D(o[827]), .CLK(clk), .RST(rst), .Q(zreg[827]) );
  DFF \zreg_reg[828]  ( .D(o[828]), .CLK(clk), .RST(rst), .Q(zreg[828]) );
  DFF \zreg_reg[829]  ( .D(o[829]), .CLK(clk), .RST(rst), .Q(zreg[829]) );
  DFF \zreg_reg[830]  ( .D(o[830]), .CLK(clk), .RST(rst), .Q(zreg[830]) );
  DFF \zreg_reg[831]  ( .D(o[831]), .CLK(clk), .RST(rst), .Q(zreg[831]) );
  DFF \zreg_reg[832]  ( .D(o[832]), .CLK(clk), .RST(rst), .Q(zreg[832]) );
  DFF \zreg_reg[833]  ( .D(o[833]), .CLK(clk), .RST(rst), .Q(zreg[833]) );
  DFF \zreg_reg[834]  ( .D(o[834]), .CLK(clk), .RST(rst), .Q(zreg[834]) );
  DFF \zreg_reg[835]  ( .D(o[835]), .CLK(clk), .RST(rst), .Q(zreg[835]) );
  DFF \zreg_reg[836]  ( .D(o[836]), .CLK(clk), .RST(rst), .Q(zreg[836]) );
  DFF \zreg_reg[837]  ( .D(o[837]), .CLK(clk), .RST(rst), .Q(zreg[837]) );
  DFF \zreg_reg[838]  ( .D(o[838]), .CLK(clk), .RST(rst), .Q(zreg[838]) );
  DFF \zreg_reg[839]  ( .D(o[839]), .CLK(clk), .RST(rst), .Q(zreg[839]) );
  DFF \zreg_reg[840]  ( .D(o[840]), .CLK(clk), .RST(rst), .Q(zreg[840]) );
  DFF \zreg_reg[841]  ( .D(o[841]), .CLK(clk), .RST(rst), .Q(zreg[841]) );
  DFF \zreg_reg[842]  ( .D(o[842]), .CLK(clk), .RST(rst), .Q(zreg[842]) );
  DFF \zreg_reg[843]  ( .D(o[843]), .CLK(clk), .RST(rst), .Q(zreg[843]) );
  DFF \zreg_reg[844]  ( .D(o[844]), .CLK(clk), .RST(rst), .Q(zreg[844]) );
  DFF \zreg_reg[845]  ( .D(o[845]), .CLK(clk), .RST(rst), .Q(zreg[845]) );
  DFF \zreg_reg[846]  ( .D(o[846]), .CLK(clk), .RST(rst), .Q(zreg[846]) );
  DFF \zreg_reg[847]  ( .D(o[847]), .CLK(clk), .RST(rst), .Q(zreg[847]) );
  DFF \zreg_reg[848]  ( .D(o[848]), .CLK(clk), .RST(rst), .Q(zreg[848]) );
  DFF \zreg_reg[849]  ( .D(o[849]), .CLK(clk), .RST(rst), .Q(zreg[849]) );
  DFF \zreg_reg[850]  ( .D(o[850]), .CLK(clk), .RST(rst), .Q(zreg[850]) );
  DFF \zreg_reg[851]  ( .D(o[851]), .CLK(clk), .RST(rst), .Q(zreg[851]) );
  DFF \zreg_reg[852]  ( .D(o[852]), .CLK(clk), .RST(rst), .Q(zreg[852]) );
  DFF \zreg_reg[853]  ( .D(o[853]), .CLK(clk), .RST(rst), .Q(zreg[853]) );
  DFF \zreg_reg[854]  ( .D(o[854]), .CLK(clk), .RST(rst), .Q(zreg[854]) );
  DFF \zreg_reg[855]  ( .D(o[855]), .CLK(clk), .RST(rst), .Q(zreg[855]) );
  DFF \zreg_reg[856]  ( .D(o[856]), .CLK(clk), .RST(rst), .Q(zreg[856]) );
  DFF \zreg_reg[857]  ( .D(o[857]), .CLK(clk), .RST(rst), .Q(zreg[857]) );
  DFF \zreg_reg[858]  ( .D(o[858]), .CLK(clk), .RST(rst), .Q(zreg[858]) );
  DFF \zreg_reg[859]  ( .D(o[859]), .CLK(clk), .RST(rst), .Q(zreg[859]) );
  DFF \zreg_reg[860]  ( .D(o[860]), .CLK(clk), .RST(rst), .Q(zreg[860]) );
  DFF \zreg_reg[861]  ( .D(o[861]), .CLK(clk), .RST(rst), .Q(zreg[861]) );
  DFF \zreg_reg[862]  ( .D(o[862]), .CLK(clk), .RST(rst), .Q(zreg[862]) );
  DFF \zreg_reg[863]  ( .D(o[863]), .CLK(clk), .RST(rst), .Q(zreg[863]) );
  DFF \zreg_reg[864]  ( .D(o[864]), .CLK(clk), .RST(rst), .Q(zreg[864]) );
  DFF \zreg_reg[865]  ( .D(o[865]), .CLK(clk), .RST(rst), .Q(zreg[865]) );
  DFF \zreg_reg[866]  ( .D(o[866]), .CLK(clk), .RST(rst), .Q(zreg[866]) );
  DFF \zreg_reg[867]  ( .D(o[867]), .CLK(clk), .RST(rst), .Q(zreg[867]) );
  DFF \zreg_reg[868]  ( .D(o[868]), .CLK(clk), .RST(rst), .Q(zreg[868]) );
  DFF \zreg_reg[869]  ( .D(o[869]), .CLK(clk), .RST(rst), .Q(zreg[869]) );
  DFF \zreg_reg[870]  ( .D(o[870]), .CLK(clk), .RST(rst), .Q(zreg[870]) );
  DFF \zreg_reg[871]  ( .D(o[871]), .CLK(clk), .RST(rst), .Q(zreg[871]) );
  DFF \zreg_reg[872]  ( .D(o[872]), .CLK(clk), .RST(rst), .Q(zreg[872]) );
  DFF \zreg_reg[873]  ( .D(o[873]), .CLK(clk), .RST(rst), .Q(zreg[873]) );
  DFF \zreg_reg[874]  ( .D(o[874]), .CLK(clk), .RST(rst), .Q(zreg[874]) );
  DFF \zreg_reg[875]  ( .D(o[875]), .CLK(clk), .RST(rst), .Q(zreg[875]) );
  DFF \zreg_reg[876]  ( .D(o[876]), .CLK(clk), .RST(rst), .Q(zreg[876]) );
  DFF \zreg_reg[877]  ( .D(o[877]), .CLK(clk), .RST(rst), .Q(zreg[877]) );
  DFF \zreg_reg[878]  ( .D(o[878]), .CLK(clk), .RST(rst), .Q(zreg[878]) );
  DFF \zreg_reg[879]  ( .D(o[879]), .CLK(clk), .RST(rst), .Q(zreg[879]) );
  DFF \zreg_reg[880]  ( .D(o[880]), .CLK(clk), .RST(rst), .Q(zreg[880]) );
  DFF \zreg_reg[881]  ( .D(o[881]), .CLK(clk), .RST(rst), .Q(zreg[881]) );
  DFF \zreg_reg[882]  ( .D(o[882]), .CLK(clk), .RST(rst), .Q(zreg[882]) );
  DFF \zreg_reg[883]  ( .D(o[883]), .CLK(clk), .RST(rst), .Q(zreg[883]) );
  DFF \zreg_reg[884]  ( .D(o[884]), .CLK(clk), .RST(rst), .Q(zreg[884]) );
  DFF \zreg_reg[885]  ( .D(o[885]), .CLK(clk), .RST(rst), .Q(zreg[885]) );
  DFF \zreg_reg[886]  ( .D(o[886]), .CLK(clk), .RST(rst), .Q(zreg[886]) );
  DFF \zreg_reg[887]  ( .D(o[887]), .CLK(clk), .RST(rst), .Q(zreg[887]) );
  DFF \zreg_reg[888]  ( .D(o[888]), .CLK(clk), .RST(rst), .Q(zreg[888]) );
  DFF \zreg_reg[889]  ( .D(o[889]), .CLK(clk), .RST(rst), .Q(zreg[889]) );
  DFF \zreg_reg[890]  ( .D(o[890]), .CLK(clk), .RST(rst), .Q(zreg[890]) );
  DFF \zreg_reg[891]  ( .D(o[891]), .CLK(clk), .RST(rst), .Q(zreg[891]) );
  DFF \zreg_reg[892]  ( .D(o[892]), .CLK(clk), .RST(rst), .Q(zreg[892]) );
  DFF \zreg_reg[893]  ( .D(o[893]), .CLK(clk), .RST(rst), .Q(zreg[893]) );
  DFF \zreg_reg[894]  ( .D(o[894]), .CLK(clk), .RST(rst), .Q(zreg[894]) );
  DFF \zreg_reg[895]  ( .D(o[895]), .CLK(clk), .RST(rst), .Q(zreg[895]) );
  DFF \zreg_reg[896]  ( .D(o[896]), .CLK(clk), .RST(rst), .Q(zreg[896]) );
  DFF \zreg_reg[897]  ( .D(o[897]), .CLK(clk), .RST(rst), .Q(zreg[897]) );
  DFF \zreg_reg[898]  ( .D(o[898]), .CLK(clk), .RST(rst), .Q(zreg[898]) );
  DFF \zreg_reg[899]  ( .D(o[899]), .CLK(clk), .RST(rst), .Q(zreg[899]) );
  DFF \zreg_reg[900]  ( .D(o[900]), .CLK(clk), .RST(rst), .Q(zreg[900]) );
  DFF \zreg_reg[901]  ( .D(o[901]), .CLK(clk), .RST(rst), .Q(zreg[901]) );
  DFF \zreg_reg[902]  ( .D(o[902]), .CLK(clk), .RST(rst), .Q(zreg[902]) );
  DFF \zreg_reg[903]  ( .D(o[903]), .CLK(clk), .RST(rst), .Q(zreg[903]) );
  DFF \zreg_reg[904]  ( .D(o[904]), .CLK(clk), .RST(rst), .Q(zreg[904]) );
  DFF \zreg_reg[905]  ( .D(o[905]), .CLK(clk), .RST(rst), .Q(zreg[905]) );
  DFF \zreg_reg[906]  ( .D(o[906]), .CLK(clk), .RST(rst), .Q(zreg[906]) );
  DFF \zreg_reg[907]  ( .D(o[907]), .CLK(clk), .RST(rst), .Q(zreg[907]) );
  DFF \zreg_reg[908]  ( .D(o[908]), .CLK(clk), .RST(rst), .Q(zreg[908]) );
  DFF \zreg_reg[909]  ( .D(o[909]), .CLK(clk), .RST(rst), .Q(zreg[909]) );
  DFF \zreg_reg[910]  ( .D(o[910]), .CLK(clk), .RST(rst), .Q(zreg[910]) );
  DFF \zreg_reg[911]  ( .D(o[911]), .CLK(clk), .RST(rst), .Q(zreg[911]) );
  DFF \zreg_reg[912]  ( .D(o[912]), .CLK(clk), .RST(rst), .Q(zreg[912]) );
  DFF \zreg_reg[913]  ( .D(o[913]), .CLK(clk), .RST(rst), .Q(zreg[913]) );
  DFF \zreg_reg[914]  ( .D(o[914]), .CLK(clk), .RST(rst), .Q(zreg[914]) );
  DFF \zreg_reg[915]  ( .D(o[915]), .CLK(clk), .RST(rst), .Q(zreg[915]) );
  DFF \zreg_reg[916]  ( .D(o[916]), .CLK(clk), .RST(rst), .Q(zreg[916]) );
  DFF \zreg_reg[917]  ( .D(o[917]), .CLK(clk), .RST(rst), .Q(zreg[917]) );
  DFF \zreg_reg[918]  ( .D(o[918]), .CLK(clk), .RST(rst), .Q(zreg[918]) );
  DFF \zreg_reg[919]  ( .D(o[919]), .CLK(clk), .RST(rst), .Q(zreg[919]) );
  DFF \zreg_reg[920]  ( .D(o[920]), .CLK(clk), .RST(rst), .Q(zreg[920]) );
  DFF \zreg_reg[921]  ( .D(o[921]), .CLK(clk), .RST(rst), .Q(zreg[921]) );
  DFF \zreg_reg[922]  ( .D(o[922]), .CLK(clk), .RST(rst), .Q(zreg[922]) );
  DFF \zreg_reg[923]  ( .D(o[923]), .CLK(clk), .RST(rst), .Q(zreg[923]) );
  DFF \zreg_reg[924]  ( .D(o[924]), .CLK(clk), .RST(rst), .Q(zreg[924]) );
  DFF \zreg_reg[925]  ( .D(o[925]), .CLK(clk), .RST(rst), .Q(zreg[925]) );
  DFF \zreg_reg[926]  ( .D(o[926]), .CLK(clk), .RST(rst), .Q(zreg[926]) );
  DFF \zreg_reg[927]  ( .D(o[927]), .CLK(clk), .RST(rst), .Q(zreg[927]) );
  DFF \zreg_reg[928]  ( .D(o[928]), .CLK(clk), .RST(rst), .Q(zreg[928]) );
  DFF \zreg_reg[929]  ( .D(o[929]), .CLK(clk), .RST(rst), .Q(zreg[929]) );
  DFF \zreg_reg[930]  ( .D(o[930]), .CLK(clk), .RST(rst), .Q(zreg[930]) );
  DFF \zreg_reg[931]  ( .D(o[931]), .CLK(clk), .RST(rst), .Q(zreg[931]) );
  DFF \zreg_reg[932]  ( .D(o[932]), .CLK(clk), .RST(rst), .Q(zreg[932]) );
  DFF \zreg_reg[933]  ( .D(o[933]), .CLK(clk), .RST(rst), .Q(zreg[933]) );
  DFF \zreg_reg[934]  ( .D(o[934]), .CLK(clk), .RST(rst), .Q(zreg[934]) );
  DFF \zreg_reg[935]  ( .D(o[935]), .CLK(clk), .RST(rst), .Q(zreg[935]) );
  DFF \zreg_reg[936]  ( .D(o[936]), .CLK(clk), .RST(rst), .Q(zreg[936]) );
  DFF \zreg_reg[937]  ( .D(o[937]), .CLK(clk), .RST(rst), .Q(zreg[937]) );
  DFF \zreg_reg[938]  ( .D(o[938]), .CLK(clk), .RST(rst), .Q(zreg[938]) );
  DFF \zreg_reg[939]  ( .D(o[939]), .CLK(clk), .RST(rst), .Q(zreg[939]) );
  DFF \zreg_reg[940]  ( .D(o[940]), .CLK(clk), .RST(rst), .Q(zreg[940]) );
  DFF \zreg_reg[941]  ( .D(o[941]), .CLK(clk), .RST(rst), .Q(zreg[941]) );
  DFF \zreg_reg[942]  ( .D(o[942]), .CLK(clk), .RST(rst), .Q(zreg[942]) );
  DFF \zreg_reg[943]  ( .D(o[943]), .CLK(clk), .RST(rst), .Q(zreg[943]) );
  DFF \zreg_reg[944]  ( .D(o[944]), .CLK(clk), .RST(rst), .Q(zreg[944]) );
  DFF \zreg_reg[945]  ( .D(o[945]), .CLK(clk), .RST(rst), .Q(zreg[945]) );
  DFF \zreg_reg[946]  ( .D(o[946]), .CLK(clk), .RST(rst), .Q(zreg[946]) );
  DFF \zreg_reg[947]  ( .D(o[947]), .CLK(clk), .RST(rst), .Q(zreg[947]) );
  DFF \zreg_reg[948]  ( .D(o[948]), .CLK(clk), .RST(rst), .Q(zreg[948]) );
  DFF \zreg_reg[949]  ( .D(o[949]), .CLK(clk), .RST(rst), .Q(zreg[949]) );
  DFF \zreg_reg[950]  ( .D(o[950]), .CLK(clk), .RST(rst), .Q(zreg[950]) );
  DFF \zreg_reg[951]  ( .D(o[951]), .CLK(clk), .RST(rst), .Q(zreg[951]) );
  DFF \zreg_reg[952]  ( .D(o[952]), .CLK(clk), .RST(rst), .Q(zreg[952]) );
  DFF \zreg_reg[953]  ( .D(o[953]), .CLK(clk), .RST(rst), .Q(zreg[953]) );
  DFF \zreg_reg[954]  ( .D(o[954]), .CLK(clk), .RST(rst), .Q(zreg[954]) );
  DFF \zreg_reg[955]  ( .D(o[955]), .CLK(clk), .RST(rst), .Q(zreg[955]) );
  DFF \zreg_reg[956]  ( .D(o[956]), .CLK(clk), .RST(rst), .Q(zreg[956]) );
  DFF \zreg_reg[957]  ( .D(o[957]), .CLK(clk), .RST(rst), .Q(zreg[957]) );
  DFF \zreg_reg[958]  ( .D(o[958]), .CLK(clk), .RST(rst), .Q(zreg[958]) );
  DFF \zreg_reg[959]  ( .D(o[959]), .CLK(clk), .RST(rst), .Q(zreg[959]) );
  DFF \zreg_reg[960]  ( .D(o[960]), .CLK(clk), .RST(rst), .Q(zreg[960]) );
  DFF \zreg_reg[961]  ( .D(o[961]), .CLK(clk), .RST(rst), .Q(zreg[961]) );
  DFF \zreg_reg[962]  ( .D(o[962]), .CLK(clk), .RST(rst), .Q(zreg[962]) );
  DFF \zreg_reg[963]  ( .D(o[963]), .CLK(clk), .RST(rst), .Q(zreg[963]) );
  DFF \zreg_reg[964]  ( .D(o[964]), .CLK(clk), .RST(rst), .Q(zreg[964]) );
  DFF \zreg_reg[965]  ( .D(o[965]), .CLK(clk), .RST(rst), .Q(zreg[965]) );
  DFF \zreg_reg[966]  ( .D(o[966]), .CLK(clk), .RST(rst), .Q(zreg[966]) );
  DFF \zreg_reg[967]  ( .D(o[967]), .CLK(clk), .RST(rst), .Q(zreg[967]) );
  DFF \zreg_reg[968]  ( .D(o[968]), .CLK(clk), .RST(rst), .Q(zreg[968]) );
  DFF \zreg_reg[969]  ( .D(o[969]), .CLK(clk), .RST(rst), .Q(zreg[969]) );
  DFF \zreg_reg[970]  ( .D(o[970]), .CLK(clk), .RST(rst), .Q(zreg[970]) );
  DFF \zreg_reg[971]  ( .D(o[971]), .CLK(clk), .RST(rst), .Q(zreg[971]) );
  DFF \zreg_reg[972]  ( .D(o[972]), .CLK(clk), .RST(rst), .Q(zreg[972]) );
  DFF \zreg_reg[973]  ( .D(o[973]), .CLK(clk), .RST(rst), .Q(zreg[973]) );
  DFF \zreg_reg[974]  ( .D(o[974]), .CLK(clk), .RST(rst), .Q(zreg[974]) );
  DFF \zreg_reg[975]  ( .D(o[975]), .CLK(clk), .RST(rst), .Q(zreg[975]) );
  DFF \zreg_reg[976]  ( .D(o[976]), .CLK(clk), .RST(rst), .Q(zreg[976]) );
  DFF \zreg_reg[977]  ( .D(o[977]), .CLK(clk), .RST(rst), .Q(zreg[977]) );
  DFF \zreg_reg[978]  ( .D(o[978]), .CLK(clk), .RST(rst), .Q(zreg[978]) );
  DFF \zreg_reg[979]  ( .D(o[979]), .CLK(clk), .RST(rst), .Q(zreg[979]) );
  DFF \zreg_reg[980]  ( .D(o[980]), .CLK(clk), .RST(rst), .Q(zreg[980]) );
  DFF \zreg_reg[981]  ( .D(o[981]), .CLK(clk), .RST(rst), .Q(zreg[981]) );
  DFF \zreg_reg[982]  ( .D(o[982]), .CLK(clk), .RST(rst), .Q(zreg[982]) );
  DFF \zreg_reg[983]  ( .D(o[983]), .CLK(clk), .RST(rst), .Q(zreg[983]) );
  DFF \zreg_reg[984]  ( .D(o[984]), .CLK(clk), .RST(rst), .Q(zreg[984]) );
  DFF \zreg_reg[985]  ( .D(o[985]), .CLK(clk), .RST(rst), .Q(zreg[985]) );
  DFF \zreg_reg[986]  ( .D(o[986]), .CLK(clk), .RST(rst), .Q(zreg[986]) );
  DFF \zreg_reg[987]  ( .D(o[987]), .CLK(clk), .RST(rst), .Q(zreg[987]) );
  DFF \zreg_reg[988]  ( .D(o[988]), .CLK(clk), .RST(rst), .Q(zreg[988]) );
  DFF \zreg_reg[989]  ( .D(o[989]), .CLK(clk), .RST(rst), .Q(zreg[989]) );
  DFF \zreg_reg[990]  ( .D(o[990]), .CLK(clk), .RST(rst), .Q(zreg[990]) );
  DFF \zreg_reg[991]  ( .D(o[991]), .CLK(clk), .RST(rst), .Q(zreg[991]) );
  DFF \zreg_reg[992]  ( .D(o[992]), .CLK(clk), .RST(rst), .Q(zreg[992]) );
  DFF \zreg_reg[993]  ( .D(o[993]), .CLK(clk), .RST(rst), .Q(zreg[993]) );
  DFF \zreg_reg[994]  ( .D(o[994]), .CLK(clk), .RST(rst), .Q(zreg[994]) );
  DFF \zreg_reg[995]  ( .D(o[995]), .CLK(clk), .RST(rst), .Q(zreg[995]) );
  DFF \zreg_reg[996]  ( .D(o[996]), .CLK(clk), .RST(rst), .Q(zreg[996]) );
  DFF \zreg_reg[997]  ( .D(o[997]), .CLK(clk), .RST(rst), .Q(zreg[997]) );
  DFF \zreg_reg[998]  ( .D(o[998]), .CLK(clk), .RST(rst), .Q(zreg[998]) );
  DFF \zreg_reg[999]  ( .D(o[999]), .CLK(clk), .RST(rst), .Q(zreg[999]) );
  DFF \zreg_reg[1000]  ( .D(o[1000]), .CLK(clk), .RST(rst), .Q(zreg[1000]) );
  DFF \zreg_reg[1001]  ( .D(o[1001]), .CLK(clk), .RST(rst), .Q(zreg[1001]) );
  DFF \zreg_reg[1002]  ( .D(o[1002]), .CLK(clk), .RST(rst), .Q(zreg[1002]) );
  DFF \zreg_reg[1003]  ( .D(o[1003]), .CLK(clk), .RST(rst), .Q(zreg[1003]) );
  DFF \zreg_reg[1004]  ( .D(o[1004]), .CLK(clk), .RST(rst), .Q(zreg[1004]) );
  DFF \zreg_reg[1005]  ( .D(o[1005]), .CLK(clk), .RST(rst), .Q(zreg[1005]) );
  DFF \zreg_reg[1006]  ( .D(o[1006]), .CLK(clk), .RST(rst), .Q(zreg[1006]) );
  DFF \zreg_reg[1007]  ( .D(o[1007]), .CLK(clk), .RST(rst), .Q(zreg[1007]) );
  DFF \zreg_reg[1008]  ( .D(o[1008]), .CLK(clk), .RST(rst), .Q(zreg[1008]) );
  DFF \zreg_reg[1009]  ( .D(o[1009]), .CLK(clk), .RST(rst), .Q(zreg[1009]) );
  DFF \zreg_reg[1010]  ( .D(o[1010]), .CLK(clk), .RST(rst), .Q(zreg[1010]) );
  DFF \zreg_reg[1011]  ( .D(o[1011]), .CLK(clk), .RST(rst), .Q(zreg[1011]) );
  DFF \zreg_reg[1012]  ( .D(o[1012]), .CLK(clk), .RST(rst), .Q(zreg[1012]) );
  DFF \zreg_reg[1013]  ( .D(o[1013]), .CLK(clk), .RST(rst), .Q(zreg[1013]) );
  DFF \zreg_reg[1014]  ( .D(o[1014]), .CLK(clk), .RST(rst), .Q(zreg[1014]) );
  DFF \zreg_reg[1015]  ( .D(o[1015]), .CLK(clk), .RST(rst), .Q(zreg[1015]) );
  DFF \zreg_reg[1016]  ( .D(o[1016]), .CLK(clk), .RST(rst), .Q(zreg[1016]) );
  DFF \zreg_reg[1017]  ( .D(o[1017]), .CLK(clk), .RST(rst), .Q(zreg[1017]) );
  DFF \zreg_reg[1018]  ( .D(o[1018]), .CLK(clk), .RST(rst), .Q(zreg[1018]) );
  DFF \zreg_reg[1019]  ( .D(o[1019]), .CLK(clk), .RST(rst), .Q(zreg[1019]) );
  DFF \zreg_reg[1020]  ( .D(o[1020]), .CLK(clk), .RST(rst), .Q(zreg[1020]) );
  DFF \zreg_reg[1021]  ( .D(o[1021]), .CLK(clk), .RST(rst), .Q(zreg[1021]) );
  DFF \zreg_reg[1022]  ( .D(o[1022]), .CLK(clk), .RST(rst), .Q(zreg[1022]) );
  DFF \zreg_reg[1023]  ( .D(o[1023]), .CLK(clk), .RST(rst), .Q(zreg[1023]) );
  DFF \zreg_reg[1024]  ( .D(\zout[0][1024] ), .CLK(clk), .RST(rst), .Q(
        zreg[1024]) );
  DFF \zreg_reg[1025]  ( .D(\zout[0][1025] ), .CLK(clk), .RST(rst), .Q(
        zreg[1025]) );
  modmult_step_N1024 \MODMULT_STEP[0].modmult_step_  ( .xregN_1(xin[1023]), 
        .y(y), .n(n), .zin({\zin[0][1025] , \zin[0][1024] , \zin[0][1023] , 
        \zin[0][1022] , \zin[0][1021] , \zin[0][1020] , \zin[0][1019] , 
        \zin[0][1018] , \zin[0][1017] , \zin[0][1016] , \zin[0][1015] , 
        \zin[0][1014] , \zin[0][1013] , \zin[0][1012] , \zin[0][1011] , 
        \zin[0][1010] , \zin[0][1009] , \zin[0][1008] , \zin[0][1007] , 
        \zin[0][1006] , \zin[0][1005] , \zin[0][1004] , \zin[0][1003] , 
        \zin[0][1002] , \zin[0][1001] , \zin[0][1000] , \zin[0][999] , 
        \zin[0][998] , \zin[0][997] , \zin[0][996] , \zin[0][995] , 
        \zin[0][994] , \zin[0][993] , \zin[0][992] , \zin[0][991] , 
        \zin[0][990] , \zin[0][989] , \zin[0][988] , \zin[0][987] , 
        \zin[0][986] , \zin[0][985] , \zin[0][984] , \zin[0][983] , 
        \zin[0][982] , \zin[0][981] , \zin[0][980] , \zin[0][979] , 
        \zin[0][978] , \zin[0][977] , \zin[0][976] , \zin[0][975] , 
        \zin[0][974] , \zin[0][973] , \zin[0][972] , \zin[0][971] , 
        \zin[0][970] , \zin[0][969] , \zin[0][968] , \zin[0][967] , 
        \zin[0][966] , \zin[0][965] , \zin[0][964] , \zin[0][963] , 
        \zin[0][962] , \zin[0][961] , \zin[0][960] , \zin[0][959] , 
        \zin[0][958] , \zin[0][957] , \zin[0][956] , \zin[0][955] , 
        \zin[0][954] , \zin[0][953] , \zin[0][952] , \zin[0][951] , 
        \zin[0][950] , \zin[0][949] , \zin[0][948] , \zin[0][947] , 
        \zin[0][946] , \zin[0][945] , \zin[0][944] , \zin[0][943] , 
        \zin[0][942] , \zin[0][941] , \zin[0][940] , \zin[0][939] , 
        \zin[0][938] , \zin[0][937] , \zin[0][936] , \zin[0][935] , 
        \zin[0][934] , \zin[0][933] , \zin[0][932] , \zin[0][931] , 
        \zin[0][930] , \zin[0][929] , \zin[0][928] , \zin[0][927] , 
        \zin[0][926] , \zin[0][925] , \zin[0][924] , \zin[0][923] , 
        \zin[0][922] , \zin[0][921] , \zin[0][920] , \zin[0][919] , 
        \zin[0][918] , \zin[0][917] , \zin[0][916] , \zin[0][915] , 
        \zin[0][914] , \zin[0][913] , \zin[0][912] , \zin[0][911] , 
        \zin[0][910] , \zin[0][909] , \zin[0][908] , \zin[0][907] , 
        \zin[0][906] , \zin[0][905] , \zin[0][904] , \zin[0][903] , 
        \zin[0][902] , \zin[0][901] , \zin[0][900] , \zin[0][899] , 
        \zin[0][898] , \zin[0][897] , \zin[0][896] , \zin[0][895] , 
        \zin[0][894] , \zin[0][893] , \zin[0][892] , \zin[0][891] , 
        \zin[0][890] , \zin[0][889] , \zin[0][888] , \zin[0][887] , 
        \zin[0][886] , \zin[0][885] , \zin[0][884] , \zin[0][883] , 
        \zin[0][882] , \zin[0][881] , \zin[0][880] , \zin[0][879] , 
        \zin[0][878] , \zin[0][877] , \zin[0][876] , \zin[0][875] , 
        \zin[0][874] , \zin[0][873] , \zin[0][872] , \zin[0][871] , 
        \zin[0][870] , \zin[0][869] , \zin[0][868] , \zin[0][867] , 
        \zin[0][866] , \zin[0][865] , \zin[0][864] , \zin[0][863] , 
        \zin[0][862] , \zin[0][861] , \zin[0][860] , \zin[0][859] , 
        \zin[0][858] , \zin[0][857] , \zin[0][856] , \zin[0][855] , 
        \zin[0][854] , \zin[0][853] , \zin[0][852] , \zin[0][851] , 
        \zin[0][850] , \zin[0][849] , \zin[0][848] , \zin[0][847] , 
        \zin[0][846] , \zin[0][845] , \zin[0][844] , \zin[0][843] , 
        \zin[0][842] , \zin[0][841] , \zin[0][840] , \zin[0][839] , 
        \zin[0][838] , \zin[0][837] , \zin[0][836] , \zin[0][835] , 
        \zin[0][834] , \zin[0][833] , \zin[0][832] , \zin[0][831] , 
        \zin[0][830] , \zin[0][829] , \zin[0][828] , \zin[0][827] , 
        \zin[0][826] , \zin[0][825] , \zin[0][824] , \zin[0][823] , 
        \zin[0][822] , \zin[0][821] , \zin[0][820] , \zin[0][819] , 
        \zin[0][818] , \zin[0][817] , \zin[0][816] , \zin[0][815] , 
        \zin[0][814] , \zin[0][813] , \zin[0][812] , \zin[0][811] , 
        \zin[0][810] , \zin[0][809] , \zin[0][808] , \zin[0][807] , 
        \zin[0][806] , \zin[0][805] , \zin[0][804] , \zin[0][803] , 
        \zin[0][802] , \zin[0][801] , \zin[0][800] , \zin[0][799] , 
        \zin[0][798] , \zin[0][797] , \zin[0][796] , \zin[0][795] , 
        \zin[0][794] , \zin[0][793] , \zin[0][792] , \zin[0][791] , 
        \zin[0][790] , \zin[0][789] , \zin[0][788] , \zin[0][787] , 
        \zin[0][786] , \zin[0][785] , \zin[0][784] , \zin[0][783] , 
        \zin[0][782] , \zin[0][781] , \zin[0][780] , \zin[0][779] , 
        \zin[0][778] , \zin[0][777] , \zin[0][776] , \zin[0][775] , 
        \zin[0][774] , \zin[0][773] , \zin[0][772] , \zin[0][771] , 
        \zin[0][770] , \zin[0][769] , \zin[0][768] , \zin[0][767] , 
        \zin[0][766] , \zin[0][765] , \zin[0][764] , \zin[0][763] , 
        \zin[0][762] , \zin[0][761] , \zin[0][760] , \zin[0][759] , 
        \zin[0][758] , \zin[0][757] , \zin[0][756] , \zin[0][755] , 
        \zin[0][754] , \zin[0][753] , \zin[0][752] , \zin[0][751] , 
        \zin[0][750] , \zin[0][749] , \zin[0][748] , \zin[0][747] , 
        \zin[0][746] , \zin[0][745] , \zin[0][744] , \zin[0][743] , 
        \zin[0][742] , \zin[0][741] , \zin[0][740] , \zin[0][739] , 
        \zin[0][738] , \zin[0][737] , \zin[0][736] , \zin[0][735] , 
        \zin[0][734] , \zin[0][733] , \zin[0][732] , \zin[0][731] , 
        \zin[0][730] , \zin[0][729] , \zin[0][728] , \zin[0][727] , 
        \zin[0][726] , \zin[0][725] , \zin[0][724] , \zin[0][723] , 
        \zin[0][722] , \zin[0][721] , \zin[0][720] , \zin[0][719] , 
        \zin[0][718] , \zin[0][717] , \zin[0][716] , \zin[0][715] , 
        \zin[0][714] , \zin[0][713] , \zin[0][712] , \zin[0][711] , 
        \zin[0][710] , \zin[0][709] , \zin[0][708] , \zin[0][707] , 
        \zin[0][706] , \zin[0][705] , \zin[0][704] , \zin[0][703] , 
        \zin[0][702] , \zin[0][701] , \zin[0][700] , \zin[0][699] , 
        \zin[0][698] , \zin[0][697] , \zin[0][696] , \zin[0][695] , 
        \zin[0][694] , \zin[0][693] , \zin[0][692] , \zin[0][691] , 
        \zin[0][690] , \zin[0][689] , \zin[0][688] , \zin[0][687] , 
        \zin[0][686] , \zin[0][685] , \zin[0][684] , \zin[0][683] , 
        \zin[0][682] , \zin[0][681] , \zin[0][680] , \zin[0][679] , 
        \zin[0][678] , \zin[0][677] , \zin[0][676] , \zin[0][675] , 
        \zin[0][674] , \zin[0][673] , \zin[0][672] , \zin[0][671] , 
        \zin[0][670] , \zin[0][669] , \zin[0][668] , \zin[0][667] , 
        \zin[0][666] , \zin[0][665] , \zin[0][664] , \zin[0][663] , 
        \zin[0][662] , \zin[0][661] , \zin[0][660] , \zin[0][659] , 
        \zin[0][658] , \zin[0][657] , \zin[0][656] , \zin[0][655] , 
        \zin[0][654] , \zin[0][653] , \zin[0][652] , \zin[0][651] , 
        \zin[0][650] , \zin[0][649] , \zin[0][648] , \zin[0][647] , 
        \zin[0][646] , \zin[0][645] , \zin[0][644] , \zin[0][643] , 
        \zin[0][642] , \zin[0][641] , \zin[0][640] , \zin[0][639] , 
        \zin[0][638] , \zin[0][637] , \zin[0][636] , \zin[0][635] , 
        \zin[0][634] , \zin[0][633] , \zin[0][632] , \zin[0][631] , 
        \zin[0][630] , \zin[0][629] , \zin[0][628] , \zin[0][627] , 
        \zin[0][626] , \zin[0][625] , \zin[0][624] , \zin[0][623] , 
        \zin[0][622] , \zin[0][621] , \zin[0][620] , \zin[0][619] , 
        \zin[0][618] , \zin[0][617] , \zin[0][616] , \zin[0][615] , 
        \zin[0][614] , \zin[0][613] , \zin[0][612] , \zin[0][611] , 
        \zin[0][610] , \zin[0][609] , \zin[0][608] , \zin[0][607] , 
        \zin[0][606] , \zin[0][605] , \zin[0][604] , \zin[0][603] , 
        \zin[0][602] , \zin[0][601] , \zin[0][600] , \zin[0][599] , 
        \zin[0][598] , \zin[0][597] , \zin[0][596] , \zin[0][595] , 
        \zin[0][594] , \zin[0][593] , \zin[0][592] , \zin[0][591] , 
        \zin[0][590] , \zin[0][589] , \zin[0][588] , \zin[0][587] , 
        \zin[0][586] , \zin[0][585] , \zin[0][584] , \zin[0][583] , 
        \zin[0][582] , \zin[0][581] , \zin[0][580] , \zin[0][579] , 
        \zin[0][578] , \zin[0][577] , \zin[0][576] , \zin[0][575] , 
        \zin[0][574] , \zin[0][573] , \zin[0][572] , \zin[0][571] , 
        \zin[0][570] , \zin[0][569] , \zin[0][568] , \zin[0][567] , 
        \zin[0][566] , \zin[0][565] , \zin[0][564] , \zin[0][563] , 
        \zin[0][562] , \zin[0][561] , \zin[0][560] , \zin[0][559] , 
        \zin[0][558] , \zin[0][557] , \zin[0][556] , \zin[0][555] , 
        \zin[0][554] , \zin[0][553] , \zin[0][552] , \zin[0][551] , 
        \zin[0][550] , \zin[0][549] , \zin[0][548] , \zin[0][547] , 
        \zin[0][546] , \zin[0][545] , \zin[0][544] , \zin[0][543] , 
        \zin[0][542] , \zin[0][541] , \zin[0][540] , \zin[0][539] , 
        \zin[0][538] , \zin[0][537] , \zin[0][536] , \zin[0][535] , 
        \zin[0][534] , \zin[0][533] , \zin[0][532] , \zin[0][531] , 
        \zin[0][530] , \zin[0][529] , \zin[0][528] , \zin[0][527] , 
        \zin[0][526] , \zin[0][525] , \zin[0][524] , \zin[0][523] , 
        \zin[0][522] , \zin[0][521] , \zin[0][520] , \zin[0][519] , 
        \zin[0][518] , \zin[0][517] , \zin[0][516] , \zin[0][515] , 
        \zin[0][514] , \zin[0][513] , \zin[0][512] , \zin[0][511] , 
        \zin[0][510] , \zin[0][509] , \zin[0][508] , \zin[0][507] , 
        \zin[0][506] , \zin[0][505] , \zin[0][504] , \zin[0][503] , 
        \zin[0][502] , \zin[0][501] , \zin[0][500] , \zin[0][499] , 
        \zin[0][498] , \zin[0][497] , \zin[0][496] , \zin[0][495] , 
        \zin[0][494] , \zin[0][493] , \zin[0][492] , \zin[0][491] , 
        \zin[0][490] , \zin[0][489] , \zin[0][488] , \zin[0][487] , 
        \zin[0][486] , \zin[0][485] , \zin[0][484] , \zin[0][483] , 
        \zin[0][482] , \zin[0][481] , \zin[0][480] , \zin[0][479] , 
        \zin[0][478] , \zin[0][477] , \zin[0][476] , \zin[0][475] , 
        \zin[0][474] , \zin[0][473] , \zin[0][472] , \zin[0][471] , 
        \zin[0][470] , \zin[0][469] , \zin[0][468] , \zin[0][467] , 
        \zin[0][466] , \zin[0][465] , \zin[0][464] , \zin[0][463] , 
        \zin[0][462] , \zin[0][461] , \zin[0][460] , \zin[0][459] , 
        \zin[0][458] , \zin[0][457] , \zin[0][456] , \zin[0][455] , 
        \zin[0][454] , \zin[0][453] , \zin[0][452] , \zin[0][451] , 
        \zin[0][450] , \zin[0][449] , \zin[0][448] , \zin[0][447] , 
        \zin[0][446] , \zin[0][445] , \zin[0][444] , \zin[0][443] , 
        \zin[0][442] , \zin[0][441] , \zin[0][440] , \zin[0][439] , 
        \zin[0][438] , \zin[0][437] , \zin[0][436] , \zin[0][435] , 
        \zin[0][434] , \zin[0][433] , \zin[0][432] , \zin[0][431] , 
        \zin[0][430] , \zin[0][429] , \zin[0][428] , \zin[0][427] , 
        \zin[0][426] , \zin[0][425] , \zin[0][424] , \zin[0][423] , 
        \zin[0][422] , \zin[0][421] , \zin[0][420] , \zin[0][419] , 
        \zin[0][418] , \zin[0][417] , \zin[0][416] , \zin[0][415] , 
        \zin[0][414] , \zin[0][413] , \zin[0][412] , \zin[0][411] , 
        \zin[0][410] , \zin[0][409] , \zin[0][408] , \zin[0][407] , 
        \zin[0][406] , \zin[0][405] , \zin[0][404] , \zin[0][403] , 
        \zin[0][402] , \zin[0][401] , \zin[0][400] , \zin[0][399] , 
        \zin[0][398] , \zin[0][397] , \zin[0][396] , \zin[0][395] , 
        \zin[0][394] , \zin[0][393] , \zin[0][392] , \zin[0][391] , 
        \zin[0][390] , \zin[0][389] , \zin[0][388] , \zin[0][387] , 
        \zin[0][386] , \zin[0][385] , \zin[0][384] , \zin[0][383] , 
        \zin[0][382] , \zin[0][381] , \zin[0][380] , \zin[0][379] , 
        \zin[0][378] , \zin[0][377] , \zin[0][376] , \zin[0][375] , 
        \zin[0][374] , \zin[0][373] , \zin[0][372] , \zin[0][371] , 
        \zin[0][370] , \zin[0][369] , \zin[0][368] , \zin[0][367] , 
        \zin[0][366] , \zin[0][365] , \zin[0][364] , \zin[0][363] , 
        \zin[0][362] , \zin[0][361] , \zin[0][360] , \zin[0][359] , 
        \zin[0][358] , \zin[0][357] , \zin[0][356] , \zin[0][355] , 
        \zin[0][354] , \zin[0][353] , \zin[0][352] , \zin[0][351] , 
        \zin[0][350] , \zin[0][349] , \zin[0][348] , \zin[0][347] , 
        \zin[0][346] , \zin[0][345] , \zin[0][344] , \zin[0][343] , 
        \zin[0][342] , \zin[0][341] , \zin[0][340] , \zin[0][339] , 
        \zin[0][338] , \zin[0][337] , \zin[0][336] , \zin[0][335] , 
        \zin[0][334] , \zin[0][333] , \zin[0][332] , \zin[0][331] , 
        \zin[0][330] , \zin[0][329] , \zin[0][328] , \zin[0][327] , 
        \zin[0][326] , \zin[0][325] , \zin[0][324] , \zin[0][323] , 
        \zin[0][322] , \zin[0][321] , \zin[0][320] , \zin[0][319] , 
        \zin[0][318] , \zin[0][317] , \zin[0][316] , \zin[0][315] , 
        \zin[0][314] , \zin[0][313] , \zin[0][312] , \zin[0][311] , 
        \zin[0][310] , \zin[0][309] , \zin[0][308] , \zin[0][307] , 
        \zin[0][306] , \zin[0][305] , \zin[0][304] , \zin[0][303] , 
        \zin[0][302] , \zin[0][301] , \zin[0][300] , \zin[0][299] , 
        \zin[0][298] , \zin[0][297] , \zin[0][296] , \zin[0][295] , 
        \zin[0][294] , \zin[0][293] , \zin[0][292] , \zin[0][291] , 
        \zin[0][290] , \zin[0][289] , \zin[0][288] , \zin[0][287] , 
        \zin[0][286] , \zin[0][285] , \zin[0][284] , \zin[0][283] , 
        \zin[0][282] , \zin[0][281] , \zin[0][280] , \zin[0][279] , 
        \zin[0][278] , \zin[0][277] , \zin[0][276] , \zin[0][275] , 
        \zin[0][274] , \zin[0][273] , \zin[0][272] , \zin[0][271] , 
        \zin[0][270] , \zin[0][269] , \zin[0][268] , \zin[0][267] , 
        \zin[0][266] , \zin[0][265] , \zin[0][264] , \zin[0][263] , 
        \zin[0][262] , \zin[0][261] , \zin[0][260] , \zin[0][259] , 
        \zin[0][258] , \zin[0][257] , \zin[0][256] , \zin[0][255] , 
        \zin[0][254] , \zin[0][253] , \zin[0][252] , \zin[0][251] , 
        \zin[0][250] , \zin[0][249] , \zin[0][248] , \zin[0][247] , 
        \zin[0][246] , \zin[0][245] , \zin[0][244] , \zin[0][243] , 
        \zin[0][242] , \zin[0][241] , \zin[0][240] , \zin[0][239] , 
        \zin[0][238] , \zin[0][237] , \zin[0][236] , \zin[0][235] , 
        \zin[0][234] , \zin[0][233] , \zin[0][232] , \zin[0][231] , 
        \zin[0][230] , \zin[0][229] , \zin[0][228] , \zin[0][227] , 
        \zin[0][226] , \zin[0][225] , \zin[0][224] , \zin[0][223] , 
        \zin[0][222] , \zin[0][221] , \zin[0][220] , \zin[0][219] , 
        \zin[0][218] , \zin[0][217] , \zin[0][216] , \zin[0][215] , 
        \zin[0][214] , \zin[0][213] , \zin[0][212] , \zin[0][211] , 
        \zin[0][210] , \zin[0][209] , \zin[0][208] , \zin[0][207] , 
        \zin[0][206] , \zin[0][205] , \zin[0][204] , \zin[0][203] , 
        \zin[0][202] , \zin[0][201] , \zin[0][200] , \zin[0][199] , 
        \zin[0][198] , \zin[0][197] , \zin[0][196] , \zin[0][195] , 
        \zin[0][194] , \zin[0][193] , \zin[0][192] , \zin[0][191] , 
        \zin[0][190] , \zin[0][189] , \zin[0][188] , \zin[0][187] , 
        \zin[0][186] , \zin[0][185] , \zin[0][184] , \zin[0][183] , 
        \zin[0][182] , \zin[0][181] , \zin[0][180] , \zin[0][179] , 
        \zin[0][178] , \zin[0][177] , \zin[0][176] , \zin[0][175] , 
        \zin[0][174] , \zin[0][173] , \zin[0][172] , \zin[0][171] , 
        \zin[0][170] , \zin[0][169] , \zin[0][168] , \zin[0][167] , 
        \zin[0][166] , \zin[0][165] , \zin[0][164] , \zin[0][163] , 
        \zin[0][162] , \zin[0][161] , \zin[0][160] , \zin[0][159] , 
        \zin[0][158] , \zin[0][157] , \zin[0][156] , \zin[0][155] , 
        \zin[0][154] , \zin[0][153] , \zin[0][152] , \zin[0][151] , 
        \zin[0][150] , \zin[0][149] , \zin[0][148] , \zin[0][147] , 
        \zin[0][146] , \zin[0][145] , \zin[0][144] , \zin[0][143] , 
        \zin[0][142] , \zin[0][141] , \zin[0][140] , \zin[0][139] , 
        \zin[0][138] , \zin[0][137] , \zin[0][136] , \zin[0][135] , 
        \zin[0][134] , \zin[0][133] , \zin[0][132] , \zin[0][131] , 
        \zin[0][130] , \zin[0][129] , \zin[0][128] , \zin[0][127] , 
        \zin[0][126] , \zin[0][125] , \zin[0][124] , \zin[0][123] , 
        \zin[0][122] , \zin[0][121] , \zin[0][120] , \zin[0][119] , 
        \zin[0][118] , \zin[0][117] , \zin[0][116] , \zin[0][115] , 
        \zin[0][114] , \zin[0][113] , \zin[0][112] , \zin[0][111] , 
        \zin[0][110] , \zin[0][109] , \zin[0][108] , \zin[0][107] , 
        \zin[0][106] , \zin[0][105] , \zin[0][104] , \zin[0][103] , 
        \zin[0][102] , \zin[0][101] , \zin[0][100] , \zin[0][99] , 
        \zin[0][98] , \zin[0][97] , \zin[0][96] , \zin[0][95] , \zin[0][94] , 
        \zin[0][93] , \zin[0][92] , \zin[0][91] , \zin[0][90] , \zin[0][89] , 
        \zin[0][88] , \zin[0][87] , \zin[0][86] , \zin[0][85] , \zin[0][84] , 
        \zin[0][83] , \zin[0][82] , \zin[0][81] , \zin[0][80] , \zin[0][79] , 
        \zin[0][78] , \zin[0][77] , \zin[0][76] , \zin[0][75] , \zin[0][74] , 
        \zin[0][73] , \zin[0][72] , \zin[0][71] , \zin[0][70] , \zin[0][69] , 
        \zin[0][68] , \zin[0][67] , \zin[0][66] , \zin[0][65] , \zin[0][64] , 
        \zin[0][63] , \zin[0][62] , \zin[0][61] , \zin[0][60] , \zin[0][59] , 
        \zin[0][58] , \zin[0][57] , \zin[0][56] , \zin[0][55] , \zin[0][54] , 
        \zin[0][53] , \zin[0][52] , \zin[0][51] , \zin[0][50] , \zin[0][49] , 
        \zin[0][48] , \zin[0][47] , \zin[0][46] , \zin[0][45] , \zin[0][44] , 
        \zin[0][43] , \zin[0][42] , \zin[0][41] , \zin[0][40] , \zin[0][39] , 
        \zin[0][38] , \zin[0][37] , \zin[0][36] , \zin[0][35] , \zin[0][34] , 
        \zin[0][33] , \zin[0][32] , \zin[0][31] , \zin[0][30] , \zin[0][29] , 
        \zin[0][28] , \zin[0][27] , \zin[0][26] , \zin[0][25] , \zin[0][24] , 
        \zin[0][23] , \zin[0][22] , \zin[0][21] , \zin[0][20] , \zin[0][19] , 
        \zin[0][18] , \zin[0][17] , \zin[0][16] , \zin[0][15] , \zin[0][14] , 
        \zin[0][13] , \zin[0][12] , \zin[0][11] , \zin[0][10] , \zin[0][9] , 
        \zin[0][8] , \zin[0][7] , \zin[0][6] , \zin[0][5] , \zin[0][4] , 
        \zin[0][3] , \zin[0][2] , \zin[0][1] , \zin[0][0] }), .zout({
        \zout[0][1025] , \zout[0][1024] , o}) );
  ANDN U3 ( .B(zreg[9]), .A(start), .Z(\zin[0][9] ) );
  ANDN U4 ( .B(zreg[99]), .A(start), .Z(\zin[0][99] ) );
  ANDN U5 ( .B(zreg[999]), .A(start), .Z(\zin[0][999] ) );
  ANDN U6 ( .B(zreg[998]), .A(start), .Z(\zin[0][998] ) );
  ANDN U7 ( .B(zreg[997]), .A(start), .Z(\zin[0][997] ) );
  ANDN U8 ( .B(zreg[996]), .A(start), .Z(\zin[0][996] ) );
  ANDN U9 ( .B(zreg[995]), .A(start), .Z(\zin[0][995] ) );
  ANDN U10 ( .B(zreg[994]), .A(start), .Z(\zin[0][994] ) );
  ANDN U11 ( .B(zreg[993]), .A(start), .Z(\zin[0][993] ) );
  ANDN U12 ( .B(zreg[992]), .A(start), .Z(\zin[0][992] ) );
  ANDN U13 ( .B(zreg[991]), .A(start), .Z(\zin[0][991] ) );
  ANDN U14 ( .B(zreg[990]), .A(start), .Z(\zin[0][990] ) );
  ANDN U15 ( .B(zreg[98]), .A(start), .Z(\zin[0][98] ) );
  ANDN U16 ( .B(zreg[989]), .A(start), .Z(\zin[0][989] ) );
  ANDN U17 ( .B(zreg[988]), .A(start), .Z(\zin[0][988] ) );
  ANDN U18 ( .B(zreg[987]), .A(start), .Z(\zin[0][987] ) );
  ANDN U19 ( .B(zreg[986]), .A(start), .Z(\zin[0][986] ) );
  ANDN U20 ( .B(zreg[985]), .A(start), .Z(\zin[0][985] ) );
  ANDN U21 ( .B(zreg[984]), .A(start), .Z(\zin[0][984] ) );
  ANDN U22 ( .B(zreg[983]), .A(start), .Z(\zin[0][983] ) );
  ANDN U23 ( .B(zreg[982]), .A(start), .Z(\zin[0][982] ) );
  ANDN U24 ( .B(zreg[981]), .A(start), .Z(\zin[0][981] ) );
  ANDN U25 ( .B(zreg[980]), .A(start), .Z(\zin[0][980] ) );
  ANDN U26 ( .B(zreg[97]), .A(start), .Z(\zin[0][97] ) );
  ANDN U27 ( .B(zreg[979]), .A(start), .Z(\zin[0][979] ) );
  ANDN U28 ( .B(zreg[978]), .A(start), .Z(\zin[0][978] ) );
  ANDN U29 ( .B(zreg[977]), .A(start), .Z(\zin[0][977] ) );
  ANDN U30 ( .B(zreg[976]), .A(start), .Z(\zin[0][976] ) );
  ANDN U31 ( .B(zreg[975]), .A(start), .Z(\zin[0][975] ) );
  ANDN U32 ( .B(zreg[974]), .A(start), .Z(\zin[0][974] ) );
  ANDN U33 ( .B(zreg[973]), .A(start), .Z(\zin[0][973] ) );
  ANDN U34 ( .B(zreg[972]), .A(start), .Z(\zin[0][972] ) );
  ANDN U35 ( .B(zreg[971]), .A(start), .Z(\zin[0][971] ) );
  ANDN U36 ( .B(zreg[970]), .A(start), .Z(\zin[0][970] ) );
  ANDN U37 ( .B(zreg[96]), .A(start), .Z(\zin[0][96] ) );
  ANDN U38 ( .B(zreg[969]), .A(start), .Z(\zin[0][969] ) );
  ANDN U39 ( .B(zreg[968]), .A(start), .Z(\zin[0][968] ) );
  ANDN U40 ( .B(zreg[967]), .A(start), .Z(\zin[0][967] ) );
  ANDN U41 ( .B(zreg[966]), .A(start), .Z(\zin[0][966] ) );
  ANDN U42 ( .B(zreg[965]), .A(start), .Z(\zin[0][965] ) );
  ANDN U43 ( .B(zreg[964]), .A(start), .Z(\zin[0][964] ) );
  ANDN U44 ( .B(zreg[963]), .A(start), .Z(\zin[0][963] ) );
  ANDN U45 ( .B(zreg[962]), .A(start), .Z(\zin[0][962] ) );
  ANDN U46 ( .B(zreg[961]), .A(start), .Z(\zin[0][961] ) );
  ANDN U47 ( .B(zreg[960]), .A(start), .Z(\zin[0][960] ) );
  ANDN U48 ( .B(zreg[95]), .A(start), .Z(\zin[0][95] ) );
  ANDN U49 ( .B(zreg[959]), .A(start), .Z(\zin[0][959] ) );
  ANDN U50 ( .B(zreg[958]), .A(start), .Z(\zin[0][958] ) );
  ANDN U51 ( .B(zreg[957]), .A(start), .Z(\zin[0][957] ) );
  ANDN U52 ( .B(zreg[956]), .A(start), .Z(\zin[0][956] ) );
  ANDN U53 ( .B(zreg[955]), .A(start), .Z(\zin[0][955] ) );
  ANDN U54 ( .B(zreg[954]), .A(start), .Z(\zin[0][954] ) );
  ANDN U55 ( .B(zreg[953]), .A(start), .Z(\zin[0][953] ) );
  ANDN U56 ( .B(zreg[952]), .A(start), .Z(\zin[0][952] ) );
  ANDN U57 ( .B(zreg[951]), .A(start), .Z(\zin[0][951] ) );
  ANDN U58 ( .B(zreg[950]), .A(start), .Z(\zin[0][950] ) );
  ANDN U59 ( .B(zreg[94]), .A(start), .Z(\zin[0][94] ) );
  ANDN U60 ( .B(zreg[949]), .A(start), .Z(\zin[0][949] ) );
  ANDN U61 ( .B(zreg[948]), .A(start), .Z(\zin[0][948] ) );
  ANDN U62 ( .B(zreg[947]), .A(start), .Z(\zin[0][947] ) );
  ANDN U63 ( .B(zreg[946]), .A(start), .Z(\zin[0][946] ) );
  ANDN U64 ( .B(zreg[945]), .A(start), .Z(\zin[0][945] ) );
  ANDN U65 ( .B(zreg[944]), .A(start), .Z(\zin[0][944] ) );
  ANDN U66 ( .B(zreg[943]), .A(start), .Z(\zin[0][943] ) );
  ANDN U67 ( .B(zreg[942]), .A(start), .Z(\zin[0][942] ) );
  ANDN U68 ( .B(zreg[941]), .A(start), .Z(\zin[0][941] ) );
  ANDN U69 ( .B(zreg[940]), .A(start), .Z(\zin[0][940] ) );
  ANDN U70 ( .B(zreg[93]), .A(start), .Z(\zin[0][93] ) );
  ANDN U71 ( .B(zreg[939]), .A(start), .Z(\zin[0][939] ) );
  ANDN U72 ( .B(zreg[938]), .A(start), .Z(\zin[0][938] ) );
  ANDN U73 ( .B(zreg[937]), .A(start), .Z(\zin[0][937] ) );
  ANDN U74 ( .B(zreg[936]), .A(start), .Z(\zin[0][936] ) );
  ANDN U75 ( .B(zreg[935]), .A(start), .Z(\zin[0][935] ) );
  ANDN U76 ( .B(zreg[934]), .A(start), .Z(\zin[0][934] ) );
  ANDN U77 ( .B(zreg[933]), .A(start), .Z(\zin[0][933] ) );
  ANDN U78 ( .B(zreg[932]), .A(start), .Z(\zin[0][932] ) );
  ANDN U79 ( .B(zreg[931]), .A(start), .Z(\zin[0][931] ) );
  ANDN U80 ( .B(zreg[930]), .A(start), .Z(\zin[0][930] ) );
  ANDN U81 ( .B(zreg[92]), .A(start), .Z(\zin[0][92] ) );
  ANDN U82 ( .B(zreg[929]), .A(start), .Z(\zin[0][929] ) );
  ANDN U83 ( .B(zreg[928]), .A(start), .Z(\zin[0][928] ) );
  ANDN U84 ( .B(zreg[927]), .A(start), .Z(\zin[0][927] ) );
  ANDN U85 ( .B(zreg[926]), .A(start), .Z(\zin[0][926] ) );
  ANDN U86 ( .B(zreg[925]), .A(start), .Z(\zin[0][925] ) );
  ANDN U87 ( .B(zreg[924]), .A(start), .Z(\zin[0][924] ) );
  ANDN U88 ( .B(zreg[923]), .A(start), .Z(\zin[0][923] ) );
  ANDN U89 ( .B(zreg[922]), .A(start), .Z(\zin[0][922] ) );
  ANDN U90 ( .B(zreg[921]), .A(start), .Z(\zin[0][921] ) );
  ANDN U91 ( .B(zreg[920]), .A(start), .Z(\zin[0][920] ) );
  ANDN U92 ( .B(zreg[91]), .A(start), .Z(\zin[0][91] ) );
  ANDN U93 ( .B(zreg[919]), .A(start), .Z(\zin[0][919] ) );
  ANDN U94 ( .B(zreg[918]), .A(start), .Z(\zin[0][918] ) );
  ANDN U95 ( .B(zreg[917]), .A(start), .Z(\zin[0][917] ) );
  ANDN U96 ( .B(zreg[916]), .A(start), .Z(\zin[0][916] ) );
  ANDN U97 ( .B(zreg[915]), .A(start), .Z(\zin[0][915] ) );
  ANDN U98 ( .B(zreg[914]), .A(start), .Z(\zin[0][914] ) );
  ANDN U99 ( .B(zreg[913]), .A(start), .Z(\zin[0][913] ) );
  ANDN U100 ( .B(zreg[912]), .A(start), .Z(\zin[0][912] ) );
  ANDN U101 ( .B(zreg[911]), .A(start), .Z(\zin[0][911] ) );
  ANDN U102 ( .B(zreg[910]), .A(start), .Z(\zin[0][910] ) );
  ANDN U103 ( .B(zreg[90]), .A(start), .Z(\zin[0][90] ) );
  ANDN U104 ( .B(zreg[909]), .A(start), .Z(\zin[0][909] ) );
  ANDN U105 ( .B(zreg[908]), .A(start), .Z(\zin[0][908] ) );
  ANDN U106 ( .B(zreg[907]), .A(start), .Z(\zin[0][907] ) );
  ANDN U107 ( .B(zreg[906]), .A(start), .Z(\zin[0][906] ) );
  ANDN U108 ( .B(zreg[905]), .A(start), .Z(\zin[0][905] ) );
  ANDN U109 ( .B(zreg[904]), .A(start), .Z(\zin[0][904] ) );
  ANDN U110 ( .B(zreg[903]), .A(start), .Z(\zin[0][903] ) );
  ANDN U111 ( .B(zreg[902]), .A(start), .Z(\zin[0][902] ) );
  ANDN U112 ( .B(zreg[901]), .A(start), .Z(\zin[0][901] ) );
  ANDN U113 ( .B(zreg[900]), .A(start), .Z(\zin[0][900] ) );
  ANDN U114 ( .B(zreg[8]), .A(start), .Z(\zin[0][8] ) );
  ANDN U115 ( .B(zreg[89]), .A(start), .Z(\zin[0][89] ) );
  ANDN U116 ( .B(zreg[899]), .A(start), .Z(\zin[0][899] ) );
  ANDN U117 ( .B(zreg[898]), .A(start), .Z(\zin[0][898] ) );
  ANDN U118 ( .B(zreg[897]), .A(start), .Z(\zin[0][897] ) );
  ANDN U119 ( .B(zreg[896]), .A(start), .Z(\zin[0][896] ) );
  ANDN U120 ( .B(zreg[895]), .A(start), .Z(\zin[0][895] ) );
  ANDN U121 ( .B(zreg[894]), .A(start), .Z(\zin[0][894] ) );
  ANDN U122 ( .B(zreg[893]), .A(start), .Z(\zin[0][893] ) );
  ANDN U123 ( .B(zreg[892]), .A(start), .Z(\zin[0][892] ) );
  ANDN U124 ( .B(zreg[891]), .A(start), .Z(\zin[0][891] ) );
  ANDN U125 ( .B(zreg[890]), .A(start), .Z(\zin[0][890] ) );
  ANDN U126 ( .B(zreg[88]), .A(start), .Z(\zin[0][88] ) );
  ANDN U127 ( .B(zreg[889]), .A(start), .Z(\zin[0][889] ) );
  ANDN U128 ( .B(zreg[888]), .A(start), .Z(\zin[0][888] ) );
  ANDN U129 ( .B(zreg[887]), .A(start), .Z(\zin[0][887] ) );
  ANDN U130 ( .B(zreg[886]), .A(start), .Z(\zin[0][886] ) );
  ANDN U131 ( .B(zreg[885]), .A(start), .Z(\zin[0][885] ) );
  ANDN U132 ( .B(zreg[884]), .A(start), .Z(\zin[0][884] ) );
  ANDN U133 ( .B(zreg[883]), .A(start), .Z(\zin[0][883] ) );
  ANDN U134 ( .B(zreg[882]), .A(start), .Z(\zin[0][882] ) );
  ANDN U135 ( .B(zreg[881]), .A(start), .Z(\zin[0][881] ) );
  ANDN U136 ( .B(zreg[880]), .A(start), .Z(\zin[0][880] ) );
  ANDN U137 ( .B(zreg[87]), .A(start), .Z(\zin[0][87] ) );
  ANDN U138 ( .B(zreg[879]), .A(start), .Z(\zin[0][879] ) );
  ANDN U139 ( .B(zreg[878]), .A(start), .Z(\zin[0][878] ) );
  ANDN U140 ( .B(zreg[877]), .A(start), .Z(\zin[0][877] ) );
  ANDN U141 ( .B(zreg[876]), .A(start), .Z(\zin[0][876] ) );
  ANDN U142 ( .B(zreg[875]), .A(start), .Z(\zin[0][875] ) );
  ANDN U143 ( .B(zreg[874]), .A(start), .Z(\zin[0][874] ) );
  ANDN U144 ( .B(zreg[873]), .A(start), .Z(\zin[0][873] ) );
  ANDN U145 ( .B(zreg[872]), .A(start), .Z(\zin[0][872] ) );
  ANDN U146 ( .B(zreg[871]), .A(start), .Z(\zin[0][871] ) );
  ANDN U147 ( .B(zreg[870]), .A(start), .Z(\zin[0][870] ) );
  ANDN U148 ( .B(zreg[86]), .A(start), .Z(\zin[0][86] ) );
  ANDN U149 ( .B(zreg[869]), .A(start), .Z(\zin[0][869] ) );
  ANDN U150 ( .B(zreg[868]), .A(start), .Z(\zin[0][868] ) );
  ANDN U151 ( .B(zreg[867]), .A(start), .Z(\zin[0][867] ) );
  ANDN U152 ( .B(zreg[866]), .A(start), .Z(\zin[0][866] ) );
  ANDN U153 ( .B(zreg[865]), .A(start), .Z(\zin[0][865] ) );
  ANDN U154 ( .B(zreg[864]), .A(start), .Z(\zin[0][864] ) );
  ANDN U155 ( .B(zreg[863]), .A(start), .Z(\zin[0][863] ) );
  ANDN U156 ( .B(zreg[862]), .A(start), .Z(\zin[0][862] ) );
  ANDN U157 ( .B(zreg[861]), .A(start), .Z(\zin[0][861] ) );
  ANDN U158 ( .B(zreg[860]), .A(start), .Z(\zin[0][860] ) );
  ANDN U159 ( .B(zreg[85]), .A(start), .Z(\zin[0][85] ) );
  ANDN U160 ( .B(zreg[859]), .A(start), .Z(\zin[0][859] ) );
  ANDN U161 ( .B(zreg[858]), .A(start), .Z(\zin[0][858] ) );
  ANDN U162 ( .B(zreg[857]), .A(start), .Z(\zin[0][857] ) );
  ANDN U163 ( .B(zreg[856]), .A(start), .Z(\zin[0][856] ) );
  ANDN U164 ( .B(zreg[855]), .A(start), .Z(\zin[0][855] ) );
  ANDN U165 ( .B(zreg[854]), .A(start), .Z(\zin[0][854] ) );
  ANDN U166 ( .B(zreg[853]), .A(start), .Z(\zin[0][853] ) );
  ANDN U167 ( .B(zreg[852]), .A(start), .Z(\zin[0][852] ) );
  ANDN U168 ( .B(zreg[851]), .A(start), .Z(\zin[0][851] ) );
  ANDN U169 ( .B(zreg[850]), .A(start), .Z(\zin[0][850] ) );
  ANDN U170 ( .B(zreg[84]), .A(start), .Z(\zin[0][84] ) );
  ANDN U171 ( .B(zreg[849]), .A(start), .Z(\zin[0][849] ) );
  ANDN U172 ( .B(zreg[848]), .A(start), .Z(\zin[0][848] ) );
  ANDN U173 ( .B(zreg[847]), .A(start), .Z(\zin[0][847] ) );
  ANDN U174 ( .B(zreg[846]), .A(start), .Z(\zin[0][846] ) );
  ANDN U175 ( .B(zreg[845]), .A(start), .Z(\zin[0][845] ) );
  ANDN U176 ( .B(zreg[844]), .A(start), .Z(\zin[0][844] ) );
  ANDN U177 ( .B(zreg[843]), .A(start), .Z(\zin[0][843] ) );
  ANDN U178 ( .B(zreg[842]), .A(start), .Z(\zin[0][842] ) );
  ANDN U179 ( .B(zreg[841]), .A(start), .Z(\zin[0][841] ) );
  ANDN U180 ( .B(zreg[840]), .A(start), .Z(\zin[0][840] ) );
  ANDN U181 ( .B(zreg[83]), .A(start), .Z(\zin[0][83] ) );
  ANDN U182 ( .B(zreg[839]), .A(start), .Z(\zin[0][839] ) );
  ANDN U183 ( .B(zreg[838]), .A(start), .Z(\zin[0][838] ) );
  ANDN U184 ( .B(zreg[837]), .A(start), .Z(\zin[0][837] ) );
  ANDN U185 ( .B(zreg[836]), .A(start), .Z(\zin[0][836] ) );
  ANDN U186 ( .B(zreg[835]), .A(start), .Z(\zin[0][835] ) );
  ANDN U187 ( .B(zreg[834]), .A(start), .Z(\zin[0][834] ) );
  ANDN U188 ( .B(zreg[833]), .A(start), .Z(\zin[0][833] ) );
  ANDN U189 ( .B(zreg[832]), .A(start), .Z(\zin[0][832] ) );
  ANDN U190 ( .B(zreg[831]), .A(start), .Z(\zin[0][831] ) );
  ANDN U191 ( .B(zreg[830]), .A(start), .Z(\zin[0][830] ) );
  ANDN U192 ( .B(zreg[82]), .A(start), .Z(\zin[0][82] ) );
  ANDN U193 ( .B(zreg[829]), .A(start), .Z(\zin[0][829] ) );
  ANDN U194 ( .B(zreg[828]), .A(start), .Z(\zin[0][828] ) );
  ANDN U195 ( .B(zreg[827]), .A(start), .Z(\zin[0][827] ) );
  ANDN U196 ( .B(zreg[826]), .A(start), .Z(\zin[0][826] ) );
  ANDN U197 ( .B(zreg[825]), .A(start), .Z(\zin[0][825] ) );
  ANDN U198 ( .B(zreg[824]), .A(start), .Z(\zin[0][824] ) );
  ANDN U199 ( .B(zreg[823]), .A(start), .Z(\zin[0][823] ) );
  ANDN U200 ( .B(zreg[822]), .A(start), .Z(\zin[0][822] ) );
  ANDN U201 ( .B(zreg[821]), .A(start), .Z(\zin[0][821] ) );
  ANDN U202 ( .B(zreg[820]), .A(start), .Z(\zin[0][820] ) );
  ANDN U203 ( .B(zreg[81]), .A(start), .Z(\zin[0][81] ) );
  ANDN U204 ( .B(zreg[819]), .A(start), .Z(\zin[0][819] ) );
  ANDN U205 ( .B(zreg[818]), .A(start), .Z(\zin[0][818] ) );
  ANDN U206 ( .B(zreg[817]), .A(start), .Z(\zin[0][817] ) );
  ANDN U207 ( .B(zreg[816]), .A(start), .Z(\zin[0][816] ) );
  ANDN U208 ( .B(zreg[815]), .A(start), .Z(\zin[0][815] ) );
  ANDN U209 ( .B(zreg[814]), .A(start), .Z(\zin[0][814] ) );
  ANDN U210 ( .B(zreg[813]), .A(start), .Z(\zin[0][813] ) );
  ANDN U211 ( .B(zreg[812]), .A(start), .Z(\zin[0][812] ) );
  ANDN U212 ( .B(zreg[811]), .A(start), .Z(\zin[0][811] ) );
  ANDN U213 ( .B(zreg[810]), .A(start), .Z(\zin[0][810] ) );
  ANDN U214 ( .B(zreg[80]), .A(start), .Z(\zin[0][80] ) );
  ANDN U215 ( .B(zreg[809]), .A(start), .Z(\zin[0][809] ) );
  ANDN U216 ( .B(zreg[808]), .A(start), .Z(\zin[0][808] ) );
  ANDN U217 ( .B(zreg[807]), .A(start), .Z(\zin[0][807] ) );
  ANDN U218 ( .B(zreg[806]), .A(start), .Z(\zin[0][806] ) );
  ANDN U219 ( .B(zreg[805]), .A(start), .Z(\zin[0][805] ) );
  ANDN U220 ( .B(zreg[804]), .A(start), .Z(\zin[0][804] ) );
  ANDN U221 ( .B(zreg[803]), .A(start), .Z(\zin[0][803] ) );
  ANDN U222 ( .B(zreg[802]), .A(start), .Z(\zin[0][802] ) );
  ANDN U223 ( .B(zreg[801]), .A(start), .Z(\zin[0][801] ) );
  ANDN U224 ( .B(zreg[800]), .A(start), .Z(\zin[0][800] ) );
  ANDN U225 ( .B(zreg[7]), .A(start), .Z(\zin[0][7] ) );
  ANDN U226 ( .B(zreg[79]), .A(start), .Z(\zin[0][79] ) );
  ANDN U227 ( .B(zreg[799]), .A(start), .Z(\zin[0][799] ) );
  ANDN U228 ( .B(zreg[798]), .A(start), .Z(\zin[0][798] ) );
  ANDN U229 ( .B(zreg[797]), .A(start), .Z(\zin[0][797] ) );
  ANDN U230 ( .B(zreg[796]), .A(start), .Z(\zin[0][796] ) );
  ANDN U231 ( .B(zreg[795]), .A(start), .Z(\zin[0][795] ) );
  ANDN U232 ( .B(zreg[794]), .A(start), .Z(\zin[0][794] ) );
  ANDN U233 ( .B(zreg[793]), .A(start), .Z(\zin[0][793] ) );
  ANDN U234 ( .B(zreg[792]), .A(start), .Z(\zin[0][792] ) );
  ANDN U235 ( .B(zreg[791]), .A(start), .Z(\zin[0][791] ) );
  ANDN U236 ( .B(zreg[790]), .A(start), .Z(\zin[0][790] ) );
  ANDN U237 ( .B(zreg[78]), .A(start), .Z(\zin[0][78] ) );
  ANDN U238 ( .B(zreg[789]), .A(start), .Z(\zin[0][789] ) );
  ANDN U239 ( .B(zreg[788]), .A(start), .Z(\zin[0][788] ) );
  ANDN U240 ( .B(zreg[787]), .A(start), .Z(\zin[0][787] ) );
  ANDN U241 ( .B(zreg[786]), .A(start), .Z(\zin[0][786] ) );
  ANDN U242 ( .B(zreg[785]), .A(start), .Z(\zin[0][785] ) );
  ANDN U243 ( .B(zreg[784]), .A(start), .Z(\zin[0][784] ) );
  ANDN U244 ( .B(zreg[783]), .A(start), .Z(\zin[0][783] ) );
  ANDN U245 ( .B(zreg[782]), .A(start), .Z(\zin[0][782] ) );
  ANDN U246 ( .B(zreg[781]), .A(start), .Z(\zin[0][781] ) );
  ANDN U247 ( .B(zreg[780]), .A(start), .Z(\zin[0][780] ) );
  ANDN U248 ( .B(zreg[77]), .A(start), .Z(\zin[0][77] ) );
  ANDN U249 ( .B(zreg[779]), .A(start), .Z(\zin[0][779] ) );
  ANDN U250 ( .B(zreg[778]), .A(start), .Z(\zin[0][778] ) );
  ANDN U251 ( .B(zreg[777]), .A(start), .Z(\zin[0][777] ) );
  ANDN U252 ( .B(zreg[776]), .A(start), .Z(\zin[0][776] ) );
  ANDN U253 ( .B(zreg[775]), .A(start), .Z(\zin[0][775] ) );
  ANDN U254 ( .B(zreg[774]), .A(start), .Z(\zin[0][774] ) );
  ANDN U255 ( .B(zreg[773]), .A(start), .Z(\zin[0][773] ) );
  ANDN U256 ( .B(zreg[772]), .A(start), .Z(\zin[0][772] ) );
  ANDN U257 ( .B(zreg[771]), .A(start), .Z(\zin[0][771] ) );
  ANDN U258 ( .B(zreg[770]), .A(start), .Z(\zin[0][770] ) );
  ANDN U259 ( .B(zreg[76]), .A(start), .Z(\zin[0][76] ) );
  ANDN U260 ( .B(zreg[769]), .A(start), .Z(\zin[0][769] ) );
  ANDN U261 ( .B(zreg[768]), .A(start), .Z(\zin[0][768] ) );
  ANDN U262 ( .B(zreg[767]), .A(start), .Z(\zin[0][767] ) );
  ANDN U263 ( .B(zreg[766]), .A(start), .Z(\zin[0][766] ) );
  ANDN U264 ( .B(zreg[765]), .A(start), .Z(\zin[0][765] ) );
  ANDN U265 ( .B(zreg[764]), .A(start), .Z(\zin[0][764] ) );
  ANDN U266 ( .B(zreg[763]), .A(start), .Z(\zin[0][763] ) );
  ANDN U267 ( .B(zreg[762]), .A(start), .Z(\zin[0][762] ) );
  ANDN U268 ( .B(zreg[761]), .A(start), .Z(\zin[0][761] ) );
  ANDN U269 ( .B(zreg[760]), .A(start), .Z(\zin[0][760] ) );
  ANDN U270 ( .B(zreg[75]), .A(start), .Z(\zin[0][75] ) );
  ANDN U271 ( .B(zreg[759]), .A(start), .Z(\zin[0][759] ) );
  ANDN U272 ( .B(zreg[758]), .A(start), .Z(\zin[0][758] ) );
  ANDN U273 ( .B(zreg[757]), .A(start), .Z(\zin[0][757] ) );
  ANDN U274 ( .B(zreg[756]), .A(start), .Z(\zin[0][756] ) );
  ANDN U275 ( .B(zreg[755]), .A(start), .Z(\zin[0][755] ) );
  ANDN U276 ( .B(zreg[754]), .A(start), .Z(\zin[0][754] ) );
  ANDN U277 ( .B(zreg[753]), .A(start), .Z(\zin[0][753] ) );
  ANDN U278 ( .B(zreg[752]), .A(start), .Z(\zin[0][752] ) );
  ANDN U279 ( .B(zreg[751]), .A(start), .Z(\zin[0][751] ) );
  ANDN U280 ( .B(zreg[750]), .A(start), .Z(\zin[0][750] ) );
  ANDN U281 ( .B(zreg[74]), .A(start), .Z(\zin[0][74] ) );
  ANDN U282 ( .B(zreg[749]), .A(start), .Z(\zin[0][749] ) );
  ANDN U283 ( .B(zreg[748]), .A(start), .Z(\zin[0][748] ) );
  ANDN U284 ( .B(zreg[747]), .A(start), .Z(\zin[0][747] ) );
  ANDN U285 ( .B(zreg[746]), .A(start), .Z(\zin[0][746] ) );
  ANDN U286 ( .B(zreg[745]), .A(start), .Z(\zin[0][745] ) );
  ANDN U287 ( .B(zreg[744]), .A(start), .Z(\zin[0][744] ) );
  ANDN U288 ( .B(zreg[743]), .A(start), .Z(\zin[0][743] ) );
  ANDN U289 ( .B(zreg[742]), .A(start), .Z(\zin[0][742] ) );
  ANDN U290 ( .B(zreg[741]), .A(start), .Z(\zin[0][741] ) );
  ANDN U291 ( .B(zreg[740]), .A(start), .Z(\zin[0][740] ) );
  ANDN U292 ( .B(zreg[73]), .A(start), .Z(\zin[0][73] ) );
  ANDN U293 ( .B(zreg[739]), .A(start), .Z(\zin[0][739] ) );
  ANDN U294 ( .B(zreg[738]), .A(start), .Z(\zin[0][738] ) );
  ANDN U295 ( .B(zreg[737]), .A(start), .Z(\zin[0][737] ) );
  ANDN U296 ( .B(zreg[736]), .A(start), .Z(\zin[0][736] ) );
  ANDN U297 ( .B(zreg[735]), .A(start), .Z(\zin[0][735] ) );
  ANDN U298 ( .B(zreg[734]), .A(start), .Z(\zin[0][734] ) );
  ANDN U299 ( .B(zreg[733]), .A(start), .Z(\zin[0][733] ) );
  ANDN U300 ( .B(zreg[732]), .A(start), .Z(\zin[0][732] ) );
  ANDN U301 ( .B(zreg[731]), .A(start), .Z(\zin[0][731] ) );
  ANDN U302 ( .B(zreg[730]), .A(start), .Z(\zin[0][730] ) );
  ANDN U303 ( .B(zreg[72]), .A(start), .Z(\zin[0][72] ) );
  ANDN U304 ( .B(zreg[729]), .A(start), .Z(\zin[0][729] ) );
  ANDN U305 ( .B(zreg[728]), .A(start), .Z(\zin[0][728] ) );
  ANDN U306 ( .B(zreg[727]), .A(start), .Z(\zin[0][727] ) );
  ANDN U307 ( .B(zreg[726]), .A(start), .Z(\zin[0][726] ) );
  ANDN U308 ( .B(zreg[725]), .A(start), .Z(\zin[0][725] ) );
  ANDN U309 ( .B(zreg[724]), .A(start), .Z(\zin[0][724] ) );
  ANDN U310 ( .B(zreg[723]), .A(start), .Z(\zin[0][723] ) );
  ANDN U311 ( .B(zreg[722]), .A(start), .Z(\zin[0][722] ) );
  ANDN U312 ( .B(zreg[721]), .A(start), .Z(\zin[0][721] ) );
  ANDN U313 ( .B(zreg[720]), .A(start), .Z(\zin[0][720] ) );
  ANDN U314 ( .B(zreg[71]), .A(start), .Z(\zin[0][71] ) );
  ANDN U315 ( .B(zreg[719]), .A(start), .Z(\zin[0][719] ) );
  ANDN U316 ( .B(zreg[718]), .A(start), .Z(\zin[0][718] ) );
  ANDN U317 ( .B(zreg[717]), .A(start), .Z(\zin[0][717] ) );
  ANDN U318 ( .B(zreg[716]), .A(start), .Z(\zin[0][716] ) );
  ANDN U319 ( .B(zreg[715]), .A(start), .Z(\zin[0][715] ) );
  ANDN U320 ( .B(zreg[714]), .A(start), .Z(\zin[0][714] ) );
  ANDN U321 ( .B(zreg[713]), .A(start), .Z(\zin[0][713] ) );
  ANDN U322 ( .B(zreg[712]), .A(start), .Z(\zin[0][712] ) );
  ANDN U323 ( .B(zreg[711]), .A(start), .Z(\zin[0][711] ) );
  ANDN U324 ( .B(zreg[710]), .A(start), .Z(\zin[0][710] ) );
  ANDN U325 ( .B(zreg[70]), .A(start), .Z(\zin[0][70] ) );
  ANDN U326 ( .B(zreg[709]), .A(start), .Z(\zin[0][709] ) );
  ANDN U327 ( .B(zreg[708]), .A(start), .Z(\zin[0][708] ) );
  ANDN U328 ( .B(zreg[707]), .A(start), .Z(\zin[0][707] ) );
  ANDN U329 ( .B(zreg[706]), .A(start), .Z(\zin[0][706] ) );
  ANDN U330 ( .B(zreg[705]), .A(start), .Z(\zin[0][705] ) );
  ANDN U331 ( .B(zreg[704]), .A(start), .Z(\zin[0][704] ) );
  ANDN U332 ( .B(zreg[703]), .A(start), .Z(\zin[0][703] ) );
  ANDN U333 ( .B(zreg[702]), .A(start), .Z(\zin[0][702] ) );
  ANDN U334 ( .B(zreg[701]), .A(start), .Z(\zin[0][701] ) );
  ANDN U335 ( .B(zreg[700]), .A(start), .Z(\zin[0][700] ) );
  ANDN U336 ( .B(zreg[6]), .A(start), .Z(\zin[0][6] ) );
  ANDN U337 ( .B(zreg[69]), .A(start), .Z(\zin[0][69] ) );
  ANDN U338 ( .B(zreg[699]), .A(start), .Z(\zin[0][699] ) );
  ANDN U339 ( .B(zreg[698]), .A(start), .Z(\zin[0][698] ) );
  ANDN U340 ( .B(zreg[697]), .A(start), .Z(\zin[0][697] ) );
  ANDN U341 ( .B(zreg[696]), .A(start), .Z(\zin[0][696] ) );
  ANDN U342 ( .B(zreg[695]), .A(start), .Z(\zin[0][695] ) );
  ANDN U343 ( .B(zreg[694]), .A(start), .Z(\zin[0][694] ) );
  ANDN U344 ( .B(zreg[693]), .A(start), .Z(\zin[0][693] ) );
  ANDN U345 ( .B(zreg[692]), .A(start), .Z(\zin[0][692] ) );
  ANDN U346 ( .B(zreg[691]), .A(start), .Z(\zin[0][691] ) );
  ANDN U347 ( .B(zreg[690]), .A(start), .Z(\zin[0][690] ) );
  ANDN U348 ( .B(zreg[68]), .A(start), .Z(\zin[0][68] ) );
  ANDN U349 ( .B(zreg[689]), .A(start), .Z(\zin[0][689] ) );
  ANDN U350 ( .B(zreg[688]), .A(start), .Z(\zin[0][688] ) );
  ANDN U351 ( .B(zreg[687]), .A(start), .Z(\zin[0][687] ) );
  ANDN U352 ( .B(zreg[686]), .A(start), .Z(\zin[0][686] ) );
  ANDN U353 ( .B(zreg[685]), .A(start), .Z(\zin[0][685] ) );
  ANDN U354 ( .B(zreg[684]), .A(start), .Z(\zin[0][684] ) );
  ANDN U355 ( .B(zreg[683]), .A(start), .Z(\zin[0][683] ) );
  ANDN U356 ( .B(zreg[682]), .A(start), .Z(\zin[0][682] ) );
  ANDN U357 ( .B(zreg[681]), .A(start), .Z(\zin[0][681] ) );
  ANDN U358 ( .B(zreg[680]), .A(start), .Z(\zin[0][680] ) );
  ANDN U359 ( .B(zreg[67]), .A(start), .Z(\zin[0][67] ) );
  ANDN U360 ( .B(zreg[679]), .A(start), .Z(\zin[0][679] ) );
  ANDN U361 ( .B(zreg[678]), .A(start), .Z(\zin[0][678] ) );
  ANDN U362 ( .B(zreg[677]), .A(start), .Z(\zin[0][677] ) );
  ANDN U363 ( .B(zreg[676]), .A(start), .Z(\zin[0][676] ) );
  ANDN U364 ( .B(zreg[675]), .A(start), .Z(\zin[0][675] ) );
  ANDN U365 ( .B(zreg[674]), .A(start), .Z(\zin[0][674] ) );
  ANDN U366 ( .B(zreg[673]), .A(start), .Z(\zin[0][673] ) );
  ANDN U367 ( .B(zreg[672]), .A(start), .Z(\zin[0][672] ) );
  ANDN U368 ( .B(zreg[671]), .A(start), .Z(\zin[0][671] ) );
  ANDN U369 ( .B(zreg[670]), .A(start), .Z(\zin[0][670] ) );
  ANDN U370 ( .B(zreg[66]), .A(start), .Z(\zin[0][66] ) );
  ANDN U371 ( .B(zreg[669]), .A(start), .Z(\zin[0][669] ) );
  ANDN U372 ( .B(zreg[668]), .A(start), .Z(\zin[0][668] ) );
  ANDN U373 ( .B(zreg[667]), .A(start), .Z(\zin[0][667] ) );
  ANDN U374 ( .B(zreg[666]), .A(start), .Z(\zin[0][666] ) );
  ANDN U375 ( .B(zreg[665]), .A(start), .Z(\zin[0][665] ) );
  ANDN U376 ( .B(zreg[664]), .A(start), .Z(\zin[0][664] ) );
  ANDN U377 ( .B(zreg[663]), .A(start), .Z(\zin[0][663] ) );
  ANDN U378 ( .B(zreg[662]), .A(start), .Z(\zin[0][662] ) );
  ANDN U379 ( .B(zreg[661]), .A(start), .Z(\zin[0][661] ) );
  ANDN U380 ( .B(zreg[660]), .A(start), .Z(\zin[0][660] ) );
  ANDN U381 ( .B(zreg[65]), .A(start), .Z(\zin[0][65] ) );
  ANDN U382 ( .B(zreg[659]), .A(start), .Z(\zin[0][659] ) );
  ANDN U383 ( .B(zreg[658]), .A(start), .Z(\zin[0][658] ) );
  ANDN U384 ( .B(zreg[657]), .A(start), .Z(\zin[0][657] ) );
  ANDN U385 ( .B(zreg[656]), .A(start), .Z(\zin[0][656] ) );
  ANDN U386 ( .B(zreg[655]), .A(start), .Z(\zin[0][655] ) );
  ANDN U387 ( .B(zreg[654]), .A(start), .Z(\zin[0][654] ) );
  ANDN U388 ( .B(zreg[653]), .A(start), .Z(\zin[0][653] ) );
  ANDN U389 ( .B(zreg[652]), .A(start), .Z(\zin[0][652] ) );
  ANDN U390 ( .B(zreg[651]), .A(start), .Z(\zin[0][651] ) );
  ANDN U391 ( .B(zreg[650]), .A(start), .Z(\zin[0][650] ) );
  ANDN U392 ( .B(zreg[64]), .A(start), .Z(\zin[0][64] ) );
  ANDN U393 ( .B(zreg[649]), .A(start), .Z(\zin[0][649] ) );
  ANDN U394 ( .B(zreg[648]), .A(start), .Z(\zin[0][648] ) );
  ANDN U395 ( .B(zreg[647]), .A(start), .Z(\zin[0][647] ) );
  ANDN U396 ( .B(zreg[646]), .A(start), .Z(\zin[0][646] ) );
  ANDN U397 ( .B(zreg[645]), .A(start), .Z(\zin[0][645] ) );
  ANDN U398 ( .B(zreg[644]), .A(start), .Z(\zin[0][644] ) );
  ANDN U399 ( .B(zreg[643]), .A(start), .Z(\zin[0][643] ) );
  ANDN U400 ( .B(zreg[642]), .A(start), .Z(\zin[0][642] ) );
  ANDN U401 ( .B(zreg[641]), .A(start), .Z(\zin[0][641] ) );
  ANDN U402 ( .B(zreg[640]), .A(start), .Z(\zin[0][640] ) );
  ANDN U403 ( .B(zreg[63]), .A(start), .Z(\zin[0][63] ) );
  ANDN U404 ( .B(zreg[639]), .A(start), .Z(\zin[0][639] ) );
  ANDN U405 ( .B(zreg[638]), .A(start), .Z(\zin[0][638] ) );
  ANDN U406 ( .B(zreg[637]), .A(start), .Z(\zin[0][637] ) );
  ANDN U407 ( .B(zreg[636]), .A(start), .Z(\zin[0][636] ) );
  ANDN U408 ( .B(zreg[635]), .A(start), .Z(\zin[0][635] ) );
  ANDN U409 ( .B(zreg[634]), .A(start), .Z(\zin[0][634] ) );
  ANDN U410 ( .B(zreg[633]), .A(start), .Z(\zin[0][633] ) );
  ANDN U411 ( .B(zreg[632]), .A(start), .Z(\zin[0][632] ) );
  ANDN U412 ( .B(zreg[631]), .A(start), .Z(\zin[0][631] ) );
  ANDN U413 ( .B(zreg[630]), .A(start), .Z(\zin[0][630] ) );
  ANDN U414 ( .B(zreg[62]), .A(start), .Z(\zin[0][62] ) );
  ANDN U415 ( .B(zreg[629]), .A(start), .Z(\zin[0][629] ) );
  ANDN U416 ( .B(zreg[628]), .A(start), .Z(\zin[0][628] ) );
  ANDN U417 ( .B(zreg[627]), .A(start), .Z(\zin[0][627] ) );
  ANDN U418 ( .B(zreg[626]), .A(start), .Z(\zin[0][626] ) );
  ANDN U419 ( .B(zreg[625]), .A(start), .Z(\zin[0][625] ) );
  ANDN U420 ( .B(zreg[624]), .A(start), .Z(\zin[0][624] ) );
  ANDN U421 ( .B(zreg[623]), .A(start), .Z(\zin[0][623] ) );
  ANDN U422 ( .B(zreg[622]), .A(start), .Z(\zin[0][622] ) );
  ANDN U423 ( .B(zreg[621]), .A(start), .Z(\zin[0][621] ) );
  ANDN U424 ( .B(zreg[620]), .A(start), .Z(\zin[0][620] ) );
  ANDN U425 ( .B(zreg[61]), .A(start), .Z(\zin[0][61] ) );
  ANDN U426 ( .B(zreg[619]), .A(start), .Z(\zin[0][619] ) );
  ANDN U427 ( .B(zreg[618]), .A(start), .Z(\zin[0][618] ) );
  ANDN U428 ( .B(zreg[617]), .A(start), .Z(\zin[0][617] ) );
  ANDN U429 ( .B(zreg[616]), .A(start), .Z(\zin[0][616] ) );
  ANDN U430 ( .B(zreg[615]), .A(start), .Z(\zin[0][615] ) );
  ANDN U431 ( .B(zreg[614]), .A(start), .Z(\zin[0][614] ) );
  ANDN U432 ( .B(zreg[613]), .A(start), .Z(\zin[0][613] ) );
  ANDN U433 ( .B(zreg[612]), .A(start), .Z(\zin[0][612] ) );
  ANDN U434 ( .B(zreg[611]), .A(start), .Z(\zin[0][611] ) );
  ANDN U435 ( .B(zreg[610]), .A(start), .Z(\zin[0][610] ) );
  ANDN U436 ( .B(zreg[60]), .A(start), .Z(\zin[0][60] ) );
  ANDN U437 ( .B(zreg[609]), .A(start), .Z(\zin[0][609] ) );
  ANDN U438 ( .B(zreg[608]), .A(start), .Z(\zin[0][608] ) );
  ANDN U439 ( .B(zreg[607]), .A(start), .Z(\zin[0][607] ) );
  ANDN U440 ( .B(zreg[606]), .A(start), .Z(\zin[0][606] ) );
  ANDN U441 ( .B(zreg[605]), .A(start), .Z(\zin[0][605] ) );
  ANDN U442 ( .B(zreg[604]), .A(start), .Z(\zin[0][604] ) );
  ANDN U443 ( .B(zreg[603]), .A(start), .Z(\zin[0][603] ) );
  ANDN U444 ( .B(zreg[602]), .A(start), .Z(\zin[0][602] ) );
  ANDN U445 ( .B(zreg[601]), .A(start), .Z(\zin[0][601] ) );
  ANDN U446 ( .B(zreg[600]), .A(start), .Z(\zin[0][600] ) );
  ANDN U447 ( .B(zreg[5]), .A(start), .Z(\zin[0][5] ) );
  ANDN U448 ( .B(zreg[59]), .A(start), .Z(\zin[0][59] ) );
  ANDN U449 ( .B(zreg[599]), .A(start), .Z(\zin[0][599] ) );
  ANDN U450 ( .B(zreg[598]), .A(start), .Z(\zin[0][598] ) );
  ANDN U451 ( .B(zreg[597]), .A(start), .Z(\zin[0][597] ) );
  ANDN U452 ( .B(zreg[596]), .A(start), .Z(\zin[0][596] ) );
  ANDN U453 ( .B(zreg[595]), .A(start), .Z(\zin[0][595] ) );
  ANDN U454 ( .B(zreg[594]), .A(start), .Z(\zin[0][594] ) );
  ANDN U455 ( .B(zreg[593]), .A(start), .Z(\zin[0][593] ) );
  ANDN U456 ( .B(zreg[592]), .A(start), .Z(\zin[0][592] ) );
  ANDN U457 ( .B(zreg[591]), .A(start), .Z(\zin[0][591] ) );
  ANDN U458 ( .B(zreg[590]), .A(start), .Z(\zin[0][590] ) );
  ANDN U459 ( .B(zreg[58]), .A(start), .Z(\zin[0][58] ) );
  ANDN U460 ( .B(zreg[589]), .A(start), .Z(\zin[0][589] ) );
  ANDN U461 ( .B(zreg[588]), .A(start), .Z(\zin[0][588] ) );
  ANDN U462 ( .B(zreg[587]), .A(start), .Z(\zin[0][587] ) );
  ANDN U463 ( .B(zreg[586]), .A(start), .Z(\zin[0][586] ) );
  ANDN U464 ( .B(zreg[585]), .A(start), .Z(\zin[0][585] ) );
  ANDN U465 ( .B(zreg[584]), .A(start), .Z(\zin[0][584] ) );
  ANDN U466 ( .B(zreg[583]), .A(start), .Z(\zin[0][583] ) );
  ANDN U467 ( .B(zreg[582]), .A(start), .Z(\zin[0][582] ) );
  ANDN U468 ( .B(zreg[581]), .A(start), .Z(\zin[0][581] ) );
  ANDN U469 ( .B(zreg[580]), .A(start), .Z(\zin[0][580] ) );
  ANDN U470 ( .B(zreg[57]), .A(start), .Z(\zin[0][57] ) );
  ANDN U471 ( .B(zreg[579]), .A(start), .Z(\zin[0][579] ) );
  ANDN U472 ( .B(zreg[578]), .A(start), .Z(\zin[0][578] ) );
  ANDN U473 ( .B(zreg[577]), .A(start), .Z(\zin[0][577] ) );
  ANDN U474 ( .B(zreg[576]), .A(start), .Z(\zin[0][576] ) );
  ANDN U475 ( .B(zreg[575]), .A(start), .Z(\zin[0][575] ) );
  ANDN U476 ( .B(zreg[574]), .A(start), .Z(\zin[0][574] ) );
  ANDN U477 ( .B(zreg[573]), .A(start), .Z(\zin[0][573] ) );
  ANDN U478 ( .B(zreg[572]), .A(start), .Z(\zin[0][572] ) );
  ANDN U479 ( .B(zreg[571]), .A(start), .Z(\zin[0][571] ) );
  ANDN U480 ( .B(zreg[570]), .A(start), .Z(\zin[0][570] ) );
  ANDN U481 ( .B(zreg[56]), .A(start), .Z(\zin[0][56] ) );
  ANDN U482 ( .B(zreg[569]), .A(start), .Z(\zin[0][569] ) );
  ANDN U483 ( .B(zreg[568]), .A(start), .Z(\zin[0][568] ) );
  ANDN U484 ( .B(zreg[567]), .A(start), .Z(\zin[0][567] ) );
  ANDN U485 ( .B(zreg[566]), .A(start), .Z(\zin[0][566] ) );
  ANDN U486 ( .B(zreg[565]), .A(start), .Z(\zin[0][565] ) );
  ANDN U487 ( .B(zreg[564]), .A(start), .Z(\zin[0][564] ) );
  ANDN U488 ( .B(zreg[563]), .A(start), .Z(\zin[0][563] ) );
  ANDN U489 ( .B(zreg[562]), .A(start), .Z(\zin[0][562] ) );
  ANDN U490 ( .B(zreg[561]), .A(start), .Z(\zin[0][561] ) );
  ANDN U491 ( .B(zreg[560]), .A(start), .Z(\zin[0][560] ) );
  ANDN U492 ( .B(zreg[55]), .A(start), .Z(\zin[0][55] ) );
  ANDN U493 ( .B(zreg[559]), .A(start), .Z(\zin[0][559] ) );
  ANDN U494 ( .B(zreg[558]), .A(start), .Z(\zin[0][558] ) );
  ANDN U495 ( .B(zreg[557]), .A(start), .Z(\zin[0][557] ) );
  ANDN U496 ( .B(zreg[556]), .A(start), .Z(\zin[0][556] ) );
  ANDN U497 ( .B(zreg[555]), .A(start), .Z(\zin[0][555] ) );
  ANDN U498 ( .B(zreg[554]), .A(start), .Z(\zin[0][554] ) );
  ANDN U499 ( .B(zreg[553]), .A(start), .Z(\zin[0][553] ) );
  ANDN U500 ( .B(zreg[552]), .A(start), .Z(\zin[0][552] ) );
  ANDN U501 ( .B(zreg[551]), .A(start), .Z(\zin[0][551] ) );
  ANDN U502 ( .B(zreg[550]), .A(start), .Z(\zin[0][550] ) );
  ANDN U503 ( .B(zreg[54]), .A(start), .Z(\zin[0][54] ) );
  ANDN U504 ( .B(zreg[549]), .A(start), .Z(\zin[0][549] ) );
  ANDN U505 ( .B(zreg[548]), .A(start), .Z(\zin[0][548] ) );
  ANDN U506 ( .B(zreg[547]), .A(start), .Z(\zin[0][547] ) );
  ANDN U507 ( .B(zreg[546]), .A(start), .Z(\zin[0][546] ) );
  ANDN U508 ( .B(zreg[545]), .A(start), .Z(\zin[0][545] ) );
  ANDN U509 ( .B(zreg[544]), .A(start), .Z(\zin[0][544] ) );
  ANDN U510 ( .B(zreg[543]), .A(start), .Z(\zin[0][543] ) );
  ANDN U511 ( .B(zreg[542]), .A(start), .Z(\zin[0][542] ) );
  ANDN U512 ( .B(zreg[541]), .A(start), .Z(\zin[0][541] ) );
  ANDN U513 ( .B(zreg[540]), .A(start), .Z(\zin[0][540] ) );
  ANDN U514 ( .B(zreg[53]), .A(start), .Z(\zin[0][53] ) );
  ANDN U515 ( .B(zreg[539]), .A(start), .Z(\zin[0][539] ) );
  ANDN U516 ( .B(zreg[538]), .A(start), .Z(\zin[0][538] ) );
  ANDN U517 ( .B(zreg[537]), .A(start), .Z(\zin[0][537] ) );
  ANDN U518 ( .B(zreg[536]), .A(start), .Z(\zin[0][536] ) );
  ANDN U519 ( .B(zreg[535]), .A(start), .Z(\zin[0][535] ) );
  ANDN U520 ( .B(zreg[534]), .A(start), .Z(\zin[0][534] ) );
  ANDN U521 ( .B(zreg[533]), .A(start), .Z(\zin[0][533] ) );
  ANDN U522 ( .B(zreg[532]), .A(start), .Z(\zin[0][532] ) );
  ANDN U523 ( .B(zreg[531]), .A(start), .Z(\zin[0][531] ) );
  ANDN U524 ( .B(zreg[530]), .A(start), .Z(\zin[0][530] ) );
  ANDN U525 ( .B(zreg[52]), .A(start), .Z(\zin[0][52] ) );
  ANDN U526 ( .B(zreg[529]), .A(start), .Z(\zin[0][529] ) );
  ANDN U527 ( .B(zreg[528]), .A(start), .Z(\zin[0][528] ) );
  ANDN U528 ( .B(zreg[527]), .A(start), .Z(\zin[0][527] ) );
  ANDN U529 ( .B(zreg[526]), .A(start), .Z(\zin[0][526] ) );
  ANDN U530 ( .B(zreg[525]), .A(start), .Z(\zin[0][525] ) );
  ANDN U531 ( .B(zreg[524]), .A(start), .Z(\zin[0][524] ) );
  ANDN U532 ( .B(zreg[523]), .A(start), .Z(\zin[0][523] ) );
  ANDN U533 ( .B(zreg[522]), .A(start), .Z(\zin[0][522] ) );
  ANDN U534 ( .B(zreg[521]), .A(start), .Z(\zin[0][521] ) );
  ANDN U535 ( .B(zreg[520]), .A(start), .Z(\zin[0][520] ) );
  ANDN U536 ( .B(zreg[51]), .A(start), .Z(\zin[0][51] ) );
  ANDN U537 ( .B(zreg[519]), .A(start), .Z(\zin[0][519] ) );
  ANDN U538 ( .B(zreg[518]), .A(start), .Z(\zin[0][518] ) );
  ANDN U539 ( .B(zreg[517]), .A(start), .Z(\zin[0][517] ) );
  ANDN U540 ( .B(zreg[516]), .A(start), .Z(\zin[0][516] ) );
  ANDN U541 ( .B(zreg[515]), .A(start), .Z(\zin[0][515] ) );
  ANDN U542 ( .B(zreg[514]), .A(start), .Z(\zin[0][514] ) );
  ANDN U543 ( .B(zreg[513]), .A(start), .Z(\zin[0][513] ) );
  ANDN U544 ( .B(zreg[512]), .A(start), .Z(\zin[0][512] ) );
  ANDN U545 ( .B(zreg[511]), .A(start), .Z(\zin[0][511] ) );
  ANDN U546 ( .B(zreg[510]), .A(start), .Z(\zin[0][510] ) );
  ANDN U547 ( .B(zreg[50]), .A(start), .Z(\zin[0][50] ) );
  ANDN U548 ( .B(zreg[509]), .A(start), .Z(\zin[0][509] ) );
  ANDN U549 ( .B(zreg[508]), .A(start), .Z(\zin[0][508] ) );
  ANDN U550 ( .B(zreg[507]), .A(start), .Z(\zin[0][507] ) );
  ANDN U551 ( .B(zreg[506]), .A(start), .Z(\zin[0][506] ) );
  ANDN U552 ( .B(zreg[505]), .A(start), .Z(\zin[0][505] ) );
  ANDN U553 ( .B(zreg[504]), .A(start), .Z(\zin[0][504] ) );
  ANDN U554 ( .B(zreg[503]), .A(start), .Z(\zin[0][503] ) );
  ANDN U555 ( .B(zreg[502]), .A(start), .Z(\zin[0][502] ) );
  ANDN U556 ( .B(zreg[501]), .A(start), .Z(\zin[0][501] ) );
  ANDN U557 ( .B(zreg[500]), .A(start), .Z(\zin[0][500] ) );
  ANDN U558 ( .B(zreg[4]), .A(start), .Z(\zin[0][4] ) );
  ANDN U559 ( .B(zreg[49]), .A(start), .Z(\zin[0][49] ) );
  ANDN U560 ( .B(zreg[499]), .A(start), .Z(\zin[0][499] ) );
  ANDN U561 ( .B(zreg[498]), .A(start), .Z(\zin[0][498] ) );
  ANDN U562 ( .B(zreg[497]), .A(start), .Z(\zin[0][497] ) );
  ANDN U563 ( .B(zreg[496]), .A(start), .Z(\zin[0][496] ) );
  ANDN U564 ( .B(zreg[495]), .A(start), .Z(\zin[0][495] ) );
  ANDN U565 ( .B(zreg[494]), .A(start), .Z(\zin[0][494] ) );
  ANDN U566 ( .B(zreg[493]), .A(start), .Z(\zin[0][493] ) );
  ANDN U567 ( .B(zreg[492]), .A(start), .Z(\zin[0][492] ) );
  ANDN U568 ( .B(zreg[491]), .A(start), .Z(\zin[0][491] ) );
  ANDN U569 ( .B(zreg[490]), .A(start), .Z(\zin[0][490] ) );
  ANDN U570 ( .B(zreg[48]), .A(start), .Z(\zin[0][48] ) );
  ANDN U571 ( .B(zreg[489]), .A(start), .Z(\zin[0][489] ) );
  ANDN U572 ( .B(zreg[488]), .A(start), .Z(\zin[0][488] ) );
  ANDN U573 ( .B(zreg[487]), .A(start), .Z(\zin[0][487] ) );
  ANDN U574 ( .B(zreg[486]), .A(start), .Z(\zin[0][486] ) );
  ANDN U575 ( .B(zreg[485]), .A(start), .Z(\zin[0][485] ) );
  ANDN U576 ( .B(zreg[484]), .A(start), .Z(\zin[0][484] ) );
  ANDN U577 ( .B(zreg[483]), .A(start), .Z(\zin[0][483] ) );
  ANDN U578 ( .B(zreg[482]), .A(start), .Z(\zin[0][482] ) );
  ANDN U579 ( .B(zreg[481]), .A(start), .Z(\zin[0][481] ) );
  ANDN U580 ( .B(zreg[480]), .A(start), .Z(\zin[0][480] ) );
  ANDN U581 ( .B(zreg[47]), .A(start), .Z(\zin[0][47] ) );
  ANDN U582 ( .B(zreg[479]), .A(start), .Z(\zin[0][479] ) );
  ANDN U583 ( .B(zreg[478]), .A(start), .Z(\zin[0][478] ) );
  ANDN U584 ( .B(zreg[477]), .A(start), .Z(\zin[0][477] ) );
  ANDN U585 ( .B(zreg[476]), .A(start), .Z(\zin[0][476] ) );
  ANDN U586 ( .B(zreg[475]), .A(start), .Z(\zin[0][475] ) );
  ANDN U587 ( .B(zreg[474]), .A(start), .Z(\zin[0][474] ) );
  ANDN U588 ( .B(zreg[473]), .A(start), .Z(\zin[0][473] ) );
  ANDN U589 ( .B(zreg[472]), .A(start), .Z(\zin[0][472] ) );
  ANDN U590 ( .B(zreg[471]), .A(start), .Z(\zin[0][471] ) );
  ANDN U591 ( .B(zreg[470]), .A(start), .Z(\zin[0][470] ) );
  ANDN U592 ( .B(zreg[46]), .A(start), .Z(\zin[0][46] ) );
  ANDN U593 ( .B(zreg[469]), .A(start), .Z(\zin[0][469] ) );
  ANDN U594 ( .B(zreg[468]), .A(start), .Z(\zin[0][468] ) );
  ANDN U595 ( .B(zreg[467]), .A(start), .Z(\zin[0][467] ) );
  ANDN U596 ( .B(zreg[466]), .A(start), .Z(\zin[0][466] ) );
  ANDN U597 ( .B(zreg[465]), .A(start), .Z(\zin[0][465] ) );
  ANDN U598 ( .B(zreg[464]), .A(start), .Z(\zin[0][464] ) );
  ANDN U599 ( .B(zreg[463]), .A(start), .Z(\zin[0][463] ) );
  ANDN U600 ( .B(zreg[462]), .A(start), .Z(\zin[0][462] ) );
  ANDN U601 ( .B(zreg[461]), .A(start), .Z(\zin[0][461] ) );
  ANDN U602 ( .B(zreg[460]), .A(start), .Z(\zin[0][460] ) );
  ANDN U603 ( .B(zreg[45]), .A(start), .Z(\zin[0][45] ) );
  ANDN U604 ( .B(zreg[459]), .A(start), .Z(\zin[0][459] ) );
  ANDN U605 ( .B(zreg[458]), .A(start), .Z(\zin[0][458] ) );
  ANDN U606 ( .B(zreg[457]), .A(start), .Z(\zin[0][457] ) );
  ANDN U607 ( .B(zreg[456]), .A(start), .Z(\zin[0][456] ) );
  ANDN U608 ( .B(zreg[455]), .A(start), .Z(\zin[0][455] ) );
  ANDN U609 ( .B(zreg[454]), .A(start), .Z(\zin[0][454] ) );
  ANDN U610 ( .B(zreg[453]), .A(start), .Z(\zin[0][453] ) );
  ANDN U611 ( .B(zreg[452]), .A(start), .Z(\zin[0][452] ) );
  ANDN U612 ( .B(zreg[451]), .A(start), .Z(\zin[0][451] ) );
  ANDN U613 ( .B(zreg[450]), .A(start), .Z(\zin[0][450] ) );
  ANDN U614 ( .B(zreg[44]), .A(start), .Z(\zin[0][44] ) );
  ANDN U615 ( .B(zreg[449]), .A(start), .Z(\zin[0][449] ) );
  ANDN U616 ( .B(zreg[448]), .A(start), .Z(\zin[0][448] ) );
  ANDN U617 ( .B(zreg[447]), .A(start), .Z(\zin[0][447] ) );
  ANDN U618 ( .B(zreg[446]), .A(start), .Z(\zin[0][446] ) );
  ANDN U619 ( .B(zreg[445]), .A(start), .Z(\zin[0][445] ) );
  ANDN U620 ( .B(zreg[444]), .A(start), .Z(\zin[0][444] ) );
  ANDN U621 ( .B(zreg[443]), .A(start), .Z(\zin[0][443] ) );
  ANDN U622 ( .B(zreg[442]), .A(start), .Z(\zin[0][442] ) );
  ANDN U623 ( .B(zreg[441]), .A(start), .Z(\zin[0][441] ) );
  ANDN U624 ( .B(zreg[440]), .A(start), .Z(\zin[0][440] ) );
  ANDN U625 ( .B(zreg[43]), .A(start), .Z(\zin[0][43] ) );
  ANDN U626 ( .B(zreg[439]), .A(start), .Z(\zin[0][439] ) );
  ANDN U627 ( .B(zreg[438]), .A(start), .Z(\zin[0][438] ) );
  ANDN U628 ( .B(zreg[437]), .A(start), .Z(\zin[0][437] ) );
  ANDN U629 ( .B(zreg[436]), .A(start), .Z(\zin[0][436] ) );
  ANDN U630 ( .B(zreg[435]), .A(start), .Z(\zin[0][435] ) );
  ANDN U631 ( .B(zreg[434]), .A(start), .Z(\zin[0][434] ) );
  ANDN U632 ( .B(zreg[433]), .A(start), .Z(\zin[0][433] ) );
  ANDN U633 ( .B(zreg[432]), .A(start), .Z(\zin[0][432] ) );
  ANDN U634 ( .B(zreg[431]), .A(start), .Z(\zin[0][431] ) );
  ANDN U635 ( .B(zreg[430]), .A(start), .Z(\zin[0][430] ) );
  ANDN U636 ( .B(zreg[42]), .A(start), .Z(\zin[0][42] ) );
  ANDN U637 ( .B(zreg[429]), .A(start), .Z(\zin[0][429] ) );
  ANDN U638 ( .B(zreg[428]), .A(start), .Z(\zin[0][428] ) );
  ANDN U639 ( .B(zreg[427]), .A(start), .Z(\zin[0][427] ) );
  ANDN U640 ( .B(zreg[426]), .A(start), .Z(\zin[0][426] ) );
  ANDN U641 ( .B(zreg[425]), .A(start), .Z(\zin[0][425] ) );
  ANDN U642 ( .B(zreg[424]), .A(start), .Z(\zin[0][424] ) );
  ANDN U643 ( .B(zreg[423]), .A(start), .Z(\zin[0][423] ) );
  ANDN U644 ( .B(zreg[422]), .A(start), .Z(\zin[0][422] ) );
  ANDN U645 ( .B(zreg[421]), .A(start), .Z(\zin[0][421] ) );
  ANDN U646 ( .B(zreg[420]), .A(start), .Z(\zin[0][420] ) );
  ANDN U647 ( .B(zreg[41]), .A(start), .Z(\zin[0][41] ) );
  ANDN U648 ( .B(zreg[419]), .A(start), .Z(\zin[0][419] ) );
  ANDN U649 ( .B(zreg[418]), .A(start), .Z(\zin[0][418] ) );
  ANDN U650 ( .B(zreg[417]), .A(start), .Z(\zin[0][417] ) );
  ANDN U651 ( .B(zreg[416]), .A(start), .Z(\zin[0][416] ) );
  ANDN U652 ( .B(zreg[415]), .A(start), .Z(\zin[0][415] ) );
  ANDN U653 ( .B(zreg[414]), .A(start), .Z(\zin[0][414] ) );
  ANDN U654 ( .B(zreg[413]), .A(start), .Z(\zin[0][413] ) );
  ANDN U655 ( .B(zreg[412]), .A(start), .Z(\zin[0][412] ) );
  ANDN U656 ( .B(zreg[411]), .A(start), .Z(\zin[0][411] ) );
  ANDN U657 ( .B(zreg[410]), .A(start), .Z(\zin[0][410] ) );
  ANDN U658 ( .B(zreg[40]), .A(start), .Z(\zin[0][40] ) );
  ANDN U659 ( .B(zreg[409]), .A(start), .Z(\zin[0][409] ) );
  ANDN U660 ( .B(zreg[408]), .A(start), .Z(\zin[0][408] ) );
  ANDN U661 ( .B(zreg[407]), .A(start), .Z(\zin[0][407] ) );
  ANDN U662 ( .B(zreg[406]), .A(start), .Z(\zin[0][406] ) );
  ANDN U663 ( .B(zreg[405]), .A(start), .Z(\zin[0][405] ) );
  ANDN U664 ( .B(zreg[404]), .A(start), .Z(\zin[0][404] ) );
  ANDN U665 ( .B(zreg[403]), .A(start), .Z(\zin[0][403] ) );
  ANDN U666 ( .B(zreg[402]), .A(start), .Z(\zin[0][402] ) );
  ANDN U667 ( .B(zreg[401]), .A(start), .Z(\zin[0][401] ) );
  ANDN U668 ( .B(zreg[400]), .A(start), .Z(\zin[0][400] ) );
  ANDN U669 ( .B(zreg[3]), .A(start), .Z(\zin[0][3] ) );
  ANDN U670 ( .B(zreg[39]), .A(start), .Z(\zin[0][39] ) );
  ANDN U671 ( .B(zreg[399]), .A(start), .Z(\zin[0][399] ) );
  ANDN U672 ( .B(zreg[398]), .A(start), .Z(\zin[0][398] ) );
  ANDN U673 ( .B(zreg[397]), .A(start), .Z(\zin[0][397] ) );
  ANDN U674 ( .B(zreg[396]), .A(start), .Z(\zin[0][396] ) );
  ANDN U675 ( .B(zreg[395]), .A(start), .Z(\zin[0][395] ) );
  ANDN U676 ( .B(zreg[394]), .A(start), .Z(\zin[0][394] ) );
  ANDN U677 ( .B(zreg[393]), .A(start), .Z(\zin[0][393] ) );
  ANDN U678 ( .B(zreg[392]), .A(start), .Z(\zin[0][392] ) );
  ANDN U679 ( .B(zreg[391]), .A(start), .Z(\zin[0][391] ) );
  ANDN U680 ( .B(zreg[390]), .A(start), .Z(\zin[0][390] ) );
  ANDN U681 ( .B(zreg[38]), .A(start), .Z(\zin[0][38] ) );
  ANDN U682 ( .B(zreg[389]), .A(start), .Z(\zin[0][389] ) );
  ANDN U683 ( .B(zreg[388]), .A(start), .Z(\zin[0][388] ) );
  ANDN U684 ( .B(zreg[387]), .A(start), .Z(\zin[0][387] ) );
  ANDN U685 ( .B(zreg[386]), .A(start), .Z(\zin[0][386] ) );
  ANDN U686 ( .B(zreg[385]), .A(start), .Z(\zin[0][385] ) );
  ANDN U687 ( .B(zreg[384]), .A(start), .Z(\zin[0][384] ) );
  ANDN U688 ( .B(zreg[383]), .A(start), .Z(\zin[0][383] ) );
  ANDN U689 ( .B(zreg[382]), .A(start), .Z(\zin[0][382] ) );
  ANDN U690 ( .B(zreg[381]), .A(start), .Z(\zin[0][381] ) );
  ANDN U691 ( .B(zreg[380]), .A(start), .Z(\zin[0][380] ) );
  ANDN U692 ( .B(zreg[37]), .A(start), .Z(\zin[0][37] ) );
  ANDN U693 ( .B(zreg[379]), .A(start), .Z(\zin[0][379] ) );
  ANDN U694 ( .B(zreg[378]), .A(start), .Z(\zin[0][378] ) );
  ANDN U695 ( .B(zreg[377]), .A(start), .Z(\zin[0][377] ) );
  ANDN U696 ( .B(zreg[376]), .A(start), .Z(\zin[0][376] ) );
  ANDN U697 ( .B(zreg[375]), .A(start), .Z(\zin[0][375] ) );
  ANDN U698 ( .B(zreg[374]), .A(start), .Z(\zin[0][374] ) );
  ANDN U699 ( .B(zreg[373]), .A(start), .Z(\zin[0][373] ) );
  ANDN U700 ( .B(zreg[372]), .A(start), .Z(\zin[0][372] ) );
  ANDN U701 ( .B(zreg[371]), .A(start), .Z(\zin[0][371] ) );
  ANDN U702 ( .B(zreg[370]), .A(start), .Z(\zin[0][370] ) );
  ANDN U703 ( .B(zreg[36]), .A(start), .Z(\zin[0][36] ) );
  ANDN U704 ( .B(zreg[369]), .A(start), .Z(\zin[0][369] ) );
  ANDN U705 ( .B(zreg[368]), .A(start), .Z(\zin[0][368] ) );
  ANDN U706 ( .B(zreg[367]), .A(start), .Z(\zin[0][367] ) );
  ANDN U707 ( .B(zreg[366]), .A(start), .Z(\zin[0][366] ) );
  ANDN U708 ( .B(zreg[365]), .A(start), .Z(\zin[0][365] ) );
  ANDN U709 ( .B(zreg[364]), .A(start), .Z(\zin[0][364] ) );
  ANDN U710 ( .B(zreg[363]), .A(start), .Z(\zin[0][363] ) );
  ANDN U711 ( .B(zreg[362]), .A(start), .Z(\zin[0][362] ) );
  ANDN U712 ( .B(zreg[361]), .A(start), .Z(\zin[0][361] ) );
  ANDN U713 ( .B(zreg[360]), .A(start), .Z(\zin[0][360] ) );
  ANDN U714 ( .B(zreg[35]), .A(start), .Z(\zin[0][35] ) );
  ANDN U715 ( .B(zreg[359]), .A(start), .Z(\zin[0][359] ) );
  ANDN U716 ( .B(zreg[358]), .A(start), .Z(\zin[0][358] ) );
  ANDN U717 ( .B(zreg[357]), .A(start), .Z(\zin[0][357] ) );
  ANDN U718 ( .B(zreg[356]), .A(start), .Z(\zin[0][356] ) );
  ANDN U719 ( .B(zreg[355]), .A(start), .Z(\zin[0][355] ) );
  ANDN U720 ( .B(zreg[354]), .A(start), .Z(\zin[0][354] ) );
  ANDN U721 ( .B(zreg[353]), .A(start), .Z(\zin[0][353] ) );
  ANDN U722 ( .B(zreg[352]), .A(start), .Z(\zin[0][352] ) );
  ANDN U723 ( .B(zreg[351]), .A(start), .Z(\zin[0][351] ) );
  ANDN U724 ( .B(zreg[350]), .A(start), .Z(\zin[0][350] ) );
  ANDN U725 ( .B(zreg[34]), .A(start), .Z(\zin[0][34] ) );
  ANDN U726 ( .B(zreg[349]), .A(start), .Z(\zin[0][349] ) );
  ANDN U727 ( .B(zreg[348]), .A(start), .Z(\zin[0][348] ) );
  ANDN U728 ( .B(zreg[347]), .A(start), .Z(\zin[0][347] ) );
  ANDN U729 ( .B(zreg[346]), .A(start), .Z(\zin[0][346] ) );
  ANDN U730 ( .B(zreg[345]), .A(start), .Z(\zin[0][345] ) );
  ANDN U731 ( .B(zreg[344]), .A(start), .Z(\zin[0][344] ) );
  ANDN U732 ( .B(zreg[343]), .A(start), .Z(\zin[0][343] ) );
  ANDN U733 ( .B(zreg[342]), .A(start), .Z(\zin[0][342] ) );
  ANDN U734 ( .B(zreg[341]), .A(start), .Z(\zin[0][341] ) );
  ANDN U735 ( .B(zreg[340]), .A(start), .Z(\zin[0][340] ) );
  ANDN U736 ( .B(zreg[33]), .A(start), .Z(\zin[0][33] ) );
  ANDN U737 ( .B(zreg[339]), .A(start), .Z(\zin[0][339] ) );
  ANDN U738 ( .B(zreg[338]), .A(start), .Z(\zin[0][338] ) );
  ANDN U739 ( .B(zreg[337]), .A(start), .Z(\zin[0][337] ) );
  ANDN U740 ( .B(zreg[336]), .A(start), .Z(\zin[0][336] ) );
  ANDN U741 ( .B(zreg[335]), .A(start), .Z(\zin[0][335] ) );
  ANDN U742 ( .B(zreg[334]), .A(start), .Z(\zin[0][334] ) );
  ANDN U743 ( .B(zreg[333]), .A(start), .Z(\zin[0][333] ) );
  ANDN U744 ( .B(zreg[332]), .A(start), .Z(\zin[0][332] ) );
  ANDN U745 ( .B(zreg[331]), .A(start), .Z(\zin[0][331] ) );
  ANDN U746 ( .B(zreg[330]), .A(start), .Z(\zin[0][330] ) );
  ANDN U747 ( .B(zreg[32]), .A(start), .Z(\zin[0][32] ) );
  ANDN U748 ( .B(zreg[329]), .A(start), .Z(\zin[0][329] ) );
  ANDN U749 ( .B(zreg[328]), .A(start), .Z(\zin[0][328] ) );
  ANDN U750 ( .B(zreg[327]), .A(start), .Z(\zin[0][327] ) );
  ANDN U751 ( .B(zreg[326]), .A(start), .Z(\zin[0][326] ) );
  ANDN U752 ( .B(zreg[325]), .A(start), .Z(\zin[0][325] ) );
  ANDN U753 ( .B(zreg[324]), .A(start), .Z(\zin[0][324] ) );
  ANDN U754 ( .B(zreg[323]), .A(start), .Z(\zin[0][323] ) );
  ANDN U755 ( .B(zreg[322]), .A(start), .Z(\zin[0][322] ) );
  ANDN U756 ( .B(zreg[321]), .A(start), .Z(\zin[0][321] ) );
  ANDN U757 ( .B(zreg[320]), .A(start), .Z(\zin[0][320] ) );
  ANDN U758 ( .B(zreg[31]), .A(start), .Z(\zin[0][31] ) );
  ANDN U759 ( .B(zreg[319]), .A(start), .Z(\zin[0][319] ) );
  ANDN U760 ( .B(zreg[318]), .A(start), .Z(\zin[0][318] ) );
  ANDN U761 ( .B(zreg[317]), .A(start), .Z(\zin[0][317] ) );
  ANDN U762 ( .B(zreg[316]), .A(start), .Z(\zin[0][316] ) );
  ANDN U763 ( .B(zreg[315]), .A(start), .Z(\zin[0][315] ) );
  ANDN U764 ( .B(zreg[314]), .A(start), .Z(\zin[0][314] ) );
  ANDN U765 ( .B(zreg[313]), .A(start), .Z(\zin[0][313] ) );
  ANDN U766 ( .B(zreg[312]), .A(start), .Z(\zin[0][312] ) );
  ANDN U767 ( .B(zreg[311]), .A(start), .Z(\zin[0][311] ) );
  ANDN U768 ( .B(zreg[310]), .A(start), .Z(\zin[0][310] ) );
  ANDN U769 ( .B(zreg[30]), .A(start), .Z(\zin[0][30] ) );
  ANDN U770 ( .B(zreg[309]), .A(start), .Z(\zin[0][309] ) );
  ANDN U771 ( .B(zreg[308]), .A(start), .Z(\zin[0][308] ) );
  ANDN U772 ( .B(zreg[307]), .A(start), .Z(\zin[0][307] ) );
  ANDN U773 ( .B(zreg[306]), .A(start), .Z(\zin[0][306] ) );
  ANDN U774 ( .B(zreg[305]), .A(start), .Z(\zin[0][305] ) );
  ANDN U775 ( .B(zreg[304]), .A(start), .Z(\zin[0][304] ) );
  ANDN U776 ( .B(zreg[303]), .A(start), .Z(\zin[0][303] ) );
  ANDN U777 ( .B(zreg[302]), .A(start), .Z(\zin[0][302] ) );
  ANDN U778 ( .B(zreg[301]), .A(start), .Z(\zin[0][301] ) );
  ANDN U779 ( .B(zreg[300]), .A(start), .Z(\zin[0][300] ) );
  ANDN U780 ( .B(zreg[2]), .A(start), .Z(\zin[0][2] ) );
  ANDN U781 ( .B(zreg[29]), .A(start), .Z(\zin[0][29] ) );
  ANDN U782 ( .B(zreg[299]), .A(start), .Z(\zin[0][299] ) );
  ANDN U783 ( .B(zreg[298]), .A(start), .Z(\zin[0][298] ) );
  ANDN U784 ( .B(zreg[297]), .A(start), .Z(\zin[0][297] ) );
  ANDN U785 ( .B(zreg[296]), .A(start), .Z(\zin[0][296] ) );
  ANDN U786 ( .B(zreg[295]), .A(start), .Z(\zin[0][295] ) );
  ANDN U787 ( .B(zreg[294]), .A(start), .Z(\zin[0][294] ) );
  ANDN U788 ( .B(zreg[293]), .A(start), .Z(\zin[0][293] ) );
  ANDN U789 ( .B(zreg[292]), .A(start), .Z(\zin[0][292] ) );
  ANDN U790 ( .B(zreg[291]), .A(start), .Z(\zin[0][291] ) );
  ANDN U791 ( .B(zreg[290]), .A(start), .Z(\zin[0][290] ) );
  ANDN U792 ( .B(zreg[28]), .A(start), .Z(\zin[0][28] ) );
  ANDN U793 ( .B(zreg[289]), .A(start), .Z(\zin[0][289] ) );
  ANDN U794 ( .B(zreg[288]), .A(start), .Z(\zin[0][288] ) );
  ANDN U795 ( .B(zreg[287]), .A(start), .Z(\zin[0][287] ) );
  ANDN U796 ( .B(zreg[286]), .A(start), .Z(\zin[0][286] ) );
  ANDN U797 ( .B(zreg[285]), .A(start), .Z(\zin[0][285] ) );
  ANDN U798 ( .B(zreg[284]), .A(start), .Z(\zin[0][284] ) );
  ANDN U799 ( .B(zreg[283]), .A(start), .Z(\zin[0][283] ) );
  ANDN U800 ( .B(zreg[282]), .A(start), .Z(\zin[0][282] ) );
  ANDN U801 ( .B(zreg[281]), .A(start), .Z(\zin[0][281] ) );
  ANDN U802 ( .B(zreg[280]), .A(start), .Z(\zin[0][280] ) );
  ANDN U803 ( .B(zreg[27]), .A(start), .Z(\zin[0][27] ) );
  ANDN U804 ( .B(zreg[279]), .A(start), .Z(\zin[0][279] ) );
  ANDN U805 ( .B(zreg[278]), .A(start), .Z(\zin[0][278] ) );
  ANDN U806 ( .B(zreg[277]), .A(start), .Z(\zin[0][277] ) );
  ANDN U807 ( .B(zreg[276]), .A(start), .Z(\zin[0][276] ) );
  ANDN U808 ( .B(zreg[275]), .A(start), .Z(\zin[0][275] ) );
  ANDN U809 ( .B(zreg[274]), .A(start), .Z(\zin[0][274] ) );
  ANDN U810 ( .B(zreg[273]), .A(start), .Z(\zin[0][273] ) );
  ANDN U811 ( .B(zreg[272]), .A(start), .Z(\zin[0][272] ) );
  ANDN U812 ( .B(zreg[271]), .A(start), .Z(\zin[0][271] ) );
  ANDN U813 ( .B(zreg[270]), .A(start), .Z(\zin[0][270] ) );
  ANDN U814 ( .B(zreg[26]), .A(start), .Z(\zin[0][26] ) );
  ANDN U815 ( .B(zreg[269]), .A(start), .Z(\zin[0][269] ) );
  ANDN U816 ( .B(zreg[268]), .A(start), .Z(\zin[0][268] ) );
  ANDN U817 ( .B(zreg[267]), .A(start), .Z(\zin[0][267] ) );
  ANDN U818 ( .B(zreg[266]), .A(start), .Z(\zin[0][266] ) );
  ANDN U819 ( .B(zreg[265]), .A(start), .Z(\zin[0][265] ) );
  ANDN U820 ( .B(zreg[264]), .A(start), .Z(\zin[0][264] ) );
  ANDN U821 ( .B(zreg[263]), .A(start), .Z(\zin[0][263] ) );
  ANDN U822 ( .B(zreg[262]), .A(start), .Z(\zin[0][262] ) );
  ANDN U823 ( .B(zreg[261]), .A(start), .Z(\zin[0][261] ) );
  ANDN U824 ( .B(zreg[260]), .A(start), .Z(\zin[0][260] ) );
  ANDN U825 ( .B(zreg[25]), .A(start), .Z(\zin[0][25] ) );
  ANDN U826 ( .B(zreg[259]), .A(start), .Z(\zin[0][259] ) );
  ANDN U827 ( .B(zreg[258]), .A(start), .Z(\zin[0][258] ) );
  ANDN U828 ( .B(zreg[257]), .A(start), .Z(\zin[0][257] ) );
  ANDN U829 ( .B(zreg[256]), .A(start), .Z(\zin[0][256] ) );
  ANDN U830 ( .B(zreg[255]), .A(start), .Z(\zin[0][255] ) );
  ANDN U831 ( .B(zreg[254]), .A(start), .Z(\zin[0][254] ) );
  ANDN U832 ( .B(zreg[253]), .A(start), .Z(\zin[0][253] ) );
  ANDN U833 ( .B(zreg[252]), .A(start), .Z(\zin[0][252] ) );
  ANDN U834 ( .B(zreg[251]), .A(start), .Z(\zin[0][251] ) );
  ANDN U835 ( .B(zreg[250]), .A(start), .Z(\zin[0][250] ) );
  ANDN U836 ( .B(zreg[24]), .A(start), .Z(\zin[0][24] ) );
  ANDN U837 ( .B(zreg[249]), .A(start), .Z(\zin[0][249] ) );
  ANDN U838 ( .B(zreg[248]), .A(start), .Z(\zin[0][248] ) );
  ANDN U839 ( .B(zreg[247]), .A(start), .Z(\zin[0][247] ) );
  ANDN U840 ( .B(zreg[246]), .A(start), .Z(\zin[0][246] ) );
  ANDN U841 ( .B(zreg[245]), .A(start), .Z(\zin[0][245] ) );
  ANDN U842 ( .B(zreg[244]), .A(start), .Z(\zin[0][244] ) );
  ANDN U843 ( .B(zreg[243]), .A(start), .Z(\zin[0][243] ) );
  ANDN U844 ( .B(zreg[242]), .A(start), .Z(\zin[0][242] ) );
  ANDN U845 ( .B(zreg[241]), .A(start), .Z(\zin[0][241] ) );
  ANDN U846 ( .B(zreg[240]), .A(start), .Z(\zin[0][240] ) );
  ANDN U847 ( .B(zreg[23]), .A(start), .Z(\zin[0][23] ) );
  ANDN U848 ( .B(zreg[239]), .A(start), .Z(\zin[0][239] ) );
  ANDN U849 ( .B(zreg[238]), .A(start), .Z(\zin[0][238] ) );
  ANDN U850 ( .B(zreg[237]), .A(start), .Z(\zin[0][237] ) );
  ANDN U851 ( .B(zreg[236]), .A(start), .Z(\zin[0][236] ) );
  ANDN U852 ( .B(zreg[235]), .A(start), .Z(\zin[0][235] ) );
  ANDN U853 ( .B(zreg[234]), .A(start), .Z(\zin[0][234] ) );
  ANDN U854 ( .B(zreg[233]), .A(start), .Z(\zin[0][233] ) );
  ANDN U855 ( .B(zreg[232]), .A(start), .Z(\zin[0][232] ) );
  ANDN U856 ( .B(zreg[231]), .A(start), .Z(\zin[0][231] ) );
  ANDN U857 ( .B(zreg[230]), .A(start), .Z(\zin[0][230] ) );
  ANDN U858 ( .B(zreg[22]), .A(start), .Z(\zin[0][22] ) );
  ANDN U859 ( .B(zreg[229]), .A(start), .Z(\zin[0][229] ) );
  ANDN U860 ( .B(zreg[228]), .A(start), .Z(\zin[0][228] ) );
  ANDN U861 ( .B(zreg[227]), .A(start), .Z(\zin[0][227] ) );
  ANDN U862 ( .B(zreg[226]), .A(start), .Z(\zin[0][226] ) );
  ANDN U863 ( .B(zreg[225]), .A(start), .Z(\zin[0][225] ) );
  ANDN U864 ( .B(zreg[224]), .A(start), .Z(\zin[0][224] ) );
  ANDN U865 ( .B(zreg[223]), .A(start), .Z(\zin[0][223] ) );
  ANDN U866 ( .B(zreg[222]), .A(start), .Z(\zin[0][222] ) );
  ANDN U867 ( .B(zreg[221]), .A(start), .Z(\zin[0][221] ) );
  ANDN U868 ( .B(zreg[220]), .A(start), .Z(\zin[0][220] ) );
  ANDN U869 ( .B(zreg[21]), .A(start), .Z(\zin[0][21] ) );
  ANDN U870 ( .B(zreg[219]), .A(start), .Z(\zin[0][219] ) );
  ANDN U871 ( .B(zreg[218]), .A(start), .Z(\zin[0][218] ) );
  ANDN U872 ( .B(zreg[217]), .A(start), .Z(\zin[0][217] ) );
  ANDN U873 ( .B(zreg[216]), .A(start), .Z(\zin[0][216] ) );
  ANDN U874 ( .B(zreg[215]), .A(start), .Z(\zin[0][215] ) );
  ANDN U875 ( .B(zreg[214]), .A(start), .Z(\zin[0][214] ) );
  ANDN U876 ( .B(zreg[213]), .A(start), .Z(\zin[0][213] ) );
  ANDN U877 ( .B(zreg[212]), .A(start), .Z(\zin[0][212] ) );
  ANDN U878 ( .B(zreg[211]), .A(start), .Z(\zin[0][211] ) );
  ANDN U879 ( .B(zreg[210]), .A(start), .Z(\zin[0][210] ) );
  ANDN U880 ( .B(zreg[20]), .A(start), .Z(\zin[0][20] ) );
  ANDN U881 ( .B(zreg[209]), .A(start), .Z(\zin[0][209] ) );
  ANDN U882 ( .B(zreg[208]), .A(start), .Z(\zin[0][208] ) );
  ANDN U883 ( .B(zreg[207]), .A(start), .Z(\zin[0][207] ) );
  ANDN U884 ( .B(zreg[206]), .A(start), .Z(\zin[0][206] ) );
  ANDN U885 ( .B(zreg[205]), .A(start), .Z(\zin[0][205] ) );
  ANDN U886 ( .B(zreg[204]), .A(start), .Z(\zin[0][204] ) );
  ANDN U887 ( .B(zreg[203]), .A(start), .Z(\zin[0][203] ) );
  ANDN U888 ( .B(zreg[202]), .A(start), .Z(\zin[0][202] ) );
  ANDN U889 ( .B(zreg[201]), .A(start), .Z(\zin[0][201] ) );
  ANDN U890 ( .B(zreg[200]), .A(start), .Z(\zin[0][200] ) );
  ANDN U891 ( .B(zreg[1]), .A(start), .Z(\zin[0][1] ) );
  ANDN U892 ( .B(zreg[19]), .A(start), .Z(\zin[0][19] ) );
  ANDN U893 ( .B(zreg[199]), .A(start), .Z(\zin[0][199] ) );
  ANDN U894 ( .B(zreg[198]), .A(start), .Z(\zin[0][198] ) );
  ANDN U895 ( .B(zreg[197]), .A(start), .Z(\zin[0][197] ) );
  ANDN U896 ( .B(zreg[196]), .A(start), .Z(\zin[0][196] ) );
  ANDN U897 ( .B(zreg[195]), .A(start), .Z(\zin[0][195] ) );
  ANDN U898 ( .B(zreg[194]), .A(start), .Z(\zin[0][194] ) );
  ANDN U899 ( .B(zreg[193]), .A(start), .Z(\zin[0][193] ) );
  ANDN U900 ( .B(zreg[192]), .A(start), .Z(\zin[0][192] ) );
  ANDN U901 ( .B(zreg[191]), .A(start), .Z(\zin[0][191] ) );
  ANDN U902 ( .B(zreg[190]), .A(start), .Z(\zin[0][190] ) );
  ANDN U903 ( .B(zreg[18]), .A(start), .Z(\zin[0][18] ) );
  ANDN U904 ( .B(zreg[189]), .A(start), .Z(\zin[0][189] ) );
  ANDN U905 ( .B(zreg[188]), .A(start), .Z(\zin[0][188] ) );
  ANDN U906 ( .B(zreg[187]), .A(start), .Z(\zin[0][187] ) );
  ANDN U907 ( .B(zreg[186]), .A(start), .Z(\zin[0][186] ) );
  ANDN U908 ( .B(zreg[185]), .A(start), .Z(\zin[0][185] ) );
  ANDN U909 ( .B(zreg[184]), .A(start), .Z(\zin[0][184] ) );
  ANDN U910 ( .B(zreg[183]), .A(start), .Z(\zin[0][183] ) );
  ANDN U911 ( .B(zreg[182]), .A(start), .Z(\zin[0][182] ) );
  ANDN U912 ( .B(zreg[181]), .A(start), .Z(\zin[0][181] ) );
  ANDN U913 ( .B(zreg[180]), .A(start), .Z(\zin[0][180] ) );
  ANDN U914 ( .B(zreg[17]), .A(start), .Z(\zin[0][17] ) );
  ANDN U915 ( .B(zreg[179]), .A(start), .Z(\zin[0][179] ) );
  ANDN U916 ( .B(zreg[178]), .A(start), .Z(\zin[0][178] ) );
  ANDN U917 ( .B(zreg[177]), .A(start), .Z(\zin[0][177] ) );
  ANDN U918 ( .B(zreg[176]), .A(start), .Z(\zin[0][176] ) );
  ANDN U919 ( .B(zreg[175]), .A(start), .Z(\zin[0][175] ) );
  ANDN U920 ( .B(zreg[174]), .A(start), .Z(\zin[0][174] ) );
  ANDN U921 ( .B(zreg[173]), .A(start), .Z(\zin[0][173] ) );
  ANDN U922 ( .B(zreg[172]), .A(start), .Z(\zin[0][172] ) );
  ANDN U923 ( .B(zreg[171]), .A(start), .Z(\zin[0][171] ) );
  ANDN U924 ( .B(zreg[170]), .A(start), .Z(\zin[0][170] ) );
  ANDN U925 ( .B(zreg[16]), .A(start), .Z(\zin[0][16] ) );
  ANDN U926 ( .B(zreg[169]), .A(start), .Z(\zin[0][169] ) );
  ANDN U927 ( .B(zreg[168]), .A(start), .Z(\zin[0][168] ) );
  ANDN U928 ( .B(zreg[167]), .A(start), .Z(\zin[0][167] ) );
  ANDN U929 ( .B(zreg[166]), .A(start), .Z(\zin[0][166] ) );
  ANDN U930 ( .B(zreg[165]), .A(start), .Z(\zin[0][165] ) );
  ANDN U931 ( .B(zreg[164]), .A(start), .Z(\zin[0][164] ) );
  ANDN U932 ( .B(zreg[163]), .A(start), .Z(\zin[0][163] ) );
  ANDN U933 ( .B(zreg[162]), .A(start), .Z(\zin[0][162] ) );
  ANDN U934 ( .B(zreg[161]), .A(start), .Z(\zin[0][161] ) );
  ANDN U935 ( .B(zreg[160]), .A(start), .Z(\zin[0][160] ) );
  ANDN U936 ( .B(zreg[15]), .A(start), .Z(\zin[0][15] ) );
  ANDN U937 ( .B(zreg[159]), .A(start), .Z(\zin[0][159] ) );
  ANDN U938 ( .B(zreg[158]), .A(start), .Z(\zin[0][158] ) );
  ANDN U939 ( .B(zreg[157]), .A(start), .Z(\zin[0][157] ) );
  ANDN U940 ( .B(zreg[156]), .A(start), .Z(\zin[0][156] ) );
  ANDN U941 ( .B(zreg[155]), .A(start), .Z(\zin[0][155] ) );
  ANDN U942 ( .B(zreg[154]), .A(start), .Z(\zin[0][154] ) );
  ANDN U943 ( .B(zreg[153]), .A(start), .Z(\zin[0][153] ) );
  ANDN U944 ( .B(zreg[152]), .A(start), .Z(\zin[0][152] ) );
  ANDN U945 ( .B(zreg[151]), .A(start), .Z(\zin[0][151] ) );
  ANDN U946 ( .B(zreg[150]), .A(start), .Z(\zin[0][150] ) );
  ANDN U947 ( .B(zreg[14]), .A(start), .Z(\zin[0][14] ) );
  ANDN U948 ( .B(zreg[149]), .A(start), .Z(\zin[0][149] ) );
  ANDN U949 ( .B(zreg[148]), .A(start), .Z(\zin[0][148] ) );
  ANDN U950 ( .B(zreg[147]), .A(start), .Z(\zin[0][147] ) );
  ANDN U951 ( .B(zreg[146]), .A(start), .Z(\zin[0][146] ) );
  ANDN U952 ( .B(zreg[145]), .A(start), .Z(\zin[0][145] ) );
  ANDN U953 ( .B(zreg[144]), .A(start), .Z(\zin[0][144] ) );
  ANDN U954 ( .B(zreg[143]), .A(start), .Z(\zin[0][143] ) );
  ANDN U955 ( .B(zreg[142]), .A(start), .Z(\zin[0][142] ) );
  ANDN U956 ( .B(zreg[141]), .A(start), .Z(\zin[0][141] ) );
  ANDN U957 ( .B(zreg[140]), .A(start), .Z(\zin[0][140] ) );
  ANDN U958 ( .B(zreg[13]), .A(start), .Z(\zin[0][13] ) );
  ANDN U959 ( .B(zreg[139]), .A(start), .Z(\zin[0][139] ) );
  ANDN U960 ( .B(zreg[138]), .A(start), .Z(\zin[0][138] ) );
  ANDN U961 ( .B(zreg[137]), .A(start), .Z(\zin[0][137] ) );
  ANDN U962 ( .B(zreg[136]), .A(start), .Z(\zin[0][136] ) );
  ANDN U963 ( .B(zreg[135]), .A(start), .Z(\zin[0][135] ) );
  ANDN U964 ( .B(zreg[134]), .A(start), .Z(\zin[0][134] ) );
  ANDN U965 ( .B(zreg[133]), .A(start), .Z(\zin[0][133] ) );
  ANDN U966 ( .B(zreg[132]), .A(start), .Z(\zin[0][132] ) );
  ANDN U967 ( .B(zreg[131]), .A(start), .Z(\zin[0][131] ) );
  ANDN U968 ( .B(zreg[130]), .A(start), .Z(\zin[0][130] ) );
  ANDN U969 ( .B(zreg[12]), .A(start), .Z(\zin[0][12] ) );
  ANDN U970 ( .B(zreg[129]), .A(start), .Z(\zin[0][129] ) );
  ANDN U971 ( .B(zreg[128]), .A(start), .Z(\zin[0][128] ) );
  ANDN U972 ( .B(zreg[127]), .A(start), .Z(\zin[0][127] ) );
  ANDN U973 ( .B(zreg[126]), .A(start), .Z(\zin[0][126] ) );
  ANDN U974 ( .B(zreg[125]), .A(start), .Z(\zin[0][125] ) );
  ANDN U975 ( .B(zreg[124]), .A(start), .Z(\zin[0][124] ) );
  ANDN U976 ( .B(zreg[123]), .A(start), .Z(\zin[0][123] ) );
  ANDN U977 ( .B(zreg[122]), .A(start), .Z(\zin[0][122] ) );
  ANDN U978 ( .B(zreg[121]), .A(start), .Z(\zin[0][121] ) );
  ANDN U979 ( .B(zreg[120]), .A(start), .Z(\zin[0][120] ) );
  ANDN U980 ( .B(zreg[11]), .A(start), .Z(\zin[0][11] ) );
  ANDN U981 ( .B(zreg[119]), .A(start), .Z(\zin[0][119] ) );
  ANDN U982 ( .B(zreg[118]), .A(start), .Z(\zin[0][118] ) );
  ANDN U983 ( .B(zreg[117]), .A(start), .Z(\zin[0][117] ) );
  ANDN U984 ( .B(zreg[116]), .A(start), .Z(\zin[0][116] ) );
  ANDN U985 ( .B(zreg[115]), .A(start), .Z(\zin[0][115] ) );
  ANDN U986 ( .B(zreg[114]), .A(start), .Z(\zin[0][114] ) );
  ANDN U987 ( .B(zreg[113]), .A(start), .Z(\zin[0][113] ) );
  ANDN U988 ( .B(zreg[112]), .A(start), .Z(\zin[0][112] ) );
  ANDN U989 ( .B(zreg[111]), .A(start), .Z(\zin[0][111] ) );
  ANDN U990 ( .B(zreg[110]), .A(start), .Z(\zin[0][110] ) );
  ANDN U991 ( .B(zreg[10]), .A(start), .Z(\zin[0][10] ) );
  ANDN U992 ( .B(zreg[109]), .A(start), .Z(\zin[0][109] ) );
  ANDN U993 ( .B(zreg[108]), .A(start), .Z(\zin[0][108] ) );
  ANDN U994 ( .B(zreg[107]), .A(start), .Z(\zin[0][107] ) );
  ANDN U995 ( .B(zreg[106]), .A(start), .Z(\zin[0][106] ) );
  ANDN U996 ( .B(zreg[105]), .A(start), .Z(\zin[0][105] ) );
  ANDN U997 ( .B(zreg[104]), .A(start), .Z(\zin[0][104] ) );
  ANDN U998 ( .B(zreg[103]), .A(start), .Z(\zin[0][103] ) );
  ANDN U999 ( .B(zreg[102]), .A(start), .Z(\zin[0][102] ) );
  ANDN U1000 ( .B(zreg[1025]), .A(start), .Z(\zin[0][1025] ) );
  ANDN U1001 ( .B(zreg[1024]), .A(start), .Z(\zin[0][1024] ) );
  ANDN U1002 ( .B(zreg[1023]), .A(start), .Z(\zin[0][1023] ) );
  ANDN U1003 ( .B(zreg[1022]), .A(start), .Z(\zin[0][1022] ) );
  ANDN U1004 ( .B(zreg[1021]), .A(start), .Z(\zin[0][1021] ) );
  ANDN U1005 ( .B(zreg[1020]), .A(start), .Z(\zin[0][1020] ) );
  ANDN U1006 ( .B(zreg[101]), .A(start), .Z(\zin[0][101] ) );
  ANDN U1007 ( .B(zreg[1019]), .A(start), .Z(\zin[0][1019] ) );
  ANDN U1008 ( .B(zreg[1018]), .A(start), .Z(\zin[0][1018] ) );
  ANDN U1009 ( .B(zreg[1017]), .A(start), .Z(\zin[0][1017] ) );
  ANDN U1010 ( .B(zreg[1016]), .A(start), .Z(\zin[0][1016] ) );
  ANDN U1011 ( .B(zreg[1015]), .A(start), .Z(\zin[0][1015] ) );
  ANDN U1012 ( .B(zreg[1014]), .A(start), .Z(\zin[0][1014] ) );
  ANDN U1013 ( .B(zreg[1013]), .A(start), .Z(\zin[0][1013] ) );
  ANDN U1014 ( .B(zreg[1012]), .A(start), .Z(\zin[0][1012] ) );
  ANDN U1015 ( .B(zreg[1011]), .A(start), .Z(\zin[0][1011] ) );
  ANDN U1016 ( .B(zreg[1010]), .A(start), .Z(\zin[0][1010] ) );
  ANDN U1017 ( .B(zreg[100]), .A(start), .Z(\zin[0][100] ) );
  ANDN U1018 ( .B(zreg[1009]), .A(start), .Z(\zin[0][1009] ) );
  ANDN U1019 ( .B(zreg[1008]), .A(start), .Z(\zin[0][1008] ) );
  ANDN U1020 ( .B(zreg[1007]), .A(start), .Z(\zin[0][1007] ) );
  ANDN U1021 ( .B(zreg[1006]), .A(start), .Z(\zin[0][1006] ) );
  ANDN U1022 ( .B(zreg[1005]), .A(start), .Z(\zin[0][1005] ) );
  ANDN U1023 ( .B(zreg[1004]), .A(start), .Z(\zin[0][1004] ) );
  ANDN U1024 ( .B(zreg[1003]), .A(start), .Z(\zin[0][1003] ) );
  ANDN U1025 ( .B(zreg[1002]), .A(start), .Z(\zin[0][1002] ) );
  ANDN U1026 ( .B(zreg[1001]), .A(start), .Z(\zin[0][1001] ) );
  ANDN U1027 ( .B(zreg[1000]), .A(start), .Z(\zin[0][1000] ) );
  ANDN U1028 ( .B(zreg[0]), .A(start), .Z(\zin[0][0] ) );
  NAND U1029 ( .A(n1), .B(n2), .Z(xin[9]) );
  NANDN U1030 ( .A(start), .B(xreg[9]), .Z(n2) );
  NAND U1031 ( .A(x[9]), .B(start), .Z(n1) );
  NAND U1032 ( .A(n3), .B(n4), .Z(xin[99]) );
  NANDN U1033 ( .A(start), .B(xreg[99]), .Z(n4) );
  NAND U1034 ( .A(x[99]), .B(start), .Z(n3) );
  NAND U1035 ( .A(n5), .B(n6), .Z(xin[999]) );
  NANDN U1036 ( .A(start), .B(xreg[999]), .Z(n6) );
  NAND U1037 ( .A(x[999]), .B(start), .Z(n5) );
  NAND U1038 ( .A(n7), .B(n8), .Z(xin[998]) );
  NANDN U1039 ( .A(start), .B(xreg[998]), .Z(n8) );
  NAND U1040 ( .A(x[998]), .B(start), .Z(n7) );
  NAND U1041 ( .A(n9), .B(n10), .Z(xin[997]) );
  NANDN U1042 ( .A(start), .B(xreg[997]), .Z(n10) );
  NAND U1043 ( .A(x[997]), .B(start), .Z(n9) );
  NAND U1044 ( .A(n11), .B(n12), .Z(xin[996]) );
  NANDN U1045 ( .A(start), .B(xreg[996]), .Z(n12) );
  NAND U1046 ( .A(x[996]), .B(start), .Z(n11) );
  NAND U1047 ( .A(n13), .B(n14), .Z(xin[995]) );
  NANDN U1048 ( .A(start), .B(xreg[995]), .Z(n14) );
  NAND U1049 ( .A(x[995]), .B(start), .Z(n13) );
  NAND U1050 ( .A(n15), .B(n16), .Z(xin[994]) );
  NANDN U1051 ( .A(start), .B(xreg[994]), .Z(n16) );
  NAND U1052 ( .A(x[994]), .B(start), .Z(n15) );
  NAND U1053 ( .A(n17), .B(n18), .Z(xin[993]) );
  NANDN U1054 ( .A(start), .B(xreg[993]), .Z(n18) );
  NAND U1055 ( .A(x[993]), .B(start), .Z(n17) );
  NAND U1056 ( .A(n19), .B(n20), .Z(xin[992]) );
  NANDN U1057 ( .A(start), .B(xreg[992]), .Z(n20) );
  NAND U1058 ( .A(x[992]), .B(start), .Z(n19) );
  NAND U1059 ( .A(n21), .B(n22), .Z(xin[991]) );
  NANDN U1060 ( .A(start), .B(xreg[991]), .Z(n22) );
  NAND U1061 ( .A(x[991]), .B(start), .Z(n21) );
  NAND U1062 ( .A(n23), .B(n24), .Z(xin[990]) );
  NANDN U1063 ( .A(start), .B(xreg[990]), .Z(n24) );
  NAND U1064 ( .A(x[990]), .B(start), .Z(n23) );
  NAND U1065 ( .A(n25), .B(n26), .Z(xin[98]) );
  NANDN U1066 ( .A(start), .B(xreg[98]), .Z(n26) );
  NAND U1067 ( .A(x[98]), .B(start), .Z(n25) );
  NAND U1068 ( .A(n27), .B(n28), .Z(xin[989]) );
  NANDN U1069 ( .A(start), .B(xreg[989]), .Z(n28) );
  NAND U1070 ( .A(x[989]), .B(start), .Z(n27) );
  NAND U1071 ( .A(n29), .B(n30), .Z(xin[988]) );
  NANDN U1072 ( .A(start), .B(xreg[988]), .Z(n30) );
  NAND U1073 ( .A(x[988]), .B(start), .Z(n29) );
  NAND U1074 ( .A(n31), .B(n32), .Z(xin[987]) );
  NANDN U1075 ( .A(start), .B(xreg[987]), .Z(n32) );
  NAND U1076 ( .A(x[987]), .B(start), .Z(n31) );
  NAND U1077 ( .A(n33), .B(n34), .Z(xin[986]) );
  NANDN U1078 ( .A(start), .B(xreg[986]), .Z(n34) );
  NAND U1079 ( .A(x[986]), .B(start), .Z(n33) );
  NAND U1080 ( .A(n35), .B(n36), .Z(xin[985]) );
  NANDN U1081 ( .A(start), .B(xreg[985]), .Z(n36) );
  NAND U1082 ( .A(x[985]), .B(start), .Z(n35) );
  NAND U1083 ( .A(n37), .B(n38), .Z(xin[984]) );
  NANDN U1084 ( .A(start), .B(xreg[984]), .Z(n38) );
  NAND U1085 ( .A(x[984]), .B(start), .Z(n37) );
  NAND U1086 ( .A(n39), .B(n40), .Z(xin[983]) );
  NANDN U1087 ( .A(start), .B(xreg[983]), .Z(n40) );
  NAND U1088 ( .A(x[983]), .B(start), .Z(n39) );
  NAND U1089 ( .A(n41), .B(n42), .Z(xin[982]) );
  NANDN U1090 ( .A(start), .B(xreg[982]), .Z(n42) );
  NAND U1091 ( .A(x[982]), .B(start), .Z(n41) );
  NAND U1092 ( .A(n43), .B(n44), .Z(xin[981]) );
  NANDN U1093 ( .A(start), .B(xreg[981]), .Z(n44) );
  NAND U1094 ( .A(x[981]), .B(start), .Z(n43) );
  NAND U1095 ( .A(n45), .B(n46), .Z(xin[980]) );
  NANDN U1096 ( .A(start), .B(xreg[980]), .Z(n46) );
  NAND U1097 ( .A(x[980]), .B(start), .Z(n45) );
  NAND U1098 ( .A(n47), .B(n48), .Z(xin[97]) );
  NANDN U1099 ( .A(start), .B(xreg[97]), .Z(n48) );
  NAND U1100 ( .A(x[97]), .B(start), .Z(n47) );
  NAND U1101 ( .A(n49), .B(n50), .Z(xin[979]) );
  NANDN U1102 ( .A(start), .B(xreg[979]), .Z(n50) );
  NAND U1103 ( .A(x[979]), .B(start), .Z(n49) );
  NAND U1104 ( .A(n51), .B(n52), .Z(xin[978]) );
  NANDN U1105 ( .A(start), .B(xreg[978]), .Z(n52) );
  NAND U1106 ( .A(x[978]), .B(start), .Z(n51) );
  NAND U1107 ( .A(n53), .B(n54), .Z(xin[977]) );
  NANDN U1108 ( .A(start), .B(xreg[977]), .Z(n54) );
  NAND U1109 ( .A(x[977]), .B(start), .Z(n53) );
  NAND U1110 ( .A(n55), .B(n56), .Z(xin[976]) );
  NANDN U1111 ( .A(start), .B(xreg[976]), .Z(n56) );
  NAND U1112 ( .A(x[976]), .B(start), .Z(n55) );
  NAND U1113 ( .A(n57), .B(n58), .Z(xin[975]) );
  NANDN U1114 ( .A(start), .B(xreg[975]), .Z(n58) );
  NAND U1115 ( .A(x[975]), .B(start), .Z(n57) );
  NAND U1116 ( .A(n59), .B(n60), .Z(xin[974]) );
  NANDN U1117 ( .A(start), .B(xreg[974]), .Z(n60) );
  NAND U1118 ( .A(x[974]), .B(start), .Z(n59) );
  NAND U1119 ( .A(n61), .B(n62), .Z(xin[973]) );
  NANDN U1120 ( .A(start), .B(xreg[973]), .Z(n62) );
  NAND U1121 ( .A(x[973]), .B(start), .Z(n61) );
  NAND U1122 ( .A(n63), .B(n64), .Z(xin[972]) );
  NANDN U1123 ( .A(start), .B(xreg[972]), .Z(n64) );
  NAND U1124 ( .A(x[972]), .B(start), .Z(n63) );
  NAND U1125 ( .A(n65), .B(n66), .Z(xin[971]) );
  NANDN U1126 ( .A(start), .B(xreg[971]), .Z(n66) );
  NAND U1127 ( .A(x[971]), .B(start), .Z(n65) );
  NAND U1128 ( .A(n67), .B(n68), .Z(xin[970]) );
  NANDN U1129 ( .A(start), .B(xreg[970]), .Z(n68) );
  NAND U1130 ( .A(x[970]), .B(start), .Z(n67) );
  NAND U1131 ( .A(n69), .B(n70), .Z(xin[96]) );
  NANDN U1132 ( .A(start), .B(xreg[96]), .Z(n70) );
  NAND U1133 ( .A(x[96]), .B(start), .Z(n69) );
  NAND U1134 ( .A(n71), .B(n72), .Z(xin[969]) );
  NANDN U1135 ( .A(start), .B(xreg[969]), .Z(n72) );
  NAND U1136 ( .A(x[969]), .B(start), .Z(n71) );
  NAND U1137 ( .A(n73), .B(n74), .Z(xin[968]) );
  NANDN U1138 ( .A(start), .B(xreg[968]), .Z(n74) );
  NAND U1139 ( .A(x[968]), .B(start), .Z(n73) );
  NAND U1140 ( .A(n75), .B(n76), .Z(xin[967]) );
  NANDN U1141 ( .A(start), .B(xreg[967]), .Z(n76) );
  NAND U1142 ( .A(x[967]), .B(start), .Z(n75) );
  NAND U1143 ( .A(n77), .B(n78), .Z(xin[966]) );
  NANDN U1144 ( .A(start), .B(xreg[966]), .Z(n78) );
  NAND U1145 ( .A(x[966]), .B(start), .Z(n77) );
  NAND U1146 ( .A(n79), .B(n80), .Z(xin[965]) );
  NANDN U1147 ( .A(start), .B(xreg[965]), .Z(n80) );
  NAND U1148 ( .A(x[965]), .B(start), .Z(n79) );
  NAND U1149 ( .A(n81), .B(n82), .Z(xin[964]) );
  NANDN U1150 ( .A(start), .B(xreg[964]), .Z(n82) );
  NAND U1151 ( .A(x[964]), .B(start), .Z(n81) );
  NAND U1152 ( .A(n83), .B(n84), .Z(xin[963]) );
  NANDN U1153 ( .A(start), .B(xreg[963]), .Z(n84) );
  NAND U1154 ( .A(x[963]), .B(start), .Z(n83) );
  NAND U1155 ( .A(n85), .B(n86), .Z(xin[962]) );
  NANDN U1156 ( .A(start), .B(xreg[962]), .Z(n86) );
  NAND U1157 ( .A(x[962]), .B(start), .Z(n85) );
  NAND U1158 ( .A(n87), .B(n88), .Z(xin[961]) );
  NANDN U1159 ( .A(start), .B(xreg[961]), .Z(n88) );
  NAND U1160 ( .A(x[961]), .B(start), .Z(n87) );
  NAND U1161 ( .A(n89), .B(n90), .Z(xin[960]) );
  NANDN U1162 ( .A(start), .B(xreg[960]), .Z(n90) );
  NAND U1163 ( .A(x[960]), .B(start), .Z(n89) );
  NAND U1164 ( .A(n91), .B(n92), .Z(xin[95]) );
  NANDN U1165 ( .A(start), .B(xreg[95]), .Z(n92) );
  NAND U1166 ( .A(x[95]), .B(start), .Z(n91) );
  NAND U1167 ( .A(n93), .B(n94), .Z(xin[959]) );
  NANDN U1168 ( .A(start), .B(xreg[959]), .Z(n94) );
  NAND U1169 ( .A(x[959]), .B(start), .Z(n93) );
  NAND U1170 ( .A(n95), .B(n96), .Z(xin[958]) );
  NANDN U1171 ( .A(start), .B(xreg[958]), .Z(n96) );
  NAND U1172 ( .A(x[958]), .B(start), .Z(n95) );
  NAND U1173 ( .A(n97), .B(n98), .Z(xin[957]) );
  NANDN U1174 ( .A(start), .B(xreg[957]), .Z(n98) );
  NAND U1175 ( .A(x[957]), .B(start), .Z(n97) );
  NAND U1176 ( .A(n99), .B(n100), .Z(xin[956]) );
  NANDN U1177 ( .A(start), .B(xreg[956]), .Z(n100) );
  NAND U1178 ( .A(x[956]), .B(start), .Z(n99) );
  NAND U1179 ( .A(n101), .B(n102), .Z(xin[955]) );
  NANDN U1180 ( .A(start), .B(xreg[955]), .Z(n102) );
  NAND U1181 ( .A(x[955]), .B(start), .Z(n101) );
  NAND U1182 ( .A(n103), .B(n104), .Z(xin[954]) );
  NANDN U1183 ( .A(start), .B(xreg[954]), .Z(n104) );
  NAND U1184 ( .A(x[954]), .B(start), .Z(n103) );
  NAND U1185 ( .A(n105), .B(n106), .Z(xin[953]) );
  NANDN U1186 ( .A(start), .B(xreg[953]), .Z(n106) );
  NAND U1187 ( .A(x[953]), .B(start), .Z(n105) );
  NAND U1188 ( .A(n107), .B(n108), .Z(xin[952]) );
  NANDN U1189 ( .A(start), .B(xreg[952]), .Z(n108) );
  NAND U1190 ( .A(x[952]), .B(start), .Z(n107) );
  NAND U1191 ( .A(n109), .B(n110), .Z(xin[951]) );
  NANDN U1192 ( .A(start), .B(xreg[951]), .Z(n110) );
  NAND U1193 ( .A(x[951]), .B(start), .Z(n109) );
  NAND U1194 ( .A(n111), .B(n112), .Z(xin[950]) );
  NANDN U1195 ( .A(start), .B(xreg[950]), .Z(n112) );
  NAND U1196 ( .A(x[950]), .B(start), .Z(n111) );
  NAND U1197 ( .A(n113), .B(n114), .Z(xin[94]) );
  NANDN U1198 ( .A(start), .B(xreg[94]), .Z(n114) );
  NAND U1199 ( .A(x[94]), .B(start), .Z(n113) );
  NAND U1200 ( .A(n115), .B(n116), .Z(xin[949]) );
  NANDN U1201 ( .A(start), .B(xreg[949]), .Z(n116) );
  NAND U1202 ( .A(x[949]), .B(start), .Z(n115) );
  NAND U1203 ( .A(n117), .B(n118), .Z(xin[948]) );
  NANDN U1204 ( .A(start), .B(xreg[948]), .Z(n118) );
  NAND U1205 ( .A(x[948]), .B(start), .Z(n117) );
  NAND U1206 ( .A(n119), .B(n120), .Z(xin[947]) );
  NANDN U1207 ( .A(start), .B(xreg[947]), .Z(n120) );
  NAND U1208 ( .A(x[947]), .B(start), .Z(n119) );
  NAND U1209 ( .A(n121), .B(n122), .Z(xin[946]) );
  NANDN U1210 ( .A(start), .B(xreg[946]), .Z(n122) );
  NAND U1211 ( .A(x[946]), .B(start), .Z(n121) );
  NAND U1212 ( .A(n123), .B(n124), .Z(xin[945]) );
  NANDN U1213 ( .A(start), .B(xreg[945]), .Z(n124) );
  NAND U1214 ( .A(x[945]), .B(start), .Z(n123) );
  NAND U1215 ( .A(n125), .B(n126), .Z(xin[944]) );
  NANDN U1216 ( .A(start), .B(xreg[944]), .Z(n126) );
  NAND U1217 ( .A(x[944]), .B(start), .Z(n125) );
  NAND U1218 ( .A(n127), .B(n128), .Z(xin[943]) );
  NANDN U1219 ( .A(start), .B(xreg[943]), .Z(n128) );
  NAND U1220 ( .A(x[943]), .B(start), .Z(n127) );
  NAND U1221 ( .A(n129), .B(n130), .Z(xin[942]) );
  NANDN U1222 ( .A(start), .B(xreg[942]), .Z(n130) );
  NAND U1223 ( .A(x[942]), .B(start), .Z(n129) );
  NAND U1224 ( .A(n131), .B(n132), .Z(xin[941]) );
  NANDN U1225 ( .A(start), .B(xreg[941]), .Z(n132) );
  NAND U1226 ( .A(x[941]), .B(start), .Z(n131) );
  NAND U1227 ( .A(n133), .B(n134), .Z(xin[940]) );
  NANDN U1228 ( .A(start), .B(xreg[940]), .Z(n134) );
  NAND U1229 ( .A(x[940]), .B(start), .Z(n133) );
  NAND U1230 ( .A(n135), .B(n136), .Z(xin[93]) );
  NANDN U1231 ( .A(start), .B(xreg[93]), .Z(n136) );
  NAND U1232 ( .A(x[93]), .B(start), .Z(n135) );
  NAND U1233 ( .A(n137), .B(n138), .Z(xin[939]) );
  NANDN U1234 ( .A(start), .B(xreg[939]), .Z(n138) );
  NAND U1235 ( .A(x[939]), .B(start), .Z(n137) );
  NAND U1236 ( .A(n139), .B(n140), .Z(xin[938]) );
  NANDN U1237 ( .A(start), .B(xreg[938]), .Z(n140) );
  NAND U1238 ( .A(x[938]), .B(start), .Z(n139) );
  NAND U1239 ( .A(n141), .B(n142), .Z(xin[937]) );
  NANDN U1240 ( .A(start), .B(xreg[937]), .Z(n142) );
  NAND U1241 ( .A(x[937]), .B(start), .Z(n141) );
  NAND U1242 ( .A(n143), .B(n144), .Z(xin[936]) );
  NANDN U1243 ( .A(start), .B(xreg[936]), .Z(n144) );
  NAND U1244 ( .A(x[936]), .B(start), .Z(n143) );
  NAND U1245 ( .A(n145), .B(n146), .Z(xin[935]) );
  NANDN U1246 ( .A(start), .B(xreg[935]), .Z(n146) );
  NAND U1247 ( .A(x[935]), .B(start), .Z(n145) );
  NAND U1248 ( .A(n147), .B(n148), .Z(xin[934]) );
  NANDN U1249 ( .A(start), .B(xreg[934]), .Z(n148) );
  NAND U1250 ( .A(x[934]), .B(start), .Z(n147) );
  NAND U1251 ( .A(n149), .B(n150), .Z(xin[933]) );
  NANDN U1252 ( .A(start), .B(xreg[933]), .Z(n150) );
  NAND U1253 ( .A(x[933]), .B(start), .Z(n149) );
  NAND U1254 ( .A(n151), .B(n152), .Z(xin[932]) );
  NANDN U1255 ( .A(start), .B(xreg[932]), .Z(n152) );
  NAND U1256 ( .A(x[932]), .B(start), .Z(n151) );
  NAND U1257 ( .A(n153), .B(n154), .Z(xin[931]) );
  NANDN U1258 ( .A(start), .B(xreg[931]), .Z(n154) );
  NAND U1259 ( .A(x[931]), .B(start), .Z(n153) );
  NAND U1260 ( .A(n155), .B(n156), .Z(xin[930]) );
  NANDN U1261 ( .A(start), .B(xreg[930]), .Z(n156) );
  NAND U1262 ( .A(x[930]), .B(start), .Z(n155) );
  NAND U1263 ( .A(n157), .B(n158), .Z(xin[92]) );
  NANDN U1264 ( .A(start), .B(xreg[92]), .Z(n158) );
  NAND U1265 ( .A(x[92]), .B(start), .Z(n157) );
  NAND U1266 ( .A(n159), .B(n160), .Z(xin[929]) );
  NANDN U1267 ( .A(start), .B(xreg[929]), .Z(n160) );
  NAND U1268 ( .A(x[929]), .B(start), .Z(n159) );
  NAND U1269 ( .A(n161), .B(n162), .Z(xin[928]) );
  NANDN U1270 ( .A(start), .B(xreg[928]), .Z(n162) );
  NAND U1271 ( .A(x[928]), .B(start), .Z(n161) );
  NAND U1272 ( .A(n163), .B(n164), .Z(xin[927]) );
  NANDN U1273 ( .A(start), .B(xreg[927]), .Z(n164) );
  NAND U1274 ( .A(x[927]), .B(start), .Z(n163) );
  NAND U1275 ( .A(n165), .B(n166), .Z(xin[926]) );
  NANDN U1276 ( .A(start), .B(xreg[926]), .Z(n166) );
  NAND U1277 ( .A(x[926]), .B(start), .Z(n165) );
  NAND U1278 ( .A(n167), .B(n168), .Z(xin[925]) );
  NANDN U1279 ( .A(start), .B(xreg[925]), .Z(n168) );
  NAND U1280 ( .A(x[925]), .B(start), .Z(n167) );
  NAND U1281 ( .A(n169), .B(n170), .Z(xin[924]) );
  NANDN U1282 ( .A(start), .B(xreg[924]), .Z(n170) );
  NAND U1283 ( .A(x[924]), .B(start), .Z(n169) );
  NAND U1284 ( .A(n171), .B(n172), .Z(xin[923]) );
  NANDN U1285 ( .A(start), .B(xreg[923]), .Z(n172) );
  NAND U1286 ( .A(x[923]), .B(start), .Z(n171) );
  NAND U1287 ( .A(n173), .B(n174), .Z(xin[922]) );
  NANDN U1288 ( .A(start), .B(xreg[922]), .Z(n174) );
  NAND U1289 ( .A(x[922]), .B(start), .Z(n173) );
  NAND U1290 ( .A(n175), .B(n176), .Z(xin[921]) );
  NANDN U1291 ( .A(start), .B(xreg[921]), .Z(n176) );
  NAND U1292 ( .A(x[921]), .B(start), .Z(n175) );
  NAND U1293 ( .A(n177), .B(n178), .Z(xin[920]) );
  NANDN U1294 ( .A(start), .B(xreg[920]), .Z(n178) );
  NAND U1295 ( .A(x[920]), .B(start), .Z(n177) );
  NAND U1296 ( .A(n179), .B(n180), .Z(xin[91]) );
  NANDN U1297 ( .A(start), .B(xreg[91]), .Z(n180) );
  NAND U1298 ( .A(x[91]), .B(start), .Z(n179) );
  NAND U1299 ( .A(n181), .B(n182), .Z(xin[919]) );
  NANDN U1300 ( .A(start), .B(xreg[919]), .Z(n182) );
  NAND U1301 ( .A(x[919]), .B(start), .Z(n181) );
  NAND U1302 ( .A(n183), .B(n184), .Z(xin[918]) );
  NANDN U1303 ( .A(start), .B(xreg[918]), .Z(n184) );
  NAND U1304 ( .A(x[918]), .B(start), .Z(n183) );
  NAND U1305 ( .A(n185), .B(n186), .Z(xin[917]) );
  NANDN U1306 ( .A(start), .B(xreg[917]), .Z(n186) );
  NAND U1307 ( .A(x[917]), .B(start), .Z(n185) );
  NAND U1308 ( .A(n187), .B(n188), .Z(xin[916]) );
  NANDN U1309 ( .A(start), .B(xreg[916]), .Z(n188) );
  NAND U1310 ( .A(x[916]), .B(start), .Z(n187) );
  NAND U1311 ( .A(n189), .B(n190), .Z(xin[915]) );
  NANDN U1312 ( .A(start), .B(xreg[915]), .Z(n190) );
  NAND U1313 ( .A(x[915]), .B(start), .Z(n189) );
  NAND U1314 ( .A(n191), .B(n192), .Z(xin[914]) );
  NANDN U1315 ( .A(start), .B(xreg[914]), .Z(n192) );
  NAND U1316 ( .A(x[914]), .B(start), .Z(n191) );
  NAND U1317 ( .A(n193), .B(n194), .Z(xin[913]) );
  NANDN U1318 ( .A(start), .B(xreg[913]), .Z(n194) );
  NAND U1319 ( .A(x[913]), .B(start), .Z(n193) );
  NAND U1320 ( .A(n195), .B(n196), .Z(xin[912]) );
  NANDN U1321 ( .A(start), .B(xreg[912]), .Z(n196) );
  NAND U1322 ( .A(x[912]), .B(start), .Z(n195) );
  NAND U1323 ( .A(n197), .B(n198), .Z(xin[911]) );
  NANDN U1324 ( .A(start), .B(xreg[911]), .Z(n198) );
  NAND U1325 ( .A(x[911]), .B(start), .Z(n197) );
  NAND U1326 ( .A(n199), .B(n200), .Z(xin[910]) );
  NANDN U1327 ( .A(start), .B(xreg[910]), .Z(n200) );
  NAND U1328 ( .A(x[910]), .B(start), .Z(n199) );
  NAND U1329 ( .A(n201), .B(n202), .Z(xin[90]) );
  NANDN U1330 ( .A(start), .B(xreg[90]), .Z(n202) );
  NAND U1331 ( .A(x[90]), .B(start), .Z(n201) );
  NAND U1332 ( .A(n203), .B(n204), .Z(xin[909]) );
  NANDN U1333 ( .A(start), .B(xreg[909]), .Z(n204) );
  NAND U1334 ( .A(x[909]), .B(start), .Z(n203) );
  NAND U1335 ( .A(n205), .B(n206), .Z(xin[908]) );
  NANDN U1336 ( .A(start), .B(xreg[908]), .Z(n206) );
  NAND U1337 ( .A(x[908]), .B(start), .Z(n205) );
  NAND U1338 ( .A(n207), .B(n208), .Z(xin[907]) );
  NANDN U1339 ( .A(start), .B(xreg[907]), .Z(n208) );
  NAND U1340 ( .A(x[907]), .B(start), .Z(n207) );
  NAND U1341 ( .A(n209), .B(n210), .Z(xin[906]) );
  NANDN U1342 ( .A(start), .B(xreg[906]), .Z(n210) );
  NAND U1343 ( .A(x[906]), .B(start), .Z(n209) );
  NAND U1344 ( .A(n211), .B(n212), .Z(xin[905]) );
  NANDN U1345 ( .A(start), .B(xreg[905]), .Z(n212) );
  NAND U1346 ( .A(x[905]), .B(start), .Z(n211) );
  NAND U1347 ( .A(n213), .B(n214), .Z(xin[904]) );
  NANDN U1348 ( .A(start), .B(xreg[904]), .Z(n214) );
  NAND U1349 ( .A(x[904]), .B(start), .Z(n213) );
  NAND U1350 ( .A(n215), .B(n216), .Z(xin[903]) );
  NANDN U1351 ( .A(start), .B(xreg[903]), .Z(n216) );
  NAND U1352 ( .A(x[903]), .B(start), .Z(n215) );
  NAND U1353 ( .A(n217), .B(n218), .Z(xin[902]) );
  NANDN U1354 ( .A(start), .B(xreg[902]), .Z(n218) );
  NAND U1355 ( .A(x[902]), .B(start), .Z(n217) );
  NAND U1356 ( .A(n219), .B(n220), .Z(xin[901]) );
  NANDN U1357 ( .A(start), .B(xreg[901]), .Z(n220) );
  NAND U1358 ( .A(x[901]), .B(start), .Z(n219) );
  NAND U1359 ( .A(n221), .B(n222), .Z(xin[900]) );
  NANDN U1360 ( .A(start), .B(xreg[900]), .Z(n222) );
  NAND U1361 ( .A(x[900]), .B(start), .Z(n221) );
  NAND U1362 ( .A(n223), .B(n224), .Z(xin[8]) );
  NANDN U1363 ( .A(start), .B(xreg[8]), .Z(n224) );
  NAND U1364 ( .A(x[8]), .B(start), .Z(n223) );
  NAND U1365 ( .A(n225), .B(n226), .Z(xin[89]) );
  NANDN U1366 ( .A(start), .B(xreg[89]), .Z(n226) );
  NAND U1367 ( .A(x[89]), .B(start), .Z(n225) );
  NAND U1368 ( .A(n227), .B(n228), .Z(xin[899]) );
  NANDN U1369 ( .A(start), .B(xreg[899]), .Z(n228) );
  NAND U1370 ( .A(x[899]), .B(start), .Z(n227) );
  NAND U1371 ( .A(n229), .B(n230), .Z(xin[898]) );
  NANDN U1372 ( .A(start), .B(xreg[898]), .Z(n230) );
  NAND U1373 ( .A(x[898]), .B(start), .Z(n229) );
  NAND U1374 ( .A(n231), .B(n232), .Z(xin[897]) );
  NANDN U1375 ( .A(start), .B(xreg[897]), .Z(n232) );
  NAND U1376 ( .A(x[897]), .B(start), .Z(n231) );
  NAND U1377 ( .A(n233), .B(n234), .Z(xin[896]) );
  NANDN U1378 ( .A(start), .B(xreg[896]), .Z(n234) );
  NAND U1379 ( .A(x[896]), .B(start), .Z(n233) );
  NAND U1380 ( .A(n235), .B(n236), .Z(xin[895]) );
  NANDN U1381 ( .A(start), .B(xreg[895]), .Z(n236) );
  NAND U1382 ( .A(x[895]), .B(start), .Z(n235) );
  NAND U1383 ( .A(n237), .B(n238), .Z(xin[894]) );
  NANDN U1384 ( .A(start), .B(xreg[894]), .Z(n238) );
  NAND U1385 ( .A(x[894]), .B(start), .Z(n237) );
  NAND U1386 ( .A(n239), .B(n240), .Z(xin[893]) );
  NANDN U1387 ( .A(start), .B(xreg[893]), .Z(n240) );
  NAND U1388 ( .A(x[893]), .B(start), .Z(n239) );
  NAND U1389 ( .A(n241), .B(n242), .Z(xin[892]) );
  NANDN U1390 ( .A(start), .B(xreg[892]), .Z(n242) );
  NAND U1391 ( .A(x[892]), .B(start), .Z(n241) );
  NAND U1392 ( .A(n243), .B(n244), .Z(xin[891]) );
  NANDN U1393 ( .A(start), .B(xreg[891]), .Z(n244) );
  NAND U1394 ( .A(x[891]), .B(start), .Z(n243) );
  NAND U1395 ( .A(n245), .B(n246), .Z(xin[890]) );
  NANDN U1396 ( .A(start), .B(xreg[890]), .Z(n246) );
  NAND U1397 ( .A(x[890]), .B(start), .Z(n245) );
  NAND U1398 ( .A(n247), .B(n248), .Z(xin[88]) );
  NANDN U1399 ( .A(start), .B(xreg[88]), .Z(n248) );
  NAND U1400 ( .A(x[88]), .B(start), .Z(n247) );
  NAND U1401 ( .A(n249), .B(n250), .Z(xin[889]) );
  NANDN U1402 ( .A(start), .B(xreg[889]), .Z(n250) );
  NAND U1403 ( .A(x[889]), .B(start), .Z(n249) );
  NAND U1404 ( .A(n251), .B(n252), .Z(xin[888]) );
  NANDN U1405 ( .A(start), .B(xreg[888]), .Z(n252) );
  NAND U1406 ( .A(x[888]), .B(start), .Z(n251) );
  NAND U1407 ( .A(n253), .B(n254), .Z(xin[887]) );
  NANDN U1408 ( .A(start), .B(xreg[887]), .Z(n254) );
  NAND U1409 ( .A(x[887]), .B(start), .Z(n253) );
  NAND U1410 ( .A(n255), .B(n256), .Z(xin[886]) );
  NANDN U1411 ( .A(start), .B(xreg[886]), .Z(n256) );
  NAND U1412 ( .A(x[886]), .B(start), .Z(n255) );
  NAND U1413 ( .A(n257), .B(n258), .Z(xin[885]) );
  NANDN U1414 ( .A(start), .B(xreg[885]), .Z(n258) );
  NAND U1415 ( .A(x[885]), .B(start), .Z(n257) );
  NAND U1416 ( .A(n259), .B(n260), .Z(xin[884]) );
  NANDN U1417 ( .A(start), .B(xreg[884]), .Z(n260) );
  NAND U1418 ( .A(x[884]), .B(start), .Z(n259) );
  NAND U1419 ( .A(n261), .B(n262), .Z(xin[883]) );
  NANDN U1420 ( .A(start), .B(xreg[883]), .Z(n262) );
  NAND U1421 ( .A(x[883]), .B(start), .Z(n261) );
  NAND U1422 ( .A(n263), .B(n264), .Z(xin[882]) );
  NANDN U1423 ( .A(start), .B(xreg[882]), .Z(n264) );
  NAND U1424 ( .A(x[882]), .B(start), .Z(n263) );
  NAND U1425 ( .A(n265), .B(n266), .Z(xin[881]) );
  NANDN U1426 ( .A(start), .B(xreg[881]), .Z(n266) );
  NAND U1427 ( .A(x[881]), .B(start), .Z(n265) );
  NAND U1428 ( .A(n267), .B(n268), .Z(xin[880]) );
  NANDN U1429 ( .A(start), .B(xreg[880]), .Z(n268) );
  NAND U1430 ( .A(x[880]), .B(start), .Z(n267) );
  NAND U1431 ( .A(n269), .B(n270), .Z(xin[87]) );
  NANDN U1432 ( .A(start), .B(xreg[87]), .Z(n270) );
  NAND U1433 ( .A(x[87]), .B(start), .Z(n269) );
  NAND U1434 ( .A(n271), .B(n272), .Z(xin[879]) );
  NANDN U1435 ( .A(start), .B(xreg[879]), .Z(n272) );
  NAND U1436 ( .A(x[879]), .B(start), .Z(n271) );
  NAND U1437 ( .A(n273), .B(n274), .Z(xin[878]) );
  NANDN U1438 ( .A(start), .B(xreg[878]), .Z(n274) );
  NAND U1439 ( .A(x[878]), .B(start), .Z(n273) );
  NAND U1440 ( .A(n275), .B(n276), .Z(xin[877]) );
  NANDN U1441 ( .A(start), .B(xreg[877]), .Z(n276) );
  NAND U1442 ( .A(x[877]), .B(start), .Z(n275) );
  NAND U1443 ( .A(n277), .B(n278), .Z(xin[876]) );
  NANDN U1444 ( .A(start), .B(xreg[876]), .Z(n278) );
  NAND U1445 ( .A(x[876]), .B(start), .Z(n277) );
  NAND U1446 ( .A(n279), .B(n280), .Z(xin[875]) );
  NANDN U1447 ( .A(start), .B(xreg[875]), .Z(n280) );
  NAND U1448 ( .A(x[875]), .B(start), .Z(n279) );
  NAND U1449 ( .A(n281), .B(n282), .Z(xin[874]) );
  NANDN U1450 ( .A(start), .B(xreg[874]), .Z(n282) );
  NAND U1451 ( .A(x[874]), .B(start), .Z(n281) );
  NAND U1452 ( .A(n283), .B(n284), .Z(xin[873]) );
  NANDN U1453 ( .A(start), .B(xreg[873]), .Z(n284) );
  NAND U1454 ( .A(x[873]), .B(start), .Z(n283) );
  NAND U1455 ( .A(n285), .B(n286), .Z(xin[872]) );
  NANDN U1456 ( .A(start), .B(xreg[872]), .Z(n286) );
  NAND U1457 ( .A(x[872]), .B(start), .Z(n285) );
  NAND U1458 ( .A(n287), .B(n288), .Z(xin[871]) );
  NANDN U1459 ( .A(start), .B(xreg[871]), .Z(n288) );
  NAND U1460 ( .A(x[871]), .B(start), .Z(n287) );
  NAND U1461 ( .A(n289), .B(n290), .Z(xin[870]) );
  NANDN U1462 ( .A(start), .B(xreg[870]), .Z(n290) );
  NAND U1463 ( .A(x[870]), .B(start), .Z(n289) );
  NAND U1464 ( .A(n291), .B(n292), .Z(xin[86]) );
  NANDN U1465 ( .A(start), .B(xreg[86]), .Z(n292) );
  NAND U1466 ( .A(x[86]), .B(start), .Z(n291) );
  NAND U1467 ( .A(n293), .B(n294), .Z(xin[869]) );
  NANDN U1468 ( .A(start), .B(xreg[869]), .Z(n294) );
  NAND U1469 ( .A(x[869]), .B(start), .Z(n293) );
  NAND U1470 ( .A(n295), .B(n296), .Z(xin[868]) );
  NANDN U1471 ( .A(start), .B(xreg[868]), .Z(n296) );
  NAND U1472 ( .A(x[868]), .B(start), .Z(n295) );
  NAND U1473 ( .A(n297), .B(n298), .Z(xin[867]) );
  NANDN U1474 ( .A(start), .B(xreg[867]), .Z(n298) );
  NAND U1475 ( .A(x[867]), .B(start), .Z(n297) );
  NAND U1476 ( .A(n299), .B(n300), .Z(xin[866]) );
  NANDN U1477 ( .A(start), .B(xreg[866]), .Z(n300) );
  NAND U1478 ( .A(x[866]), .B(start), .Z(n299) );
  NAND U1479 ( .A(n301), .B(n302), .Z(xin[865]) );
  NANDN U1480 ( .A(start), .B(xreg[865]), .Z(n302) );
  NAND U1481 ( .A(x[865]), .B(start), .Z(n301) );
  NAND U1482 ( .A(n303), .B(n304), .Z(xin[864]) );
  NANDN U1483 ( .A(start), .B(xreg[864]), .Z(n304) );
  NAND U1484 ( .A(x[864]), .B(start), .Z(n303) );
  NAND U1485 ( .A(n305), .B(n306), .Z(xin[863]) );
  NANDN U1486 ( .A(start), .B(xreg[863]), .Z(n306) );
  NAND U1487 ( .A(x[863]), .B(start), .Z(n305) );
  NAND U1488 ( .A(n307), .B(n308), .Z(xin[862]) );
  NANDN U1489 ( .A(start), .B(xreg[862]), .Z(n308) );
  NAND U1490 ( .A(x[862]), .B(start), .Z(n307) );
  NAND U1491 ( .A(n309), .B(n310), .Z(xin[861]) );
  NANDN U1492 ( .A(start), .B(xreg[861]), .Z(n310) );
  NAND U1493 ( .A(x[861]), .B(start), .Z(n309) );
  NAND U1494 ( .A(n311), .B(n312), .Z(xin[860]) );
  NANDN U1495 ( .A(start), .B(xreg[860]), .Z(n312) );
  NAND U1496 ( .A(x[860]), .B(start), .Z(n311) );
  NAND U1497 ( .A(n313), .B(n314), .Z(xin[85]) );
  NANDN U1498 ( .A(start), .B(xreg[85]), .Z(n314) );
  NAND U1499 ( .A(x[85]), .B(start), .Z(n313) );
  NAND U1500 ( .A(n315), .B(n316), .Z(xin[859]) );
  NANDN U1501 ( .A(start), .B(xreg[859]), .Z(n316) );
  NAND U1502 ( .A(x[859]), .B(start), .Z(n315) );
  NAND U1503 ( .A(n317), .B(n318), .Z(xin[858]) );
  NANDN U1504 ( .A(start), .B(xreg[858]), .Z(n318) );
  NAND U1505 ( .A(x[858]), .B(start), .Z(n317) );
  NAND U1506 ( .A(n319), .B(n320), .Z(xin[857]) );
  NANDN U1507 ( .A(start), .B(xreg[857]), .Z(n320) );
  NAND U1508 ( .A(x[857]), .B(start), .Z(n319) );
  NAND U1509 ( .A(n321), .B(n322), .Z(xin[856]) );
  NANDN U1510 ( .A(start), .B(xreg[856]), .Z(n322) );
  NAND U1511 ( .A(x[856]), .B(start), .Z(n321) );
  NAND U1512 ( .A(n323), .B(n324), .Z(xin[855]) );
  NANDN U1513 ( .A(start), .B(xreg[855]), .Z(n324) );
  NAND U1514 ( .A(x[855]), .B(start), .Z(n323) );
  NAND U1515 ( .A(n325), .B(n326), .Z(xin[854]) );
  NANDN U1516 ( .A(start), .B(xreg[854]), .Z(n326) );
  NAND U1517 ( .A(x[854]), .B(start), .Z(n325) );
  NAND U1518 ( .A(n327), .B(n328), .Z(xin[853]) );
  NANDN U1519 ( .A(start), .B(xreg[853]), .Z(n328) );
  NAND U1520 ( .A(x[853]), .B(start), .Z(n327) );
  NAND U1521 ( .A(n329), .B(n330), .Z(xin[852]) );
  NANDN U1522 ( .A(start), .B(xreg[852]), .Z(n330) );
  NAND U1523 ( .A(x[852]), .B(start), .Z(n329) );
  NAND U1524 ( .A(n331), .B(n332), .Z(xin[851]) );
  NANDN U1525 ( .A(start), .B(xreg[851]), .Z(n332) );
  NAND U1526 ( .A(x[851]), .B(start), .Z(n331) );
  NAND U1527 ( .A(n333), .B(n334), .Z(xin[850]) );
  NANDN U1528 ( .A(start), .B(xreg[850]), .Z(n334) );
  NAND U1529 ( .A(x[850]), .B(start), .Z(n333) );
  NAND U1530 ( .A(n335), .B(n336), .Z(xin[84]) );
  NANDN U1531 ( .A(start), .B(xreg[84]), .Z(n336) );
  NAND U1532 ( .A(x[84]), .B(start), .Z(n335) );
  NAND U1533 ( .A(n337), .B(n338), .Z(xin[849]) );
  NANDN U1534 ( .A(start), .B(xreg[849]), .Z(n338) );
  NAND U1535 ( .A(x[849]), .B(start), .Z(n337) );
  NAND U1536 ( .A(n339), .B(n340), .Z(xin[848]) );
  NANDN U1537 ( .A(start), .B(xreg[848]), .Z(n340) );
  NAND U1538 ( .A(x[848]), .B(start), .Z(n339) );
  NAND U1539 ( .A(n341), .B(n342), .Z(xin[847]) );
  NANDN U1540 ( .A(start), .B(xreg[847]), .Z(n342) );
  NAND U1541 ( .A(x[847]), .B(start), .Z(n341) );
  NAND U1542 ( .A(n343), .B(n344), .Z(xin[846]) );
  NANDN U1543 ( .A(start), .B(xreg[846]), .Z(n344) );
  NAND U1544 ( .A(x[846]), .B(start), .Z(n343) );
  NAND U1545 ( .A(n345), .B(n346), .Z(xin[845]) );
  NANDN U1546 ( .A(start), .B(xreg[845]), .Z(n346) );
  NAND U1547 ( .A(x[845]), .B(start), .Z(n345) );
  NAND U1548 ( .A(n347), .B(n348), .Z(xin[844]) );
  NANDN U1549 ( .A(start), .B(xreg[844]), .Z(n348) );
  NAND U1550 ( .A(x[844]), .B(start), .Z(n347) );
  NAND U1551 ( .A(n349), .B(n350), .Z(xin[843]) );
  NANDN U1552 ( .A(start), .B(xreg[843]), .Z(n350) );
  NAND U1553 ( .A(x[843]), .B(start), .Z(n349) );
  NAND U1554 ( .A(n351), .B(n352), .Z(xin[842]) );
  NANDN U1555 ( .A(start), .B(xreg[842]), .Z(n352) );
  NAND U1556 ( .A(x[842]), .B(start), .Z(n351) );
  NAND U1557 ( .A(n353), .B(n354), .Z(xin[841]) );
  NANDN U1558 ( .A(start), .B(xreg[841]), .Z(n354) );
  NAND U1559 ( .A(x[841]), .B(start), .Z(n353) );
  NAND U1560 ( .A(n355), .B(n356), .Z(xin[840]) );
  NANDN U1561 ( .A(start), .B(xreg[840]), .Z(n356) );
  NAND U1562 ( .A(x[840]), .B(start), .Z(n355) );
  NAND U1563 ( .A(n357), .B(n358), .Z(xin[83]) );
  NANDN U1564 ( .A(start), .B(xreg[83]), .Z(n358) );
  NAND U1565 ( .A(x[83]), .B(start), .Z(n357) );
  NAND U1566 ( .A(n359), .B(n360), .Z(xin[839]) );
  NANDN U1567 ( .A(start), .B(xreg[839]), .Z(n360) );
  NAND U1568 ( .A(x[839]), .B(start), .Z(n359) );
  NAND U1569 ( .A(n361), .B(n362), .Z(xin[838]) );
  NANDN U1570 ( .A(start), .B(xreg[838]), .Z(n362) );
  NAND U1571 ( .A(x[838]), .B(start), .Z(n361) );
  NAND U1572 ( .A(n363), .B(n364), .Z(xin[837]) );
  NANDN U1573 ( .A(start), .B(xreg[837]), .Z(n364) );
  NAND U1574 ( .A(x[837]), .B(start), .Z(n363) );
  NAND U1575 ( .A(n365), .B(n366), .Z(xin[836]) );
  NANDN U1576 ( .A(start), .B(xreg[836]), .Z(n366) );
  NAND U1577 ( .A(x[836]), .B(start), .Z(n365) );
  NAND U1578 ( .A(n367), .B(n368), .Z(xin[835]) );
  NANDN U1579 ( .A(start), .B(xreg[835]), .Z(n368) );
  NAND U1580 ( .A(x[835]), .B(start), .Z(n367) );
  NAND U1581 ( .A(n369), .B(n370), .Z(xin[834]) );
  NANDN U1582 ( .A(start), .B(xreg[834]), .Z(n370) );
  NAND U1583 ( .A(x[834]), .B(start), .Z(n369) );
  NAND U1584 ( .A(n371), .B(n372), .Z(xin[833]) );
  NANDN U1585 ( .A(start), .B(xreg[833]), .Z(n372) );
  NAND U1586 ( .A(x[833]), .B(start), .Z(n371) );
  NAND U1587 ( .A(n373), .B(n374), .Z(xin[832]) );
  NANDN U1588 ( .A(start), .B(xreg[832]), .Z(n374) );
  NAND U1589 ( .A(x[832]), .B(start), .Z(n373) );
  NAND U1590 ( .A(n375), .B(n376), .Z(xin[831]) );
  NANDN U1591 ( .A(start), .B(xreg[831]), .Z(n376) );
  NAND U1592 ( .A(x[831]), .B(start), .Z(n375) );
  NAND U1593 ( .A(n377), .B(n378), .Z(xin[830]) );
  NANDN U1594 ( .A(start), .B(xreg[830]), .Z(n378) );
  NAND U1595 ( .A(x[830]), .B(start), .Z(n377) );
  NAND U1596 ( .A(n379), .B(n380), .Z(xin[82]) );
  NANDN U1597 ( .A(start), .B(xreg[82]), .Z(n380) );
  NAND U1598 ( .A(x[82]), .B(start), .Z(n379) );
  NAND U1599 ( .A(n381), .B(n382), .Z(xin[829]) );
  NANDN U1600 ( .A(start), .B(xreg[829]), .Z(n382) );
  NAND U1601 ( .A(x[829]), .B(start), .Z(n381) );
  NAND U1602 ( .A(n383), .B(n384), .Z(xin[828]) );
  NANDN U1603 ( .A(start), .B(xreg[828]), .Z(n384) );
  NAND U1604 ( .A(x[828]), .B(start), .Z(n383) );
  NAND U1605 ( .A(n385), .B(n386), .Z(xin[827]) );
  NANDN U1606 ( .A(start), .B(xreg[827]), .Z(n386) );
  NAND U1607 ( .A(x[827]), .B(start), .Z(n385) );
  NAND U1608 ( .A(n387), .B(n388), .Z(xin[826]) );
  NANDN U1609 ( .A(start), .B(xreg[826]), .Z(n388) );
  NAND U1610 ( .A(x[826]), .B(start), .Z(n387) );
  NAND U1611 ( .A(n389), .B(n390), .Z(xin[825]) );
  NANDN U1612 ( .A(start), .B(xreg[825]), .Z(n390) );
  NAND U1613 ( .A(x[825]), .B(start), .Z(n389) );
  NAND U1614 ( .A(n391), .B(n392), .Z(xin[824]) );
  NANDN U1615 ( .A(start), .B(xreg[824]), .Z(n392) );
  NAND U1616 ( .A(x[824]), .B(start), .Z(n391) );
  NAND U1617 ( .A(n393), .B(n394), .Z(xin[823]) );
  NANDN U1618 ( .A(start), .B(xreg[823]), .Z(n394) );
  NAND U1619 ( .A(x[823]), .B(start), .Z(n393) );
  NAND U1620 ( .A(n395), .B(n396), .Z(xin[822]) );
  NANDN U1621 ( .A(start), .B(xreg[822]), .Z(n396) );
  NAND U1622 ( .A(x[822]), .B(start), .Z(n395) );
  NAND U1623 ( .A(n397), .B(n398), .Z(xin[821]) );
  NANDN U1624 ( .A(start), .B(xreg[821]), .Z(n398) );
  NAND U1625 ( .A(x[821]), .B(start), .Z(n397) );
  NAND U1626 ( .A(n399), .B(n400), .Z(xin[820]) );
  NANDN U1627 ( .A(start), .B(xreg[820]), .Z(n400) );
  NAND U1628 ( .A(x[820]), .B(start), .Z(n399) );
  NAND U1629 ( .A(n401), .B(n402), .Z(xin[81]) );
  NANDN U1630 ( .A(start), .B(xreg[81]), .Z(n402) );
  NAND U1631 ( .A(x[81]), .B(start), .Z(n401) );
  NAND U1632 ( .A(n403), .B(n404), .Z(xin[819]) );
  NANDN U1633 ( .A(start), .B(xreg[819]), .Z(n404) );
  NAND U1634 ( .A(x[819]), .B(start), .Z(n403) );
  NAND U1635 ( .A(n405), .B(n406), .Z(xin[818]) );
  NANDN U1636 ( .A(start), .B(xreg[818]), .Z(n406) );
  NAND U1637 ( .A(x[818]), .B(start), .Z(n405) );
  NAND U1638 ( .A(n407), .B(n408), .Z(xin[817]) );
  NANDN U1639 ( .A(start), .B(xreg[817]), .Z(n408) );
  NAND U1640 ( .A(x[817]), .B(start), .Z(n407) );
  NAND U1641 ( .A(n409), .B(n410), .Z(xin[816]) );
  NANDN U1642 ( .A(start), .B(xreg[816]), .Z(n410) );
  NAND U1643 ( .A(x[816]), .B(start), .Z(n409) );
  NAND U1644 ( .A(n411), .B(n412), .Z(xin[815]) );
  NANDN U1645 ( .A(start), .B(xreg[815]), .Z(n412) );
  NAND U1646 ( .A(x[815]), .B(start), .Z(n411) );
  NAND U1647 ( .A(n413), .B(n414), .Z(xin[814]) );
  NANDN U1648 ( .A(start), .B(xreg[814]), .Z(n414) );
  NAND U1649 ( .A(x[814]), .B(start), .Z(n413) );
  NAND U1650 ( .A(n415), .B(n416), .Z(xin[813]) );
  NANDN U1651 ( .A(start), .B(xreg[813]), .Z(n416) );
  NAND U1652 ( .A(x[813]), .B(start), .Z(n415) );
  NAND U1653 ( .A(n417), .B(n418), .Z(xin[812]) );
  NANDN U1654 ( .A(start), .B(xreg[812]), .Z(n418) );
  NAND U1655 ( .A(x[812]), .B(start), .Z(n417) );
  NAND U1656 ( .A(n419), .B(n420), .Z(xin[811]) );
  NANDN U1657 ( .A(start), .B(xreg[811]), .Z(n420) );
  NAND U1658 ( .A(x[811]), .B(start), .Z(n419) );
  NAND U1659 ( .A(n421), .B(n422), .Z(xin[810]) );
  NANDN U1660 ( .A(start), .B(xreg[810]), .Z(n422) );
  NAND U1661 ( .A(x[810]), .B(start), .Z(n421) );
  NAND U1662 ( .A(n423), .B(n424), .Z(xin[80]) );
  NANDN U1663 ( .A(start), .B(xreg[80]), .Z(n424) );
  NAND U1664 ( .A(x[80]), .B(start), .Z(n423) );
  NAND U1665 ( .A(n425), .B(n426), .Z(xin[809]) );
  NANDN U1666 ( .A(start), .B(xreg[809]), .Z(n426) );
  NAND U1667 ( .A(x[809]), .B(start), .Z(n425) );
  NAND U1668 ( .A(n427), .B(n428), .Z(xin[808]) );
  NANDN U1669 ( .A(start), .B(xreg[808]), .Z(n428) );
  NAND U1670 ( .A(x[808]), .B(start), .Z(n427) );
  NAND U1671 ( .A(n429), .B(n430), .Z(xin[807]) );
  NANDN U1672 ( .A(start), .B(xreg[807]), .Z(n430) );
  NAND U1673 ( .A(x[807]), .B(start), .Z(n429) );
  NAND U1674 ( .A(n431), .B(n432), .Z(xin[806]) );
  NANDN U1675 ( .A(start), .B(xreg[806]), .Z(n432) );
  NAND U1676 ( .A(x[806]), .B(start), .Z(n431) );
  NAND U1677 ( .A(n433), .B(n434), .Z(xin[805]) );
  NANDN U1678 ( .A(start), .B(xreg[805]), .Z(n434) );
  NAND U1679 ( .A(x[805]), .B(start), .Z(n433) );
  NAND U1680 ( .A(n435), .B(n436), .Z(xin[804]) );
  NANDN U1681 ( .A(start), .B(xreg[804]), .Z(n436) );
  NAND U1682 ( .A(x[804]), .B(start), .Z(n435) );
  NAND U1683 ( .A(n437), .B(n438), .Z(xin[803]) );
  NANDN U1684 ( .A(start), .B(xreg[803]), .Z(n438) );
  NAND U1685 ( .A(x[803]), .B(start), .Z(n437) );
  NAND U1686 ( .A(n439), .B(n440), .Z(xin[802]) );
  NANDN U1687 ( .A(start), .B(xreg[802]), .Z(n440) );
  NAND U1688 ( .A(x[802]), .B(start), .Z(n439) );
  NAND U1689 ( .A(n441), .B(n442), .Z(xin[801]) );
  NANDN U1690 ( .A(start), .B(xreg[801]), .Z(n442) );
  NAND U1691 ( .A(x[801]), .B(start), .Z(n441) );
  NAND U1692 ( .A(n443), .B(n444), .Z(xin[800]) );
  NANDN U1693 ( .A(start), .B(xreg[800]), .Z(n444) );
  NAND U1694 ( .A(x[800]), .B(start), .Z(n443) );
  NAND U1695 ( .A(n445), .B(n446), .Z(xin[7]) );
  NANDN U1696 ( .A(start), .B(xreg[7]), .Z(n446) );
  NAND U1697 ( .A(x[7]), .B(start), .Z(n445) );
  NAND U1698 ( .A(n447), .B(n448), .Z(xin[79]) );
  NANDN U1699 ( .A(start), .B(xreg[79]), .Z(n448) );
  NAND U1700 ( .A(x[79]), .B(start), .Z(n447) );
  NAND U1701 ( .A(n449), .B(n450), .Z(xin[799]) );
  NANDN U1702 ( .A(start), .B(xreg[799]), .Z(n450) );
  NAND U1703 ( .A(x[799]), .B(start), .Z(n449) );
  NAND U1704 ( .A(n451), .B(n452), .Z(xin[798]) );
  NANDN U1705 ( .A(start), .B(xreg[798]), .Z(n452) );
  NAND U1706 ( .A(x[798]), .B(start), .Z(n451) );
  NAND U1707 ( .A(n453), .B(n454), .Z(xin[797]) );
  NANDN U1708 ( .A(start), .B(xreg[797]), .Z(n454) );
  NAND U1709 ( .A(x[797]), .B(start), .Z(n453) );
  NAND U1710 ( .A(n455), .B(n456), .Z(xin[796]) );
  NANDN U1711 ( .A(start), .B(xreg[796]), .Z(n456) );
  NAND U1712 ( .A(x[796]), .B(start), .Z(n455) );
  NAND U1713 ( .A(n457), .B(n458), .Z(xin[795]) );
  NANDN U1714 ( .A(start), .B(xreg[795]), .Z(n458) );
  NAND U1715 ( .A(x[795]), .B(start), .Z(n457) );
  NAND U1716 ( .A(n459), .B(n460), .Z(xin[794]) );
  NANDN U1717 ( .A(start), .B(xreg[794]), .Z(n460) );
  NAND U1718 ( .A(x[794]), .B(start), .Z(n459) );
  NAND U1719 ( .A(n461), .B(n462), .Z(xin[793]) );
  NANDN U1720 ( .A(start), .B(xreg[793]), .Z(n462) );
  NAND U1721 ( .A(x[793]), .B(start), .Z(n461) );
  NAND U1722 ( .A(n463), .B(n464), .Z(xin[792]) );
  NANDN U1723 ( .A(start), .B(xreg[792]), .Z(n464) );
  NAND U1724 ( .A(x[792]), .B(start), .Z(n463) );
  NAND U1725 ( .A(n465), .B(n466), .Z(xin[791]) );
  NANDN U1726 ( .A(start), .B(xreg[791]), .Z(n466) );
  NAND U1727 ( .A(x[791]), .B(start), .Z(n465) );
  NAND U1728 ( .A(n467), .B(n468), .Z(xin[790]) );
  NANDN U1729 ( .A(start), .B(xreg[790]), .Z(n468) );
  NAND U1730 ( .A(x[790]), .B(start), .Z(n467) );
  NAND U1731 ( .A(n469), .B(n470), .Z(xin[78]) );
  NANDN U1732 ( .A(start), .B(xreg[78]), .Z(n470) );
  NAND U1733 ( .A(x[78]), .B(start), .Z(n469) );
  NAND U1734 ( .A(n471), .B(n472), .Z(xin[789]) );
  NANDN U1735 ( .A(start), .B(xreg[789]), .Z(n472) );
  NAND U1736 ( .A(x[789]), .B(start), .Z(n471) );
  NAND U1737 ( .A(n473), .B(n474), .Z(xin[788]) );
  NANDN U1738 ( .A(start), .B(xreg[788]), .Z(n474) );
  NAND U1739 ( .A(x[788]), .B(start), .Z(n473) );
  NAND U1740 ( .A(n475), .B(n476), .Z(xin[787]) );
  NANDN U1741 ( .A(start), .B(xreg[787]), .Z(n476) );
  NAND U1742 ( .A(x[787]), .B(start), .Z(n475) );
  NAND U1743 ( .A(n477), .B(n478), .Z(xin[786]) );
  NANDN U1744 ( .A(start), .B(xreg[786]), .Z(n478) );
  NAND U1745 ( .A(x[786]), .B(start), .Z(n477) );
  NAND U1746 ( .A(n479), .B(n480), .Z(xin[785]) );
  NANDN U1747 ( .A(start), .B(xreg[785]), .Z(n480) );
  NAND U1748 ( .A(x[785]), .B(start), .Z(n479) );
  NAND U1749 ( .A(n481), .B(n482), .Z(xin[784]) );
  NANDN U1750 ( .A(start), .B(xreg[784]), .Z(n482) );
  NAND U1751 ( .A(x[784]), .B(start), .Z(n481) );
  NAND U1752 ( .A(n483), .B(n484), .Z(xin[783]) );
  NANDN U1753 ( .A(start), .B(xreg[783]), .Z(n484) );
  NAND U1754 ( .A(x[783]), .B(start), .Z(n483) );
  NAND U1755 ( .A(n485), .B(n486), .Z(xin[782]) );
  NANDN U1756 ( .A(start), .B(xreg[782]), .Z(n486) );
  NAND U1757 ( .A(x[782]), .B(start), .Z(n485) );
  NAND U1758 ( .A(n487), .B(n488), .Z(xin[781]) );
  NANDN U1759 ( .A(start), .B(xreg[781]), .Z(n488) );
  NAND U1760 ( .A(x[781]), .B(start), .Z(n487) );
  NAND U1761 ( .A(n489), .B(n490), .Z(xin[780]) );
  NANDN U1762 ( .A(start), .B(xreg[780]), .Z(n490) );
  NAND U1763 ( .A(x[780]), .B(start), .Z(n489) );
  NAND U1764 ( .A(n491), .B(n492), .Z(xin[77]) );
  NANDN U1765 ( .A(start), .B(xreg[77]), .Z(n492) );
  NAND U1766 ( .A(x[77]), .B(start), .Z(n491) );
  NAND U1767 ( .A(n493), .B(n494), .Z(xin[779]) );
  NANDN U1768 ( .A(start), .B(xreg[779]), .Z(n494) );
  NAND U1769 ( .A(x[779]), .B(start), .Z(n493) );
  NAND U1770 ( .A(n495), .B(n496), .Z(xin[778]) );
  NANDN U1771 ( .A(start), .B(xreg[778]), .Z(n496) );
  NAND U1772 ( .A(x[778]), .B(start), .Z(n495) );
  NAND U1773 ( .A(n497), .B(n498), .Z(xin[777]) );
  NANDN U1774 ( .A(start), .B(xreg[777]), .Z(n498) );
  NAND U1775 ( .A(x[777]), .B(start), .Z(n497) );
  NAND U1776 ( .A(n499), .B(n500), .Z(xin[776]) );
  NANDN U1777 ( .A(start), .B(xreg[776]), .Z(n500) );
  NAND U1778 ( .A(x[776]), .B(start), .Z(n499) );
  NAND U1779 ( .A(n501), .B(n502), .Z(xin[775]) );
  NANDN U1780 ( .A(start), .B(xreg[775]), .Z(n502) );
  NAND U1781 ( .A(x[775]), .B(start), .Z(n501) );
  NAND U1782 ( .A(n503), .B(n504), .Z(xin[774]) );
  NANDN U1783 ( .A(start), .B(xreg[774]), .Z(n504) );
  NAND U1784 ( .A(x[774]), .B(start), .Z(n503) );
  NAND U1785 ( .A(n505), .B(n506), .Z(xin[773]) );
  NANDN U1786 ( .A(start), .B(xreg[773]), .Z(n506) );
  NAND U1787 ( .A(x[773]), .B(start), .Z(n505) );
  NAND U1788 ( .A(n507), .B(n508), .Z(xin[772]) );
  NANDN U1789 ( .A(start), .B(xreg[772]), .Z(n508) );
  NAND U1790 ( .A(x[772]), .B(start), .Z(n507) );
  NAND U1791 ( .A(n509), .B(n510), .Z(xin[771]) );
  NANDN U1792 ( .A(start), .B(xreg[771]), .Z(n510) );
  NAND U1793 ( .A(x[771]), .B(start), .Z(n509) );
  NAND U1794 ( .A(n511), .B(n512), .Z(xin[770]) );
  NANDN U1795 ( .A(start), .B(xreg[770]), .Z(n512) );
  NAND U1796 ( .A(x[770]), .B(start), .Z(n511) );
  NAND U1797 ( .A(n513), .B(n514), .Z(xin[76]) );
  NANDN U1798 ( .A(start), .B(xreg[76]), .Z(n514) );
  NAND U1799 ( .A(x[76]), .B(start), .Z(n513) );
  NAND U1800 ( .A(n515), .B(n516), .Z(xin[769]) );
  NANDN U1801 ( .A(start), .B(xreg[769]), .Z(n516) );
  NAND U1802 ( .A(x[769]), .B(start), .Z(n515) );
  NAND U1803 ( .A(n517), .B(n518), .Z(xin[768]) );
  NANDN U1804 ( .A(start), .B(xreg[768]), .Z(n518) );
  NAND U1805 ( .A(x[768]), .B(start), .Z(n517) );
  NAND U1806 ( .A(n519), .B(n520), .Z(xin[767]) );
  NANDN U1807 ( .A(start), .B(xreg[767]), .Z(n520) );
  NAND U1808 ( .A(x[767]), .B(start), .Z(n519) );
  NAND U1809 ( .A(n521), .B(n522), .Z(xin[766]) );
  NANDN U1810 ( .A(start), .B(xreg[766]), .Z(n522) );
  NAND U1811 ( .A(x[766]), .B(start), .Z(n521) );
  NAND U1812 ( .A(n523), .B(n524), .Z(xin[765]) );
  NANDN U1813 ( .A(start), .B(xreg[765]), .Z(n524) );
  NAND U1814 ( .A(x[765]), .B(start), .Z(n523) );
  NAND U1815 ( .A(n525), .B(n526), .Z(xin[764]) );
  NANDN U1816 ( .A(start), .B(xreg[764]), .Z(n526) );
  NAND U1817 ( .A(x[764]), .B(start), .Z(n525) );
  NAND U1818 ( .A(n527), .B(n528), .Z(xin[763]) );
  NANDN U1819 ( .A(start), .B(xreg[763]), .Z(n528) );
  NAND U1820 ( .A(x[763]), .B(start), .Z(n527) );
  NAND U1821 ( .A(n529), .B(n530), .Z(xin[762]) );
  NANDN U1822 ( .A(start), .B(xreg[762]), .Z(n530) );
  NAND U1823 ( .A(x[762]), .B(start), .Z(n529) );
  NAND U1824 ( .A(n531), .B(n532), .Z(xin[761]) );
  NANDN U1825 ( .A(start), .B(xreg[761]), .Z(n532) );
  NAND U1826 ( .A(x[761]), .B(start), .Z(n531) );
  NAND U1827 ( .A(n533), .B(n534), .Z(xin[760]) );
  NANDN U1828 ( .A(start), .B(xreg[760]), .Z(n534) );
  NAND U1829 ( .A(x[760]), .B(start), .Z(n533) );
  NAND U1830 ( .A(n535), .B(n536), .Z(xin[75]) );
  NANDN U1831 ( .A(start), .B(xreg[75]), .Z(n536) );
  NAND U1832 ( .A(x[75]), .B(start), .Z(n535) );
  NAND U1833 ( .A(n537), .B(n538), .Z(xin[759]) );
  NANDN U1834 ( .A(start), .B(xreg[759]), .Z(n538) );
  NAND U1835 ( .A(x[759]), .B(start), .Z(n537) );
  NAND U1836 ( .A(n539), .B(n540), .Z(xin[758]) );
  NANDN U1837 ( .A(start), .B(xreg[758]), .Z(n540) );
  NAND U1838 ( .A(x[758]), .B(start), .Z(n539) );
  NAND U1839 ( .A(n541), .B(n542), .Z(xin[757]) );
  NANDN U1840 ( .A(start), .B(xreg[757]), .Z(n542) );
  NAND U1841 ( .A(x[757]), .B(start), .Z(n541) );
  NAND U1842 ( .A(n543), .B(n544), .Z(xin[756]) );
  NANDN U1843 ( .A(start), .B(xreg[756]), .Z(n544) );
  NAND U1844 ( .A(x[756]), .B(start), .Z(n543) );
  NAND U1845 ( .A(n545), .B(n546), .Z(xin[755]) );
  NANDN U1846 ( .A(start), .B(xreg[755]), .Z(n546) );
  NAND U1847 ( .A(x[755]), .B(start), .Z(n545) );
  NAND U1848 ( .A(n547), .B(n548), .Z(xin[754]) );
  NANDN U1849 ( .A(start), .B(xreg[754]), .Z(n548) );
  NAND U1850 ( .A(x[754]), .B(start), .Z(n547) );
  NAND U1851 ( .A(n549), .B(n550), .Z(xin[753]) );
  NANDN U1852 ( .A(start), .B(xreg[753]), .Z(n550) );
  NAND U1853 ( .A(x[753]), .B(start), .Z(n549) );
  NAND U1854 ( .A(n551), .B(n552), .Z(xin[752]) );
  NANDN U1855 ( .A(start), .B(xreg[752]), .Z(n552) );
  NAND U1856 ( .A(x[752]), .B(start), .Z(n551) );
  NAND U1857 ( .A(n553), .B(n554), .Z(xin[751]) );
  NANDN U1858 ( .A(start), .B(xreg[751]), .Z(n554) );
  NAND U1859 ( .A(x[751]), .B(start), .Z(n553) );
  NAND U1860 ( .A(n555), .B(n556), .Z(xin[750]) );
  NANDN U1861 ( .A(start), .B(xreg[750]), .Z(n556) );
  NAND U1862 ( .A(x[750]), .B(start), .Z(n555) );
  NAND U1863 ( .A(n557), .B(n558), .Z(xin[74]) );
  NANDN U1864 ( .A(start), .B(xreg[74]), .Z(n558) );
  NAND U1865 ( .A(x[74]), .B(start), .Z(n557) );
  NAND U1866 ( .A(n559), .B(n560), .Z(xin[749]) );
  NANDN U1867 ( .A(start), .B(xreg[749]), .Z(n560) );
  NAND U1868 ( .A(x[749]), .B(start), .Z(n559) );
  NAND U1869 ( .A(n561), .B(n562), .Z(xin[748]) );
  NANDN U1870 ( .A(start), .B(xreg[748]), .Z(n562) );
  NAND U1871 ( .A(x[748]), .B(start), .Z(n561) );
  NAND U1872 ( .A(n563), .B(n564), .Z(xin[747]) );
  NANDN U1873 ( .A(start), .B(xreg[747]), .Z(n564) );
  NAND U1874 ( .A(x[747]), .B(start), .Z(n563) );
  NAND U1875 ( .A(n565), .B(n566), .Z(xin[746]) );
  NANDN U1876 ( .A(start), .B(xreg[746]), .Z(n566) );
  NAND U1877 ( .A(x[746]), .B(start), .Z(n565) );
  NAND U1878 ( .A(n567), .B(n568), .Z(xin[745]) );
  NANDN U1879 ( .A(start), .B(xreg[745]), .Z(n568) );
  NAND U1880 ( .A(x[745]), .B(start), .Z(n567) );
  NAND U1881 ( .A(n569), .B(n570), .Z(xin[744]) );
  NANDN U1882 ( .A(start), .B(xreg[744]), .Z(n570) );
  NAND U1883 ( .A(x[744]), .B(start), .Z(n569) );
  NAND U1884 ( .A(n571), .B(n572), .Z(xin[743]) );
  NANDN U1885 ( .A(start), .B(xreg[743]), .Z(n572) );
  NAND U1886 ( .A(x[743]), .B(start), .Z(n571) );
  NAND U1887 ( .A(n573), .B(n574), .Z(xin[742]) );
  NANDN U1888 ( .A(start), .B(xreg[742]), .Z(n574) );
  NAND U1889 ( .A(x[742]), .B(start), .Z(n573) );
  NAND U1890 ( .A(n575), .B(n576), .Z(xin[741]) );
  NANDN U1891 ( .A(start), .B(xreg[741]), .Z(n576) );
  NAND U1892 ( .A(x[741]), .B(start), .Z(n575) );
  NAND U1893 ( .A(n577), .B(n578), .Z(xin[740]) );
  NANDN U1894 ( .A(start), .B(xreg[740]), .Z(n578) );
  NAND U1895 ( .A(x[740]), .B(start), .Z(n577) );
  NAND U1896 ( .A(n579), .B(n580), .Z(xin[73]) );
  NANDN U1897 ( .A(start), .B(xreg[73]), .Z(n580) );
  NAND U1898 ( .A(x[73]), .B(start), .Z(n579) );
  NAND U1899 ( .A(n581), .B(n582), .Z(xin[739]) );
  NANDN U1900 ( .A(start), .B(xreg[739]), .Z(n582) );
  NAND U1901 ( .A(x[739]), .B(start), .Z(n581) );
  NAND U1902 ( .A(n583), .B(n584), .Z(xin[738]) );
  NANDN U1903 ( .A(start), .B(xreg[738]), .Z(n584) );
  NAND U1904 ( .A(x[738]), .B(start), .Z(n583) );
  NAND U1905 ( .A(n585), .B(n586), .Z(xin[737]) );
  NANDN U1906 ( .A(start), .B(xreg[737]), .Z(n586) );
  NAND U1907 ( .A(x[737]), .B(start), .Z(n585) );
  NAND U1908 ( .A(n587), .B(n588), .Z(xin[736]) );
  NANDN U1909 ( .A(start), .B(xreg[736]), .Z(n588) );
  NAND U1910 ( .A(x[736]), .B(start), .Z(n587) );
  NAND U1911 ( .A(n589), .B(n590), .Z(xin[735]) );
  NANDN U1912 ( .A(start), .B(xreg[735]), .Z(n590) );
  NAND U1913 ( .A(x[735]), .B(start), .Z(n589) );
  NAND U1914 ( .A(n591), .B(n592), .Z(xin[734]) );
  NANDN U1915 ( .A(start), .B(xreg[734]), .Z(n592) );
  NAND U1916 ( .A(x[734]), .B(start), .Z(n591) );
  NAND U1917 ( .A(n593), .B(n594), .Z(xin[733]) );
  NANDN U1918 ( .A(start), .B(xreg[733]), .Z(n594) );
  NAND U1919 ( .A(x[733]), .B(start), .Z(n593) );
  NAND U1920 ( .A(n595), .B(n596), .Z(xin[732]) );
  NANDN U1921 ( .A(start), .B(xreg[732]), .Z(n596) );
  NAND U1922 ( .A(x[732]), .B(start), .Z(n595) );
  NAND U1923 ( .A(n597), .B(n598), .Z(xin[731]) );
  NANDN U1924 ( .A(start), .B(xreg[731]), .Z(n598) );
  NAND U1925 ( .A(x[731]), .B(start), .Z(n597) );
  NAND U1926 ( .A(n599), .B(n600), .Z(xin[730]) );
  NANDN U1927 ( .A(start), .B(xreg[730]), .Z(n600) );
  NAND U1928 ( .A(x[730]), .B(start), .Z(n599) );
  NAND U1929 ( .A(n601), .B(n602), .Z(xin[72]) );
  NANDN U1930 ( .A(start), .B(xreg[72]), .Z(n602) );
  NAND U1931 ( .A(x[72]), .B(start), .Z(n601) );
  NAND U1932 ( .A(n603), .B(n604), .Z(xin[729]) );
  NANDN U1933 ( .A(start), .B(xreg[729]), .Z(n604) );
  NAND U1934 ( .A(x[729]), .B(start), .Z(n603) );
  NAND U1935 ( .A(n605), .B(n606), .Z(xin[728]) );
  NANDN U1936 ( .A(start), .B(xreg[728]), .Z(n606) );
  NAND U1937 ( .A(x[728]), .B(start), .Z(n605) );
  NAND U1938 ( .A(n607), .B(n608), .Z(xin[727]) );
  NANDN U1939 ( .A(start), .B(xreg[727]), .Z(n608) );
  NAND U1940 ( .A(x[727]), .B(start), .Z(n607) );
  NAND U1941 ( .A(n609), .B(n610), .Z(xin[726]) );
  NANDN U1942 ( .A(start), .B(xreg[726]), .Z(n610) );
  NAND U1943 ( .A(x[726]), .B(start), .Z(n609) );
  NAND U1944 ( .A(n611), .B(n612), .Z(xin[725]) );
  NANDN U1945 ( .A(start), .B(xreg[725]), .Z(n612) );
  NAND U1946 ( .A(x[725]), .B(start), .Z(n611) );
  NAND U1947 ( .A(n613), .B(n614), .Z(xin[724]) );
  NANDN U1948 ( .A(start), .B(xreg[724]), .Z(n614) );
  NAND U1949 ( .A(x[724]), .B(start), .Z(n613) );
  NAND U1950 ( .A(n615), .B(n616), .Z(xin[723]) );
  NANDN U1951 ( .A(start), .B(xreg[723]), .Z(n616) );
  NAND U1952 ( .A(x[723]), .B(start), .Z(n615) );
  NAND U1953 ( .A(n617), .B(n618), .Z(xin[722]) );
  NANDN U1954 ( .A(start), .B(xreg[722]), .Z(n618) );
  NAND U1955 ( .A(x[722]), .B(start), .Z(n617) );
  NAND U1956 ( .A(n619), .B(n620), .Z(xin[721]) );
  NANDN U1957 ( .A(start), .B(xreg[721]), .Z(n620) );
  NAND U1958 ( .A(x[721]), .B(start), .Z(n619) );
  NAND U1959 ( .A(n621), .B(n622), .Z(xin[720]) );
  NANDN U1960 ( .A(start), .B(xreg[720]), .Z(n622) );
  NAND U1961 ( .A(x[720]), .B(start), .Z(n621) );
  NAND U1962 ( .A(n623), .B(n624), .Z(xin[71]) );
  NANDN U1963 ( .A(start), .B(xreg[71]), .Z(n624) );
  NAND U1964 ( .A(x[71]), .B(start), .Z(n623) );
  NAND U1965 ( .A(n625), .B(n626), .Z(xin[719]) );
  NANDN U1966 ( .A(start), .B(xreg[719]), .Z(n626) );
  NAND U1967 ( .A(x[719]), .B(start), .Z(n625) );
  NAND U1968 ( .A(n627), .B(n628), .Z(xin[718]) );
  NANDN U1969 ( .A(start), .B(xreg[718]), .Z(n628) );
  NAND U1970 ( .A(x[718]), .B(start), .Z(n627) );
  NAND U1971 ( .A(n629), .B(n630), .Z(xin[717]) );
  NANDN U1972 ( .A(start), .B(xreg[717]), .Z(n630) );
  NAND U1973 ( .A(x[717]), .B(start), .Z(n629) );
  NAND U1974 ( .A(n631), .B(n632), .Z(xin[716]) );
  NANDN U1975 ( .A(start), .B(xreg[716]), .Z(n632) );
  NAND U1976 ( .A(x[716]), .B(start), .Z(n631) );
  NAND U1977 ( .A(n633), .B(n634), .Z(xin[715]) );
  NANDN U1978 ( .A(start), .B(xreg[715]), .Z(n634) );
  NAND U1979 ( .A(x[715]), .B(start), .Z(n633) );
  NAND U1980 ( .A(n635), .B(n636), .Z(xin[714]) );
  NANDN U1981 ( .A(start), .B(xreg[714]), .Z(n636) );
  NAND U1982 ( .A(x[714]), .B(start), .Z(n635) );
  NAND U1983 ( .A(n637), .B(n638), .Z(xin[713]) );
  NANDN U1984 ( .A(start), .B(xreg[713]), .Z(n638) );
  NAND U1985 ( .A(x[713]), .B(start), .Z(n637) );
  NAND U1986 ( .A(n639), .B(n640), .Z(xin[712]) );
  NANDN U1987 ( .A(start), .B(xreg[712]), .Z(n640) );
  NAND U1988 ( .A(x[712]), .B(start), .Z(n639) );
  NAND U1989 ( .A(n641), .B(n642), .Z(xin[711]) );
  NANDN U1990 ( .A(start), .B(xreg[711]), .Z(n642) );
  NAND U1991 ( .A(x[711]), .B(start), .Z(n641) );
  NAND U1992 ( .A(n643), .B(n644), .Z(xin[710]) );
  NANDN U1993 ( .A(start), .B(xreg[710]), .Z(n644) );
  NAND U1994 ( .A(x[710]), .B(start), .Z(n643) );
  NAND U1995 ( .A(n645), .B(n646), .Z(xin[70]) );
  NANDN U1996 ( .A(start), .B(xreg[70]), .Z(n646) );
  NAND U1997 ( .A(x[70]), .B(start), .Z(n645) );
  NAND U1998 ( .A(n647), .B(n648), .Z(xin[709]) );
  NANDN U1999 ( .A(start), .B(xreg[709]), .Z(n648) );
  NAND U2000 ( .A(x[709]), .B(start), .Z(n647) );
  NAND U2001 ( .A(n649), .B(n650), .Z(xin[708]) );
  NANDN U2002 ( .A(start), .B(xreg[708]), .Z(n650) );
  NAND U2003 ( .A(x[708]), .B(start), .Z(n649) );
  NAND U2004 ( .A(n651), .B(n652), .Z(xin[707]) );
  NANDN U2005 ( .A(start), .B(xreg[707]), .Z(n652) );
  NAND U2006 ( .A(x[707]), .B(start), .Z(n651) );
  NAND U2007 ( .A(n653), .B(n654), .Z(xin[706]) );
  NANDN U2008 ( .A(start), .B(xreg[706]), .Z(n654) );
  NAND U2009 ( .A(x[706]), .B(start), .Z(n653) );
  NAND U2010 ( .A(n655), .B(n656), .Z(xin[705]) );
  NANDN U2011 ( .A(start), .B(xreg[705]), .Z(n656) );
  NAND U2012 ( .A(x[705]), .B(start), .Z(n655) );
  NAND U2013 ( .A(n657), .B(n658), .Z(xin[704]) );
  NANDN U2014 ( .A(start), .B(xreg[704]), .Z(n658) );
  NAND U2015 ( .A(x[704]), .B(start), .Z(n657) );
  NAND U2016 ( .A(n659), .B(n660), .Z(xin[703]) );
  NANDN U2017 ( .A(start), .B(xreg[703]), .Z(n660) );
  NAND U2018 ( .A(x[703]), .B(start), .Z(n659) );
  NAND U2019 ( .A(n661), .B(n662), .Z(xin[702]) );
  NANDN U2020 ( .A(start), .B(xreg[702]), .Z(n662) );
  NAND U2021 ( .A(x[702]), .B(start), .Z(n661) );
  NAND U2022 ( .A(n663), .B(n664), .Z(xin[701]) );
  NANDN U2023 ( .A(start), .B(xreg[701]), .Z(n664) );
  NAND U2024 ( .A(x[701]), .B(start), .Z(n663) );
  NAND U2025 ( .A(n665), .B(n666), .Z(xin[700]) );
  NANDN U2026 ( .A(start), .B(xreg[700]), .Z(n666) );
  NAND U2027 ( .A(x[700]), .B(start), .Z(n665) );
  NAND U2028 ( .A(n667), .B(n668), .Z(xin[6]) );
  NANDN U2029 ( .A(start), .B(xreg[6]), .Z(n668) );
  NAND U2030 ( .A(x[6]), .B(start), .Z(n667) );
  NAND U2031 ( .A(n669), .B(n670), .Z(xin[69]) );
  NANDN U2032 ( .A(start), .B(xreg[69]), .Z(n670) );
  NAND U2033 ( .A(x[69]), .B(start), .Z(n669) );
  NAND U2034 ( .A(n671), .B(n672), .Z(xin[699]) );
  NANDN U2035 ( .A(start), .B(xreg[699]), .Z(n672) );
  NAND U2036 ( .A(x[699]), .B(start), .Z(n671) );
  NAND U2037 ( .A(n673), .B(n674), .Z(xin[698]) );
  NANDN U2038 ( .A(start), .B(xreg[698]), .Z(n674) );
  NAND U2039 ( .A(x[698]), .B(start), .Z(n673) );
  NAND U2040 ( .A(n675), .B(n676), .Z(xin[697]) );
  NANDN U2041 ( .A(start), .B(xreg[697]), .Z(n676) );
  NAND U2042 ( .A(x[697]), .B(start), .Z(n675) );
  NAND U2043 ( .A(n677), .B(n678), .Z(xin[696]) );
  NANDN U2044 ( .A(start), .B(xreg[696]), .Z(n678) );
  NAND U2045 ( .A(x[696]), .B(start), .Z(n677) );
  NAND U2046 ( .A(n679), .B(n680), .Z(xin[695]) );
  NANDN U2047 ( .A(start), .B(xreg[695]), .Z(n680) );
  NAND U2048 ( .A(x[695]), .B(start), .Z(n679) );
  NAND U2049 ( .A(n681), .B(n682), .Z(xin[694]) );
  NANDN U2050 ( .A(start), .B(xreg[694]), .Z(n682) );
  NAND U2051 ( .A(x[694]), .B(start), .Z(n681) );
  NAND U2052 ( .A(n683), .B(n684), .Z(xin[693]) );
  NANDN U2053 ( .A(start), .B(xreg[693]), .Z(n684) );
  NAND U2054 ( .A(x[693]), .B(start), .Z(n683) );
  NAND U2055 ( .A(n685), .B(n686), .Z(xin[692]) );
  NANDN U2056 ( .A(start), .B(xreg[692]), .Z(n686) );
  NAND U2057 ( .A(x[692]), .B(start), .Z(n685) );
  NAND U2058 ( .A(n687), .B(n688), .Z(xin[691]) );
  NANDN U2059 ( .A(start), .B(xreg[691]), .Z(n688) );
  NAND U2060 ( .A(x[691]), .B(start), .Z(n687) );
  NAND U2061 ( .A(n689), .B(n690), .Z(xin[690]) );
  NANDN U2062 ( .A(start), .B(xreg[690]), .Z(n690) );
  NAND U2063 ( .A(x[690]), .B(start), .Z(n689) );
  NAND U2064 ( .A(n691), .B(n692), .Z(xin[68]) );
  NANDN U2065 ( .A(start), .B(xreg[68]), .Z(n692) );
  NAND U2066 ( .A(x[68]), .B(start), .Z(n691) );
  NAND U2067 ( .A(n693), .B(n694), .Z(xin[689]) );
  NANDN U2068 ( .A(start), .B(xreg[689]), .Z(n694) );
  NAND U2069 ( .A(x[689]), .B(start), .Z(n693) );
  NAND U2070 ( .A(n695), .B(n696), .Z(xin[688]) );
  NANDN U2071 ( .A(start), .B(xreg[688]), .Z(n696) );
  NAND U2072 ( .A(x[688]), .B(start), .Z(n695) );
  NAND U2073 ( .A(n697), .B(n698), .Z(xin[687]) );
  NANDN U2074 ( .A(start), .B(xreg[687]), .Z(n698) );
  NAND U2075 ( .A(x[687]), .B(start), .Z(n697) );
  NAND U2076 ( .A(n699), .B(n700), .Z(xin[686]) );
  NANDN U2077 ( .A(start), .B(xreg[686]), .Z(n700) );
  NAND U2078 ( .A(x[686]), .B(start), .Z(n699) );
  NAND U2079 ( .A(n701), .B(n702), .Z(xin[685]) );
  NANDN U2080 ( .A(start), .B(xreg[685]), .Z(n702) );
  NAND U2081 ( .A(x[685]), .B(start), .Z(n701) );
  NAND U2082 ( .A(n703), .B(n704), .Z(xin[684]) );
  NANDN U2083 ( .A(start), .B(xreg[684]), .Z(n704) );
  NAND U2084 ( .A(x[684]), .B(start), .Z(n703) );
  NAND U2085 ( .A(n705), .B(n706), .Z(xin[683]) );
  NANDN U2086 ( .A(start), .B(xreg[683]), .Z(n706) );
  NAND U2087 ( .A(x[683]), .B(start), .Z(n705) );
  NAND U2088 ( .A(n707), .B(n708), .Z(xin[682]) );
  NANDN U2089 ( .A(start), .B(xreg[682]), .Z(n708) );
  NAND U2090 ( .A(x[682]), .B(start), .Z(n707) );
  NAND U2091 ( .A(n709), .B(n710), .Z(xin[681]) );
  NANDN U2092 ( .A(start), .B(xreg[681]), .Z(n710) );
  NAND U2093 ( .A(x[681]), .B(start), .Z(n709) );
  NAND U2094 ( .A(n711), .B(n712), .Z(xin[680]) );
  NANDN U2095 ( .A(start), .B(xreg[680]), .Z(n712) );
  NAND U2096 ( .A(x[680]), .B(start), .Z(n711) );
  NAND U2097 ( .A(n713), .B(n714), .Z(xin[67]) );
  NANDN U2098 ( .A(start), .B(xreg[67]), .Z(n714) );
  NAND U2099 ( .A(x[67]), .B(start), .Z(n713) );
  NAND U2100 ( .A(n715), .B(n716), .Z(xin[679]) );
  NANDN U2101 ( .A(start), .B(xreg[679]), .Z(n716) );
  NAND U2102 ( .A(x[679]), .B(start), .Z(n715) );
  NAND U2103 ( .A(n717), .B(n718), .Z(xin[678]) );
  NANDN U2104 ( .A(start), .B(xreg[678]), .Z(n718) );
  NAND U2105 ( .A(x[678]), .B(start), .Z(n717) );
  NAND U2106 ( .A(n719), .B(n720), .Z(xin[677]) );
  NANDN U2107 ( .A(start), .B(xreg[677]), .Z(n720) );
  NAND U2108 ( .A(x[677]), .B(start), .Z(n719) );
  NAND U2109 ( .A(n721), .B(n722), .Z(xin[676]) );
  NANDN U2110 ( .A(start), .B(xreg[676]), .Z(n722) );
  NAND U2111 ( .A(x[676]), .B(start), .Z(n721) );
  NAND U2112 ( .A(n723), .B(n724), .Z(xin[675]) );
  NANDN U2113 ( .A(start), .B(xreg[675]), .Z(n724) );
  NAND U2114 ( .A(x[675]), .B(start), .Z(n723) );
  NAND U2115 ( .A(n725), .B(n726), .Z(xin[674]) );
  NANDN U2116 ( .A(start), .B(xreg[674]), .Z(n726) );
  NAND U2117 ( .A(x[674]), .B(start), .Z(n725) );
  NAND U2118 ( .A(n727), .B(n728), .Z(xin[673]) );
  NANDN U2119 ( .A(start), .B(xreg[673]), .Z(n728) );
  NAND U2120 ( .A(x[673]), .B(start), .Z(n727) );
  NAND U2121 ( .A(n729), .B(n730), .Z(xin[672]) );
  NANDN U2122 ( .A(start), .B(xreg[672]), .Z(n730) );
  NAND U2123 ( .A(x[672]), .B(start), .Z(n729) );
  NAND U2124 ( .A(n731), .B(n732), .Z(xin[671]) );
  NANDN U2125 ( .A(start), .B(xreg[671]), .Z(n732) );
  NAND U2126 ( .A(x[671]), .B(start), .Z(n731) );
  NAND U2127 ( .A(n733), .B(n734), .Z(xin[670]) );
  NANDN U2128 ( .A(start), .B(xreg[670]), .Z(n734) );
  NAND U2129 ( .A(x[670]), .B(start), .Z(n733) );
  NAND U2130 ( .A(n735), .B(n736), .Z(xin[66]) );
  NANDN U2131 ( .A(start), .B(xreg[66]), .Z(n736) );
  NAND U2132 ( .A(x[66]), .B(start), .Z(n735) );
  NAND U2133 ( .A(n737), .B(n738), .Z(xin[669]) );
  NANDN U2134 ( .A(start), .B(xreg[669]), .Z(n738) );
  NAND U2135 ( .A(x[669]), .B(start), .Z(n737) );
  NAND U2136 ( .A(n739), .B(n740), .Z(xin[668]) );
  NANDN U2137 ( .A(start), .B(xreg[668]), .Z(n740) );
  NAND U2138 ( .A(x[668]), .B(start), .Z(n739) );
  NAND U2139 ( .A(n741), .B(n742), .Z(xin[667]) );
  NANDN U2140 ( .A(start), .B(xreg[667]), .Z(n742) );
  NAND U2141 ( .A(x[667]), .B(start), .Z(n741) );
  NAND U2142 ( .A(n743), .B(n744), .Z(xin[666]) );
  NANDN U2143 ( .A(start), .B(xreg[666]), .Z(n744) );
  NAND U2144 ( .A(x[666]), .B(start), .Z(n743) );
  NAND U2145 ( .A(n745), .B(n746), .Z(xin[665]) );
  NANDN U2146 ( .A(start), .B(xreg[665]), .Z(n746) );
  NAND U2147 ( .A(x[665]), .B(start), .Z(n745) );
  NAND U2148 ( .A(n747), .B(n748), .Z(xin[664]) );
  NANDN U2149 ( .A(start), .B(xreg[664]), .Z(n748) );
  NAND U2150 ( .A(x[664]), .B(start), .Z(n747) );
  NAND U2151 ( .A(n749), .B(n750), .Z(xin[663]) );
  NANDN U2152 ( .A(start), .B(xreg[663]), .Z(n750) );
  NAND U2153 ( .A(x[663]), .B(start), .Z(n749) );
  NAND U2154 ( .A(n751), .B(n752), .Z(xin[662]) );
  NANDN U2155 ( .A(start), .B(xreg[662]), .Z(n752) );
  NAND U2156 ( .A(x[662]), .B(start), .Z(n751) );
  NAND U2157 ( .A(n753), .B(n754), .Z(xin[661]) );
  NANDN U2158 ( .A(start), .B(xreg[661]), .Z(n754) );
  NAND U2159 ( .A(x[661]), .B(start), .Z(n753) );
  NAND U2160 ( .A(n755), .B(n756), .Z(xin[660]) );
  NANDN U2161 ( .A(start), .B(xreg[660]), .Z(n756) );
  NAND U2162 ( .A(x[660]), .B(start), .Z(n755) );
  NAND U2163 ( .A(n757), .B(n758), .Z(xin[65]) );
  NANDN U2164 ( .A(start), .B(xreg[65]), .Z(n758) );
  NAND U2165 ( .A(x[65]), .B(start), .Z(n757) );
  NAND U2166 ( .A(n759), .B(n760), .Z(xin[659]) );
  NANDN U2167 ( .A(start), .B(xreg[659]), .Z(n760) );
  NAND U2168 ( .A(x[659]), .B(start), .Z(n759) );
  NAND U2169 ( .A(n761), .B(n762), .Z(xin[658]) );
  NANDN U2170 ( .A(start), .B(xreg[658]), .Z(n762) );
  NAND U2171 ( .A(x[658]), .B(start), .Z(n761) );
  NAND U2172 ( .A(n763), .B(n764), .Z(xin[657]) );
  NANDN U2173 ( .A(start), .B(xreg[657]), .Z(n764) );
  NAND U2174 ( .A(x[657]), .B(start), .Z(n763) );
  NAND U2175 ( .A(n765), .B(n766), .Z(xin[656]) );
  NANDN U2176 ( .A(start), .B(xreg[656]), .Z(n766) );
  NAND U2177 ( .A(x[656]), .B(start), .Z(n765) );
  NAND U2178 ( .A(n767), .B(n768), .Z(xin[655]) );
  NANDN U2179 ( .A(start), .B(xreg[655]), .Z(n768) );
  NAND U2180 ( .A(x[655]), .B(start), .Z(n767) );
  NAND U2181 ( .A(n769), .B(n770), .Z(xin[654]) );
  NANDN U2182 ( .A(start), .B(xreg[654]), .Z(n770) );
  NAND U2183 ( .A(x[654]), .B(start), .Z(n769) );
  NAND U2184 ( .A(n771), .B(n772), .Z(xin[653]) );
  NANDN U2185 ( .A(start), .B(xreg[653]), .Z(n772) );
  NAND U2186 ( .A(x[653]), .B(start), .Z(n771) );
  NAND U2187 ( .A(n773), .B(n774), .Z(xin[652]) );
  NANDN U2188 ( .A(start), .B(xreg[652]), .Z(n774) );
  NAND U2189 ( .A(x[652]), .B(start), .Z(n773) );
  NAND U2190 ( .A(n775), .B(n776), .Z(xin[651]) );
  NANDN U2191 ( .A(start), .B(xreg[651]), .Z(n776) );
  NAND U2192 ( .A(x[651]), .B(start), .Z(n775) );
  NAND U2193 ( .A(n777), .B(n778), .Z(xin[650]) );
  NANDN U2194 ( .A(start), .B(xreg[650]), .Z(n778) );
  NAND U2195 ( .A(x[650]), .B(start), .Z(n777) );
  NAND U2196 ( .A(n779), .B(n780), .Z(xin[64]) );
  NANDN U2197 ( .A(start), .B(xreg[64]), .Z(n780) );
  NAND U2198 ( .A(x[64]), .B(start), .Z(n779) );
  NAND U2199 ( .A(n781), .B(n782), .Z(xin[649]) );
  NANDN U2200 ( .A(start), .B(xreg[649]), .Z(n782) );
  NAND U2201 ( .A(x[649]), .B(start), .Z(n781) );
  NAND U2202 ( .A(n783), .B(n784), .Z(xin[648]) );
  NANDN U2203 ( .A(start), .B(xreg[648]), .Z(n784) );
  NAND U2204 ( .A(x[648]), .B(start), .Z(n783) );
  NAND U2205 ( .A(n785), .B(n786), .Z(xin[647]) );
  NANDN U2206 ( .A(start), .B(xreg[647]), .Z(n786) );
  NAND U2207 ( .A(x[647]), .B(start), .Z(n785) );
  NAND U2208 ( .A(n787), .B(n788), .Z(xin[646]) );
  NANDN U2209 ( .A(start), .B(xreg[646]), .Z(n788) );
  NAND U2210 ( .A(x[646]), .B(start), .Z(n787) );
  NAND U2211 ( .A(n789), .B(n790), .Z(xin[645]) );
  NANDN U2212 ( .A(start), .B(xreg[645]), .Z(n790) );
  NAND U2213 ( .A(x[645]), .B(start), .Z(n789) );
  NAND U2214 ( .A(n791), .B(n792), .Z(xin[644]) );
  NANDN U2215 ( .A(start), .B(xreg[644]), .Z(n792) );
  NAND U2216 ( .A(x[644]), .B(start), .Z(n791) );
  NAND U2217 ( .A(n793), .B(n794), .Z(xin[643]) );
  NANDN U2218 ( .A(start), .B(xreg[643]), .Z(n794) );
  NAND U2219 ( .A(x[643]), .B(start), .Z(n793) );
  NAND U2220 ( .A(n795), .B(n796), .Z(xin[642]) );
  NANDN U2221 ( .A(start), .B(xreg[642]), .Z(n796) );
  NAND U2222 ( .A(x[642]), .B(start), .Z(n795) );
  NAND U2223 ( .A(n797), .B(n798), .Z(xin[641]) );
  NANDN U2224 ( .A(start), .B(xreg[641]), .Z(n798) );
  NAND U2225 ( .A(x[641]), .B(start), .Z(n797) );
  NAND U2226 ( .A(n799), .B(n800), .Z(xin[640]) );
  NANDN U2227 ( .A(start), .B(xreg[640]), .Z(n800) );
  NAND U2228 ( .A(x[640]), .B(start), .Z(n799) );
  NAND U2229 ( .A(n801), .B(n802), .Z(xin[63]) );
  NANDN U2230 ( .A(start), .B(xreg[63]), .Z(n802) );
  NAND U2231 ( .A(x[63]), .B(start), .Z(n801) );
  NAND U2232 ( .A(n803), .B(n804), .Z(xin[639]) );
  NANDN U2233 ( .A(start), .B(xreg[639]), .Z(n804) );
  NAND U2234 ( .A(x[639]), .B(start), .Z(n803) );
  NAND U2235 ( .A(n805), .B(n806), .Z(xin[638]) );
  NANDN U2236 ( .A(start), .B(xreg[638]), .Z(n806) );
  NAND U2237 ( .A(x[638]), .B(start), .Z(n805) );
  NAND U2238 ( .A(n807), .B(n808), .Z(xin[637]) );
  NANDN U2239 ( .A(start), .B(xreg[637]), .Z(n808) );
  NAND U2240 ( .A(x[637]), .B(start), .Z(n807) );
  NAND U2241 ( .A(n809), .B(n810), .Z(xin[636]) );
  NANDN U2242 ( .A(start), .B(xreg[636]), .Z(n810) );
  NAND U2243 ( .A(x[636]), .B(start), .Z(n809) );
  NAND U2244 ( .A(n811), .B(n812), .Z(xin[635]) );
  NANDN U2245 ( .A(start), .B(xreg[635]), .Z(n812) );
  NAND U2246 ( .A(x[635]), .B(start), .Z(n811) );
  NAND U2247 ( .A(n813), .B(n814), .Z(xin[634]) );
  NANDN U2248 ( .A(start), .B(xreg[634]), .Z(n814) );
  NAND U2249 ( .A(x[634]), .B(start), .Z(n813) );
  NAND U2250 ( .A(n815), .B(n816), .Z(xin[633]) );
  NANDN U2251 ( .A(start), .B(xreg[633]), .Z(n816) );
  NAND U2252 ( .A(x[633]), .B(start), .Z(n815) );
  NAND U2253 ( .A(n817), .B(n818), .Z(xin[632]) );
  NANDN U2254 ( .A(start), .B(xreg[632]), .Z(n818) );
  NAND U2255 ( .A(x[632]), .B(start), .Z(n817) );
  NAND U2256 ( .A(n819), .B(n820), .Z(xin[631]) );
  NANDN U2257 ( .A(start), .B(xreg[631]), .Z(n820) );
  NAND U2258 ( .A(x[631]), .B(start), .Z(n819) );
  NAND U2259 ( .A(n821), .B(n822), .Z(xin[630]) );
  NANDN U2260 ( .A(start), .B(xreg[630]), .Z(n822) );
  NAND U2261 ( .A(x[630]), .B(start), .Z(n821) );
  NAND U2262 ( .A(n823), .B(n824), .Z(xin[62]) );
  NANDN U2263 ( .A(start), .B(xreg[62]), .Z(n824) );
  NAND U2264 ( .A(x[62]), .B(start), .Z(n823) );
  NAND U2265 ( .A(n825), .B(n826), .Z(xin[629]) );
  NANDN U2266 ( .A(start), .B(xreg[629]), .Z(n826) );
  NAND U2267 ( .A(x[629]), .B(start), .Z(n825) );
  NAND U2268 ( .A(n827), .B(n828), .Z(xin[628]) );
  NANDN U2269 ( .A(start), .B(xreg[628]), .Z(n828) );
  NAND U2270 ( .A(x[628]), .B(start), .Z(n827) );
  NAND U2271 ( .A(n829), .B(n830), .Z(xin[627]) );
  NANDN U2272 ( .A(start), .B(xreg[627]), .Z(n830) );
  NAND U2273 ( .A(x[627]), .B(start), .Z(n829) );
  NAND U2274 ( .A(n831), .B(n832), .Z(xin[626]) );
  NANDN U2275 ( .A(start), .B(xreg[626]), .Z(n832) );
  NAND U2276 ( .A(x[626]), .B(start), .Z(n831) );
  NAND U2277 ( .A(n833), .B(n834), .Z(xin[625]) );
  NANDN U2278 ( .A(start), .B(xreg[625]), .Z(n834) );
  NAND U2279 ( .A(x[625]), .B(start), .Z(n833) );
  NAND U2280 ( .A(n835), .B(n836), .Z(xin[624]) );
  NANDN U2281 ( .A(start), .B(xreg[624]), .Z(n836) );
  NAND U2282 ( .A(x[624]), .B(start), .Z(n835) );
  NAND U2283 ( .A(n837), .B(n838), .Z(xin[623]) );
  NANDN U2284 ( .A(start), .B(xreg[623]), .Z(n838) );
  NAND U2285 ( .A(x[623]), .B(start), .Z(n837) );
  NAND U2286 ( .A(n839), .B(n840), .Z(xin[622]) );
  NANDN U2287 ( .A(start), .B(xreg[622]), .Z(n840) );
  NAND U2288 ( .A(x[622]), .B(start), .Z(n839) );
  NAND U2289 ( .A(n841), .B(n842), .Z(xin[621]) );
  NANDN U2290 ( .A(start), .B(xreg[621]), .Z(n842) );
  NAND U2291 ( .A(x[621]), .B(start), .Z(n841) );
  NAND U2292 ( .A(n843), .B(n844), .Z(xin[620]) );
  NANDN U2293 ( .A(start), .B(xreg[620]), .Z(n844) );
  NAND U2294 ( .A(x[620]), .B(start), .Z(n843) );
  NAND U2295 ( .A(n845), .B(n846), .Z(xin[61]) );
  NANDN U2296 ( .A(start), .B(xreg[61]), .Z(n846) );
  NAND U2297 ( .A(x[61]), .B(start), .Z(n845) );
  NAND U2298 ( .A(n847), .B(n848), .Z(xin[619]) );
  NANDN U2299 ( .A(start), .B(xreg[619]), .Z(n848) );
  NAND U2300 ( .A(x[619]), .B(start), .Z(n847) );
  NAND U2301 ( .A(n849), .B(n850), .Z(xin[618]) );
  NANDN U2302 ( .A(start), .B(xreg[618]), .Z(n850) );
  NAND U2303 ( .A(x[618]), .B(start), .Z(n849) );
  NAND U2304 ( .A(n851), .B(n852), .Z(xin[617]) );
  NANDN U2305 ( .A(start), .B(xreg[617]), .Z(n852) );
  NAND U2306 ( .A(x[617]), .B(start), .Z(n851) );
  NAND U2307 ( .A(n853), .B(n854), .Z(xin[616]) );
  NANDN U2308 ( .A(start), .B(xreg[616]), .Z(n854) );
  NAND U2309 ( .A(x[616]), .B(start), .Z(n853) );
  NAND U2310 ( .A(n855), .B(n856), .Z(xin[615]) );
  NANDN U2311 ( .A(start), .B(xreg[615]), .Z(n856) );
  NAND U2312 ( .A(x[615]), .B(start), .Z(n855) );
  NAND U2313 ( .A(n857), .B(n858), .Z(xin[614]) );
  NANDN U2314 ( .A(start), .B(xreg[614]), .Z(n858) );
  NAND U2315 ( .A(x[614]), .B(start), .Z(n857) );
  NAND U2316 ( .A(n859), .B(n860), .Z(xin[613]) );
  NANDN U2317 ( .A(start), .B(xreg[613]), .Z(n860) );
  NAND U2318 ( .A(x[613]), .B(start), .Z(n859) );
  NAND U2319 ( .A(n861), .B(n862), .Z(xin[612]) );
  NANDN U2320 ( .A(start), .B(xreg[612]), .Z(n862) );
  NAND U2321 ( .A(x[612]), .B(start), .Z(n861) );
  NAND U2322 ( .A(n863), .B(n864), .Z(xin[611]) );
  NANDN U2323 ( .A(start), .B(xreg[611]), .Z(n864) );
  NAND U2324 ( .A(x[611]), .B(start), .Z(n863) );
  NAND U2325 ( .A(n865), .B(n866), .Z(xin[610]) );
  NANDN U2326 ( .A(start), .B(xreg[610]), .Z(n866) );
  NAND U2327 ( .A(x[610]), .B(start), .Z(n865) );
  NAND U2328 ( .A(n867), .B(n868), .Z(xin[60]) );
  NANDN U2329 ( .A(start), .B(xreg[60]), .Z(n868) );
  NAND U2330 ( .A(x[60]), .B(start), .Z(n867) );
  NAND U2331 ( .A(n869), .B(n870), .Z(xin[609]) );
  NANDN U2332 ( .A(start), .B(xreg[609]), .Z(n870) );
  NAND U2333 ( .A(x[609]), .B(start), .Z(n869) );
  NAND U2334 ( .A(n871), .B(n872), .Z(xin[608]) );
  NANDN U2335 ( .A(start), .B(xreg[608]), .Z(n872) );
  NAND U2336 ( .A(x[608]), .B(start), .Z(n871) );
  NAND U2337 ( .A(n873), .B(n874), .Z(xin[607]) );
  NANDN U2338 ( .A(start), .B(xreg[607]), .Z(n874) );
  NAND U2339 ( .A(x[607]), .B(start), .Z(n873) );
  NAND U2340 ( .A(n875), .B(n876), .Z(xin[606]) );
  NANDN U2341 ( .A(start), .B(xreg[606]), .Z(n876) );
  NAND U2342 ( .A(x[606]), .B(start), .Z(n875) );
  NAND U2343 ( .A(n877), .B(n878), .Z(xin[605]) );
  NANDN U2344 ( .A(start), .B(xreg[605]), .Z(n878) );
  NAND U2345 ( .A(x[605]), .B(start), .Z(n877) );
  NAND U2346 ( .A(n879), .B(n880), .Z(xin[604]) );
  NANDN U2347 ( .A(start), .B(xreg[604]), .Z(n880) );
  NAND U2348 ( .A(x[604]), .B(start), .Z(n879) );
  NAND U2349 ( .A(n881), .B(n882), .Z(xin[603]) );
  NANDN U2350 ( .A(start), .B(xreg[603]), .Z(n882) );
  NAND U2351 ( .A(x[603]), .B(start), .Z(n881) );
  NAND U2352 ( .A(n883), .B(n884), .Z(xin[602]) );
  NANDN U2353 ( .A(start), .B(xreg[602]), .Z(n884) );
  NAND U2354 ( .A(x[602]), .B(start), .Z(n883) );
  NAND U2355 ( .A(n885), .B(n886), .Z(xin[601]) );
  NANDN U2356 ( .A(start), .B(xreg[601]), .Z(n886) );
  NAND U2357 ( .A(x[601]), .B(start), .Z(n885) );
  NAND U2358 ( .A(n887), .B(n888), .Z(xin[600]) );
  NANDN U2359 ( .A(start), .B(xreg[600]), .Z(n888) );
  NAND U2360 ( .A(x[600]), .B(start), .Z(n887) );
  NAND U2361 ( .A(n889), .B(n890), .Z(xin[5]) );
  NANDN U2362 ( .A(start), .B(xreg[5]), .Z(n890) );
  NAND U2363 ( .A(x[5]), .B(start), .Z(n889) );
  NAND U2364 ( .A(n891), .B(n892), .Z(xin[59]) );
  NANDN U2365 ( .A(start), .B(xreg[59]), .Z(n892) );
  NAND U2366 ( .A(x[59]), .B(start), .Z(n891) );
  NAND U2367 ( .A(n893), .B(n894), .Z(xin[599]) );
  NANDN U2368 ( .A(start), .B(xreg[599]), .Z(n894) );
  NAND U2369 ( .A(x[599]), .B(start), .Z(n893) );
  NAND U2370 ( .A(n895), .B(n896), .Z(xin[598]) );
  NANDN U2371 ( .A(start), .B(xreg[598]), .Z(n896) );
  NAND U2372 ( .A(x[598]), .B(start), .Z(n895) );
  NAND U2373 ( .A(n897), .B(n898), .Z(xin[597]) );
  NANDN U2374 ( .A(start), .B(xreg[597]), .Z(n898) );
  NAND U2375 ( .A(x[597]), .B(start), .Z(n897) );
  NAND U2376 ( .A(n899), .B(n900), .Z(xin[596]) );
  NANDN U2377 ( .A(start), .B(xreg[596]), .Z(n900) );
  NAND U2378 ( .A(x[596]), .B(start), .Z(n899) );
  NAND U2379 ( .A(n901), .B(n902), .Z(xin[595]) );
  NANDN U2380 ( .A(start), .B(xreg[595]), .Z(n902) );
  NAND U2381 ( .A(x[595]), .B(start), .Z(n901) );
  NAND U2382 ( .A(n903), .B(n904), .Z(xin[594]) );
  NANDN U2383 ( .A(start), .B(xreg[594]), .Z(n904) );
  NAND U2384 ( .A(x[594]), .B(start), .Z(n903) );
  NAND U2385 ( .A(n905), .B(n906), .Z(xin[593]) );
  NANDN U2386 ( .A(start), .B(xreg[593]), .Z(n906) );
  NAND U2387 ( .A(x[593]), .B(start), .Z(n905) );
  NAND U2388 ( .A(n907), .B(n908), .Z(xin[592]) );
  NANDN U2389 ( .A(start), .B(xreg[592]), .Z(n908) );
  NAND U2390 ( .A(x[592]), .B(start), .Z(n907) );
  NAND U2391 ( .A(n909), .B(n910), .Z(xin[591]) );
  NANDN U2392 ( .A(start), .B(xreg[591]), .Z(n910) );
  NAND U2393 ( .A(x[591]), .B(start), .Z(n909) );
  NAND U2394 ( .A(n911), .B(n912), .Z(xin[590]) );
  NANDN U2395 ( .A(start), .B(xreg[590]), .Z(n912) );
  NAND U2396 ( .A(x[590]), .B(start), .Z(n911) );
  NAND U2397 ( .A(n913), .B(n914), .Z(xin[58]) );
  NANDN U2398 ( .A(start), .B(xreg[58]), .Z(n914) );
  NAND U2399 ( .A(x[58]), .B(start), .Z(n913) );
  NAND U2400 ( .A(n915), .B(n916), .Z(xin[589]) );
  NANDN U2401 ( .A(start), .B(xreg[589]), .Z(n916) );
  NAND U2402 ( .A(x[589]), .B(start), .Z(n915) );
  NAND U2403 ( .A(n917), .B(n918), .Z(xin[588]) );
  NANDN U2404 ( .A(start), .B(xreg[588]), .Z(n918) );
  NAND U2405 ( .A(x[588]), .B(start), .Z(n917) );
  NAND U2406 ( .A(n919), .B(n920), .Z(xin[587]) );
  NANDN U2407 ( .A(start), .B(xreg[587]), .Z(n920) );
  NAND U2408 ( .A(x[587]), .B(start), .Z(n919) );
  NAND U2409 ( .A(n921), .B(n922), .Z(xin[586]) );
  NANDN U2410 ( .A(start), .B(xreg[586]), .Z(n922) );
  NAND U2411 ( .A(x[586]), .B(start), .Z(n921) );
  NAND U2412 ( .A(n923), .B(n924), .Z(xin[585]) );
  NANDN U2413 ( .A(start), .B(xreg[585]), .Z(n924) );
  NAND U2414 ( .A(x[585]), .B(start), .Z(n923) );
  NAND U2415 ( .A(n925), .B(n926), .Z(xin[584]) );
  NANDN U2416 ( .A(start), .B(xreg[584]), .Z(n926) );
  NAND U2417 ( .A(x[584]), .B(start), .Z(n925) );
  NAND U2418 ( .A(n927), .B(n928), .Z(xin[583]) );
  NANDN U2419 ( .A(start), .B(xreg[583]), .Z(n928) );
  NAND U2420 ( .A(x[583]), .B(start), .Z(n927) );
  NAND U2421 ( .A(n929), .B(n930), .Z(xin[582]) );
  NANDN U2422 ( .A(start), .B(xreg[582]), .Z(n930) );
  NAND U2423 ( .A(x[582]), .B(start), .Z(n929) );
  NAND U2424 ( .A(n931), .B(n932), .Z(xin[581]) );
  NANDN U2425 ( .A(start), .B(xreg[581]), .Z(n932) );
  NAND U2426 ( .A(x[581]), .B(start), .Z(n931) );
  NAND U2427 ( .A(n933), .B(n934), .Z(xin[580]) );
  NANDN U2428 ( .A(start), .B(xreg[580]), .Z(n934) );
  NAND U2429 ( .A(x[580]), .B(start), .Z(n933) );
  NAND U2430 ( .A(n935), .B(n936), .Z(xin[57]) );
  NANDN U2431 ( .A(start), .B(xreg[57]), .Z(n936) );
  NAND U2432 ( .A(x[57]), .B(start), .Z(n935) );
  NAND U2433 ( .A(n937), .B(n938), .Z(xin[579]) );
  NANDN U2434 ( .A(start), .B(xreg[579]), .Z(n938) );
  NAND U2435 ( .A(x[579]), .B(start), .Z(n937) );
  NAND U2436 ( .A(n939), .B(n940), .Z(xin[578]) );
  NANDN U2437 ( .A(start), .B(xreg[578]), .Z(n940) );
  NAND U2438 ( .A(x[578]), .B(start), .Z(n939) );
  NAND U2439 ( .A(n941), .B(n942), .Z(xin[577]) );
  NANDN U2440 ( .A(start), .B(xreg[577]), .Z(n942) );
  NAND U2441 ( .A(x[577]), .B(start), .Z(n941) );
  NAND U2442 ( .A(n943), .B(n944), .Z(xin[576]) );
  NANDN U2443 ( .A(start), .B(xreg[576]), .Z(n944) );
  NAND U2444 ( .A(x[576]), .B(start), .Z(n943) );
  NAND U2445 ( .A(n945), .B(n946), .Z(xin[575]) );
  NANDN U2446 ( .A(start), .B(xreg[575]), .Z(n946) );
  NAND U2447 ( .A(x[575]), .B(start), .Z(n945) );
  NAND U2448 ( .A(n947), .B(n948), .Z(xin[574]) );
  NANDN U2449 ( .A(start), .B(xreg[574]), .Z(n948) );
  NAND U2450 ( .A(x[574]), .B(start), .Z(n947) );
  NAND U2451 ( .A(n949), .B(n950), .Z(xin[573]) );
  NANDN U2452 ( .A(start), .B(xreg[573]), .Z(n950) );
  NAND U2453 ( .A(x[573]), .B(start), .Z(n949) );
  NAND U2454 ( .A(n951), .B(n952), .Z(xin[572]) );
  NANDN U2455 ( .A(start), .B(xreg[572]), .Z(n952) );
  NAND U2456 ( .A(x[572]), .B(start), .Z(n951) );
  NAND U2457 ( .A(n953), .B(n954), .Z(xin[571]) );
  NANDN U2458 ( .A(start), .B(xreg[571]), .Z(n954) );
  NAND U2459 ( .A(x[571]), .B(start), .Z(n953) );
  NAND U2460 ( .A(n955), .B(n956), .Z(xin[570]) );
  NANDN U2461 ( .A(start), .B(xreg[570]), .Z(n956) );
  NAND U2462 ( .A(x[570]), .B(start), .Z(n955) );
  NAND U2463 ( .A(n957), .B(n958), .Z(xin[56]) );
  NANDN U2464 ( .A(start), .B(xreg[56]), .Z(n958) );
  NAND U2465 ( .A(x[56]), .B(start), .Z(n957) );
  NAND U2466 ( .A(n959), .B(n960), .Z(xin[569]) );
  NANDN U2467 ( .A(start), .B(xreg[569]), .Z(n960) );
  NAND U2468 ( .A(x[569]), .B(start), .Z(n959) );
  NAND U2469 ( .A(n961), .B(n962), .Z(xin[568]) );
  NANDN U2470 ( .A(start), .B(xreg[568]), .Z(n962) );
  NAND U2471 ( .A(x[568]), .B(start), .Z(n961) );
  NAND U2472 ( .A(n963), .B(n964), .Z(xin[567]) );
  NANDN U2473 ( .A(start), .B(xreg[567]), .Z(n964) );
  NAND U2474 ( .A(x[567]), .B(start), .Z(n963) );
  NAND U2475 ( .A(n965), .B(n966), .Z(xin[566]) );
  NANDN U2476 ( .A(start), .B(xreg[566]), .Z(n966) );
  NAND U2477 ( .A(x[566]), .B(start), .Z(n965) );
  NAND U2478 ( .A(n967), .B(n968), .Z(xin[565]) );
  NANDN U2479 ( .A(start), .B(xreg[565]), .Z(n968) );
  NAND U2480 ( .A(x[565]), .B(start), .Z(n967) );
  NAND U2481 ( .A(n969), .B(n970), .Z(xin[564]) );
  NANDN U2482 ( .A(start), .B(xreg[564]), .Z(n970) );
  NAND U2483 ( .A(x[564]), .B(start), .Z(n969) );
  NAND U2484 ( .A(n971), .B(n972), .Z(xin[563]) );
  NANDN U2485 ( .A(start), .B(xreg[563]), .Z(n972) );
  NAND U2486 ( .A(x[563]), .B(start), .Z(n971) );
  NAND U2487 ( .A(n973), .B(n974), .Z(xin[562]) );
  NANDN U2488 ( .A(start), .B(xreg[562]), .Z(n974) );
  NAND U2489 ( .A(x[562]), .B(start), .Z(n973) );
  NAND U2490 ( .A(n975), .B(n976), .Z(xin[561]) );
  NANDN U2491 ( .A(start), .B(xreg[561]), .Z(n976) );
  NAND U2492 ( .A(x[561]), .B(start), .Z(n975) );
  NAND U2493 ( .A(n977), .B(n978), .Z(xin[560]) );
  NANDN U2494 ( .A(start), .B(xreg[560]), .Z(n978) );
  NAND U2495 ( .A(x[560]), .B(start), .Z(n977) );
  NAND U2496 ( .A(n979), .B(n980), .Z(xin[55]) );
  NANDN U2497 ( .A(start), .B(xreg[55]), .Z(n980) );
  NAND U2498 ( .A(x[55]), .B(start), .Z(n979) );
  NAND U2499 ( .A(n981), .B(n982), .Z(xin[559]) );
  NANDN U2500 ( .A(start), .B(xreg[559]), .Z(n982) );
  NAND U2501 ( .A(x[559]), .B(start), .Z(n981) );
  NAND U2502 ( .A(n983), .B(n984), .Z(xin[558]) );
  NANDN U2503 ( .A(start), .B(xreg[558]), .Z(n984) );
  NAND U2504 ( .A(x[558]), .B(start), .Z(n983) );
  NAND U2505 ( .A(n985), .B(n986), .Z(xin[557]) );
  NANDN U2506 ( .A(start), .B(xreg[557]), .Z(n986) );
  NAND U2507 ( .A(x[557]), .B(start), .Z(n985) );
  NAND U2508 ( .A(n987), .B(n988), .Z(xin[556]) );
  NANDN U2509 ( .A(start), .B(xreg[556]), .Z(n988) );
  NAND U2510 ( .A(x[556]), .B(start), .Z(n987) );
  NAND U2511 ( .A(n989), .B(n990), .Z(xin[555]) );
  NANDN U2512 ( .A(start), .B(xreg[555]), .Z(n990) );
  NAND U2513 ( .A(x[555]), .B(start), .Z(n989) );
  NAND U2514 ( .A(n991), .B(n992), .Z(xin[554]) );
  NANDN U2515 ( .A(start), .B(xreg[554]), .Z(n992) );
  NAND U2516 ( .A(x[554]), .B(start), .Z(n991) );
  NAND U2517 ( .A(n993), .B(n994), .Z(xin[553]) );
  NANDN U2518 ( .A(start), .B(xreg[553]), .Z(n994) );
  NAND U2519 ( .A(x[553]), .B(start), .Z(n993) );
  NAND U2520 ( .A(n995), .B(n996), .Z(xin[552]) );
  NANDN U2521 ( .A(start), .B(xreg[552]), .Z(n996) );
  NAND U2522 ( .A(x[552]), .B(start), .Z(n995) );
  NAND U2523 ( .A(n997), .B(n998), .Z(xin[551]) );
  NANDN U2524 ( .A(start), .B(xreg[551]), .Z(n998) );
  NAND U2525 ( .A(x[551]), .B(start), .Z(n997) );
  NAND U2526 ( .A(n999), .B(n1000), .Z(xin[550]) );
  NANDN U2527 ( .A(start), .B(xreg[550]), .Z(n1000) );
  NAND U2528 ( .A(x[550]), .B(start), .Z(n999) );
  NAND U2529 ( .A(n1001), .B(n1002), .Z(xin[54]) );
  NANDN U2530 ( .A(start), .B(xreg[54]), .Z(n1002) );
  NAND U2531 ( .A(x[54]), .B(start), .Z(n1001) );
  NAND U2532 ( .A(n1003), .B(n1004), .Z(xin[549]) );
  NANDN U2533 ( .A(start), .B(xreg[549]), .Z(n1004) );
  NAND U2534 ( .A(x[549]), .B(start), .Z(n1003) );
  NAND U2535 ( .A(n1005), .B(n1006), .Z(xin[548]) );
  NANDN U2536 ( .A(start), .B(xreg[548]), .Z(n1006) );
  NAND U2537 ( .A(x[548]), .B(start), .Z(n1005) );
  NAND U2538 ( .A(n1007), .B(n1008), .Z(xin[547]) );
  NANDN U2539 ( .A(start), .B(xreg[547]), .Z(n1008) );
  NAND U2540 ( .A(x[547]), .B(start), .Z(n1007) );
  NAND U2541 ( .A(n1009), .B(n1010), .Z(xin[546]) );
  NANDN U2542 ( .A(start), .B(xreg[546]), .Z(n1010) );
  NAND U2543 ( .A(x[546]), .B(start), .Z(n1009) );
  NAND U2544 ( .A(n1011), .B(n1012), .Z(xin[545]) );
  NANDN U2545 ( .A(start), .B(xreg[545]), .Z(n1012) );
  NAND U2546 ( .A(x[545]), .B(start), .Z(n1011) );
  NAND U2547 ( .A(n1013), .B(n1014), .Z(xin[544]) );
  NANDN U2548 ( .A(start), .B(xreg[544]), .Z(n1014) );
  NAND U2549 ( .A(x[544]), .B(start), .Z(n1013) );
  NAND U2550 ( .A(n1015), .B(n1016), .Z(xin[543]) );
  NANDN U2551 ( .A(start), .B(xreg[543]), .Z(n1016) );
  NAND U2552 ( .A(x[543]), .B(start), .Z(n1015) );
  NAND U2553 ( .A(n1017), .B(n1018), .Z(xin[542]) );
  NANDN U2554 ( .A(start), .B(xreg[542]), .Z(n1018) );
  NAND U2555 ( .A(x[542]), .B(start), .Z(n1017) );
  NAND U2556 ( .A(n1019), .B(n1020), .Z(xin[541]) );
  NANDN U2557 ( .A(start), .B(xreg[541]), .Z(n1020) );
  NAND U2558 ( .A(x[541]), .B(start), .Z(n1019) );
  NAND U2559 ( .A(n1021), .B(n1022), .Z(xin[540]) );
  NANDN U2560 ( .A(start), .B(xreg[540]), .Z(n1022) );
  NAND U2561 ( .A(x[540]), .B(start), .Z(n1021) );
  NAND U2562 ( .A(n1023), .B(n1024), .Z(xin[53]) );
  NANDN U2563 ( .A(start), .B(xreg[53]), .Z(n1024) );
  NAND U2564 ( .A(x[53]), .B(start), .Z(n1023) );
  NAND U2565 ( .A(n1025), .B(n1026), .Z(xin[539]) );
  NANDN U2566 ( .A(start), .B(xreg[539]), .Z(n1026) );
  NAND U2567 ( .A(x[539]), .B(start), .Z(n1025) );
  NAND U2568 ( .A(n1027), .B(n1028), .Z(xin[538]) );
  NANDN U2569 ( .A(start), .B(xreg[538]), .Z(n1028) );
  NAND U2570 ( .A(x[538]), .B(start), .Z(n1027) );
  NAND U2571 ( .A(n1029), .B(n1030), .Z(xin[537]) );
  NANDN U2572 ( .A(start), .B(xreg[537]), .Z(n1030) );
  NAND U2573 ( .A(x[537]), .B(start), .Z(n1029) );
  NAND U2574 ( .A(n1031), .B(n1032), .Z(xin[536]) );
  NANDN U2575 ( .A(start), .B(xreg[536]), .Z(n1032) );
  NAND U2576 ( .A(x[536]), .B(start), .Z(n1031) );
  NAND U2577 ( .A(n1033), .B(n1034), .Z(xin[535]) );
  NANDN U2578 ( .A(start), .B(xreg[535]), .Z(n1034) );
  NAND U2579 ( .A(x[535]), .B(start), .Z(n1033) );
  NAND U2580 ( .A(n1035), .B(n1036), .Z(xin[534]) );
  NANDN U2581 ( .A(start), .B(xreg[534]), .Z(n1036) );
  NAND U2582 ( .A(x[534]), .B(start), .Z(n1035) );
  NAND U2583 ( .A(n1037), .B(n1038), .Z(xin[533]) );
  NANDN U2584 ( .A(start), .B(xreg[533]), .Z(n1038) );
  NAND U2585 ( .A(x[533]), .B(start), .Z(n1037) );
  NAND U2586 ( .A(n1039), .B(n1040), .Z(xin[532]) );
  NANDN U2587 ( .A(start), .B(xreg[532]), .Z(n1040) );
  NAND U2588 ( .A(x[532]), .B(start), .Z(n1039) );
  NAND U2589 ( .A(n1041), .B(n1042), .Z(xin[531]) );
  NANDN U2590 ( .A(start), .B(xreg[531]), .Z(n1042) );
  NAND U2591 ( .A(x[531]), .B(start), .Z(n1041) );
  NAND U2592 ( .A(n1043), .B(n1044), .Z(xin[530]) );
  NANDN U2593 ( .A(start), .B(xreg[530]), .Z(n1044) );
  NAND U2594 ( .A(x[530]), .B(start), .Z(n1043) );
  NAND U2595 ( .A(n1045), .B(n1046), .Z(xin[52]) );
  NANDN U2596 ( .A(start), .B(xreg[52]), .Z(n1046) );
  NAND U2597 ( .A(x[52]), .B(start), .Z(n1045) );
  NAND U2598 ( .A(n1047), .B(n1048), .Z(xin[529]) );
  NANDN U2599 ( .A(start), .B(xreg[529]), .Z(n1048) );
  NAND U2600 ( .A(x[529]), .B(start), .Z(n1047) );
  NAND U2601 ( .A(n1049), .B(n1050), .Z(xin[528]) );
  NANDN U2602 ( .A(start), .B(xreg[528]), .Z(n1050) );
  NAND U2603 ( .A(x[528]), .B(start), .Z(n1049) );
  NAND U2604 ( .A(n1051), .B(n1052), .Z(xin[527]) );
  NANDN U2605 ( .A(start), .B(xreg[527]), .Z(n1052) );
  NAND U2606 ( .A(x[527]), .B(start), .Z(n1051) );
  NAND U2607 ( .A(n1053), .B(n1054), .Z(xin[526]) );
  NANDN U2608 ( .A(start), .B(xreg[526]), .Z(n1054) );
  NAND U2609 ( .A(x[526]), .B(start), .Z(n1053) );
  NAND U2610 ( .A(n1055), .B(n1056), .Z(xin[525]) );
  NANDN U2611 ( .A(start), .B(xreg[525]), .Z(n1056) );
  NAND U2612 ( .A(x[525]), .B(start), .Z(n1055) );
  NAND U2613 ( .A(n1057), .B(n1058), .Z(xin[524]) );
  NANDN U2614 ( .A(start), .B(xreg[524]), .Z(n1058) );
  NAND U2615 ( .A(x[524]), .B(start), .Z(n1057) );
  NAND U2616 ( .A(n1059), .B(n1060), .Z(xin[523]) );
  NANDN U2617 ( .A(start), .B(xreg[523]), .Z(n1060) );
  NAND U2618 ( .A(x[523]), .B(start), .Z(n1059) );
  NAND U2619 ( .A(n1061), .B(n1062), .Z(xin[522]) );
  NANDN U2620 ( .A(start), .B(xreg[522]), .Z(n1062) );
  NAND U2621 ( .A(x[522]), .B(start), .Z(n1061) );
  NAND U2622 ( .A(n1063), .B(n1064), .Z(xin[521]) );
  NANDN U2623 ( .A(start), .B(xreg[521]), .Z(n1064) );
  NAND U2624 ( .A(x[521]), .B(start), .Z(n1063) );
  NAND U2625 ( .A(n1065), .B(n1066), .Z(xin[520]) );
  NANDN U2626 ( .A(start), .B(xreg[520]), .Z(n1066) );
  NAND U2627 ( .A(x[520]), .B(start), .Z(n1065) );
  NAND U2628 ( .A(n1067), .B(n1068), .Z(xin[51]) );
  NANDN U2629 ( .A(start), .B(xreg[51]), .Z(n1068) );
  NAND U2630 ( .A(x[51]), .B(start), .Z(n1067) );
  NAND U2631 ( .A(n1069), .B(n1070), .Z(xin[519]) );
  NANDN U2632 ( .A(start), .B(xreg[519]), .Z(n1070) );
  NAND U2633 ( .A(x[519]), .B(start), .Z(n1069) );
  NAND U2634 ( .A(n1071), .B(n1072), .Z(xin[518]) );
  NANDN U2635 ( .A(start), .B(xreg[518]), .Z(n1072) );
  NAND U2636 ( .A(x[518]), .B(start), .Z(n1071) );
  NAND U2637 ( .A(n1073), .B(n1074), .Z(xin[517]) );
  NANDN U2638 ( .A(start), .B(xreg[517]), .Z(n1074) );
  NAND U2639 ( .A(x[517]), .B(start), .Z(n1073) );
  NAND U2640 ( .A(n1075), .B(n1076), .Z(xin[516]) );
  NANDN U2641 ( .A(start), .B(xreg[516]), .Z(n1076) );
  NAND U2642 ( .A(x[516]), .B(start), .Z(n1075) );
  NAND U2643 ( .A(n1077), .B(n1078), .Z(xin[515]) );
  NANDN U2644 ( .A(start), .B(xreg[515]), .Z(n1078) );
  NAND U2645 ( .A(x[515]), .B(start), .Z(n1077) );
  NAND U2646 ( .A(n1079), .B(n1080), .Z(xin[514]) );
  NANDN U2647 ( .A(start), .B(xreg[514]), .Z(n1080) );
  NAND U2648 ( .A(x[514]), .B(start), .Z(n1079) );
  NAND U2649 ( .A(n1081), .B(n1082), .Z(xin[513]) );
  NANDN U2650 ( .A(start), .B(xreg[513]), .Z(n1082) );
  NAND U2651 ( .A(x[513]), .B(start), .Z(n1081) );
  NAND U2652 ( .A(n1083), .B(n1084), .Z(xin[512]) );
  NANDN U2653 ( .A(start), .B(xreg[512]), .Z(n1084) );
  NAND U2654 ( .A(x[512]), .B(start), .Z(n1083) );
  NAND U2655 ( .A(n1085), .B(n1086), .Z(xin[511]) );
  NANDN U2656 ( .A(start), .B(xreg[511]), .Z(n1086) );
  NAND U2657 ( .A(x[511]), .B(start), .Z(n1085) );
  NAND U2658 ( .A(n1087), .B(n1088), .Z(xin[510]) );
  NANDN U2659 ( .A(start), .B(xreg[510]), .Z(n1088) );
  NAND U2660 ( .A(x[510]), .B(start), .Z(n1087) );
  NAND U2661 ( .A(n1089), .B(n1090), .Z(xin[50]) );
  NANDN U2662 ( .A(start), .B(xreg[50]), .Z(n1090) );
  NAND U2663 ( .A(x[50]), .B(start), .Z(n1089) );
  NAND U2664 ( .A(n1091), .B(n1092), .Z(xin[509]) );
  NANDN U2665 ( .A(start), .B(xreg[509]), .Z(n1092) );
  NAND U2666 ( .A(x[509]), .B(start), .Z(n1091) );
  NAND U2667 ( .A(n1093), .B(n1094), .Z(xin[508]) );
  NANDN U2668 ( .A(start), .B(xreg[508]), .Z(n1094) );
  NAND U2669 ( .A(x[508]), .B(start), .Z(n1093) );
  NAND U2670 ( .A(n1095), .B(n1096), .Z(xin[507]) );
  NANDN U2671 ( .A(start), .B(xreg[507]), .Z(n1096) );
  NAND U2672 ( .A(x[507]), .B(start), .Z(n1095) );
  NAND U2673 ( .A(n1097), .B(n1098), .Z(xin[506]) );
  NANDN U2674 ( .A(start), .B(xreg[506]), .Z(n1098) );
  NAND U2675 ( .A(x[506]), .B(start), .Z(n1097) );
  NAND U2676 ( .A(n1099), .B(n1100), .Z(xin[505]) );
  NANDN U2677 ( .A(start), .B(xreg[505]), .Z(n1100) );
  NAND U2678 ( .A(x[505]), .B(start), .Z(n1099) );
  NAND U2679 ( .A(n1101), .B(n1102), .Z(xin[504]) );
  NANDN U2680 ( .A(start), .B(xreg[504]), .Z(n1102) );
  NAND U2681 ( .A(x[504]), .B(start), .Z(n1101) );
  NAND U2682 ( .A(n1103), .B(n1104), .Z(xin[503]) );
  NANDN U2683 ( .A(start), .B(xreg[503]), .Z(n1104) );
  NAND U2684 ( .A(x[503]), .B(start), .Z(n1103) );
  NAND U2685 ( .A(n1105), .B(n1106), .Z(xin[502]) );
  NANDN U2686 ( .A(start), .B(xreg[502]), .Z(n1106) );
  NAND U2687 ( .A(x[502]), .B(start), .Z(n1105) );
  NAND U2688 ( .A(n1107), .B(n1108), .Z(xin[501]) );
  NANDN U2689 ( .A(start), .B(xreg[501]), .Z(n1108) );
  NAND U2690 ( .A(x[501]), .B(start), .Z(n1107) );
  NAND U2691 ( .A(n1109), .B(n1110), .Z(xin[500]) );
  NANDN U2692 ( .A(start), .B(xreg[500]), .Z(n1110) );
  NAND U2693 ( .A(x[500]), .B(start), .Z(n1109) );
  NAND U2694 ( .A(n1111), .B(n1112), .Z(xin[4]) );
  NANDN U2695 ( .A(start), .B(xreg[4]), .Z(n1112) );
  NAND U2696 ( .A(x[4]), .B(start), .Z(n1111) );
  NAND U2697 ( .A(n1113), .B(n1114), .Z(xin[49]) );
  NANDN U2698 ( .A(start), .B(xreg[49]), .Z(n1114) );
  NAND U2699 ( .A(x[49]), .B(start), .Z(n1113) );
  NAND U2700 ( .A(n1115), .B(n1116), .Z(xin[499]) );
  NANDN U2701 ( .A(start), .B(xreg[499]), .Z(n1116) );
  NAND U2702 ( .A(x[499]), .B(start), .Z(n1115) );
  NAND U2703 ( .A(n1117), .B(n1118), .Z(xin[498]) );
  NANDN U2704 ( .A(start), .B(xreg[498]), .Z(n1118) );
  NAND U2705 ( .A(x[498]), .B(start), .Z(n1117) );
  NAND U2706 ( .A(n1119), .B(n1120), .Z(xin[497]) );
  NANDN U2707 ( .A(start), .B(xreg[497]), .Z(n1120) );
  NAND U2708 ( .A(x[497]), .B(start), .Z(n1119) );
  NAND U2709 ( .A(n1121), .B(n1122), .Z(xin[496]) );
  NANDN U2710 ( .A(start), .B(xreg[496]), .Z(n1122) );
  NAND U2711 ( .A(x[496]), .B(start), .Z(n1121) );
  NAND U2712 ( .A(n1123), .B(n1124), .Z(xin[495]) );
  NANDN U2713 ( .A(start), .B(xreg[495]), .Z(n1124) );
  NAND U2714 ( .A(x[495]), .B(start), .Z(n1123) );
  NAND U2715 ( .A(n1125), .B(n1126), .Z(xin[494]) );
  NANDN U2716 ( .A(start), .B(xreg[494]), .Z(n1126) );
  NAND U2717 ( .A(x[494]), .B(start), .Z(n1125) );
  NAND U2718 ( .A(n1127), .B(n1128), .Z(xin[493]) );
  NANDN U2719 ( .A(start), .B(xreg[493]), .Z(n1128) );
  NAND U2720 ( .A(x[493]), .B(start), .Z(n1127) );
  NAND U2721 ( .A(n1129), .B(n1130), .Z(xin[492]) );
  NANDN U2722 ( .A(start), .B(xreg[492]), .Z(n1130) );
  NAND U2723 ( .A(x[492]), .B(start), .Z(n1129) );
  NAND U2724 ( .A(n1131), .B(n1132), .Z(xin[491]) );
  NANDN U2725 ( .A(start), .B(xreg[491]), .Z(n1132) );
  NAND U2726 ( .A(x[491]), .B(start), .Z(n1131) );
  NAND U2727 ( .A(n1133), .B(n1134), .Z(xin[490]) );
  NANDN U2728 ( .A(start), .B(xreg[490]), .Z(n1134) );
  NAND U2729 ( .A(x[490]), .B(start), .Z(n1133) );
  NAND U2730 ( .A(n1135), .B(n1136), .Z(xin[48]) );
  NANDN U2731 ( .A(start), .B(xreg[48]), .Z(n1136) );
  NAND U2732 ( .A(x[48]), .B(start), .Z(n1135) );
  NAND U2733 ( .A(n1137), .B(n1138), .Z(xin[489]) );
  NANDN U2734 ( .A(start), .B(xreg[489]), .Z(n1138) );
  NAND U2735 ( .A(x[489]), .B(start), .Z(n1137) );
  NAND U2736 ( .A(n1139), .B(n1140), .Z(xin[488]) );
  NANDN U2737 ( .A(start), .B(xreg[488]), .Z(n1140) );
  NAND U2738 ( .A(x[488]), .B(start), .Z(n1139) );
  NAND U2739 ( .A(n1141), .B(n1142), .Z(xin[487]) );
  NANDN U2740 ( .A(start), .B(xreg[487]), .Z(n1142) );
  NAND U2741 ( .A(x[487]), .B(start), .Z(n1141) );
  NAND U2742 ( .A(n1143), .B(n1144), .Z(xin[486]) );
  NANDN U2743 ( .A(start), .B(xreg[486]), .Z(n1144) );
  NAND U2744 ( .A(x[486]), .B(start), .Z(n1143) );
  NAND U2745 ( .A(n1145), .B(n1146), .Z(xin[485]) );
  NANDN U2746 ( .A(start), .B(xreg[485]), .Z(n1146) );
  NAND U2747 ( .A(x[485]), .B(start), .Z(n1145) );
  NAND U2748 ( .A(n1147), .B(n1148), .Z(xin[484]) );
  NANDN U2749 ( .A(start), .B(xreg[484]), .Z(n1148) );
  NAND U2750 ( .A(x[484]), .B(start), .Z(n1147) );
  NAND U2751 ( .A(n1149), .B(n1150), .Z(xin[483]) );
  NANDN U2752 ( .A(start), .B(xreg[483]), .Z(n1150) );
  NAND U2753 ( .A(x[483]), .B(start), .Z(n1149) );
  NAND U2754 ( .A(n1151), .B(n1152), .Z(xin[482]) );
  NANDN U2755 ( .A(start), .B(xreg[482]), .Z(n1152) );
  NAND U2756 ( .A(x[482]), .B(start), .Z(n1151) );
  NAND U2757 ( .A(n1153), .B(n1154), .Z(xin[481]) );
  NANDN U2758 ( .A(start), .B(xreg[481]), .Z(n1154) );
  NAND U2759 ( .A(x[481]), .B(start), .Z(n1153) );
  NAND U2760 ( .A(n1155), .B(n1156), .Z(xin[480]) );
  NANDN U2761 ( .A(start), .B(xreg[480]), .Z(n1156) );
  NAND U2762 ( .A(x[480]), .B(start), .Z(n1155) );
  NAND U2763 ( .A(n1157), .B(n1158), .Z(xin[47]) );
  NANDN U2764 ( .A(start), .B(xreg[47]), .Z(n1158) );
  NAND U2765 ( .A(x[47]), .B(start), .Z(n1157) );
  NAND U2766 ( .A(n1159), .B(n1160), .Z(xin[479]) );
  NANDN U2767 ( .A(start), .B(xreg[479]), .Z(n1160) );
  NAND U2768 ( .A(x[479]), .B(start), .Z(n1159) );
  NAND U2769 ( .A(n1161), .B(n1162), .Z(xin[478]) );
  NANDN U2770 ( .A(start), .B(xreg[478]), .Z(n1162) );
  NAND U2771 ( .A(x[478]), .B(start), .Z(n1161) );
  NAND U2772 ( .A(n1163), .B(n1164), .Z(xin[477]) );
  NANDN U2773 ( .A(start), .B(xreg[477]), .Z(n1164) );
  NAND U2774 ( .A(x[477]), .B(start), .Z(n1163) );
  NAND U2775 ( .A(n1165), .B(n1166), .Z(xin[476]) );
  NANDN U2776 ( .A(start), .B(xreg[476]), .Z(n1166) );
  NAND U2777 ( .A(x[476]), .B(start), .Z(n1165) );
  NAND U2778 ( .A(n1167), .B(n1168), .Z(xin[475]) );
  NANDN U2779 ( .A(start), .B(xreg[475]), .Z(n1168) );
  NAND U2780 ( .A(x[475]), .B(start), .Z(n1167) );
  NAND U2781 ( .A(n1169), .B(n1170), .Z(xin[474]) );
  NANDN U2782 ( .A(start), .B(xreg[474]), .Z(n1170) );
  NAND U2783 ( .A(x[474]), .B(start), .Z(n1169) );
  NAND U2784 ( .A(n1171), .B(n1172), .Z(xin[473]) );
  NANDN U2785 ( .A(start), .B(xreg[473]), .Z(n1172) );
  NAND U2786 ( .A(x[473]), .B(start), .Z(n1171) );
  NAND U2787 ( .A(n1173), .B(n1174), .Z(xin[472]) );
  NANDN U2788 ( .A(start), .B(xreg[472]), .Z(n1174) );
  NAND U2789 ( .A(x[472]), .B(start), .Z(n1173) );
  NAND U2790 ( .A(n1175), .B(n1176), .Z(xin[471]) );
  NANDN U2791 ( .A(start), .B(xreg[471]), .Z(n1176) );
  NAND U2792 ( .A(x[471]), .B(start), .Z(n1175) );
  NAND U2793 ( .A(n1177), .B(n1178), .Z(xin[470]) );
  NANDN U2794 ( .A(start), .B(xreg[470]), .Z(n1178) );
  NAND U2795 ( .A(x[470]), .B(start), .Z(n1177) );
  NAND U2796 ( .A(n1179), .B(n1180), .Z(xin[46]) );
  NANDN U2797 ( .A(start), .B(xreg[46]), .Z(n1180) );
  NAND U2798 ( .A(x[46]), .B(start), .Z(n1179) );
  NAND U2799 ( .A(n1181), .B(n1182), .Z(xin[469]) );
  NANDN U2800 ( .A(start), .B(xreg[469]), .Z(n1182) );
  NAND U2801 ( .A(x[469]), .B(start), .Z(n1181) );
  NAND U2802 ( .A(n1183), .B(n1184), .Z(xin[468]) );
  NANDN U2803 ( .A(start), .B(xreg[468]), .Z(n1184) );
  NAND U2804 ( .A(x[468]), .B(start), .Z(n1183) );
  NAND U2805 ( .A(n1185), .B(n1186), .Z(xin[467]) );
  NANDN U2806 ( .A(start), .B(xreg[467]), .Z(n1186) );
  NAND U2807 ( .A(x[467]), .B(start), .Z(n1185) );
  NAND U2808 ( .A(n1187), .B(n1188), .Z(xin[466]) );
  NANDN U2809 ( .A(start), .B(xreg[466]), .Z(n1188) );
  NAND U2810 ( .A(x[466]), .B(start), .Z(n1187) );
  NAND U2811 ( .A(n1189), .B(n1190), .Z(xin[465]) );
  NANDN U2812 ( .A(start), .B(xreg[465]), .Z(n1190) );
  NAND U2813 ( .A(x[465]), .B(start), .Z(n1189) );
  NAND U2814 ( .A(n1191), .B(n1192), .Z(xin[464]) );
  NANDN U2815 ( .A(start), .B(xreg[464]), .Z(n1192) );
  NAND U2816 ( .A(x[464]), .B(start), .Z(n1191) );
  NAND U2817 ( .A(n1193), .B(n1194), .Z(xin[463]) );
  NANDN U2818 ( .A(start), .B(xreg[463]), .Z(n1194) );
  NAND U2819 ( .A(x[463]), .B(start), .Z(n1193) );
  NAND U2820 ( .A(n1195), .B(n1196), .Z(xin[462]) );
  NANDN U2821 ( .A(start), .B(xreg[462]), .Z(n1196) );
  NAND U2822 ( .A(x[462]), .B(start), .Z(n1195) );
  NAND U2823 ( .A(n1197), .B(n1198), .Z(xin[461]) );
  NANDN U2824 ( .A(start), .B(xreg[461]), .Z(n1198) );
  NAND U2825 ( .A(x[461]), .B(start), .Z(n1197) );
  NAND U2826 ( .A(n1199), .B(n1200), .Z(xin[460]) );
  NANDN U2827 ( .A(start), .B(xreg[460]), .Z(n1200) );
  NAND U2828 ( .A(x[460]), .B(start), .Z(n1199) );
  NAND U2829 ( .A(n1201), .B(n1202), .Z(xin[45]) );
  NANDN U2830 ( .A(start), .B(xreg[45]), .Z(n1202) );
  NAND U2831 ( .A(x[45]), .B(start), .Z(n1201) );
  NAND U2832 ( .A(n1203), .B(n1204), .Z(xin[459]) );
  NANDN U2833 ( .A(start), .B(xreg[459]), .Z(n1204) );
  NAND U2834 ( .A(x[459]), .B(start), .Z(n1203) );
  NAND U2835 ( .A(n1205), .B(n1206), .Z(xin[458]) );
  NANDN U2836 ( .A(start), .B(xreg[458]), .Z(n1206) );
  NAND U2837 ( .A(x[458]), .B(start), .Z(n1205) );
  NAND U2838 ( .A(n1207), .B(n1208), .Z(xin[457]) );
  NANDN U2839 ( .A(start), .B(xreg[457]), .Z(n1208) );
  NAND U2840 ( .A(x[457]), .B(start), .Z(n1207) );
  NAND U2841 ( .A(n1209), .B(n1210), .Z(xin[456]) );
  NANDN U2842 ( .A(start), .B(xreg[456]), .Z(n1210) );
  NAND U2843 ( .A(x[456]), .B(start), .Z(n1209) );
  NAND U2844 ( .A(n1211), .B(n1212), .Z(xin[455]) );
  NANDN U2845 ( .A(start), .B(xreg[455]), .Z(n1212) );
  NAND U2846 ( .A(x[455]), .B(start), .Z(n1211) );
  NAND U2847 ( .A(n1213), .B(n1214), .Z(xin[454]) );
  NANDN U2848 ( .A(start), .B(xreg[454]), .Z(n1214) );
  NAND U2849 ( .A(x[454]), .B(start), .Z(n1213) );
  NAND U2850 ( .A(n1215), .B(n1216), .Z(xin[453]) );
  NANDN U2851 ( .A(start), .B(xreg[453]), .Z(n1216) );
  NAND U2852 ( .A(x[453]), .B(start), .Z(n1215) );
  NAND U2853 ( .A(n1217), .B(n1218), .Z(xin[452]) );
  NANDN U2854 ( .A(start), .B(xreg[452]), .Z(n1218) );
  NAND U2855 ( .A(x[452]), .B(start), .Z(n1217) );
  NAND U2856 ( .A(n1219), .B(n1220), .Z(xin[451]) );
  NANDN U2857 ( .A(start), .B(xreg[451]), .Z(n1220) );
  NAND U2858 ( .A(x[451]), .B(start), .Z(n1219) );
  NAND U2859 ( .A(n1221), .B(n1222), .Z(xin[450]) );
  NANDN U2860 ( .A(start), .B(xreg[450]), .Z(n1222) );
  NAND U2861 ( .A(x[450]), .B(start), .Z(n1221) );
  NAND U2862 ( .A(n1223), .B(n1224), .Z(xin[44]) );
  NANDN U2863 ( .A(start), .B(xreg[44]), .Z(n1224) );
  NAND U2864 ( .A(x[44]), .B(start), .Z(n1223) );
  NAND U2865 ( .A(n1225), .B(n1226), .Z(xin[449]) );
  NANDN U2866 ( .A(start), .B(xreg[449]), .Z(n1226) );
  NAND U2867 ( .A(x[449]), .B(start), .Z(n1225) );
  NAND U2868 ( .A(n1227), .B(n1228), .Z(xin[448]) );
  NANDN U2869 ( .A(start), .B(xreg[448]), .Z(n1228) );
  NAND U2870 ( .A(x[448]), .B(start), .Z(n1227) );
  NAND U2871 ( .A(n1229), .B(n1230), .Z(xin[447]) );
  NANDN U2872 ( .A(start), .B(xreg[447]), .Z(n1230) );
  NAND U2873 ( .A(x[447]), .B(start), .Z(n1229) );
  NAND U2874 ( .A(n1231), .B(n1232), .Z(xin[446]) );
  NANDN U2875 ( .A(start), .B(xreg[446]), .Z(n1232) );
  NAND U2876 ( .A(x[446]), .B(start), .Z(n1231) );
  NAND U2877 ( .A(n1233), .B(n1234), .Z(xin[445]) );
  NANDN U2878 ( .A(start), .B(xreg[445]), .Z(n1234) );
  NAND U2879 ( .A(x[445]), .B(start), .Z(n1233) );
  NAND U2880 ( .A(n1235), .B(n1236), .Z(xin[444]) );
  NANDN U2881 ( .A(start), .B(xreg[444]), .Z(n1236) );
  NAND U2882 ( .A(x[444]), .B(start), .Z(n1235) );
  NAND U2883 ( .A(n1237), .B(n1238), .Z(xin[443]) );
  NANDN U2884 ( .A(start), .B(xreg[443]), .Z(n1238) );
  NAND U2885 ( .A(x[443]), .B(start), .Z(n1237) );
  NAND U2886 ( .A(n1239), .B(n1240), .Z(xin[442]) );
  NANDN U2887 ( .A(start), .B(xreg[442]), .Z(n1240) );
  NAND U2888 ( .A(x[442]), .B(start), .Z(n1239) );
  NAND U2889 ( .A(n1241), .B(n1242), .Z(xin[441]) );
  NANDN U2890 ( .A(start), .B(xreg[441]), .Z(n1242) );
  NAND U2891 ( .A(x[441]), .B(start), .Z(n1241) );
  NAND U2892 ( .A(n1243), .B(n1244), .Z(xin[440]) );
  NANDN U2893 ( .A(start), .B(xreg[440]), .Z(n1244) );
  NAND U2894 ( .A(x[440]), .B(start), .Z(n1243) );
  NAND U2895 ( .A(n1245), .B(n1246), .Z(xin[43]) );
  NANDN U2896 ( .A(start), .B(xreg[43]), .Z(n1246) );
  NAND U2897 ( .A(x[43]), .B(start), .Z(n1245) );
  NAND U2898 ( .A(n1247), .B(n1248), .Z(xin[439]) );
  NANDN U2899 ( .A(start), .B(xreg[439]), .Z(n1248) );
  NAND U2900 ( .A(x[439]), .B(start), .Z(n1247) );
  NAND U2901 ( .A(n1249), .B(n1250), .Z(xin[438]) );
  NANDN U2902 ( .A(start), .B(xreg[438]), .Z(n1250) );
  NAND U2903 ( .A(x[438]), .B(start), .Z(n1249) );
  NAND U2904 ( .A(n1251), .B(n1252), .Z(xin[437]) );
  NANDN U2905 ( .A(start), .B(xreg[437]), .Z(n1252) );
  NAND U2906 ( .A(x[437]), .B(start), .Z(n1251) );
  NAND U2907 ( .A(n1253), .B(n1254), .Z(xin[436]) );
  NANDN U2908 ( .A(start), .B(xreg[436]), .Z(n1254) );
  NAND U2909 ( .A(x[436]), .B(start), .Z(n1253) );
  NAND U2910 ( .A(n1255), .B(n1256), .Z(xin[435]) );
  NANDN U2911 ( .A(start), .B(xreg[435]), .Z(n1256) );
  NAND U2912 ( .A(x[435]), .B(start), .Z(n1255) );
  NAND U2913 ( .A(n1257), .B(n1258), .Z(xin[434]) );
  NANDN U2914 ( .A(start), .B(xreg[434]), .Z(n1258) );
  NAND U2915 ( .A(x[434]), .B(start), .Z(n1257) );
  NAND U2916 ( .A(n1259), .B(n1260), .Z(xin[433]) );
  NANDN U2917 ( .A(start), .B(xreg[433]), .Z(n1260) );
  NAND U2918 ( .A(x[433]), .B(start), .Z(n1259) );
  NAND U2919 ( .A(n1261), .B(n1262), .Z(xin[432]) );
  NANDN U2920 ( .A(start), .B(xreg[432]), .Z(n1262) );
  NAND U2921 ( .A(x[432]), .B(start), .Z(n1261) );
  NAND U2922 ( .A(n1263), .B(n1264), .Z(xin[431]) );
  NANDN U2923 ( .A(start), .B(xreg[431]), .Z(n1264) );
  NAND U2924 ( .A(x[431]), .B(start), .Z(n1263) );
  NAND U2925 ( .A(n1265), .B(n1266), .Z(xin[430]) );
  NANDN U2926 ( .A(start), .B(xreg[430]), .Z(n1266) );
  NAND U2927 ( .A(x[430]), .B(start), .Z(n1265) );
  NAND U2928 ( .A(n1267), .B(n1268), .Z(xin[42]) );
  NANDN U2929 ( .A(start), .B(xreg[42]), .Z(n1268) );
  NAND U2930 ( .A(x[42]), .B(start), .Z(n1267) );
  NAND U2931 ( .A(n1269), .B(n1270), .Z(xin[429]) );
  NANDN U2932 ( .A(start), .B(xreg[429]), .Z(n1270) );
  NAND U2933 ( .A(x[429]), .B(start), .Z(n1269) );
  NAND U2934 ( .A(n1271), .B(n1272), .Z(xin[428]) );
  NANDN U2935 ( .A(start), .B(xreg[428]), .Z(n1272) );
  NAND U2936 ( .A(x[428]), .B(start), .Z(n1271) );
  NAND U2937 ( .A(n1273), .B(n1274), .Z(xin[427]) );
  NANDN U2938 ( .A(start), .B(xreg[427]), .Z(n1274) );
  NAND U2939 ( .A(x[427]), .B(start), .Z(n1273) );
  NAND U2940 ( .A(n1275), .B(n1276), .Z(xin[426]) );
  NANDN U2941 ( .A(start), .B(xreg[426]), .Z(n1276) );
  NAND U2942 ( .A(x[426]), .B(start), .Z(n1275) );
  NAND U2943 ( .A(n1277), .B(n1278), .Z(xin[425]) );
  NANDN U2944 ( .A(start), .B(xreg[425]), .Z(n1278) );
  NAND U2945 ( .A(x[425]), .B(start), .Z(n1277) );
  NAND U2946 ( .A(n1279), .B(n1280), .Z(xin[424]) );
  NANDN U2947 ( .A(start), .B(xreg[424]), .Z(n1280) );
  NAND U2948 ( .A(x[424]), .B(start), .Z(n1279) );
  NAND U2949 ( .A(n1281), .B(n1282), .Z(xin[423]) );
  NANDN U2950 ( .A(start), .B(xreg[423]), .Z(n1282) );
  NAND U2951 ( .A(x[423]), .B(start), .Z(n1281) );
  NAND U2952 ( .A(n1283), .B(n1284), .Z(xin[422]) );
  NANDN U2953 ( .A(start), .B(xreg[422]), .Z(n1284) );
  NAND U2954 ( .A(x[422]), .B(start), .Z(n1283) );
  NAND U2955 ( .A(n1285), .B(n1286), .Z(xin[421]) );
  NANDN U2956 ( .A(start), .B(xreg[421]), .Z(n1286) );
  NAND U2957 ( .A(x[421]), .B(start), .Z(n1285) );
  NAND U2958 ( .A(n1287), .B(n1288), .Z(xin[420]) );
  NANDN U2959 ( .A(start), .B(xreg[420]), .Z(n1288) );
  NAND U2960 ( .A(x[420]), .B(start), .Z(n1287) );
  NAND U2961 ( .A(n1289), .B(n1290), .Z(xin[41]) );
  NANDN U2962 ( .A(start), .B(xreg[41]), .Z(n1290) );
  NAND U2963 ( .A(x[41]), .B(start), .Z(n1289) );
  NAND U2964 ( .A(n1291), .B(n1292), .Z(xin[419]) );
  NANDN U2965 ( .A(start), .B(xreg[419]), .Z(n1292) );
  NAND U2966 ( .A(x[419]), .B(start), .Z(n1291) );
  NAND U2967 ( .A(n1293), .B(n1294), .Z(xin[418]) );
  NANDN U2968 ( .A(start), .B(xreg[418]), .Z(n1294) );
  NAND U2969 ( .A(x[418]), .B(start), .Z(n1293) );
  NAND U2970 ( .A(n1295), .B(n1296), .Z(xin[417]) );
  NANDN U2971 ( .A(start), .B(xreg[417]), .Z(n1296) );
  NAND U2972 ( .A(x[417]), .B(start), .Z(n1295) );
  NAND U2973 ( .A(n1297), .B(n1298), .Z(xin[416]) );
  NANDN U2974 ( .A(start), .B(xreg[416]), .Z(n1298) );
  NAND U2975 ( .A(x[416]), .B(start), .Z(n1297) );
  NAND U2976 ( .A(n1299), .B(n1300), .Z(xin[415]) );
  NANDN U2977 ( .A(start), .B(xreg[415]), .Z(n1300) );
  NAND U2978 ( .A(x[415]), .B(start), .Z(n1299) );
  NAND U2979 ( .A(n1301), .B(n1302), .Z(xin[414]) );
  NANDN U2980 ( .A(start), .B(xreg[414]), .Z(n1302) );
  NAND U2981 ( .A(x[414]), .B(start), .Z(n1301) );
  NAND U2982 ( .A(n1303), .B(n1304), .Z(xin[413]) );
  NANDN U2983 ( .A(start), .B(xreg[413]), .Z(n1304) );
  NAND U2984 ( .A(x[413]), .B(start), .Z(n1303) );
  NAND U2985 ( .A(n1305), .B(n1306), .Z(xin[412]) );
  NANDN U2986 ( .A(start), .B(xreg[412]), .Z(n1306) );
  NAND U2987 ( .A(x[412]), .B(start), .Z(n1305) );
  NAND U2988 ( .A(n1307), .B(n1308), .Z(xin[411]) );
  NANDN U2989 ( .A(start), .B(xreg[411]), .Z(n1308) );
  NAND U2990 ( .A(x[411]), .B(start), .Z(n1307) );
  NAND U2991 ( .A(n1309), .B(n1310), .Z(xin[410]) );
  NANDN U2992 ( .A(start), .B(xreg[410]), .Z(n1310) );
  NAND U2993 ( .A(x[410]), .B(start), .Z(n1309) );
  NAND U2994 ( .A(n1311), .B(n1312), .Z(xin[40]) );
  NANDN U2995 ( .A(start), .B(xreg[40]), .Z(n1312) );
  NAND U2996 ( .A(x[40]), .B(start), .Z(n1311) );
  NAND U2997 ( .A(n1313), .B(n1314), .Z(xin[409]) );
  NANDN U2998 ( .A(start), .B(xreg[409]), .Z(n1314) );
  NAND U2999 ( .A(x[409]), .B(start), .Z(n1313) );
  NAND U3000 ( .A(n1315), .B(n1316), .Z(xin[408]) );
  NANDN U3001 ( .A(start), .B(xreg[408]), .Z(n1316) );
  NAND U3002 ( .A(x[408]), .B(start), .Z(n1315) );
  NAND U3003 ( .A(n1317), .B(n1318), .Z(xin[407]) );
  NANDN U3004 ( .A(start), .B(xreg[407]), .Z(n1318) );
  NAND U3005 ( .A(x[407]), .B(start), .Z(n1317) );
  NAND U3006 ( .A(n1319), .B(n1320), .Z(xin[406]) );
  NANDN U3007 ( .A(start), .B(xreg[406]), .Z(n1320) );
  NAND U3008 ( .A(x[406]), .B(start), .Z(n1319) );
  NAND U3009 ( .A(n1321), .B(n1322), .Z(xin[405]) );
  NANDN U3010 ( .A(start), .B(xreg[405]), .Z(n1322) );
  NAND U3011 ( .A(x[405]), .B(start), .Z(n1321) );
  NAND U3012 ( .A(n1323), .B(n1324), .Z(xin[404]) );
  NANDN U3013 ( .A(start), .B(xreg[404]), .Z(n1324) );
  NAND U3014 ( .A(x[404]), .B(start), .Z(n1323) );
  NAND U3015 ( .A(n1325), .B(n1326), .Z(xin[403]) );
  NANDN U3016 ( .A(start), .B(xreg[403]), .Z(n1326) );
  NAND U3017 ( .A(x[403]), .B(start), .Z(n1325) );
  NAND U3018 ( .A(n1327), .B(n1328), .Z(xin[402]) );
  NANDN U3019 ( .A(start), .B(xreg[402]), .Z(n1328) );
  NAND U3020 ( .A(x[402]), .B(start), .Z(n1327) );
  NAND U3021 ( .A(n1329), .B(n1330), .Z(xin[401]) );
  NANDN U3022 ( .A(start), .B(xreg[401]), .Z(n1330) );
  NAND U3023 ( .A(x[401]), .B(start), .Z(n1329) );
  NAND U3024 ( .A(n1331), .B(n1332), .Z(xin[400]) );
  NANDN U3025 ( .A(start), .B(xreg[400]), .Z(n1332) );
  NAND U3026 ( .A(x[400]), .B(start), .Z(n1331) );
  NAND U3027 ( .A(n1333), .B(n1334), .Z(xin[3]) );
  NANDN U3028 ( .A(start), .B(xreg[3]), .Z(n1334) );
  NAND U3029 ( .A(x[3]), .B(start), .Z(n1333) );
  NAND U3030 ( .A(n1335), .B(n1336), .Z(xin[39]) );
  NANDN U3031 ( .A(start), .B(xreg[39]), .Z(n1336) );
  NAND U3032 ( .A(x[39]), .B(start), .Z(n1335) );
  NAND U3033 ( .A(n1337), .B(n1338), .Z(xin[399]) );
  NANDN U3034 ( .A(start), .B(xreg[399]), .Z(n1338) );
  NAND U3035 ( .A(x[399]), .B(start), .Z(n1337) );
  NAND U3036 ( .A(n1339), .B(n1340), .Z(xin[398]) );
  NANDN U3037 ( .A(start), .B(xreg[398]), .Z(n1340) );
  NAND U3038 ( .A(x[398]), .B(start), .Z(n1339) );
  NAND U3039 ( .A(n1341), .B(n1342), .Z(xin[397]) );
  NANDN U3040 ( .A(start), .B(xreg[397]), .Z(n1342) );
  NAND U3041 ( .A(x[397]), .B(start), .Z(n1341) );
  NAND U3042 ( .A(n1343), .B(n1344), .Z(xin[396]) );
  NANDN U3043 ( .A(start), .B(xreg[396]), .Z(n1344) );
  NAND U3044 ( .A(x[396]), .B(start), .Z(n1343) );
  NAND U3045 ( .A(n1345), .B(n1346), .Z(xin[395]) );
  NANDN U3046 ( .A(start), .B(xreg[395]), .Z(n1346) );
  NAND U3047 ( .A(x[395]), .B(start), .Z(n1345) );
  NAND U3048 ( .A(n1347), .B(n1348), .Z(xin[394]) );
  NANDN U3049 ( .A(start), .B(xreg[394]), .Z(n1348) );
  NAND U3050 ( .A(x[394]), .B(start), .Z(n1347) );
  NAND U3051 ( .A(n1349), .B(n1350), .Z(xin[393]) );
  NANDN U3052 ( .A(start), .B(xreg[393]), .Z(n1350) );
  NAND U3053 ( .A(x[393]), .B(start), .Z(n1349) );
  NAND U3054 ( .A(n1351), .B(n1352), .Z(xin[392]) );
  NANDN U3055 ( .A(start), .B(xreg[392]), .Z(n1352) );
  NAND U3056 ( .A(x[392]), .B(start), .Z(n1351) );
  NAND U3057 ( .A(n1353), .B(n1354), .Z(xin[391]) );
  NANDN U3058 ( .A(start), .B(xreg[391]), .Z(n1354) );
  NAND U3059 ( .A(x[391]), .B(start), .Z(n1353) );
  NAND U3060 ( .A(n1355), .B(n1356), .Z(xin[390]) );
  NANDN U3061 ( .A(start), .B(xreg[390]), .Z(n1356) );
  NAND U3062 ( .A(x[390]), .B(start), .Z(n1355) );
  NAND U3063 ( .A(n1357), .B(n1358), .Z(xin[38]) );
  NANDN U3064 ( .A(start), .B(xreg[38]), .Z(n1358) );
  NAND U3065 ( .A(x[38]), .B(start), .Z(n1357) );
  NAND U3066 ( .A(n1359), .B(n1360), .Z(xin[389]) );
  NANDN U3067 ( .A(start), .B(xreg[389]), .Z(n1360) );
  NAND U3068 ( .A(x[389]), .B(start), .Z(n1359) );
  NAND U3069 ( .A(n1361), .B(n1362), .Z(xin[388]) );
  NANDN U3070 ( .A(start), .B(xreg[388]), .Z(n1362) );
  NAND U3071 ( .A(x[388]), .B(start), .Z(n1361) );
  NAND U3072 ( .A(n1363), .B(n1364), .Z(xin[387]) );
  NANDN U3073 ( .A(start), .B(xreg[387]), .Z(n1364) );
  NAND U3074 ( .A(x[387]), .B(start), .Z(n1363) );
  NAND U3075 ( .A(n1365), .B(n1366), .Z(xin[386]) );
  NANDN U3076 ( .A(start), .B(xreg[386]), .Z(n1366) );
  NAND U3077 ( .A(x[386]), .B(start), .Z(n1365) );
  NAND U3078 ( .A(n1367), .B(n1368), .Z(xin[385]) );
  NANDN U3079 ( .A(start), .B(xreg[385]), .Z(n1368) );
  NAND U3080 ( .A(x[385]), .B(start), .Z(n1367) );
  NAND U3081 ( .A(n1369), .B(n1370), .Z(xin[384]) );
  NANDN U3082 ( .A(start), .B(xreg[384]), .Z(n1370) );
  NAND U3083 ( .A(x[384]), .B(start), .Z(n1369) );
  NAND U3084 ( .A(n1371), .B(n1372), .Z(xin[383]) );
  NANDN U3085 ( .A(start), .B(xreg[383]), .Z(n1372) );
  NAND U3086 ( .A(x[383]), .B(start), .Z(n1371) );
  NAND U3087 ( .A(n1373), .B(n1374), .Z(xin[382]) );
  NANDN U3088 ( .A(start), .B(xreg[382]), .Z(n1374) );
  NAND U3089 ( .A(x[382]), .B(start), .Z(n1373) );
  NAND U3090 ( .A(n1375), .B(n1376), .Z(xin[381]) );
  NANDN U3091 ( .A(start), .B(xreg[381]), .Z(n1376) );
  NAND U3092 ( .A(x[381]), .B(start), .Z(n1375) );
  NAND U3093 ( .A(n1377), .B(n1378), .Z(xin[380]) );
  NANDN U3094 ( .A(start), .B(xreg[380]), .Z(n1378) );
  NAND U3095 ( .A(x[380]), .B(start), .Z(n1377) );
  NAND U3096 ( .A(n1379), .B(n1380), .Z(xin[37]) );
  NANDN U3097 ( .A(start), .B(xreg[37]), .Z(n1380) );
  NAND U3098 ( .A(x[37]), .B(start), .Z(n1379) );
  NAND U3099 ( .A(n1381), .B(n1382), .Z(xin[379]) );
  NANDN U3100 ( .A(start), .B(xreg[379]), .Z(n1382) );
  NAND U3101 ( .A(x[379]), .B(start), .Z(n1381) );
  NAND U3102 ( .A(n1383), .B(n1384), .Z(xin[378]) );
  NANDN U3103 ( .A(start), .B(xreg[378]), .Z(n1384) );
  NAND U3104 ( .A(x[378]), .B(start), .Z(n1383) );
  NAND U3105 ( .A(n1385), .B(n1386), .Z(xin[377]) );
  NANDN U3106 ( .A(start), .B(xreg[377]), .Z(n1386) );
  NAND U3107 ( .A(x[377]), .B(start), .Z(n1385) );
  NAND U3108 ( .A(n1387), .B(n1388), .Z(xin[376]) );
  NANDN U3109 ( .A(start), .B(xreg[376]), .Z(n1388) );
  NAND U3110 ( .A(x[376]), .B(start), .Z(n1387) );
  NAND U3111 ( .A(n1389), .B(n1390), .Z(xin[375]) );
  NANDN U3112 ( .A(start), .B(xreg[375]), .Z(n1390) );
  NAND U3113 ( .A(x[375]), .B(start), .Z(n1389) );
  NAND U3114 ( .A(n1391), .B(n1392), .Z(xin[374]) );
  NANDN U3115 ( .A(start), .B(xreg[374]), .Z(n1392) );
  NAND U3116 ( .A(x[374]), .B(start), .Z(n1391) );
  NAND U3117 ( .A(n1393), .B(n1394), .Z(xin[373]) );
  NANDN U3118 ( .A(start), .B(xreg[373]), .Z(n1394) );
  NAND U3119 ( .A(x[373]), .B(start), .Z(n1393) );
  NAND U3120 ( .A(n1395), .B(n1396), .Z(xin[372]) );
  NANDN U3121 ( .A(start), .B(xreg[372]), .Z(n1396) );
  NAND U3122 ( .A(x[372]), .B(start), .Z(n1395) );
  NAND U3123 ( .A(n1397), .B(n1398), .Z(xin[371]) );
  NANDN U3124 ( .A(start), .B(xreg[371]), .Z(n1398) );
  NAND U3125 ( .A(x[371]), .B(start), .Z(n1397) );
  NAND U3126 ( .A(n1399), .B(n1400), .Z(xin[370]) );
  NANDN U3127 ( .A(start), .B(xreg[370]), .Z(n1400) );
  NAND U3128 ( .A(x[370]), .B(start), .Z(n1399) );
  NAND U3129 ( .A(n1401), .B(n1402), .Z(xin[36]) );
  NANDN U3130 ( .A(start), .B(xreg[36]), .Z(n1402) );
  NAND U3131 ( .A(x[36]), .B(start), .Z(n1401) );
  NAND U3132 ( .A(n1403), .B(n1404), .Z(xin[369]) );
  NANDN U3133 ( .A(start), .B(xreg[369]), .Z(n1404) );
  NAND U3134 ( .A(x[369]), .B(start), .Z(n1403) );
  NAND U3135 ( .A(n1405), .B(n1406), .Z(xin[368]) );
  NANDN U3136 ( .A(start), .B(xreg[368]), .Z(n1406) );
  NAND U3137 ( .A(x[368]), .B(start), .Z(n1405) );
  NAND U3138 ( .A(n1407), .B(n1408), .Z(xin[367]) );
  NANDN U3139 ( .A(start), .B(xreg[367]), .Z(n1408) );
  NAND U3140 ( .A(x[367]), .B(start), .Z(n1407) );
  NAND U3141 ( .A(n1409), .B(n1410), .Z(xin[366]) );
  NANDN U3142 ( .A(start), .B(xreg[366]), .Z(n1410) );
  NAND U3143 ( .A(x[366]), .B(start), .Z(n1409) );
  NAND U3144 ( .A(n1411), .B(n1412), .Z(xin[365]) );
  NANDN U3145 ( .A(start), .B(xreg[365]), .Z(n1412) );
  NAND U3146 ( .A(x[365]), .B(start), .Z(n1411) );
  NAND U3147 ( .A(n1413), .B(n1414), .Z(xin[364]) );
  NANDN U3148 ( .A(start), .B(xreg[364]), .Z(n1414) );
  NAND U3149 ( .A(x[364]), .B(start), .Z(n1413) );
  NAND U3150 ( .A(n1415), .B(n1416), .Z(xin[363]) );
  NANDN U3151 ( .A(start), .B(xreg[363]), .Z(n1416) );
  NAND U3152 ( .A(x[363]), .B(start), .Z(n1415) );
  NAND U3153 ( .A(n1417), .B(n1418), .Z(xin[362]) );
  NANDN U3154 ( .A(start), .B(xreg[362]), .Z(n1418) );
  NAND U3155 ( .A(x[362]), .B(start), .Z(n1417) );
  NAND U3156 ( .A(n1419), .B(n1420), .Z(xin[361]) );
  NANDN U3157 ( .A(start), .B(xreg[361]), .Z(n1420) );
  NAND U3158 ( .A(x[361]), .B(start), .Z(n1419) );
  NAND U3159 ( .A(n1421), .B(n1422), .Z(xin[360]) );
  NANDN U3160 ( .A(start), .B(xreg[360]), .Z(n1422) );
  NAND U3161 ( .A(x[360]), .B(start), .Z(n1421) );
  NAND U3162 ( .A(n1423), .B(n1424), .Z(xin[35]) );
  NANDN U3163 ( .A(start), .B(xreg[35]), .Z(n1424) );
  NAND U3164 ( .A(x[35]), .B(start), .Z(n1423) );
  NAND U3165 ( .A(n1425), .B(n1426), .Z(xin[359]) );
  NANDN U3166 ( .A(start), .B(xreg[359]), .Z(n1426) );
  NAND U3167 ( .A(x[359]), .B(start), .Z(n1425) );
  NAND U3168 ( .A(n1427), .B(n1428), .Z(xin[358]) );
  NANDN U3169 ( .A(start), .B(xreg[358]), .Z(n1428) );
  NAND U3170 ( .A(x[358]), .B(start), .Z(n1427) );
  NAND U3171 ( .A(n1429), .B(n1430), .Z(xin[357]) );
  NANDN U3172 ( .A(start), .B(xreg[357]), .Z(n1430) );
  NAND U3173 ( .A(x[357]), .B(start), .Z(n1429) );
  NAND U3174 ( .A(n1431), .B(n1432), .Z(xin[356]) );
  NANDN U3175 ( .A(start), .B(xreg[356]), .Z(n1432) );
  NAND U3176 ( .A(x[356]), .B(start), .Z(n1431) );
  NAND U3177 ( .A(n1433), .B(n1434), .Z(xin[355]) );
  NANDN U3178 ( .A(start), .B(xreg[355]), .Z(n1434) );
  NAND U3179 ( .A(x[355]), .B(start), .Z(n1433) );
  NAND U3180 ( .A(n1435), .B(n1436), .Z(xin[354]) );
  NANDN U3181 ( .A(start), .B(xreg[354]), .Z(n1436) );
  NAND U3182 ( .A(x[354]), .B(start), .Z(n1435) );
  NAND U3183 ( .A(n1437), .B(n1438), .Z(xin[353]) );
  NANDN U3184 ( .A(start), .B(xreg[353]), .Z(n1438) );
  NAND U3185 ( .A(x[353]), .B(start), .Z(n1437) );
  NAND U3186 ( .A(n1439), .B(n1440), .Z(xin[352]) );
  NANDN U3187 ( .A(start), .B(xreg[352]), .Z(n1440) );
  NAND U3188 ( .A(x[352]), .B(start), .Z(n1439) );
  NAND U3189 ( .A(n1441), .B(n1442), .Z(xin[351]) );
  NANDN U3190 ( .A(start), .B(xreg[351]), .Z(n1442) );
  NAND U3191 ( .A(x[351]), .B(start), .Z(n1441) );
  NAND U3192 ( .A(n1443), .B(n1444), .Z(xin[350]) );
  NANDN U3193 ( .A(start), .B(xreg[350]), .Z(n1444) );
  NAND U3194 ( .A(x[350]), .B(start), .Z(n1443) );
  NAND U3195 ( .A(n1445), .B(n1446), .Z(xin[34]) );
  NANDN U3196 ( .A(start), .B(xreg[34]), .Z(n1446) );
  NAND U3197 ( .A(x[34]), .B(start), .Z(n1445) );
  NAND U3198 ( .A(n1447), .B(n1448), .Z(xin[349]) );
  NANDN U3199 ( .A(start), .B(xreg[349]), .Z(n1448) );
  NAND U3200 ( .A(x[349]), .B(start), .Z(n1447) );
  NAND U3201 ( .A(n1449), .B(n1450), .Z(xin[348]) );
  NANDN U3202 ( .A(start), .B(xreg[348]), .Z(n1450) );
  NAND U3203 ( .A(x[348]), .B(start), .Z(n1449) );
  NAND U3204 ( .A(n1451), .B(n1452), .Z(xin[347]) );
  NANDN U3205 ( .A(start), .B(xreg[347]), .Z(n1452) );
  NAND U3206 ( .A(x[347]), .B(start), .Z(n1451) );
  NAND U3207 ( .A(n1453), .B(n1454), .Z(xin[346]) );
  NANDN U3208 ( .A(start), .B(xreg[346]), .Z(n1454) );
  NAND U3209 ( .A(x[346]), .B(start), .Z(n1453) );
  NAND U3210 ( .A(n1455), .B(n1456), .Z(xin[345]) );
  NANDN U3211 ( .A(start), .B(xreg[345]), .Z(n1456) );
  NAND U3212 ( .A(x[345]), .B(start), .Z(n1455) );
  NAND U3213 ( .A(n1457), .B(n1458), .Z(xin[344]) );
  NANDN U3214 ( .A(start), .B(xreg[344]), .Z(n1458) );
  NAND U3215 ( .A(x[344]), .B(start), .Z(n1457) );
  NAND U3216 ( .A(n1459), .B(n1460), .Z(xin[343]) );
  NANDN U3217 ( .A(start), .B(xreg[343]), .Z(n1460) );
  NAND U3218 ( .A(x[343]), .B(start), .Z(n1459) );
  NAND U3219 ( .A(n1461), .B(n1462), .Z(xin[342]) );
  NANDN U3220 ( .A(start), .B(xreg[342]), .Z(n1462) );
  NAND U3221 ( .A(x[342]), .B(start), .Z(n1461) );
  NAND U3222 ( .A(n1463), .B(n1464), .Z(xin[341]) );
  NANDN U3223 ( .A(start), .B(xreg[341]), .Z(n1464) );
  NAND U3224 ( .A(x[341]), .B(start), .Z(n1463) );
  NAND U3225 ( .A(n1465), .B(n1466), .Z(xin[340]) );
  NANDN U3226 ( .A(start), .B(xreg[340]), .Z(n1466) );
  NAND U3227 ( .A(x[340]), .B(start), .Z(n1465) );
  NAND U3228 ( .A(n1467), .B(n1468), .Z(xin[33]) );
  NANDN U3229 ( .A(start), .B(xreg[33]), .Z(n1468) );
  NAND U3230 ( .A(x[33]), .B(start), .Z(n1467) );
  NAND U3231 ( .A(n1469), .B(n1470), .Z(xin[339]) );
  NANDN U3232 ( .A(start), .B(xreg[339]), .Z(n1470) );
  NAND U3233 ( .A(x[339]), .B(start), .Z(n1469) );
  NAND U3234 ( .A(n1471), .B(n1472), .Z(xin[338]) );
  NANDN U3235 ( .A(start), .B(xreg[338]), .Z(n1472) );
  NAND U3236 ( .A(x[338]), .B(start), .Z(n1471) );
  NAND U3237 ( .A(n1473), .B(n1474), .Z(xin[337]) );
  NANDN U3238 ( .A(start), .B(xreg[337]), .Z(n1474) );
  NAND U3239 ( .A(x[337]), .B(start), .Z(n1473) );
  NAND U3240 ( .A(n1475), .B(n1476), .Z(xin[336]) );
  NANDN U3241 ( .A(start), .B(xreg[336]), .Z(n1476) );
  NAND U3242 ( .A(x[336]), .B(start), .Z(n1475) );
  NAND U3243 ( .A(n1477), .B(n1478), .Z(xin[335]) );
  NANDN U3244 ( .A(start), .B(xreg[335]), .Z(n1478) );
  NAND U3245 ( .A(x[335]), .B(start), .Z(n1477) );
  NAND U3246 ( .A(n1479), .B(n1480), .Z(xin[334]) );
  NANDN U3247 ( .A(start), .B(xreg[334]), .Z(n1480) );
  NAND U3248 ( .A(x[334]), .B(start), .Z(n1479) );
  NAND U3249 ( .A(n1481), .B(n1482), .Z(xin[333]) );
  NANDN U3250 ( .A(start), .B(xreg[333]), .Z(n1482) );
  NAND U3251 ( .A(x[333]), .B(start), .Z(n1481) );
  NAND U3252 ( .A(n1483), .B(n1484), .Z(xin[332]) );
  NANDN U3253 ( .A(start), .B(xreg[332]), .Z(n1484) );
  NAND U3254 ( .A(x[332]), .B(start), .Z(n1483) );
  NAND U3255 ( .A(n1485), .B(n1486), .Z(xin[331]) );
  NANDN U3256 ( .A(start), .B(xreg[331]), .Z(n1486) );
  NAND U3257 ( .A(x[331]), .B(start), .Z(n1485) );
  NAND U3258 ( .A(n1487), .B(n1488), .Z(xin[330]) );
  NANDN U3259 ( .A(start), .B(xreg[330]), .Z(n1488) );
  NAND U3260 ( .A(x[330]), .B(start), .Z(n1487) );
  NAND U3261 ( .A(n1489), .B(n1490), .Z(xin[32]) );
  NANDN U3262 ( .A(start), .B(xreg[32]), .Z(n1490) );
  NAND U3263 ( .A(x[32]), .B(start), .Z(n1489) );
  NAND U3264 ( .A(n1491), .B(n1492), .Z(xin[329]) );
  NANDN U3265 ( .A(start), .B(xreg[329]), .Z(n1492) );
  NAND U3266 ( .A(x[329]), .B(start), .Z(n1491) );
  NAND U3267 ( .A(n1493), .B(n1494), .Z(xin[328]) );
  NANDN U3268 ( .A(start), .B(xreg[328]), .Z(n1494) );
  NAND U3269 ( .A(x[328]), .B(start), .Z(n1493) );
  NAND U3270 ( .A(n1495), .B(n1496), .Z(xin[327]) );
  NANDN U3271 ( .A(start), .B(xreg[327]), .Z(n1496) );
  NAND U3272 ( .A(x[327]), .B(start), .Z(n1495) );
  NAND U3273 ( .A(n1497), .B(n1498), .Z(xin[326]) );
  NANDN U3274 ( .A(start), .B(xreg[326]), .Z(n1498) );
  NAND U3275 ( .A(x[326]), .B(start), .Z(n1497) );
  NAND U3276 ( .A(n1499), .B(n1500), .Z(xin[325]) );
  NANDN U3277 ( .A(start), .B(xreg[325]), .Z(n1500) );
  NAND U3278 ( .A(x[325]), .B(start), .Z(n1499) );
  NAND U3279 ( .A(n1501), .B(n1502), .Z(xin[324]) );
  NANDN U3280 ( .A(start), .B(xreg[324]), .Z(n1502) );
  NAND U3281 ( .A(x[324]), .B(start), .Z(n1501) );
  NAND U3282 ( .A(n1503), .B(n1504), .Z(xin[323]) );
  NANDN U3283 ( .A(start), .B(xreg[323]), .Z(n1504) );
  NAND U3284 ( .A(x[323]), .B(start), .Z(n1503) );
  NAND U3285 ( .A(n1505), .B(n1506), .Z(xin[322]) );
  NANDN U3286 ( .A(start), .B(xreg[322]), .Z(n1506) );
  NAND U3287 ( .A(x[322]), .B(start), .Z(n1505) );
  NAND U3288 ( .A(n1507), .B(n1508), .Z(xin[321]) );
  NANDN U3289 ( .A(start), .B(xreg[321]), .Z(n1508) );
  NAND U3290 ( .A(x[321]), .B(start), .Z(n1507) );
  NAND U3291 ( .A(n1509), .B(n1510), .Z(xin[320]) );
  NANDN U3292 ( .A(start), .B(xreg[320]), .Z(n1510) );
  NAND U3293 ( .A(x[320]), .B(start), .Z(n1509) );
  NAND U3294 ( .A(n1511), .B(n1512), .Z(xin[31]) );
  NANDN U3295 ( .A(start), .B(xreg[31]), .Z(n1512) );
  NAND U3296 ( .A(x[31]), .B(start), .Z(n1511) );
  NAND U3297 ( .A(n1513), .B(n1514), .Z(xin[319]) );
  NANDN U3298 ( .A(start), .B(xreg[319]), .Z(n1514) );
  NAND U3299 ( .A(x[319]), .B(start), .Z(n1513) );
  NAND U3300 ( .A(n1515), .B(n1516), .Z(xin[318]) );
  NANDN U3301 ( .A(start), .B(xreg[318]), .Z(n1516) );
  NAND U3302 ( .A(x[318]), .B(start), .Z(n1515) );
  NAND U3303 ( .A(n1517), .B(n1518), .Z(xin[317]) );
  NANDN U3304 ( .A(start), .B(xreg[317]), .Z(n1518) );
  NAND U3305 ( .A(x[317]), .B(start), .Z(n1517) );
  NAND U3306 ( .A(n1519), .B(n1520), .Z(xin[316]) );
  NANDN U3307 ( .A(start), .B(xreg[316]), .Z(n1520) );
  NAND U3308 ( .A(x[316]), .B(start), .Z(n1519) );
  NAND U3309 ( .A(n1521), .B(n1522), .Z(xin[315]) );
  NANDN U3310 ( .A(start), .B(xreg[315]), .Z(n1522) );
  NAND U3311 ( .A(x[315]), .B(start), .Z(n1521) );
  NAND U3312 ( .A(n1523), .B(n1524), .Z(xin[314]) );
  NANDN U3313 ( .A(start), .B(xreg[314]), .Z(n1524) );
  NAND U3314 ( .A(x[314]), .B(start), .Z(n1523) );
  NAND U3315 ( .A(n1525), .B(n1526), .Z(xin[313]) );
  NANDN U3316 ( .A(start), .B(xreg[313]), .Z(n1526) );
  NAND U3317 ( .A(x[313]), .B(start), .Z(n1525) );
  NAND U3318 ( .A(n1527), .B(n1528), .Z(xin[312]) );
  NANDN U3319 ( .A(start), .B(xreg[312]), .Z(n1528) );
  NAND U3320 ( .A(x[312]), .B(start), .Z(n1527) );
  NAND U3321 ( .A(n1529), .B(n1530), .Z(xin[311]) );
  NANDN U3322 ( .A(start), .B(xreg[311]), .Z(n1530) );
  NAND U3323 ( .A(x[311]), .B(start), .Z(n1529) );
  NAND U3324 ( .A(n1531), .B(n1532), .Z(xin[310]) );
  NANDN U3325 ( .A(start), .B(xreg[310]), .Z(n1532) );
  NAND U3326 ( .A(x[310]), .B(start), .Z(n1531) );
  NAND U3327 ( .A(n1533), .B(n1534), .Z(xin[30]) );
  NANDN U3328 ( .A(start), .B(xreg[30]), .Z(n1534) );
  NAND U3329 ( .A(x[30]), .B(start), .Z(n1533) );
  NAND U3330 ( .A(n1535), .B(n1536), .Z(xin[309]) );
  NANDN U3331 ( .A(start), .B(xreg[309]), .Z(n1536) );
  NAND U3332 ( .A(x[309]), .B(start), .Z(n1535) );
  NAND U3333 ( .A(n1537), .B(n1538), .Z(xin[308]) );
  NANDN U3334 ( .A(start), .B(xreg[308]), .Z(n1538) );
  NAND U3335 ( .A(x[308]), .B(start), .Z(n1537) );
  NAND U3336 ( .A(n1539), .B(n1540), .Z(xin[307]) );
  NANDN U3337 ( .A(start), .B(xreg[307]), .Z(n1540) );
  NAND U3338 ( .A(x[307]), .B(start), .Z(n1539) );
  NAND U3339 ( .A(n1541), .B(n1542), .Z(xin[306]) );
  NANDN U3340 ( .A(start), .B(xreg[306]), .Z(n1542) );
  NAND U3341 ( .A(x[306]), .B(start), .Z(n1541) );
  NAND U3342 ( .A(n1543), .B(n1544), .Z(xin[305]) );
  NANDN U3343 ( .A(start), .B(xreg[305]), .Z(n1544) );
  NAND U3344 ( .A(x[305]), .B(start), .Z(n1543) );
  NAND U3345 ( .A(n1545), .B(n1546), .Z(xin[304]) );
  NANDN U3346 ( .A(start), .B(xreg[304]), .Z(n1546) );
  NAND U3347 ( .A(x[304]), .B(start), .Z(n1545) );
  NAND U3348 ( .A(n1547), .B(n1548), .Z(xin[303]) );
  NANDN U3349 ( .A(start), .B(xreg[303]), .Z(n1548) );
  NAND U3350 ( .A(x[303]), .B(start), .Z(n1547) );
  NAND U3351 ( .A(n1549), .B(n1550), .Z(xin[302]) );
  NANDN U3352 ( .A(start), .B(xreg[302]), .Z(n1550) );
  NAND U3353 ( .A(x[302]), .B(start), .Z(n1549) );
  NAND U3354 ( .A(n1551), .B(n1552), .Z(xin[301]) );
  NANDN U3355 ( .A(start), .B(xreg[301]), .Z(n1552) );
  NAND U3356 ( .A(x[301]), .B(start), .Z(n1551) );
  NAND U3357 ( .A(n1553), .B(n1554), .Z(xin[300]) );
  NANDN U3358 ( .A(start), .B(xreg[300]), .Z(n1554) );
  NAND U3359 ( .A(x[300]), .B(start), .Z(n1553) );
  NAND U3360 ( .A(n1555), .B(n1556), .Z(xin[2]) );
  NANDN U3361 ( .A(start), .B(xreg[2]), .Z(n1556) );
  NAND U3362 ( .A(x[2]), .B(start), .Z(n1555) );
  NAND U3363 ( .A(n1557), .B(n1558), .Z(xin[29]) );
  NANDN U3364 ( .A(start), .B(xreg[29]), .Z(n1558) );
  NAND U3365 ( .A(x[29]), .B(start), .Z(n1557) );
  NAND U3366 ( .A(n1559), .B(n1560), .Z(xin[299]) );
  NANDN U3367 ( .A(start), .B(xreg[299]), .Z(n1560) );
  NAND U3368 ( .A(x[299]), .B(start), .Z(n1559) );
  NAND U3369 ( .A(n1561), .B(n1562), .Z(xin[298]) );
  NANDN U3370 ( .A(start), .B(xreg[298]), .Z(n1562) );
  NAND U3371 ( .A(x[298]), .B(start), .Z(n1561) );
  NAND U3372 ( .A(n1563), .B(n1564), .Z(xin[297]) );
  NANDN U3373 ( .A(start), .B(xreg[297]), .Z(n1564) );
  NAND U3374 ( .A(x[297]), .B(start), .Z(n1563) );
  NAND U3375 ( .A(n1565), .B(n1566), .Z(xin[296]) );
  NANDN U3376 ( .A(start), .B(xreg[296]), .Z(n1566) );
  NAND U3377 ( .A(x[296]), .B(start), .Z(n1565) );
  NAND U3378 ( .A(n1567), .B(n1568), .Z(xin[295]) );
  NANDN U3379 ( .A(start), .B(xreg[295]), .Z(n1568) );
  NAND U3380 ( .A(x[295]), .B(start), .Z(n1567) );
  NAND U3381 ( .A(n1569), .B(n1570), .Z(xin[294]) );
  NANDN U3382 ( .A(start), .B(xreg[294]), .Z(n1570) );
  NAND U3383 ( .A(x[294]), .B(start), .Z(n1569) );
  NAND U3384 ( .A(n1571), .B(n1572), .Z(xin[293]) );
  NANDN U3385 ( .A(start), .B(xreg[293]), .Z(n1572) );
  NAND U3386 ( .A(x[293]), .B(start), .Z(n1571) );
  NAND U3387 ( .A(n1573), .B(n1574), .Z(xin[292]) );
  NANDN U3388 ( .A(start), .B(xreg[292]), .Z(n1574) );
  NAND U3389 ( .A(x[292]), .B(start), .Z(n1573) );
  NAND U3390 ( .A(n1575), .B(n1576), .Z(xin[291]) );
  NANDN U3391 ( .A(start), .B(xreg[291]), .Z(n1576) );
  NAND U3392 ( .A(x[291]), .B(start), .Z(n1575) );
  NAND U3393 ( .A(n1577), .B(n1578), .Z(xin[290]) );
  NANDN U3394 ( .A(start), .B(xreg[290]), .Z(n1578) );
  NAND U3395 ( .A(x[290]), .B(start), .Z(n1577) );
  NAND U3396 ( .A(n1579), .B(n1580), .Z(xin[28]) );
  NANDN U3397 ( .A(start), .B(xreg[28]), .Z(n1580) );
  NAND U3398 ( .A(x[28]), .B(start), .Z(n1579) );
  NAND U3399 ( .A(n1581), .B(n1582), .Z(xin[289]) );
  NANDN U3400 ( .A(start), .B(xreg[289]), .Z(n1582) );
  NAND U3401 ( .A(x[289]), .B(start), .Z(n1581) );
  NAND U3402 ( .A(n1583), .B(n1584), .Z(xin[288]) );
  NANDN U3403 ( .A(start), .B(xreg[288]), .Z(n1584) );
  NAND U3404 ( .A(x[288]), .B(start), .Z(n1583) );
  NAND U3405 ( .A(n1585), .B(n1586), .Z(xin[287]) );
  NANDN U3406 ( .A(start), .B(xreg[287]), .Z(n1586) );
  NAND U3407 ( .A(x[287]), .B(start), .Z(n1585) );
  NAND U3408 ( .A(n1587), .B(n1588), .Z(xin[286]) );
  NANDN U3409 ( .A(start), .B(xreg[286]), .Z(n1588) );
  NAND U3410 ( .A(x[286]), .B(start), .Z(n1587) );
  NAND U3411 ( .A(n1589), .B(n1590), .Z(xin[285]) );
  NANDN U3412 ( .A(start), .B(xreg[285]), .Z(n1590) );
  NAND U3413 ( .A(x[285]), .B(start), .Z(n1589) );
  NAND U3414 ( .A(n1591), .B(n1592), .Z(xin[284]) );
  NANDN U3415 ( .A(start), .B(xreg[284]), .Z(n1592) );
  NAND U3416 ( .A(x[284]), .B(start), .Z(n1591) );
  NAND U3417 ( .A(n1593), .B(n1594), .Z(xin[283]) );
  NANDN U3418 ( .A(start), .B(xreg[283]), .Z(n1594) );
  NAND U3419 ( .A(x[283]), .B(start), .Z(n1593) );
  NAND U3420 ( .A(n1595), .B(n1596), .Z(xin[282]) );
  NANDN U3421 ( .A(start), .B(xreg[282]), .Z(n1596) );
  NAND U3422 ( .A(x[282]), .B(start), .Z(n1595) );
  NAND U3423 ( .A(n1597), .B(n1598), .Z(xin[281]) );
  NANDN U3424 ( .A(start), .B(xreg[281]), .Z(n1598) );
  NAND U3425 ( .A(x[281]), .B(start), .Z(n1597) );
  NAND U3426 ( .A(n1599), .B(n1600), .Z(xin[280]) );
  NANDN U3427 ( .A(start), .B(xreg[280]), .Z(n1600) );
  NAND U3428 ( .A(x[280]), .B(start), .Z(n1599) );
  NAND U3429 ( .A(n1601), .B(n1602), .Z(xin[27]) );
  NANDN U3430 ( .A(start), .B(xreg[27]), .Z(n1602) );
  NAND U3431 ( .A(x[27]), .B(start), .Z(n1601) );
  NAND U3432 ( .A(n1603), .B(n1604), .Z(xin[279]) );
  NANDN U3433 ( .A(start), .B(xreg[279]), .Z(n1604) );
  NAND U3434 ( .A(x[279]), .B(start), .Z(n1603) );
  NAND U3435 ( .A(n1605), .B(n1606), .Z(xin[278]) );
  NANDN U3436 ( .A(start), .B(xreg[278]), .Z(n1606) );
  NAND U3437 ( .A(x[278]), .B(start), .Z(n1605) );
  NAND U3438 ( .A(n1607), .B(n1608), .Z(xin[277]) );
  NANDN U3439 ( .A(start), .B(xreg[277]), .Z(n1608) );
  NAND U3440 ( .A(x[277]), .B(start), .Z(n1607) );
  NAND U3441 ( .A(n1609), .B(n1610), .Z(xin[276]) );
  NANDN U3442 ( .A(start), .B(xreg[276]), .Z(n1610) );
  NAND U3443 ( .A(x[276]), .B(start), .Z(n1609) );
  NAND U3444 ( .A(n1611), .B(n1612), .Z(xin[275]) );
  NANDN U3445 ( .A(start), .B(xreg[275]), .Z(n1612) );
  NAND U3446 ( .A(x[275]), .B(start), .Z(n1611) );
  NAND U3447 ( .A(n1613), .B(n1614), .Z(xin[274]) );
  NANDN U3448 ( .A(start), .B(xreg[274]), .Z(n1614) );
  NAND U3449 ( .A(x[274]), .B(start), .Z(n1613) );
  NAND U3450 ( .A(n1615), .B(n1616), .Z(xin[273]) );
  NANDN U3451 ( .A(start), .B(xreg[273]), .Z(n1616) );
  NAND U3452 ( .A(x[273]), .B(start), .Z(n1615) );
  NAND U3453 ( .A(n1617), .B(n1618), .Z(xin[272]) );
  NANDN U3454 ( .A(start), .B(xreg[272]), .Z(n1618) );
  NAND U3455 ( .A(x[272]), .B(start), .Z(n1617) );
  NAND U3456 ( .A(n1619), .B(n1620), .Z(xin[271]) );
  NANDN U3457 ( .A(start), .B(xreg[271]), .Z(n1620) );
  NAND U3458 ( .A(x[271]), .B(start), .Z(n1619) );
  NAND U3459 ( .A(n1621), .B(n1622), .Z(xin[270]) );
  NANDN U3460 ( .A(start), .B(xreg[270]), .Z(n1622) );
  NAND U3461 ( .A(x[270]), .B(start), .Z(n1621) );
  NAND U3462 ( .A(n1623), .B(n1624), .Z(xin[26]) );
  NANDN U3463 ( .A(start), .B(xreg[26]), .Z(n1624) );
  NAND U3464 ( .A(x[26]), .B(start), .Z(n1623) );
  NAND U3465 ( .A(n1625), .B(n1626), .Z(xin[269]) );
  NANDN U3466 ( .A(start), .B(xreg[269]), .Z(n1626) );
  NAND U3467 ( .A(x[269]), .B(start), .Z(n1625) );
  NAND U3468 ( .A(n1627), .B(n1628), .Z(xin[268]) );
  NANDN U3469 ( .A(start), .B(xreg[268]), .Z(n1628) );
  NAND U3470 ( .A(x[268]), .B(start), .Z(n1627) );
  NAND U3471 ( .A(n1629), .B(n1630), .Z(xin[267]) );
  NANDN U3472 ( .A(start), .B(xreg[267]), .Z(n1630) );
  NAND U3473 ( .A(x[267]), .B(start), .Z(n1629) );
  NAND U3474 ( .A(n1631), .B(n1632), .Z(xin[266]) );
  NANDN U3475 ( .A(start), .B(xreg[266]), .Z(n1632) );
  NAND U3476 ( .A(x[266]), .B(start), .Z(n1631) );
  NAND U3477 ( .A(n1633), .B(n1634), .Z(xin[265]) );
  NANDN U3478 ( .A(start), .B(xreg[265]), .Z(n1634) );
  NAND U3479 ( .A(x[265]), .B(start), .Z(n1633) );
  NAND U3480 ( .A(n1635), .B(n1636), .Z(xin[264]) );
  NANDN U3481 ( .A(start), .B(xreg[264]), .Z(n1636) );
  NAND U3482 ( .A(x[264]), .B(start), .Z(n1635) );
  NAND U3483 ( .A(n1637), .B(n1638), .Z(xin[263]) );
  NANDN U3484 ( .A(start), .B(xreg[263]), .Z(n1638) );
  NAND U3485 ( .A(x[263]), .B(start), .Z(n1637) );
  NAND U3486 ( .A(n1639), .B(n1640), .Z(xin[262]) );
  NANDN U3487 ( .A(start), .B(xreg[262]), .Z(n1640) );
  NAND U3488 ( .A(x[262]), .B(start), .Z(n1639) );
  NAND U3489 ( .A(n1641), .B(n1642), .Z(xin[261]) );
  NANDN U3490 ( .A(start), .B(xreg[261]), .Z(n1642) );
  NAND U3491 ( .A(x[261]), .B(start), .Z(n1641) );
  NAND U3492 ( .A(n1643), .B(n1644), .Z(xin[260]) );
  NANDN U3493 ( .A(start), .B(xreg[260]), .Z(n1644) );
  NAND U3494 ( .A(x[260]), .B(start), .Z(n1643) );
  NAND U3495 ( .A(n1645), .B(n1646), .Z(xin[25]) );
  NANDN U3496 ( .A(start), .B(xreg[25]), .Z(n1646) );
  NAND U3497 ( .A(x[25]), .B(start), .Z(n1645) );
  NAND U3498 ( .A(n1647), .B(n1648), .Z(xin[259]) );
  NANDN U3499 ( .A(start), .B(xreg[259]), .Z(n1648) );
  NAND U3500 ( .A(x[259]), .B(start), .Z(n1647) );
  NAND U3501 ( .A(n1649), .B(n1650), .Z(xin[258]) );
  NANDN U3502 ( .A(start), .B(xreg[258]), .Z(n1650) );
  NAND U3503 ( .A(x[258]), .B(start), .Z(n1649) );
  NAND U3504 ( .A(n1651), .B(n1652), .Z(xin[257]) );
  NANDN U3505 ( .A(start), .B(xreg[257]), .Z(n1652) );
  NAND U3506 ( .A(x[257]), .B(start), .Z(n1651) );
  NAND U3507 ( .A(n1653), .B(n1654), .Z(xin[256]) );
  NANDN U3508 ( .A(start), .B(xreg[256]), .Z(n1654) );
  NAND U3509 ( .A(x[256]), .B(start), .Z(n1653) );
  NAND U3510 ( .A(n1655), .B(n1656), .Z(xin[255]) );
  NANDN U3511 ( .A(start), .B(xreg[255]), .Z(n1656) );
  NAND U3512 ( .A(x[255]), .B(start), .Z(n1655) );
  NAND U3513 ( .A(n1657), .B(n1658), .Z(xin[254]) );
  NANDN U3514 ( .A(start), .B(xreg[254]), .Z(n1658) );
  NAND U3515 ( .A(x[254]), .B(start), .Z(n1657) );
  NAND U3516 ( .A(n1659), .B(n1660), .Z(xin[253]) );
  NANDN U3517 ( .A(start), .B(xreg[253]), .Z(n1660) );
  NAND U3518 ( .A(x[253]), .B(start), .Z(n1659) );
  NAND U3519 ( .A(n1661), .B(n1662), .Z(xin[252]) );
  NANDN U3520 ( .A(start), .B(xreg[252]), .Z(n1662) );
  NAND U3521 ( .A(x[252]), .B(start), .Z(n1661) );
  NAND U3522 ( .A(n1663), .B(n1664), .Z(xin[251]) );
  NANDN U3523 ( .A(start), .B(xreg[251]), .Z(n1664) );
  NAND U3524 ( .A(x[251]), .B(start), .Z(n1663) );
  NAND U3525 ( .A(n1665), .B(n1666), .Z(xin[250]) );
  NANDN U3526 ( .A(start), .B(xreg[250]), .Z(n1666) );
  NAND U3527 ( .A(x[250]), .B(start), .Z(n1665) );
  NAND U3528 ( .A(n1667), .B(n1668), .Z(xin[24]) );
  NANDN U3529 ( .A(start), .B(xreg[24]), .Z(n1668) );
  NAND U3530 ( .A(x[24]), .B(start), .Z(n1667) );
  NAND U3531 ( .A(n1669), .B(n1670), .Z(xin[249]) );
  NANDN U3532 ( .A(start), .B(xreg[249]), .Z(n1670) );
  NAND U3533 ( .A(x[249]), .B(start), .Z(n1669) );
  NAND U3534 ( .A(n1671), .B(n1672), .Z(xin[248]) );
  NANDN U3535 ( .A(start), .B(xreg[248]), .Z(n1672) );
  NAND U3536 ( .A(x[248]), .B(start), .Z(n1671) );
  NAND U3537 ( .A(n1673), .B(n1674), .Z(xin[247]) );
  NANDN U3538 ( .A(start), .B(xreg[247]), .Z(n1674) );
  NAND U3539 ( .A(x[247]), .B(start), .Z(n1673) );
  NAND U3540 ( .A(n1675), .B(n1676), .Z(xin[246]) );
  NANDN U3541 ( .A(start), .B(xreg[246]), .Z(n1676) );
  NAND U3542 ( .A(x[246]), .B(start), .Z(n1675) );
  NAND U3543 ( .A(n1677), .B(n1678), .Z(xin[245]) );
  NANDN U3544 ( .A(start), .B(xreg[245]), .Z(n1678) );
  NAND U3545 ( .A(x[245]), .B(start), .Z(n1677) );
  NAND U3546 ( .A(n1679), .B(n1680), .Z(xin[244]) );
  NANDN U3547 ( .A(start), .B(xreg[244]), .Z(n1680) );
  NAND U3548 ( .A(x[244]), .B(start), .Z(n1679) );
  NAND U3549 ( .A(n1681), .B(n1682), .Z(xin[243]) );
  NANDN U3550 ( .A(start), .B(xreg[243]), .Z(n1682) );
  NAND U3551 ( .A(x[243]), .B(start), .Z(n1681) );
  NAND U3552 ( .A(n1683), .B(n1684), .Z(xin[242]) );
  NANDN U3553 ( .A(start), .B(xreg[242]), .Z(n1684) );
  NAND U3554 ( .A(x[242]), .B(start), .Z(n1683) );
  NAND U3555 ( .A(n1685), .B(n1686), .Z(xin[241]) );
  NANDN U3556 ( .A(start), .B(xreg[241]), .Z(n1686) );
  NAND U3557 ( .A(x[241]), .B(start), .Z(n1685) );
  NAND U3558 ( .A(n1687), .B(n1688), .Z(xin[240]) );
  NANDN U3559 ( .A(start), .B(xreg[240]), .Z(n1688) );
  NAND U3560 ( .A(x[240]), .B(start), .Z(n1687) );
  NAND U3561 ( .A(n1689), .B(n1690), .Z(xin[23]) );
  NANDN U3562 ( .A(start), .B(xreg[23]), .Z(n1690) );
  NAND U3563 ( .A(x[23]), .B(start), .Z(n1689) );
  NAND U3564 ( .A(n1691), .B(n1692), .Z(xin[239]) );
  NANDN U3565 ( .A(start), .B(xreg[239]), .Z(n1692) );
  NAND U3566 ( .A(x[239]), .B(start), .Z(n1691) );
  NAND U3567 ( .A(n1693), .B(n1694), .Z(xin[238]) );
  NANDN U3568 ( .A(start), .B(xreg[238]), .Z(n1694) );
  NAND U3569 ( .A(x[238]), .B(start), .Z(n1693) );
  NAND U3570 ( .A(n1695), .B(n1696), .Z(xin[237]) );
  NANDN U3571 ( .A(start), .B(xreg[237]), .Z(n1696) );
  NAND U3572 ( .A(x[237]), .B(start), .Z(n1695) );
  NAND U3573 ( .A(n1697), .B(n1698), .Z(xin[236]) );
  NANDN U3574 ( .A(start), .B(xreg[236]), .Z(n1698) );
  NAND U3575 ( .A(x[236]), .B(start), .Z(n1697) );
  NAND U3576 ( .A(n1699), .B(n1700), .Z(xin[235]) );
  NANDN U3577 ( .A(start), .B(xreg[235]), .Z(n1700) );
  NAND U3578 ( .A(x[235]), .B(start), .Z(n1699) );
  NAND U3579 ( .A(n1701), .B(n1702), .Z(xin[234]) );
  NANDN U3580 ( .A(start), .B(xreg[234]), .Z(n1702) );
  NAND U3581 ( .A(x[234]), .B(start), .Z(n1701) );
  NAND U3582 ( .A(n1703), .B(n1704), .Z(xin[233]) );
  NANDN U3583 ( .A(start), .B(xreg[233]), .Z(n1704) );
  NAND U3584 ( .A(x[233]), .B(start), .Z(n1703) );
  NAND U3585 ( .A(n1705), .B(n1706), .Z(xin[232]) );
  NANDN U3586 ( .A(start), .B(xreg[232]), .Z(n1706) );
  NAND U3587 ( .A(x[232]), .B(start), .Z(n1705) );
  NAND U3588 ( .A(n1707), .B(n1708), .Z(xin[231]) );
  NANDN U3589 ( .A(start), .B(xreg[231]), .Z(n1708) );
  NAND U3590 ( .A(x[231]), .B(start), .Z(n1707) );
  NAND U3591 ( .A(n1709), .B(n1710), .Z(xin[230]) );
  NANDN U3592 ( .A(start), .B(xreg[230]), .Z(n1710) );
  NAND U3593 ( .A(x[230]), .B(start), .Z(n1709) );
  NAND U3594 ( .A(n1711), .B(n1712), .Z(xin[22]) );
  NANDN U3595 ( .A(start), .B(xreg[22]), .Z(n1712) );
  NAND U3596 ( .A(x[22]), .B(start), .Z(n1711) );
  NAND U3597 ( .A(n1713), .B(n1714), .Z(xin[229]) );
  NANDN U3598 ( .A(start), .B(xreg[229]), .Z(n1714) );
  NAND U3599 ( .A(x[229]), .B(start), .Z(n1713) );
  NAND U3600 ( .A(n1715), .B(n1716), .Z(xin[228]) );
  NANDN U3601 ( .A(start), .B(xreg[228]), .Z(n1716) );
  NAND U3602 ( .A(x[228]), .B(start), .Z(n1715) );
  NAND U3603 ( .A(n1717), .B(n1718), .Z(xin[227]) );
  NANDN U3604 ( .A(start), .B(xreg[227]), .Z(n1718) );
  NAND U3605 ( .A(x[227]), .B(start), .Z(n1717) );
  NAND U3606 ( .A(n1719), .B(n1720), .Z(xin[226]) );
  NANDN U3607 ( .A(start), .B(xreg[226]), .Z(n1720) );
  NAND U3608 ( .A(x[226]), .B(start), .Z(n1719) );
  NAND U3609 ( .A(n1721), .B(n1722), .Z(xin[225]) );
  NANDN U3610 ( .A(start), .B(xreg[225]), .Z(n1722) );
  NAND U3611 ( .A(x[225]), .B(start), .Z(n1721) );
  NAND U3612 ( .A(n1723), .B(n1724), .Z(xin[224]) );
  NANDN U3613 ( .A(start), .B(xreg[224]), .Z(n1724) );
  NAND U3614 ( .A(x[224]), .B(start), .Z(n1723) );
  NAND U3615 ( .A(n1725), .B(n1726), .Z(xin[223]) );
  NANDN U3616 ( .A(start), .B(xreg[223]), .Z(n1726) );
  NAND U3617 ( .A(x[223]), .B(start), .Z(n1725) );
  NAND U3618 ( .A(n1727), .B(n1728), .Z(xin[222]) );
  NANDN U3619 ( .A(start), .B(xreg[222]), .Z(n1728) );
  NAND U3620 ( .A(x[222]), .B(start), .Z(n1727) );
  NAND U3621 ( .A(n1729), .B(n1730), .Z(xin[221]) );
  NANDN U3622 ( .A(start), .B(xreg[221]), .Z(n1730) );
  NAND U3623 ( .A(x[221]), .B(start), .Z(n1729) );
  NAND U3624 ( .A(n1731), .B(n1732), .Z(xin[220]) );
  NANDN U3625 ( .A(start), .B(xreg[220]), .Z(n1732) );
  NAND U3626 ( .A(x[220]), .B(start), .Z(n1731) );
  NAND U3627 ( .A(n1733), .B(n1734), .Z(xin[21]) );
  NANDN U3628 ( .A(start), .B(xreg[21]), .Z(n1734) );
  NAND U3629 ( .A(x[21]), .B(start), .Z(n1733) );
  NAND U3630 ( .A(n1735), .B(n1736), .Z(xin[219]) );
  NANDN U3631 ( .A(start), .B(xreg[219]), .Z(n1736) );
  NAND U3632 ( .A(x[219]), .B(start), .Z(n1735) );
  NAND U3633 ( .A(n1737), .B(n1738), .Z(xin[218]) );
  NANDN U3634 ( .A(start), .B(xreg[218]), .Z(n1738) );
  NAND U3635 ( .A(x[218]), .B(start), .Z(n1737) );
  NAND U3636 ( .A(n1739), .B(n1740), .Z(xin[217]) );
  NANDN U3637 ( .A(start), .B(xreg[217]), .Z(n1740) );
  NAND U3638 ( .A(x[217]), .B(start), .Z(n1739) );
  NAND U3639 ( .A(n1741), .B(n1742), .Z(xin[216]) );
  NANDN U3640 ( .A(start), .B(xreg[216]), .Z(n1742) );
  NAND U3641 ( .A(x[216]), .B(start), .Z(n1741) );
  NAND U3642 ( .A(n1743), .B(n1744), .Z(xin[215]) );
  NANDN U3643 ( .A(start), .B(xreg[215]), .Z(n1744) );
  NAND U3644 ( .A(x[215]), .B(start), .Z(n1743) );
  NAND U3645 ( .A(n1745), .B(n1746), .Z(xin[214]) );
  NANDN U3646 ( .A(start), .B(xreg[214]), .Z(n1746) );
  NAND U3647 ( .A(x[214]), .B(start), .Z(n1745) );
  NAND U3648 ( .A(n1747), .B(n1748), .Z(xin[213]) );
  NANDN U3649 ( .A(start), .B(xreg[213]), .Z(n1748) );
  NAND U3650 ( .A(x[213]), .B(start), .Z(n1747) );
  NAND U3651 ( .A(n1749), .B(n1750), .Z(xin[212]) );
  NANDN U3652 ( .A(start), .B(xreg[212]), .Z(n1750) );
  NAND U3653 ( .A(x[212]), .B(start), .Z(n1749) );
  NAND U3654 ( .A(n1751), .B(n1752), .Z(xin[211]) );
  NANDN U3655 ( .A(start), .B(xreg[211]), .Z(n1752) );
  NAND U3656 ( .A(x[211]), .B(start), .Z(n1751) );
  NAND U3657 ( .A(n1753), .B(n1754), .Z(xin[210]) );
  NANDN U3658 ( .A(start), .B(xreg[210]), .Z(n1754) );
  NAND U3659 ( .A(x[210]), .B(start), .Z(n1753) );
  NAND U3660 ( .A(n1755), .B(n1756), .Z(xin[20]) );
  NANDN U3661 ( .A(start), .B(xreg[20]), .Z(n1756) );
  NAND U3662 ( .A(x[20]), .B(start), .Z(n1755) );
  NAND U3663 ( .A(n1757), .B(n1758), .Z(xin[209]) );
  NANDN U3664 ( .A(start), .B(xreg[209]), .Z(n1758) );
  NAND U3665 ( .A(x[209]), .B(start), .Z(n1757) );
  NAND U3666 ( .A(n1759), .B(n1760), .Z(xin[208]) );
  NANDN U3667 ( .A(start), .B(xreg[208]), .Z(n1760) );
  NAND U3668 ( .A(x[208]), .B(start), .Z(n1759) );
  NAND U3669 ( .A(n1761), .B(n1762), .Z(xin[207]) );
  NANDN U3670 ( .A(start), .B(xreg[207]), .Z(n1762) );
  NAND U3671 ( .A(x[207]), .B(start), .Z(n1761) );
  NAND U3672 ( .A(n1763), .B(n1764), .Z(xin[206]) );
  NANDN U3673 ( .A(start), .B(xreg[206]), .Z(n1764) );
  NAND U3674 ( .A(x[206]), .B(start), .Z(n1763) );
  NAND U3675 ( .A(n1765), .B(n1766), .Z(xin[205]) );
  NANDN U3676 ( .A(start), .B(xreg[205]), .Z(n1766) );
  NAND U3677 ( .A(x[205]), .B(start), .Z(n1765) );
  NAND U3678 ( .A(n1767), .B(n1768), .Z(xin[204]) );
  NANDN U3679 ( .A(start), .B(xreg[204]), .Z(n1768) );
  NAND U3680 ( .A(x[204]), .B(start), .Z(n1767) );
  NAND U3681 ( .A(n1769), .B(n1770), .Z(xin[203]) );
  NANDN U3682 ( .A(start), .B(xreg[203]), .Z(n1770) );
  NAND U3683 ( .A(x[203]), .B(start), .Z(n1769) );
  NAND U3684 ( .A(n1771), .B(n1772), .Z(xin[202]) );
  NANDN U3685 ( .A(start), .B(xreg[202]), .Z(n1772) );
  NAND U3686 ( .A(x[202]), .B(start), .Z(n1771) );
  NAND U3687 ( .A(n1773), .B(n1774), .Z(xin[201]) );
  NANDN U3688 ( .A(start), .B(xreg[201]), .Z(n1774) );
  NAND U3689 ( .A(x[201]), .B(start), .Z(n1773) );
  NAND U3690 ( .A(n1775), .B(n1776), .Z(xin[200]) );
  NANDN U3691 ( .A(start), .B(xreg[200]), .Z(n1776) );
  NAND U3692 ( .A(x[200]), .B(start), .Z(n1775) );
  NAND U3693 ( .A(n1777), .B(n1778), .Z(xin[1]) );
  NANDN U3694 ( .A(start), .B(xreg[1]), .Z(n1778) );
  NAND U3695 ( .A(x[1]), .B(start), .Z(n1777) );
  NAND U3696 ( .A(n1779), .B(n1780), .Z(xin[19]) );
  NANDN U3697 ( .A(start), .B(xreg[19]), .Z(n1780) );
  NAND U3698 ( .A(x[19]), .B(start), .Z(n1779) );
  NAND U3699 ( .A(n1781), .B(n1782), .Z(xin[199]) );
  NANDN U3700 ( .A(start), .B(xreg[199]), .Z(n1782) );
  NAND U3701 ( .A(x[199]), .B(start), .Z(n1781) );
  NAND U3702 ( .A(n1783), .B(n1784), .Z(xin[198]) );
  NANDN U3703 ( .A(start), .B(xreg[198]), .Z(n1784) );
  NAND U3704 ( .A(x[198]), .B(start), .Z(n1783) );
  NAND U3705 ( .A(n1785), .B(n1786), .Z(xin[197]) );
  NANDN U3706 ( .A(start), .B(xreg[197]), .Z(n1786) );
  NAND U3707 ( .A(x[197]), .B(start), .Z(n1785) );
  NAND U3708 ( .A(n1787), .B(n1788), .Z(xin[196]) );
  NANDN U3709 ( .A(start), .B(xreg[196]), .Z(n1788) );
  NAND U3710 ( .A(x[196]), .B(start), .Z(n1787) );
  NAND U3711 ( .A(n1789), .B(n1790), .Z(xin[195]) );
  NANDN U3712 ( .A(start), .B(xreg[195]), .Z(n1790) );
  NAND U3713 ( .A(x[195]), .B(start), .Z(n1789) );
  NAND U3714 ( .A(n1791), .B(n1792), .Z(xin[194]) );
  NANDN U3715 ( .A(start), .B(xreg[194]), .Z(n1792) );
  NAND U3716 ( .A(x[194]), .B(start), .Z(n1791) );
  NAND U3717 ( .A(n1793), .B(n1794), .Z(xin[193]) );
  NANDN U3718 ( .A(start), .B(xreg[193]), .Z(n1794) );
  NAND U3719 ( .A(x[193]), .B(start), .Z(n1793) );
  NAND U3720 ( .A(n1795), .B(n1796), .Z(xin[192]) );
  NANDN U3721 ( .A(start), .B(xreg[192]), .Z(n1796) );
  NAND U3722 ( .A(x[192]), .B(start), .Z(n1795) );
  NAND U3723 ( .A(n1797), .B(n1798), .Z(xin[191]) );
  NANDN U3724 ( .A(start), .B(xreg[191]), .Z(n1798) );
  NAND U3725 ( .A(x[191]), .B(start), .Z(n1797) );
  NAND U3726 ( .A(n1799), .B(n1800), .Z(xin[190]) );
  NANDN U3727 ( .A(start), .B(xreg[190]), .Z(n1800) );
  NAND U3728 ( .A(x[190]), .B(start), .Z(n1799) );
  NAND U3729 ( .A(n1801), .B(n1802), .Z(xin[18]) );
  NANDN U3730 ( .A(start), .B(xreg[18]), .Z(n1802) );
  NAND U3731 ( .A(x[18]), .B(start), .Z(n1801) );
  NAND U3732 ( .A(n1803), .B(n1804), .Z(xin[189]) );
  NANDN U3733 ( .A(start), .B(xreg[189]), .Z(n1804) );
  NAND U3734 ( .A(x[189]), .B(start), .Z(n1803) );
  NAND U3735 ( .A(n1805), .B(n1806), .Z(xin[188]) );
  NANDN U3736 ( .A(start), .B(xreg[188]), .Z(n1806) );
  NAND U3737 ( .A(x[188]), .B(start), .Z(n1805) );
  NAND U3738 ( .A(n1807), .B(n1808), .Z(xin[187]) );
  NANDN U3739 ( .A(start), .B(xreg[187]), .Z(n1808) );
  NAND U3740 ( .A(x[187]), .B(start), .Z(n1807) );
  NAND U3741 ( .A(n1809), .B(n1810), .Z(xin[186]) );
  NANDN U3742 ( .A(start), .B(xreg[186]), .Z(n1810) );
  NAND U3743 ( .A(x[186]), .B(start), .Z(n1809) );
  NAND U3744 ( .A(n1811), .B(n1812), .Z(xin[185]) );
  NANDN U3745 ( .A(start), .B(xreg[185]), .Z(n1812) );
  NAND U3746 ( .A(x[185]), .B(start), .Z(n1811) );
  NAND U3747 ( .A(n1813), .B(n1814), .Z(xin[184]) );
  NANDN U3748 ( .A(start), .B(xreg[184]), .Z(n1814) );
  NAND U3749 ( .A(x[184]), .B(start), .Z(n1813) );
  NAND U3750 ( .A(n1815), .B(n1816), .Z(xin[183]) );
  NANDN U3751 ( .A(start), .B(xreg[183]), .Z(n1816) );
  NAND U3752 ( .A(x[183]), .B(start), .Z(n1815) );
  NAND U3753 ( .A(n1817), .B(n1818), .Z(xin[182]) );
  NANDN U3754 ( .A(start), .B(xreg[182]), .Z(n1818) );
  NAND U3755 ( .A(x[182]), .B(start), .Z(n1817) );
  NAND U3756 ( .A(n1819), .B(n1820), .Z(xin[181]) );
  NANDN U3757 ( .A(start), .B(xreg[181]), .Z(n1820) );
  NAND U3758 ( .A(x[181]), .B(start), .Z(n1819) );
  NAND U3759 ( .A(n1821), .B(n1822), .Z(xin[180]) );
  NANDN U3760 ( .A(start), .B(xreg[180]), .Z(n1822) );
  NAND U3761 ( .A(x[180]), .B(start), .Z(n1821) );
  NAND U3762 ( .A(n1823), .B(n1824), .Z(xin[17]) );
  NANDN U3763 ( .A(start), .B(xreg[17]), .Z(n1824) );
  NAND U3764 ( .A(x[17]), .B(start), .Z(n1823) );
  NAND U3765 ( .A(n1825), .B(n1826), .Z(xin[179]) );
  NANDN U3766 ( .A(start), .B(xreg[179]), .Z(n1826) );
  NAND U3767 ( .A(x[179]), .B(start), .Z(n1825) );
  NAND U3768 ( .A(n1827), .B(n1828), .Z(xin[178]) );
  NANDN U3769 ( .A(start), .B(xreg[178]), .Z(n1828) );
  NAND U3770 ( .A(x[178]), .B(start), .Z(n1827) );
  NAND U3771 ( .A(n1829), .B(n1830), .Z(xin[177]) );
  NANDN U3772 ( .A(start), .B(xreg[177]), .Z(n1830) );
  NAND U3773 ( .A(x[177]), .B(start), .Z(n1829) );
  NAND U3774 ( .A(n1831), .B(n1832), .Z(xin[176]) );
  NANDN U3775 ( .A(start), .B(xreg[176]), .Z(n1832) );
  NAND U3776 ( .A(x[176]), .B(start), .Z(n1831) );
  NAND U3777 ( .A(n1833), .B(n1834), .Z(xin[175]) );
  NANDN U3778 ( .A(start), .B(xreg[175]), .Z(n1834) );
  NAND U3779 ( .A(x[175]), .B(start), .Z(n1833) );
  NAND U3780 ( .A(n1835), .B(n1836), .Z(xin[174]) );
  NANDN U3781 ( .A(start), .B(xreg[174]), .Z(n1836) );
  NAND U3782 ( .A(x[174]), .B(start), .Z(n1835) );
  NAND U3783 ( .A(n1837), .B(n1838), .Z(xin[173]) );
  NANDN U3784 ( .A(start), .B(xreg[173]), .Z(n1838) );
  NAND U3785 ( .A(x[173]), .B(start), .Z(n1837) );
  NAND U3786 ( .A(n1839), .B(n1840), .Z(xin[172]) );
  NANDN U3787 ( .A(start), .B(xreg[172]), .Z(n1840) );
  NAND U3788 ( .A(x[172]), .B(start), .Z(n1839) );
  NAND U3789 ( .A(n1841), .B(n1842), .Z(xin[171]) );
  NANDN U3790 ( .A(start), .B(xreg[171]), .Z(n1842) );
  NAND U3791 ( .A(x[171]), .B(start), .Z(n1841) );
  NAND U3792 ( .A(n1843), .B(n1844), .Z(xin[170]) );
  NANDN U3793 ( .A(start), .B(xreg[170]), .Z(n1844) );
  NAND U3794 ( .A(x[170]), .B(start), .Z(n1843) );
  NAND U3795 ( .A(n1845), .B(n1846), .Z(xin[16]) );
  NANDN U3796 ( .A(start), .B(xreg[16]), .Z(n1846) );
  NAND U3797 ( .A(x[16]), .B(start), .Z(n1845) );
  NAND U3798 ( .A(n1847), .B(n1848), .Z(xin[169]) );
  NANDN U3799 ( .A(start), .B(xreg[169]), .Z(n1848) );
  NAND U3800 ( .A(x[169]), .B(start), .Z(n1847) );
  NAND U3801 ( .A(n1849), .B(n1850), .Z(xin[168]) );
  NANDN U3802 ( .A(start), .B(xreg[168]), .Z(n1850) );
  NAND U3803 ( .A(x[168]), .B(start), .Z(n1849) );
  NAND U3804 ( .A(n1851), .B(n1852), .Z(xin[167]) );
  NANDN U3805 ( .A(start), .B(xreg[167]), .Z(n1852) );
  NAND U3806 ( .A(x[167]), .B(start), .Z(n1851) );
  NAND U3807 ( .A(n1853), .B(n1854), .Z(xin[166]) );
  NANDN U3808 ( .A(start), .B(xreg[166]), .Z(n1854) );
  NAND U3809 ( .A(x[166]), .B(start), .Z(n1853) );
  NAND U3810 ( .A(n1855), .B(n1856), .Z(xin[165]) );
  NANDN U3811 ( .A(start), .B(xreg[165]), .Z(n1856) );
  NAND U3812 ( .A(x[165]), .B(start), .Z(n1855) );
  NAND U3813 ( .A(n1857), .B(n1858), .Z(xin[164]) );
  NANDN U3814 ( .A(start), .B(xreg[164]), .Z(n1858) );
  NAND U3815 ( .A(x[164]), .B(start), .Z(n1857) );
  NAND U3816 ( .A(n1859), .B(n1860), .Z(xin[163]) );
  NANDN U3817 ( .A(start), .B(xreg[163]), .Z(n1860) );
  NAND U3818 ( .A(x[163]), .B(start), .Z(n1859) );
  NAND U3819 ( .A(n1861), .B(n1862), .Z(xin[162]) );
  NANDN U3820 ( .A(start), .B(xreg[162]), .Z(n1862) );
  NAND U3821 ( .A(x[162]), .B(start), .Z(n1861) );
  NAND U3822 ( .A(n1863), .B(n1864), .Z(xin[161]) );
  NANDN U3823 ( .A(start), .B(xreg[161]), .Z(n1864) );
  NAND U3824 ( .A(x[161]), .B(start), .Z(n1863) );
  NAND U3825 ( .A(n1865), .B(n1866), .Z(xin[160]) );
  NANDN U3826 ( .A(start), .B(xreg[160]), .Z(n1866) );
  NAND U3827 ( .A(x[160]), .B(start), .Z(n1865) );
  NAND U3828 ( .A(n1867), .B(n1868), .Z(xin[15]) );
  NANDN U3829 ( .A(start), .B(xreg[15]), .Z(n1868) );
  NAND U3830 ( .A(x[15]), .B(start), .Z(n1867) );
  NAND U3831 ( .A(n1869), .B(n1870), .Z(xin[159]) );
  NANDN U3832 ( .A(start), .B(xreg[159]), .Z(n1870) );
  NAND U3833 ( .A(x[159]), .B(start), .Z(n1869) );
  NAND U3834 ( .A(n1871), .B(n1872), .Z(xin[158]) );
  NANDN U3835 ( .A(start), .B(xreg[158]), .Z(n1872) );
  NAND U3836 ( .A(x[158]), .B(start), .Z(n1871) );
  NAND U3837 ( .A(n1873), .B(n1874), .Z(xin[157]) );
  NANDN U3838 ( .A(start), .B(xreg[157]), .Z(n1874) );
  NAND U3839 ( .A(x[157]), .B(start), .Z(n1873) );
  NAND U3840 ( .A(n1875), .B(n1876), .Z(xin[156]) );
  NANDN U3841 ( .A(start), .B(xreg[156]), .Z(n1876) );
  NAND U3842 ( .A(x[156]), .B(start), .Z(n1875) );
  NAND U3843 ( .A(n1877), .B(n1878), .Z(xin[155]) );
  NANDN U3844 ( .A(start), .B(xreg[155]), .Z(n1878) );
  NAND U3845 ( .A(x[155]), .B(start), .Z(n1877) );
  NAND U3846 ( .A(n1879), .B(n1880), .Z(xin[154]) );
  NANDN U3847 ( .A(start), .B(xreg[154]), .Z(n1880) );
  NAND U3848 ( .A(x[154]), .B(start), .Z(n1879) );
  NAND U3849 ( .A(n1881), .B(n1882), .Z(xin[153]) );
  NANDN U3850 ( .A(start), .B(xreg[153]), .Z(n1882) );
  NAND U3851 ( .A(x[153]), .B(start), .Z(n1881) );
  NAND U3852 ( .A(n1883), .B(n1884), .Z(xin[152]) );
  NANDN U3853 ( .A(start), .B(xreg[152]), .Z(n1884) );
  NAND U3854 ( .A(x[152]), .B(start), .Z(n1883) );
  NAND U3855 ( .A(n1885), .B(n1886), .Z(xin[151]) );
  NANDN U3856 ( .A(start), .B(xreg[151]), .Z(n1886) );
  NAND U3857 ( .A(x[151]), .B(start), .Z(n1885) );
  NAND U3858 ( .A(n1887), .B(n1888), .Z(xin[150]) );
  NANDN U3859 ( .A(start), .B(xreg[150]), .Z(n1888) );
  NAND U3860 ( .A(x[150]), .B(start), .Z(n1887) );
  NAND U3861 ( .A(n1889), .B(n1890), .Z(xin[14]) );
  NANDN U3862 ( .A(start), .B(xreg[14]), .Z(n1890) );
  NAND U3863 ( .A(x[14]), .B(start), .Z(n1889) );
  NAND U3864 ( .A(n1891), .B(n1892), .Z(xin[149]) );
  NANDN U3865 ( .A(start), .B(xreg[149]), .Z(n1892) );
  NAND U3866 ( .A(x[149]), .B(start), .Z(n1891) );
  NAND U3867 ( .A(n1893), .B(n1894), .Z(xin[148]) );
  NANDN U3868 ( .A(start), .B(xreg[148]), .Z(n1894) );
  NAND U3869 ( .A(x[148]), .B(start), .Z(n1893) );
  NAND U3870 ( .A(n1895), .B(n1896), .Z(xin[147]) );
  NANDN U3871 ( .A(start), .B(xreg[147]), .Z(n1896) );
  NAND U3872 ( .A(x[147]), .B(start), .Z(n1895) );
  NAND U3873 ( .A(n1897), .B(n1898), .Z(xin[146]) );
  NANDN U3874 ( .A(start), .B(xreg[146]), .Z(n1898) );
  NAND U3875 ( .A(x[146]), .B(start), .Z(n1897) );
  NAND U3876 ( .A(n1899), .B(n1900), .Z(xin[145]) );
  NANDN U3877 ( .A(start), .B(xreg[145]), .Z(n1900) );
  NAND U3878 ( .A(x[145]), .B(start), .Z(n1899) );
  NAND U3879 ( .A(n1901), .B(n1902), .Z(xin[144]) );
  NANDN U3880 ( .A(start), .B(xreg[144]), .Z(n1902) );
  NAND U3881 ( .A(x[144]), .B(start), .Z(n1901) );
  NAND U3882 ( .A(n1903), .B(n1904), .Z(xin[143]) );
  NANDN U3883 ( .A(start), .B(xreg[143]), .Z(n1904) );
  NAND U3884 ( .A(x[143]), .B(start), .Z(n1903) );
  NAND U3885 ( .A(n1905), .B(n1906), .Z(xin[142]) );
  NANDN U3886 ( .A(start), .B(xreg[142]), .Z(n1906) );
  NAND U3887 ( .A(x[142]), .B(start), .Z(n1905) );
  NAND U3888 ( .A(n1907), .B(n1908), .Z(xin[141]) );
  NANDN U3889 ( .A(start), .B(xreg[141]), .Z(n1908) );
  NAND U3890 ( .A(x[141]), .B(start), .Z(n1907) );
  NAND U3891 ( .A(n1909), .B(n1910), .Z(xin[140]) );
  NANDN U3892 ( .A(start), .B(xreg[140]), .Z(n1910) );
  NAND U3893 ( .A(x[140]), .B(start), .Z(n1909) );
  NAND U3894 ( .A(n1911), .B(n1912), .Z(xin[13]) );
  NANDN U3895 ( .A(start), .B(xreg[13]), .Z(n1912) );
  NAND U3896 ( .A(x[13]), .B(start), .Z(n1911) );
  NAND U3897 ( .A(n1913), .B(n1914), .Z(xin[139]) );
  NANDN U3898 ( .A(start), .B(xreg[139]), .Z(n1914) );
  NAND U3899 ( .A(x[139]), .B(start), .Z(n1913) );
  NAND U3900 ( .A(n1915), .B(n1916), .Z(xin[138]) );
  NANDN U3901 ( .A(start), .B(xreg[138]), .Z(n1916) );
  NAND U3902 ( .A(x[138]), .B(start), .Z(n1915) );
  NAND U3903 ( .A(n1917), .B(n1918), .Z(xin[137]) );
  NANDN U3904 ( .A(start), .B(xreg[137]), .Z(n1918) );
  NAND U3905 ( .A(x[137]), .B(start), .Z(n1917) );
  NAND U3906 ( .A(n1919), .B(n1920), .Z(xin[136]) );
  NANDN U3907 ( .A(start), .B(xreg[136]), .Z(n1920) );
  NAND U3908 ( .A(x[136]), .B(start), .Z(n1919) );
  NAND U3909 ( .A(n1921), .B(n1922), .Z(xin[135]) );
  NANDN U3910 ( .A(start), .B(xreg[135]), .Z(n1922) );
  NAND U3911 ( .A(x[135]), .B(start), .Z(n1921) );
  NAND U3912 ( .A(n1923), .B(n1924), .Z(xin[134]) );
  NANDN U3913 ( .A(start), .B(xreg[134]), .Z(n1924) );
  NAND U3914 ( .A(x[134]), .B(start), .Z(n1923) );
  NAND U3915 ( .A(n1925), .B(n1926), .Z(xin[133]) );
  NANDN U3916 ( .A(start), .B(xreg[133]), .Z(n1926) );
  NAND U3917 ( .A(x[133]), .B(start), .Z(n1925) );
  NAND U3918 ( .A(n1927), .B(n1928), .Z(xin[132]) );
  NANDN U3919 ( .A(start), .B(xreg[132]), .Z(n1928) );
  NAND U3920 ( .A(x[132]), .B(start), .Z(n1927) );
  NAND U3921 ( .A(n1929), .B(n1930), .Z(xin[131]) );
  NANDN U3922 ( .A(start), .B(xreg[131]), .Z(n1930) );
  NAND U3923 ( .A(x[131]), .B(start), .Z(n1929) );
  NAND U3924 ( .A(n1931), .B(n1932), .Z(xin[130]) );
  NANDN U3925 ( .A(start), .B(xreg[130]), .Z(n1932) );
  NAND U3926 ( .A(x[130]), .B(start), .Z(n1931) );
  NAND U3927 ( .A(n1933), .B(n1934), .Z(xin[12]) );
  NANDN U3928 ( .A(start), .B(xreg[12]), .Z(n1934) );
  NAND U3929 ( .A(x[12]), .B(start), .Z(n1933) );
  NAND U3930 ( .A(n1935), .B(n1936), .Z(xin[129]) );
  NANDN U3931 ( .A(start), .B(xreg[129]), .Z(n1936) );
  NAND U3932 ( .A(x[129]), .B(start), .Z(n1935) );
  NAND U3933 ( .A(n1937), .B(n1938), .Z(xin[128]) );
  NANDN U3934 ( .A(start), .B(xreg[128]), .Z(n1938) );
  NAND U3935 ( .A(x[128]), .B(start), .Z(n1937) );
  NAND U3936 ( .A(n1939), .B(n1940), .Z(xin[127]) );
  NANDN U3937 ( .A(start), .B(xreg[127]), .Z(n1940) );
  NAND U3938 ( .A(x[127]), .B(start), .Z(n1939) );
  NAND U3939 ( .A(n1941), .B(n1942), .Z(xin[126]) );
  NANDN U3940 ( .A(start), .B(xreg[126]), .Z(n1942) );
  NAND U3941 ( .A(x[126]), .B(start), .Z(n1941) );
  NAND U3942 ( .A(n1943), .B(n1944), .Z(xin[125]) );
  NANDN U3943 ( .A(start), .B(xreg[125]), .Z(n1944) );
  NAND U3944 ( .A(x[125]), .B(start), .Z(n1943) );
  NAND U3945 ( .A(n1945), .B(n1946), .Z(xin[124]) );
  NANDN U3946 ( .A(start), .B(xreg[124]), .Z(n1946) );
  NAND U3947 ( .A(x[124]), .B(start), .Z(n1945) );
  NAND U3948 ( .A(n1947), .B(n1948), .Z(xin[123]) );
  NANDN U3949 ( .A(start), .B(xreg[123]), .Z(n1948) );
  NAND U3950 ( .A(x[123]), .B(start), .Z(n1947) );
  NAND U3951 ( .A(n1949), .B(n1950), .Z(xin[122]) );
  NANDN U3952 ( .A(start), .B(xreg[122]), .Z(n1950) );
  NAND U3953 ( .A(x[122]), .B(start), .Z(n1949) );
  NAND U3954 ( .A(n1951), .B(n1952), .Z(xin[121]) );
  NANDN U3955 ( .A(start), .B(xreg[121]), .Z(n1952) );
  NAND U3956 ( .A(x[121]), .B(start), .Z(n1951) );
  NAND U3957 ( .A(n1953), .B(n1954), .Z(xin[120]) );
  NANDN U3958 ( .A(start), .B(xreg[120]), .Z(n1954) );
  NAND U3959 ( .A(x[120]), .B(start), .Z(n1953) );
  NAND U3960 ( .A(n1955), .B(n1956), .Z(xin[11]) );
  NANDN U3961 ( .A(start), .B(xreg[11]), .Z(n1956) );
  NAND U3962 ( .A(x[11]), .B(start), .Z(n1955) );
  NAND U3963 ( .A(n1957), .B(n1958), .Z(xin[119]) );
  NANDN U3964 ( .A(start), .B(xreg[119]), .Z(n1958) );
  NAND U3965 ( .A(x[119]), .B(start), .Z(n1957) );
  NAND U3966 ( .A(n1959), .B(n1960), .Z(xin[118]) );
  NANDN U3967 ( .A(start), .B(xreg[118]), .Z(n1960) );
  NAND U3968 ( .A(x[118]), .B(start), .Z(n1959) );
  NAND U3969 ( .A(n1961), .B(n1962), .Z(xin[117]) );
  NANDN U3970 ( .A(start), .B(xreg[117]), .Z(n1962) );
  NAND U3971 ( .A(x[117]), .B(start), .Z(n1961) );
  NAND U3972 ( .A(n1963), .B(n1964), .Z(xin[116]) );
  NANDN U3973 ( .A(start), .B(xreg[116]), .Z(n1964) );
  NAND U3974 ( .A(x[116]), .B(start), .Z(n1963) );
  NAND U3975 ( .A(n1965), .B(n1966), .Z(xin[115]) );
  NANDN U3976 ( .A(start), .B(xreg[115]), .Z(n1966) );
  NAND U3977 ( .A(x[115]), .B(start), .Z(n1965) );
  NAND U3978 ( .A(n1967), .B(n1968), .Z(xin[114]) );
  NANDN U3979 ( .A(start), .B(xreg[114]), .Z(n1968) );
  NAND U3980 ( .A(x[114]), .B(start), .Z(n1967) );
  NAND U3981 ( .A(n1969), .B(n1970), .Z(xin[113]) );
  NANDN U3982 ( .A(start), .B(xreg[113]), .Z(n1970) );
  NAND U3983 ( .A(x[113]), .B(start), .Z(n1969) );
  NAND U3984 ( .A(n1971), .B(n1972), .Z(xin[112]) );
  NANDN U3985 ( .A(start), .B(xreg[112]), .Z(n1972) );
  NAND U3986 ( .A(x[112]), .B(start), .Z(n1971) );
  NAND U3987 ( .A(n1973), .B(n1974), .Z(xin[111]) );
  NANDN U3988 ( .A(start), .B(xreg[111]), .Z(n1974) );
  NAND U3989 ( .A(x[111]), .B(start), .Z(n1973) );
  NAND U3990 ( .A(n1975), .B(n1976), .Z(xin[110]) );
  NANDN U3991 ( .A(start), .B(xreg[110]), .Z(n1976) );
  NAND U3992 ( .A(x[110]), .B(start), .Z(n1975) );
  NAND U3993 ( .A(n1977), .B(n1978), .Z(xin[10]) );
  NANDN U3994 ( .A(start), .B(xreg[10]), .Z(n1978) );
  NAND U3995 ( .A(x[10]), .B(start), .Z(n1977) );
  NAND U3996 ( .A(n1979), .B(n1980), .Z(xin[109]) );
  NANDN U3997 ( .A(start), .B(xreg[109]), .Z(n1980) );
  NAND U3998 ( .A(x[109]), .B(start), .Z(n1979) );
  NAND U3999 ( .A(n1981), .B(n1982), .Z(xin[108]) );
  NANDN U4000 ( .A(start), .B(xreg[108]), .Z(n1982) );
  NAND U4001 ( .A(x[108]), .B(start), .Z(n1981) );
  NAND U4002 ( .A(n1983), .B(n1984), .Z(xin[107]) );
  NANDN U4003 ( .A(start), .B(xreg[107]), .Z(n1984) );
  NAND U4004 ( .A(x[107]), .B(start), .Z(n1983) );
  NAND U4005 ( .A(n1985), .B(n1986), .Z(xin[106]) );
  NANDN U4006 ( .A(start), .B(xreg[106]), .Z(n1986) );
  NAND U4007 ( .A(x[106]), .B(start), .Z(n1985) );
  NAND U4008 ( .A(n1987), .B(n1988), .Z(xin[105]) );
  NANDN U4009 ( .A(start), .B(xreg[105]), .Z(n1988) );
  NAND U4010 ( .A(x[105]), .B(start), .Z(n1987) );
  NAND U4011 ( .A(n1989), .B(n1990), .Z(xin[104]) );
  NANDN U4012 ( .A(start), .B(xreg[104]), .Z(n1990) );
  NAND U4013 ( .A(x[104]), .B(start), .Z(n1989) );
  NAND U4014 ( .A(n1991), .B(n1992), .Z(xin[103]) );
  NANDN U4015 ( .A(start), .B(xreg[103]), .Z(n1992) );
  NAND U4016 ( .A(x[103]), .B(start), .Z(n1991) );
  NAND U4017 ( .A(n1993), .B(n1994), .Z(xin[102]) );
  NANDN U4018 ( .A(start), .B(xreg[102]), .Z(n1994) );
  NAND U4019 ( .A(x[102]), .B(start), .Z(n1993) );
  NAND U4020 ( .A(n1995), .B(n1996), .Z(xin[1023]) );
  NANDN U4021 ( .A(start), .B(xreg[1023]), .Z(n1996) );
  NAND U4022 ( .A(x[1023]), .B(start), .Z(n1995) );
  NAND U4023 ( .A(n1997), .B(n1998), .Z(xin[1022]) );
  NANDN U4024 ( .A(start), .B(xreg[1022]), .Z(n1998) );
  NAND U4025 ( .A(x[1022]), .B(start), .Z(n1997) );
  NAND U4026 ( .A(n1999), .B(n2000), .Z(xin[1021]) );
  NANDN U4027 ( .A(start), .B(xreg[1021]), .Z(n2000) );
  NAND U4028 ( .A(x[1021]), .B(start), .Z(n1999) );
  NAND U4029 ( .A(n2001), .B(n2002), .Z(xin[1020]) );
  NANDN U4030 ( .A(start), .B(xreg[1020]), .Z(n2002) );
  NAND U4031 ( .A(x[1020]), .B(start), .Z(n2001) );
  NAND U4032 ( .A(n2003), .B(n2004), .Z(xin[101]) );
  NANDN U4033 ( .A(start), .B(xreg[101]), .Z(n2004) );
  NAND U4034 ( .A(x[101]), .B(start), .Z(n2003) );
  NAND U4035 ( .A(n2005), .B(n2006), .Z(xin[1019]) );
  NANDN U4036 ( .A(start), .B(xreg[1019]), .Z(n2006) );
  NAND U4037 ( .A(x[1019]), .B(start), .Z(n2005) );
  NAND U4038 ( .A(n2007), .B(n2008), .Z(xin[1018]) );
  NANDN U4039 ( .A(start), .B(xreg[1018]), .Z(n2008) );
  NAND U4040 ( .A(x[1018]), .B(start), .Z(n2007) );
  NAND U4041 ( .A(n2009), .B(n2010), .Z(xin[1017]) );
  NANDN U4042 ( .A(start), .B(xreg[1017]), .Z(n2010) );
  NAND U4043 ( .A(x[1017]), .B(start), .Z(n2009) );
  NAND U4044 ( .A(n2011), .B(n2012), .Z(xin[1016]) );
  NANDN U4045 ( .A(start), .B(xreg[1016]), .Z(n2012) );
  NAND U4046 ( .A(x[1016]), .B(start), .Z(n2011) );
  NAND U4047 ( .A(n2013), .B(n2014), .Z(xin[1015]) );
  NANDN U4048 ( .A(start), .B(xreg[1015]), .Z(n2014) );
  NAND U4049 ( .A(x[1015]), .B(start), .Z(n2013) );
  NAND U4050 ( .A(n2015), .B(n2016), .Z(xin[1014]) );
  NANDN U4051 ( .A(start), .B(xreg[1014]), .Z(n2016) );
  NAND U4052 ( .A(x[1014]), .B(start), .Z(n2015) );
  NAND U4053 ( .A(n2017), .B(n2018), .Z(xin[1013]) );
  NANDN U4054 ( .A(start), .B(xreg[1013]), .Z(n2018) );
  NAND U4055 ( .A(x[1013]), .B(start), .Z(n2017) );
  NAND U4056 ( .A(n2019), .B(n2020), .Z(xin[1012]) );
  NANDN U4057 ( .A(start), .B(xreg[1012]), .Z(n2020) );
  NAND U4058 ( .A(x[1012]), .B(start), .Z(n2019) );
  NAND U4059 ( .A(n2021), .B(n2022), .Z(xin[1011]) );
  NANDN U4060 ( .A(start), .B(xreg[1011]), .Z(n2022) );
  NAND U4061 ( .A(x[1011]), .B(start), .Z(n2021) );
  NAND U4062 ( .A(n2023), .B(n2024), .Z(xin[1010]) );
  NANDN U4063 ( .A(start), .B(xreg[1010]), .Z(n2024) );
  NAND U4064 ( .A(x[1010]), .B(start), .Z(n2023) );
  NAND U4065 ( .A(n2025), .B(n2026), .Z(xin[100]) );
  NANDN U4066 ( .A(start), .B(xreg[100]), .Z(n2026) );
  NAND U4067 ( .A(x[100]), .B(start), .Z(n2025) );
  NAND U4068 ( .A(n2027), .B(n2028), .Z(xin[1009]) );
  NANDN U4069 ( .A(start), .B(xreg[1009]), .Z(n2028) );
  NAND U4070 ( .A(x[1009]), .B(start), .Z(n2027) );
  NAND U4071 ( .A(n2029), .B(n2030), .Z(xin[1008]) );
  NANDN U4072 ( .A(start), .B(xreg[1008]), .Z(n2030) );
  NAND U4073 ( .A(x[1008]), .B(start), .Z(n2029) );
  NAND U4074 ( .A(n2031), .B(n2032), .Z(xin[1007]) );
  NANDN U4075 ( .A(start), .B(xreg[1007]), .Z(n2032) );
  NAND U4076 ( .A(x[1007]), .B(start), .Z(n2031) );
  NAND U4077 ( .A(n2033), .B(n2034), .Z(xin[1006]) );
  NANDN U4078 ( .A(start), .B(xreg[1006]), .Z(n2034) );
  NAND U4079 ( .A(x[1006]), .B(start), .Z(n2033) );
  NAND U4080 ( .A(n2035), .B(n2036), .Z(xin[1005]) );
  NANDN U4081 ( .A(start), .B(xreg[1005]), .Z(n2036) );
  NAND U4082 ( .A(x[1005]), .B(start), .Z(n2035) );
  NAND U4083 ( .A(n2037), .B(n2038), .Z(xin[1004]) );
  NANDN U4084 ( .A(start), .B(xreg[1004]), .Z(n2038) );
  NAND U4085 ( .A(x[1004]), .B(start), .Z(n2037) );
  NAND U4086 ( .A(n2039), .B(n2040), .Z(xin[1003]) );
  NANDN U4087 ( .A(start), .B(xreg[1003]), .Z(n2040) );
  NAND U4088 ( .A(x[1003]), .B(start), .Z(n2039) );
  NAND U4089 ( .A(n2041), .B(n2042), .Z(xin[1002]) );
  NANDN U4090 ( .A(start), .B(xreg[1002]), .Z(n2042) );
  NAND U4091 ( .A(x[1002]), .B(start), .Z(n2041) );
  NAND U4092 ( .A(n2043), .B(n2044), .Z(xin[1001]) );
  NANDN U4093 ( .A(start), .B(xreg[1001]), .Z(n2044) );
  NAND U4094 ( .A(x[1001]), .B(start), .Z(n2043) );
  NAND U4095 ( .A(n2045), .B(n2046), .Z(xin[1000]) );
  NANDN U4096 ( .A(start), .B(xreg[1000]), .Z(n2046) );
  NAND U4097 ( .A(x[1000]), .B(start), .Z(n2045) );
  AND U4098 ( .A(x[0]), .B(start), .Z(n2047) );
endmodule


module modexp_2N_NN_N1024_CC2097152 ( clk, rst, m, e, n, c );
  input [1023:0] m;
  input [1023:0] e;
  input [1023:0] n;
  output [1023:0] c;
  input clk, rst;
  wire   init, mul_pow, first_one, n13329, n13330, n13331, n13332, n13333,
         n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341,
         n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349,
         n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357,
         n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365,
         n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373,
         n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381,
         n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389,
         n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397,
         n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405,
         n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413,
         n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421,
         n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429,
         n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437,
         n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445,
         n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453,
         n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461,
         n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469,
         n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477,
         n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485,
         n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493,
         n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501,
         n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509,
         n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517,
         n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525,
         n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533,
         n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541,
         n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549,
         n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557,
         n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565,
         n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573,
         n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581,
         n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589,
         n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597,
         n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605,
         n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613,
         n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621,
         n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629,
         n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637,
         n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645,
         n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653,
         n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661,
         n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669,
         n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677,
         n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685,
         n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693,
         n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701,
         n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709,
         n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717,
         n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725,
         n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733,
         n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741,
         n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749,
         n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757,
         n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765,
         n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773,
         n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781,
         n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789,
         n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797,
         n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805,
         n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813,
         n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821,
         n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829,
         n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837,
         n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845,
         n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853,
         n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861,
         n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869,
         n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877,
         n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885,
         n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893,
         n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901,
         n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909,
         n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917,
         n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925,
         n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933,
         n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941,
         n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949,
         n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957,
         n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965,
         n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973,
         n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981,
         n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989,
         n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997,
         n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005,
         n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013,
         n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021,
         n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029,
         n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037,
         n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045,
         n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053,
         n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061,
         n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069,
         n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077,
         n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085,
         n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093,
         n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101,
         n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109,
         n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117,
         n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125,
         n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133,
         n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141,
         n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149,
         n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157,
         n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165,
         n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
         n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181,
         n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189,
         n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197,
         n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205,
         n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213,
         n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221,
         n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229,
         n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237,
         n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245,
         n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253,
         n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261,
         n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269,
         n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277,
         n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285,
         n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293,
         n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301,
         n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309,
         n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317,
         n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325,
         n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333,
         n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341,
         n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349,
         n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357,
         n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365,
         n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373,
         n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381,
         n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389,
         n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397,
         n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405,
         n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413,
         n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421,
         n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429,
         n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437,
         n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445,
         n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453,
         n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461,
         n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469,
         n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477,
         n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485,
         n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493,
         n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501,
         n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509,
         n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517,
         n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525,
         n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533,
         n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541,
         n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549,
         n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557,
         n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565,
         n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573,
         n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581,
         n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589,
         n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597,
         n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605,
         n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613,
         n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621,
         n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629,
         n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637,
         n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645,
         n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653,
         n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661,
         n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669,
         n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677,
         n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685,
         n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693,
         n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701,
         n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709,
         n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717,
         n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725,
         n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733,
         n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741,
         n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749,
         n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757,
         n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765,
         n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773,
         n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781,
         n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789,
         n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797,
         n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805,
         n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813,
         n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821,
         n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829,
         n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837,
         n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845,
         n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853,
         n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861,
         n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869,
         n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877,
         n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885,
         n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893,
         n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901,
         n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909,
         n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917,
         n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925,
         n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933,
         n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941,
         n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949,
         n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957,
         n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965,
         n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973,
         n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981,
         n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989,
         n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997,
         n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005,
         n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013,
         n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021,
         n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029,
         n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037,
         n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045,
         n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053,
         n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061,
         n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069,
         n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077,
         n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085,
         n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093,
         n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101,
         n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109,
         n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117,
         n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125,
         n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133,
         n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141,
         n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149,
         n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157,
         n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165,
         n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173,
         n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181,
         n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189,
         n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197,
         n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205,
         n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213,
         n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221,
         n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229,
         n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237,
         n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245,
         n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253,
         n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261,
         n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269,
         n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277,
         n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285,
         n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293,
         n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301,
         n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309,
         n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317,
         n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325,
         n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333,
         n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341,
         n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349,
         n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357,
         n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365,
         n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373,
         n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381,
         n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389,
         n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397,
         n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405,
         n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413,
         n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421,
         n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429,
         n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437,
         n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445,
         n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453,
         n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461,
         n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469,
         n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477,
         n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485,
         n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493,
         n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501,
         n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509,
         n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517,
         n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525,
         n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533,
         n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541,
         n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549,
         n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557,
         n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565,
         n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573,
         n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581,
         n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589,
         n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597,
         n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605,
         n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613,
         n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621,
         n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629,
         n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637,
         n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645,
         n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653,
         n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661,
         n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669,
         n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677,
         n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685,
         n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693,
         n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701,
         n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709,
         n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717,
         n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725,
         n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733,
         n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741,
         n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749,
         n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757,
         n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765,
         n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773,
         n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781,
         n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789,
         n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797,
         n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805,
         n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813,
         n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821,
         n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829,
         n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837,
         n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845,
         n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853,
         n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861,
         n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869,
         n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877,
         n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885,
         n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893,
         n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901,
         n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909,
         n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917,
         n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925,
         n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933,
         n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941,
         n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949,
         n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957,
         n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965,
         n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973,
         n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981,
         n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989,
         n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997,
         n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005,
         n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013,
         n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021,
         n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029,
         n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037,
         n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045,
         n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053,
         n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061,
         n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069,
         n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077,
         n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085,
         n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093,
         n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101,
         n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109,
         n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117,
         n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125,
         n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133,
         n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141,
         n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149,
         n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157,
         n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165,
         n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173,
         n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181,
         n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189,
         n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197,
         n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205,
         n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213,
         n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221,
         n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229,
         n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237,
         n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245,
         n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253,
         n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261,
         n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269,
         n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277,
         n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285,
         n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293,
         n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301,
         n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309,
         n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317,
         n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325,
         n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333,
         n16334, n16335, n16336, n16337, n16338, n16339, n16340, n16341,
         n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349,
         n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357,
         n16358, n16359, n16360, n16361, n16362, n16363, n16364, n16365,
         n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373,
         n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381,
         n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389,
         n16390, n16391, n16392, n16393, n16394, n16395, n16396, n16397,
         n16398, n16399, n16400, n16401, n16402, n16403, n16404, n16405,
         n16406, n16407, n16408, n16409, n16410, n16411, n16412, n16413,
         n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16421,
         n16422, n16423, n16424, n16425, n16426, n16427, n16428, n16429,
         n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437,
         n16438, n16439, n16440, n16441, n16442, n16443, n16444, n16445,
         n16446, n16447, n16448, n16449, n16450, n16451, n16452, n16453,
         n16454, n16455, n16456, n16457, n16458, n16459, n16460, n16461,
         n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469,
         n16470, n16471, n16472, n16473, n16474, n16475, n16476, n16477,
         n16478, n16479, n16480, n16481, n16482, n16483, n16484, n16485,
         n16486, n16487, n16488, n16489, n16490, n16491, n16492, n16493,
         n16494, n16495, n16496, n16497, n16498, n16499, n16500, n16501,
         n16502, n16503, n16504, n16505, n16506, n16507, n16508, n16509,
         n16510, n16511, n16512, n16513, n16514, n16515, n16516, n16517,
         n16518, n16519, n16520, n16521, n16522, n16523, n16524, n16525,
         n16526, n16527, n16528, n16529, n16530, n16531, n16532, n16533,
         n16534, n16535, n16536, n16537, n16538, n16539, n16540, n16541,
         n16542, n16543, n16544, n16545, n16546, n16547, n16548, n16549,
         n16550, n16551, n16552, n16553, n16554, n16555, n16556, n16557,
         n16558, n16559, n16560, n16561, n16562, n16563, n16564, n16565,
         n16566, n16567, n16568, n16569, n16570, n16571, n16572, n16573,
         n16574, n16575, n16576, n16577, n16578, n16579, n16580, n16581,
         n16582, n16583, n16584, n16585, n16586, n16587, n16588, n16589,
         n16590, n16591, n16592, n16593, n16594, n16595, n16596, n16597,
         n16598, n16599, n16600, n16601, n16602, n16603, n16604, n16605,
         n16606, n16607, n16608, n16609, n16610, n16611, n16612, n16613,
         n16614, n16615, n16616, n16617, n16618, n16619, n16620, n16621,
         n16622, n16623, n16624, n16625, n16626, n16627, n16628, n16629,
         n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16637,
         n16638, n16639, n16640, n16641, n16642, n16643, n16644, n16645,
         n16646, n16647, n16648, n16649, n16650, n16651, n16652, n16653,
         n16654, n16655, n16656, n16657, n16658, n16659, n16660, n16661,
         n16662, n16663, n16664, n16665, n16666, n16667, n16668, n16669,
         n16670, n16671, n16672, n16673, n16674, n16675, n16676, n16677,
         n16678, n16679, n16680, n16681, n16682, n16683, n16684, n16685,
         n16686, n16687, n16688, n16689, n16690, n16691, n16692, n16693,
         n16694, n16695, n16696, n16697, n16698, n16699, n16700, n16701,
         n16702, n16703, n16704, n16705, n16706, n16707, n16708, n16709,
         n16710, n16711, n16712, n16713, n16714, n16715, n16716, n16717,
         n16718, n16719, n16720, n16721, n16722, n16723, n16724, n16725,
         n16726, n16727, n16728, n16729, n16730, n16731, n16732, n16733,
         n16734, n16735, n16736, n16737, n16738, n16739, n16740, n16741,
         n16742, n16743, n16744, n16745, n16746, n16747, n16748, n16749,
         n16750, n16751, n16752, n16753, n16754, n16755, n16756, n16757,
         n16758, n16759, n16760, n16761, n16762, n16763, n16764, n16765,
         n16766, n16767, n16768, n16769, n16770, n16771, n16772, n16773,
         n16774, n16775, n16776, n16777, n16778, n16779, n16780, n16781,
         n16782, n16783, n16784, n16785, n16786, n16787, n16788, n16789,
         n16790, n16791, n16792, n16793, n16794, n16795, n16796, n16797,
         n16798, n16799, n16800, n16801, n16802, n16803, n16804, n16805,
         n16806, n16807, n16808, n16809, n16810, n16811, n16812, n16813,
         n16814, n16815, n16816, n16817, n16818, n16819, n16820, n16821,
         n16822, n16823, n16824, n16825, n16826, n16827, n16828, n16829,
         n16830, n16831, n16832, n16833, n16834, n16835, n16836, n16837,
         n16838, n16839, n16840, n16841, n16842, n16843, n16844, n16845,
         n16846, n16847, n16848, n16849, n16850, n16851, n16852, n16853,
         n16854, n16855, n16856, n16857, n16858, n16859, n16860, n16861,
         n16862, n16863, n16864, n16865, n16866, n16867, n16868, n16869,
         n16870, n16871, n16872, n16873, n16874, n16875, n16876, n16877,
         n16878, n16879, n16880, n16881, n16882, n16883, n16884, n16885,
         n16886, n16887, n16888, n16889, n16890, n16891, n16892, n16893,
         n16894, n16895, n16896, n16897, n16898, n16899, n16900, n16901,
         n16902, n16903, n16904, n16905, n16906, n16907, n16908, n16909,
         n16910, n16911, n16912, n16913, n16914, n16915, n16916, n16917,
         n16918, n16919, n16920, n16921, n16922, n16923, n16924, n16925,
         n16926, n16927, n16928, n16929, n16930, n16931, n16932, n16933,
         n16934, n16935, n16936, n16937, n16938, n16939, n16940, n16941,
         n16942, n16943, n16944, n16945, n16946, n16947, n16948, n16949,
         n16950, n16951, n16952, n16953, n16954, n16955, n16956, n16957,
         n16958, n16959, n16960, n16961, n16962, n16963, n16964, n16965,
         n16966, n16967, n16968, n16969, n16970, n16971, n16972, n16973,
         n16974, n16975, n16976, n16977, n16978, n16979, n16980, n16981,
         n16982, n16983, n16984, n16985, n16986, n16987, n16988, n16989,
         n16990, n16991, n16992, n16993, n16994, n16995, n16996, n16997,
         n16998, n16999, n17000, n17001, n17002, n17003, n17004, n17005,
         n17006, n17007, n17008, n17009, n17010, n17011, n17012, n17013,
         n17014, n17015, n17016, n17017, n17018, n17019, n17020, n17021,
         n17022, n17023, n17024, n17025, n17026, n17027, n17028, n17029,
         n17030, n17031, n17032, n17033, n17034, n17035, n17036, n17037,
         n17038, n17039, n17040, n17041, n17042, n17043, n17044, n17045,
         n17046, n17047, n17048, n17049, n17050, n17051, n17052, n17053,
         n17054, n17055, n17056, n17057, n17058, n17059, n17060, n17061,
         n17062, n17063, n17064, n17065, n17066, n17067, n17068, n17069,
         n17070, n17071, n17072, n17073, n17074, n17075, n17076, n17077,
         n17078, n17079, n17080, n17081, n17082, n17083, n17084, n17085,
         n17086, n17087, n17088, n17089, n17090, n17091, n17092, n17093,
         n17094, n17095, n17096, n17097, n17098, n17099, n17100, n17101,
         n17102, n17103, n17104, n17105, n17106, n17107, n17108, n17109,
         n17110, n17111, n17112, n17113, n17114, n17115, n17116, n17117,
         n17118, n17119, n17120, n17121, n17122, n17123, n17124, n17125,
         n17126, n17127, n17128, n17129, n17130, n17131, n17132, n17133,
         n17134, n17135, n17136, n17137, n17138, n17139, n17140, n17141,
         n17142, n17143, n17144, n17145, n17146, n17147, n17148, n17149,
         n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17157,
         n17158, n17159, n17160, n17161, n17162, n17163, n17164, n17165,
         n17166, n17167, n17168, n17169, n17170, n17171, n17172, n17173,
         n17174, n17175, n17176, n17177, n17178, n17179, n17180, n17181,
         n17182, n17183, n17184, n17185, n17186, n17187, n17188, n17189,
         n17190, n17191, n17192, n17193, n17194, n17195, n17196, n17197,
         n17198, n17199, n17200, n17201, n17202, n17203, n17204, n17205,
         n17206, n17207, n17208, n17209, n17210, n17211, n17212, n17213,
         n17214, n17215, n17216, n17217, n17218, n17219, n17220, n17221,
         n17222, n17223, n17224, n17225, n17226, n17227, n17228, n17229,
         n17230, n17231, n17232, n17233, n17234, n17235, n17236, n17237,
         n17238, n17239, n17240, n17241, n17242, n17243, n17244, n17245,
         n17246, n17247, n17248, n17249, n17250, n17251, n17252, n17253,
         n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261,
         n17262, n17263, n17264, n17265, n17266, n17267, n17268, n17269,
         n17270, n17271, n17272, n17273, n17274, n17275, n17276, n17277,
         n17278, n17279, n17280, n17281, n17282, n17283, n17284, n17285,
         n17286, n17287, n17288, n17289, n17290, n17291, n17292, n17293,
         n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17301,
         n17302, n17303, n17304, n17305, n17306, n17307, n17308, n17309,
         n17310, n17311, n17312, n17313, n17314, n17315, n17316, n17317,
         n17318, n17319, n17320, n17321, n17322, n17323, n17324, n17325,
         n17326, n17327, n17328, n17329, n17330, n17331, n17332, n17333,
         n17334, n17335, n17336, n17337, n17338, n17339, n17340, n17341,
         n17342, n17343, n17344, n17345, n17346, n17347, n17348, n17349,
         n17350, n17351, n17352, n17353, n17354, n17355, n17356, n17357,
         n17358, n17359, n17360, n17361, n17362, n17363, n17364, n17365,
         n17366, n17367, n17368, n17369, n17370, n17371, n17372, n17373,
         n17374, n17375, n17376, n17377, n17378, n17379, n17380, n17381,
         n17382, n17383, n17384, n17385, n17386, n17387, n17388, n17389,
         n17390, n17391, n17392, n17393, n17394, n17395, n17396, n17397,
         n17398, n17399, n17400, n17401, n17402, n17403, n17404, n17405,
         n17406, n17407, n17408, n17409, n17410, n17411, n17412, n17413,
         n17414, n17415, n17416, n17417, n17418, n17419, n17420, n17421,
         n17422, n17423, n17424, n17425, n17426, n17427, n17428, n17429,
         n17430, n17431, n17432, n17433, n17434, n17435, n17436, n17437,
         n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445,
         n17446, n17447, n17448, n17449, n17450, n17451, n17452, n17453,
         n17454, n17455, n17456, n17457, n17458, n17459, n17460, n17461,
         n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469,
         n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477,
         n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485,
         n17486, n17487, n17488, n17489, n17490, n17491, n17492, n17493,
         n17494, n17495, n17496, n17497, n17498, n17499, n17500, n17501,
         n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509,
         n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517,
         n17518, n17519, n17520, n17521, n17522, n17523, n17524, n17525,
         n17526, n17527, n17528, n17529, n17530, n17531, n17532, n17533,
         n17534, n17535, n17536, n17537, n17538, n17539, n17540, n17541,
         n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549,
         n17550, n17551, n17552, n17553, n17554, n17555, n17556, n17557,
         n17558, n17559, n17560, n17561, n17562, n17563, n17564, n17565,
         n17566, n17567, n17568, n17569, n17570, n17571, n17572, n17573,
         n17574, n17575, n17576, n17577, n17578, n17579, n17580, n17581,
         n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589,
         n17590, n17591, n17592, n17593, n17594, n17595, n17596, n17597,
         n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605,
         n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613,
         n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621,
         n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17629,
         n17630, n17631, n17632, n17633, n17634, n17635, n17636, n17637,
         n17638, n17639, n17640, n17641, n17642, n17643, n17644, n17645,
         n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653,
         n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661,
         n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669,
         n17670, n17671, n17672, n17673, n17674, n17675, n17676, n17677,
         n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685,
         n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693,
         n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701,
         n17702, n17703, n17704, n17705, n17706, n17707, n17708, n17709,
         n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17717,
         n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725,
         n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733,
         n17734, n17735, n17736, n17737, n17738, n17739, n17740, n17741,
         n17742, n17743, n17744, n17745, n17746, n17747, n17748, n17749,
         n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757,
         n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765,
         n17766, n17767, n17768, n17769, n17770, n17771, n17772, n17773,
         n17774, n17775, n17776, n17777, n17778, n17779, n17780, n17781,
         n17782, n17783, n17784, n17785, n17786, n17787, n17788, n17789,
         n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797,
         n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805,
         n17806, n17807, n17808, n17809, n17810, n17811, n17812, n17813,
         n17814, n17815, n17816, n17817, n17818, n17819, n17820, n17821,
         n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829,
         n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17837,
         n17838, n17839, n17840, n17841, n17842, n17843, n17844, n17845,
         n17846, n17847, n17848, n17849, n17850, n17851, n17852, n17853,
         n17854, n17855, n17856, n17857, n17858, n17859, n17860, n17861,
         n17862, n17863, n17864, n17865, n17866, n17867, n17868, n17869,
         n17870, n17871, n17872, n17873, n17874, n17875, n17876, n17877,
         n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17885,
         n17886, n17887, n17888, n17889, n17890, n17891, n17892, n17893,
         n17894, n17895, n17896, n17897, n17898, n17899, n17900, n17901,
         n17902, n17903, n17904, n17905, n17906, n17907, n17908, n17909,
         n17910, n17911, n17912, n17913, n17914, n17915, n17916, n17917,
         n17918, n17919, n17920, n17921, n17922, n17923, n17924, n17925,
         n17926, n17927, n17928, n17929, n17930, n17931, n17932, n17933,
         n17934, n17935, n17936, n17937, n17938, n17939, n17940, n17941,
         n17942, n17943, n17944, n17945, n17946, n17947, n17948, n17949,
         n17950, n17951, n17952, n17953, n17954, n17955, n17956, n17957,
         n17958, n17959, n17960, n17961, n17962, n17963, n17964, n17965,
         n17966, n17967, n17968, n17969, n17970, n17971, n17972, n17973,
         n17974, n17975, n17976, n17977, n17978, n17979, n17980, n17981,
         n17982, n17983, n17984, n17985, n17986, n17987, n17988, n17989,
         n17990, n17991, n17992, n17993, n17994, n17995, n17996, n17997,
         n17998, n17999, n18000, n18001, n18002, n18003, n18004, n18005,
         n18006, n18007, n18008, n18009, n18010, n18011, n18012, n18013,
         n18014, n18015, n18016, n18017, n18018, n18019, n18020, n18021,
         n18022, n18023, n18024, n18025, n18026, n18027, n18028, n18029,
         n18030, n18031, n18032, n18033, n18034, n18035, n18036, n18037,
         n18038, n18039, n18040, n18041, n18042, n18043, n18044, n18045,
         n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053,
         n18054, n18055, n18056, n18057, n18058, n18059, n18060, n18061,
         n18062, n18063, n18064, n18065, n18066, n18067, n18068, n18069,
         n18070, n18071, n18072, n18073, n18074, n18075, n18076, n18077,
         n18078, n18079, n18080, n18081, n18082, n18083, n18084, n18085,
         n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093,
         n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101,
         n18102, n18103, n18104, n18105, n18106, n18107, n18108, n18109,
         n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117,
         n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125,
         n18126, n18127, n18128, n18129, n18130, n18131, n18132, n18133,
         n18134, n18135, n18136, n18137, n18138, n18139, n18140, n18141,
         n18142, n18143, n18144, n18145, n18146, n18147, n18148, n18149,
         n18150, n18151, n18152, n18153, n18154, n18155, n18156, n18157,
         n18158, n18159, n18160, n18161, n18162, n18163, n18164, n18165,
         n18166, n18167, n18168, n18169, n18170, n18171, n18172, n18173,
         n18174, n18175, n18176, n18177, n18178, n18179, n18180, n18181,
         n18182, n18183, n18184, n18185, n18186, n18187, n18188, n18189,
         n18190, n18191, n18192, n18193, n18194, n18195, n18196, n18197,
         n18198, n18199, n18200, n18201, n18202, n18203, n18204, n18205,
         n18206, n18207, n18208, n18209, n18210, n18211, n18212, n18213,
         n18214, n18215, n18216, n18217, n18218, n18219, n18220, n18221,
         n18222, n18223, n18224, n18225, n18226, n18227, n18228, n18229,
         n18230, n18231, n18232, n18233, n18234, n18235, n18236, n18237,
         n18238, n18239, n18240, n18241, n18242, n18243, n18244, n18245,
         n18246, n18247, n18248, n18249, n18250, n18251, n18252, n18253,
         n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18261,
         n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18269,
         n18270, n18271, n18272, n18273, n18274, n18275, n18276, n18277,
         n18278, n18279, n18280, n18281, n18282, n18283, n18284, n18285,
         n18286, n18287, n18288, n18289, n18290, n18291, n18292, n18293,
         n18294, n18295, n18296, n18297, n18298, n18299, n18300, n18301,
         n18302, n18303, n18304, n18305, n18306, n18307, n18308, n18309,
         n18310, n18311, n18312, n18313, n18314, n18315, n18316, n18317,
         n18318, n18319, n18320, n18321, n18322, n18323, n18324, n18325,
         n18326, n18327, n18328, n18329, n18330, n18331, n18332, n18333,
         n18334, n18335, n18336, n18337, n18338, n18339, n18340, n18341,
         n18342, n18343, n18344, n18345, n18346, n18347, n18348, n18349,
         n18350, n18351, n18352, n18353, n18354, n18355, n18356, n18357,
         n18358, n18359, n18360, n18361, n18362, n18363, n18364, n18365,
         n18366, n18367, n18368, n18369, n18370, n18371, n18372, n18373,
         n18374, n18375, n18376, n18377, n18378, n18379, n18380, n18381,
         n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389,
         n18390, n18391, n18392, n18393, n18394, n18395, n18396, n18397,
         n18398, n18399, n18400, n18401, n18402, n18403, n18404, n18405,
         n18406, n18407, n18408, n18409, n18410, n18411, n18412, n18413,
         n18414, n18415, n18416, n18417, n18418, n18419, n18420, n18421,
         n18422, n18423, n18424, n18425, n18426, n18427, n18428, n18429,
         n18430, n18431, n18432, n18433, n18434, n18435, n18436, n18437,
         n18438, n18439, n18440, n18441, n18442, n18443, n18444, n18445,
         n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453,
         n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18461,
         n18462, n18463, n18464, n18465, n18466, n18467, n18468, n18469,
         n18470, n18471, n18472, n18473, n18474, n18475, n18476, n18477,
         n18478, n18479, n18480, n18481, n18482, n18483, n18484, n18485,
         n18486, n18487, n18488, n18489, n18490, n18491, n18492, n18493,
         n18494, n18495, n18496, n18497, n18498, n18499, n18500, n18501,
         n18502, n18503, n18504, n18505, n18506, n18507, n18508, n18509,
         n18510, n18511, n18512, n18513, n18514, n18515, n18516, n18517,
         n18518, n18519, n18520, n18521, n18522, n18523, n18524, n18525,
         n18526, n18527, n18528, n18529, n18530, n18531, n18532, n18533,
         n18534, n18535, n18536, n18537, n18538, n18539, n18540, n18541,
         n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549,
         n18550, n18551, n18552, n18553, n18554, n18555, n18556, n18557,
         n18558, n18559, n18560, n18561, n18562, n18563, n18564, n18565,
         n18566, n18567, n18568, n18569, n18570, n18571, n18572, n18573,
         n18574, n18575, n18576, n18577, n18578, n18579, n18580, n18581,
         n18582, n18583, n18584, n18585, n18586, n18587, n18588, n18589,
         n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597,
         n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605,
         n18606, n18607, n18608, n18609, n18610, n18611, n18612, n18613,
         n18614, n18615, n18616, n18617, n18618, n18619, n18620, n18621,
         n18622, n18623, n18624, n18625, n18626, n18627, n18628, n18629,
         n18630, n18631, n18632, n18633, n18634, n18635, n18636, n18637,
         n18638, n18639, n18640, n18641, n18642, n18643, n18644, n18645,
         n18646, n18647, n18648, n18649, n18650, n18651, n18652, n18653,
         n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18661,
         n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669,
         n18670, n18671, n18672, n18673, n18674, n18675, n18676, n18677,
         n18678, n18679, n18680, n18681, n18682, n18683, n18684, n18685,
         n18686, n18687, n18688, n18689, n18690, n18691, n18692, n18693,
         n18694, n18695, n18696, n18697, n18698, n18699, n18700, n18701,
         n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709,
         n18710, n18711, n18712, n18713, n18714, n18715, n18716, n18717,
         n18718, n18719, n18720, n18721, n18722, n18723, n18724, n18725,
         n18726, n18727, n18728, n18729, n18730, n18731, n18732, n18733,
         n18734, n18735, n18736, n18737, n18738, n18739, n18740, n18741,
         n18742, n18743, n18744, n18745, n18746, n18747, n18748, n18749,
         n18750, n18751, n18752, n18753, n18754, n18755, n18756, n18757,
         n18758, n18759, n18760, n18761, n18762, n18763, n18764, n18765,
         n18766, n18767, n18768, n18769, n18770, n18771, n18772, n18773,
         n18774, n18775, n18776, n18777, n18778, n18779, n18780, n18781,
         n18782, n18783, n18784, n18785, n18786, n18787, n18788, n18789,
         n18790, n18791, n18792, n18793, n18794, n18795, n18796, n18797,
         n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18805,
         n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813,
         n18814, n18815, n18816, n18817, n18818, n18819, n18820, n18821,
         n18822, n18823, n18824, n18825, n18826, n18827, n18828, n18829,
         n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837,
         n18838, n18839, n18840, n18841, n18842, n18843, n18844, n18845,
         n18846, n18847, n18848, n18849, n18850, n18851, n18852, n18853,
         n18854, n18855, n18856, n18857, n18858, n18859, n18860, n18861,
         n18862, n18863, n18864, n18865, n18866, n18867, n18868, n18869,
         n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877,
         n18878, n18879, n18880, n18881, n18882, n18883, n18884, n18885,
         n18886, n18887, n18888, n18889, n18890, n18891, n18892, n18893,
         n18894, n18895, n18896, n18897, n18898, n18899, n18900, n18901,
         n18902, n18903, n18904, n18905, n18906, n18907, n18908, n18909,
         n18910, n18911, n18912, n18913, n18914, n18915, n18916, n18917,
         n18918, n18919, n18920, n18921, n18922, n18923, n18924, n18925,
         n18926, n18927, n18928, n18929, n18930, n18931, n18932, n18933,
         n18934, n18935, n18936, n18937, n18938, n18939, n18940, n18941,
         n18942, n18943, n18944, n18945, n18946, n18947, n18948, n18949,
         n18950, n18951, n18952, n18953, n18954, n18955, n18956, n18957,
         n18958, n18959, n18960, n18961, n18962, n18963, n18964, n18965,
         n18966, n18967, n18968, n18969, n18970, n18971, n18972, n18973,
         n18974, n18975, n18976, n18977, n18978, n18979, n18980, n18981,
         n18982, n18983, n18984, n18985, n18986, n18987, n18988, n18989,
         n18990, n18991, n18992, n18993, n18994, n18995, n18996, n18997,
         n18998, n18999, n19000, n19001, n19002, n19003, n19004, n19005,
         n19006, n19007, n19008, n19009, n19010, n19011, n19012, n19013,
         n19014, n19015, n19016, n19017, n19018, n19019, n19020, n19021,
         n19022, n19023, n19024, n19025, n19026, n19027, n19028, n19029,
         n19030, n19031, n19032, n19033, n19034, n19035, n19036, n19037,
         n19038, n19039, n19040, n19041, n19042, n19043, n19044, n19045,
         n19046, n19047, n19048, n19049, n19050, n19051, n19052, n19053,
         n19054, n19055, n19056, n19057, n19058, n19059, n19060, n19061,
         n19062, n19063, n19064, n19065, n19066, n19067, n19068, n19069,
         n19070, n19071, n19072, n19073, n19074, n19075, n19076, n19077,
         n19078, n19079, n19080, n19081, n19082, n19083, n19084, n19085,
         n19086, n19087, n19088, n19089, n19090, n19091, n19092, n19093,
         n19094, n19095, n19096, n19097, n19098, n19099, n19100, n19101,
         n19102, n19103, n19104, n19105, n19106, n19107, n19108, n19109,
         n19110, n19111, n19112, n19113, n19114, n19115, n19116, n19117,
         n19118, n19119, n19120, n19121, n19122, n19123, n19124, n19125,
         n19126, n19127, n19128, n19129, n19130, n19131, n19132, n19133,
         n19134, n19135, n19136, n19137, n19138, n19139, n19140, n19141,
         n19142, n19143, n19144, n19145, n19146, n19147, n19148, n19149,
         n19150, n19151, n19152, n19153, n19154, n19155, n19156, n19157,
         n19158, n19159, n19160, n19161, n19162, n19163, n19164, n19165,
         n19166, n19167, n19168, n19169, n19170, n19171, n19172, n19173,
         n19174, n19175, n19176, n19177, n19178, n19179, n19180, n19181,
         n19182, n19183, n19184, n19185, n19186, n19187, n19188, n19189,
         n19190, n19191, n19192, n19193, n19194, n19195, n19196, n19197,
         n19198, n19199, n19200, n19201, n19202, n19203, n19204, n19205,
         n19206, n19207, n19208, n19209, n19210, n19211, n19212, n19213,
         n19214, n19215, n19216, n19217, n19218, n19219, n19220, n19221,
         n19222, n19223, n19224, n19225, n19226, n19227, n19228, n19229,
         n19230, n19231, n19232, n19233, n19234, n19235, n19236, n19237,
         n19238, n19239, n19240, n19241, n19242, n19243, n19244, n19245,
         n19246, n19247, n19248, n19249, n19250, n19251, n19252, n19253,
         n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261,
         n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269,
         n19270, n19271, n19272, n19273, n19274, n19275, n19276, n19277,
         n19278, n19279, n19280, n19281, n19282, n19283, n19284, n19285,
         n19286, n19287, n19288, n19289, n19290, n19291, n19292, n19293,
         n19294, n19295, n19296, n19297, n19298, n19299, n19300, n19301,
         n19302, n19303, n19304, n19305, n19306, n19307, n19308, n19309,
         n19310, n19311, n19312, n19313, n19314, n19315, n19316, n19317,
         n19318, n19319, n19320, n19321, n19322, n19323, n19324, n19325,
         n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333,
         n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341,
         n19342, n19343, n19344, n19345, n19346, n19347, n19348, n19349,
         n19350, n19351, n19352, n19353, n19354, n19355, n19356, n19357,
         n19358, n19359, n19360, n19361, n19362, n19363, n19364, n19365,
         n19366, n19367, n19368, n19369, n19370, n19371, n19372, n19373,
         n19374, n19375, n19376, n19377, n19378, n19379, n19380, n19381,
         n19382, n19383, n19384, n19385, n19386, n19387, n19388, n19389,
         n19390, n19391, n19392, n19393, n19394, n19395, n19396, n19397,
         n19398, n19399, n19400, n19401, n19402, n19403, n19404, n19405,
         n19406, n19407, n19408, n19409, n19410, n19411, n19412, n19413,
         n19414, n19415, n19416, n19417, n19418, n19419, n19420, n19421,
         n19422, n19423, n19424, n19425, n19426, n19427, n19428, n19429,
         n19430, n19431, n19432, n19433, n19434, n19435, n19436, n19437,
         n19438, n19439, n19440, n19441, n19442, n19443, n19444, n19445,
         n19446, n19447, n19448, n19449, n19450, n19451, n19452, n19453,
         n19454, n19455, n19456, n19457, n19458, n19459, n19460, n19461,
         n19462, n19463, n19464, n19465, n19466, n19467, n19468, n19469,
         n19470, n19471, n19472, n19473, n19474, n19475, n19476, n19477,
         n19478, n19479, n19480, n19481, n19482, n19483, n19484, n19485,
         n19486, n19487, n19488, n19489, n19490, n19491, n19492, n19493,
         n19494, n19495, n19496, n19497, n19498, n19499, n19500, n19501,
         n19502, n19503, n19504, n19505, n19506, n19507, n19508, n19509,
         n19510, n19511, n19512, n19513, n19514, n19515, n19516, n19517,
         n19518, n19519, n19520, n19521, n19522, n19523, n19524, n19525,
         n19526, n19527, n19528, n19529, n19530, n19531, n19532, n19533,
         n19534, n19535, n19536, n19537, n19538, n19539, n19540, n19541,
         n19542, n19543, n19544, n19545, n19546, n19547, n19548, n19549,
         n19550, n19551, n19552, n19553, n19554, n19555, n19556, n19557,
         n19558, n19559, n19560, n19561, n19562, n19563, n19564, n19565,
         n19566, n19567, n19568, n19569, n19570, n19571, n19572, n19573,
         n19574, n19575, n19576, n19577, n19578, n19579, n19580, n19581,
         n19582, n19583, n19584, n19585, n19586, n19587, n19588, n19589,
         n19590, n19591, n19592, n19593, n19594, n19595, n19596, n19597,
         n19598, n19599, n19600, n19601, n19602, n19603, n19604, n19605,
         n19606, n19607, n19608, n19609, n19610, n19611, n19612, n19613,
         n19614, n19615, n19616, n19617, n19618, n19619, n19620, n19621,
         n19622, n19623, n19624, n19625, n19626, n19627, n19628, n19629,
         n19630, n19631, n19632, n19633, n19634, n19635, n19636, n19637,
         n19638, n19639, n19640, n19641, n19642, n19643, n19644, n19645,
         n19646, n19647, n19648, n19649, n19650, n19651, n19652, n19653,
         n19654, n19655, n19656, n19657, n19658, n19659, n19660, n19661,
         n19662, n19663, n19664, n19665, n19666, n19667, n19668, n19669,
         n19670, n19671, n19672, n19673, n19674, n19675, n19676, n19677,
         n19678, n19679, n19680, n19681, n19682, n19683, n19684, n19685,
         n19686, n19687, n19688, n19689, n19690, n19691, n19692, n19693,
         n19694, n19695, n19696, n19697, n19698, n19699, n19700, n19701,
         n19702, n19703, n19704, n19705, n19706, n19707, n19708, n19709,
         n19710, n19711, n19712, n19713, n19714, n19715, n19716, n19717,
         n19718, n19719, n19720, n19721, n19722, n19723, n19724, n19725,
         n19726, n19727, n19728, n19729, n19730, n19731, n19732, n19733,
         n19734, n19735, n19736, n19737, n19738, n19739, n19740, n19741,
         n19742, n19743, n19744, n19745, n19746, n19747, n19748, n19749,
         n19750, n19751, n19752, n19753, n19754, n19755, n19756, n19757,
         n19758, n19759, n19760, n19761, n19762, n19763, n19764, n19765,
         n19766, n19767, n19768, n19769, n19770, n19771, n19772, n19773,
         n19774, n19775, n19776, n19777, n19778, n19779, n19780, n19781,
         n19782, n19783, n19784, n19785, n19786, n19787, n19788, n19789,
         n19790, n19791, n19792, n19793, n19794, n19795, n19796, n19797,
         n19798, n19799, n19800, n19801, n19802, n19803, n19804, n19805,
         n19806, n19807, n19808, n19809, n19810, n19811, n19812, n19813,
         n19814, n19815, n19816, n19817, n19818, n19819, n19820, n19821,
         n19822, n19823, n19824, n19825, n19826, n19827, n19828, n19829,
         n19830, n19831, n19832, n19833, n19834, n19835, n19836, n19837,
         n19838, n19839, n19840, n19841, n19842, n19843, n19844, n19845,
         n19846, n19847, n19848, n19849, n19850, n19851, n19852, n19853,
         n19854, n19855, n19856, n19857, n19858, n19859, n19860, n19861,
         n19862, n19863, n19864, n19865, n19866, n19867, n19868, n19869,
         n19870, n19871, n19872, n19873, n19874, n19875, n19876, n19877,
         n19878, n19879, n19880, n19881, n19882, n19883, n19884, n19885,
         n19886, n19887, n19888, n19889, n19890, n19891, n19892, n19893,
         n19894, n19895, n19896, n19897, n19898, n19899, n19900, n19901,
         n19902, n19903, n19904, n19905, n19906, n19907, n19908, n19909,
         n19910, n19911, n19912, n19913, n19914, n19915, n19916, n19917,
         n19918, n19919, n19920, n19921, n19922, n19923, n19924, n19925,
         n19926, n19927, n19928, n19929, n19930, n19931, n19932, n19933,
         n19934, n19935, n19936, n19937, n19938, n19939, n19940, n19941,
         n19942, n19943, n19944, n19945, n19946, n19947, n19948, n19949,
         n19950, n19951, n19952, n19953, n19954, n19955, n19956, n19957,
         n19958, n19959, n19960, n19961, n19962, n19963, n19964, n19965,
         n19966, n19967, n19968, n19969, n19970, n19971, n19972, n19973,
         n19974, n19975, n19976, n19977, n19978, n19979, n19980, n19981,
         n19982, n19983, n19984, n19985, n19986, n19987, n19988, n19989,
         n19990, n19991, n19992, n19993, n19994, n19995, n19996, n19997,
         n19998, n19999, n20000, n20001, n20002, n20003, n20004, n20005,
         n20006, n20007, n20008, n20009, n20010, n20011, n20012, n20013,
         n20014, n20015, n20016, n20017, n20018, n20019, n20020, n20021,
         n20022, n20023, n20024, n20025, n20026, n20027, n20028, n20029,
         n20030, n20031, n20032, n20033, n20034, n20035, n20036, n20037,
         n20038, n20039, n20040, n20041, n20042, n20043, n20044, n20045,
         n20046, n20047, n20048, n20049, n20050, n20051, n20052, n20053,
         n20054, n20055, n20056, n20057, n20058, n20059, n20060, n20061,
         n20062, n20063, n20064, n20065, n20066, n20067, n20068, n20069,
         n20070, n20071, n20072, n20073, n20074, n20075, n20076, n20077,
         n20078, n20079, n20080, n20081, n20082, n20083, n20084, n20085,
         n20086, n20087, n20088, n20089, n20090, n20091, n20092, n20093,
         n20094, n20095, n20096, n20097, n20098, n20099, n20100, n20101,
         n20102, n20103, n20104, n20105, n20106, n20107, n20108, n20109,
         n20110, n20111, n20112, n20113, n20114, n20115, n20116, n20117,
         n20118, n20119, n20120, n20121, n20122, n20123, n20124, n20125,
         n20126, n20127, n20128, n20129, n20130, n20131, n20132, n20133,
         n20134, n20135, n20136, n20137, n20138, n20139, n20140, n20141,
         n20142, n20143, n20144, n20145, n20146, n20147, n20148, n20149,
         n20150, n20151, n20152, n20153, n20154, n20155, n20156, n20157,
         n20158, n20159, n20160, n20161, n20162, n20163, n20164, n20165,
         n20166, n20167, n20168, n20169, n20170, n20171, n20172, n20173,
         n20174, n20175, n20176, n20177, n20178, n20179, n20180, n20181,
         n20182, n20183, n20184, n20185, n20186, n20187, n20188, n20189,
         n20190, n20191, n20192, n20193, n20194, n20195, n20196, n20197,
         n20198, n20199, n20200, n20201, n20202, n20203, n20204, n20205,
         n20206, n20207, n20208, n20209, n20210, n20211, n20212, n20213,
         n20214, n20215, n20216, n20217, n20218, n20219, n20220, n20221,
         n20222, n20223, n20224, n20225, n20226, n20227, n20228, n20229,
         n20230, n20231, n20232, n20233, n20234, n20235, n20236, n20237,
         n20238, n20239, n20240, n20241, n20242, n20243, n20244, n20245,
         n20246, n20247, n20248, n20249, n20250, n20251, n20252, n20253,
         n20254, n20255, n20256, n20257, n20258, n20259, n20260, n20261,
         n20262, n20263, n20264, n20265, n20266, n20267, n20268, n20269,
         n20270, n20271, n20272, n20273, n20274, n20275, n20276, n20277,
         n20278, n20279, n20280, n20281, n20282, n20283, n20284, n20285,
         n20286, n20287, n20288, n20289, n20290, n20291, n20292, n20293,
         n20294, n20295, n20296, n20297, n20298, n20299, n20300, n20301,
         n20302, n20303, n20304, n20305, n20306, n20307, n20308, n20309,
         n20310, n20311, n20312, n20313, n20314, n20315, n20316, n20317,
         n20318, n20319, n20320, n20321, n20322, n20323, n20324, n20325,
         n20326, n20327, n20328, n20329, n20330, n20331, n20332, n20333,
         n20334, n20335, n20336, n20337, n20338, n20339, n20340, n20341,
         n20342, n20343, n20344, n20345, n20346, n20347, n20348, n20349,
         n20350, n20351, n20352, n20353, n20354, n20355, n20356, n20357,
         n20358, n20359, n20360, n20361, n20362, n20363, n20364, n20365,
         n20366, n20367, n20368, n20369, n20370, n20371, n20372, n20373,
         n20374, n20375, n20376, n20377, n20378, n20379, n20380, n20381,
         n20382, n20383, n20384, n20385, n20386, n20387, n20388, n20389,
         n20390, n20391, n20392, n20393, n20394, n20395, n20396, n20397,
         n20398, n20399, n20400, n20401, n20402, n20403, n20404, n20405,
         n20406, n20407, n20408, n20409, n20410, n20411, n20412, n20413,
         n20414, n20415, n20416, n20417, n20418, n20419, n20420, n20421,
         n20422, n20423, n20424, n20425, n20426, n20427, n20428, n20429,
         n20430, n20431, n20432, n20433, n20434, n20435, n20436, n20437,
         n20438, n20439, n20440, n20441, n20442, n20443, n20444, n20445,
         n20446, n20447, n20448, n20449, n20450, n20451, n20452, n20453,
         n20454, n20455, n20456, n20457, n20458, n20459, n20460, n20461,
         n20462, n20463, n20464, n20465, n20466, n20467, n20468, n20469,
         n20470, n20471, n20472, n20473, n20474, n20475, n20476, n20477,
         n20478, n20479, n20480, n20481, n20482, n20483, n20484, n20485,
         n20486, n20487, n20488, n20489, n20490, n20491, n20492, n20493,
         n20494, n20495, n20496, n20497, n20498, n20499, n20500, n20501,
         n20502, n20503, n20504, n20505, n20506, n20507, n20508, n20509,
         n20510, n20511, n20512, n20513, n20514, n20515, n20516, n20517,
         n20518, n20519, n20520, n20521, n20522, n20523, n20524, n20525,
         n20526, n20527, n20528, n20529, n20530, n20531, n20532, n20533,
         n20534, n20535, n20536, n20537, n20538, n20539, n20540, n20541,
         n20542, n20543, n20544, n20545, n20546, n20547, n20548, n20549,
         n20550, n20551, n20552, n20553, n20554, n20555, n20556, n20557,
         n20558, n20559, n20560, n20561, n20562, n20563, n20564, n20565,
         n20566, n20567, n20568, n20569, n20570, n20571, n20572, n20573,
         n20574, n20575, n20576, n20577, n20578, n20579, n20580, n20581,
         n20582, n20583, n20584, n20585, n20586, n20587, n20588, n20589,
         n20590, n20591, n20592, n20593, n20594, n20595, n20596, n20597,
         n20598, n20599, n20600, n20601, n20602, n20603, n20604, n20605,
         n20606, n20607, n20608, n20609, n20610, n20611, n20612, n20613,
         n20614, n20615, n20616, n20617, n20618, n20619, n20620, n20621,
         n20622, n20623, n20624, n20625, n20626, n20627, n20628, n20629,
         n20630, n20631, n20632, n20633, n20634, n20635, n20636, n20637,
         n20638, n20639, n20640, n20641, n20642, n20643, n20644, n20645,
         n20646, n20647, n20648, n20649, n20650, n20651, n20652, n20653,
         n20654, n20655, n20656, n20657, n20658, n20659, n20660, n20661,
         n20662, n20663, n20664, n20665, n20666, n20667, n20668, n20669,
         n20670, n20671, n20672, n20673, n20674, n20675, n20676, n20677,
         n20678, n20679, n20680, n20681, n20682, n20683, n20684, n20685,
         n20686, n20687, n20688, n20689, n20690, n20691, n20692, n20693,
         n20694, n20695, n20696, n20697, n20698, n20699, n20700, n20701,
         n20702, n20703, n20704, n20705, n20706, n20707, n20708, n20709,
         n20710, n20711, n20712, n20713, n20714, n20715, n20716, n20717,
         n20718, n20719, n20720, n20721, n20722, n20723, n20724, n20725,
         n20726, n20727, n20728, n20729, n20730, n20731, n20732, n20733,
         n20734, n20735, n20736, n20737, n20738, n20739, n20740, n20741,
         n20742, n20743, n20744, n20745, n20746, n20747, n20748, n20749,
         n20750, n20751, n20752, n20753, n20754, n20755, n20756, n20757,
         n20758, n20759, n20760, n20761, n20762, n20763, n20764, n20765,
         n20766, n20767, n20768, n20769, n20770, n20771, n20772, n20773,
         n20774, n20775, n20776, n20777, n20778, n20779, n20780, n20781,
         n20782, n20783, n20784, n20785, n20786, n20787, n20788, n20789,
         n20790, n20791, n20792, n20793, n20794, n20795, n20796, n20797,
         n20798, n20799, n20800, n20801, n20802, n20803, n20804, n20805,
         n20806, n20807, n20808, n20809, n20810, n20811, n20812, n20813,
         n20814, n20815, n20816, n20817, n20818, n20819, n20820, n20821,
         n20822, n20823, n20824, n20825, n20826, n20827, n20828, n20829,
         n20830, n20831, n20832, n20833, n20834, n20835, n20836, n20837,
         n20838, n20839, n20840, n20841, n20842, n20843, n20844, n20845,
         n20846, n20847, n20848, n20849, n20850, n20851, n20852, n20853,
         n20854, n20855, n20856, n20857, n20858, n20859, n20860, n20861,
         n20862, n20863, n20864, n20865, n20866, n20867, n20868, n20869,
         n20870, n20871, n20872, n20873, n20874, n20875, n20876, n20877,
         n20878, n20879, n20880, n20881, n20882, n20883, n20884, n20885,
         n20886, n20887, n20888, n20889, n20890, n20891, n20892, n20893,
         n20894, n20895, n20896, n20897, n20898, n20899, n20900, n20901,
         n20902, n20903, n20904, n20905, n20906, n20907, n20908, n20909,
         n20910, n20911, n20912, n20913, n20914, n20915, n20916, n20917,
         n20918, n20919, n20920, n20921, n20922, n20923, n20924, n20925,
         n20926, n20927, n20928, n20929, n20930, n20931, n20932, n20933,
         n20934, n20935, n20936, n20937, n20938, n20939, n20940, n20941,
         n20942, n20943, n20944, n20945, n20946, n20947, n20948, n20949,
         n20950, n20951, n20952, n20953, n20954, n20955, n20956, n20957,
         n20958, n20959, n20960, n20961, n20962, n20963, n20964, n20965,
         n20966, n20967, n20968, n20969, n20970, n20971, n20972, n20973,
         n20974, n20975, n20976, n20977, n20978, n20979, n20980, n20981,
         n20982, n20983, n20984, n20985, n20986, n20987, n20988, n20989,
         n20990, n20991, n20992, n20993, n20994, n20995, n20996, n20997,
         n20998, n20999, n21000, n21001, n21002, n21003, n21004, n21005,
         n21006, n21007, n21008, n21009, n21010, n21011, n21012, n21013,
         n21014, n21015, n21016, n21017, n21018, n21019, n21020, n21021,
         n21022, n21023, n21024, n21025, n21026, n21027, n21028, n21029,
         n21030, n21031, n21032, n21033, n21034, n21035, n21036, n21037,
         n21038, n21039, n21040, n21041, n21042, n21043, n21044, n21045,
         n21046, n21047, n21048, n21049, n21050, n21051, n21052, n21053,
         n21054, n21055, n21056, n21057, n21058, n21059, n21060, n21061,
         n21062, n21063, n21064, n21065, n21066, n21067, n21068, n21069,
         n21070, n21071, n21072, n21073, n21074, n21075, n21076, n21077,
         n21078, n21079, n21080, n21081, n21082, n21083, n21084, n21085,
         n21086, n21087, n21088, n21089, n21090, n21091, n21092, n21093,
         n21094, n21095, n21096, n21097, n21098, n21099, n21100, n21101,
         n21102, n21103, n21104, n21105, n21106, n21107, n21108, n21109,
         n21110, n21111, n21112, n21113, n21114, n21115, n21116, n21117,
         n21118, n21119, n21120, n21121, n21122, n21123, n21124, n21125,
         n21126, n21127, n21128, n21129, n21130, n21131, n21132, n21133,
         n21134, n21135, n21136, n21137, n21138, n21139, n21140, n21141,
         n21142, n21143, n21144, n21145, n21146, n21147, n21148, n21149,
         n21150, n21151, n21152, n21153, n21154, n21155, n21156, n21157,
         n21158, n21159, n21160, n21161, n21162, n21163, n21164, n21165,
         n21166, n21167, n21168, n21169, n21170, n21171, n21172, n21173,
         n21174, n21175, n21176, n21177, n21178, n21179, n21180, n21181,
         n21182, n21183, n21184, n21185, n21186, n21187, n21188, n21189,
         n21190, n21191, n21192, n21193, n21194, n21195, n21196, n21197,
         n21198, n21199, n21200, n21201, n21202, n21203, n21204, n21205,
         n21206, n21207, n21208, n21209, n21210, n21211, n21212, n21213,
         n21214, n21215, n21216, n21217, n21218, n21219, n21220, n21221,
         n21222, n21223, n21224, n21225, n21226, n21227, n21228, n21229,
         n21230, n21231, n21232, n21233, n21234, n21235, n21236, n21237,
         n21238, n21239, n21240, n21241, n21242, n21243, n21244, n21245,
         n21246, n21247, n21248, n21249, n21250, n21251, n21252, n21253,
         n21254, n21255, n21256, n21257, n21258, n21259, n21260, n21261,
         n21262, n21263, n21264, n21265, n21266, n21267, n21268, n21269,
         n21270, n21271, n21272, n21273, n21274, n21275, n21276, n21277,
         n21278, n21279, n21280, n21281, n21282, n21283, n21284, n21285,
         n21286, n21287, n21288, n21289, n21290, n21291, n21292, n21293,
         n21294, n21295, n21296, n21297, n21298, n21299, n21300, n21301,
         n21302, n21303, n21304, n21305, n21306, n21307, n21308, n21309,
         n21310, n21311, n21312, n21313, n21314, n21315, n21316, n21317,
         n21318, n21319, n21320, n21321, n21322, n21323, n21324, n21325,
         n21326, n21327, n21328, n21329, n21330, n21331, n21332, n21333,
         n21334, n21335, n21336, n21337, n21338, n21339, n21340, n21341,
         n21342, n21343, n21344, n21345, n21346, n21347, n21348, n21349,
         n21350, n21351, n21352, n21353, n21354, n21355, n21356, n21357,
         n21358, n21359, n21360, n21361, n21362, n21363, n21364, n21365,
         n21366, n21367, n21368, n21369, n21370, n21371, n21372, n21373,
         n21374, n21375, n21376, n21377, n21378, n21379, n21380, n21381,
         n21382, n21383, n21384, n21385, n21386, n21387, n21388, n21389,
         n21390, n21391, n21392, n21393, n21394, n21395, n21396, n21397,
         n21398, n21399, n21400, n21401, n21402, n21403, n21404, n21405,
         n21406, n21407, n21408, n21409, n21410, n21411, n21412, n21413,
         n21414, n21415, n21416, n21417, n21418, n21419, n21420, n21421,
         n21422, n21423, n21424, n21425, n21426, n21427, n21428, n21429,
         n21430, n21431, n21432, n21433, n21434, n21435, n21436, n21437,
         n21438, n21439, n21440, n21441, n21442, n21443, n21444, n21445,
         n21446, n21447, n21448, n21449, n21450, n21451, n21452, n21453,
         n21454, n21455, n21456, n21457, n21458, n21459, n21460, n21461,
         n21462, n21463, n21464, n21465, n21466, n21467, n21468, n21469,
         n21470, n21471, n21472, n21473, n21474, n21475, n21476, n21477,
         n21478, n21479, n21480, n21481, n21482, n21483, n21484, n21485,
         n21486, n21487, n21488, n21489, n21490, n21491, n21492, n21493,
         n21494, n21495, n21496, n21497, n21498, n21499, n21500, n21501,
         n21502, n21503, n21504, n21505, n21506, n21507, n21508, n21509,
         n21510, n21511, n21512, n21513, n21514, n21515, n21516, n21517,
         n21518, n21519, n21520, n21521, n21522, n21523, n21524, n21525,
         n21526, n21527, n21528, n21529, n21530, n21531, n21532, n21533,
         n21534, n21535, n21536, n21537, n21538, n21539, n21540, n21541,
         n21542, n21543, n21544, n21545, n21546, n21547, n21548, n21549,
         n21550, n21551, n21552, n21553, n21554, n21555, n21556, n21557,
         n21558, n21559, n21560, n21561, n21562, n21563, n21564, n21565,
         n21566, n21567, n21568, n21569, n21570, n21571, n21572, n21573,
         n21574, n21575, n21576, n21577, n21578, n21579, n21580, n21581,
         n21582, n21583, n21584, n21585, n21586, n21587, n21588, n21589,
         n21590, n21591, n21592, n21593, n21594, n21595, n21596, n21597,
         n21598, n21599, n21600, n21601, n21602, n21603, n21604, n21605,
         n21606, n21607, n21608, n21609, n21610, n21611, n21612, n21613,
         n21614, n21615, n21616, n21617, n21618, n21619, n21620, n21621,
         n21622, n21623, n21624, n21625, n21626, n21627, n21628, n21629,
         n21630, n21631, n21632, n21633, n21634, n21635, n21636, n21637,
         n21638, n21639, n21640, n21641, n21642, n21643, n21644, n21645,
         n21646, n21647, n21648, n21649, n21650, n21651, n21652, n21653,
         n21654, n21655, n21656, n21657, n21658, n21659, n21660, n21661,
         n21662, n21663, n21664, n21665, n21666, n21667, n21668, n21669,
         n21670, n21671, n21672, n21673, n21674, n21675, n21676, n21677,
         n21678, n21679, n21680, n21681, n21682, n21683, n21684, n21685,
         n21686, n21687, n21688, n21689, n21690, n21691, n21692, n21693,
         n21694, n21695, n21696, n21697, n21698, n21699, n21700, n21701,
         n21702, n21703, n21704, n21705, n21706, n21707, n21708, n21709,
         n21710, n21711, n21712, n21713, n21714, n21715, n21716, n21717,
         n21718, n21719, n21720, n21721, n21722, n21723, n21724, n21725,
         n21726, n21727, n21728, n21729, n21730, n21731, n21732, n21733,
         n21734, n21735, n21736, n21737, n21738, n21739, n21740, n21741,
         n21742, n21743, n21744, n21745, n21746, n21747, n21748, n21749,
         n21750, n21751, n21752, n21753, n21754, n21755, n21756, n21757,
         n21758, n21759, n21760, n21761, n21762, n21763, n21764, n21765,
         n21766, n21767, n21768, n21769, n21770, n21771, n21772, n21773,
         n21774, n21775, n21776, n21777, n21778, n21779, n21780, n21781,
         n21782, n21783, n21784, n21785, n21786, n21787, n21788, n21789,
         n21790, n21791, n21792, n21793, n21794, n21795, n21796, n21797,
         n21798, n21799, n21800, n21801, n21802, n21803, n21804, n21805,
         n21806, n21807, n21808, n21809, n21810, n21811, n21812, n21813,
         n21814, n21815, n21816, n21817, n21818, n21819, n21820, n21821,
         n21822, n21823, n21824, n21825, n21826, n21827, n21828, n21829,
         n21830, n21831, n21832, n21833, n21834, n21835, n21836, n21837,
         n21838, n21839, n21840, n21841, n21842, n21843, n21844, n21845,
         n21846, n21847, n21848, n21849, n21850, n21851, n21852, n21853,
         n21854, n21855, n21856, n21857, n21858, n21859, n21860, n21861,
         n21862, n21863, n21864, n21865, n21866, n21867, n21868, n21869,
         n21870, n21871, n21872, n21873, n21874, n21875, n21876, n21877,
         n21878, n21879, n21880, n21881, n21882, n21883, n21884, n21885,
         n21886, n21887, n21888, n21889, n21890, n21891, n21892, n21893,
         n21894, n21895, n21896, n21897, n21898, n21899, n21900, n21901,
         n21902, n21903, n21904, n21905, n21906, n21907, n21908, n21909,
         n21910, n21911, n21912, n21913, n21914, n21915, n21916, n21917,
         n21918, n21919, n21920, n21921, n21922, n21923, n21924, n21925,
         n21926, n21927, n21928, n21929, n21930, n21931, n21932, n21933,
         n21934, n21935, n21936, n21937, n21938, n21939, n21940, n21941,
         n21942, n21943, n21944, n21945, n21946, n21947, n21948, n21949,
         n21950, n21951, n21952, n21953, n21954, n21955, n21956, n21957,
         n21958, n21959, n21960, n21961, n21962, n21963, n21964, n21965,
         n21966, n21967, n21968, n21969, n21970, n21971, n21972, n21973,
         n21974, n21975, n21976, n21977, n21978, n21979, n21980, n21981,
         n21982, n21983, n21984, n21985, n21986, n21987, n21988, n21989,
         n21990, n21991, n21992, n21993, n21994, n21995, n21996, n21997,
         n21998, n21999, n22000, n22001, n22002, n22003, n22004, n22005,
         n22006, n22007, n22008, n22009, n22010, n22011, n22012, n22013,
         n22014, n22015, n22016, n22017, n22018, n22019, n22020, n22021,
         n22022, n22023, n22024, n22025, n22026, n22027, n22028, n22029,
         n22030, n22031, n22032, n22033, n22034, n22035, n22036, n22037,
         n22038, n22039, n22040, n22041, n22042, n22043, n22044, n22045,
         n22046, n22047, n22048, n22049, n22050, n22051, n22052, n22053,
         n22054, n22055, n22056, n22057, n22058, n22059, n22060, n22061,
         n22062, n22063, n22064, n22065, n22066, n22067, n22068, n22069,
         n22070, n22071, n22072, n22073, n22074, n22075, n22076, n22077,
         n22078, n22079, n22080, n22081, n22082, n22083, n22084, n22085,
         n22086, n22087, n22088, n22089, n22090, n22091, n22092, n22093,
         n22094, n22095, n22096, n22097, n22098, n22099, n22100, n22101,
         n22102, n22103, n22104, n22105, n22106, n22107, n22108, n22109,
         n22110, n22111, n22112, n22113, n22114, n22115, n22116, n22117,
         n22118, n22119, n22120, n22121, n22122, n22123, n22124, n22125,
         n22126, n22127, n22128, n22129, n22130, n22131, n22132, n22133,
         n22134, n22135, n22136, n22137, n22138, n22139, n22140, n22141,
         n22142, n22143, n22144, n22145, n22146, n22147, n22148, n22149,
         n22150, n22151, n22152, n22153, n22154, n22155, n22156, n22157,
         n22158, n22159, n22160, n22161, n22162, n22163, n22164, n22165,
         n22166, n22167, n22168, n22169, n22170, n22171, n22172, n22173,
         n22174, n22175, n22176, n22177, n22178, n22179, n22180, n22181,
         n22182, n22183, n22184, n22185, n22186, n22187, n22188, n22189,
         n22190, n22191, n22192, n22193, n22194, n22195, n22196, n22197,
         n22198, n22199, n22200, n22201, n22202, n22203, n22204, n22205,
         n22206, n22207, n22208, n22209, n22210, n22211, n22212, n22213,
         n22214, n22215, n22216, n22217, n22218, n22219, n22220, n22221,
         n22222, n22223, n22224, n22225, n22226, n22227, n22228, n22229,
         n22230, n22231, n22232, n22233, n22234, n22235, n22236, n22237,
         n22238, n22239, n22240, n22241, n22242, n22243, n22244, n22245,
         n22246, n22247, n22248, n22249, n22250, n22251, n22252, n22253,
         n22254, n22255, n22256, n22257, n22258, n22259, n22260, n22261,
         n22262, n22263, n22264, n22265, n22266, n22267, n22268, n22269,
         n22270, n22271, n22272, n22273, n22274, n22275, n22276, n22277,
         n22278, n22279, n22280, n22281, n22282, n22283, n22284, n22285,
         n22286, n22287, n22288, n22289, n22290, n22291, n22292, n22293,
         n22294, n22295, n22296, n22297, n22298, n22299, n22300, n22301,
         n22302, n22303, n22304, n22305, n22306, n22307, n22308, n22309,
         n22310, n22311, n22312, n22313, n22314, n22315, n22316, n22317,
         n22318, n22319, n22320, n22321, n22322, n22323, n22324, n22325,
         n22326, n22327, n22328, n22329, n22330, n22331, n22332, n22333,
         n22334, n22335, n22336, n22337, n22338, n22339, n22340, n22341,
         n22342, n22343, n22344, n22345, n22346, n22347, n22348, n22349,
         n22350, n22351, n22352, n22353, n22354, n22355, n22356, n22357,
         n22358, n22359, n22360, n22361, n22362, n22363, n22364, n22365,
         n22366, n22367, n22368, n22369, n22370, n22371, n22372, n22373,
         n22374, n22375, n22376, n22377, n22378, n22379, n22380, n22381,
         n22382, n22383, n22384, n22385, n22386, n22387, n22388, n22389,
         n22390, n22391, n22392, n22393, n22394, n22395, n22396, n22397,
         n22398, n22399, n22400, n22401, n22402, n22403, n22404, n22405,
         n22406, n22407, n22408, n22409, n22410, n22411, n22412, n22413,
         n22414, n22415, n22416, n22417, n22418, n22419, n22420, n22421,
         n22422, n22423, n22424, n22425, n22426, n22427, n22428, n22429,
         n22430, n22431, n22432, n22433, n22434, n22435, n22436, n22437,
         n22438, n22439, n22440, n22441, n22442, n22443, n22444, n22445,
         n22446, n22447, n22448, n22449, n22450, n22451, n22452, n22453,
         n22454, n22455, n22456, n22457, n22458, n22459, n22460, n22461,
         n22462, n22463, n22464, n22465, n22466, n22467, n22468, n22469,
         n22470, n22471, n22472, n22473, n22474, n22475, n22476, n22477,
         n22478, n22479, n22480, n22481, n22482, n22483, n22484, n22485,
         n22486, n22487, n22488, n22489, n22490, n22491, n22492, n22493,
         n22494, n22495, n22496, n22497, n22498, n22499, n22500, n22501,
         n22502, n22503, n22504, n22505, n22506, n22507, n22508, n22509,
         n22510, n22511, n22512, n22513, n22514, n22515, n22516, n22517,
         n22518, n22519, n22520, n22521, n22522, n22523, n22524, n22525,
         n22526, n22527, n22528, n22529, n22530, n22531, n22532, n22533,
         n22534, n22535, n22536, n22537, n22538, n22539, n22540, n22541,
         n22542, n22543, n22544, n22545, n22546, n22547, n22548, n22549,
         n22550, n22551, n22552, n22553, n22554, n22555, n22556, n22557,
         n22558, n22559, n22560, n22561, n22562, n22563, n22564, n22565,
         n22566, n22567, n22568, n22569, n22570, n22571, n22572, n22573,
         n22574, n22575, n22576, n22577, n22578, n22579, n22580, n22581,
         n22582, n22583, n22584, n22585, n22586, n22587, n22588, n22589,
         n22590, n22591, n22592, n22593, n22594, n22595, n22596, n22597,
         n22598, n22599, n22600, n22601, n22602, n22603, n22604, n22605,
         n22606, n22607, n22608, n22609, n22610, n22611, n22612, n22613,
         n22614, n22615, n22616, n22617, n22618, n22619, n22620, n22621,
         n22622, n22623, n22624, n22625, n22626, n22627, n22628, n22629,
         n22630, n22631, n22632, n22633, n22634, n22635, n22636, n22637,
         n22638, n22639, n22640, n22641, n22642, n22643, n22644, n22645,
         n22646, n22647, n22648, n22649, n22650, n22651, n22652, n22653,
         n22654, n22655, n22656, n22657, n22658, n22659, n22660, n22661,
         n22662, n22663, n22664, n22665, n22666, n22667, n22668, n22669,
         n22670, n22671, n22672, n22673, n22674, n22675, n22676, n22677,
         n22678, n22679, n22680, n22681, n22682, n22683, n22684, n22685,
         n22686, n22687, n22688, n22689, n22690, n22691, n22692, n22693,
         n22694, n22695, n22696, n22697, n22698, n22699, n22700, n22701,
         n22702, n22703, n22704, n22705, n22706, n22707, n22708, n22709,
         n22710, n22711, n22712, n22713, n22714, n22715, n22716, n22717,
         n22718, n22719, n22720, n22721, n22722, n22723, n22724, n22725,
         n22726, n22727, n22728, n22729, n22730, n22731, n22732, n22733,
         n22734, n22735, n22736, n22737, n22738, n22739, n22740, n22741,
         n22742, n22743, n22744, n22745, n22746, n22747, n22748, n22749,
         n22750, n22751, n22752, n22753, n22754, n22755, n22756, n22757,
         n22758, n22759, n22760, n22761, n22762, n22763, n22764, n22765,
         n22766, n22767, n22768, n22769, n22770, n22771, n22772, n22773,
         n22774, n22775, n22776, n22777, n22778, n22779, n22780, n22781,
         n22782, n22783, n22784, n22785, n22786, n22787, n22788, n22789,
         n22790, n22791, n22792, n22793, n22794, n22795, n22796, n22797,
         n22798, n22799, n22800, n22801, n22802, n22803, n22804, n22805,
         n22806, n22807, n22808, n22809, n22810, n22811, n22812, n22813,
         n22814, n22815, n22816, n22817, n22818, n22819, n22820, n22821,
         n22822, n22823, n22824, n22825, n22826, n22827, n22828, n22829,
         n22830, n22831, n22832, n22833, n22834, n22835, n22836, n22837,
         n22838, n22839, n22840, n22841, n22842, n22843, n22844, n22845,
         n22846, n22847, n22848, n22849, n22850, n22851, n22852, n22853,
         n22854, n22855, n22856, n22857, n22858, n22859, n22860, n22861,
         n22862, n22863, n22864, n22865, n22866, n22867, n22868, n22869,
         n22870, n22871, n22872, n22873, n22874, n22875, n22876, n22877,
         n22878, n22879, n22880, n22881, n22882, n22883, n22884, n22885,
         n22886, n22887, n22888, n22889, n22890, n22891, n22892, n22893,
         n22894, n22895, n22896, n22897, n22898, n22899, n22900, n22901,
         n22902, n22903, n22904, n22905, n22906, n22907, n22908, n22909,
         n22910, n22911, n22912, n22913, n22914, n22915, n22916, n22917,
         n22918, n22919, n22920, n22921, n22922, n22923, n22924, n22925,
         n22926, n22927, n22928, n22929, n22930, n22931, n22932, n22933,
         n22934, n22935, n22936, n22937, n22938, n22939, n22940, n22941,
         n22942, n22943, n22944, n22945, n22946, n22947, n22948, n22949,
         n22950, n22951, n22952, n22953, n22954, n22955, n22956, n22957,
         n22958, n22959, n22960, n22961, n22962, n22963, n22964, n22965,
         n22966, n22967, n22968, n22969, n22970, n22971, n22972, n22973,
         n22974, n22975, n22976, n22977, n22978, n22979, n22980, n22981,
         n22982, n22983, n22984, n22985, n22986, n22987, n22988, n22989,
         n22990, n22991, n22992, n22993, n22994, n22995, n22996, n22997,
         n22998, n22999, n23000, n23001, n23002, n23003, n23004, n23005,
         n23006, n23007, n23008, n23009, n23010, n23011, n23012, n23013,
         n23014, n23015, n23016, n23017, n23018, n23019, n23020, n23021,
         n23022, n23023, n23024, n23025, n23026, n23027, n23028, n23029,
         n23030, n23031, n23032, n23033, n23034, n23035, n23036, n23037,
         n23038, n23039, n23040, n23041, n23042, n23043, n23044, n23045,
         n23046, n23047, n23048, n23049, n23050, n23051, n23052, n23053,
         n23054, n23055, n23056, n23057, n23058, n23059, n23060, n23061,
         n23062, n23063, n23064, n23065, n23066, n23067, n23068, n23069,
         n23070, n23071, n23072, n23073, n23074, n23075, n23076, n23077,
         n23078, n23079, n23080, n23081, n23082, n23083, n23084, n23085,
         n23086, n23087, n23088, n23089, n23090, n23091, n23092, n23093,
         n23094, n23095, n23096, n23097, n23098, n23099, n23100, n23101,
         n23102, n23103, n23104, n23105, n23106, n23107, n23108, n23109,
         n23110, n23111, n23112, n23113, n23114, n23115, n23116, n23117,
         n23118, n23119, n23120, n23121, n23122, n23123, n23124, n23125,
         n23126, n23127, n23128, n23129, n23130, n23131, n23132, n23133,
         n23134, n23135, n23136, n23137, n23138, n23139, n23140, n23141,
         n23142, n23143, n23144, n23145, n23146, n23147, n23148, n23149,
         n23150, n23151, n23152, n23153, n23154, n23155, n23156, n23157,
         n23158, n23159, n23160, n23161, n23162, n23163, n23164, n23165,
         n23166, n23167, n23168, n23169, n23170, n23171, n23172, n23173,
         n23174, n23175, n23176, n23177, n23178, n23179, n23180, n23181,
         n23182, n23183, n23184, n23185, n23186, n23187, n23188, n23189,
         n23190, n23191, n23192, n23193, n23194, n23195, n23196, n23197,
         n23198, n23199, n23200, n23201, n23202, n23203, n23204, n23205,
         n23206, n23207, n23208, n23209, n23210, n23211, n23212, n23213,
         n23214, n23215, n23216, n23217, n23218, n23219, n23220, n23221,
         n23222, n23223, n23224, n23225, n23226, n23227, n23228, n23229,
         n23230, n23231, n23232, n23233, n23234, n23235, n23236, n23237,
         n23238, n23239, n23240, n23241, n23242, n23243, n23244, n23245,
         n23246, n23247, n23248, n23249, n23250, n23251, n23252, n23253,
         n23254, n23255, n23256, n23257, n23258, n23259, n23260, n23261,
         n23262, n23263, n23264, n23265, n23266, n23267, n23268, n23269,
         n23270, n23271, n23272, n23273, n23274, n23275, n23276, n23277,
         n23278, n23279, n23280, n23281, n23282, n23283, n23284, n23285,
         n23286, n23287, n23288, n23289, n23290, n23291, n23292, n23293,
         n23294, n23295, n23296, n23297, n23298, n23299, n23300, n23301,
         n23302, n23303, n23304, n23305, n23306, n23307, n23308, n23309,
         n23310, n23311, n23312, n23313, n23314, n23315, n23316, n23317,
         n23318, n23319, n23320, n23321, n23322, n23323, n23324, n23325,
         n23326, n23327, n23328, n23329, n23330, n23331, n23332, n23333,
         n23334, n23335, n23336, n23337, n23338, n23339, n23340, n23341,
         n23342, n23343, n23344, n23345, n23346, n23347, n23348, n23349,
         n23350, n23351, n23352, n23353, n23354, n23355, n23356, n23357,
         n23358, n23359, n23360, n23361, n23362, n23363, n23364, n23365,
         n23366, n23367, n23368, n23369, n23370, n23371, n23372, n23373,
         n23374, n23375, n23376, n23377, n23378, n23379, n23380, n23381,
         n23382, n23383, n23384, n23385, n23386, n23387, n23388, n23389,
         n23390, n23391, n23392, n23393, n23394, n23395, n23396, n23397,
         n23398, n23399, n23400, n23401, n23402, n23403, n23404, n23405,
         n23406, n23407, n23408, n23409, n23410, n23411, n23412, n23413,
         n23414, n23415, n23416, n23417, n23418, n23419, n23420, n23421,
         n23422, n23423, n23424, n23425, n23426, n23427, n23428, n23429,
         n23430, n23431, n23432, n23433, n23434, n23435, n23436, n23437,
         n23438, n23439, n23440, n23441, n23442, n23443, n23444, n23445,
         n23446, n23447, n23448, n23449, n23450, n23451, n23452, n23453,
         n23454, n23455, n23456, n23457, n23458, n23459, n23460, n23461,
         n23462, n23463, n23464, n23465, n23466, n23467, n23468, n23469,
         n23470, n23471, n23472, n23473, n23474, n23475, n23476, n23477,
         n23478, n23479, n23480, n23481, n23482, n23483, n23484, n23485,
         n23486, n23487, n23488, n23489, n23490, n23491, n23492, n23493,
         n23494, n23495, n23496, n23497, n23498, n23499, n23500, n23501,
         n23502, n23503, n23504, n23505, n23506, n23507, n23508, n23509,
         n23510, n23511, n23512, n23513, n23514, n23515, n23516, n23517,
         n23518, n23519, n23520, n23521, n23522, n23523, n23524, n23525,
         n23526, n23527, n23528, n23529, n23530, n23531, n23532, n23533,
         n23534, n23535, n23536, n23537, n23538, n23539, n23540, n23541,
         n23542, n23543, n23544, n23545, n23546, n23547, n23548, n23549,
         n23550, n23551, n23552, n23553, n23554, n23555, n23556, n23557,
         n23558, n23559, n23560, n23561, n23562, n23563, n23564, n23565,
         n23566, n23567, n23568, n23569, n23570, n23571, n23572, n23573,
         n23574, n23575, n23576, n23577, n23578, n23579, n23580, n23581,
         n23582, n23583, n23584, n23585, n23586, n23587, n23588, n23589,
         n23590, n23591, n23592, n23593, n23594, n23595, n23596, n23597,
         n23598, n23599, n23600, n23601, n23602, n23603, n23604, n23605,
         n23606, n23607, n23608, n23609, n23610, n23611, n23612, n23613,
         n23614, n23615, n23616, n23617, n23618, n23619, n23620, n23621,
         n23622, n23623, n23624, n23625, n23626, n23627, n23628, n23629,
         n23630, n23631, n23632, n23633, n23634, n23635, n23636, n23637,
         n23638, n23639, n23640, n23641, n23642, n23643, n23644, n23645,
         n23646, n23647, n23648, n23649, n23650, n23651, n23652, n23653,
         n23654, n23655, n23656, n23657, n23658, n23659, n23660, n23661,
         n23662, n23663, n23664, n23665, n23666, n23667, n23668, n23669,
         n23670, n23671, n23672, n23673, n23674, n23675, n23676, n23677,
         n23678, n23679, n23680, n23681, n23682, n23683, n23684, n23685,
         n23686, n23687, n23688, n23689, n23690, n23691, n23692, n23693,
         n23694, n23695, n23696, n23697, n23698, n23699, n23700, n23701,
         n23702, n23703, n23704, n23705, n23706, n23707, n23708, n23709,
         n23710, n23711, n23712, n23713, n23714, n23715, n23716, n23717,
         n23718, n23719, n23720, n23721, n23722, n23723, n23724, n23725,
         n23726, n23727, n23728, n23729, n23730, n23731, n23732, n23733,
         n23734, n23735, n23736, n23737, n23738, n23739, n23740, n23741,
         n23742, n23743, n23744, n23745, n23746, n23747, n23748, n23749,
         n23750, n23751, n23752, n23753, n23754, n23755, n23756, n23757,
         n23758, n23759, n23760, n23761, n23762, n23763, n23764, n23765,
         n23766, n23767, n23768, n23769, n23770, n23771, n23772, n23773,
         n23774, n23775, n23776, n23777, n23778, n23779, n23780, n23781,
         n23782, n23783, n23784, n23785, n23786, n23787, n23788, n23789,
         n23790, n23791, n23792, n23793, n23794, n23795, n23796, n23797,
         n23798, n23799, n23800, n23801, n23802, n23803, n23804, n23805,
         n23806, n23807, n23808, n23809, n23810, n23811, n23812, n23813,
         n23814, n23815, n23816, n23817, n23818, n23819, n23820, n23821,
         n23822, n23823, n23824, n23825, n23826, n23827, n23828, n23829,
         n23830, n23831, n23832, n23833, n23834, n23835, n23836, n23837,
         n23838, n23839, n23840, n23841, n23842, n23843, n23844, n23845,
         n23846, n23847, n23848, n23849, n23850, n23851, n23852, n23853,
         n23854, n23855, n23856, n23857, n23858, n23859, n23860, n23861,
         n23862, n23863, n23864, n23865, n23866, n23867, n23868, n23869,
         n23870, n23871, n23872, n23873, n23874, n23875, n23876, n23877,
         n23878, n23879, n23880, n23881, n23882, n23883, n23884, n23885,
         n23886, n23887, n23888, n23889, n23890, n23891, n23892, n23893,
         n23894, n23895, n23896, n23897, n23898, n23899, n23900, n23901,
         n23902, n23903, n23904, n23905, n23906, n23907, n23908, n23909,
         n23910, n23911, n23912, n23913, n23914, n23915, n23916, n23917,
         n23918, n23919, n23920, n23921, n23922, n23923, n23924, n23925,
         n23926, n23927, n23928, n23929, n23930, n23931, n23932, n23933,
         n23934, n23935, n23936, n23937, n23938, n23939, n23940, n23941,
         n23942, n23943, n23944, n23945, n23946, n23947, n23948, n23949,
         n23950, n23951, n23952, n23953, n23954, n23955, n23956, n23957,
         n23958, n23959, n23960, n23961, n23962, n23963, n23964, n23965,
         n23966, n23967, n23968, n23969, n23970, n23971, n23972, n23973,
         n23974, n23975, n23976, n23977, n23978, n23979, n23980, n23981,
         n23982, n23983, n23984, n23985, n23986, n23987, n23988, n23989,
         n23990, n23991, n23992, n23993, n23994, n23995, n23996, n23997,
         n23998, n23999, n24000, n24001, n24002, n24003, n24004, n24005,
         n24006, n24007, n24008, n24009, n24010, n24011, n24012, n24013,
         n24014, n24015, n24016, n24017, n24018, n24019, n24020, n24021,
         n24022, n24023, n24024, n24025, n24026, n24027, n24028, n24029,
         n24030, n24031, n24032, n24033, n24034, n24035, n24036, n24037,
         n24038, n24039, n24040, n24041, n24042, n24043, n24044, n24045,
         n24046, n24047, n24048, n24049, n24050, n24051, n24052, n24053,
         n24054, n24055, n24056, n24057, n24058, n24059, n24060, n24061,
         n24062, n24063, n24064, n24065, n24066, n24067, n24068, n24069,
         n24070, n24071, n24072, n24073, n24074, n24075, n24076, n24077,
         n24078, n24079, n24080, n24081, n24082, n24083, n24084, n24085,
         n24086, n24087, n24088, n24089, n24090, n24091, n24092, n24093,
         n24094, n24095, n24096, n24097, n24098, n24099, n24100, n24101,
         n24102, n24103, n24104, n24105, n24106, n24107, n24108, n24109,
         n24110, n24111, n24112, n24113, n24114, n24115, n24116, n24117,
         n24118, n24119, n24120, n24121, n24122, n24123, n24124, n24125,
         n24126, n24127, n24128, n24129, n24130, n24131, n24132, n24133,
         n24134, n24135, n24136, n24137, n24138, n24139, n24140, n24141,
         n24142, n24143, n24144, n24145, n24146, n24147, n24148, n24149,
         n24150, n24151, n24152, n24153, n24154, n24155, n24156, n24157,
         n24158, n24159, n24160, n24161, n24162, n24163, n24164, n24165,
         n24166, n24167, n24168, n24169, n24170, n24171, n24172, n24173,
         n24174, n24175, n24176, n24177, n24178, n24179, n24180, n24181,
         n24182, n24183, n24184, n24185, n24186, n24187, n24188, n24189,
         n24190, n24191, n24192, n24193, n24194, n24195, n24196, n24197,
         n24198, n24199, n24200, n24201, n24202, n24203, n24204, n24205,
         n24206, n24207, n24208, n24209, n24210, n24211, n24212, n24213,
         n24214, n24215, n24216, n24217, n24218, n24219, n24220, n24221,
         n24222, n24223, n24224, n24225, n24226, n24227, n24228, n24229,
         n24230, n24231, n24232, n24233, n24234, n24235, n24236, n24237,
         n24238, n24239, n24240, n24241, n24242, n24243, n24244, n24245,
         n24246, n24247, n24248, n24249, n24250, n24251, n24252, n24253,
         n24254, n24255, n24256, n24257, n24258, n24259, n24260, n24261,
         n24262, n24263, n24264, n24265, n24266, n24267, n24268, n24269,
         n24270, n24271, n24272, n24273, n24274, n24275, n24276, n24277,
         n24278, n24279, n24280, n24281, n24282, n24283, n24284, n24285,
         n24286, n24287, n24288, n24289, n24290, n24291, n24292, n24293,
         n24294, n24295, n24296, n24297, n24298, n24299, n24300, n24301,
         n24302, n24303, n24304, n24305, n24306, n24307, n24308, n24309,
         n24310, n24311, n24312, n24313, n24314, n24315, n24316, n24317,
         n24318, n24319, n24320, n24321, n24322, n24323, n24324, n24325,
         n24326, n24327, n24328, n24329, n24330, n24331, n24332, n24333,
         n24334, n24335, n24336, n24337, n24338, n24339, n24340, n24341,
         n24342, n24343, n24344, n24345, n24346, n24347, n24348, n24349,
         n24350, n24351, n24352, n24353, n24354, n24355, n24356, n24357,
         n24358, n24359, n24360, n24361, n24362, n24363, n24364, n24365,
         n24366, n24367, n24368, n24369, n24370, n24371, n24372, n24373,
         n24374, n24375, n24376, n24377, n24378, n24379, n24380, n24381,
         n24382, n24383, n24384, n24385, n24386, n24387, n24388, n24389,
         n24390, n24391, n24392, n24393, n24394, n24395, n24396, n24397,
         n24398, n24399, n24400, n24401, n24402, n24403, n24404, n24405,
         n24406, n24407, n24408, n24409, n24410, n24411, n24412, n24413,
         n24414, n24415, n24416, n24417, n24418, n24419, n24420, n24421,
         n24422, n24423, n24424, n24425, n24426, n24427, n24428, n24429,
         n24430, n24431, n24432, n24433, n24434, n24435, n24436, n24437,
         n24438, n24439, n24440, n24441, n24442, n24443, n24444, n24445,
         n24446, n24447, n24448, n24449, n24450, n24451, n24452, n24453,
         n24454, n24455, n24456, n24457, n24458, n24459, n24460, n24461,
         n24462, n24463, n24464, n24465, n24466, n24467, n24468, n24469,
         n24470, n24471, n24472, n24473, n24474, n24475, n24476, n24477,
         n24478, n24479, n24480, n24481, n24482, n24483, n24484, n24485,
         n24486, n24487, n24488, n24489, n24490, n24491, n24492, n24493,
         n24494, n24495, n24496, n24497, n24498, n24499, n24500, n24501,
         n24502, n24503, n24504, n24505, n24506, n24507, n24508, n24509,
         n24510, n24511, n24512, n24513, n24514, n24515, n24516, n24517,
         n24518, n24519, n24520, n24521, n24522, n24523, n24524, n24525,
         n24526, n24527, n24528, n24529, n24530, n24531, n24532, n24533,
         n24534, n24535, n24536, n24537, n24538, n24539, n24540, n24541,
         n24542, n24543, n24544, n24545, n24546, n24547, n24548, n24549,
         n24550, n24551, n24552, n24553, n24554, n24555, n24556, n24557,
         n24558, n24559, n24560, n24561, n24562, n24563, n24564, n24565,
         n24566, n24567, n24568, n24569, n24570, n24571, n24572, n24573,
         n24574, n24575, n24576, n24577, n24578, n24579, n24580, n24581,
         n24582, n24583, n24584, n24585, n24586, n24587, n24588, n24589,
         n24590, n24591, n24592, n24593, n24594, n24595, n24596, n24597,
         n24598, n24599, n24600, n24601, n24602, n24603, n24604, n24605,
         n24606, n24607, n24608, n24609, n24610, n24611, n24612, n24613,
         n24614, n24615, n24616, n24617, n24618, n24619, n24620, n24621,
         n24622, n24623, n24624, n24625, n24626, n24627, n24628, n24629,
         n24630, n24631, n24632, n24633, n24634, n24635, n24636, n24637,
         n24638, n24639, n24640, n24641, n24642, n24643, n24644, n24645,
         n24646, n24647, n24648, n24649, n24650, n24651, n24652, n24653,
         n24654, n24655, n24656, n24657, n24658, n24659, n24660, n24661,
         n24662, n24663, n24664, n24665, n24666, n24667, n24668, n24669,
         n24670, n24671, n24672, n24673, n24674, n24675, n24676, n24677,
         n24678, n24679, n24680, n24681, n24682, n24683, n24684, n24685,
         n24686, n24687, n24688, n24689, n24690, n24691, n24692, n24693,
         n24694, n24695, n24696, n24697, n24698, n24699, n24700, n24701,
         n24702, n24703, n24704, n24705, n24706, n24707, n24708, n24709,
         n24710, n24711, n24712, n24713, n24714, n24715, n24716, n24717,
         n24718, n24719, n24720, n24721, n24722, n24723, n24724, n24725,
         n24726, n24727, n24728, n24729, n24730, n24731, n24732, n24733,
         n24734, n24735, n24736, n24737, n24738, n24739, n24740, n24741,
         n24742, n24743, n24744, n24745, n24746, n24747, n24748, n24749,
         n24750, n24751, n24752, n24753, n24754, n24755, n24756, n24757,
         n24758, n24759, n24760, n24761, n24762, n24763, n24764, n24765,
         n24766, n24767, n24768, n24769, n24770, n24771, n24772, n24773,
         n24774, n24775, n24776, n24777, n24778, n24779, n24780, n24781,
         n24782, n24783, n24784, n24785, n24786, n24787, n24788, n24789,
         n24790, n24791, n24792, n24793, n24794, n24795, n24796, n24797,
         n24798, n24799, n24800, n24801, n24802, n24803, n24804, n24805,
         n24806, n24807, n24808, n24809, n24810, n24811, n24812, n24813,
         n24814, n24815, n24816, n24817, n24818, n24819, n24820, n24821,
         n24822, n24823, n24824, n24825, n24826, n24827, n24828, n24829,
         n24830, n24831, n24832, n24833, n24834, n24835, n24836, n24837,
         n24838, n24839, n24840, n24841, n24842, n24843, n24844, n24845,
         n24846, n24847, n24848, n24849, n24850, n24851, n24852, n24853,
         n24854, n24855, n24856, n24857, n24858, n24859, n24860, n24861,
         n24862, n24863, n24864, n24865, n24866, n24867, n24868, n24869,
         n24870, n24871, n24872, n24873, n24874, n24875, n24876, n24877,
         n24878, n24879, n24880, n24881, n24882, n24883, n24884, n24885,
         n24886, n24887, n24888, n24889, n24890, n24891, n24892, n24893,
         n24894, n24895, n24896, n24897, n24898, n24899, n24900, n24901,
         n24902, n24903, n24904, n24905, n24906, n24907, n24908, n24909,
         n24910, n24911, n24912, n24913, n24914, n24915, n24916, n24917,
         n24918, n24919, n24920, n24921, n24922, n24923, n24924, n24925,
         n24926, n24927, n24928, n24929, n24930, n24931, n24932, n24933,
         n24934, n24935, n24936, n24937, n24938, n24939, n24940, n24941,
         n24942, n24943, n24944, n24945, n24946, n24947, n24948, n24949,
         n24950, n24951, n24952, n24953, n24954, n24955, n24956, n24957,
         n24958, n24959, n24960, n24961, n24962, n24963, n24964, n24965,
         n24966, n24967, n24968, n24969, n24970, n24971, n24972, n24973,
         n24974, n24975, n24976, n24977, n24978, n24979, n24980, n24981,
         n24982, n24983, n24984, n24985, n24986, n24987, n24988, n24989,
         n24990, n24991, n24992, n24993, n24994, n24995, n24996, n24997,
         n24998, n24999, n25000, n25001, n25002, n25003, n25004, n25005,
         n25006, n25007, n25008, n25009, n25010, n25011, n25012, n25013,
         n25014, n25015, n25016, n25017, n25018, n25019, n25020, n25021,
         n25022, n25023, n25024, n25025, n25026, n25027, n25028, n25029,
         n25030, n25031, n25032, n25033, n25034, n25035, n25036, n25037,
         n25038, n25039, n25040, n25041, n25042, n25043, n25044, n25045,
         n25046, n25047, n25048, n25049, n25050, n25051, n25052, n25053,
         n25054, n25055, n25056, n25057, n25058, n25059, n25060, n25061,
         n25062, n25063, n25064, n25065, n25066, n25067, n25068, n25069,
         n25070, n25071, n25072, n25073, n25074, n25075, n25076, n25077,
         n25078, n25079, n25080, n25081, n25082, n25083, n25084, n25085,
         n25086, n25087, n25088, n25089, n25090, n25091, n25092, n25093,
         n25094, n25095, n25096, n25097, n25098, n25099, n25100, n25101,
         n25102, n25103, n25104, n25105, n25106, n25107, n25108, n25109,
         n25110, n25111, n25112, n25113, n25114, n25115, n25116, n25117,
         n25118, n25119, n25120, n25121, n25122, n25123, n25124, n25125,
         n25126, n25127, n25128, n25129, n25130, n25131, n25132, n25133,
         n25134, n25135, n25136, n25137, n25138, n25139, n25140, n25141,
         n25142, n25143, n25144, n25145, n25146, n25147, n25148, n25149,
         n25150, n25151, n25152, n25153, n25154, n25155, n25156, n25157,
         n25158, n25159, n25160, n25161, n25162, n25163, n25164, n25165,
         n25166, n25167, n25168, n25169, n25170, n25171, n25172, n25173,
         n25174, n25175, n25176, n25177, n25178, n25179, n25180, n25181,
         n25182, n25183, n25184, n25185, n25186, n25187, n25188, n25189,
         n25190, n25191, n25192, n25193, n25194, n25195, n25196, n25197,
         n25198, n25199, n25200, n25201, n25202, n25203, n25204, n25205,
         n25206, n25207, n25208, n25209, n25210, n25211, n25212, n25213,
         n25214, n25215, n25216, n25217, n25218, n25219, n25220, n25221,
         n25222, n25223, n25224, n25225, n25226, n25227, n25228, n25229,
         n25230, n25231, n25232, n25233, n25234, n25235, n25236, n25237,
         n25238, n25239, n25240, n25241, n25242, n25243, n25244, n25245,
         n25246, n25247, n25248, n25249, n25250, n25251, n25252, n25253,
         n25254, n25255, n25256, n25257, n25258, n25259, n25260, n25261,
         n25262, n25263, n25264, n25265, n25266, n25267, n25268, n25269,
         n25270, n25271, n25272, n25273, n25274, n25275, n25276, n25277,
         n25278, n25279, n25280, n25281, n25282, n25283, n25284, n25285,
         n25286, n25287, n25288, n25289, n25290, n25291, n25292, n25293,
         n25294, n25295, n25296, n25297, n25298, n25299, n25300, n25301,
         n25302, n25303, n25304, n25305, n25306, n25307, n25308, n25309,
         n25310, n25311, n25312, n25313, n25314, n25315, n25316, n25317,
         n25318, n25319, n25320, n25321, n25322, n25323, n25324, n25325,
         n25326, n25327, n25328, n25329, n25330, n25331, n25332, n25333,
         n25334, n25335, n25336, n25337, n25338, n25339, n25340, n25341,
         n25342, n25343, n25344, n25345, n25346, n25347, n25348, n25349,
         n25350, n25351, n25352, n25353, n25354, n25355, n25356, n25357,
         n25358, n25359, n25360, n25361, n25362, n25363, n25364, n25365,
         n25366, n25367, n25368, n25369, n25370, n25371, n25372, n25373,
         n25374, n25375, n25376, n25377, n25378, n25379, n25380, n25381,
         n25382, n25383, n25384, n25385, n25386, n25387, n25388, n25389,
         n25390, n25391, n25392, n25393, n25394, n25395, n25396, n25397,
         n25398, n25399, n25400, n25401, n25402, n25403, n25404, n25405,
         n25406, n25407, n25408, n25409, n25410, n25411, n25412, n25413,
         n25414, n25415, n25416, n25417, n25418, n25419, n25420, n25421,
         n25422, n25423, n25424, n25425, n25426, n25427, n25428, n25429,
         n25430, n25431, n25432, n25433, n25434, n25435, n25436, n25437,
         n25438, n25439, n25440, n25441, n25442, n25443, n25444, n25445,
         n25446, n25447, n25448, n25449, n25450, n25451, n25452, n25453,
         n25454, n25455, n25456, n25457, n25458, n25459, n25460, n25461,
         n25462, n25463, n25464, n25465, n25466, n25467, n25468, n25469,
         n25470, n25471, n25472, n25473, n25474, n25475, n25476, n25477,
         n25478, n25479, n25480, n25481, n25482, n25483, n25484, n25485,
         n25486, n25487, n25488, n25489, n25490, n25491, n25492, n25493,
         n25494, n25495, n25496, n25497, n25498, n25499, n25500, n25501,
         n25502, n25503, n25504, n25505, n25506, n25507, n25508, n25509,
         n25510, n25511, n25512, n25513, n25514, n25515, n25516, n25517,
         n25518, n25519, n25520, n25521, n25522, n25523, n25524, n25525,
         n25526, n25527, n25528, n25529, n25530, n25531, n25532, n25533,
         n25534, n25535, n25536, n25537, n25538, n25539, n25540, n25541,
         n25542, n25543, n25544, n25545, n25546, n25547, n25548, n25549,
         n25550, n25551, n25552, n25553, n25554, n25555, n25556, n25557,
         n25558, n25559, n25560, n25561, n25562, n25563, n25564, n25565,
         n25566, n25567, n25568, n25569, n25570, n25571, n25572, n25573,
         n25574, n25575, n25576, n25577, n25578, n25579, n25580, n25581,
         n25582, n25583, n25584, n25585, n25586, n25587, n25588, n25589,
         n25590, n25591, n25592, n25593, n25594, n25595, n25596, n25597,
         n25598, n25599, n25600, n25601, n25602, n25603, n25604, n25605,
         n25606, n25607, n25608, n25609, n25610, n25611, n25612, n25613,
         n25614, n25615, n25616, n25617, n25618, n25619, n25620, n25621,
         n25622, n25623, n25624, n25625, n25626, n25627, n25628, n25629,
         n25630, n25631, n25632, n25633, n25634, n25635, n25636, n25637,
         n25638, n25639, n25640, n25641, n25642, n25643, n25644, n25645,
         n25646, n25647, n25648, n25649, n25650, n25651, n25652, n25653,
         n25654, n25655, n25656, n25657, n25658, n25659, n25660, n25661,
         n25662, n25663, n25664, n25665, n25666, n25667, n25668, n25669,
         n25670, n25671, n25672, n25673, n25674, n25675, n25676, n25677,
         n25678, n25679, n25680, n25681, n25682, n25683, n25684, n25685,
         n25686, n25687, n25688, n25689, n25690, n25691, n25692, n25693,
         n25694, n25695, n25696, n25697, n25698, n25699, n25700, n25701,
         n25702, n25703, n25704, n25705, n25706, n25707, n25708, n25709,
         n25710, n25711, n25712, n25713, n25714, n25715, n25716, n25717,
         n25718, n25719, n25720, n25721, n25722, n25723, n25724, n25725,
         n25726, n25727, n25728, n25729, n25730, n25731, n25732, n25733,
         n25734, n25735, n25736, n25737, n25738, n25739, n25740, n25741,
         n25742, n25743, n25744, n25745, n25746, n25747, n25748, n25749,
         n25750, n25751, n25752, n25753, n25754, n25755, n25756, n25757,
         n25758, n25759, n25760, n25761, n25762, n25763, n25764, n25765,
         n25766, n25767, n25768, n25769, n25770, n25771, n25772, n25773,
         n25774, n25775, n25776, n25777, n25778, n25779, n25780, n25781,
         n25782, n25783, n25784, n25785, n25786, n25787, n25788, n25789,
         n25790, n25791, n25792, n25793, n25794, n25795, n25796, n25797,
         n25798, n25799, n25800, n25801, n25802, n25803, n25804, n25805,
         n25806, n25807, n25808, n25809, n25810, n25811, n25812, n25813,
         n25814, n25815, n25816, n25817, n25818, n25819, n25820, n25821,
         n25822, n25823, n25824, n25825, n25826, n25827, n25828, n25829,
         n25830, n25831, n25832, n25833, n25834, n25835, n25836, n25837,
         n25838, n25839, n25840, n25841, n25842, n25843, n25844, n25845,
         n25846, n25847, n25848, n25849, n25850, n25851, n25852, n25853,
         n25854, n25855, n25856, n25857, n25858, n25859, n25860, n25861,
         n25862, n25863, n25864, n25865, n25866, n25867, n25868, n25869,
         n25870, n25871, n25872, n25873, n25874, n25875, n25876, n25877,
         n25878, n25879, n25880, n25881, n25882, n25883, n25884, n25885,
         n25886, n25887, n25888, n25889, n25890, n25891, n25892, n25893,
         n25894, n25895, n25896, n25897, n25898, n25899, n25900, n25901,
         n25902, n25903, n25904, n25905, n25906, n25907, n25908, n25909,
         n25910, n25911, n25912, n25913, n25914, n25915, n25916, n25917,
         n25918, n25919, n25920, n25921, n25922, n25923, n25924, n25925,
         n25926, n25927, n25928, n25929, n25930, n25931, n25932, n25933,
         n25934, n25935, n25936, n25937, n25938, n25939, n25940, n25941,
         n25942, n25943, n25944, n25945, n25946, n25947, n25948, n25949,
         n25950, n25951, n25952, n25953, n25954, n25955, n25956, n25957,
         n25958, n25959, n25960, n25961, n25962, n25963, n25964, n25965,
         n25966, n25967, n25968, n25969, n25970, n25971, n25972, n25973,
         n25974, n25975, n25976, n25977, n25978, n25979, n25980, n25981,
         n25982, n25983, n25984, n25985, n25986, n25987, n25988, n25989,
         n25990, n25991, n25992, n25993, n25994, n25995, n25996, n25997,
         n25998, n25999, n26000, n26001, n26002, n26003, n26004, n26005,
         n26006, n26007, n26008, n26009, n26010, n26011, n26012, n26013,
         n26014, n26015, n26016, n26017, n26018, n26019, n26020, n26021,
         n26022, n26023, n26024, n26025, n26026, n26027, n26028, n26029,
         n26030, n26031, n26032, n26033, n26034, n26035, n26036, n26037,
         n26038, n26039, n26040, n26041, n26042, n26043, n26044, n26045,
         n26046, n26047, n26048, n26049, n26050, n26051, n26052, n26053,
         n26054, n26055, n26056, n26057, n26058, n26059, n26060, n26061,
         n26062, n26063, n26064, n26065, n26066, n26067, n26068, n26069,
         n26070, n26071, n26072, n26073, n26074, n26075, n26076, n26077,
         n26078, n26079, n26080, n26081, n26082, n26083, n26084, n26085,
         n26086, n26087, n26088, n26089, n26090, n26091, n26092, n26093,
         n26094, n26095, n26096, n26097, n26098, n26099, n26100, n26101,
         n26102, n26103, n26104, n26105, n26106, n26107, n26108, n26109,
         n26110, n26111, n26112, n26113, n26114, n26115, n26116, n26117,
         n26118, n26119, n26120, n26121, n26122, n26123, n26124, n26125,
         n26126, n26127, n26128, n26129, n26130, n26131, n26132, n26133,
         n26134, n26135, n26136, n26137, n26138, n26139, n26140, n26141,
         n26142, n26143, n26144, n26145, n26146, n26147, n26148, n26149,
         n26150, n26151, n26152, n26153, n26154, n26155, n26156, n26157,
         n26158, n26159, n26160, n26161, n26162, n26163, n26164, n26165,
         n26166, n26167, n26168, n26169, n26170, n26171, n26172, n26173,
         n26174, n26175, n26176, n26177, n26178, n26179, n26180, n26181,
         n26182, n26183, n26184, n26185, n26186, n26187, n26188, n26189,
         n26190, n26191, n26192, n26193, n26194, n26195, n26196, n26197,
         n26198, n26199, n26200, n26201, n26202, n26203, n26204, n26205,
         n26206, n26207, n26208, n26209, n26210, n26211, n26212, n26213,
         n26214, n26215, n26216, n26217, n26218, n26219, n26220, n26221,
         n26222, n26223, n26224, n26225, n26226, n26227, n26228, n26229,
         n26230, n26231, n26232, n26233, n26234, n26235, n26236, n26237,
         n26238, n26239, n26240, n26241, n26242, n26243, n26244, n26245,
         n26246, n26247, n26248, n26249, n26250, n26251, n26252, n26253,
         n26254, n26255, n26256, n26257, n26258, n26259, n26260, n26261,
         n26262, n26263, n26264, n26265, n26266, n26267, n26268, n26269,
         n26270, n26271, n26272, n26273, n26274, n26275, n26276, n26277,
         n26278, n26279, n26280, n26281, n26282, n26283, n26284, n26285,
         n26286, n26287, n26288, n26289, n26290, n26291, n26292, n26293,
         n26294, n26295, n26296, n26297, n26298, n26299, n26300, n26301,
         n26302, n26303, n26304, n26305, n26306, n26307, n26308, n26309,
         n26310, n26311, n26312, n26313, n26314, n26315, n26316, n26317,
         n26318, n26319, n26320, n26321, n26322, n26323, n26324, n26325,
         n26326, n26327, n26328, n26329, n26330, n26331, n26332, n26333,
         n26334, n26335, n26336, n26337, n26338, n26339, n26340, n26341,
         n26342, n26343, n26344, n26345, n26346, n26347, n26348, n26349,
         n26350, n26351, n26352, n26353, n26354, n26355, n26356, n26357,
         n26358, n26359, n26360, n26361, n26362, n26363, n26364, n26365,
         n26366, n26367, n26368, n26369, n26370, n26371, n26372, n26373,
         n26374, n26375, n26376, n26377, n26378, n26379, n26380, n26381,
         n26382, n26383, n26384, n26385, n26386, n26387, n26388, n26389,
         n26390, n26391, n26392, n26393, n26394, n26395, n26396, n26397,
         n26398, n26399, n26400, n26401, n26402, n26403, n26404, n26405,
         n26406, n26407, n26408, n26409, n26410, n26411, n26412, n26413,
         n26414, n26415, n26416, n26417, n26418, n26419, n26420, n26421,
         n26422, n26423, n26424, n26425, n26426, n26427, n26428, n26429,
         n26430, n26431, n26432, n26433, n26434, n26435, n26436, n26437,
         n26438, n26439, n26440, n26441, n26442, n26443, n26444, n26445,
         n26446, n26447, n26448, n26449, n26450, n26451, n26452, n26453,
         n26454, n26455, n26456, n26457, n26458, n26459, n26460, n26461,
         n26462, n26463, n26464, n26465, n26466, n26467, n26468, n26469,
         n26470, n26471, n26472, n26473, n26474, n26475, n26476, n26477,
         n26478, n26479, n26480, n26481, n26482, n26483, n26484, n26485,
         n26486, n26487, n26488, n26489, n26490, n26491, n26492, n26493,
         n26494, n26495, n26496, n26497, n26498, n26499, n26500, n26501,
         n26502, n26503, n26504, n26505, n26506, n26507, n26508, n26509,
         n26510, n26511, n26512, n26513, n26514, n26515, n26516, n26517,
         n26518, n26519, n26520, n26521, n26522, n26523, n26524, n26525,
         n26526, n26527, n26528, n26529, n26530, n26531, n26532, n26533,
         n26534, n26535, n26536, n26537, n26538, n26539, n26540, n26541,
         n26542, n26543, n26544, n26545, n26546, n26547, n26548, n26549,
         n26550, n26551, n26552, n26553, n26554, n26555, n26556, n26557,
         n26558, n26559, n26560, n26561, n26562, n26563, n26564, n26565,
         n26566, n26567, n26568, n26569, n26570, n26571, n26572, n26573,
         n26574, n26575, n26576, n26577, n26578, n26579, n26580, n26581,
         n26582, n26583, n26584, n26585, n26586, n26587, n26588, n26589,
         n26590, n26591, n26592, n26593, n26594, n26595, n26596, n26597,
         n26598, n26599, n26600, n26601, n26602, n26603, n26604, n26605,
         n26606, n26607, n26608, n26609, n26610, n26611, n26612, n26613,
         n26614, n26615, n26616, n26617, n26618, n26619, n26620, n26621,
         n26622, n26623, n26624, n26625, n26626, n26627, n26628, n26629,
         n26630, n26631, n26632, n26633, n26634, n26635, n26636, n26637,
         n26638, n26639, n26640, n26641, n26642, n26643, n26644, n26645,
         n26646, n26647, n26648, n26649, n26650, n26651, n26652, n26653,
         n26654, n26655, n26656, n26657, n26658, n26659, n26660, n26661,
         n26662, n26663, n26664, n26665, n26666, n26667, n26668, n26669,
         n26670, n26671, n26672, n26673, n26674, n26675, n26676, n26677,
         n26678, n26679, n26680, n26681, n26682, n26683, n26684, n26685,
         n26686, n26687, n26688, n26689, n26690, n26691, n26692, n26693,
         n26694, n26695, n26696, n26697, n26698, n26699, n26700, n26701,
         n26702, n26703, n26704, n26705, n26706, n26707, n26708, n26709,
         n26710, n26711, n26712, n26713, n26714, n26715, n26716, n26717,
         n26718, n26719, n26720, n26721, n26722, n26723, n26724, n26725,
         n26726, n26727, n26728, n26729, n26730, n26731, n26732, n26733,
         n26734, n26735, n26736, n26737, n26738, n26739, n26740, n26741,
         n26742, n26743, n26744, n26745, n26746, n26747, n26748, n26749,
         n26750, n26751, n26752, n26753, n26754, n26755, n26756, n26757,
         n26758, n26759, n26760, n26761, n26762, n26763, n26764, n26765,
         n26766, n26767, n26768, n26769, n26770, n26771, n26772, n26773,
         n26774, n26775, n26776, n26777, n26778, n26779, n26780, n26781,
         n26782, n26783, n26784, n26785, n26786, n26787, n26788, n26789,
         n26790, n26791, n26792, n26793, n26794, n26795, n26796, n26797,
         n26798, n26799, n26800, n26801, n26802, n26803, n26804, n26805,
         n26806, n26807, n26808, n26809, n26810, n26811, n26812, n26813,
         n26814, n26815, n26816, n26817, n26818, n26819, n26820, n26821,
         n26822, n26823, n26824, n26825, n26826, n26827, n26828, n26829,
         n26830, n26831, n26832, n26833, n26834, n26835, n26836, n26837,
         n26838, n26839, n26840, n26841, n26842, n26843, n26844, n26845,
         n26846, n26847, n26848, n26849, n26850, n26851, n26852, n26853,
         n26854, n26855, n26856, n26857, n26858, n26859, n26860, n26861,
         n26862, n26863, n26864, n26865, n26866, n26867, n26868, n26869,
         n26870, n26871, n26872, n26873, n26874, n26875, n26876, n26877,
         n26878, n26879, n26880, n26881, n26882, n26883, n26884, n26885,
         n26886, n26887, n26888, n26889, n26890, n26891, n26892, n26893,
         n26894, n26895, n26896, n26897, n26898, n26899, n26900, n26901,
         n26902, n26903, n26904, n26905, n26906, n26907, n26908, n26909,
         n26910, n26911, n26912, n26913, n26914, n26915, n26916, n26917,
         n26918, n26919, n26920, n26921, n26922, n26923, n26924, n26925,
         n26926, n26927, n26928, n26929, n26930, n26931, n26932, n26933,
         n26934, n26935, n26936, n26937, n26938, n26939, n26940, n26941,
         n26942, n26943, n26944, n26945, n26946, n26947, n26948, n26949,
         n26950, n26951, n26952, n26953, n26954, n26955, n26956, n26957,
         n26958, n26959, n26960, n26961, n26962, n26963, n26964, n26965,
         n26966, n26967, n26968, n26969, n26970, n26971, n26972, n26973,
         n26974, n26975, n26976, n26977, n26978, n26979, n26980, n26981,
         n26982, n26983, n26984, n26985, n26986, n26987, n26988, n26989,
         n26990, n26991, n26992, n26993, n26994, n26995, n26996, n26997,
         n26998, n26999, n27000, n27001, n27002, n27003, n27004, n27005,
         n27006, n27007, n27008, n27009, n27010, n27011, n27012, n27013,
         n27014, n27015, n27016, n27017, n27018, n27019, n27020, n27021,
         n27022, n27023, n27024, n27025, n27026, n27027, n27028, n27029,
         n27030, n27031, n27032, n27033, n27034, n27035, n27036, n27037,
         n27038, n27039, n27040, n27041, n27042, n27043, n27044, n27045,
         n27046, n27047, n27048, n27049, n27050, n27051, n27052, n27053,
         n27054, n27055, n27056, n27057, n27058, n27059, n27060, n27061,
         n27062, n27063, n27064, n27065, n27066, n27067, n27068, n27069,
         n27070, n27071, n27072, n27073, n27074, n27075, n27076, n27077,
         n27078, n27079, n27080, n27081, n27082, n27083, n27084, n27085,
         n27086, n27087, n27088, n27089, n27090, n27091, n27092, n27093,
         n27094, n27095, n27096, n27097, n27098, n27099, n27100, n27101,
         n27102, n27103, n27104, n27105, n27106, n27107, n27108, n27109,
         n27110, n27111, n27112, n27113, n27114, n27115, n27116, n27117,
         n27118, n27119, n27120, n27121, n27122, n27123, n27124, n27125,
         n27126, n27127, n27128, n27129, n27130, n27131, n27132, n27133,
         n27134, n27135, n27136, n27137, n27138, n27139, n27140, n27141,
         n27142, n27143, n27144, n27145, n27146, n27147, n27148, n27149,
         n27150, n27151, n27152, n27153, n27154, n27155, n27156, n27157,
         n27158, n27159, n27160, n27161, n27162, n27163, n27164, n27165,
         n27166, n27167, n27168, n27169, n27170, n27171, n27172, n27173,
         n27174, n27175, n27176, n27177, n27178, n27179, n27180, n27181,
         n27182, n27183, n27184, n27185, n27186, n27187, n27188, n27189,
         n27190, n27191, n27192, n27193, n27194, n27195, n27196, n27197,
         n27198, n27199, n27200, n27201, n27202, n27203, n27204, n27205,
         n27206, n27207, n27208, n27209, n27210, n27211, n27212, n27213,
         n27214, n27215, n27216, n27217, n27218, n27219, n27220, n27221,
         n27222, n27223, n27224, n27225, n27226, n27227, n27228, n27229,
         n27230, n27231, n27232, n27233, n27234, n27235, n27236, n27237,
         n27238, n27239, n27240, n27241, n27242, n27243, n27244, n27245,
         n27246, n27247, n27248, n27249, n27250, n27251, n27252, n27253,
         n27254, n27255, n27256, n27257, n27258, n27259, n27260, n27261,
         n27262, n27263, n27264, n27265, n27266, n27267, n27268, n27269,
         n27270, n27271, n27272, n27273, n27274, n27275, n27276, n27277,
         n27278, n27279, n27280, n27281, n27282, n27283, n27284, n27285,
         n27286, n27287, n27288, n27289, n27290, n27291, n27292, n27293,
         n27294, n27295, n27296, n27297, n27298, n27299, n27300, n27301,
         n27302, n27303, n27304, n27305, n27306, n27307, n27308, n27309,
         n27310, n27311, n27312, n27313, n27314, n27315, n27316, n27317,
         n27318, n27319, n27320, n27321, n27322, n27323, n27324, n27325,
         n27326, n27327, n27328, n27329, n27330, n27331, n27332, n27333,
         n27334, n27335, n27336, n27337, n27338, n27339, n27340, n27341,
         n27342, n27343, n27344, n27345, n27346, n27347, n27348, n27349,
         n27350, n27351, n27352, n27353, n27354, n27355, n27356, n27357,
         n27358, n27359, n27360, n27361, n27362, n27363, n27364, n27365,
         n27366, n27367, n27368, n27369, n27370, n27371, n27372, n27373,
         n27374, n27375, n27376, n27377, n27378, n27379, n27380, n27381,
         n27382, n27383, n27384, n27385, n27386, n27387, n27388, n27389,
         n27390, n27391, n27392, n27393, n27394, n27395, n27396, n27397,
         n27398, n27399, n27400, n27401, n27402, n27403, n27404, n27405,
         n27406, n27407, n27408, n27409, n27410, n27411, n27412, n27413,
         n27414, n27415, n27416, n27417, n27418, n27419, n27420, n27421,
         n27422, n27423, n27424, n27425, n27426, n27427, n27428, n27429,
         n27430, n27431, n27432, n27433, n27434, n27435, n27436, n27437,
         n27438, n27439, n27440, n27441, n27442, n27443, n27444, n27445,
         n27446, n27447, n27448, n27449, n27450, n27451, n27452, n27453,
         n27454, n27455, n27456, n27457, n27458, n27459, n27460, n27461,
         n27462, n27463, n27464, n27465, n27466, n27467, n27468, n27469,
         n27470, n27471, n27472, n27473, n27474, n27475, n27476, n27477,
         n27478, n27479, n27480, n27481, n27482, n27483, n27484, n27485,
         n27486, n27487, n27488, n27489, n27490, n27491, n27492, n27493,
         n27494, n27495, n27496, n27497, n27498, n27499, n27500, n27501,
         n27502, n27503, n27504, n27505, n27506, n27507, n27508, n27509,
         n27510, n27511, n27512, n27513, n27514, n27515, n27516, n27517,
         n27518, n27519, n27520, n27521, n27522, n27523, n27524, n27525,
         n27526, n27527, n27528, n27529, n27530, n27531, n27532, n27533,
         n27534, n27535, n27536, n27537, n27538, n27539, n27540, n27541,
         n27542, n27543, n27544, n27545, n27546, n27547, n27548, n27549,
         n27550, n27551, n27552, n27553, n27554, n27555, n27556, n27557,
         n27558, n27559, n27560, n27561, n27562, n27563, n27564, n27565,
         n27566, n27567, n27568, n27569, n27570, n27571, n27572, n27573,
         n27574, n27575, n27576, n27577, n27578, n27579, n27580, n27581,
         n27582, n27583, n27584, n27585, n27586, n27587, n27588, n27589,
         n27590, n27591, n27592, n27593, n27594, n27595, n27596, n27597,
         n27598, n27599, n27600, n27601, n27602, n27603, n27604, n27605,
         n27606, n27607, n27608, n27609, n27610, n27611, n27612, n27613,
         n27614, n27615, n27616, n27617, n27618, n27619, n27620, n27621,
         n27622, n27623, n27624, n27625, n27626, n27627, n27628, n27629,
         n27630, n27631, n27632, n27633, n27634, n27635, n27636, n27637,
         n27638, n27639, n27640, n27641, n27642, n27643, n27644, n27645,
         n27646, n27647, n27648, n27649, n27650, n27651, n27652, n27653,
         n27654, n27655, n27656, n27657, n27658, n27659, n27660, n27661,
         n27662, n27663, n27664, n27665, n27666, n27667, n27668, n27669,
         n27670, n27671, n27672, n27673, n27674, n27675, n27676, n27677,
         n27678, n27679, n27680, n27681, n27682, n27683, n27684, n27685,
         n27686, n27687, n27688, n27689, n27690, n27691, n27692, n27693,
         n27694, n27695, n27696, n27697, n27698, n27699, n27700, n27701,
         n27702, n27703, n27704, n27705, n27706, n27707, n27708, n27709,
         n27710, n27711, n27712, n27713, n27714, n27715, n27716, n27717,
         n27718, n27719, n27720, n27721, n27722, n27723, n27724, n27725,
         n27726, n27727, n27728, n27729, n27730, n27731, n27732, n27733,
         n27734, n27735, n27736, n27737, n27738, n27739, n27740, n27741,
         n27742, n27743, n27744, n27745, n27746, n27747, n27748, n27749,
         n27750, n27751, n27752, n27753, n27754, n27755, n27756, n27757,
         n27758, n27759, n27760, n27761, n27762, n27763, n27764, n27765,
         n27766, n27767, n27768, n27769, n27770, n27771, n27772, n27773,
         n27774, n27775, n27776, n27777, n27778, n27779, n27780, n27781,
         n27782, n27783, n27784, n27785, n27786, n27787, n27788, n27789,
         n27790, n27791, n27792, n27793, n27794, n27795, n27796, n27797,
         n27798, n27799, n27800, n27801, n27802, n27803, n27804, n27805,
         n27806, n27807, n27808, n27809, n27810, n27811, n27812, n27813,
         n27814, n27815, n27816, n27817, n27818, n27819, n27820, n27821,
         n27822, n27823, n27824, n27825, n27826, n27827, n27828, n27829,
         n27830, n27831, n27832, n27833, n27834, n27835, n27836, n27837,
         n27838, n27839, n27840, n27841, n27842, n27843, n27844, n27845,
         n27846, n27847, n27848, n27849, n27850, n27851, n27852, n27853,
         n27854, n27855, n27856, n27857, n27858, n27859, n27860, n27861,
         n27862, n27863, n27864, n27865, n27866, n27867, n27868, n27869,
         n27870, n27871, n27872, n27873, n27874, n27875, n27876, n27877,
         n27878, n27879, n27880, n27881, n27882, n27883, n27884, n27885,
         n27886, n27887, n27888, n27889, n27890, n27891, n27892, n27893,
         n27894, n27895, n27896, n27897, n27898, n27899, n27900, n27901,
         n27902, n27903, n27904, n27905, n27906, n27907, n27908, n27909,
         n27910, n27911, n27912, n27913, n27914, n27915, n27916, n27917,
         n27918, n27919, n27920, n27921, n27922, n27923, n27924, n27925,
         n27926, n27927, n27928, n27929, n27930, n27931, n27932, n27933,
         n27934, n27935, n27936, n27937, n27938, n27939, n27940, n27941,
         n27942, n27943, n27944, n27945, n27946, n27947, n27948, n27949,
         n27950, n27951, n27952, n27953, n27954, n27955, n27956, n27957,
         n27958, n27959, n27960, n27961, n27962, n27963, n27964, n27965,
         n27966, n27967, n27968, n27969, n27970, n27971, n27972, n27973,
         n27974, n27975, n27976, n27977, n27978, n27979, n27980, n27981,
         n27982, n27983, n27984, n27985, n27986, n27987, n27988, n27989,
         n27990, n27991, n27992, n27993, n27994, n27995, n27996, n27997,
         n27998, n27999, n28000, n28001, n28002, n28003, n28004, n28005,
         n28006, n28007, n28008, n28009, n28010, n28011, n28012, n28013,
         n28014, n28015, n28016, n28017, n28018, n28019, n28020, n28021,
         n28022, n28023, n28024, n28025, n28026, n28027, n28028, n28029,
         n28030, n28031, n28032, n28033, n28034, n28035, n28036, n28037,
         n28038, n28039, n28040, n28041, n28042, n28043, n28044, n28045,
         n28046, n28047, n28048, n28049, n28050, n28051, n28052, n28053,
         n28054, n28055, n28056, n28057, n28058, n28059, n28060, n28061,
         n28062, n28063, n28064, n28065, n28066, n28067, n28068, n28069,
         n28070, n28071, n28072, n28073, n28074, n28075, n28076, n28077,
         n28078, n28079, n28080, n28081, n28082, n28083, n28084, n28085,
         n28086, n28087, n28088, n28089, n28090, n28091, n28092, n28093,
         n28094, n28095, n28096, n28097, n28098, n28099, n28100, n28101,
         n28102, n28103, n28104, n28105, n28106, n28107, n28108, n28109,
         n28110, n28111, n28112, n28113, n28114, n28115, n28116, n28117,
         n28118, n28119, n28120, n28121, n28122, n28123, n28124, n28125,
         n28126, n28127, n28128, n28129, n28130, n28131, n28132, n28133,
         n28134, n28135, n28136, n28137, n28138, n28139, n28140, n28141,
         n28142, n28143, n28144, n28145, n28146, n28147, n28148, n28149,
         n28150, n28151, n28152, n28153, n28154, n28155, n28156, n28157,
         n28158, n28159, n28160, n28161, n28162, n28163, n28164, n28165,
         n28166, n28167, n28168, n28169, n28170, n28171, n28172, n28173,
         n28174, n28175, n28176, n28177, n28178, n28179, n28180, n28181,
         n28182, n28183, n28184, n28185, n28186, n28187, n28188, n28189,
         n28190, n28191, n28192, n28193, n28194, n28195, n28196, n28197,
         n28198, n28199, n28200, n28201, n28202, n28203, n28204, n28205,
         n28206, n28207, n28208, n28209, n28210, n28211, n28212, n28213,
         n28214, n28215, n28216, n28217, n28218, n28219, n28220, n28221,
         n28222, n28223, n28224, n28225, n28226, n28227, n28228, n28229,
         n28230, n28231, n28232, n28233, n28234, n28235, n28236, n28237,
         n28238, n28239, n28240, n28241, n28242, n28243, n28244, n28245,
         n28246, n28247, n28248, n28249, n28250, n28251, n28252, n28253,
         n28254, n28255, n28256, n28257, n28258, n28259, n28260, n28261,
         n28262, n28263, n28264, n28265, n28266, n28267, n28268, n28269,
         n28270, n28271, n28272, n28273, n28274, n28275, n28276, n28277,
         n28278, n28279, n28280, n28281, n28282, n28283, n28284, n28285,
         n28286, n28287, n28288, n28289, n28290, n28291, n28292, n28293,
         n28294, n28295, n28296, n28297, n28298, n28299, n28300, n28301,
         n28302, n28303, n28304, n28305, n28306, n28307, n28308, n28309,
         n28310, n28311, n28312, n28313, n28314, n28315, n28316, n28317,
         n28318, n28319, n28320, n28321, n28322, n28323, n28324, n28325,
         n28326, n28327, n28328, n28329, n28330, n28331, n28332, n28333,
         n28334, n28335, n28336, n28337, n28338, n28339, n28340, n28341,
         n28342, n28343, n28344, n28345, n28346, n28347, n28348, n28349,
         n28350, n28351, n28352, n28353, n28354, n28355, n28356, n28357,
         n28358, n28359, n28360, n28361, n28362, n28363, n28364, n28365,
         n28366, n28367, n28368, n28369, n28370, n28371, n28372, n28373,
         n28374, n28375, n28376, n28377, n28378, n28379, n28380, n28381,
         n28382, n28383, n28384, n28385, n28386, n28387, n28388, n28389,
         n28390, n28391, n28392, n28393, n28394, n28395, n28396, n28397,
         n28398, n28399, n28400, n28401, n28402, n28403, n28404, n28405,
         n28406, n28407, n28408, n28409, n28410, n28411, n28412, n28413,
         n28414, n28415, n28416, n28417, n28418, n28419, n28420, n28421,
         n28422, n28423, n28424, n28425, n28426, n28427, n28428, n28429,
         n28430, n28431, n28432, n28433, n28434, n28435, n28436, n28437,
         n28438, n28439, n28440, n28441, n28442, n28443, n28444, n28445,
         n28446, n28447, n28448, n28449, n28450, n28451, n28452, n28453,
         n28454, n28455, n28456, n28457, n28458, n28459, n28460, n28461,
         n28462, n28463, n28464, n28465, n28466, n28467, n28468, n28469,
         n28470, n28471, n28472, n28473, n28474, n28475, n28476, n28477,
         n28478, n28479, n28480, n28481, n28482, n28483, n28484, n28485,
         n28486, n28487, n28488, n28489, n28490, n28491, n28492, n28493,
         n28494, n28495, n28496, n28497, n28498, n28499, n28500, n28501,
         n28502, n28503, n28504, n28505, n28506, n28507, n28508, n28509,
         n28510, n28511, n28512, n28513, n28514, n28515, n28516, n28517,
         n28518, n28519, n28520, n28521, n28522, n28523, n28524, n28525,
         n28526, n28527, n28528, n28529, n28530, n28531, n28532, n28533,
         n28534, n28535, n28536, n28537, n28538, n28539, n28540, n28541,
         n28542, n28543, n28544, n28545, n28546, n28547, n28548, n28549,
         n28550, n28551, n28552, n28553, n28554, n28555, n28556, n28557,
         n28558, n28559, n28560, n28561, n28562, n28563, n28564, n28565,
         n28566, n28567, n28568, n28569, n28570, n28571, n28572, n28573,
         n28574, n28575, n28576, n28577, n28578, n28579, n28580, n28581,
         n28582, n28583, n28584, n28585, n28586, n28587, n28588, n28589,
         n28590, n28591, n28592, n28593, n28594, n28595, n28596, n28597,
         n28598, n28599, n28600, n28601, n28602, n28603, n28604, n28605,
         n28606, n28607, n28608, n28609, n28610, n28611, n28612, n28613,
         n28614, n28615, n28616, n28617, n28618, n28619, n28620, n28621,
         n28622, n28623, n28624, n28625, n28626, n28627, n28628, n28629,
         n28630, n28631, n28632, n28633, n28634, n28635, n28636, n28637,
         n28638, n28639, n28640, n28641, n28642, n28643, n28644, n28645,
         n28646, n28647, n28648, n28649, n28650, n28651, n28652, n28653,
         n28654, n28655, n28656, n28657, n28658, n28659, n28660, n28661,
         n28662, n28663, n28664, n28665, n28666, n28667, n28668, n28669,
         n28670, n28671, n28672, n28673, n28674, n28675, n28676, n28677,
         n28678, n28679, n28680, n28681, n28682, n28683, n28684, n28685,
         n28686, n28687, n28688, n28689, n28690, n28691, n28692, n28693,
         n28694, n28695, n28696, n28697, n28698, n28699, n28700, n28701,
         n28702, n28703, n28704, n28705, n28706;
  wire   [1023:0] start_in;
  wire   [1023:0] start_reg;
  wire   [1023:0] ereg;
  wire   [1023:0] o;
  wire   [1023:0] creg;
  wire   [1023:0] x;
  wire   [1023:0] y;

  DFF init_reg ( .D(1'b1), .CLK(clk), .RST(rst), .Q(init) );
  DFF \start_reg_reg[0]  ( .D(start_in[1023]), .CLK(clk), .RST(rst), .Q(
        start_reg[0]) );
  DFF \start_reg_reg[1]  ( .D(start_in[0]), .CLK(clk), .RST(rst), .Q(
        start_reg[1]) );
  DFF \start_reg_reg[2]  ( .D(start_in[1]), .CLK(clk), .RST(rst), .Q(
        start_reg[2]) );
  DFF \start_reg_reg[3]  ( .D(start_in[2]), .CLK(clk), .RST(rst), .Q(
        start_reg[3]) );
  DFF \start_reg_reg[4]  ( .D(start_in[3]), .CLK(clk), .RST(rst), .Q(
        start_reg[4]) );
  DFF \start_reg_reg[5]  ( .D(start_in[4]), .CLK(clk), .RST(rst), .Q(
        start_reg[5]) );
  DFF \start_reg_reg[6]  ( .D(start_in[5]), .CLK(clk), .RST(rst), .Q(
        start_reg[6]) );
  DFF \start_reg_reg[7]  ( .D(start_in[6]), .CLK(clk), .RST(rst), .Q(
        start_reg[7]) );
  DFF \start_reg_reg[8]  ( .D(start_in[7]), .CLK(clk), .RST(rst), .Q(
        start_reg[8]) );
  DFF \start_reg_reg[9]  ( .D(start_in[8]), .CLK(clk), .RST(rst), .Q(
        start_reg[9]) );
  DFF \start_reg_reg[10]  ( .D(start_in[9]), .CLK(clk), .RST(rst), .Q(
        start_reg[10]) );
  DFF \start_reg_reg[11]  ( .D(start_in[10]), .CLK(clk), .RST(rst), .Q(
        start_reg[11]) );
  DFF \start_reg_reg[12]  ( .D(start_in[11]), .CLK(clk), .RST(rst), .Q(
        start_reg[12]) );
  DFF \start_reg_reg[13]  ( .D(start_in[12]), .CLK(clk), .RST(rst), .Q(
        start_reg[13]) );
  DFF \start_reg_reg[14]  ( .D(start_in[13]), .CLK(clk), .RST(rst), .Q(
        start_reg[14]) );
  DFF \start_reg_reg[15]  ( .D(start_in[14]), .CLK(clk), .RST(rst), .Q(
        start_reg[15]) );
  DFF \start_reg_reg[16]  ( .D(start_in[15]), .CLK(clk), .RST(rst), .Q(
        start_reg[16]) );
  DFF \start_reg_reg[17]  ( .D(start_in[16]), .CLK(clk), .RST(rst), .Q(
        start_reg[17]) );
  DFF \start_reg_reg[18]  ( .D(start_in[17]), .CLK(clk), .RST(rst), .Q(
        start_reg[18]) );
  DFF \start_reg_reg[19]  ( .D(start_in[18]), .CLK(clk), .RST(rst), .Q(
        start_reg[19]) );
  DFF \start_reg_reg[20]  ( .D(start_in[19]), .CLK(clk), .RST(rst), .Q(
        start_reg[20]) );
  DFF \start_reg_reg[21]  ( .D(start_in[20]), .CLK(clk), .RST(rst), .Q(
        start_reg[21]) );
  DFF \start_reg_reg[22]  ( .D(start_in[21]), .CLK(clk), .RST(rst), .Q(
        start_reg[22]) );
  DFF \start_reg_reg[23]  ( .D(start_in[22]), .CLK(clk), .RST(rst), .Q(
        start_reg[23]) );
  DFF \start_reg_reg[24]  ( .D(start_in[23]), .CLK(clk), .RST(rst), .Q(
        start_reg[24]) );
  DFF \start_reg_reg[25]  ( .D(start_in[24]), .CLK(clk), .RST(rst), .Q(
        start_reg[25]) );
  DFF \start_reg_reg[26]  ( .D(start_in[25]), .CLK(clk), .RST(rst), .Q(
        start_reg[26]) );
  DFF \start_reg_reg[27]  ( .D(start_in[26]), .CLK(clk), .RST(rst), .Q(
        start_reg[27]) );
  DFF \start_reg_reg[28]  ( .D(start_in[27]), .CLK(clk), .RST(rst), .Q(
        start_reg[28]) );
  DFF \start_reg_reg[29]  ( .D(start_in[28]), .CLK(clk), .RST(rst), .Q(
        start_reg[29]) );
  DFF \start_reg_reg[30]  ( .D(start_in[29]), .CLK(clk), .RST(rst), .Q(
        start_reg[30]) );
  DFF \start_reg_reg[31]  ( .D(start_in[30]), .CLK(clk), .RST(rst), .Q(
        start_reg[31]) );
  DFF \start_reg_reg[32]  ( .D(start_in[31]), .CLK(clk), .RST(rst), .Q(
        start_reg[32]) );
  DFF \start_reg_reg[33]  ( .D(start_in[32]), .CLK(clk), .RST(rst), .Q(
        start_reg[33]) );
  DFF \start_reg_reg[34]  ( .D(start_in[33]), .CLK(clk), .RST(rst), .Q(
        start_reg[34]) );
  DFF \start_reg_reg[35]  ( .D(start_in[34]), .CLK(clk), .RST(rst), .Q(
        start_reg[35]) );
  DFF \start_reg_reg[36]  ( .D(start_in[35]), .CLK(clk), .RST(rst), .Q(
        start_reg[36]) );
  DFF \start_reg_reg[37]  ( .D(start_in[36]), .CLK(clk), .RST(rst), .Q(
        start_reg[37]) );
  DFF \start_reg_reg[38]  ( .D(start_in[37]), .CLK(clk), .RST(rst), .Q(
        start_reg[38]) );
  DFF \start_reg_reg[39]  ( .D(start_in[38]), .CLK(clk), .RST(rst), .Q(
        start_reg[39]) );
  DFF \start_reg_reg[40]  ( .D(start_in[39]), .CLK(clk), .RST(rst), .Q(
        start_reg[40]) );
  DFF \start_reg_reg[41]  ( .D(start_in[40]), .CLK(clk), .RST(rst), .Q(
        start_reg[41]) );
  DFF \start_reg_reg[42]  ( .D(start_in[41]), .CLK(clk), .RST(rst), .Q(
        start_reg[42]) );
  DFF \start_reg_reg[43]  ( .D(start_in[42]), .CLK(clk), .RST(rst), .Q(
        start_reg[43]) );
  DFF \start_reg_reg[44]  ( .D(start_in[43]), .CLK(clk), .RST(rst), .Q(
        start_reg[44]) );
  DFF \start_reg_reg[45]  ( .D(start_in[44]), .CLK(clk), .RST(rst), .Q(
        start_reg[45]) );
  DFF \start_reg_reg[46]  ( .D(start_in[45]), .CLK(clk), .RST(rst), .Q(
        start_reg[46]) );
  DFF \start_reg_reg[47]  ( .D(start_in[46]), .CLK(clk), .RST(rst), .Q(
        start_reg[47]) );
  DFF \start_reg_reg[48]  ( .D(start_in[47]), .CLK(clk), .RST(rst), .Q(
        start_reg[48]) );
  DFF \start_reg_reg[49]  ( .D(start_in[48]), .CLK(clk), .RST(rst), .Q(
        start_reg[49]) );
  DFF \start_reg_reg[50]  ( .D(start_in[49]), .CLK(clk), .RST(rst), .Q(
        start_reg[50]) );
  DFF \start_reg_reg[51]  ( .D(start_in[50]), .CLK(clk), .RST(rst), .Q(
        start_reg[51]) );
  DFF \start_reg_reg[52]  ( .D(start_in[51]), .CLK(clk), .RST(rst), .Q(
        start_reg[52]) );
  DFF \start_reg_reg[53]  ( .D(start_in[52]), .CLK(clk), .RST(rst), .Q(
        start_reg[53]) );
  DFF \start_reg_reg[54]  ( .D(start_in[53]), .CLK(clk), .RST(rst), .Q(
        start_reg[54]) );
  DFF \start_reg_reg[55]  ( .D(start_in[54]), .CLK(clk), .RST(rst), .Q(
        start_reg[55]) );
  DFF \start_reg_reg[56]  ( .D(start_in[55]), .CLK(clk), .RST(rst), .Q(
        start_reg[56]) );
  DFF \start_reg_reg[57]  ( .D(start_in[56]), .CLK(clk), .RST(rst), .Q(
        start_reg[57]) );
  DFF \start_reg_reg[58]  ( .D(start_in[57]), .CLK(clk), .RST(rst), .Q(
        start_reg[58]) );
  DFF \start_reg_reg[59]  ( .D(start_in[58]), .CLK(clk), .RST(rst), .Q(
        start_reg[59]) );
  DFF \start_reg_reg[60]  ( .D(start_in[59]), .CLK(clk), .RST(rst), .Q(
        start_reg[60]) );
  DFF \start_reg_reg[61]  ( .D(start_in[60]), .CLK(clk), .RST(rst), .Q(
        start_reg[61]) );
  DFF \start_reg_reg[62]  ( .D(start_in[61]), .CLK(clk), .RST(rst), .Q(
        start_reg[62]) );
  DFF \start_reg_reg[63]  ( .D(start_in[62]), .CLK(clk), .RST(rst), .Q(
        start_reg[63]) );
  DFF \start_reg_reg[64]  ( .D(start_in[63]), .CLK(clk), .RST(rst), .Q(
        start_reg[64]) );
  DFF \start_reg_reg[65]  ( .D(start_in[64]), .CLK(clk), .RST(rst), .Q(
        start_reg[65]) );
  DFF \start_reg_reg[66]  ( .D(start_in[65]), .CLK(clk), .RST(rst), .Q(
        start_reg[66]) );
  DFF \start_reg_reg[67]  ( .D(start_in[66]), .CLK(clk), .RST(rst), .Q(
        start_reg[67]) );
  DFF \start_reg_reg[68]  ( .D(start_in[67]), .CLK(clk), .RST(rst), .Q(
        start_reg[68]) );
  DFF \start_reg_reg[69]  ( .D(start_in[68]), .CLK(clk), .RST(rst), .Q(
        start_reg[69]) );
  DFF \start_reg_reg[70]  ( .D(start_in[69]), .CLK(clk), .RST(rst), .Q(
        start_reg[70]) );
  DFF \start_reg_reg[71]  ( .D(start_in[70]), .CLK(clk), .RST(rst), .Q(
        start_reg[71]) );
  DFF \start_reg_reg[72]  ( .D(start_in[71]), .CLK(clk), .RST(rst), .Q(
        start_reg[72]) );
  DFF \start_reg_reg[73]  ( .D(start_in[72]), .CLK(clk), .RST(rst), .Q(
        start_reg[73]) );
  DFF \start_reg_reg[74]  ( .D(start_in[73]), .CLK(clk), .RST(rst), .Q(
        start_reg[74]) );
  DFF \start_reg_reg[75]  ( .D(start_in[74]), .CLK(clk), .RST(rst), .Q(
        start_reg[75]) );
  DFF \start_reg_reg[76]  ( .D(start_in[75]), .CLK(clk), .RST(rst), .Q(
        start_reg[76]) );
  DFF \start_reg_reg[77]  ( .D(start_in[76]), .CLK(clk), .RST(rst), .Q(
        start_reg[77]) );
  DFF \start_reg_reg[78]  ( .D(start_in[77]), .CLK(clk), .RST(rst), .Q(
        start_reg[78]) );
  DFF \start_reg_reg[79]  ( .D(start_in[78]), .CLK(clk), .RST(rst), .Q(
        start_reg[79]) );
  DFF \start_reg_reg[80]  ( .D(start_in[79]), .CLK(clk), .RST(rst), .Q(
        start_reg[80]) );
  DFF \start_reg_reg[81]  ( .D(start_in[80]), .CLK(clk), .RST(rst), .Q(
        start_reg[81]) );
  DFF \start_reg_reg[82]  ( .D(start_in[81]), .CLK(clk), .RST(rst), .Q(
        start_reg[82]) );
  DFF \start_reg_reg[83]  ( .D(start_in[82]), .CLK(clk), .RST(rst), .Q(
        start_reg[83]) );
  DFF \start_reg_reg[84]  ( .D(start_in[83]), .CLK(clk), .RST(rst), .Q(
        start_reg[84]) );
  DFF \start_reg_reg[85]  ( .D(start_in[84]), .CLK(clk), .RST(rst), .Q(
        start_reg[85]) );
  DFF \start_reg_reg[86]  ( .D(start_in[85]), .CLK(clk), .RST(rst), .Q(
        start_reg[86]) );
  DFF \start_reg_reg[87]  ( .D(start_in[86]), .CLK(clk), .RST(rst), .Q(
        start_reg[87]) );
  DFF \start_reg_reg[88]  ( .D(start_in[87]), .CLK(clk), .RST(rst), .Q(
        start_reg[88]) );
  DFF \start_reg_reg[89]  ( .D(start_in[88]), .CLK(clk), .RST(rst), .Q(
        start_reg[89]) );
  DFF \start_reg_reg[90]  ( .D(start_in[89]), .CLK(clk), .RST(rst), .Q(
        start_reg[90]) );
  DFF \start_reg_reg[91]  ( .D(start_in[90]), .CLK(clk), .RST(rst), .Q(
        start_reg[91]) );
  DFF \start_reg_reg[92]  ( .D(start_in[91]), .CLK(clk), .RST(rst), .Q(
        start_reg[92]) );
  DFF \start_reg_reg[93]  ( .D(start_in[92]), .CLK(clk), .RST(rst), .Q(
        start_reg[93]) );
  DFF \start_reg_reg[94]  ( .D(start_in[93]), .CLK(clk), .RST(rst), .Q(
        start_reg[94]) );
  DFF \start_reg_reg[95]  ( .D(start_in[94]), .CLK(clk), .RST(rst), .Q(
        start_reg[95]) );
  DFF \start_reg_reg[96]  ( .D(start_in[95]), .CLK(clk), .RST(rst), .Q(
        start_reg[96]) );
  DFF \start_reg_reg[97]  ( .D(start_in[96]), .CLK(clk), .RST(rst), .Q(
        start_reg[97]) );
  DFF \start_reg_reg[98]  ( .D(start_in[97]), .CLK(clk), .RST(rst), .Q(
        start_reg[98]) );
  DFF \start_reg_reg[99]  ( .D(start_in[98]), .CLK(clk), .RST(rst), .Q(
        start_reg[99]) );
  DFF \start_reg_reg[100]  ( .D(start_in[99]), .CLK(clk), .RST(rst), .Q(
        start_reg[100]) );
  DFF \start_reg_reg[101]  ( .D(start_in[100]), .CLK(clk), .RST(rst), .Q(
        start_reg[101]) );
  DFF \start_reg_reg[102]  ( .D(start_in[101]), .CLK(clk), .RST(rst), .Q(
        start_reg[102]) );
  DFF \start_reg_reg[103]  ( .D(start_in[102]), .CLK(clk), .RST(rst), .Q(
        start_reg[103]) );
  DFF \start_reg_reg[104]  ( .D(start_in[103]), .CLK(clk), .RST(rst), .Q(
        start_reg[104]) );
  DFF \start_reg_reg[105]  ( .D(start_in[104]), .CLK(clk), .RST(rst), .Q(
        start_reg[105]) );
  DFF \start_reg_reg[106]  ( .D(start_in[105]), .CLK(clk), .RST(rst), .Q(
        start_reg[106]) );
  DFF \start_reg_reg[107]  ( .D(start_in[106]), .CLK(clk), .RST(rst), .Q(
        start_reg[107]) );
  DFF \start_reg_reg[108]  ( .D(start_in[107]), .CLK(clk), .RST(rst), .Q(
        start_reg[108]) );
  DFF \start_reg_reg[109]  ( .D(start_in[108]), .CLK(clk), .RST(rst), .Q(
        start_reg[109]) );
  DFF \start_reg_reg[110]  ( .D(start_in[109]), .CLK(clk), .RST(rst), .Q(
        start_reg[110]) );
  DFF \start_reg_reg[111]  ( .D(start_in[110]), .CLK(clk), .RST(rst), .Q(
        start_reg[111]) );
  DFF \start_reg_reg[112]  ( .D(start_in[111]), .CLK(clk), .RST(rst), .Q(
        start_reg[112]) );
  DFF \start_reg_reg[113]  ( .D(start_in[112]), .CLK(clk), .RST(rst), .Q(
        start_reg[113]) );
  DFF \start_reg_reg[114]  ( .D(start_in[113]), .CLK(clk), .RST(rst), .Q(
        start_reg[114]) );
  DFF \start_reg_reg[115]  ( .D(start_in[114]), .CLK(clk), .RST(rst), .Q(
        start_reg[115]) );
  DFF \start_reg_reg[116]  ( .D(start_in[115]), .CLK(clk), .RST(rst), .Q(
        start_reg[116]) );
  DFF \start_reg_reg[117]  ( .D(start_in[116]), .CLK(clk), .RST(rst), .Q(
        start_reg[117]) );
  DFF \start_reg_reg[118]  ( .D(start_in[117]), .CLK(clk), .RST(rst), .Q(
        start_reg[118]) );
  DFF \start_reg_reg[119]  ( .D(start_in[118]), .CLK(clk), .RST(rst), .Q(
        start_reg[119]) );
  DFF \start_reg_reg[120]  ( .D(start_in[119]), .CLK(clk), .RST(rst), .Q(
        start_reg[120]) );
  DFF \start_reg_reg[121]  ( .D(start_in[120]), .CLK(clk), .RST(rst), .Q(
        start_reg[121]) );
  DFF \start_reg_reg[122]  ( .D(start_in[121]), .CLK(clk), .RST(rst), .Q(
        start_reg[122]) );
  DFF \start_reg_reg[123]  ( .D(start_in[122]), .CLK(clk), .RST(rst), .Q(
        start_reg[123]) );
  DFF \start_reg_reg[124]  ( .D(start_in[123]), .CLK(clk), .RST(rst), .Q(
        start_reg[124]) );
  DFF \start_reg_reg[125]  ( .D(start_in[124]), .CLK(clk), .RST(rst), .Q(
        start_reg[125]) );
  DFF \start_reg_reg[126]  ( .D(start_in[125]), .CLK(clk), .RST(rst), .Q(
        start_reg[126]) );
  DFF \start_reg_reg[127]  ( .D(start_in[126]), .CLK(clk), .RST(rst), .Q(
        start_reg[127]) );
  DFF \start_reg_reg[128]  ( .D(start_in[127]), .CLK(clk), .RST(rst), .Q(
        start_reg[128]) );
  DFF \start_reg_reg[129]  ( .D(start_in[128]), .CLK(clk), .RST(rst), .Q(
        start_reg[129]) );
  DFF \start_reg_reg[130]  ( .D(start_in[129]), .CLK(clk), .RST(rst), .Q(
        start_reg[130]) );
  DFF \start_reg_reg[131]  ( .D(start_in[130]), .CLK(clk), .RST(rst), .Q(
        start_reg[131]) );
  DFF \start_reg_reg[132]  ( .D(start_in[131]), .CLK(clk), .RST(rst), .Q(
        start_reg[132]) );
  DFF \start_reg_reg[133]  ( .D(start_in[132]), .CLK(clk), .RST(rst), .Q(
        start_reg[133]) );
  DFF \start_reg_reg[134]  ( .D(start_in[133]), .CLK(clk), .RST(rst), .Q(
        start_reg[134]) );
  DFF \start_reg_reg[135]  ( .D(start_in[134]), .CLK(clk), .RST(rst), .Q(
        start_reg[135]) );
  DFF \start_reg_reg[136]  ( .D(start_in[135]), .CLK(clk), .RST(rst), .Q(
        start_reg[136]) );
  DFF \start_reg_reg[137]  ( .D(start_in[136]), .CLK(clk), .RST(rst), .Q(
        start_reg[137]) );
  DFF \start_reg_reg[138]  ( .D(start_in[137]), .CLK(clk), .RST(rst), .Q(
        start_reg[138]) );
  DFF \start_reg_reg[139]  ( .D(start_in[138]), .CLK(clk), .RST(rst), .Q(
        start_reg[139]) );
  DFF \start_reg_reg[140]  ( .D(start_in[139]), .CLK(clk), .RST(rst), .Q(
        start_reg[140]) );
  DFF \start_reg_reg[141]  ( .D(start_in[140]), .CLK(clk), .RST(rst), .Q(
        start_reg[141]) );
  DFF \start_reg_reg[142]  ( .D(start_in[141]), .CLK(clk), .RST(rst), .Q(
        start_reg[142]) );
  DFF \start_reg_reg[143]  ( .D(start_in[142]), .CLK(clk), .RST(rst), .Q(
        start_reg[143]) );
  DFF \start_reg_reg[144]  ( .D(start_in[143]), .CLK(clk), .RST(rst), .Q(
        start_reg[144]) );
  DFF \start_reg_reg[145]  ( .D(start_in[144]), .CLK(clk), .RST(rst), .Q(
        start_reg[145]) );
  DFF \start_reg_reg[146]  ( .D(start_in[145]), .CLK(clk), .RST(rst), .Q(
        start_reg[146]) );
  DFF \start_reg_reg[147]  ( .D(start_in[146]), .CLK(clk), .RST(rst), .Q(
        start_reg[147]) );
  DFF \start_reg_reg[148]  ( .D(start_in[147]), .CLK(clk), .RST(rst), .Q(
        start_reg[148]) );
  DFF \start_reg_reg[149]  ( .D(start_in[148]), .CLK(clk), .RST(rst), .Q(
        start_reg[149]) );
  DFF \start_reg_reg[150]  ( .D(start_in[149]), .CLK(clk), .RST(rst), .Q(
        start_reg[150]) );
  DFF \start_reg_reg[151]  ( .D(start_in[150]), .CLK(clk), .RST(rst), .Q(
        start_reg[151]) );
  DFF \start_reg_reg[152]  ( .D(start_in[151]), .CLK(clk), .RST(rst), .Q(
        start_reg[152]) );
  DFF \start_reg_reg[153]  ( .D(start_in[152]), .CLK(clk), .RST(rst), .Q(
        start_reg[153]) );
  DFF \start_reg_reg[154]  ( .D(start_in[153]), .CLK(clk), .RST(rst), .Q(
        start_reg[154]) );
  DFF \start_reg_reg[155]  ( .D(start_in[154]), .CLK(clk), .RST(rst), .Q(
        start_reg[155]) );
  DFF \start_reg_reg[156]  ( .D(start_in[155]), .CLK(clk), .RST(rst), .Q(
        start_reg[156]) );
  DFF \start_reg_reg[157]  ( .D(start_in[156]), .CLK(clk), .RST(rst), .Q(
        start_reg[157]) );
  DFF \start_reg_reg[158]  ( .D(start_in[157]), .CLK(clk), .RST(rst), .Q(
        start_reg[158]) );
  DFF \start_reg_reg[159]  ( .D(start_in[158]), .CLK(clk), .RST(rst), .Q(
        start_reg[159]) );
  DFF \start_reg_reg[160]  ( .D(start_in[159]), .CLK(clk), .RST(rst), .Q(
        start_reg[160]) );
  DFF \start_reg_reg[161]  ( .D(start_in[160]), .CLK(clk), .RST(rst), .Q(
        start_reg[161]) );
  DFF \start_reg_reg[162]  ( .D(start_in[161]), .CLK(clk), .RST(rst), .Q(
        start_reg[162]) );
  DFF \start_reg_reg[163]  ( .D(start_in[162]), .CLK(clk), .RST(rst), .Q(
        start_reg[163]) );
  DFF \start_reg_reg[164]  ( .D(start_in[163]), .CLK(clk), .RST(rst), .Q(
        start_reg[164]) );
  DFF \start_reg_reg[165]  ( .D(start_in[164]), .CLK(clk), .RST(rst), .Q(
        start_reg[165]) );
  DFF \start_reg_reg[166]  ( .D(start_in[165]), .CLK(clk), .RST(rst), .Q(
        start_reg[166]) );
  DFF \start_reg_reg[167]  ( .D(start_in[166]), .CLK(clk), .RST(rst), .Q(
        start_reg[167]) );
  DFF \start_reg_reg[168]  ( .D(start_in[167]), .CLK(clk), .RST(rst), .Q(
        start_reg[168]) );
  DFF \start_reg_reg[169]  ( .D(start_in[168]), .CLK(clk), .RST(rst), .Q(
        start_reg[169]) );
  DFF \start_reg_reg[170]  ( .D(start_in[169]), .CLK(clk), .RST(rst), .Q(
        start_reg[170]) );
  DFF \start_reg_reg[171]  ( .D(start_in[170]), .CLK(clk), .RST(rst), .Q(
        start_reg[171]) );
  DFF \start_reg_reg[172]  ( .D(start_in[171]), .CLK(clk), .RST(rst), .Q(
        start_reg[172]) );
  DFF \start_reg_reg[173]  ( .D(start_in[172]), .CLK(clk), .RST(rst), .Q(
        start_reg[173]) );
  DFF \start_reg_reg[174]  ( .D(start_in[173]), .CLK(clk), .RST(rst), .Q(
        start_reg[174]) );
  DFF \start_reg_reg[175]  ( .D(start_in[174]), .CLK(clk), .RST(rst), .Q(
        start_reg[175]) );
  DFF \start_reg_reg[176]  ( .D(start_in[175]), .CLK(clk), .RST(rst), .Q(
        start_reg[176]) );
  DFF \start_reg_reg[177]  ( .D(start_in[176]), .CLK(clk), .RST(rst), .Q(
        start_reg[177]) );
  DFF \start_reg_reg[178]  ( .D(start_in[177]), .CLK(clk), .RST(rst), .Q(
        start_reg[178]) );
  DFF \start_reg_reg[179]  ( .D(start_in[178]), .CLK(clk), .RST(rst), .Q(
        start_reg[179]) );
  DFF \start_reg_reg[180]  ( .D(start_in[179]), .CLK(clk), .RST(rst), .Q(
        start_reg[180]) );
  DFF \start_reg_reg[181]  ( .D(start_in[180]), .CLK(clk), .RST(rst), .Q(
        start_reg[181]) );
  DFF \start_reg_reg[182]  ( .D(start_in[181]), .CLK(clk), .RST(rst), .Q(
        start_reg[182]) );
  DFF \start_reg_reg[183]  ( .D(start_in[182]), .CLK(clk), .RST(rst), .Q(
        start_reg[183]) );
  DFF \start_reg_reg[184]  ( .D(start_in[183]), .CLK(clk), .RST(rst), .Q(
        start_reg[184]) );
  DFF \start_reg_reg[185]  ( .D(start_in[184]), .CLK(clk), .RST(rst), .Q(
        start_reg[185]) );
  DFF \start_reg_reg[186]  ( .D(start_in[185]), .CLK(clk), .RST(rst), .Q(
        start_reg[186]) );
  DFF \start_reg_reg[187]  ( .D(start_in[186]), .CLK(clk), .RST(rst), .Q(
        start_reg[187]) );
  DFF \start_reg_reg[188]  ( .D(start_in[187]), .CLK(clk), .RST(rst), .Q(
        start_reg[188]) );
  DFF \start_reg_reg[189]  ( .D(start_in[188]), .CLK(clk), .RST(rst), .Q(
        start_reg[189]) );
  DFF \start_reg_reg[190]  ( .D(start_in[189]), .CLK(clk), .RST(rst), .Q(
        start_reg[190]) );
  DFF \start_reg_reg[191]  ( .D(start_in[190]), .CLK(clk), .RST(rst), .Q(
        start_reg[191]) );
  DFF \start_reg_reg[192]  ( .D(start_in[191]), .CLK(clk), .RST(rst), .Q(
        start_reg[192]) );
  DFF \start_reg_reg[193]  ( .D(start_in[192]), .CLK(clk), .RST(rst), .Q(
        start_reg[193]) );
  DFF \start_reg_reg[194]  ( .D(start_in[193]), .CLK(clk), .RST(rst), .Q(
        start_reg[194]) );
  DFF \start_reg_reg[195]  ( .D(start_in[194]), .CLK(clk), .RST(rst), .Q(
        start_reg[195]) );
  DFF \start_reg_reg[196]  ( .D(start_in[195]), .CLK(clk), .RST(rst), .Q(
        start_reg[196]) );
  DFF \start_reg_reg[197]  ( .D(start_in[196]), .CLK(clk), .RST(rst), .Q(
        start_reg[197]) );
  DFF \start_reg_reg[198]  ( .D(start_in[197]), .CLK(clk), .RST(rst), .Q(
        start_reg[198]) );
  DFF \start_reg_reg[199]  ( .D(start_in[198]), .CLK(clk), .RST(rst), .Q(
        start_reg[199]) );
  DFF \start_reg_reg[200]  ( .D(start_in[199]), .CLK(clk), .RST(rst), .Q(
        start_reg[200]) );
  DFF \start_reg_reg[201]  ( .D(start_in[200]), .CLK(clk), .RST(rst), .Q(
        start_reg[201]) );
  DFF \start_reg_reg[202]  ( .D(start_in[201]), .CLK(clk), .RST(rst), .Q(
        start_reg[202]) );
  DFF \start_reg_reg[203]  ( .D(start_in[202]), .CLK(clk), .RST(rst), .Q(
        start_reg[203]) );
  DFF \start_reg_reg[204]  ( .D(start_in[203]), .CLK(clk), .RST(rst), .Q(
        start_reg[204]) );
  DFF \start_reg_reg[205]  ( .D(start_in[204]), .CLK(clk), .RST(rst), .Q(
        start_reg[205]) );
  DFF \start_reg_reg[206]  ( .D(start_in[205]), .CLK(clk), .RST(rst), .Q(
        start_reg[206]) );
  DFF \start_reg_reg[207]  ( .D(start_in[206]), .CLK(clk), .RST(rst), .Q(
        start_reg[207]) );
  DFF \start_reg_reg[208]  ( .D(start_in[207]), .CLK(clk), .RST(rst), .Q(
        start_reg[208]) );
  DFF \start_reg_reg[209]  ( .D(start_in[208]), .CLK(clk), .RST(rst), .Q(
        start_reg[209]) );
  DFF \start_reg_reg[210]  ( .D(start_in[209]), .CLK(clk), .RST(rst), .Q(
        start_reg[210]) );
  DFF \start_reg_reg[211]  ( .D(start_in[210]), .CLK(clk), .RST(rst), .Q(
        start_reg[211]) );
  DFF \start_reg_reg[212]  ( .D(start_in[211]), .CLK(clk), .RST(rst), .Q(
        start_reg[212]) );
  DFF \start_reg_reg[213]  ( .D(start_in[212]), .CLK(clk), .RST(rst), .Q(
        start_reg[213]) );
  DFF \start_reg_reg[214]  ( .D(start_in[213]), .CLK(clk), .RST(rst), .Q(
        start_reg[214]) );
  DFF \start_reg_reg[215]  ( .D(start_in[214]), .CLK(clk), .RST(rst), .Q(
        start_reg[215]) );
  DFF \start_reg_reg[216]  ( .D(start_in[215]), .CLK(clk), .RST(rst), .Q(
        start_reg[216]) );
  DFF \start_reg_reg[217]  ( .D(start_in[216]), .CLK(clk), .RST(rst), .Q(
        start_reg[217]) );
  DFF \start_reg_reg[218]  ( .D(start_in[217]), .CLK(clk), .RST(rst), .Q(
        start_reg[218]) );
  DFF \start_reg_reg[219]  ( .D(start_in[218]), .CLK(clk), .RST(rst), .Q(
        start_reg[219]) );
  DFF \start_reg_reg[220]  ( .D(start_in[219]), .CLK(clk), .RST(rst), .Q(
        start_reg[220]) );
  DFF \start_reg_reg[221]  ( .D(start_in[220]), .CLK(clk), .RST(rst), .Q(
        start_reg[221]) );
  DFF \start_reg_reg[222]  ( .D(start_in[221]), .CLK(clk), .RST(rst), .Q(
        start_reg[222]) );
  DFF \start_reg_reg[223]  ( .D(start_in[222]), .CLK(clk), .RST(rst), .Q(
        start_reg[223]) );
  DFF \start_reg_reg[224]  ( .D(start_in[223]), .CLK(clk), .RST(rst), .Q(
        start_reg[224]) );
  DFF \start_reg_reg[225]  ( .D(start_in[224]), .CLK(clk), .RST(rst), .Q(
        start_reg[225]) );
  DFF \start_reg_reg[226]  ( .D(start_in[225]), .CLK(clk), .RST(rst), .Q(
        start_reg[226]) );
  DFF \start_reg_reg[227]  ( .D(start_in[226]), .CLK(clk), .RST(rst), .Q(
        start_reg[227]) );
  DFF \start_reg_reg[228]  ( .D(start_in[227]), .CLK(clk), .RST(rst), .Q(
        start_reg[228]) );
  DFF \start_reg_reg[229]  ( .D(start_in[228]), .CLK(clk), .RST(rst), .Q(
        start_reg[229]) );
  DFF \start_reg_reg[230]  ( .D(start_in[229]), .CLK(clk), .RST(rst), .Q(
        start_reg[230]) );
  DFF \start_reg_reg[231]  ( .D(start_in[230]), .CLK(clk), .RST(rst), .Q(
        start_reg[231]) );
  DFF \start_reg_reg[232]  ( .D(start_in[231]), .CLK(clk), .RST(rst), .Q(
        start_reg[232]) );
  DFF \start_reg_reg[233]  ( .D(start_in[232]), .CLK(clk), .RST(rst), .Q(
        start_reg[233]) );
  DFF \start_reg_reg[234]  ( .D(start_in[233]), .CLK(clk), .RST(rst), .Q(
        start_reg[234]) );
  DFF \start_reg_reg[235]  ( .D(start_in[234]), .CLK(clk), .RST(rst), .Q(
        start_reg[235]) );
  DFF \start_reg_reg[236]  ( .D(start_in[235]), .CLK(clk), .RST(rst), .Q(
        start_reg[236]) );
  DFF \start_reg_reg[237]  ( .D(start_in[236]), .CLK(clk), .RST(rst), .Q(
        start_reg[237]) );
  DFF \start_reg_reg[238]  ( .D(start_in[237]), .CLK(clk), .RST(rst), .Q(
        start_reg[238]) );
  DFF \start_reg_reg[239]  ( .D(start_in[238]), .CLK(clk), .RST(rst), .Q(
        start_reg[239]) );
  DFF \start_reg_reg[240]  ( .D(start_in[239]), .CLK(clk), .RST(rst), .Q(
        start_reg[240]) );
  DFF \start_reg_reg[241]  ( .D(start_in[240]), .CLK(clk), .RST(rst), .Q(
        start_reg[241]) );
  DFF \start_reg_reg[242]  ( .D(start_in[241]), .CLK(clk), .RST(rst), .Q(
        start_reg[242]) );
  DFF \start_reg_reg[243]  ( .D(start_in[242]), .CLK(clk), .RST(rst), .Q(
        start_reg[243]) );
  DFF \start_reg_reg[244]  ( .D(start_in[243]), .CLK(clk), .RST(rst), .Q(
        start_reg[244]) );
  DFF \start_reg_reg[245]  ( .D(start_in[244]), .CLK(clk), .RST(rst), .Q(
        start_reg[245]) );
  DFF \start_reg_reg[246]  ( .D(start_in[245]), .CLK(clk), .RST(rst), .Q(
        start_reg[246]) );
  DFF \start_reg_reg[247]  ( .D(start_in[246]), .CLK(clk), .RST(rst), .Q(
        start_reg[247]) );
  DFF \start_reg_reg[248]  ( .D(start_in[247]), .CLK(clk), .RST(rst), .Q(
        start_reg[248]) );
  DFF \start_reg_reg[249]  ( .D(start_in[248]), .CLK(clk), .RST(rst), .Q(
        start_reg[249]) );
  DFF \start_reg_reg[250]  ( .D(start_in[249]), .CLK(clk), .RST(rst), .Q(
        start_reg[250]) );
  DFF \start_reg_reg[251]  ( .D(start_in[250]), .CLK(clk), .RST(rst), .Q(
        start_reg[251]) );
  DFF \start_reg_reg[252]  ( .D(start_in[251]), .CLK(clk), .RST(rst), .Q(
        start_reg[252]) );
  DFF \start_reg_reg[253]  ( .D(start_in[252]), .CLK(clk), .RST(rst), .Q(
        start_reg[253]) );
  DFF \start_reg_reg[254]  ( .D(start_in[253]), .CLK(clk), .RST(rst), .Q(
        start_reg[254]) );
  DFF \start_reg_reg[255]  ( .D(start_in[254]), .CLK(clk), .RST(rst), .Q(
        start_reg[255]) );
  DFF \start_reg_reg[256]  ( .D(start_in[255]), .CLK(clk), .RST(rst), .Q(
        start_reg[256]) );
  DFF \start_reg_reg[257]  ( .D(start_in[256]), .CLK(clk), .RST(rst), .Q(
        start_reg[257]) );
  DFF \start_reg_reg[258]  ( .D(start_in[257]), .CLK(clk), .RST(rst), .Q(
        start_reg[258]) );
  DFF \start_reg_reg[259]  ( .D(start_in[258]), .CLK(clk), .RST(rst), .Q(
        start_reg[259]) );
  DFF \start_reg_reg[260]  ( .D(start_in[259]), .CLK(clk), .RST(rst), .Q(
        start_reg[260]) );
  DFF \start_reg_reg[261]  ( .D(start_in[260]), .CLK(clk), .RST(rst), .Q(
        start_reg[261]) );
  DFF \start_reg_reg[262]  ( .D(start_in[261]), .CLK(clk), .RST(rst), .Q(
        start_reg[262]) );
  DFF \start_reg_reg[263]  ( .D(start_in[262]), .CLK(clk), .RST(rst), .Q(
        start_reg[263]) );
  DFF \start_reg_reg[264]  ( .D(start_in[263]), .CLK(clk), .RST(rst), .Q(
        start_reg[264]) );
  DFF \start_reg_reg[265]  ( .D(start_in[264]), .CLK(clk), .RST(rst), .Q(
        start_reg[265]) );
  DFF \start_reg_reg[266]  ( .D(start_in[265]), .CLK(clk), .RST(rst), .Q(
        start_reg[266]) );
  DFF \start_reg_reg[267]  ( .D(start_in[266]), .CLK(clk), .RST(rst), .Q(
        start_reg[267]) );
  DFF \start_reg_reg[268]  ( .D(start_in[267]), .CLK(clk), .RST(rst), .Q(
        start_reg[268]) );
  DFF \start_reg_reg[269]  ( .D(start_in[268]), .CLK(clk), .RST(rst), .Q(
        start_reg[269]) );
  DFF \start_reg_reg[270]  ( .D(start_in[269]), .CLK(clk), .RST(rst), .Q(
        start_reg[270]) );
  DFF \start_reg_reg[271]  ( .D(start_in[270]), .CLK(clk), .RST(rst), .Q(
        start_reg[271]) );
  DFF \start_reg_reg[272]  ( .D(start_in[271]), .CLK(clk), .RST(rst), .Q(
        start_reg[272]) );
  DFF \start_reg_reg[273]  ( .D(start_in[272]), .CLK(clk), .RST(rst), .Q(
        start_reg[273]) );
  DFF \start_reg_reg[274]  ( .D(start_in[273]), .CLK(clk), .RST(rst), .Q(
        start_reg[274]) );
  DFF \start_reg_reg[275]  ( .D(start_in[274]), .CLK(clk), .RST(rst), .Q(
        start_reg[275]) );
  DFF \start_reg_reg[276]  ( .D(start_in[275]), .CLK(clk), .RST(rst), .Q(
        start_reg[276]) );
  DFF \start_reg_reg[277]  ( .D(start_in[276]), .CLK(clk), .RST(rst), .Q(
        start_reg[277]) );
  DFF \start_reg_reg[278]  ( .D(start_in[277]), .CLK(clk), .RST(rst), .Q(
        start_reg[278]) );
  DFF \start_reg_reg[279]  ( .D(start_in[278]), .CLK(clk), .RST(rst), .Q(
        start_reg[279]) );
  DFF \start_reg_reg[280]  ( .D(start_in[279]), .CLK(clk), .RST(rst), .Q(
        start_reg[280]) );
  DFF \start_reg_reg[281]  ( .D(start_in[280]), .CLK(clk), .RST(rst), .Q(
        start_reg[281]) );
  DFF \start_reg_reg[282]  ( .D(start_in[281]), .CLK(clk), .RST(rst), .Q(
        start_reg[282]) );
  DFF \start_reg_reg[283]  ( .D(start_in[282]), .CLK(clk), .RST(rst), .Q(
        start_reg[283]) );
  DFF \start_reg_reg[284]  ( .D(start_in[283]), .CLK(clk), .RST(rst), .Q(
        start_reg[284]) );
  DFF \start_reg_reg[285]  ( .D(start_in[284]), .CLK(clk), .RST(rst), .Q(
        start_reg[285]) );
  DFF \start_reg_reg[286]  ( .D(start_in[285]), .CLK(clk), .RST(rst), .Q(
        start_reg[286]) );
  DFF \start_reg_reg[287]  ( .D(start_in[286]), .CLK(clk), .RST(rst), .Q(
        start_reg[287]) );
  DFF \start_reg_reg[288]  ( .D(start_in[287]), .CLK(clk), .RST(rst), .Q(
        start_reg[288]) );
  DFF \start_reg_reg[289]  ( .D(start_in[288]), .CLK(clk), .RST(rst), .Q(
        start_reg[289]) );
  DFF \start_reg_reg[290]  ( .D(start_in[289]), .CLK(clk), .RST(rst), .Q(
        start_reg[290]) );
  DFF \start_reg_reg[291]  ( .D(start_in[290]), .CLK(clk), .RST(rst), .Q(
        start_reg[291]) );
  DFF \start_reg_reg[292]  ( .D(start_in[291]), .CLK(clk), .RST(rst), .Q(
        start_reg[292]) );
  DFF \start_reg_reg[293]  ( .D(start_in[292]), .CLK(clk), .RST(rst), .Q(
        start_reg[293]) );
  DFF \start_reg_reg[294]  ( .D(start_in[293]), .CLK(clk), .RST(rst), .Q(
        start_reg[294]) );
  DFF \start_reg_reg[295]  ( .D(start_in[294]), .CLK(clk), .RST(rst), .Q(
        start_reg[295]) );
  DFF \start_reg_reg[296]  ( .D(start_in[295]), .CLK(clk), .RST(rst), .Q(
        start_reg[296]) );
  DFF \start_reg_reg[297]  ( .D(start_in[296]), .CLK(clk), .RST(rst), .Q(
        start_reg[297]) );
  DFF \start_reg_reg[298]  ( .D(start_in[297]), .CLK(clk), .RST(rst), .Q(
        start_reg[298]) );
  DFF \start_reg_reg[299]  ( .D(start_in[298]), .CLK(clk), .RST(rst), .Q(
        start_reg[299]) );
  DFF \start_reg_reg[300]  ( .D(start_in[299]), .CLK(clk), .RST(rst), .Q(
        start_reg[300]) );
  DFF \start_reg_reg[301]  ( .D(start_in[300]), .CLK(clk), .RST(rst), .Q(
        start_reg[301]) );
  DFF \start_reg_reg[302]  ( .D(start_in[301]), .CLK(clk), .RST(rst), .Q(
        start_reg[302]) );
  DFF \start_reg_reg[303]  ( .D(start_in[302]), .CLK(clk), .RST(rst), .Q(
        start_reg[303]) );
  DFF \start_reg_reg[304]  ( .D(start_in[303]), .CLK(clk), .RST(rst), .Q(
        start_reg[304]) );
  DFF \start_reg_reg[305]  ( .D(start_in[304]), .CLK(clk), .RST(rst), .Q(
        start_reg[305]) );
  DFF \start_reg_reg[306]  ( .D(start_in[305]), .CLK(clk), .RST(rst), .Q(
        start_reg[306]) );
  DFF \start_reg_reg[307]  ( .D(start_in[306]), .CLK(clk), .RST(rst), .Q(
        start_reg[307]) );
  DFF \start_reg_reg[308]  ( .D(start_in[307]), .CLK(clk), .RST(rst), .Q(
        start_reg[308]) );
  DFF \start_reg_reg[309]  ( .D(start_in[308]), .CLK(clk), .RST(rst), .Q(
        start_reg[309]) );
  DFF \start_reg_reg[310]  ( .D(start_in[309]), .CLK(clk), .RST(rst), .Q(
        start_reg[310]) );
  DFF \start_reg_reg[311]  ( .D(start_in[310]), .CLK(clk), .RST(rst), .Q(
        start_reg[311]) );
  DFF \start_reg_reg[312]  ( .D(start_in[311]), .CLK(clk), .RST(rst), .Q(
        start_reg[312]) );
  DFF \start_reg_reg[313]  ( .D(start_in[312]), .CLK(clk), .RST(rst), .Q(
        start_reg[313]) );
  DFF \start_reg_reg[314]  ( .D(start_in[313]), .CLK(clk), .RST(rst), .Q(
        start_reg[314]) );
  DFF \start_reg_reg[315]  ( .D(start_in[314]), .CLK(clk), .RST(rst), .Q(
        start_reg[315]) );
  DFF \start_reg_reg[316]  ( .D(start_in[315]), .CLK(clk), .RST(rst), .Q(
        start_reg[316]) );
  DFF \start_reg_reg[317]  ( .D(start_in[316]), .CLK(clk), .RST(rst), .Q(
        start_reg[317]) );
  DFF \start_reg_reg[318]  ( .D(start_in[317]), .CLK(clk), .RST(rst), .Q(
        start_reg[318]) );
  DFF \start_reg_reg[319]  ( .D(start_in[318]), .CLK(clk), .RST(rst), .Q(
        start_reg[319]) );
  DFF \start_reg_reg[320]  ( .D(start_in[319]), .CLK(clk), .RST(rst), .Q(
        start_reg[320]) );
  DFF \start_reg_reg[321]  ( .D(start_in[320]), .CLK(clk), .RST(rst), .Q(
        start_reg[321]) );
  DFF \start_reg_reg[322]  ( .D(start_in[321]), .CLK(clk), .RST(rst), .Q(
        start_reg[322]) );
  DFF \start_reg_reg[323]  ( .D(start_in[322]), .CLK(clk), .RST(rst), .Q(
        start_reg[323]) );
  DFF \start_reg_reg[324]  ( .D(start_in[323]), .CLK(clk), .RST(rst), .Q(
        start_reg[324]) );
  DFF \start_reg_reg[325]  ( .D(start_in[324]), .CLK(clk), .RST(rst), .Q(
        start_reg[325]) );
  DFF \start_reg_reg[326]  ( .D(start_in[325]), .CLK(clk), .RST(rst), .Q(
        start_reg[326]) );
  DFF \start_reg_reg[327]  ( .D(start_in[326]), .CLK(clk), .RST(rst), .Q(
        start_reg[327]) );
  DFF \start_reg_reg[328]  ( .D(start_in[327]), .CLK(clk), .RST(rst), .Q(
        start_reg[328]) );
  DFF \start_reg_reg[329]  ( .D(start_in[328]), .CLK(clk), .RST(rst), .Q(
        start_reg[329]) );
  DFF \start_reg_reg[330]  ( .D(start_in[329]), .CLK(clk), .RST(rst), .Q(
        start_reg[330]) );
  DFF \start_reg_reg[331]  ( .D(start_in[330]), .CLK(clk), .RST(rst), .Q(
        start_reg[331]) );
  DFF \start_reg_reg[332]  ( .D(start_in[331]), .CLK(clk), .RST(rst), .Q(
        start_reg[332]) );
  DFF \start_reg_reg[333]  ( .D(start_in[332]), .CLK(clk), .RST(rst), .Q(
        start_reg[333]) );
  DFF \start_reg_reg[334]  ( .D(start_in[333]), .CLK(clk), .RST(rst), .Q(
        start_reg[334]) );
  DFF \start_reg_reg[335]  ( .D(start_in[334]), .CLK(clk), .RST(rst), .Q(
        start_reg[335]) );
  DFF \start_reg_reg[336]  ( .D(start_in[335]), .CLK(clk), .RST(rst), .Q(
        start_reg[336]) );
  DFF \start_reg_reg[337]  ( .D(start_in[336]), .CLK(clk), .RST(rst), .Q(
        start_reg[337]) );
  DFF \start_reg_reg[338]  ( .D(start_in[337]), .CLK(clk), .RST(rst), .Q(
        start_reg[338]) );
  DFF \start_reg_reg[339]  ( .D(start_in[338]), .CLK(clk), .RST(rst), .Q(
        start_reg[339]) );
  DFF \start_reg_reg[340]  ( .D(start_in[339]), .CLK(clk), .RST(rst), .Q(
        start_reg[340]) );
  DFF \start_reg_reg[341]  ( .D(start_in[340]), .CLK(clk), .RST(rst), .Q(
        start_reg[341]) );
  DFF \start_reg_reg[342]  ( .D(start_in[341]), .CLK(clk), .RST(rst), .Q(
        start_reg[342]) );
  DFF \start_reg_reg[343]  ( .D(start_in[342]), .CLK(clk), .RST(rst), .Q(
        start_reg[343]) );
  DFF \start_reg_reg[344]  ( .D(start_in[343]), .CLK(clk), .RST(rst), .Q(
        start_reg[344]) );
  DFF \start_reg_reg[345]  ( .D(start_in[344]), .CLK(clk), .RST(rst), .Q(
        start_reg[345]) );
  DFF \start_reg_reg[346]  ( .D(start_in[345]), .CLK(clk), .RST(rst), .Q(
        start_reg[346]) );
  DFF \start_reg_reg[347]  ( .D(start_in[346]), .CLK(clk), .RST(rst), .Q(
        start_reg[347]) );
  DFF \start_reg_reg[348]  ( .D(start_in[347]), .CLK(clk), .RST(rst), .Q(
        start_reg[348]) );
  DFF \start_reg_reg[349]  ( .D(start_in[348]), .CLK(clk), .RST(rst), .Q(
        start_reg[349]) );
  DFF \start_reg_reg[350]  ( .D(start_in[349]), .CLK(clk), .RST(rst), .Q(
        start_reg[350]) );
  DFF \start_reg_reg[351]  ( .D(start_in[350]), .CLK(clk), .RST(rst), .Q(
        start_reg[351]) );
  DFF \start_reg_reg[352]  ( .D(start_in[351]), .CLK(clk), .RST(rst), .Q(
        start_reg[352]) );
  DFF \start_reg_reg[353]  ( .D(start_in[352]), .CLK(clk), .RST(rst), .Q(
        start_reg[353]) );
  DFF \start_reg_reg[354]  ( .D(start_in[353]), .CLK(clk), .RST(rst), .Q(
        start_reg[354]) );
  DFF \start_reg_reg[355]  ( .D(start_in[354]), .CLK(clk), .RST(rst), .Q(
        start_reg[355]) );
  DFF \start_reg_reg[356]  ( .D(start_in[355]), .CLK(clk), .RST(rst), .Q(
        start_reg[356]) );
  DFF \start_reg_reg[357]  ( .D(start_in[356]), .CLK(clk), .RST(rst), .Q(
        start_reg[357]) );
  DFF \start_reg_reg[358]  ( .D(start_in[357]), .CLK(clk), .RST(rst), .Q(
        start_reg[358]) );
  DFF \start_reg_reg[359]  ( .D(start_in[358]), .CLK(clk), .RST(rst), .Q(
        start_reg[359]) );
  DFF \start_reg_reg[360]  ( .D(start_in[359]), .CLK(clk), .RST(rst), .Q(
        start_reg[360]) );
  DFF \start_reg_reg[361]  ( .D(start_in[360]), .CLK(clk), .RST(rst), .Q(
        start_reg[361]) );
  DFF \start_reg_reg[362]  ( .D(start_in[361]), .CLK(clk), .RST(rst), .Q(
        start_reg[362]) );
  DFF \start_reg_reg[363]  ( .D(start_in[362]), .CLK(clk), .RST(rst), .Q(
        start_reg[363]) );
  DFF \start_reg_reg[364]  ( .D(start_in[363]), .CLK(clk), .RST(rst), .Q(
        start_reg[364]) );
  DFF \start_reg_reg[365]  ( .D(start_in[364]), .CLK(clk), .RST(rst), .Q(
        start_reg[365]) );
  DFF \start_reg_reg[366]  ( .D(start_in[365]), .CLK(clk), .RST(rst), .Q(
        start_reg[366]) );
  DFF \start_reg_reg[367]  ( .D(start_in[366]), .CLK(clk), .RST(rst), .Q(
        start_reg[367]) );
  DFF \start_reg_reg[368]  ( .D(start_in[367]), .CLK(clk), .RST(rst), .Q(
        start_reg[368]) );
  DFF \start_reg_reg[369]  ( .D(start_in[368]), .CLK(clk), .RST(rst), .Q(
        start_reg[369]) );
  DFF \start_reg_reg[370]  ( .D(start_in[369]), .CLK(clk), .RST(rst), .Q(
        start_reg[370]) );
  DFF \start_reg_reg[371]  ( .D(start_in[370]), .CLK(clk), .RST(rst), .Q(
        start_reg[371]) );
  DFF \start_reg_reg[372]  ( .D(start_in[371]), .CLK(clk), .RST(rst), .Q(
        start_reg[372]) );
  DFF \start_reg_reg[373]  ( .D(start_in[372]), .CLK(clk), .RST(rst), .Q(
        start_reg[373]) );
  DFF \start_reg_reg[374]  ( .D(start_in[373]), .CLK(clk), .RST(rst), .Q(
        start_reg[374]) );
  DFF \start_reg_reg[375]  ( .D(start_in[374]), .CLK(clk), .RST(rst), .Q(
        start_reg[375]) );
  DFF \start_reg_reg[376]  ( .D(start_in[375]), .CLK(clk), .RST(rst), .Q(
        start_reg[376]) );
  DFF \start_reg_reg[377]  ( .D(start_in[376]), .CLK(clk), .RST(rst), .Q(
        start_reg[377]) );
  DFF \start_reg_reg[378]  ( .D(start_in[377]), .CLK(clk), .RST(rst), .Q(
        start_reg[378]) );
  DFF \start_reg_reg[379]  ( .D(start_in[378]), .CLK(clk), .RST(rst), .Q(
        start_reg[379]) );
  DFF \start_reg_reg[380]  ( .D(start_in[379]), .CLK(clk), .RST(rst), .Q(
        start_reg[380]) );
  DFF \start_reg_reg[381]  ( .D(start_in[380]), .CLK(clk), .RST(rst), .Q(
        start_reg[381]) );
  DFF \start_reg_reg[382]  ( .D(start_in[381]), .CLK(clk), .RST(rst), .Q(
        start_reg[382]) );
  DFF \start_reg_reg[383]  ( .D(start_in[382]), .CLK(clk), .RST(rst), .Q(
        start_reg[383]) );
  DFF \start_reg_reg[384]  ( .D(start_in[383]), .CLK(clk), .RST(rst), .Q(
        start_reg[384]) );
  DFF \start_reg_reg[385]  ( .D(start_in[384]), .CLK(clk), .RST(rst), .Q(
        start_reg[385]) );
  DFF \start_reg_reg[386]  ( .D(start_in[385]), .CLK(clk), .RST(rst), .Q(
        start_reg[386]) );
  DFF \start_reg_reg[387]  ( .D(start_in[386]), .CLK(clk), .RST(rst), .Q(
        start_reg[387]) );
  DFF \start_reg_reg[388]  ( .D(start_in[387]), .CLK(clk), .RST(rst), .Q(
        start_reg[388]) );
  DFF \start_reg_reg[389]  ( .D(start_in[388]), .CLK(clk), .RST(rst), .Q(
        start_reg[389]) );
  DFF \start_reg_reg[390]  ( .D(start_in[389]), .CLK(clk), .RST(rst), .Q(
        start_reg[390]) );
  DFF \start_reg_reg[391]  ( .D(start_in[390]), .CLK(clk), .RST(rst), .Q(
        start_reg[391]) );
  DFF \start_reg_reg[392]  ( .D(start_in[391]), .CLK(clk), .RST(rst), .Q(
        start_reg[392]) );
  DFF \start_reg_reg[393]  ( .D(start_in[392]), .CLK(clk), .RST(rst), .Q(
        start_reg[393]) );
  DFF \start_reg_reg[394]  ( .D(start_in[393]), .CLK(clk), .RST(rst), .Q(
        start_reg[394]) );
  DFF \start_reg_reg[395]  ( .D(start_in[394]), .CLK(clk), .RST(rst), .Q(
        start_reg[395]) );
  DFF \start_reg_reg[396]  ( .D(start_in[395]), .CLK(clk), .RST(rst), .Q(
        start_reg[396]) );
  DFF \start_reg_reg[397]  ( .D(start_in[396]), .CLK(clk), .RST(rst), .Q(
        start_reg[397]) );
  DFF \start_reg_reg[398]  ( .D(start_in[397]), .CLK(clk), .RST(rst), .Q(
        start_reg[398]) );
  DFF \start_reg_reg[399]  ( .D(start_in[398]), .CLK(clk), .RST(rst), .Q(
        start_reg[399]) );
  DFF \start_reg_reg[400]  ( .D(start_in[399]), .CLK(clk), .RST(rst), .Q(
        start_reg[400]) );
  DFF \start_reg_reg[401]  ( .D(start_in[400]), .CLK(clk), .RST(rst), .Q(
        start_reg[401]) );
  DFF \start_reg_reg[402]  ( .D(start_in[401]), .CLK(clk), .RST(rst), .Q(
        start_reg[402]) );
  DFF \start_reg_reg[403]  ( .D(start_in[402]), .CLK(clk), .RST(rst), .Q(
        start_reg[403]) );
  DFF \start_reg_reg[404]  ( .D(start_in[403]), .CLK(clk), .RST(rst), .Q(
        start_reg[404]) );
  DFF \start_reg_reg[405]  ( .D(start_in[404]), .CLK(clk), .RST(rst), .Q(
        start_reg[405]) );
  DFF \start_reg_reg[406]  ( .D(start_in[405]), .CLK(clk), .RST(rst), .Q(
        start_reg[406]) );
  DFF \start_reg_reg[407]  ( .D(start_in[406]), .CLK(clk), .RST(rst), .Q(
        start_reg[407]) );
  DFF \start_reg_reg[408]  ( .D(start_in[407]), .CLK(clk), .RST(rst), .Q(
        start_reg[408]) );
  DFF \start_reg_reg[409]  ( .D(start_in[408]), .CLK(clk), .RST(rst), .Q(
        start_reg[409]) );
  DFF \start_reg_reg[410]  ( .D(start_in[409]), .CLK(clk), .RST(rst), .Q(
        start_reg[410]) );
  DFF \start_reg_reg[411]  ( .D(start_in[410]), .CLK(clk), .RST(rst), .Q(
        start_reg[411]) );
  DFF \start_reg_reg[412]  ( .D(start_in[411]), .CLK(clk), .RST(rst), .Q(
        start_reg[412]) );
  DFF \start_reg_reg[413]  ( .D(start_in[412]), .CLK(clk), .RST(rst), .Q(
        start_reg[413]) );
  DFF \start_reg_reg[414]  ( .D(start_in[413]), .CLK(clk), .RST(rst), .Q(
        start_reg[414]) );
  DFF \start_reg_reg[415]  ( .D(start_in[414]), .CLK(clk), .RST(rst), .Q(
        start_reg[415]) );
  DFF \start_reg_reg[416]  ( .D(start_in[415]), .CLK(clk), .RST(rst), .Q(
        start_reg[416]) );
  DFF \start_reg_reg[417]  ( .D(start_in[416]), .CLK(clk), .RST(rst), .Q(
        start_reg[417]) );
  DFF \start_reg_reg[418]  ( .D(start_in[417]), .CLK(clk), .RST(rst), .Q(
        start_reg[418]) );
  DFF \start_reg_reg[419]  ( .D(start_in[418]), .CLK(clk), .RST(rst), .Q(
        start_reg[419]) );
  DFF \start_reg_reg[420]  ( .D(start_in[419]), .CLK(clk), .RST(rst), .Q(
        start_reg[420]) );
  DFF \start_reg_reg[421]  ( .D(start_in[420]), .CLK(clk), .RST(rst), .Q(
        start_reg[421]) );
  DFF \start_reg_reg[422]  ( .D(start_in[421]), .CLK(clk), .RST(rst), .Q(
        start_reg[422]) );
  DFF \start_reg_reg[423]  ( .D(start_in[422]), .CLK(clk), .RST(rst), .Q(
        start_reg[423]) );
  DFF \start_reg_reg[424]  ( .D(start_in[423]), .CLK(clk), .RST(rst), .Q(
        start_reg[424]) );
  DFF \start_reg_reg[425]  ( .D(start_in[424]), .CLK(clk), .RST(rst), .Q(
        start_reg[425]) );
  DFF \start_reg_reg[426]  ( .D(start_in[425]), .CLK(clk), .RST(rst), .Q(
        start_reg[426]) );
  DFF \start_reg_reg[427]  ( .D(start_in[426]), .CLK(clk), .RST(rst), .Q(
        start_reg[427]) );
  DFF \start_reg_reg[428]  ( .D(start_in[427]), .CLK(clk), .RST(rst), .Q(
        start_reg[428]) );
  DFF \start_reg_reg[429]  ( .D(start_in[428]), .CLK(clk), .RST(rst), .Q(
        start_reg[429]) );
  DFF \start_reg_reg[430]  ( .D(start_in[429]), .CLK(clk), .RST(rst), .Q(
        start_reg[430]) );
  DFF \start_reg_reg[431]  ( .D(start_in[430]), .CLK(clk), .RST(rst), .Q(
        start_reg[431]) );
  DFF \start_reg_reg[432]  ( .D(start_in[431]), .CLK(clk), .RST(rst), .Q(
        start_reg[432]) );
  DFF \start_reg_reg[433]  ( .D(start_in[432]), .CLK(clk), .RST(rst), .Q(
        start_reg[433]) );
  DFF \start_reg_reg[434]  ( .D(start_in[433]), .CLK(clk), .RST(rst), .Q(
        start_reg[434]) );
  DFF \start_reg_reg[435]  ( .D(start_in[434]), .CLK(clk), .RST(rst), .Q(
        start_reg[435]) );
  DFF \start_reg_reg[436]  ( .D(start_in[435]), .CLK(clk), .RST(rst), .Q(
        start_reg[436]) );
  DFF \start_reg_reg[437]  ( .D(start_in[436]), .CLK(clk), .RST(rst), .Q(
        start_reg[437]) );
  DFF \start_reg_reg[438]  ( .D(start_in[437]), .CLK(clk), .RST(rst), .Q(
        start_reg[438]) );
  DFF \start_reg_reg[439]  ( .D(start_in[438]), .CLK(clk), .RST(rst), .Q(
        start_reg[439]) );
  DFF \start_reg_reg[440]  ( .D(start_in[439]), .CLK(clk), .RST(rst), .Q(
        start_reg[440]) );
  DFF \start_reg_reg[441]  ( .D(start_in[440]), .CLK(clk), .RST(rst), .Q(
        start_reg[441]) );
  DFF \start_reg_reg[442]  ( .D(start_in[441]), .CLK(clk), .RST(rst), .Q(
        start_reg[442]) );
  DFF \start_reg_reg[443]  ( .D(start_in[442]), .CLK(clk), .RST(rst), .Q(
        start_reg[443]) );
  DFF \start_reg_reg[444]  ( .D(start_in[443]), .CLK(clk), .RST(rst), .Q(
        start_reg[444]) );
  DFF \start_reg_reg[445]  ( .D(start_in[444]), .CLK(clk), .RST(rst), .Q(
        start_reg[445]) );
  DFF \start_reg_reg[446]  ( .D(start_in[445]), .CLK(clk), .RST(rst), .Q(
        start_reg[446]) );
  DFF \start_reg_reg[447]  ( .D(start_in[446]), .CLK(clk), .RST(rst), .Q(
        start_reg[447]) );
  DFF \start_reg_reg[448]  ( .D(start_in[447]), .CLK(clk), .RST(rst), .Q(
        start_reg[448]) );
  DFF \start_reg_reg[449]  ( .D(start_in[448]), .CLK(clk), .RST(rst), .Q(
        start_reg[449]) );
  DFF \start_reg_reg[450]  ( .D(start_in[449]), .CLK(clk), .RST(rst), .Q(
        start_reg[450]) );
  DFF \start_reg_reg[451]  ( .D(start_in[450]), .CLK(clk), .RST(rst), .Q(
        start_reg[451]) );
  DFF \start_reg_reg[452]  ( .D(start_in[451]), .CLK(clk), .RST(rst), .Q(
        start_reg[452]) );
  DFF \start_reg_reg[453]  ( .D(start_in[452]), .CLK(clk), .RST(rst), .Q(
        start_reg[453]) );
  DFF \start_reg_reg[454]  ( .D(start_in[453]), .CLK(clk), .RST(rst), .Q(
        start_reg[454]) );
  DFF \start_reg_reg[455]  ( .D(start_in[454]), .CLK(clk), .RST(rst), .Q(
        start_reg[455]) );
  DFF \start_reg_reg[456]  ( .D(start_in[455]), .CLK(clk), .RST(rst), .Q(
        start_reg[456]) );
  DFF \start_reg_reg[457]  ( .D(start_in[456]), .CLK(clk), .RST(rst), .Q(
        start_reg[457]) );
  DFF \start_reg_reg[458]  ( .D(start_in[457]), .CLK(clk), .RST(rst), .Q(
        start_reg[458]) );
  DFF \start_reg_reg[459]  ( .D(start_in[458]), .CLK(clk), .RST(rst), .Q(
        start_reg[459]) );
  DFF \start_reg_reg[460]  ( .D(start_in[459]), .CLK(clk), .RST(rst), .Q(
        start_reg[460]) );
  DFF \start_reg_reg[461]  ( .D(start_in[460]), .CLK(clk), .RST(rst), .Q(
        start_reg[461]) );
  DFF \start_reg_reg[462]  ( .D(start_in[461]), .CLK(clk), .RST(rst), .Q(
        start_reg[462]) );
  DFF \start_reg_reg[463]  ( .D(start_in[462]), .CLK(clk), .RST(rst), .Q(
        start_reg[463]) );
  DFF \start_reg_reg[464]  ( .D(start_in[463]), .CLK(clk), .RST(rst), .Q(
        start_reg[464]) );
  DFF \start_reg_reg[465]  ( .D(start_in[464]), .CLK(clk), .RST(rst), .Q(
        start_reg[465]) );
  DFF \start_reg_reg[466]  ( .D(start_in[465]), .CLK(clk), .RST(rst), .Q(
        start_reg[466]) );
  DFF \start_reg_reg[467]  ( .D(start_in[466]), .CLK(clk), .RST(rst), .Q(
        start_reg[467]) );
  DFF \start_reg_reg[468]  ( .D(start_in[467]), .CLK(clk), .RST(rst), .Q(
        start_reg[468]) );
  DFF \start_reg_reg[469]  ( .D(start_in[468]), .CLK(clk), .RST(rst), .Q(
        start_reg[469]) );
  DFF \start_reg_reg[470]  ( .D(start_in[469]), .CLK(clk), .RST(rst), .Q(
        start_reg[470]) );
  DFF \start_reg_reg[471]  ( .D(start_in[470]), .CLK(clk), .RST(rst), .Q(
        start_reg[471]) );
  DFF \start_reg_reg[472]  ( .D(start_in[471]), .CLK(clk), .RST(rst), .Q(
        start_reg[472]) );
  DFF \start_reg_reg[473]  ( .D(start_in[472]), .CLK(clk), .RST(rst), .Q(
        start_reg[473]) );
  DFF \start_reg_reg[474]  ( .D(start_in[473]), .CLK(clk), .RST(rst), .Q(
        start_reg[474]) );
  DFF \start_reg_reg[475]  ( .D(start_in[474]), .CLK(clk), .RST(rst), .Q(
        start_reg[475]) );
  DFF \start_reg_reg[476]  ( .D(start_in[475]), .CLK(clk), .RST(rst), .Q(
        start_reg[476]) );
  DFF \start_reg_reg[477]  ( .D(start_in[476]), .CLK(clk), .RST(rst), .Q(
        start_reg[477]) );
  DFF \start_reg_reg[478]  ( .D(start_in[477]), .CLK(clk), .RST(rst), .Q(
        start_reg[478]) );
  DFF \start_reg_reg[479]  ( .D(start_in[478]), .CLK(clk), .RST(rst), .Q(
        start_reg[479]) );
  DFF \start_reg_reg[480]  ( .D(start_in[479]), .CLK(clk), .RST(rst), .Q(
        start_reg[480]) );
  DFF \start_reg_reg[481]  ( .D(start_in[480]), .CLK(clk), .RST(rst), .Q(
        start_reg[481]) );
  DFF \start_reg_reg[482]  ( .D(start_in[481]), .CLK(clk), .RST(rst), .Q(
        start_reg[482]) );
  DFF \start_reg_reg[483]  ( .D(start_in[482]), .CLK(clk), .RST(rst), .Q(
        start_reg[483]) );
  DFF \start_reg_reg[484]  ( .D(start_in[483]), .CLK(clk), .RST(rst), .Q(
        start_reg[484]) );
  DFF \start_reg_reg[485]  ( .D(start_in[484]), .CLK(clk), .RST(rst), .Q(
        start_reg[485]) );
  DFF \start_reg_reg[486]  ( .D(start_in[485]), .CLK(clk), .RST(rst), .Q(
        start_reg[486]) );
  DFF \start_reg_reg[487]  ( .D(start_in[486]), .CLK(clk), .RST(rst), .Q(
        start_reg[487]) );
  DFF \start_reg_reg[488]  ( .D(start_in[487]), .CLK(clk), .RST(rst), .Q(
        start_reg[488]) );
  DFF \start_reg_reg[489]  ( .D(start_in[488]), .CLK(clk), .RST(rst), .Q(
        start_reg[489]) );
  DFF \start_reg_reg[490]  ( .D(start_in[489]), .CLK(clk), .RST(rst), .Q(
        start_reg[490]) );
  DFF \start_reg_reg[491]  ( .D(start_in[490]), .CLK(clk), .RST(rst), .Q(
        start_reg[491]) );
  DFF \start_reg_reg[492]  ( .D(start_in[491]), .CLK(clk), .RST(rst), .Q(
        start_reg[492]) );
  DFF \start_reg_reg[493]  ( .D(start_in[492]), .CLK(clk), .RST(rst), .Q(
        start_reg[493]) );
  DFF \start_reg_reg[494]  ( .D(start_in[493]), .CLK(clk), .RST(rst), .Q(
        start_reg[494]) );
  DFF \start_reg_reg[495]  ( .D(start_in[494]), .CLK(clk), .RST(rst), .Q(
        start_reg[495]) );
  DFF \start_reg_reg[496]  ( .D(start_in[495]), .CLK(clk), .RST(rst), .Q(
        start_reg[496]) );
  DFF \start_reg_reg[497]  ( .D(start_in[496]), .CLK(clk), .RST(rst), .Q(
        start_reg[497]) );
  DFF \start_reg_reg[498]  ( .D(start_in[497]), .CLK(clk), .RST(rst), .Q(
        start_reg[498]) );
  DFF \start_reg_reg[499]  ( .D(start_in[498]), .CLK(clk), .RST(rst), .Q(
        start_reg[499]) );
  DFF \start_reg_reg[500]  ( .D(start_in[499]), .CLK(clk), .RST(rst), .Q(
        start_reg[500]) );
  DFF \start_reg_reg[501]  ( .D(start_in[500]), .CLK(clk), .RST(rst), .Q(
        start_reg[501]) );
  DFF \start_reg_reg[502]  ( .D(start_in[501]), .CLK(clk), .RST(rst), .Q(
        start_reg[502]) );
  DFF \start_reg_reg[503]  ( .D(start_in[502]), .CLK(clk), .RST(rst), .Q(
        start_reg[503]) );
  DFF \start_reg_reg[504]  ( .D(start_in[503]), .CLK(clk), .RST(rst), .Q(
        start_reg[504]) );
  DFF \start_reg_reg[505]  ( .D(start_in[504]), .CLK(clk), .RST(rst), .Q(
        start_reg[505]) );
  DFF \start_reg_reg[506]  ( .D(start_in[505]), .CLK(clk), .RST(rst), .Q(
        start_reg[506]) );
  DFF \start_reg_reg[507]  ( .D(start_in[506]), .CLK(clk), .RST(rst), .Q(
        start_reg[507]) );
  DFF \start_reg_reg[508]  ( .D(start_in[507]), .CLK(clk), .RST(rst), .Q(
        start_reg[508]) );
  DFF \start_reg_reg[509]  ( .D(start_in[508]), .CLK(clk), .RST(rst), .Q(
        start_reg[509]) );
  DFF \start_reg_reg[510]  ( .D(start_in[509]), .CLK(clk), .RST(rst), .Q(
        start_reg[510]) );
  DFF \start_reg_reg[511]  ( .D(start_in[510]), .CLK(clk), .RST(rst), .Q(
        start_reg[511]) );
  DFF \start_reg_reg[512]  ( .D(start_in[511]), .CLK(clk), .RST(rst), .Q(
        start_reg[512]) );
  DFF \start_reg_reg[513]  ( .D(start_in[512]), .CLK(clk), .RST(rst), .Q(
        start_reg[513]) );
  DFF \start_reg_reg[514]  ( .D(start_in[513]), .CLK(clk), .RST(rst), .Q(
        start_reg[514]) );
  DFF \start_reg_reg[515]  ( .D(start_in[514]), .CLK(clk), .RST(rst), .Q(
        start_reg[515]) );
  DFF \start_reg_reg[516]  ( .D(start_in[515]), .CLK(clk), .RST(rst), .Q(
        start_reg[516]) );
  DFF \start_reg_reg[517]  ( .D(start_in[516]), .CLK(clk), .RST(rst), .Q(
        start_reg[517]) );
  DFF \start_reg_reg[518]  ( .D(start_in[517]), .CLK(clk), .RST(rst), .Q(
        start_reg[518]) );
  DFF \start_reg_reg[519]  ( .D(start_in[518]), .CLK(clk), .RST(rst), .Q(
        start_reg[519]) );
  DFF \start_reg_reg[520]  ( .D(start_in[519]), .CLK(clk), .RST(rst), .Q(
        start_reg[520]) );
  DFF \start_reg_reg[521]  ( .D(start_in[520]), .CLK(clk), .RST(rst), .Q(
        start_reg[521]) );
  DFF \start_reg_reg[522]  ( .D(start_in[521]), .CLK(clk), .RST(rst), .Q(
        start_reg[522]) );
  DFF \start_reg_reg[523]  ( .D(start_in[522]), .CLK(clk), .RST(rst), .Q(
        start_reg[523]) );
  DFF \start_reg_reg[524]  ( .D(start_in[523]), .CLK(clk), .RST(rst), .Q(
        start_reg[524]) );
  DFF \start_reg_reg[525]  ( .D(start_in[524]), .CLK(clk), .RST(rst), .Q(
        start_reg[525]) );
  DFF \start_reg_reg[526]  ( .D(start_in[525]), .CLK(clk), .RST(rst), .Q(
        start_reg[526]) );
  DFF \start_reg_reg[527]  ( .D(start_in[526]), .CLK(clk), .RST(rst), .Q(
        start_reg[527]) );
  DFF \start_reg_reg[528]  ( .D(start_in[527]), .CLK(clk), .RST(rst), .Q(
        start_reg[528]) );
  DFF \start_reg_reg[529]  ( .D(start_in[528]), .CLK(clk), .RST(rst), .Q(
        start_reg[529]) );
  DFF \start_reg_reg[530]  ( .D(start_in[529]), .CLK(clk), .RST(rst), .Q(
        start_reg[530]) );
  DFF \start_reg_reg[531]  ( .D(start_in[530]), .CLK(clk), .RST(rst), .Q(
        start_reg[531]) );
  DFF \start_reg_reg[532]  ( .D(start_in[531]), .CLK(clk), .RST(rst), .Q(
        start_reg[532]) );
  DFF \start_reg_reg[533]  ( .D(start_in[532]), .CLK(clk), .RST(rst), .Q(
        start_reg[533]) );
  DFF \start_reg_reg[534]  ( .D(start_in[533]), .CLK(clk), .RST(rst), .Q(
        start_reg[534]) );
  DFF \start_reg_reg[535]  ( .D(start_in[534]), .CLK(clk), .RST(rst), .Q(
        start_reg[535]) );
  DFF \start_reg_reg[536]  ( .D(start_in[535]), .CLK(clk), .RST(rst), .Q(
        start_reg[536]) );
  DFF \start_reg_reg[537]  ( .D(start_in[536]), .CLK(clk), .RST(rst), .Q(
        start_reg[537]) );
  DFF \start_reg_reg[538]  ( .D(start_in[537]), .CLK(clk), .RST(rst), .Q(
        start_reg[538]) );
  DFF \start_reg_reg[539]  ( .D(start_in[538]), .CLK(clk), .RST(rst), .Q(
        start_reg[539]) );
  DFF \start_reg_reg[540]  ( .D(start_in[539]), .CLK(clk), .RST(rst), .Q(
        start_reg[540]) );
  DFF \start_reg_reg[541]  ( .D(start_in[540]), .CLK(clk), .RST(rst), .Q(
        start_reg[541]) );
  DFF \start_reg_reg[542]  ( .D(start_in[541]), .CLK(clk), .RST(rst), .Q(
        start_reg[542]) );
  DFF \start_reg_reg[543]  ( .D(start_in[542]), .CLK(clk), .RST(rst), .Q(
        start_reg[543]) );
  DFF \start_reg_reg[544]  ( .D(start_in[543]), .CLK(clk), .RST(rst), .Q(
        start_reg[544]) );
  DFF \start_reg_reg[545]  ( .D(start_in[544]), .CLK(clk), .RST(rst), .Q(
        start_reg[545]) );
  DFF \start_reg_reg[546]  ( .D(start_in[545]), .CLK(clk), .RST(rst), .Q(
        start_reg[546]) );
  DFF \start_reg_reg[547]  ( .D(start_in[546]), .CLK(clk), .RST(rst), .Q(
        start_reg[547]) );
  DFF \start_reg_reg[548]  ( .D(start_in[547]), .CLK(clk), .RST(rst), .Q(
        start_reg[548]) );
  DFF \start_reg_reg[549]  ( .D(start_in[548]), .CLK(clk), .RST(rst), .Q(
        start_reg[549]) );
  DFF \start_reg_reg[550]  ( .D(start_in[549]), .CLK(clk), .RST(rst), .Q(
        start_reg[550]) );
  DFF \start_reg_reg[551]  ( .D(start_in[550]), .CLK(clk), .RST(rst), .Q(
        start_reg[551]) );
  DFF \start_reg_reg[552]  ( .D(start_in[551]), .CLK(clk), .RST(rst), .Q(
        start_reg[552]) );
  DFF \start_reg_reg[553]  ( .D(start_in[552]), .CLK(clk), .RST(rst), .Q(
        start_reg[553]) );
  DFF \start_reg_reg[554]  ( .D(start_in[553]), .CLK(clk), .RST(rst), .Q(
        start_reg[554]) );
  DFF \start_reg_reg[555]  ( .D(start_in[554]), .CLK(clk), .RST(rst), .Q(
        start_reg[555]) );
  DFF \start_reg_reg[556]  ( .D(start_in[555]), .CLK(clk), .RST(rst), .Q(
        start_reg[556]) );
  DFF \start_reg_reg[557]  ( .D(start_in[556]), .CLK(clk), .RST(rst), .Q(
        start_reg[557]) );
  DFF \start_reg_reg[558]  ( .D(start_in[557]), .CLK(clk), .RST(rst), .Q(
        start_reg[558]) );
  DFF \start_reg_reg[559]  ( .D(start_in[558]), .CLK(clk), .RST(rst), .Q(
        start_reg[559]) );
  DFF \start_reg_reg[560]  ( .D(start_in[559]), .CLK(clk), .RST(rst), .Q(
        start_reg[560]) );
  DFF \start_reg_reg[561]  ( .D(start_in[560]), .CLK(clk), .RST(rst), .Q(
        start_reg[561]) );
  DFF \start_reg_reg[562]  ( .D(start_in[561]), .CLK(clk), .RST(rst), .Q(
        start_reg[562]) );
  DFF \start_reg_reg[563]  ( .D(start_in[562]), .CLK(clk), .RST(rst), .Q(
        start_reg[563]) );
  DFF \start_reg_reg[564]  ( .D(start_in[563]), .CLK(clk), .RST(rst), .Q(
        start_reg[564]) );
  DFF \start_reg_reg[565]  ( .D(start_in[564]), .CLK(clk), .RST(rst), .Q(
        start_reg[565]) );
  DFF \start_reg_reg[566]  ( .D(start_in[565]), .CLK(clk), .RST(rst), .Q(
        start_reg[566]) );
  DFF \start_reg_reg[567]  ( .D(start_in[566]), .CLK(clk), .RST(rst), .Q(
        start_reg[567]) );
  DFF \start_reg_reg[568]  ( .D(start_in[567]), .CLK(clk), .RST(rst), .Q(
        start_reg[568]) );
  DFF \start_reg_reg[569]  ( .D(start_in[568]), .CLK(clk), .RST(rst), .Q(
        start_reg[569]) );
  DFF \start_reg_reg[570]  ( .D(start_in[569]), .CLK(clk), .RST(rst), .Q(
        start_reg[570]) );
  DFF \start_reg_reg[571]  ( .D(start_in[570]), .CLK(clk), .RST(rst), .Q(
        start_reg[571]) );
  DFF \start_reg_reg[572]  ( .D(start_in[571]), .CLK(clk), .RST(rst), .Q(
        start_reg[572]) );
  DFF \start_reg_reg[573]  ( .D(start_in[572]), .CLK(clk), .RST(rst), .Q(
        start_reg[573]) );
  DFF \start_reg_reg[574]  ( .D(start_in[573]), .CLK(clk), .RST(rst), .Q(
        start_reg[574]) );
  DFF \start_reg_reg[575]  ( .D(start_in[574]), .CLK(clk), .RST(rst), .Q(
        start_reg[575]) );
  DFF \start_reg_reg[576]  ( .D(start_in[575]), .CLK(clk), .RST(rst), .Q(
        start_reg[576]) );
  DFF \start_reg_reg[577]  ( .D(start_in[576]), .CLK(clk), .RST(rst), .Q(
        start_reg[577]) );
  DFF \start_reg_reg[578]  ( .D(start_in[577]), .CLK(clk), .RST(rst), .Q(
        start_reg[578]) );
  DFF \start_reg_reg[579]  ( .D(start_in[578]), .CLK(clk), .RST(rst), .Q(
        start_reg[579]) );
  DFF \start_reg_reg[580]  ( .D(start_in[579]), .CLK(clk), .RST(rst), .Q(
        start_reg[580]) );
  DFF \start_reg_reg[581]  ( .D(start_in[580]), .CLK(clk), .RST(rst), .Q(
        start_reg[581]) );
  DFF \start_reg_reg[582]  ( .D(start_in[581]), .CLK(clk), .RST(rst), .Q(
        start_reg[582]) );
  DFF \start_reg_reg[583]  ( .D(start_in[582]), .CLK(clk), .RST(rst), .Q(
        start_reg[583]) );
  DFF \start_reg_reg[584]  ( .D(start_in[583]), .CLK(clk), .RST(rst), .Q(
        start_reg[584]) );
  DFF \start_reg_reg[585]  ( .D(start_in[584]), .CLK(clk), .RST(rst), .Q(
        start_reg[585]) );
  DFF \start_reg_reg[586]  ( .D(start_in[585]), .CLK(clk), .RST(rst), .Q(
        start_reg[586]) );
  DFF \start_reg_reg[587]  ( .D(start_in[586]), .CLK(clk), .RST(rst), .Q(
        start_reg[587]) );
  DFF \start_reg_reg[588]  ( .D(start_in[587]), .CLK(clk), .RST(rst), .Q(
        start_reg[588]) );
  DFF \start_reg_reg[589]  ( .D(start_in[588]), .CLK(clk), .RST(rst), .Q(
        start_reg[589]) );
  DFF \start_reg_reg[590]  ( .D(start_in[589]), .CLK(clk), .RST(rst), .Q(
        start_reg[590]) );
  DFF \start_reg_reg[591]  ( .D(start_in[590]), .CLK(clk), .RST(rst), .Q(
        start_reg[591]) );
  DFF \start_reg_reg[592]  ( .D(start_in[591]), .CLK(clk), .RST(rst), .Q(
        start_reg[592]) );
  DFF \start_reg_reg[593]  ( .D(start_in[592]), .CLK(clk), .RST(rst), .Q(
        start_reg[593]) );
  DFF \start_reg_reg[594]  ( .D(start_in[593]), .CLK(clk), .RST(rst), .Q(
        start_reg[594]) );
  DFF \start_reg_reg[595]  ( .D(start_in[594]), .CLK(clk), .RST(rst), .Q(
        start_reg[595]) );
  DFF \start_reg_reg[596]  ( .D(start_in[595]), .CLK(clk), .RST(rst), .Q(
        start_reg[596]) );
  DFF \start_reg_reg[597]  ( .D(start_in[596]), .CLK(clk), .RST(rst), .Q(
        start_reg[597]) );
  DFF \start_reg_reg[598]  ( .D(start_in[597]), .CLK(clk), .RST(rst), .Q(
        start_reg[598]) );
  DFF \start_reg_reg[599]  ( .D(start_in[598]), .CLK(clk), .RST(rst), .Q(
        start_reg[599]) );
  DFF \start_reg_reg[600]  ( .D(start_in[599]), .CLK(clk), .RST(rst), .Q(
        start_reg[600]) );
  DFF \start_reg_reg[601]  ( .D(start_in[600]), .CLK(clk), .RST(rst), .Q(
        start_reg[601]) );
  DFF \start_reg_reg[602]  ( .D(start_in[601]), .CLK(clk), .RST(rst), .Q(
        start_reg[602]) );
  DFF \start_reg_reg[603]  ( .D(start_in[602]), .CLK(clk), .RST(rst), .Q(
        start_reg[603]) );
  DFF \start_reg_reg[604]  ( .D(start_in[603]), .CLK(clk), .RST(rst), .Q(
        start_reg[604]) );
  DFF \start_reg_reg[605]  ( .D(start_in[604]), .CLK(clk), .RST(rst), .Q(
        start_reg[605]) );
  DFF \start_reg_reg[606]  ( .D(start_in[605]), .CLK(clk), .RST(rst), .Q(
        start_reg[606]) );
  DFF \start_reg_reg[607]  ( .D(start_in[606]), .CLK(clk), .RST(rst), .Q(
        start_reg[607]) );
  DFF \start_reg_reg[608]  ( .D(start_in[607]), .CLK(clk), .RST(rst), .Q(
        start_reg[608]) );
  DFF \start_reg_reg[609]  ( .D(start_in[608]), .CLK(clk), .RST(rst), .Q(
        start_reg[609]) );
  DFF \start_reg_reg[610]  ( .D(start_in[609]), .CLK(clk), .RST(rst), .Q(
        start_reg[610]) );
  DFF \start_reg_reg[611]  ( .D(start_in[610]), .CLK(clk), .RST(rst), .Q(
        start_reg[611]) );
  DFF \start_reg_reg[612]  ( .D(start_in[611]), .CLK(clk), .RST(rst), .Q(
        start_reg[612]) );
  DFF \start_reg_reg[613]  ( .D(start_in[612]), .CLK(clk), .RST(rst), .Q(
        start_reg[613]) );
  DFF \start_reg_reg[614]  ( .D(start_in[613]), .CLK(clk), .RST(rst), .Q(
        start_reg[614]) );
  DFF \start_reg_reg[615]  ( .D(start_in[614]), .CLK(clk), .RST(rst), .Q(
        start_reg[615]) );
  DFF \start_reg_reg[616]  ( .D(start_in[615]), .CLK(clk), .RST(rst), .Q(
        start_reg[616]) );
  DFF \start_reg_reg[617]  ( .D(start_in[616]), .CLK(clk), .RST(rst), .Q(
        start_reg[617]) );
  DFF \start_reg_reg[618]  ( .D(start_in[617]), .CLK(clk), .RST(rst), .Q(
        start_reg[618]) );
  DFF \start_reg_reg[619]  ( .D(start_in[618]), .CLK(clk), .RST(rst), .Q(
        start_reg[619]) );
  DFF \start_reg_reg[620]  ( .D(start_in[619]), .CLK(clk), .RST(rst), .Q(
        start_reg[620]) );
  DFF \start_reg_reg[621]  ( .D(start_in[620]), .CLK(clk), .RST(rst), .Q(
        start_reg[621]) );
  DFF \start_reg_reg[622]  ( .D(start_in[621]), .CLK(clk), .RST(rst), .Q(
        start_reg[622]) );
  DFF \start_reg_reg[623]  ( .D(start_in[622]), .CLK(clk), .RST(rst), .Q(
        start_reg[623]) );
  DFF \start_reg_reg[624]  ( .D(start_in[623]), .CLK(clk), .RST(rst), .Q(
        start_reg[624]) );
  DFF \start_reg_reg[625]  ( .D(start_in[624]), .CLK(clk), .RST(rst), .Q(
        start_reg[625]) );
  DFF \start_reg_reg[626]  ( .D(start_in[625]), .CLK(clk), .RST(rst), .Q(
        start_reg[626]) );
  DFF \start_reg_reg[627]  ( .D(start_in[626]), .CLK(clk), .RST(rst), .Q(
        start_reg[627]) );
  DFF \start_reg_reg[628]  ( .D(start_in[627]), .CLK(clk), .RST(rst), .Q(
        start_reg[628]) );
  DFF \start_reg_reg[629]  ( .D(start_in[628]), .CLK(clk), .RST(rst), .Q(
        start_reg[629]) );
  DFF \start_reg_reg[630]  ( .D(start_in[629]), .CLK(clk), .RST(rst), .Q(
        start_reg[630]) );
  DFF \start_reg_reg[631]  ( .D(start_in[630]), .CLK(clk), .RST(rst), .Q(
        start_reg[631]) );
  DFF \start_reg_reg[632]  ( .D(start_in[631]), .CLK(clk), .RST(rst), .Q(
        start_reg[632]) );
  DFF \start_reg_reg[633]  ( .D(start_in[632]), .CLK(clk), .RST(rst), .Q(
        start_reg[633]) );
  DFF \start_reg_reg[634]  ( .D(start_in[633]), .CLK(clk), .RST(rst), .Q(
        start_reg[634]) );
  DFF \start_reg_reg[635]  ( .D(start_in[634]), .CLK(clk), .RST(rst), .Q(
        start_reg[635]) );
  DFF \start_reg_reg[636]  ( .D(start_in[635]), .CLK(clk), .RST(rst), .Q(
        start_reg[636]) );
  DFF \start_reg_reg[637]  ( .D(start_in[636]), .CLK(clk), .RST(rst), .Q(
        start_reg[637]) );
  DFF \start_reg_reg[638]  ( .D(start_in[637]), .CLK(clk), .RST(rst), .Q(
        start_reg[638]) );
  DFF \start_reg_reg[639]  ( .D(start_in[638]), .CLK(clk), .RST(rst), .Q(
        start_reg[639]) );
  DFF \start_reg_reg[640]  ( .D(start_in[639]), .CLK(clk), .RST(rst), .Q(
        start_reg[640]) );
  DFF \start_reg_reg[641]  ( .D(start_in[640]), .CLK(clk), .RST(rst), .Q(
        start_reg[641]) );
  DFF \start_reg_reg[642]  ( .D(start_in[641]), .CLK(clk), .RST(rst), .Q(
        start_reg[642]) );
  DFF \start_reg_reg[643]  ( .D(start_in[642]), .CLK(clk), .RST(rst), .Q(
        start_reg[643]) );
  DFF \start_reg_reg[644]  ( .D(start_in[643]), .CLK(clk), .RST(rst), .Q(
        start_reg[644]) );
  DFF \start_reg_reg[645]  ( .D(start_in[644]), .CLK(clk), .RST(rst), .Q(
        start_reg[645]) );
  DFF \start_reg_reg[646]  ( .D(start_in[645]), .CLK(clk), .RST(rst), .Q(
        start_reg[646]) );
  DFF \start_reg_reg[647]  ( .D(start_in[646]), .CLK(clk), .RST(rst), .Q(
        start_reg[647]) );
  DFF \start_reg_reg[648]  ( .D(start_in[647]), .CLK(clk), .RST(rst), .Q(
        start_reg[648]) );
  DFF \start_reg_reg[649]  ( .D(start_in[648]), .CLK(clk), .RST(rst), .Q(
        start_reg[649]) );
  DFF \start_reg_reg[650]  ( .D(start_in[649]), .CLK(clk), .RST(rst), .Q(
        start_reg[650]) );
  DFF \start_reg_reg[651]  ( .D(start_in[650]), .CLK(clk), .RST(rst), .Q(
        start_reg[651]) );
  DFF \start_reg_reg[652]  ( .D(start_in[651]), .CLK(clk), .RST(rst), .Q(
        start_reg[652]) );
  DFF \start_reg_reg[653]  ( .D(start_in[652]), .CLK(clk), .RST(rst), .Q(
        start_reg[653]) );
  DFF \start_reg_reg[654]  ( .D(start_in[653]), .CLK(clk), .RST(rst), .Q(
        start_reg[654]) );
  DFF \start_reg_reg[655]  ( .D(start_in[654]), .CLK(clk), .RST(rst), .Q(
        start_reg[655]) );
  DFF \start_reg_reg[656]  ( .D(start_in[655]), .CLK(clk), .RST(rst), .Q(
        start_reg[656]) );
  DFF \start_reg_reg[657]  ( .D(start_in[656]), .CLK(clk), .RST(rst), .Q(
        start_reg[657]) );
  DFF \start_reg_reg[658]  ( .D(start_in[657]), .CLK(clk), .RST(rst), .Q(
        start_reg[658]) );
  DFF \start_reg_reg[659]  ( .D(start_in[658]), .CLK(clk), .RST(rst), .Q(
        start_reg[659]) );
  DFF \start_reg_reg[660]  ( .D(start_in[659]), .CLK(clk), .RST(rst), .Q(
        start_reg[660]) );
  DFF \start_reg_reg[661]  ( .D(start_in[660]), .CLK(clk), .RST(rst), .Q(
        start_reg[661]) );
  DFF \start_reg_reg[662]  ( .D(start_in[661]), .CLK(clk), .RST(rst), .Q(
        start_reg[662]) );
  DFF \start_reg_reg[663]  ( .D(start_in[662]), .CLK(clk), .RST(rst), .Q(
        start_reg[663]) );
  DFF \start_reg_reg[664]  ( .D(start_in[663]), .CLK(clk), .RST(rst), .Q(
        start_reg[664]) );
  DFF \start_reg_reg[665]  ( .D(start_in[664]), .CLK(clk), .RST(rst), .Q(
        start_reg[665]) );
  DFF \start_reg_reg[666]  ( .D(start_in[665]), .CLK(clk), .RST(rst), .Q(
        start_reg[666]) );
  DFF \start_reg_reg[667]  ( .D(start_in[666]), .CLK(clk), .RST(rst), .Q(
        start_reg[667]) );
  DFF \start_reg_reg[668]  ( .D(start_in[667]), .CLK(clk), .RST(rst), .Q(
        start_reg[668]) );
  DFF \start_reg_reg[669]  ( .D(start_in[668]), .CLK(clk), .RST(rst), .Q(
        start_reg[669]) );
  DFF \start_reg_reg[670]  ( .D(start_in[669]), .CLK(clk), .RST(rst), .Q(
        start_reg[670]) );
  DFF \start_reg_reg[671]  ( .D(start_in[670]), .CLK(clk), .RST(rst), .Q(
        start_reg[671]) );
  DFF \start_reg_reg[672]  ( .D(start_in[671]), .CLK(clk), .RST(rst), .Q(
        start_reg[672]) );
  DFF \start_reg_reg[673]  ( .D(start_in[672]), .CLK(clk), .RST(rst), .Q(
        start_reg[673]) );
  DFF \start_reg_reg[674]  ( .D(start_in[673]), .CLK(clk), .RST(rst), .Q(
        start_reg[674]) );
  DFF \start_reg_reg[675]  ( .D(start_in[674]), .CLK(clk), .RST(rst), .Q(
        start_reg[675]) );
  DFF \start_reg_reg[676]  ( .D(start_in[675]), .CLK(clk), .RST(rst), .Q(
        start_reg[676]) );
  DFF \start_reg_reg[677]  ( .D(start_in[676]), .CLK(clk), .RST(rst), .Q(
        start_reg[677]) );
  DFF \start_reg_reg[678]  ( .D(start_in[677]), .CLK(clk), .RST(rst), .Q(
        start_reg[678]) );
  DFF \start_reg_reg[679]  ( .D(start_in[678]), .CLK(clk), .RST(rst), .Q(
        start_reg[679]) );
  DFF \start_reg_reg[680]  ( .D(start_in[679]), .CLK(clk), .RST(rst), .Q(
        start_reg[680]) );
  DFF \start_reg_reg[681]  ( .D(start_in[680]), .CLK(clk), .RST(rst), .Q(
        start_reg[681]) );
  DFF \start_reg_reg[682]  ( .D(start_in[681]), .CLK(clk), .RST(rst), .Q(
        start_reg[682]) );
  DFF \start_reg_reg[683]  ( .D(start_in[682]), .CLK(clk), .RST(rst), .Q(
        start_reg[683]) );
  DFF \start_reg_reg[684]  ( .D(start_in[683]), .CLK(clk), .RST(rst), .Q(
        start_reg[684]) );
  DFF \start_reg_reg[685]  ( .D(start_in[684]), .CLK(clk), .RST(rst), .Q(
        start_reg[685]) );
  DFF \start_reg_reg[686]  ( .D(start_in[685]), .CLK(clk), .RST(rst), .Q(
        start_reg[686]) );
  DFF \start_reg_reg[687]  ( .D(start_in[686]), .CLK(clk), .RST(rst), .Q(
        start_reg[687]) );
  DFF \start_reg_reg[688]  ( .D(start_in[687]), .CLK(clk), .RST(rst), .Q(
        start_reg[688]) );
  DFF \start_reg_reg[689]  ( .D(start_in[688]), .CLK(clk), .RST(rst), .Q(
        start_reg[689]) );
  DFF \start_reg_reg[690]  ( .D(start_in[689]), .CLK(clk), .RST(rst), .Q(
        start_reg[690]) );
  DFF \start_reg_reg[691]  ( .D(start_in[690]), .CLK(clk), .RST(rst), .Q(
        start_reg[691]) );
  DFF \start_reg_reg[692]  ( .D(start_in[691]), .CLK(clk), .RST(rst), .Q(
        start_reg[692]) );
  DFF \start_reg_reg[693]  ( .D(start_in[692]), .CLK(clk), .RST(rst), .Q(
        start_reg[693]) );
  DFF \start_reg_reg[694]  ( .D(start_in[693]), .CLK(clk), .RST(rst), .Q(
        start_reg[694]) );
  DFF \start_reg_reg[695]  ( .D(start_in[694]), .CLK(clk), .RST(rst), .Q(
        start_reg[695]) );
  DFF \start_reg_reg[696]  ( .D(start_in[695]), .CLK(clk), .RST(rst), .Q(
        start_reg[696]) );
  DFF \start_reg_reg[697]  ( .D(start_in[696]), .CLK(clk), .RST(rst), .Q(
        start_reg[697]) );
  DFF \start_reg_reg[698]  ( .D(start_in[697]), .CLK(clk), .RST(rst), .Q(
        start_reg[698]) );
  DFF \start_reg_reg[699]  ( .D(start_in[698]), .CLK(clk), .RST(rst), .Q(
        start_reg[699]) );
  DFF \start_reg_reg[700]  ( .D(start_in[699]), .CLK(clk), .RST(rst), .Q(
        start_reg[700]) );
  DFF \start_reg_reg[701]  ( .D(start_in[700]), .CLK(clk), .RST(rst), .Q(
        start_reg[701]) );
  DFF \start_reg_reg[702]  ( .D(start_in[701]), .CLK(clk), .RST(rst), .Q(
        start_reg[702]) );
  DFF \start_reg_reg[703]  ( .D(start_in[702]), .CLK(clk), .RST(rst), .Q(
        start_reg[703]) );
  DFF \start_reg_reg[704]  ( .D(start_in[703]), .CLK(clk), .RST(rst), .Q(
        start_reg[704]) );
  DFF \start_reg_reg[705]  ( .D(start_in[704]), .CLK(clk), .RST(rst), .Q(
        start_reg[705]) );
  DFF \start_reg_reg[706]  ( .D(start_in[705]), .CLK(clk), .RST(rst), .Q(
        start_reg[706]) );
  DFF \start_reg_reg[707]  ( .D(start_in[706]), .CLK(clk), .RST(rst), .Q(
        start_reg[707]) );
  DFF \start_reg_reg[708]  ( .D(start_in[707]), .CLK(clk), .RST(rst), .Q(
        start_reg[708]) );
  DFF \start_reg_reg[709]  ( .D(start_in[708]), .CLK(clk), .RST(rst), .Q(
        start_reg[709]) );
  DFF \start_reg_reg[710]  ( .D(start_in[709]), .CLK(clk), .RST(rst), .Q(
        start_reg[710]) );
  DFF \start_reg_reg[711]  ( .D(start_in[710]), .CLK(clk), .RST(rst), .Q(
        start_reg[711]) );
  DFF \start_reg_reg[712]  ( .D(start_in[711]), .CLK(clk), .RST(rst), .Q(
        start_reg[712]) );
  DFF \start_reg_reg[713]  ( .D(start_in[712]), .CLK(clk), .RST(rst), .Q(
        start_reg[713]) );
  DFF \start_reg_reg[714]  ( .D(start_in[713]), .CLK(clk), .RST(rst), .Q(
        start_reg[714]) );
  DFF \start_reg_reg[715]  ( .D(start_in[714]), .CLK(clk), .RST(rst), .Q(
        start_reg[715]) );
  DFF \start_reg_reg[716]  ( .D(start_in[715]), .CLK(clk), .RST(rst), .Q(
        start_reg[716]) );
  DFF \start_reg_reg[717]  ( .D(start_in[716]), .CLK(clk), .RST(rst), .Q(
        start_reg[717]) );
  DFF \start_reg_reg[718]  ( .D(start_in[717]), .CLK(clk), .RST(rst), .Q(
        start_reg[718]) );
  DFF \start_reg_reg[719]  ( .D(start_in[718]), .CLK(clk), .RST(rst), .Q(
        start_reg[719]) );
  DFF \start_reg_reg[720]  ( .D(start_in[719]), .CLK(clk), .RST(rst), .Q(
        start_reg[720]) );
  DFF \start_reg_reg[721]  ( .D(start_in[720]), .CLK(clk), .RST(rst), .Q(
        start_reg[721]) );
  DFF \start_reg_reg[722]  ( .D(start_in[721]), .CLK(clk), .RST(rst), .Q(
        start_reg[722]) );
  DFF \start_reg_reg[723]  ( .D(start_in[722]), .CLK(clk), .RST(rst), .Q(
        start_reg[723]) );
  DFF \start_reg_reg[724]  ( .D(start_in[723]), .CLK(clk), .RST(rst), .Q(
        start_reg[724]) );
  DFF \start_reg_reg[725]  ( .D(start_in[724]), .CLK(clk), .RST(rst), .Q(
        start_reg[725]) );
  DFF \start_reg_reg[726]  ( .D(start_in[725]), .CLK(clk), .RST(rst), .Q(
        start_reg[726]) );
  DFF \start_reg_reg[727]  ( .D(start_in[726]), .CLK(clk), .RST(rst), .Q(
        start_reg[727]) );
  DFF \start_reg_reg[728]  ( .D(start_in[727]), .CLK(clk), .RST(rst), .Q(
        start_reg[728]) );
  DFF \start_reg_reg[729]  ( .D(start_in[728]), .CLK(clk), .RST(rst), .Q(
        start_reg[729]) );
  DFF \start_reg_reg[730]  ( .D(start_in[729]), .CLK(clk), .RST(rst), .Q(
        start_reg[730]) );
  DFF \start_reg_reg[731]  ( .D(start_in[730]), .CLK(clk), .RST(rst), .Q(
        start_reg[731]) );
  DFF \start_reg_reg[732]  ( .D(start_in[731]), .CLK(clk), .RST(rst), .Q(
        start_reg[732]) );
  DFF \start_reg_reg[733]  ( .D(start_in[732]), .CLK(clk), .RST(rst), .Q(
        start_reg[733]) );
  DFF \start_reg_reg[734]  ( .D(start_in[733]), .CLK(clk), .RST(rst), .Q(
        start_reg[734]) );
  DFF \start_reg_reg[735]  ( .D(start_in[734]), .CLK(clk), .RST(rst), .Q(
        start_reg[735]) );
  DFF \start_reg_reg[736]  ( .D(start_in[735]), .CLK(clk), .RST(rst), .Q(
        start_reg[736]) );
  DFF \start_reg_reg[737]  ( .D(start_in[736]), .CLK(clk), .RST(rst), .Q(
        start_reg[737]) );
  DFF \start_reg_reg[738]  ( .D(start_in[737]), .CLK(clk), .RST(rst), .Q(
        start_reg[738]) );
  DFF \start_reg_reg[739]  ( .D(start_in[738]), .CLK(clk), .RST(rst), .Q(
        start_reg[739]) );
  DFF \start_reg_reg[740]  ( .D(start_in[739]), .CLK(clk), .RST(rst), .Q(
        start_reg[740]) );
  DFF \start_reg_reg[741]  ( .D(start_in[740]), .CLK(clk), .RST(rst), .Q(
        start_reg[741]) );
  DFF \start_reg_reg[742]  ( .D(start_in[741]), .CLK(clk), .RST(rst), .Q(
        start_reg[742]) );
  DFF \start_reg_reg[743]  ( .D(start_in[742]), .CLK(clk), .RST(rst), .Q(
        start_reg[743]) );
  DFF \start_reg_reg[744]  ( .D(start_in[743]), .CLK(clk), .RST(rst), .Q(
        start_reg[744]) );
  DFF \start_reg_reg[745]  ( .D(start_in[744]), .CLK(clk), .RST(rst), .Q(
        start_reg[745]) );
  DFF \start_reg_reg[746]  ( .D(start_in[745]), .CLK(clk), .RST(rst), .Q(
        start_reg[746]) );
  DFF \start_reg_reg[747]  ( .D(start_in[746]), .CLK(clk), .RST(rst), .Q(
        start_reg[747]) );
  DFF \start_reg_reg[748]  ( .D(start_in[747]), .CLK(clk), .RST(rst), .Q(
        start_reg[748]) );
  DFF \start_reg_reg[749]  ( .D(start_in[748]), .CLK(clk), .RST(rst), .Q(
        start_reg[749]) );
  DFF \start_reg_reg[750]  ( .D(start_in[749]), .CLK(clk), .RST(rst), .Q(
        start_reg[750]) );
  DFF \start_reg_reg[751]  ( .D(start_in[750]), .CLK(clk), .RST(rst), .Q(
        start_reg[751]) );
  DFF \start_reg_reg[752]  ( .D(start_in[751]), .CLK(clk), .RST(rst), .Q(
        start_reg[752]) );
  DFF \start_reg_reg[753]  ( .D(start_in[752]), .CLK(clk), .RST(rst), .Q(
        start_reg[753]) );
  DFF \start_reg_reg[754]  ( .D(start_in[753]), .CLK(clk), .RST(rst), .Q(
        start_reg[754]) );
  DFF \start_reg_reg[755]  ( .D(start_in[754]), .CLK(clk), .RST(rst), .Q(
        start_reg[755]) );
  DFF \start_reg_reg[756]  ( .D(start_in[755]), .CLK(clk), .RST(rst), .Q(
        start_reg[756]) );
  DFF \start_reg_reg[757]  ( .D(start_in[756]), .CLK(clk), .RST(rst), .Q(
        start_reg[757]) );
  DFF \start_reg_reg[758]  ( .D(start_in[757]), .CLK(clk), .RST(rst), .Q(
        start_reg[758]) );
  DFF \start_reg_reg[759]  ( .D(start_in[758]), .CLK(clk), .RST(rst), .Q(
        start_reg[759]) );
  DFF \start_reg_reg[760]  ( .D(start_in[759]), .CLK(clk), .RST(rst), .Q(
        start_reg[760]) );
  DFF \start_reg_reg[761]  ( .D(start_in[760]), .CLK(clk), .RST(rst), .Q(
        start_reg[761]) );
  DFF \start_reg_reg[762]  ( .D(start_in[761]), .CLK(clk), .RST(rst), .Q(
        start_reg[762]) );
  DFF \start_reg_reg[763]  ( .D(start_in[762]), .CLK(clk), .RST(rst), .Q(
        start_reg[763]) );
  DFF \start_reg_reg[764]  ( .D(start_in[763]), .CLK(clk), .RST(rst), .Q(
        start_reg[764]) );
  DFF \start_reg_reg[765]  ( .D(start_in[764]), .CLK(clk), .RST(rst), .Q(
        start_reg[765]) );
  DFF \start_reg_reg[766]  ( .D(start_in[765]), .CLK(clk), .RST(rst), .Q(
        start_reg[766]) );
  DFF \start_reg_reg[767]  ( .D(start_in[766]), .CLK(clk), .RST(rst), .Q(
        start_reg[767]) );
  DFF \start_reg_reg[768]  ( .D(start_in[767]), .CLK(clk), .RST(rst), .Q(
        start_reg[768]) );
  DFF \start_reg_reg[769]  ( .D(start_in[768]), .CLK(clk), .RST(rst), .Q(
        start_reg[769]) );
  DFF \start_reg_reg[770]  ( .D(start_in[769]), .CLK(clk), .RST(rst), .Q(
        start_reg[770]) );
  DFF \start_reg_reg[771]  ( .D(start_in[770]), .CLK(clk), .RST(rst), .Q(
        start_reg[771]) );
  DFF \start_reg_reg[772]  ( .D(start_in[771]), .CLK(clk), .RST(rst), .Q(
        start_reg[772]) );
  DFF \start_reg_reg[773]  ( .D(start_in[772]), .CLK(clk), .RST(rst), .Q(
        start_reg[773]) );
  DFF \start_reg_reg[774]  ( .D(start_in[773]), .CLK(clk), .RST(rst), .Q(
        start_reg[774]) );
  DFF \start_reg_reg[775]  ( .D(start_in[774]), .CLK(clk), .RST(rst), .Q(
        start_reg[775]) );
  DFF \start_reg_reg[776]  ( .D(start_in[775]), .CLK(clk), .RST(rst), .Q(
        start_reg[776]) );
  DFF \start_reg_reg[777]  ( .D(start_in[776]), .CLK(clk), .RST(rst), .Q(
        start_reg[777]) );
  DFF \start_reg_reg[778]  ( .D(start_in[777]), .CLK(clk), .RST(rst), .Q(
        start_reg[778]) );
  DFF \start_reg_reg[779]  ( .D(start_in[778]), .CLK(clk), .RST(rst), .Q(
        start_reg[779]) );
  DFF \start_reg_reg[780]  ( .D(start_in[779]), .CLK(clk), .RST(rst), .Q(
        start_reg[780]) );
  DFF \start_reg_reg[781]  ( .D(start_in[780]), .CLK(clk), .RST(rst), .Q(
        start_reg[781]) );
  DFF \start_reg_reg[782]  ( .D(start_in[781]), .CLK(clk), .RST(rst), .Q(
        start_reg[782]) );
  DFF \start_reg_reg[783]  ( .D(start_in[782]), .CLK(clk), .RST(rst), .Q(
        start_reg[783]) );
  DFF \start_reg_reg[784]  ( .D(start_in[783]), .CLK(clk), .RST(rst), .Q(
        start_reg[784]) );
  DFF \start_reg_reg[785]  ( .D(start_in[784]), .CLK(clk), .RST(rst), .Q(
        start_reg[785]) );
  DFF \start_reg_reg[786]  ( .D(start_in[785]), .CLK(clk), .RST(rst), .Q(
        start_reg[786]) );
  DFF \start_reg_reg[787]  ( .D(start_in[786]), .CLK(clk), .RST(rst), .Q(
        start_reg[787]) );
  DFF \start_reg_reg[788]  ( .D(start_in[787]), .CLK(clk), .RST(rst), .Q(
        start_reg[788]) );
  DFF \start_reg_reg[789]  ( .D(start_in[788]), .CLK(clk), .RST(rst), .Q(
        start_reg[789]) );
  DFF \start_reg_reg[790]  ( .D(start_in[789]), .CLK(clk), .RST(rst), .Q(
        start_reg[790]) );
  DFF \start_reg_reg[791]  ( .D(start_in[790]), .CLK(clk), .RST(rst), .Q(
        start_reg[791]) );
  DFF \start_reg_reg[792]  ( .D(start_in[791]), .CLK(clk), .RST(rst), .Q(
        start_reg[792]) );
  DFF \start_reg_reg[793]  ( .D(start_in[792]), .CLK(clk), .RST(rst), .Q(
        start_reg[793]) );
  DFF \start_reg_reg[794]  ( .D(start_in[793]), .CLK(clk), .RST(rst), .Q(
        start_reg[794]) );
  DFF \start_reg_reg[795]  ( .D(start_in[794]), .CLK(clk), .RST(rst), .Q(
        start_reg[795]) );
  DFF \start_reg_reg[796]  ( .D(start_in[795]), .CLK(clk), .RST(rst), .Q(
        start_reg[796]) );
  DFF \start_reg_reg[797]  ( .D(start_in[796]), .CLK(clk), .RST(rst), .Q(
        start_reg[797]) );
  DFF \start_reg_reg[798]  ( .D(start_in[797]), .CLK(clk), .RST(rst), .Q(
        start_reg[798]) );
  DFF \start_reg_reg[799]  ( .D(start_in[798]), .CLK(clk), .RST(rst), .Q(
        start_reg[799]) );
  DFF \start_reg_reg[800]  ( .D(start_in[799]), .CLK(clk), .RST(rst), .Q(
        start_reg[800]) );
  DFF \start_reg_reg[801]  ( .D(start_in[800]), .CLK(clk), .RST(rst), .Q(
        start_reg[801]) );
  DFF \start_reg_reg[802]  ( .D(start_in[801]), .CLK(clk), .RST(rst), .Q(
        start_reg[802]) );
  DFF \start_reg_reg[803]  ( .D(start_in[802]), .CLK(clk), .RST(rst), .Q(
        start_reg[803]) );
  DFF \start_reg_reg[804]  ( .D(start_in[803]), .CLK(clk), .RST(rst), .Q(
        start_reg[804]) );
  DFF \start_reg_reg[805]  ( .D(start_in[804]), .CLK(clk), .RST(rst), .Q(
        start_reg[805]) );
  DFF \start_reg_reg[806]  ( .D(start_in[805]), .CLK(clk), .RST(rst), .Q(
        start_reg[806]) );
  DFF \start_reg_reg[807]  ( .D(start_in[806]), .CLK(clk), .RST(rst), .Q(
        start_reg[807]) );
  DFF \start_reg_reg[808]  ( .D(start_in[807]), .CLK(clk), .RST(rst), .Q(
        start_reg[808]) );
  DFF \start_reg_reg[809]  ( .D(start_in[808]), .CLK(clk), .RST(rst), .Q(
        start_reg[809]) );
  DFF \start_reg_reg[810]  ( .D(start_in[809]), .CLK(clk), .RST(rst), .Q(
        start_reg[810]) );
  DFF \start_reg_reg[811]  ( .D(start_in[810]), .CLK(clk), .RST(rst), .Q(
        start_reg[811]) );
  DFF \start_reg_reg[812]  ( .D(start_in[811]), .CLK(clk), .RST(rst), .Q(
        start_reg[812]) );
  DFF \start_reg_reg[813]  ( .D(start_in[812]), .CLK(clk), .RST(rst), .Q(
        start_reg[813]) );
  DFF \start_reg_reg[814]  ( .D(start_in[813]), .CLK(clk), .RST(rst), .Q(
        start_reg[814]) );
  DFF \start_reg_reg[815]  ( .D(start_in[814]), .CLK(clk), .RST(rst), .Q(
        start_reg[815]) );
  DFF \start_reg_reg[816]  ( .D(start_in[815]), .CLK(clk), .RST(rst), .Q(
        start_reg[816]) );
  DFF \start_reg_reg[817]  ( .D(start_in[816]), .CLK(clk), .RST(rst), .Q(
        start_reg[817]) );
  DFF \start_reg_reg[818]  ( .D(start_in[817]), .CLK(clk), .RST(rst), .Q(
        start_reg[818]) );
  DFF \start_reg_reg[819]  ( .D(start_in[818]), .CLK(clk), .RST(rst), .Q(
        start_reg[819]) );
  DFF \start_reg_reg[820]  ( .D(start_in[819]), .CLK(clk), .RST(rst), .Q(
        start_reg[820]) );
  DFF \start_reg_reg[821]  ( .D(start_in[820]), .CLK(clk), .RST(rst), .Q(
        start_reg[821]) );
  DFF \start_reg_reg[822]  ( .D(start_in[821]), .CLK(clk), .RST(rst), .Q(
        start_reg[822]) );
  DFF \start_reg_reg[823]  ( .D(start_in[822]), .CLK(clk), .RST(rst), .Q(
        start_reg[823]) );
  DFF \start_reg_reg[824]  ( .D(start_in[823]), .CLK(clk), .RST(rst), .Q(
        start_reg[824]) );
  DFF \start_reg_reg[825]  ( .D(start_in[824]), .CLK(clk), .RST(rst), .Q(
        start_reg[825]) );
  DFF \start_reg_reg[826]  ( .D(start_in[825]), .CLK(clk), .RST(rst), .Q(
        start_reg[826]) );
  DFF \start_reg_reg[827]  ( .D(start_in[826]), .CLK(clk), .RST(rst), .Q(
        start_reg[827]) );
  DFF \start_reg_reg[828]  ( .D(start_in[827]), .CLK(clk), .RST(rst), .Q(
        start_reg[828]) );
  DFF \start_reg_reg[829]  ( .D(start_in[828]), .CLK(clk), .RST(rst), .Q(
        start_reg[829]) );
  DFF \start_reg_reg[830]  ( .D(start_in[829]), .CLK(clk), .RST(rst), .Q(
        start_reg[830]) );
  DFF \start_reg_reg[831]  ( .D(start_in[830]), .CLK(clk), .RST(rst), .Q(
        start_reg[831]) );
  DFF \start_reg_reg[832]  ( .D(start_in[831]), .CLK(clk), .RST(rst), .Q(
        start_reg[832]) );
  DFF \start_reg_reg[833]  ( .D(start_in[832]), .CLK(clk), .RST(rst), .Q(
        start_reg[833]) );
  DFF \start_reg_reg[834]  ( .D(start_in[833]), .CLK(clk), .RST(rst), .Q(
        start_reg[834]) );
  DFF \start_reg_reg[835]  ( .D(start_in[834]), .CLK(clk), .RST(rst), .Q(
        start_reg[835]) );
  DFF \start_reg_reg[836]  ( .D(start_in[835]), .CLK(clk), .RST(rst), .Q(
        start_reg[836]) );
  DFF \start_reg_reg[837]  ( .D(start_in[836]), .CLK(clk), .RST(rst), .Q(
        start_reg[837]) );
  DFF \start_reg_reg[838]  ( .D(start_in[837]), .CLK(clk), .RST(rst), .Q(
        start_reg[838]) );
  DFF \start_reg_reg[839]  ( .D(start_in[838]), .CLK(clk), .RST(rst), .Q(
        start_reg[839]) );
  DFF \start_reg_reg[840]  ( .D(start_in[839]), .CLK(clk), .RST(rst), .Q(
        start_reg[840]) );
  DFF \start_reg_reg[841]  ( .D(start_in[840]), .CLK(clk), .RST(rst), .Q(
        start_reg[841]) );
  DFF \start_reg_reg[842]  ( .D(start_in[841]), .CLK(clk), .RST(rst), .Q(
        start_reg[842]) );
  DFF \start_reg_reg[843]  ( .D(start_in[842]), .CLK(clk), .RST(rst), .Q(
        start_reg[843]) );
  DFF \start_reg_reg[844]  ( .D(start_in[843]), .CLK(clk), .RST(rst), .Q(
        start_reg[844]) );
  DFF \start_reg_reg[845]  ( .D(start_in[844]), .CLK(clk), .RST(rst), .Q(
        start_reg[845]) );
  DFF \start_reg_reg[846]  ( .D(start_in[845]), .CLK(clk), .RST(rst), .Q(
        start_reg[846]) );
  DFF \start_reg_reg[847]  ( .D(start_in[846]), .CLK(clk), .RST(rst), .Q(
        start_reg[847]) );
  DFF \start_reg_reg[848]  ( .D(start_in[847]), .CLK(clk), .RST(rst), .Q(
        start_reg[848]) );
  DFF \start_reg_reg[849]  ( .D(start_in[848]), .CLK(clk), .RST(rst), .Q(
        start_reg[849]) );
  DFF \start_reg_reg[850]  ( .D(start_in[849]), .CLK(clk), .RST(rst), .Q(
        start_reg[850]) );
  DFF \start_reg_reg[851]  ( .D(start_in[850]), .CLK(clk), .RST(rst), .Q(
        start_reg[851]) );
  DFF \start_reg_reg[852]  ( .D(start_in[851]), .CLK(clk), .RST(rst), .Q(
        start_reg[852]) );
  DFF \start_reg_reg[853]  ( .D(start_in[852]), .CLK(clk), .RST(rst), .Q(
        start_reg[853]) );
  DFF \start_reg_reg[854]  ( .D(start_in[853]), .CLK(clk), .RST(rst), .Q(
        start_reg[854]) );
  DFF \start_reg_reg[855]  ( .D(start_in[854]), .CLK(clk), .RST(rst), .Q(
        start_reg[855]) );
  DFF \start_reg_reg[856]  ( .D(start_in[855]), .CLK(clk), .RST(rst), .Q(
        start_reg[856]) );
  DFF \start_reg_reg[857]  ( .D(start_in[856]), .CLK(clk), .RST(rst), .Q(
        start_reg[857]) );
  DFF \start_reg_reg[858]  ( .D(start_in[857]), .CLK(clk), .RST(rst), .Q(
        start_reg[858]) );
  DFF \start_reg_reg[859]  ( .D(start_in[858]), .CLK(clk), .RST(rst), .Q(
        start_reg[859]) );
  DFF \start_reg_reg[860]  ( .D(start_in[859]), .CLK(clk), .RST(rst), .Q(
        start_reg[860]) );
  DFF \start_reg_reg[861]  ( .D(start_in[860]), .CLK(clk), .RST(rst), .Q(
        start_reg[861]) );
  DFF \start_reg_reg[862]  ( .D(start_in[861]), .CLK(clk), .RST(rst), .Q(
        start_reg[862]) );
  DFF \start_reg_reg[863]  ( .D(start_in[862]), .CLK(clk), .RST(rst), .Q(
        start_reg[863]) );
  DFF \start_reg_reg[864]  ( .D(start_in[863]), .CLK(clk), .RST(rst), .Q(
        start_reg[864]) );
  DFF \start_reg_reg[865]  ( .D(start_in[864]), .CLK(clk), .RST(rst), .Q(
        start_reg[865]) );
  DFF \start_reg_reg[866]  ( .D(start_in[865]), .CLK(clk), .RST(rst), .Q(
        start_reg[866]) );
  DFF \start_reg_reg[867]  ( .D(start_in[866]), .CLK(clk), .RST(rst), .Q(
        start_reg[867]) );
  DFF \start_reg_reg[868]  ( .D(start_in[867]), .CLK(clk), .RST(rst), .Q(
        start_reg[868]) );
  DFF \start_reg_reg[869]  ( .D(start_in[868]), .CLK(clk), .RST(rst), .Q(
        start_reg[869]) );
  DFF \start_reg_reg[870]  ( .D(start_in[869]), .CLK(clk), .RST(rst), .Q(
        start_reg[870]) );
  DFF \start_reg_reg[871]  ( .D(start_in[870]), .CLK(clk), .RST(rst), .Q(
        start_reg[871]) );
  DFF \start_reg_reg[872]  ( .D(start_in[871]), .CLK(clk), .RST(rst), .Q(
        start_reg[872]) );
  DFF \start_reg_reg[873]  ( .D(start_in[872]), .CLK(clk), .RST(rst), .Q(
        start_reg[873]) );
  DFF \start_reg_reg[874]  ( .D(start_in[873]), .CLK(clk), .RST(rst), .Q(
        start_reg[874]) );
  DFF \start_reg_reg[875]  ( .D(start_in[874]), .CLK(clk), .RST(rst), .Q(
        start_reg[875]) );
  DFF \start_reg_reg[876]  ( .D(start_in[875]), .CLK(clk), .RST(rst), .Q(
        start_reg[876]) );
  DFF \start_reg_reg[877]  ( .D(start_in[876]), .CLK(clk), .RST(rst), .Q(
        start_reg[877]) );
  DFF \start_reg_reg[878]  ( .D(start_in[877]), .CLK(clk), .RST(rst), .Q(
        start_reg[878]) );
  DFF \start_reg_reg[879]  ( .D(start_in[878]), .CLK(clk), .RST(rst), .Q(
        start_reg[879]) );
  DFF \start_reg_reg[880]  ( .D(start_in[879]), .CLK(clk), .RST(rst), .Q(
        start_reg[880]) );
  DFF \start_reg_reg[881]  ( .D(start_in[880]), .CLK(clk), .RST(rst), .Q(
        start_reg[881]) );
  DFF \start_reg_reg[882]  ( .D(start_in[881]), .CLK(clk), .RST(rst), .Q(
        start_reg[882]) );
  DFF \start_reg_reg[883]  ( .D(start_in[882]), .CLK(clk), .RST(rst), .Q(
        start_reg[883]) );
  DFF \start_reg_reg[884]  ( .D(start_in[883]), .CLK(clk), .RST(rst), .Q(
        start_reg[884]) );
  DFF \start_reg_reg[885]  ( .D(start_in[884]), .CLK(clk), .RST(rst), .Q(
        start_reg[885]) );
  DFF \start_reg_reg[886]  ( .D(start_in[885]), .CLK(clk), .RST(rst), .Q(
        start_reg[886]) );
  DFF \start_reg_reg[887]  ( .D(start_in[886]), .CLK(clk), .RST(rst), .Q(
        start_reg[887]) );
  DFF \start_reg_reg[888]  ( .D(start_in[887]), .CLK(clk), .RST(rst), .Q(
        start_reg[888]) );
  DFF \start_reg_reg[889]  ( .D(start_in[888]), .CLK(clk), .RST(rst), .Q(
        start_reg[889]) );
  DFF \start_reg_reg[890]  ( .D(start_in[889]), .CLK(clk), .RST(rst), .Q(
        start_reg[890]) );
  DFF \start_reg_reg[891]  ( .D(start_in[890]), .CLK(clk), .RST(rst), .Q(
        start_reg[891]) );
  DFF \start_reg_reg[892]  ( .D(start_in[891]), .CLK(clk), .RST(rst), .Q(
        start_reg[892]) );
  DFF \start_reg_reg[893]  ( .D(start_in[892]), .CLK(clk), .RST(rst), .Q(
        start_reg[893]) );
  DFF \start_reg_reg[894]  ( .D(start_in[893]), .CLK(clk), .RST(rst), .Q(
        start_reg[894]) );
  DFF \start_reg_reg[895]  ( .D(start_in[894]), .CLK(clk), .RST(rst), .Q(
        start_reg[895]) );
  DFF \start_reg_reg[896]  ( .D(start_in[895]), .CLK(clk), .RST(rst), .Q(
        start_reg[896]) );
  DFF \start_reg_reg[897]  ( .D(start_in[896]), .CLK(clk), .RST(rst), .Q(
        start_reg[897]) );
  DFF \start_reg_reg[898]  ( .D(start_in[897]), .CLK(clk), .RST(rst), .Q(
        start_reg[898]) );
  DFF \start_reg_reg[899]  ( .D(start_in[898]), .CLK(clk), .RST(rst), .Q(
        start_reg[899]) );
  DFF \start_reg_reg[900]  ( .D(start_in[899]), .CLK(clk), .RST(rst), .Q(
        start_reg[900]) );
  DFF \start_reg_reg[901]  ( .D(start_in[900]), .CLK(clk), .RST(rst), .Q(
        start_reg[901]) );
  DFF \start_reg_reg[902]  ( .D(start_in[901]), .CLK(clk), .RST(rst), .Q(
        start_reg[902]) );
  DFF \start_reg_reg[903]  ( .D(start_in[902]), .CLK(clk), .RST(rst), .Q(
        start_reg[903]) );
  DFF \start_reg_reg[904]  ( .D(start_in[903]), .CLK(clk), .RST(rst), .Q(
        start_reg[904]) );
  DFF \start_reg_reg[905]  ( .D(start_in[904]), .CLK(clk), .RST(rst), .Q(
        start_reg[905]) );
  DFF \start_reg_reg[906]  ( .D(start_in[905]), .CLK(clk), .RST(rst), .Q(
        start_reg[906]) );
  DFF \start_reg_reg[907]  ( .D(start_in[906]), .CLK(clk), .RST(rst), .Q(
        start_reg[907]) );
  DFF \start_reg_reg[908]  ( .D(start_in[907]), .CLK(clk), .RST(rst), .Q(
        start_reg[908]) );
  DFF \start_reg_reg[909]  ( .D(start_in[908]), .CLK(clk), .RST(rst), .Q(
        start_reg[909]) );
  DFF \start_reg_reg[910]  ( .D(start_in[909]), .CLK(clk), .RST(rst), .Q(
        start_reg[910]) );
  DFF \start_reg_reg[911]  ( .D(start_in[910]), .CLK(clk), .RST(rst), .Q(
        start_reg[911]) );
  DFF \start_reg_reg[912]  ( .D(start_in[911]), .CLK(clk), .RST(rst), .Q(
        start_reg[912]) );
  DFF \start_reg_reg[913]  ( .D(start_in[912]), .CLK(clk), .RST(rst), .Q(
        start_reg[913]) );
  DFF \start_reg_reg[914]  ( .D(start_in[913]), .CLK(clk), .RST(rst), .Q(
        start_reg[914]) );
  DFF \start_reg_reg[915]  ( .D(start_in[914]), .CLK(clk), .RST(rst), .Q(
        start_reg[915]) );
  DFF \start_reg_reg[916]  ( .D(start_in[915]), .CLK(clk), .RST(rst), .Q(
        start_reg[916]) );
  DFF \start_reg_reg[917]  ( .D(start_in[916]), .CLK(clk), .RST(rst), .Q(
        start_reg[917]) );
  DFF \start_reg_reg[918]  ( .D(start_in[917]), .CLK(clk), .RST(rst), .Q(
        start_reg[918]) );
  DFF \start_reg_reg[919]  ( .D(start_in[918]), .CLK(clk), .RST(rst), .Q(
        start_reg[919]) );
  DFF \start_reg_reg[920]  ( .D(start_in[919]), .CLK(clk), .RST(rst), .Q(
        start_reg[920]) );
  DFF \start_reg_reg[921]  ( .D(start_in[920]), .CLK(clk), .RST(rst), .Q(
        start_reg[921]) );
  DFF \start_reg_reg[922]  ( .D(start_in[921]), .CLK(clk), .RST(rst), .Q(
        start_reg[922]) );
  DFF \start_reg_reg[923]  ( .D(start_in[922]), .CLK(clk), .RST(rst), .Q(
        start_reg[923]) );
  DFF \start_reg_reg[924]  ( .D(start_in[923]), .CLK(clk), .RST(rst), .Q(
        start_reg[924]) );
  DFF \start_reg_reg[925]  ( .D(start_in[924]), .CLK(clk), .RST(rst), .Q(
        start_reg[925]) );
  DFF \start_reg_reg[926]  ( .D(start_in[925]), .CLK(clk), .RST(rst), .Q(
        start_reg[926]) );
  DFF \start_reg_reg[927]  ( .D(start_in[926]), .CLK(clk), .RST(rst), .Q(
        start_reg[927]) );
  DFF \start_reg_reg[928]  ( .D(start_in[927]), .CLK(clk), .RST(rst), .Q(
        start_reg[928]) );
  DFF \start_reg_reg[929]  ( .D(start_in[928]), .CLK(clk), .RST(rst), .Q(
        start_reg[929]) );
  DFF \start_reg_reg[930]  ( .D(start_in[929]), .CLK(clk), .RST(rst), .Q(
        start_reg[930]) );
  DFF \start_reg_reg[931]  ( .D(start_in[930]), .CLK(clk), .RST(rst), .Q(
        start_reg[931]) );
  DFF \start_reg_reg[932]  ( .D(start_in[931]), .CLK(clk), .RST(rst), .Q(
        start_reg[932]) );
  DFF \start_reg_reg[933]  ( .D(start_in[932]), .CLK(clk), .RST(rst), .Q(
        start_reg[933]) );
  DFF \start_reg_reg[934]  ( .D(start_in[933]), .CLK(clk), .RST(rst), .Q(
        start_reg[934]) );
  DFF \start_reg_reg[935]  ( .D(start_in[934]), .CLK(clk), .RST(rst), .Q(
        start_reg[935]) );
  DFF \start_reg_reg[936]  ( .D(start_in[935]), .CLK(clk), .RST(rst), .Q(
        start_reg[936]) );
  DFF \start_reg_reg[937]  ( .D(start_in[936]), .CLK(clk), .RST(rst), .Q(
        start_reg[937]) );
  DFF \start_reg_reg[938]  ( .D(start_in[937]), .CLK(clk), .RST(rst), .Q(
        start_reg[938]) );
  DFF \start_reg_reg[939]  ( .D(start_in[938]), .CLK(clk), .RST(rst), .Q(
        start_reg[939]) );
  DFF \start_reg_reg[940]  ( .D(start_in[939]), .CLK(clk), .RST(rst), .Q(
        start_reg[940]) );
  DFF \start_reg_reg[941]  ( .D(start_in[940]), .CLK(clk), .RST(rst), .Q(
        start_reg[941]) );
  DFF \start_reg_reg[942]  ( .D(start_in[941]), .CLK(clk), .RST(rst), .Q(
        start_reg[942]) );
  DFF \start_reg_reg[943]  ( .D(start_in[942]), .CLK(clk), .RST(rst), .Q(
        start_reg[943]) );
  DFF \start_reg_reg[944]  ( .D(start_in[943]), .CLK(clk), .RST(rst), .Q(
        start_reg[944]) );
  DFF \start_reg_reg[945]  ( .D(start_in[944]), .CLK(clk), .RST(rst), .Q(
        start_reg[945]) );
  DFF \start_reg_reg[946]  ( .D(start_in[945]), .CLK(clk), .RST(rst), .Q(
        start_reg[946]) );
  DFF \start_reg_reg[947]  ( .D(start_in[946]), .CLK(clk), .RST(rst), .Q(
        start_reg[947]) );
  DFF \start_reg_reg[948]  ( .D(start_in[947]), .CLK(clk), .RST(rst), .Q(
        start_reg[948]) );
  DFF \start_reg_reg[949]  ( .D(start_in[948]), .CLK(clk), .RST(rst), .Q(
        start_reg[949]) );
  DFF \start_reg_reg[950]  ( .D(start_in[949]), .CLK(clk), .RST(rst), .Q(
        start_reg[950]) );
  DFF \start_reg_reg[951]  ( .D(start_in[950]), .CLK(clk), .RST(rst), .Q(
        start_reg[951]) );
  DFF \start_reg_reg[952]  ( .D(start_in[951]), .CLK(clk), .RST(rst), .Q(
        start_reg[952]) );
  DFF \start_reg_reg[953]  ( .D(start_in[952]), .CLK(clk), .RST(rst), .Q(
        start_reg[953]) );
  DFF \start_reg_reg[954]  ( .D(start_in[953]), .CLK(clk), .RST(rst), .Q(
        start_reg[954]) );
  DFF \start_reg_reg[955]  ( .D(start_in[954]), .CLK(clk), .RST(rst), .Q(
        start_reg[955]) );
  DFF \start_reg_reg[956]  ( .D(start_in[955]), .CLK(clk), .RST(rst), .Q(
        start_reg[956]) );
  DFF \start_reg_reg[957]  ( .D(start_in[956]), .CLK(clk), .RST(rst), .Q(
        start_reg[957]) );
  DFF \start_reg_reg[958]  ( .D(start_in[957]), .CLK(clk), .RST(rst), .Q(
        start_reg[958]) );
  DFF \start_reg_reg[959]  ( .D(start_in[958]), .CLK(clk), .RST(rst), .Q(
        start_reg[959]) );
  DFF \start_reg_reg[960]  ( .D(start_in[959]), .CLK(clk), .RST(rst), .Q(
        start_reg[960]) );
  DFF \start_reg_reg[961]  ( .D(start_in[960]), .CLK(clk), .RST(rst), .Q(
        start_reg[961]) );
  DFF \start_reg_reg[962]  ( .D(start_in[961]), .CLK(clk), .RST(rst), .Q(
        start_reg[962]) );
  DFF \start_reg_reg[963]  ( .D(start_in[962]), .CLK(clk), .RST(rst), .Q(
        start_reg[963]) );
  DFF \start_reg_reg[964]  ( .D(start_in[963]), .CLK(clk), .RST(rst), .Q(
        start_reg[964]) );
  DFF \start_reg_reg[965]  ( .D(start_in[964]), .CLK(clk), .RST(rst), .Q(
        start_reg[965]) );
  DFF \start_reg_reg[966]  ( .D(start_in[965]), .CLK(clk), .RST(rst), .Q(
        start_reg[966]) );
  DFF \start_reg_reg[967]  ( .D(start_in[966]), .CLK(clk), .RST(rst), .Q(
        start_reg[967]) );
  DFF \start_reg_reg[968]  ( .D(start_in[967]), .CLK(clk), .RST(rst), .Q(
        start_reg[968]) );
  DFF \start_reg_reg[969]  ( .D(start_in[968]), .CLK(clk), .RST(rst), .Q(
        start_reg[969]) );
  DFF \start_reg_reg[970]  ( .D(start_in[969]), .CLK(clk), .RST(rst), .Q(
        start_reg[970]) );
  DFF \start_reg_reg[971]  ( .D(start_in[970]), .CLK(clk), .RST(rst), .Q(
        start_reg[971]) );
  DFF \start_reg_reg[972]  ( .D(start_in[971]), .CLK(clk), .RST(rst), .Q(
        start_reg[972]) );
  DFF \start_reg_reg[973]  ( .D(start_in[972]), .CLK(clk), .RST(rst), .Q(
        start_reg[973]) );
  DFF \start_reg_reg[974]  ( .D(start_in[973]), .CLK(clk), .RST(rst), .Q(
        start_reg[974]) );
  DFF \start_reg_reg[975]  ( .D(start_in[974]), .CLK(clk), .RST(rst), .Q(
        start_reg[975]) );
  DFF \start_reg_reg[976]  ( .D(start_in[975]), .CLK(clk), .RST(rst), .Q(
        start_reg[976]) );
  DFF \start_reg_reg[977]  ( .D(start_in[976]), .CLK(clk), .RST(rst), .Q(
        start_reg[977]) );
  DFF \start_reg_reg[978]  ( .D(start_in[977]), .CLK(clk), .RST(rst), .Q(
        start_reg[978]) );
  DFF \start_reg_reg[979]  ( .D(start_in[978]), .CLK(clk), .RST(rst), .Q(
        start_reg[979]) );
  DFF \start_reg_reg[980]  ( .D(start_in[979]), .CLK(clk), .RST(rst), .Q(
        start_reg[980]) );
  DFF \start_reg_reg[981]  ( .D(start_in[980]), .CLK(clk), .RST(rst), .Q(
        start_reg[981]) );
  DFF \start_reg_reg[982]  ( .D(start_in[981]), .CLK(clk), .RST(rst), .Q(
        start_reg[982]) );
  DFF \start_reg_reg[983]  ( .D(start_in[982]), .CLK(clk), .RST(rst), .Q(
        start_reg[983]) );
  DFF \start_reg_reg[984]  ( .D(start_in[983]), .CLK(clk), .RST(rst), .Q(
        start_reg[984]) );
  DFF \start_reg_reg[985]  ( .D(start_in[984]), .CLK(clk), .RST(rst), .Q(
        start_reg[985]) );
  DFF \start_reg_reg[986]  ( .D(start_in[985]), .CLK(clk), .RST(rst), .Q(
        start_reg[986]) );
  DFF \start_reg_reg[987]  ( .D(start_in[986]), .CLK(clk), .RST(rst), .Q(
        start_reg[987]) );
  DFF \start_reg_reg[988]  ( .D(start_in[987]), .CLK(clk), .RST(rst), .Q(
        start_reg[988]) );
  DFF \start_reg_reg[989]  ( .D(start_in[988]), .CLK(clk), .RST(rst), .Q(
        start_reg[989]) );
  DFF \start_reg_reg[990]  ( .D(start_in[989]), .CLK(clk), .RST(rst), .Q(
        start_reg[990]) );
  DFF \start_reg_reg[991]  ( .D(start_in[990]), .CLK(clk), .RST(rst), .Q(
        start_reg[991]) );
  DFF \start_reg_reg[992]  ( .D(start_in[991]), .CLK(clk), .RST(rst), .Q(
        start_reg[992]) );
  DFF \start_reg_reg[993]  ( .D(start_in[992]), .CLK(clk), .RST(rst), .Q(
        start_reg[993]) );
  DFF \start_reg_reg[994]  ( .D(start_in[993]), .CLK(clk), .RST(rst), .Q(
        start_reg[994]) );
  DFF \start_reg_reg[995]  ( .D(start_in[994]), .CLK(clk), .RST(rst), .Q(
        start_reg[995]) );
  DFF \start_reg_reg[996]  ( .D(start_in[995]), .CLK(clk), .RST(rst), .Q(
        start_reg[996]) );
  DFF \start_reg_reg[997]  ( .D(start_in[996]), .CLK(clk), .RST(rst), .Q(
        start_reg[997]) );
  DFF \start_reg_reg[998]  ( .D(start_in[997]), .CLK(clk), .RST(rst), .Q(
        start_reg[998]) );
  DFF \start_reg_reg[999]  ( .D(start_in[998]), .CLK(clk), .RST(rst), .Q(
        start_reg[999]) );
  DFF \start_reg_reg[1000]  ( .D(start_in[999]), .CLK(clk), .RST(rst), .Q(
        start_reg[1000]) );
  DFF \start_reg_reg[1001]  ( .D(start_in[1000]), .CLK(clk), .RST(rst), .Q(
        start_reg[1001]) );
  DFF \start_reg_reg[1002]  ( .D(start_in[1001]), .CLK(clk), .RST(rst), .Q(
        start_reg[1002]) );
  DFF \start_reg_reg[1003]  ( .D(start_in[1002]), .CLK(clk), .RST(rst), .Q(
        start_reg[1003]) );
  DFF \start_reg_reg[1004]  ( .D(start_in[1003]), .CLK(clk), .RST(rst), .Q(
        start_reg[1004]) );
  DFF \start_reg_reg[1005]  ( .D(start_in[1004]), .CLK(clk), .RST(rst), .Q(
        start_reg[1005]) );
  DFF \start_reg_reg[1006]  ( .D(start_in[1005]), .CLK(clk), .RST(rst), .Q(
        start_reg[1006]) );
  DFF \start_reg_reg[1007]  ( .D(start_in[1006]), .CLK(clk), .RST(rst), .Q(
        start_reg[1007]) );
  DFF \start_reg_reg[1008]  ( .D(start_in[1007]), .CLK(clk), .RST(rst), .Q(
        start_reg[1008]) );
  DFF \start_reg_reg[1009]  ( .D(start_in[1008]), .CLK(clk), .RST(rst), .Q(
        start_reg[1009]) );
  DFF \start_reg_reg[1010]  ( .D(start_in[1009]), .CLK(clk), .RST(rst), .Q(
        start_reg[1010]) );
  DFF \start_reg_reg[1011]  ( .D(start_in[1010]), .CLK(clk), .RST(rst), .Q(
        start_reg[1011]) );
  DFF \start_reg_reg[1012]  ( .D(start_in[1011]), .CLK(clk), .RST(rst), .Q(
        start_reg[1012]) );
  DFF \start_reg_reg[1013]  ( .D(start_in[1012]), .CLK(clk), .RST(rst), .Q(
        start_reg[1013]) );
  DFF \start_reg_reg[1014]  ( .D(start_in[1013]), .CLK(clk), .RST(rst), .Q(
        start_reg[1014]) );
  DFF \start_reg_reg[1015]  ( .D(start_in[1014]), .CLK(clk), .RST(rst), .Q(
        start_reg[1015]) );
  DFF \start_reg_reg[1016]  ( .D(start_in[1015]), .CLK(clk), .RST(rst), .Q(
        start_reg[1016]) );
  DFF \start_reg_reg[1017]  ( .D(start_in[1016]), .CLK(clk), .RST(rst), .Q(
        start_reg[1017]) );
  DFF \start_reg_reg[1018]  ( .D(start_in[1017]), .CLK(clk), .RST(rst), .Q(
        start_reg[1018]) );
  DFF \start_reg_reg[1019]  ( .D(start_in[1018]), .CLK(clk), .RST(rst), .Q(
        start_reg[1019]) );
  DFF \start_reg_reg[1020]  ( .D(start_in[1019]), .CLK(clk), .RST(rst), .Q(
        start_reg[1020]) );
  DFF \start_reg_reg[1021]  ( .D(start_in[1020]), .CLK(clk), .RST(rst), .Q(
        start_reg[1021]) );
  DFF \start_reg_reg[1022]  ( .D(start_in[1021]), .CLK(clk), .RST(rst), .Q(
        start_reg[1022]) );
  DFF \start_reg_reg[1023]  ( .D(start_in[1022]), .CLK(clk), .RST(rst), .Q(
        start_reg[1023]) );
  DFF mul_pow_reg ( .D(n15378), .CLK(clk), .RST(rst), .Q(mul_pow) );
  DFF \ereg_reg[0]  ( .D(n15377), .CLK(clk), .RST(rst), .Q(ereg[0]) );
  DFF \ereg_reg[1]  ( .D(n15376), .CLK(clk), .RST(rst), .Q(ereg[1]) );
  DFF \ereg_reg[2]  ( .D(n15375), .CLK(clk), .RST(rst), .Q(ereg[2]) );
  DFF \ereg_reg[3]  ( .D(n15374), .CLK(clk), .RST(rst), .Q(ereg[3]) );
  DFF \ereg_reg[4]  ( .D(n15373), .CLK(clk), .RST(rst), .Q(ereg[4]) );
  DFF \ereg_reg[5]  ( .D(n15372), .CLK(clk), .RST(rst), .Q(ereg[5]) );
  DFF \ereg_reg[6]  ( .D(n15371), .CLK(clk), .RST(rst), .Q(ereg[6]) );
  DFF \ereg_reg[7]  ( .D(n15370), .CLK(clk), .RST(rst), .Q(ereg[7]) );
  DFF \ereg_reg[8]  ( .D(n15369), .CLK(clk), .RST(rst), .Q(ereg[8]) );
  DFF \ereg_reg[9]  ( .D(n15368), .CLK(clk), .RST(rst), .Q(ereg[9]) );
  DFF \ereg_reg[10]  ( .D(n15367), .CLK(clk), .RST(rst), .Q(ereg[10]) );
  DFF \ereg_reg[11]  ( .D(n15366), .CLK(clk), .RST(rst), .Q(ereg[11]) );
  DFF \ereg_reg[12]  ( .D(n15365), .CLK(clk), .RST(rst), .Q(ereg[12]) );
  DFF \ereg_reg[13]  ( .D(n15364), .CLK(clk), .RST(rst), .Q(ereg[13]) );
  DFF \ereg_reg[14]  ( .D(n15363), .CLK(clk), .RST(rst), .Q(ereg[14]) );
  DFF \ereg_reg[15]  ( .D(n15362), .CLK(clk), .RST(rst), .Q(ereg[15]) );
  DFF \ereg_reg[16]  ( .D(n15361), .CLK(clk), .RST(rst), .Q(ereg[16]) );
  DFF \ereg_reg[17]  ( .D(n15360), .CLK(clk), .RST(rst), .Q(ereg[17]) );
  DFF \ereg_reg[18]  ( .D(n15359), .CLK(clk), .RST(rst), .Q(ereg[18]) );
  DFF \ereg_reg[19]  ( .D(n15358), .CLK(clk), .RST(rst), .Q(ereg[19]) );
  DFF \ereg_reg[20]  ( .D(n15357), .CLK(clk), .RST(rst), .Q(ereg[20]) );
  DFF \ereg_reg[21]  ( .D(n15356), .CLK(clk), .RST(rst), .Q(ereg[21]) );
  DFF \ereg_reg[22]  ( .D(n15355), .CLK(clk), .RST(rst), .Q(ereg[22]) );
  DFF \ereg_reg[23]  ( .D(n15354), .CLK(clk), .RST(rst), .Q(ereg[23]) );
  DFF \ereg_reg[24]  ( .D(n15353), .CLK(clk), .RST(rst), .Q(ereg[24]) );
  DFF \ereg_reg[25]  ( .D(n15352), .CLK(clk), .RST(rst), .Q(ereg[25]) );
  DFF \ereg_reg[26]  ( .D(n15351), .CLK(clk), .RST(rst), .Q(ereg[26]) );
  DFF \ereg_reg[27]  ( .D(n15350), .CLK(clk), .RST(rst), .Q(ereg[27]) );
  DFF \ereg_reg[28]  ( .D(n15349), .CLK(clk), .RST(rst), .Q(ereg[28]) );
  DFF \ereg_reg[29]  ( .D(n15348), .CLK(clk), .RST(rst), .Q(ereg[29]) );
  DFF \ereg_reg[30]  ( .D(n15347), .CLK(clk), .RST(rst), .Q(ereg[30]) );
  DFF \ereg_reg[31]  ( .D(n15346), .CLK(clk), .RST(rst), .Q(ereg[31]) );
  DFF \ereg_reg[32]  ( .D(n15345), .CLK(clk), .RST(rst), .Q(ereg[32]) );
  DFF \ereg_reg[33]  ( .D(n15344), .CLK(clk), .RST(rst), .Q(ereg[33]) );
  DFF \ereg_reg[34]  ( .D(n15343), .CLK(clk), .RST(rst), .Q(ereg[34]) );
  DFF \ereg_reg[35]  ( .D(n15342), .CLK(clk), .RST(rst), .Q(ereg[35]) );
  DFF \ereg_reg[36]  ( .D(n15341), .CLK(clk), .RST(rst), .Q(ereg[36]) );
  DFF \ereg_reg[37]  ( .D(n15340), .CLK(clk), .RST(rst), .Q(ereg[37]) );
  DFF \ereg_reg[38]  ( .D(n15339), .CLK(clk), .RST(rst), .Q(ereg[38]) );
  DFF \ereg_reg[39]  ( .D(n15338), .CLK(clk), .RST(rst), .Q(ereg[39]) );
  DFF \ereg_reg[40]  ( .D(n15337), .CLK(clk), .RST(rst), .Q(ereg[40]) );
  DFF \ereg_reg[41]  ( .D(n15336), .CLK(clk), .RST(rst), .Q(ereg[41]) );
  DFF \ereg_reg[42]  ( .D(n15335), .CLK(clk), .RST(rst), .Q(ereg[42]) );
  DFF \ereg_reg[43]  ( .D(n15334), .CLK(clk), .RST(rst), .Q(ereg[43]) );
  DFF \ereg_reg[44]  ( .D(n15333), .CLK(clk), .RST(rst), .Q(ereg[44]) );
  DFF \ereg_reg[45]  ( .D(n15332), .CLK(clk), .RST(rst), .Q(ereg[45]) );
  DFF \ereg_reg[46]  ( .D(n15331), .CLK(clk), .RST(rst), .Q(ereg[46]) );
  DFF \ereg_reg[47]  ( .D(n15330), .CLK(clk), .RST(rst), .Q(ereg[47]) );
  DFF \ereg_reg[48]  ( .D(n15329), .CLK(clk), .RST(rst), .Q(ereg[48]) );
  DFF \ereg_reg[49]  ( .D(n15328), .CLK(clk), .RST(rst), .Q(ereg[49]) );
  DFF \ereg_reg[50]  ( .D(n15327), .CLK(clk), .RST(rst), .Q(ereg[50]) );
  DFF \ereg_reg[51]  ( .D(n15326), .CLK(clk), .RST(rst), .Q(ereg[51]) );
  DFF \ereg_reg[52]  ( .D(n15325), .CLK(clk), .RST(rst), .Q(ereg[52]) );
  DFF \ereg_reg[53]  ( .D(n15324), .CLK(clk), .RST(rst), .Q(ereg[53]) );
  DFF \ereg_reg[54]  ( .D(n15323), .CLK(clk), .RST(rst), .Q(ereg[54]) );
  DFF \ereg_reg[55]  ( .D(n15322), .CLK(clk), .RST(rst), .Q(ereg[55]) );
  DFF \ereg_reg[56]  ( .D(n15321), .CLK(clk), .RST(rst), .Q(ereg[56]) );
  DFF \ereg_reg[57]  ( .D(n15320), .CLK(clk), .RST(rst), .Q(ereg[57]) );
  DFF \ereg_reg[58]  ( .D(n15319), .CLK(clk), .RST(rst), .Q(ereg[58]) );
  DFF \ereg_reg[59]  ( .D(n15318), .CLK(clk), .RST(rst), .Q(ereg[59]) );
  DFF \ereg_reg[60]  ( .D(n15317), .CLK(clk), .RST(rst), .Q(ereg[60]) );
  DFF \ereg_reg[61]  ( .D(n15316), .CLK(clk), .RST(rst), .Q(ereg[61]) );
  DFF \ereg_reg[62]  ( .D(n15315), .CLK(clk), .RST(rst), .Q(ereg[62]) );
  DFF \ereg_reg[63]  ( .D(n15314), .CLK(clk), .RST(rst), .Q(ereg[63]) );
  DFF \ereg_reg[64]  ( .D(n15313), .CLK(clk), .RST(rst), .Q(ereg[64]) );
  DFF \ereg_reg[65]  ( .D(n15312), .CLK(clk), .RST(rst), .Q(ereg[65]) );
  DFF \ereg_reg[66]  ( .D(n15311), .CLK(clk), .RST(rst), .Q(ereg[66]) );
  DFF \ereg_reg[67]  ( .D(n15310), .CLK(clk), .RST(rst), .Q(ereg[67]) );
  DFF \ereg_reg[68]  ( .D(n15309), .CLK(clk), .RST(rst), .Q(ereg[68]) );
  DFF \ereg_reg[69]  ( .D(n15308), .CLK(clk), .RST(rst), .Q(ereg[69]) );
  DFF \ereg_reg[70]  ( .D(n15307), .CLK(clk), .RST(rst), .Q(ereg[70]) );
  DFF \ereg_reg[71]  ( .D(n15306), .CLK(clk), .RST(rst), .Q(ereg[71]) );
  DFF \ereg_reg[72]  ( .D(n15305), .CLK(clk), .RST(rst), .Q(ereg[72]) );
  DFF \ereg_reg[73]  ( .D(n15304), .CLK(clk), .RST(rst), .Q(ereg[73]) );
  DFF \ereg_reg[74]  ( .D(n15303), .CLK(clk), .RST(rst), .Q(ereg[74]) );
  DFF \ereg_reg[75]  ( .D(n15302), .CLK(clk), .RST(rst), .Q(ereg[75]) );
  DFF \ereg_reg[76]  ( .D(n15301), .CLK(clk), .RST(rst), .Q(ereg[76]) );
  DFF \ereg_reg[77]  ( .D(n15300), .CLK(clk), .RST(rst), .Q(ereg[77]) );
  DFF \ereg_reg[78]  ( .D(n15299), .CLK(clk), .RST(rst), .Q(ereg[78]) );
  DFF \ereg_reg[79]  ( .D(n15298), .CLK(clk), .RST(rst), .Q(ereg[79]) );
  DFF \ereg_reg[80]  ( .D(n15297), .CLK(clk), .RST(rst), .Q(ereg[80]) );
  DFF \ereg_reg[81]  ( .D(n15296), .CLK(clk), .RST(rst), .Q(ereg[81]) );
  DFF \ereg_reg[82]  ( .D(n15295), .CLK(clk), .RST(rst), .Q(ereg[82]) );
  DFF \ereg_reg[83]  ( .D(n15294), .CLK(clk), .RST(rst), .Q(ereg[83]) );
  DFF \ereg_reg[84]  ( .D(n15293), .CLK(clk), .RST(rst), .Q(ereg[84]) );
  DFF \ereg_reg[85]  ( .D(n15292), .CLK(clk), .RST(rst), .Q(ereg[85]) );
  DFF \ereg_reg[86]  ( .D(n15291), .CLK(clk), .RST(rst), .Q(ereg[86]) );
  DFF \ereg_reg[87]  ( .D(n15290), .CLK(clk), .RST(rst), .Q(ereg[87]) );
  DFF \ereg_reg[88]  ( .D(n15289), .CLK(clk), .RST(rst), .Q(ereg[88]) );
  DFF \ereg_reg[89]  ( .D(n15288), .CLK(clk), .RST(rst), .Q(ereg[89]) );
  DFF \ereg_reg[90]  ( .D(n15287), .CLK(clk), .RST(rst), .Q(ereg[90]) );
  DFF \ereg_reg[91]  ( .D(n15286), .CLK(clk), .RST(rst), .Q(ereg[91]) );
  DFF \ereg_reg[92]  ( .D(n15285), .CLK(clk), .RST(rst), .Q(ereg[92]) );
  DFF \ereg_reg[93]  ( .D(n15284), .CLK(clk), .RST(rst), .Q(ereg[93]) );
  DFF \ereg_reg[94]  ( .D(n15283), .CLK(clk), .RST(rst), .Q(ereg[94]) );
  DFF \ereg_reg[95]  ( .D(n15282), .CLK(clk), .RST(rst), .Q(ereg[95]) );
  DFF \ereg_reg[96]  ( .D(n15281), .CLK(clk), .RST(rst), .Q(ereg[96]) );
  DFF \ereg_reg[97]  ( .D(n15280), .CLK(clk), .RST(rst), .Q(ereg[97]) );
  DFF \ereg_reg[98]  ( .D(n15279), .CLK(clk), .RST(rst), .Q(ereg[98]) );
  DFF \ereg_reg[99]  ( .D(n15278), .CLK(clk), .RST(rst), .Q(ereg[99]) );
  DFF \ereg_reg[100]  ( .D(n15277), .CLK(clk), .RST(rst), .Q(ereg[100]) );
  DFF \ereg_reg[101]  ( .D(n15276), .CLK(clk), .RST(rst), .Q(ereg[101]) );
  DFF \ereg_reg[102]  ( .D(n15275), .CLK(clk), .RST(rst), .Q(ereg[102]) );
  DFF \ereg_reg[103]  ( .D(n15274), .CLK(clk), .RST(rst), .Q(ereg[103]) );
  DFF \ereg_reg[104]  ( .D(n15273), .CLK(clk), .RST(rst), .Q(ereg[104]) );
  DFF \ereg_reg[105]  ( .D(n15272), .CLK(clk), .RST(rst), .Q(ereg[105]) );
  DFF \ereg_reg[106]  ( .D(n15271), .CLK(clk), .RST(rst), .Q(ereg[106]) );
  DFF \ereg_reg[107]  ( .D(n15270), .CLK(clk), .RST(rst), .Q(ereg[107]) );
  DFF \ereg_reg[108]  ( .D(n15269), .CLK(clk), .RST(rst), .Q(ereg[108]) );
  DFF \ereg_reg[109]  ( .D(n15268), .CLK(clk), .RST(rst), .Q(ereg[109]) );
  DFF \ereg_reg[110]  ( .D(n15267), .CLK(clk), .RST(rst), .Q(ereg[110]) );
  DFF \ereg_reg[111]  ( .D(n15266), .CLK(clk), .RST(rst), .Q(ereg[111]) );
  DFF \ereg_reg[112]  ( .D(n15265), .CLK(clk), .RST(rst), .Q(ereg[112]) );
  DFF \ereg_reg[113]  ( .D(n15264), .CLK(clk), .RST(rst), .Q(ereg[113]) );
  DFF \ereg_reg[114]  ( .D(n15263), .CLK(clk), .RST(rst), .Q(ereg[114]) );
  DFF \ereg_reg[115]  ( .D(n15262), .CLK(clk), .RST(rst), .Q(ereg[115]) );
  DFF \ereg_reg[116]  ( .D(n15261), .CLK(clk), .RST(rst), .Q(ereg[116]) );
  DFF \ereg_reg[117]  ( .D(n15260), .CLK(clk), .RST(rst), .Q(ereg[117]) );
  DFF \ereg_reg[118]  ( .D(n15259), .CLK(clk), .RST(rst), .Q(ereg[118]) );
  DFF \ereg_reg[119]  ( .D(n15258), .CLK(clk), .RST(rst), .Q(ereg[119]) );
  DFF \ereg_reg[120]  ( .D(n15257), .CLK(clk), .RST(rst), .Q(ereg[120]) );
  DFF \ereg_reg[121]  ( .D(n15256), .CLK(clk), .RST(rst), .Q(ereg[121]) );
  DFF \ereg_reg[122]  ( .D(n15255), .CLK(clk), .RST(rst), .Q(ereg[122]) );
  DFF \ereg_reg[123]  ( .D(n15254), .CLK(clk), .RST(rst), .Q(ereg[123]) );
  DFF \ereg_reg[124]  ( .D(n15253), .CLK(clk), .RST(rst), .Q(ereg[124]) );
  DFF \ereg_reg[125]  ( .D(n15252), .CLK(clk), .RST(rst), .Q(ereg[125]) );
  DFF \ereg_reg[126]  ( .D(n15251), .CLK(clk), .RST(rst), .Q(ereg[126]) );
  DFF \ereg_reg[127]  ( .D(n15250), .CLK(clk), .RST(rst), .Q(ereg[127]) );
  DFF \ereg_reg[128]  ( .D(n15249), .CLK(clk), .RST(rst), .Q(ereg[128]) );
  DFF \ereg_reg[129]  ( .D(n15248), .CLK(clk), .RST(rst), .Q(ereg[129]) );
  DFF \ereg_reg[130]  ( .D(n15247), .CLK(clk), .RST(rst), .Q(ereg[130]) );
  DFF \ereg_reg[131]  ( .D(n15246), .CLK(clk), .RST(rst), .Q(ereg[131]) );
  DFF \ereg_reg[132]  ( .D(n15245), .CLK(clk), .RST(rst), .Q(ereg[132]) );
  DFF \ereg_reg[133]  ( .D(n15244), .CLK(clk), .RST(rst), .Q(ereg[133]) );
  DFF \ereg_reg[134]  ( .D(n15243), .CLK(clk), .RST(rst), .Q(ereg[134]) );
  DFF \ereg_reg[135]  ( .D(n15242), .CLK(clk), .RST(rst), .Q(ereg[135]) );
  DFF \ereg_reg[136]  ( .D(n15241), .CLK(clk), .RST(rst), .Q(ereg[136]) );
  DFF \ereg_reg[137]  ( .D(n15240), .CLK(clk), .RST(rst), .Q(ereg[137]) );
  DFF \ereg_reg[138]  ( .D(n15239), .CLK(clk), .RST(rst), .Q(ereg[138]) );
  DFF \ereg_reg[139]  ( .D(n15238), .CLK(clk), .RST(rst), .Q(ereg[139]) );
  DFF \ereg_reg[140]  ( .D(n15237), .CLK(clk), .RST(rst), .Q(ereg[140]) );
  DFF \ereg_reg[141]  ( .D(n15236), .CLK(clk), .RST(rst), .Q(ereg[141]) );
  DFF \ereg_reg[142]  ( .D(n15235), .CLK(clk), .RST(rst), .Q(ereg[142]) );
  DFF \ereg_reg[143]  ( .D(n15234), .CLK(clk), .RST(rst), .Q(ereg[143]) );
  DFF \ereg_reg[144]  ( .D(n15233), .CLK(clk), .RST(rst), .Q(ereg[144]) );
  DFF \ereg_reg[145]  ( .D(n15232), .CLK(clk), .RST(rst), .Q(ereg[145]) );
  DFF \ereg_reg[146]  ( .D(n15231), .CLK(clk), .RST(rst), .Q(ereg[146]) );
  DFF \ereg_reg[147]  ( .D(n15230), .CLK(clk), .RST(rst), .Q(ereg[147]) );
  DFF \ereg_reg[148]  ( .D(n15229), .CLK(clk), .RST(rst), .Q(ereg[148]) );
  DFF \ereg_reg[149]  ( .D(n15228), .CLK(clk), .RST(rst), .Q(ereg[149]) );
  DFF \ereg_reg[150]  ( .D(n15227), .CLK(clk), .RST(rst), .Q(ereg[150]) );
  DFF \ereg_reg[151]  ( .D(n15226), .CLK(clk), .RST(rst), .Q(ereg[151]) );
  DFF \ereg_reg[152]  ( .D(n15225), .CLK(clk), .RST(rst), .Q(ereg[152]) );
  DFF \ereg_reg[153]  ( .D(n15224), .CLK(clk), .RST(rst), .Q(ereg[153]) );
  DFF \ereg_reg[154]  ( .D(n15223), .CLK(clk), .RST(rst), .Q(ereg[154]) );
  DFF \ereg_reg[155]  ( .D(n15222), .CLK(clk), .RST(rst), .Q(ereg[155]) );
  DFF \ereg_reg[156]  ( .D(n15221), .CLK(clk), .RST(rst), .Q(ereg[156]) );
  DFF \ereg_reg[157]  ( .D(n15220), .CLK(clk), .RST(rst), .Q(ereg[157]) );
  DFF \ereg_reg[158]  ( .D(n15219), .CLK(clk), .RST(rst), .Q(ereg[158]) );
  DFF \ereg_reg[159]  ( .D(n15218), .CLK(clk), .RST(rst), .Q(ereg[159]) );
  DFF \ereg_reg[160]  ( .D(n15217), .CLK(clk), .RST(rst), .Q(ereg[160]) );
  DFF \ereg_reg[161]  ( .D(n15216), .CLK(clk), .RST(rst), .Q(ereg[161]) );
  DFF \ereg_reg[162]  ( .D(n15215), .CLK(clk), .RST(rst), .Q(ereg[162]) );
  DFF \ereg_reg[163]  ( .D(n15214), .CLK(clk), .RST(rst), .Q(ereg[163]) );
  DFF \ereg_reg[164]  ( .D(n15213), .CLK(clk), .RST(rst), .Q(ereg[164]) );
  DFF \ereg_reg[165]  ( .D(n15212), .CLK(clk), .RST(rst), .Q(ereg[165]) );
  DFF \ereg_reg[166]  ( .D(n15211), .CLK(clk), .RST(rst), .Q(ereg[166]) );
  DFF \ereg_reg[167]  ( .D(n15210), .CLK(clk), .RST(rst), .Q(ereg[167]) );
  DFF \ereg_reg[168]  ( .D(n15209), .CLK(clk), .RST(rst), .Q(ereg[168]) );
  DFF \ereg_reg[169]  ( .D(n15208), .CLK(clk), .RST(rst), .Q(ereg[169]) );
  DFF \ereg_reg[170]  ( .D(n15207), .CLK(clk), .RST(rst), .Q(ereg[170]) );
  DFF \ereg_reg[171]  ( .D(n15206), .CLK(clk), .RST(rst), .Q(ereg[171]) );
  DFF \ereg_reg[172]  ( .D(n15205), .CLK(clk), .RST(rst), .Q(ereg[172]) );
  DFF \ereg_reg[173]  ( .D(n15204), .CLK(clk), .RST(rst), .Q(ereg[173]) );
  DFF \ereg_reg[174]  ( .D(n15203), .CLK(clk), .RST(rst), .Q(ereg[174]) );
  DFF \ereg_reg[175]  ( .D(n15202), .CLK(clk), .RST(rst), .Q(ereg[175]) );
  DFF \ereg_reg[176]  ( .D(n15201), .CLK(clk), .RST(rst), .Q(ereg[176]) );
  DFF \ereg_reg[177]  ( .D(n15200), .CLK(clk), .RST(rst), .Q(ereg[177]) );
  DFF \ereg_reg[178]  ( .D(n15199), .CLK(clk), .RST(rst), .Q(ereg[178]) );
  DFF \ereg_reg[179]  ( .D(n15198), .CLK(clk), .RST(rst), .Q(ereg[179]) );
  DFF \ereg_reg[180]  ( .D(n15197), .CLK(clk), .RST(rst), .Q(ereg[180]) );
  DFF \ereg_reg[181]  ( .D(n15196), .CLK(clk), .RST(rst), .Q(ereg[181]) );
  DFF \ereg_reg[182]  ( .D(n15195), .CLK(clk), .RST(rst), .Q(ereg[182]) );
  DFF \ereg_reg[183]  ( .D(n15194), .CLK(clk), .RST(rst), .Q(ereg[183]) );
  DFF \ereg_reg[184]  ( .D(n15193), .CLK(clk), .RST(rst), .Q(ereg[184]) );
  DFF \ereg_reg[185]  ( .D(n15192), .CLK(clk), .RST(rst), .Q(ereg[185]) );
  DFF \ereg_reg[186]  ( .D(n15191), .CLK(clk), .RST(rst), .Q(ereg[186]) );
  DFF \ereg_reg[187]  ( .D(n15190), .CLK(clk), .RST(rst), .Q(ereg[187]) );
  DFF \ereg_reg[188]  ( .D(n15189), .CLK(clk), .RST(rst), .Q(ereg[188]) );
  DFF \ereg_reg[189]  ( .D(n15188), .CLK(clk), .RST(rst), .Q(ereg[189]) );
  DFF \ereg_reg[190]  ( .D(n15187), .CLK(clk), .RST(rst), .Q(ereg[190]) );
  DFF \ereg_reg[191]  ( .D(n15186), .CLK(clk), .RST(rst), .Q(ereg[191]) );
  DFF \ereg_reg[192]  ( .D(n15185), .CLK(clk), .RST(rst), .Q(ereg[192]) );
  DFF \ereg_reg[193]  ( .D(n15184), .CLK(clk), .RST(rst), .Q(ereg[193]) );
  DFF \ereg_reg[194]  ( .D(n15183), .CLK(clk), .RST(rst), .Q(ereg[194]) );
  DFF \ereg_reg[195]  ( .D(n15182), .CLK(clk), .RST(rst), .Q(ereg[195]) );
  DFF \ereg_reg[196]  ( .D(n15181), .CLK(clk), .RST(rst), .Q(ereg[196]) );
  DFF \ereg_reg[197]  ( .D(n15180), .CLK(clk), .RST(rst), .Q(ereg[197]) );
  DFF \ereg_reg[198]  ( .D(n15179), .CLK(clk), .RST(rst), .Q(ereg[198]) );
  DFF \ereg_reg[199]  ( .D(n15178), .CLK(clk), .RST(rst), .Q(ereg[199]) );
  DFF \ereg_reg[200]  ( .D(n15177), .CLK(clk), .RST(rst), .Q(ereg[200]) );
  DFF \ereg_reg[201]  ( .D(n15176), .CLK(clk), .RST(rst), .Q(ereg[201]) );
  DFF \ereg_reg[202]  ( .D(n15175), .CLK(clk), .RST(rst), .Q(ereg[202]) );
  DFF \ereg_reg[203]  ( .D(n15174), .CLK(clk), .RST(rst), .Q(ereg[203]) );
  DFF \ereg_reg[204]  ( .D(n15173), .CLK(clk), .RST(rst), .Q(ereg[204]) );
  DFF \ereg_reg[205]  ( .D(n15172), .CLK(clk), .RST(rst), .Q(ereg[205]) );
  DFF \ereg_reg[206]  ( .D(n15171), .CLK(clk), .RST(rst), .Q(ereg[206]) );
  DFF \ereg_reg[207]  ( .D(n15170), .CLK(clk), .RST(rst), .Q(ereg[207]) );
  DFF \ereg_reg[208]  ( .D(n15169), .CLK(clk), .RST(rst), .Q(ereg[208]) );
  DFF \ereg_reg[209]  ( .D(n15168), .CLK(clk), .RST(rst), .Q(ereg[209]) );
  DFF \ereg_reg[210]  ( .D(n15167), .CLK(clk), .RST(rst), .Q(ereg[210]) );
  DFF \ereg_reg[211]  ( .D(n15166), .CLK(clk), .RST(rst), .Q(ereg[211]) );
  DFF \ereg_reg[212]  ( .D(n15165), .CLK(clk), .RST(rst), .Q(ereg[212]) );
  DFF \ereg_reg[213]  ( .D(n15164), .CLK(clk), .RST(rst), .Q(ereg[213]) );
  DFF \ereg_reg[214]  ( .D(n15163), .CLK(clk), .RST(rst), .Q(ereg[214]) );
  DFF \ereg_reg[215]  ( .D(n15162), .CLK(clk), .RST(rst), .Q(ereg[215]) );
  DFF \ereg_reg[216]  ( .D(n15161), .CLK(clk), .RST(rst), .Q(ereg[216]) );
  DFF \ereg_reg[217]  ( .D(n15160), .CLK(clk), .RST(rst), .Q(ereg[217]) );
  DFF \ereg_reg[218]  ( .D(n15159), .CLK(clk), .RST(rst), .Q(ereg[218]) );
  DFF \ereg_reg[219]  ( .D(n15158), .CLK(clk), .RST(rst), .Q(ereg[219]) );
  DFF \ereg_reg[220]  ( .D(n15157), .CLK(clk), .RST(rst), .Q(ereg[220]) );
  DFF \ereg_reg[221]  ( .D(n15156), .CLK(clk), .RST(rst), .Q(ereg[221]) );
  DFF \ereg_reg[222]  ( .D(n15155), .CLK(clk), .RST(rst), .Q(ereg[222]) );
  DFF \ereg_reg[223]  ( .D(n15154), .CLK(clk), .RST(rst), .Q(ereg[223]) );
  DFF \ereg_reg[224]  ( .D(n15153), .CLK(clk), .RST(rst), .Q(ereg[224]) );
  DFF \ereg_reg[225]  ( .D(n15152), .CLK(clk), .RST(rst), .Q(ereg[225]) );
  DFF \ereg_reg[226]  ( .D(n15151), .CLK(clk), .RST(rst), .Q(ereg[226]) );
  DFF \ereg_reg[227]  ( .D(n15150), .CLK(clk), .RST(rst), .Q(ereg[227]) );
  DFF \ereg_reg[228]  ( .D(n15149), .CLK(clk), .RST(rst), .Q(ereg[228]) );
  DFF \ereg_reg[229]  ( .D(n15148), .CLK(clk), .RST(rst), .Q(ereg[229]) );
  DFF \ereg_reg[230]  ( .D(n15147), .CLK(clk), .RST(rst), .Q(ereg[230]) );
  DFF \ereg_reg[231]  ( .D(n15146), .CLK(clk), .RST(rst), .Q(ereg[231]) );
  DFF \ereg_reg[232]  ( .D(n15145), .CLK(clk), .RST(rst), .Q(ereg[232]) );
  DFF \ereg_reg[233]  ( .D(n15144), .CLK(clk), .RST(rst), .Q(ereg[233]) );
  DFF \ereg_reg[234]  ( .D(n15143), .CLK(clk), .RST(rst), .Q(ereg[234]) );
  DFF \ereg_reg[235]  ( .D(n15142), .CLK(clk), .RST(rst), .Q(ereg[235]) );
  DFF \ereg_reg[236]  ( .D(n15141), .CLK(clk), .RST(rst), .Q(ereg[236]) );
  DFF \ereg_reg[237]  ( .D(n15140), .CLK(clk), .RST(rst), .Q(ereg[237]) );
  DFF \ereg_reg[238]  ( .D(n15139), .CLK(clk), .RST(rst), .Q(ereg[238]) );
  DFF \ereg_reg[239]  ( .D(n15138), .CLK(clk), .RST(rst), .Q(ereg[239]) );
  DFF \ereg_reg[240]  ( .D(n15137), .CLK(clk), .RST(rst), .Q(ereg[240]) );
  DFF \ereg_reg[241]  ( .D(n15136), .CLK(clk), .RST(rst), .Q(ereg[241]) );
  DFF \ereg_reg[242]  ( .D(n15135), .CLK(clk), .RST(rst), .Q(ereg[242]) );
  DFF \ereg_reg[243]  ( .D(n15134), .CLK(clk), .RST(rst), .Q(ereg[243]) );
  DFF \ereg_reg[244]  ( .D(n15133), .CLK(clk), .RST(rst), .Q(ereg[244]) );
  DFF \ereg_reg[245]  ( .D(n15132), .CLK(clk), .RST(rst), .Q(ereg[245]) );
  DFF \ereg_reg[246]  ( .D(n15131), .CLK(clk), .RST(rst), .Q(ereg[246]) );
  DFF \ereg_reg[247]  ( .D(n15130), .CLK(clk), .RST(rst), .Q(ereg[247]) );
  DFF \ereg_reg[248]  ( .D(n15129), .CLK(clk), .RST(rst), .Q(ereg[248]) );
  DFF \ereg_reg[249]  ( .D(n15128), .CLK(clk), .RST(rst), .Q(ereg[249]) );
  DFF \ereg_reg[250]  ( .D(n15127), .CLK(clk), .RST(rst), .Q(ereg[250]) );
  DFF \ereg_reg[251]  ( .D(n15126), .CLK(clk), .RST(rst), .Q(ereg[251]) );
  DFF \ereg_reg[252]  ( .D(n15125), .CLK(clk), .RST(rst), .Q(ereg[252]) );
  DFF \ereg_reg[253]  ( .D(n15124), .CLK(clk), .RST(rst), .Q(ereg[253]) );
  DFF \ereg_reg[254]  ( .D(n15123), .CLK(clk), .RST(rst), .Q(ereg[254]) );
  DFF \ereg_reg[255]  ( .D(n15122), .CLK(clk), .RST(rst), .Q(ereg[255]) );
  DFF \ereg_reg[256]  ( .D(n15121), .CLK(clk), .RST(rst), .Q(ereg[256]) );
  DFF \ereg_reg[257]  ( .D(n15120), .CLK(clk), .RST(rst), .Q(ereg[257]) );
  DFF \ereg_reg[258]  ( .D(n15119), .CLK(clk), .RST(rst), .Q(ereg[258]) );
  DFF \ereg_reg[259]  ( .D(n15118), .CLK(clk), .RST(rst), .Q(ereg[259]) );
  DFF \ereg_reg[260]  ( .D(n15117), .CLK(clk), .RST(rst), .Q(ereg[260]) );
  DFF \ereg_reg[261]  ( .D(n15116), .CLK(clk), .RST(rst), .Q(ereg[261]) );
  DFF \ereg_reg[262]  ( .D(n15115), .CLK(clk), .RST(rst), .Q(ereg[262]) );
  DFF \ereg_reg[263]  ( .D(n15114), .CLK(clk), .RST(rst), .Q(ereg[263]) );
  DFF \ereg_reg[264]  ( .D(n15113), .CLK(clk), .RST(rst), .Q(ereg[264]) );
  DFF \ereg_reg[265]  ( .D(n15112), .CLK(clk), .RST(rst), .Q(ereg[265]) );
  DFF \ereg_reg[266]  ( .D(n15111), .CLK(clk), .RST(rst), .Q(ereg[266]) );
  DFF \ereg_reg[267]  ( .D(n15110), .CLK(clk), .RST(rst), .Q(ereg[267]) );
  DFF \ereg_reg[268]  ( .D(n15109), .CLK(clk), .RST(rst), .Q(ereg[268]) );
  DFF \ereg_reg[269]  ( .D(n15108), .CLK(clk), .RST(rst), .Q(ereg[269]) );
  DFF \ereg_reg[270]  ( .D(n15107), .CLK(clk), .RST(rst), .Q(ereg[270]) );
  DFF \ereg_reg[271]  ( .D(n15106), .CLK(clk), .RST(rst), .Q(ereg[271]) );
  DFF \ereg_reg[272]  ( .D(n15105), .CLK(clk), .RST(rst), .Q(ereg[272]) );
  DFF \ereg_reg[273]  ( .D(n15104), .CLK(clk), .RST(rst), .Q(ereg[273]) );
  DFF \ereg_reg[274]  ( .D(n15103), .CLK(clk), .RST(rst), .Q(ereg[274]) );
  DFF \ereg_reg[275]  ( .D(n15102), .CLK(clk), .RST(rst), .Q(ereg[275]) );
  DFF \ereg_reg[276]  ( .D(n15101), .CLK(clk), .RST(rst), .Q(ereg[276]) );
  DFF \ereg_reg[277]  ( .D(n15100), .CLK(clk), .RST(rst), .Q(ereg[277]) );
  DFF \ereg_reg[278]  ( .D(n15099), .CLK(clk), .RST(rst), .Q(ereg[278]) );
  DFF \ereg_reg[279]  ( .D(n15098), .CLK(clk), .RST(rst), .Q(ereg[279]) );
  DFF \ereg_reg[280]  ( .D(n15097), .CLK(clk), .RST(rst), .Q(ereg[280]) );
  DFF \ereg_reg[281]  ( .D(n15096), .CLK(clk), .RST(rst), .Q(ereg[281]) );
  DFF \ereg_reg[282]  ( .D(n15095), .CLK(clk), .RST(rst), .Q(ereg[282]) );
  DFF \ereg_reg[283]  ( .D(n15094), .CLK(clk), .RST(rst), .Q(ereg[283]) );
  DFF \ereg_reg[284]  ( .D(n15093), .CLK(clk), .RST(rst), .Q(ereg[284]) );
  DFF \ereg_reg[285]  ( .D(n15092), .CLK(clk), .RST(rst), .Q(ereg[285]) );
  DFF \ereg_reg[286]  ( .D(n15091), .CLK(clk), .RST(rst), .Q(ereg[286]) );
  DFF \ereg_reg[287]  ( .D(n15090), .CLK(clk), .RST(rst), .Q(ereg[287]) );
  DFF \ereg_reg[288]  ( .D(n15089), .CLK(clk), .RST(rst), .Q(ereg[288]) );
  DFF \ereg_reg[289]  ( .D(n15088), .CLK(clk), .RST(rst), .Q(ereg[289]) );
  DFF \ereg_reg[290]  ( .D(n15087), .CLK(clk), .RST(rst), .Q(ereg[290]) );
  DFF \ereg_reg[291]  ( .D(n15086), .CLK(clk), .RST(rst), .Q(ereg[291]) );
  DFF \ereg_reg[292]  ( .D(n15085), .CLK(clk), .RST(rst), .Q(ereg[292]) );
  DFF \ereg_reg[293]  ( .D(n15084), .CLK(clk), .RST(rst), .Q(ereg[293]) );
  DFF \ereg_reg[294]  ( .D(n15083), .CLK(clk), .RST(rst), .Q(ereg[294]) );
  DFF \ereg_reg[295]  ( .D(n15082), .CLK(clk), .RST(rst), .Q(ereg[295]) );
  DFF \ereg_reg[296]  ( .D(n15081), .CLK(clk), .RST(rst), .Q(ereg[296]) );
  DFF \ereg_reg[297]  ( .D(n15080), .CLK(clk), .RST(rst), .Q(ereg[297]) );
  DFF \ereg_reg[298]  ( .D(n15079), .CLK(clk), .RST(rst), .Q(ereg[298]) );
  DFF \ereg_reg[299]  ( .D(n15078), .CLK(clk), .RST(rst), .Q(ereg[299]) );
  DFF \ereg_reg[300]  ( .D(n15077), .CLK(clk), .RST(rst), .Q(ereg[300]) );
  DFF \ereg_reg[301]  ( .D(n15076), .CLK(clk), .RST(rst), .Q(ereg[301]) );
  DFF \ereg_reg[302]  ( .D(n15075), .CLK(clk), .RST(rst), .Q(ereg[302]) );
  DFF \ereg_reg[303]  ( .D(n15074), .CLK(clk), .RST(rst), .Q(ereg[303]) );
  DFF \ereg_reg[304]  ( .D(n15073), .CLK(clk), .RST(rst), .Q(ereg[304]) );
  DFF \ereg_reg[305]  ( .D(n15072), .CLK(clk), .RST(rst), .Q(ereg[305]) );
  DFF \ereg_reg[306]  ( .D(n15071), .CLK(clk), .RST(rst), .Q(ereg[306]) );
  DFF \ereg_reg[307]  ( .D(n15070), .CLK(clk), .RST(rst), .Q(ereg[307]) );
  DFF \ereg_reg[308]  ( .D(n15069), .CLK(clk), .RST(rst), .Q(ereg[308]) );
  DFF \ereg_reg[309]  ( .D(n15068), .CLK(clk), .RST(rst), .Q(ereg[309]) );
  DFF \ereg_reg[310]  ( .D(n15067), .CLK(clk), .RST(rst), .Q(ereg[310]) );
  DFF \ereg_reg[311]  ( .D(n15066), .CLK(clk), .RST(rst), .Q(ereg[311]) );
  DFF \ereg_reg[312]  ( .D(n15065), .CLK(clk), .RST(rst), .Q(ereg[312]) );
  DFF \ereg_reg[313]  ( .D(n15064), .CLK(clk), .RST(rst), .Q(ereg[313]) );
  DFF \ereg_reg[314]  ( .D(n15063), .CLK(clk), .RST(rst), .Q(ereg[314]) );
  DFF \ereg_reg[315]  ( .D(n15062), .CLK(clk), .RST(rst), .Q(ereg[315]) );
  DFF \ereg_reg[316]  ( .D(n15061), .CLK(clk), .RST(rst), .Q(ereg[316]) );
  DFF \ereg_reg[317]  ( .D(n15060), .CLK(clk), .RST(rst), .Q(ereg[317]) );
  DFF \ereg_reg[318]  ( .D(n15059), .CLK(clk), .RST(rst), .Q(ereg[318]) );
  DFF \ereg_reg[319]  ( .D(n15058), .CLK(clk), .RST(rst), .Q(ereg[319]) );
  DFF \ereg_reg[320]  ( .D(n15057), .CLK(clk), .RST(rst), .Q(ereg[320]) );
  DFF \ereg_reg[321]  ( .D(n15056), .CLK(clk), .RST(rst), .Q(ereg[321]) );
  DFF \ereg_reg[322]  ( .D(n15055), .CLK(clk), .RST(rst), .Q(ereg[322]) );
  DFF \ereg_reg[323]  ( .D(n15054), .CLK(clk), .RST(rst), .Q(ereg[323]) );
  DFF \ereg_reg[324]  ( .D(n15053), .CLK(clk), .RST(rst), .Q(ereg[324]) );
  DFF \ereg_reg[325]  ( .D(n15052), .CLK(clk), .RST(rst), .Q(ereg[325]) );
  DFF \ereg_reg[326]  ( .D(n15051), .CLK(clk), .RST(rst), .Q(ereg[326]) );
  DFF \ereg_reg[327]  ( .D(n15050), .CLK(clk), .RST(rst), .Q(ereg[327]) );
  DFF \ereg_reg[328]  ( .D(n15049), .CLK(clk), .RST(rst), .Q(ereg[328]) );
  DFF \ereg_reg[329]  ( .D(n15048), .CLK(clk), .RST(rst), .Q(ereg[329]) );
  DFF \ereg_reg[330]  ( .D(n15047), .CLK(clk), .RST(rst), .Q(ereg[330]) );
  DFF \ereg_reg[331]  ( .D(n15046), .CLK(clk), .RST(rst), .Q(ereg[331]) );
  DFF \ereg_reg[332]  ( .D(n15045), .CLK(clk), .RST(rst), .Q(ereg[332]) );
  DFF \ereg_reg[333]  ( .D(n15044), .CLK(clk), .RST(rst), .Q(ereg[333]) );
  DFF \ereg_reg[334]  ( .D(n15043), .CLK(clk), .RST(rst), .Q(ereg[334]) );
  DFF \ereg_reg[335]  ( .D(n15042), .CLK(clk), .RST(rst), .Q(ereg[335]) );
  DFF \ereg_reg[336]  ( .D(n15041), .CLK(clk), .RST(rst), .Q(ereg[336]) );
  DFF \ereg_reg[337]  ( .D(n15040), .CLK(clk), .RST(rst), .Q(ereg[337]) );
  DFF \ereg_reg[338]  ( .D(n15039), .CLK(clk), .RST(rst), .Q(ereg[338]) );
  DFF \ereg_reg[339]  ( .D(n15038), .CLK(clk), .RST(rst), .Q(ereg[339]) );
  DFF \ereg_reg[340]  ( .D(n15037), .CLK(clk), .RST(rst), .Q(ereg[340]) );
  DFF \ereg_reg[341]  ( .D(n15036), .CLK(clk), .RST(rst), .Q(ereg[341]) );
  DFF \ereg_reg[342]  ( .D(n15035), .CLK(clk), .RST(rst), .Q(ereg[342]) );
  DFF \ereg_reg[343]  ( .D(n15034), .CLK(clk), .RST(rst), .Q(ereg[343]) );
  DFF \ereg_reg[344]  ( .D(n15033), .CLK(clk), .RST(rst), .Q(ereg[344]) );
  DFF \ereg_reg[345]  ( .D(n15032), .CLK(clk), .RST(rst), .Q(ereg[345]) );
  DFF \ereg_reg[346]  ( .D(n15031), .CLK(clk), .RST(rst), .Q(ereg[346]) );
  DFF \ereg_reg[347]  ( .D(n15030), .CLK(clk), .RST(rst), .Q(ereg[347]) );
  DFF \ereg_reg[348]  ( .D(n15029), .CLK(clk), .RST(rst), .Q(ereg[348]) );
  DFF \ereg_reg[349]  ( .D(n15028), .CLK(clk), .RST(rst), .Q(ereg[349]) );
  DFF \ereg_reg[350]  ( .D(n15027), .CLK(clk), .RST(rst), .Q(ereg[350]) );
  DFF \ereg_reg[351]  ( .D(n15026), .CLK(clk), .RST(rst), .Q(ereg[351]) );
  DFF \ereg_reg[352]  ( .D(n15025), .CLK(clk), .RST(rst), .Q(ereg[352]) );
  DFF \ereg_reg[353]  ( .D(n15024), .CLK(clk), .RST(rst), .Q(ereg[353]) );
  DFF \ereg_reg[354]  ( .D(n15023), .CLK(clk), .RST(rst), .Q(ereg[354]) );
  DFF \ereg_reg[355]  ( .D(n15022), .CLK(clk), .RST(rst), .Q(ereg[355]) );
  DFF \ereg_reg[356]  ( .D(n15021), .CLK(clk), .RST(rst), .Q(ereg[356]) );
  DFF \ereg_reg[357]  ( .D(n15020), .CLK(clk), .RST(rst), .Q(ereg[357]) );
  DFF \ereg_reg[358]  ( .D(n15019), .CLK(clk), .RST(rst), .Q(ereg[358]) );
  DFF \ereg_reg[359]  ( .D(n15018), .CLK(clk), .RST(rst), .Q(ereg[359]) );
  DFF \ereg_reg[360]  ( .D(n15017), .CLK(clk), .RST(rst), .Q(ereg[360]) );
  DFF \ereg_reg[361]  ( .D(n15016), .CLK(clk), .RST(rst), .Q(ereg[361]) );
  DFF \ereg_reg[362]  ( .D(n15015), .CLK(clk), .RST(rst), .Q(ereg[362]) );
  DFF \ereg_reg[363]  ( .D(n15014), .CLK(clk), .RST(rst), .Q(ereg[363]) );
  DFF \ereg_reg[364]  ( .D(n15013), .CLK(clk), .RST(rst), .Q(ereg[364]) );
  DFF \ereg_reg[365]  ( .D(n15012), .CLK(clk), .RST(rst), .Q(ereg[365]) );
  DFF \ereg_reg[366]  ( .D(n15011), .CLK(clk), .RST(rst), .Q(ereg[366]) );
  DFF \ereg_reg[367]  ( .D(n15010), .CLK(clk), .RST(rst), .Q(ereg[367]) );
  DFF \ereg_reg[368]  ( .D(n15009), .CLK(clk), .RST(rst), .Q(ereg[368]) );
  DFF \ereg_reg[369]  ( .D(n15008), .CLK(clk), .RST(rst), .Q(ereg[369]) );
  DFF \ereg_reg[370]  ( .D(n15007), .CLK(clk), .RST(rst), .Q(ereg[370]) );
  DFF \ereg_reg[371]  ( .D(n15006), .CLK(clk), .RST(rst), .Q(ereg[371]) );
  DFF \ereg_reg[372]  ( .D(n15005), .CLK(clk), .RST(rst), .Q(ereg[372]) );
  DFF \ereg_reg[373]  ( .D(n15004), .CLK(clk), .RST(rst), .Q(ereg[373]) );
  DFF \ereg_reg[374]  ( .D(n15003), .CLK(clk), .RST(rst), .Q(ereg[374]) );
  DFF \ereg_reg[375]  ( .D(n15002), .CLK(clk), .RST(rst), .Q(ereg[375]) );
  DFF \ereg_reg[376]  ( .D(n15001), .CLK(clk), .RST(rst), .Q(ereg[376]) );
  DFF \ereg_reg[377]  ( .D(n15000), .CLK(clk), .RST(rst), .Q(ereg[377]) );
  DFF \ereg_reg[378]  ( .D(n14999), .CLK(clk), .RST(rst), .Q(ereg[378]) );
  DFF \ereg_reg[379]  ( .D(n14998), .CLK(clk), .RST(rst), .Q(ereg[379]) );
  DFF \ereg_reg[380]  ( .D(n14997), .CLK(clk), .RST(rst), .Q(ereg[380]) );
  DFF \ereg_reg[381]  ( .D(n14996), .CLK(clk), .RST(rst), .Q(ereg[381]) );
  DFF \ereg_reg[382]  ( .D(n14995), .CLK(clk), .RST(rst), .Q(ereg[382]) );
  DFF \ereg_reg[383]  ( .D(n14994), .CLK(clk), .RST(rst), .Q(ereg[383]) );
  DFF \ereg_reg[384]  ( .D(n14993), .CLK(clk), .RST(rst), .Q(ereg[384]) );
  DFF \ereg_reg[385]  ( .D(n14992), .CLK(clk), .RST(rst), .Q(ereg[385]) );
  DFF \ereg_reg[386]  ( .D(n14991), .CLK(clk), .RST(rst), .Q(ereg[386]) );
  DFF \ereg_reg[387]  ( .D(n14990), .CLK(clk), .RST(rst), .Q(ereg[387]) );
  DFF \ereg_reg[388]  ( .D(n14989), .CLK(clk), .RST(rst), .Q(ereg[388]) );
  DFF \ereg_reg[389]  ( .D(n14988), .CLK(clk), .RST(rst), .Q(ereg[389]) );
  DFF \ereg_reg[390]  ( .D(n14987), .CLK(clk), .RST(rst), .Q(ereg[390]) );
  DFF \ereg_reg[391]  ( .D(n14986), .CLK(clk), .RST(rst), .Q(ereg[391]) );
  DFF \ereg_reg[392]  ( .D(n14985), .CLK(clk), .RST(rst), .Q(ereg[392]) );
  DFF \ereg_reg[393]  ( .D(n14984), .CLK(clk), .RST(rst), .Q(ereg[393]) );
  DFF \ereg_reg[394]  ( .D(n14983), .CLK(clk), .RST(rst), .Q(ereg[394]) );
  DFF \ereg_reg[395]  ( .D(n14982), .CLK(clk), .RST(rst), .Q(ereg[395]) );
  DFF \ereg_reg[396]  ( .D(n14981), .CLK(clk), .RST(rst), .Q(ereg[396]) );
  DFF \ereg_reg[397]  ( .D(n14980), .CLK(clk), .RST(rst), .Q(ereg[397]) );
  DFF \ereg_reg[398]  ( .D(n14979), .CLK(clk), .RST(rst), .Q(ereg[398]) );
  DFF \ereg_reg[399]  ( .D(n14978), .CLK(clk), .RST(rst), .Q(ereg[399]) );
  DFF \ereg_reg[400]  ( .D(n14977), .CLK(clk), .RST(rst), .Q(ereg[400]) );
  DFF \ereg_reg[401]  ( .D(n14976), .CLK(clk), .RST(rst), .Q(ereg[401]) );
  DFF \ereg_reg[402]  ( .D(n14975), .CLK(clk), .RST(rst), .Q(ereg[402]) );
  DFF \ereg_reg[403]  ( .D(n14974), .CLK(clk), .RST(rst), .Q(ereg[403]) );
  DFF \ereg_reg[404]  ( .D(n14973), .CLK(clk), .RST(rst), .Q(ereg[404]) );
  DFF \ereg_reg[405]  ( .D(n14972), .CLK(clk), .RST(rst), .Q(ereg[405]) );
  DFF \ereg_reg[406]  ( .D(n14971), .CLK(clk), .RST(rst), .Q(ereg[406]) );
  DFF \ereg_reg[407]  ( .D(n14970), .CLK(clk), .RST(rst), .Q(ereg[407]) );
  DFF \ereg_reg[408]  ( .D(n14969), .CLK(clk), .RST(rst), .Q(ereg[408]) );
  DFF \ereg_reg[409]  ( .D(n14968), .CLK(clk), .RST(rst), .Q(ereg[409]) );
  DFF \ereg_reg[410]  ( .D(n14967), .CLK(clk), .RST(rst), .Q(ereg[410]) );
  DFF \ereg_reg[411]  ( .D(n14966), .CLK(clk), .RST(rst), .Q(ereg[411]) );
  DFF \ereg_reg[412]  ( .D(n14965), .CLK(clk), .RST(rst), .Q(ereg[412]) );
  DFF \ereg_reg[413]  ( .D(n14964), .CLK(clk), .RST(rst), .Q(ereg[413]) );
  DFF \ereg_reg[414]  ( .D(n14963), .CLK(clk), .RST(rst), .Q(ereg[414]) );
  DFF \ereg_reg[415]  ( .D(n14962), .CLK(clk), .RST(rst), .Q(ereg[415]) );
  DFF \ereg_reg[416]  ( .D(n14961), .CLK(clk), .RST(rst), .Q(ereg[416]) );
  DFF \ereg_reg[417]  ( .D(n14960), .CLK(clk), .RST(rst), .Q(ereg[417]) );
  DFF \ereg_reg[418]  ( .D(n14959), .CLK(clk), .RST(rst), .Q(ereg[418]) );
  DFF \ereg_reg[419]  ( .D(n14958), .CLK(clk), .RST(rst), .Q(ereg[419]) );
  DFF \ereg_reg[420]  ( .D(n14957), .CLK(clk), .RST(rst), .Q(ereg[420]) );
  DFF \ereg_reg[421]  ( .D(n14956), .CLK(clk), .RST(rst), .Q(ereg[421]) );
  DFF \ereg_reg[422]  ( .D(n14955), .CLK(clk), .RST(rst), .Q(ereg[422]) );
  DFF \ereg_reg[423]  ( .D(n14954), .CLK(clk), .RST(rst), .Q(ereg[423]) );
  DFF \ereg_reg[424]  ( .D(n14953), .CLK(clk), .RST(rst), .Q(ereg[424]) );
  DFF \ereg_reg[425]  ( .D(n14952), .CLK(clk), .RST(rst), .Q(ereg[425]) );
  DFF \ereg_reg[426]  ( .D(n14951), .CLK(clk), .RST(rst), .Q(ereg[426]) );
  DFF \ereg_reg[427]  ( .D(n14950), .CLK(clk), .RST(rst), .Q(ereg[427]) );
  DFF \ereg_reg[428]  ( .D(n14949), .CLK(clk), .RST(rst), .Q(ereg[428]) );
  DFF \ereg_reg[429]  ( .D(n14948), .CLK(clk), .RST(rst), .Q(ereg[429]) );
  DFF \ereg_reg[430]  ( .D(n14947), .CLK(clk), .RST(rst), .Q(ereg[430]) );
  DFF \ereg_reg[431]  ( .D(n14946), .CLK(clk), .RST(rst), .Q(ereg[431]) );
  DFF \ereg_reg[432]  ( .D(n14945), .CLK(clk), .RST(rst), .Q(ereg[432]) );
  DFF \ereg_reg[433]  ( .D(n14944), .CLK(clk), .RST(rst), .Q(ereg[433]) );
  DFF \ereg_reg[434]  ( .D(n14943), .CLK(clk), .RST(rst), .Q(ereg[434]) );
  DFF \ereg_reg[435]  ( .D(n14942), .CLK(clk), .RST(rst), .Q(ereg[435]) );
  DFF \ereg_reg[436]  ( .D(n14941), .CLK(clk), .RST(rst), .Q(ereg[436]) );
  DFF \ereg_reg[437]  ( .D(n14940), .CLK(clk), .RST(rst), .Q(ereg[437]) );
  DFF \ereg_reg[438]  ( .D(n14939), .CLK(clk), .RST(rst), .Q(ereg[438]) );
  DFF \ereg_reg[439]  ( .D(n14938), .CLK(clk), .RST(rst), .Q(ereg[439]) );
  DFF \ereg_reg[440]  ( .D(n14937), .CLK(clk), .RST(rst), .Q(ereg[440]) );
  DFF \ereg_reg[441]  ( .D(n14936), .CLK(clk), .RST(rst), .Q(ereg[441]) );
  DFF \ereg_reg[442]  ( .D(n14935), .CLK(clk), .RST(rst), .Q(ereg[442]) );
  DFF \ereg_reg[443]  ( .D(n14934), .CLK(clk), .RST(rst), .Q(ereg[443]) );
  DFF \ereg_reg[444]  ( .D(n14933), .CLK(clk), .RST(rst), .Q(ereg[444]) );
  DFF \ereg_reg[445]  ( .D(n14932), .CLK(clk), .RST(rst), .Q(ereg[445]) );
  DFF \ereg_reg[446]  ( .D(n14931), .CLK(clk), .RST(rst), .Q(ereg[446]) );
  DFF \ereg_reg[447]  ( .D(n14930), .CLK(clk), .RST(rst), .Q(ereg[447]) );
  DFF \ereg_reg[448]  ( .D(n14929), .CLK(clk), .RST(rst), .Q(ereg[448]) );
  DFF \ereg_reg[449]  ( .D(n14928), .CLK(clk), .RST(rst), .Q(ereg[449]) );
  DFF \ereg_reg[450]  ( .D(n14927), .CLK(clk), .RST(rst), .Q(ereg[450]) );
  DFF \ereg_reg[451]  ( .D(n14926), .CLK(clk), .RST(rst), .Q(ereg[451]) );
  DFF \ereg_reg[452]  ( .D(n14925), .CLK(clk), .RST(rst), .Q(ereg[452]) );
  DFF \ereg_reg[453]  ( .D(n14924), .CLK(clk), .RST(rst), .Q(ereg[453]) );
  DFF \ereg_reg[454]  ( .D(n14923), .CLK(clk), .RST(rst), .Q(ereg[454]) );
  DFF \ereg_reg[455]  ( .D(n14922), .CLK(clk), .RST(rst), .Q(ereg[455]) );
  DFF \ereg_reg[456]  ( .D(n14921), .CLK(clk), .RST(rst), .Q(ereg[456]) );
  DFF \ereg_reg[457]  ( .D(n14920), .CLK(clk), .RST(rst), .Q(ereg[457]) );
  DFF \ereg_reg[458]  ( .D(n14919), .CLK(clk), .RST(rst), .Q(ereg[458]) );
  DFF \ereg_reg[459]  ( .D(n14918), .CLK(clk), .RST(rst), .Q(ereg[459]) );
  DFF \ereg_reg[460]  ( .D(n14917), .CLK(clk), .RST(rst), .Q(ereg[460]) );
  DFF \ereg_reg[461]  ( .D(n14916), .CLK(clk), .RST(rst), .Q(ereg[461]) );
  DFF \ereg_reg[462]  ( .D(n14915), .CLK(clk), .RST(rst), .Q(ereg[462]) );
  DFF \ereg_reg[463]  ( .D(n14914), .CLK(clk), .RST(rst), .Q(ereg[463]) );
  DFF \ereg_reg[464]  ( .D(n14913), .CLK(clk), .RST(rst), .Q(ereg[464]) );
  DFF \ereg_reg[465]  ( .D(n14912), .CLK(clk), .RST(rst), .Q(ereg[465]) );
  DFF \ereg_reg[466]  ( .D(n14911), .CLK(clk), .RST(rst), .Q(ereg[466]) );
  DFF \ereg_reg[467]  ( .D(n14910), .CLK(clk), .RST(rst), .Q(ereg[467]) );
  DFF \ereg_reg[468]  ( .D(n14909), .CLK(clk), .RST(rst), .Q(ereg[468]) );
  DFF \ereg_reg[469]  ( .D(n14908), .CLK(clk), .RST(rst), .Q(ereg[469]) );
  DFF \ereg_reg[470]  ( .D(n14907), .CLK(clk), .RST(rst), .Q(ereg[470]) );
  DFF \ereg_reg[471]  ( .D(n14906), .CLK(clk), .RST(rst), .Q(ereg[471]) );
  DFF \ereg_reg[472]  ( .D(n14905), .CLK(clk), .RST(rst), .Q(ereg[472]) );
  DFF \ereg_reg[473]  ( .D(n14904), .CLK(clk), .RST(rst), .Q(ereg[473]) );
  DFF \ereg_reg[474]  ( .D(n14903), .CLK(clk), .RST(rst), .Q(ereg[474]) );
  DFF \ereg_reg[475]  ( .D(n14902), .CLK(clk), .RST(rst), .Q(ereg[475]) );
  DFF \ereg_reg[476]  ( .D(n14901), .CLK(clk), .RST(rst), .Q(ereg[476]) );
  DFF \ereg_reg[477]  ( .D(n14900), .CLK(clk), .RST(rst), .Q(ereg[477]) );
  DFF \ereg_reg[478]  ( .D(n14899), .CLK(clk), .RST(rst), .Q(ereg[478]) );
  DFF \ereg_reg[479]  ( .D(n14898), .CLK(clk), .RST(rst), .Q(ereg[479]) );
  DFF \ereg_reg[480]  ( .D(n14897), .CLK(clk), .RST(rst), .Q(ereg[480]) );
  DFF \ereg_reg[481]  ( .D(n14896), .CLK(clk), .RST(rst), .Q(ereg[481]) );
  DFF \ereg_reg[482]  ( .D(n14895), .CLK(clk), .RST(rst), .Q(ereg[482]) );
  DFF \ereg_reg[483]  ( .D(n14894), .CLK(clk), .RST(rst), .Q(ereg[483]) );
  DFF \ereg_reg[484]  ( .D(n14893), .CLK(clk), .RST(rst), .Q(ereg[484]) );
  DFF \ereg_reg[485]  ( .D(n14892), .CLK(clk), .RST(rst), .Q(ereg[485]) );
  DFF \ereg_reg[486]  ( .D(n14891), .CLK(clk), .RST(rst), .Q(ereg[486]) );
  DFF \ereg_reg[487]  ( .D(n14890), .CLK(clk), .RST(rst), .Q(ereg[487]) );
  DFF \ereg_reg[488]  ( .D(n14889), .CLK(clk), .RST(rst), .Q(ereg[488]) );
  DFF \ereg_reg[489]  ( .D(n14888), .CLK(clk), .RST(rst), .Q(ereg[489]) );
  DFF \ereg_reg[490]  ( .D(n14887), .CLK(clk), .RST(rst), .Q(ereg[490]) );
  DFF \ereg_reg[491]  ( .D(n14886), .CLK(clk), .RST(rst), .Q(ereg[491]) );
  DFF \ereg_reg[492]  ( .D(n14885), .CLK(clk), .RST(rst), .Q(ereg[492]) );
  DFF \ereg_reg[493]  ( .D(n14884), .CLK(clk), .RST(rst), .Q(ereg[493]) );
  DFF \ereg_reg[494]  ( .D(n14883), .CLK(clk), .RST(rst), .Q(ereg[494]) );
  DFF \ereg_reg[495]  ( .D(n14882), .CLK(clk), .RST(rst), .Q(ereg[495]) );
  DFF \ereg_reg[496]  ( .D(n14881), .CLK(clk), .RST(rst), .Q(ereg[496]) );
  DFF \ereg_reg[497]  ( .D(n14880), .CLK(clk), .RST(rst), .Q(ereg[497]) );
  DFF \ereg_reg[498]  ( .D(n14879), .CLK(clk), .RST(rst), .Q(ereg[498]) );
  DFF \ereg_reg[499]  ( .D(n14878), .CLK(clk), .RST(rst), .Q(ereg[499]) );
  DFF \ereg_reg[500]  ( .D(n14877), .CLK(clk), .RST(rst), .Q(ereg[500]) );
  DFF \ereg_reg[501]  ( .D(n14876), .CLK(clk), .RST(rst), .Q(ereg[501]) );
  DFF \ereg_reg[502]  ( .D(n14875), .CLK(clk), .RST(rst), .Q(ereg[502]) );
  DFF \ereg_reg[503]  ( .D(n14874), .CLK(clk), .RST(rst), .Q(ereg[503]) );
  DFF \ereg_reg[504]  ( .D(n14873), .CLK(clk), .RST(rst), .Q(ereg[504]) );
  DFF \ereg_reg[505]  ( .D(n14872), .CLK(clk), .RST(rst), .Q(ereg[505]) );
  DFF \ereg_reg[506]  ( .D(n14871), .CLK(clk), .RST(rst), .Q(ereg[506]) );
  DFF \ereg_reg[507]  ( .D(n14870), .CLK(clk), .RST(rst), .Q(ereg[507]) );
  DFF \ereg_reg[508]  ( .D(n14869), .CLK(clk), .RST(rst), .Q(ereg[508]) );
  DFF \ereg_reg[509]  ( .D(n14868), .CLK(clk), .RST(rst), .Q(ereg[509]) );
  DFF \ereg_reg[510]  ( .D(n14867), .CLK(clk), .RST(rst), .Q(ereg[510]) );
  DFF \ereg_reg[511]  ( .D(n14866), .CLK(clk), .RST(rst), .Q(ereg[511]) );
  DFF \ereg_reg[512]  ( .D(n14865), .CLK(clk), .RST(rst), .Q(ereg[512]) );
  DFF \ereg_reg[513]  ( .D(n14864), .CLK(clk), .RST(rst), .Q(ereg[513]) );
  DFF \ereg_reg[514]  ( .D(n14863), .CLK(clk), .RST(rst), .Q(ereg[514]) );
  DFF \ereg_reg[515]  ( .D(n14862), .CLK(clk), .RST(rst), .Q(ereg[515]) );
  DFF \ereg_reg[516]  ( .D(n14861), .CLK(clk), .RST(rst), .Q(ereg[516]) );
  DFF \ereg_reg[517]  ( .D(n14860), .CLK(clk), .RST(rst), .Q(ereg[517]) );
  DFF \ereg_reg[518]  ( .D(n14859), .CLK(clk), .RST(rst), .Q(ereg[518]) );
  DFF \ereg_reg[519]  ( .D(n14858), .CLK(clk), .RST(rst), .Q(ereg[519]) );
  DFF \ereg_reg[520]  ( .D(n14857), .CLK(clk), .RST(rst), .Q(ereg[520]) );
  DFF \ereg_reg[521]  ( .D(n14856), .CLK(clk), .RST(rst), .Q(ereg[521]) );
  DFF \ereg_reg[522]  ( .D(n14855), .CLK(clk), .RST(rst), .Q(ereg[522]) );
  DFF \ereg_reg[523]  ( .D(n14854), .CLK(clk), .RST(rst), .Q(ereg[523]) );
  DFF \ereg_reg[524]  ( .D(n14853), .CLK(clk), .RST(rst), .Q(ereg[524]) );
  DFF \ereg_reg[525]  ( .D(n14852), .CLK(clk), .RST(rst), .Q(ereg[525]) );
  DFF \ereg_reg[526]  ( .D(n14851), .CLK(clk), .RST(rst), .Q(ereg[526]) );
  DFF \ereg_reg[527]  ( .D(n14850), .CLK(clk), .RST(rst), .Q(ereg[527]) );
  DFF \ereg_reg[528]  ( .D(n14849), .CLK(clk), .RST(rst), .Q(ereg[528]) );
  DFF \ereg_reg[529]  ( .D(n14848), .CLK(clk), .RST(rst), .Q(ereg[529]) );
  DFF \ereg_reg[530]  ( .D(n14847), .CLK(clk), .RST(rst), .Q(ereg[530]) );
  DFF \ereg_reg[531]  ( .D(n14846), .CLK(clk), .RST(rst), .Q(ereg[531]) );
  DFF \ereg_reg[532]  ( .D(n14845), .CLK(clk), .RST(rst), .Q(ereg[532]) );
  DFF \ereg_reg[533]  ( .D(n14844), .CLK(clk), .RST(rst), .Q(ereg[533]) );
  DFF \ereg_reg[534]  ( .D(n14843), .CLK(clk), .RST(rst), .Q(ereg[534]) );
  DFF \ereg_reg[535]  ( .D(n14842), .CLK(clk), .RST(rst), .Q(ereg[535]) );
  DFF \ereg_reg[536]  ( .D(n14841), .CLK(clk), .RST(rst), .Q(ereg[536]) );
  DFF \ereg_reg[537]  ( .D(n14840), .CLK(clk), .RST(rst), .Q(ereg[537]) );
  DFF \ereg_reg[538]  ( .D(n14839), .CLK(clk), .RST(rst), .Q(ereg[538]) );
  DFF \ereg_reg[539]  ( .D(n14838), .CLK(clk), .RST(rst), .Q(ereg[539]) );
  DFF \ereg_reg[540]  ( .D(n14837), .CLK(clk), .RST(rst), .Q(ereg[540]) );
  DFF \ereg_reg[541]  ( .D(n14836), .CLK(clk), .RST(rst), .Q(ereg[541]) );
  DFF \ereg_reg[542]  ( .D(n14835), .CLK(clk), .RST(rst), .Q(ereg[542]) );
  DFF \ereg_reg[543]  ( .D(n14834), .CLK(clk), .RST(rst), .Q(ereg[543]) );
  DFF \ereg_reg[544]  ( .D(n14833), .CLK(clk), .RST(rst), .Q(ereg[544]) );
  DFF \ereg_reg[545]  ( .D(n14832), .CLK(clk), .RST(rst), .Q(ereg[545]) );
  DFF \ereg_reg[546]  ( .D(n14831), .CLK(clk), .RST(rst), .Q(ereg[546]) );
  DFF \ereg_reg[547]  ( .D(n14830), .CLK(clk), .RST(rst), .Q(ereg[547]) );
  DFF \ereg_reg[548]  ( .D(n14829), .CLK(clk), .RST(rst), .Q(ereg[548]) );
  DFF \ereg_reg[549]  ( .D(n14828), .CLK(clk), .RST(rst), .Q(ereg[549]) );
  DFF \ereg_reg[550]  ( .D(n14827), .CLK(clk), .RST(rst), .Q(ereg[550]) );
  DFF \ereg_reg[551]  ( .D(n14826), .CLK(clk), .RST(rst), .Q(ereg[551]) );
  DFF \ereg_reg[552]  ( .D(n14825), .CLK(clk), .RST(rst), .Q(ereg[552]) );
  DFF \ereg_reg[553]  ( .D(n14824), .CLK(clk), .RST(rst), .Q(ereg[553]) );
  DFF \ereg_reg[554]  ( .D(n14823), .CLK(clk), .RST(rst), .Q(ereg[554]) );
  DFF \ereg_reg[555]  ( .D(n14822), .CLK(clk), .RST(rst), .Q(ereg[555]) );
  DFF \ereg_reg[556]  ( .D(n14821), .CLK(clk), .RST(rst), .Q(ereg[556]) );
  DFF \ereg_reg[557]  ( .D(n14820), .CLK(clk), .RST(rst), .Q(ereg[557]) );
  DFF \ereg_reg[558]  ( .D(n14819), .CLK(clk), .RST(rst), .Q(ereg[558]) );
  DFF \ereg_reg[559]  ( .D(n14818), .CLK(clk), .RST(rst), .Q(ereg[559]) );
  DFF \ereg_reg[560]  ( .D(n14817), .CLK(clk), .RST(rst), .Q(ereg[560]) );
  DFF \ereg_reg[561]  ( .D(n14816), .CLK(clk), .RST(rst), .Q(ereg[561]) );
  DFF \ereg_reg[562]  ( .D(n14815), .CLK(clk), .RST(rst), .Q(ereg[562]) );
  DFF \ereg_reg[563]  ( .D(n14814), .CLK(clk), .RST(rst), .Q(ereg[563]) );
  DFF \ereg_reg[564]  ( .D(n14813), .CLK(clk), .RST(rst), .Q(ereg[564]) );
  DFF \ereg_reg[565]  ( .D(n14812), .CLK(clk), .RST(rst), .Q(ereg[565]) );
  DFF \ereg_reg[566]  ( .D(n14811), .CLK(clk), .RST(rst), .Q(ereg[566]) );
  DFF \ereg_reg[567]  ( .D(n14810), .CLK(clk), .RST(rst), .Q(ereg[567]) );
  DFF \ereg_reg[568]  ( .D(n14809), .CLK(clk), .RST(rst), .Q(ereg[568]) );
  DFF \ereg_reg[569]  ( .D(n14808), .CLK(clk), .RST(rst), .Q(ereg[569]) );
  DFF \ereg_reg[570]  ( .D(n14807), .CLK(clk), .RST(rst), .Q(ereg[570]) );
  DFF \ereg_reg[571]  ( .D(n14806), .CLK(clk), .RST(rst), .Q(ereg[571]) );
  DFF \ereg_reg[572]  ( .D(n14805), .CLK(clk), .RST(rst), .Q(ereg[572]) );
  DFF \ereg_reg[573]  ( .D(n14804), .CLK(clk), .RST(rst), .Q(ereg[573]) );
  DFF \ereg_reg[574]  ( .D(n14803), .CLK(clk), .RST(rst), .Q(ereg[574]) );
  DFF \ereg_reg[575]  ( .D(n14802), .CLK(clk), .RST(rst), .Q(ereg[575]) );
  DFF \ereg_reg[576]  ( .D(n14801), .CLK(clk), .RST(rst), .Q(ereg[576]) );
  DFF \ereg_reg[577]  ( .D(n14800), .CLK(clk), .RST(rst), .Q(ereg[577]) );
  DFF \ereg_reg[578]  ( .D(n14799), .CLK(clk), .RST(rst), .Q(ereg[578]) );
  DFF \ereg_reg[579]  ( .D(n14798), .CLK(clk), .RST(rst), .Q(ereg[579]) );
  DFF \ereg_reg[580]  ( .D(n14797), .CLK(clk), .RST(rst), .Q(ereg[580]) );
  DFF \ereg_reg[581]  ( .D(n14796), .CLK(clk), .RST(rst), .Q(ereg[581]) );
  DFF \ereg_reg[582]  ( .D(n14795), .CLK(clk), .RST(rst), .Q(ereg[582]) );
  DFF \ereg_reg[583]  ( .D(n14794), .CLK(clk), .RST(rst), .Q(ereg[583]) );
  DFF \ereg_reg[584]  ( .D(n14793), .CLK(clk), .RST(rst), .Q(ereg[584]) );
  DFF \ereg_reg[585]  ( .D(n14792), .CLK(clk), .RST(rst), .Q(ereg[585]) );
  DFF \ereg_reg[586]  ( .D(n14791), .CLK(clk), .RST(rst), .Q(ereg[586]) );
  DFF \ereg_reg[587]  ( .D(n14790), .CLK(clk), .RST(rst), .Q(ereg[587]) );
  DFF \ereg_reg[588]  ( .D(n14789), .CLK(clk), .RST(rst), .Q(ereg[588]) );
  DFF \ereg_reg[589]  ( .D(n14788), .CLK(clk), .RST(rst), .Q(ereg[589]) );
  DFF \ereg_reg[590]  ( .D(n14787), .CLK(clk), .RST(rst), .Q(ereg[590]) );
  DFF \ereg_reg[591]  ( .D(n14786), .CLK(clk), .RST(rst), .Q(ereg[591]) );
  DFF \ereg_reg[592]  ( .D(n14785), .CLK(clk), .RST(rst), .Q(ereg[592]) );
  DFF \ereg_reg[593]  ( .D(n14784), .CLK(clk), .RST(rst), .Q(ereg[593]) );
  DFF \ereg_reg[594]  ( .D(n14783), .CLK(clk), .RST(rst), .Q(ereg[594]) );
  DFF \ereg_reg[595]  ( .D(n14782), .CLK(clk), .RST(rst), .Q(ereg[595]) );
  DFF \ereg_reg[596]  ( .D(n14781), .CLK(clk), .RST(rst), .Q(ereg[596]) );
  DFF \ereg_reg[597]  ( .D(n14780), .CLK(clk), .RST(rst), .Q(ereg[597]) );
  DFF \ereg_reg[598]  ( .D(n14779), .CLK(clk), .RST(rst), .Q(ereg[598]) );
  DFF \ereg_reg[599]  ( .D(n14778), .CLK(clk), .RST(rst), .Q(ereg[599]) );
  DFF \ereg_reg[600]  ( .D(n14777), .CLK(clk), .RST(rst), .Q(ereg[600]) );
  DFF \ereg_reg[601]  ( .D(n14776), .CLK(clk), .RST(rst), .Q(ereg[601]) );
  DFF \ereg_reg[602]  ( .D(n14775), .CLK(clk), .RST(rst), .Q(ereg[602]) );
  DFF \ereg_reg[603]  ( .D(n14774), .CLK(clk), .RST(rst), .Q(ereg[603]) );
  DFF \ereg_reg[604]  ( .D(n14773), .CLK(clk), .RST(rst), .Q(ereg[604]) );
  DFF \ereg_reg[605]  ( .D(n14772), .CLK(clk), .RST(rst), .Q(ereg[605]) );
  DFF \ereg_reg[606]  ( .D(n14771), .CLK(clk), .RST(rst), .Q(ereg[606]) );
  DFF \ereg_reg[607]  ( .D(n14770), .CLK(clk), .RST(rst), .Q(ereg[607]) );
  DFF \ereg_reg[608]  ( .D(n14769), .CLK(clk), .RST(rst), .Q(ereg[608]) );
  DFF \ereg_reg[609]  ( .D(n14768), .CLK(clk), .RST(rst), .Q(ereg[609]) );
  DFF \ereg_reg[610]  ( .D(n14767), .CLK(clk), .RST(rst), .Q(ereg[610]) );
  DFF \ereg_reg[611]  ( .D(n14766), .CLK(clk), .RST(rst), .Q(ereg[611]) );
  DFF \ereg_reg[612]  ( .D(n14765), .CLK(clk), .RST(rst), .Q(ereg[612]) );
  DFF \ereg_reg[613]  ( .D(n14764), .CLK(clk), .RST(rst), .Q(ereg[613]) );
  DFF \ereg_reg[614]  ( .D(n14763), .CLK(clk), .RST(rst), .Q(ereg[614]) );
  DFF \ereg_reg[615]  ( .D(n14762), .CLK(clk), .RST(rst), .Q(ereg[615]) );
  DFF \ereg_reg[616]  ( .D(n14761), .CLK(clk), .RST(rst), .Q(ereg[616]) );
  DFF \ereg_reg[617]  ( .D(n14760), .CLK(clk), .RST(rst), .Q(ereg[617]) );
  DFF \ereg_reg[618]  ( .D(n14759), .CLK(clk), .RST(rst), .Q(ereg[618]) );
  DFF \ereg_reg[619]  ( .D(n14758), .CLK(clk), .RST(rst), .Q(ereg[619]) );
  DFF \ereg_reg[620]  ( .D(n14757), .CLK(clk), .RST(rst), .Q(ereg[620]) );
  DFF \ereg_reg[621]  ( .D(n14756), .CLK(clk), .RST(rst), .Q(ereg[621]) );
  DFF \ereg_reg[622]  ( .D(n14755), .CLK(clk), .RST(rst), .Q(ereg[622]) );
  DFF \ereg_reg[623]  ( .D(n14754), .CLK(clk), .RST(rst), .Q(ereg[623]) );
  DFF \ereg_reg[624]  ( .D(n14753), .CLK(clk), .RST(rst), .Q(ereg[624]) );
  DFF \ereg_reg[625]  ( .D(n14752), .CLK(clk), .RST(rst), .Q(ereg[625]) );
  DFF \ereg_reg[626]  ( .D(n14751), .CLK(clk), .RST(rst), .Q(ereg[626]) );
  DFF \ereg_reg[627]  ( .D(n14750), .CLK(clk), .RST(rst), .Q(ereg[627]) );
  DFF \ereg_reg[628]  ( .D(n14749), .CLK(clk), .RST(rst), .Q(ereg[628]) );
  DFF \ereg_reg[629]  ( .D(n14748), .CLK(clk), .RST(rst), .Q(ereg[629]) );
  DFF \ereg_reg[630]  ( .D(n14747), .CLK(clk), .RST(rst), .Q(ereg[630]) );
  DFF \ereg_reg[631]  ( .D(n14746), .CLK(clk), .RST(rst), .Q(ereg[631]) );
  DFF \ereg_reg[632]  ( .D(n14745), .CLK(clk), .RST(rst), .Q(ereg[632]) );
  DFF \ereg_reg[633]  ( .D(n14744), .CLK(clk), .RST(rst), .Q(ereg[633]) );
  DFF \ereg_reg[634]  ( .D(n14743), .CLK(clk), .RST(rst), .Q(ereg[634]) );
  DFF \ereg_reg[635]  ( .D(n14742), .CLK(clk), .RST(rst), .Q(ereg[635]) );
  DFF \ereg_reg[636]  ( .D(n14741), .CLK(clk), .RST(rst), .Q(ereg[636]) );
  DFF \ereg_reg[637]  ( .D(n14740), .CLK(clk), .RST(rst), .Q(ereg[637]) );
  DFF \ereg_reg[638]  ( .D(n14739), .CLK(clk), .RST(rst), .Q(ereg[638]) );
  DFF \ereg_reg[639]  ( .D(n14738), .CLK(clk), .RST(rst), .Q(ereg[639]) );
  DFF \ereg_reg[640]  ( .D(n14737), .CLK(clk), .RST(rst), .Q(ereg[640]) );
  DFF \ereg_reg[641]  ( .D(n14736), .CLK(clk), .RST(rst), .Q(ereg[641]) );
  DFF \ereg_reg[642]  ( .D(n14735), .CLK(clk), .RST(rst), .Q(ereg[642]) );
  DFF \ereg_reg[643]  ( .D(n14734), .CLK(clk), .RST(rst), .Q(ereg[643]) );
  DFF \ereg_reg[644]  ( .D(n14733), .CLK(clk), .RST(rst), .Q(ereg[644]) );
  DFF \ereg_reg[645]  ( .D(n14732), .CLK(clk), .RST(rst), .Q(ereg[645]) );
  DFF \ereg_reg[646]  ( .D(n14731), .CLK(clk), .RST(rst), .Q(ereg[646]) );
  DFF \ereg_reg[647]  ( .D(n14730), .CLK(clk), .RST(rst), .Q(ereg[647]) );
  DFF \ereg_reg[648]  ( .D(n14729), .CLK(clk), .RST(rst), .Q(ereg[648]) );
  DFF \ereg_reg[649]  ( .D(n14728), .CLK(clk), .RST(rst), .Q(ereg[649]) );
  DFF \ereg_reg[650]  ( .D(n14727), .CLK(clk), .RST(rst), .Q(ereg[650]) );
  DFF \ereg_reg[651]  ( .D(n14726), .CLK(clk), .RST(rst), .Q(ereg[651]) );
  DFF \ereg_reg[652]  ( .D(n14725), .CLK(clk), .RST(rst), .Q(ereg[652]) );
  DFF \ereg_reg[653]  ( .D(n14724), .CLK(clk), .RST(rst), .Q(ereg[653]) );
  DFF \ereg_reg[654]  ( .D(n14723), .CLK(clk), .RST(rst), .Q(ereg[654]) );
  DFF \ereg_reg[655]  ( .D(n14722), .CLK(clk), .RST(rst), .Q(ereg[655]) );
  DFF \ereg_reg[656]  ( .D(n14721), .CLK(clk), .RST(rst), .Q(ereg[656]) );
  DFF \ereg_reg[657]  ( .D(n14720), .CLK(clk), .RST(rst), .Q(ereg[657]) );
  DFF \ereg_reg[658]  ( .D(n14719), .CLK(clk), .RST(rst), .Q(ereg[658]) );
  DFF \ereg_reg[659]  ( .D(n14718), .CLK(clk), .RST(rst), .Q(ereg[659]) );
  DFF \ereg_reg[660]  ( .D(n14717), .CLK(clk), .RST(rst), .Q(ereg[660]) );
  DFF \ereg_reg[661]  ( .D(n14716), .CLK(clk), .RST(rst), .Q(ereg[661]) );
  DFF \ereg_reg[662]  ( .D(n14715), .CLK(clk), .RST(rst), .Q(ereg[662]) );
  DFF \ereg_reg[663]  ( .D(n14714), .CLK(clk), .RST(rst), .Q(ereg[663]) );
  DFF \ereg_reg[664]  ( .D(n14713), .CLK(clk), .RST(rst), .Q(ereg[664]) );
  DFF \ereg_reg[665]  ( .D(n14712), .CLK(clk), .RST(rst), .Q(ereg[665]) );
  DFF \ereg_reg[666]  ( .D(n14711), .CLK(clk), .RST(rst), .Q(ereg[666]) );
  DFF \ereg_reg[667]  ( .D(n14710), .CLK(clk), .RST(rst), .Q(ereg[667]) );
  DFF \ereg_reg[668]  ( .D(n14709), .CLK(clk), .RST(rst), .Q(ereg[668]) );
  DFF \ereg_reg[669]  ( .D(n14708), .CLK(clk), .RST(rst), .Q(ereg[669]) );
  DFF \ereg_reg[670]  ( .D(n14707), .CLK(clk), .RST(rst), .Q(ereg[670]) );
  DFF \ereg_reg[671]  ( .D(n14706), .CLK(clk), .RST(rst), .Q(ereg[671]) );
  DFF \ereg_reg[672]  ( .D(n14705), .CLK(clk), .RST(rst), .Q(ereg[672]) );
  DFF \ereg_reg[673]  ( .D(n14704), .CLK(clk), .RST(rst), .Q(ereg[673]) );
  DFF \ereg_reg[674]  ( .D(n14703), .CLK(clk), .RST(rst), .Q(ereg[674]) );
  DFF \ereg_reg[675]  ( .D(n14702), .CLK(clk), .RST(rst), .Q(ereg[675]) );
  DFF \ereg_reg[676]  ( .D(n14701), .CLK(clk), .RST(rst), .Q(ereg[676]) );
  DFF \ereg_reg[677]  ( .D(n14700), .CLK(clk), .RST(rst), .Q(ereg[677]) );
  DFF \ereg_reg[678]  ( .D(n14699), .CLK(clk), .RST(rst), .Q(ereg[678]) );
  DFF \ereg_reg[679]  ( .D(n14698), .CLK(clk), .RST(rst), .Q(ereg[679]) );
  DFF \ereg_reg[680]  ( .D(n14697), .CLK(clk), .RST(rst), .Q(ereg[680]) );
  DFF \ereg_reg[681]  ( .D(n14696), .CLK(clk), .RST(rst), .Q(ereg[681]) );
  DFF \ereg_reg[682]  ( .D(n14695), .CLK(clk), .RST(rst), .Q(ereg[682]) );
  DFF \ereg_reg[683]  ( .D(n14694), .CLK(clk), .RST(rst), .Q(ereg[683]) );
  DFF \ereg_reg[684]  ( .D(n14693), .CLK(clk), .RST(rst), .Q(ereg[684]) );
  DFF \ereg_reg[685]  ( .D(n14692), .CLK(clk), .RST(rst), .Q(ereg[685]) );
  DFF \ereg_reg[686]  ( .D(n14691), .CLK(clk), .RST(rst), .Q(ereg[686]) );
  DFF \ereg_reg[687]  ( .D(n14690), .CLK(clk), .RST(rst), .Q(ereg[687]) );
  DFF \ereg_reg[688]  ( .D(n14689), .CLK(clk), .RST(rst), .Q(ereg[688]) );
  DFF \ereg_reg[689]  ( .D(n14688), .CLK(clk), .RST(rst), .Q(ereg[689]) );
  DFF \ereg_reg[690]  ( .D(n14687), .CLK(clk), .RST(rst), .Q(ereg[690]) );
  DFF \ereg_reg[691]  ( .D(n14686), .CLK(clk), .RST(rst), .Q(ereg[691]) );
  DFF \ereg_reg[692]  ( .D(n14685), .CLK(clk), .RST(rst), .Q(ereg[692]) );
  DFF \ereg_reg[693]  ( .D(n14684), .CLK(clk), .RST(rst), .Q(ereg[693]) );
  DFF \ereg_reg[694]  ( .D(n14683), .CLK(clk), .RST(rst), .Q(ereg[694]) );
  DFF \ereg_reg[695]  ( .D(n14682), .CLK(clk), .RST(rst), .Q(ereg[695]) );
  DFF \ereg_reg[696]  ( .D(n14681), .CLK(clk), .RST(rst), .Q(ereg[696]) );
  DFF \ereg_reg[697]  ( .D(n14680), .CLK(clk), .RST(rst), .Q(ereg[697]) );
  DFF \ereg_reg[698]  ( .D(n14679), .CLK(clk), .RST(rst), .Q(ereg[698]) );
  DFF \ereg_reg[699]  ( .D(n14678), .CLK(clk), .RST(rst), .Q(ereg[699]) );
  DFF \ereg_reg[700]  ( .D(n14677), .CLK(clk), .RST(rst), .Q(ereg[700]) );
  DFF \ereg_reg[701]  ( .D(n14676), .CLK(clk), .RST(rst), .Q(ereg[701]) );
  DFF \ereg_reg[702]  ( .D(n14675), .CLK(clk), .RST(rst), .Q(ereg[702]) );
  DFF \ereg_reg[703]  ( .D(n14674), .CLK(clk), .RST(rst), .Q(ereg[703]) );
  DFF \ereg_reg[704]  ( .D(n14673), .CLK(clk), .RST(rst), .Q(ereg[704]) );
  DFF \ereg_reg[705]  ( .D(n14672), .CLK(clk), .RST(rst), .Q(ereg[705]) );
  DFF \ereg_reg[706]  ( .D(n14671), .CLK(clk), .RST(rst), .Q(ereg[706]) );
  DFF \ereg_reg[707]  ( .D(n14670), .CLK(clk), .RST(rst), .Q(ereg[707]) );
  DFF \ereg_reg[708]  ( .D(n14669), .CLK(clk), .RST(rst), .Q(ereg[708]) );
  DFF \ereg_reg[709]  ( .D(n14668), .CLK(clk), .RST(rst), .Q(ereg[709]) );
  DFF \ereg_reg[710]  ( .D(n14667), .CLK(clk), .RST(rst), .Q(ereg[710]) );
  DFF \ereg_reg[711]  ( .D(n14666), .CLK(clk), .RST(rst), .Q(ereg[711]) );
  DFF \ereg_reg[712]  ( .D(n14665), .CLK(clk), .RST(rst), .Q(ereg[712]) );
  DFF \ereg_reg[713]  ( .D(n14664), .CLK(clk), .RST(rst), .Q(ereg[713]) );
  DFF \ereg_reg[714]  ( .D(n14663), .CLK(clk), .RST(rst), .Q(ereg[714]) );
  DFF \ereg_reg[715]  ( .D(n14662), .CLK(clk), .RST(rst), .Q(ereg[715]) );
  DFF \ereg_reg[716]  ( .D(n14661), .CLK(clk), .RST(rst), .Q(ereg[716]) );
  DFF \ereg_reg[717]  ( .D(n14660), .CLK(clk), .RST(rst), .Q(ereg[717]) );
  DFF \ereg_reg[718]  ( .D(n14659), .CLK(clk), .RST(rst), .Q(ereg[718]) );
  DFF \ereg_reg[719]  ( .D(n14658), .CLK(clk), .RST(rst), .Q(ereg[719]) );
  DFF \ereg_reg[720]  ( .D(n14657), .CLK(clk), .RST(rst), .Q(ereg[720]) );
  DFF \ereg_reg[721]  ( .D(n14656), .CLK(clk), .RST(rst), .Q(ereg[721]) );
  DFF \ereg_reg[722]  ( .D(n14655), .CLK(clk), .RST(rst), .Q(ereg[722]) );
  DFF \ereg_reg[723]  ( .D(n14654), .CLK(clk), .RST(rst), .Q(ereg[723]) );
  DFF \ereg_reg[724]  ( .D(n14653), .CLK(clk), .RST(rst), .Q(ereg[724]) );
  DFF \ereg_reg[725]  ( .D(n14652), .CLK(clk), .RST(rst), .Q(ereg[725]) );
  DFF \ereg_reg[726]  ( .D(n14651), .CLK(clk), .RST(rst), .Q(ereg[726]) );
  DFF \ereg_reg[727]  ( .D(n14650), .CLK(clk), .RST(rst), .Q(ereg[727]) );
  DFF \ereg_reg[728]  ( .D(n14649), .CLK(clk), .RST(rst), .Q(ereg[728]) );
  DFF \ereg_reg[729]  ( .D(n14648), .CLK(clk), .RST(rst), .Q(ereg[729]) );
  DFF \ereg_reg[730]  ( .D(n14647), .CLK(clk), .RST(rst), .Q(ereg[730]) );
  DFF \ereg_reg[731]  ( .D(n14646), .CLK(clk), .RST(rst), .Q(ereg[731]) );
  DFF \ereg_reg[732]  ( .D(n14645), .CLK(clk), .RST(rst), .Q(ereg[732]) );
  DFF \ereg_reg[733]  ( .D(n14644), .CLK(clk), .RST(rst), .Q(ereg[733]) );
  DFF \ereg_reg[734]  ( .D(n14643), .CLK(clk), .RST(rst), .Q(ereg[734]) );
  DFF \ereg_reg[735]  ( .D(n14642), .CLK(clk), .RST(rst), .Q(ereg[735]) );
  DFF \ereg_reg[736]  ( .D(n14641), .CLK(clk), .RST(rst), .Q(ereg[736]) );
  DFF \ereg_reg[737]  ( .D(n14640), .CLK(clk), .RST(rst), .Q(ereg[737]) );
  DFF \ereg_reg[738]  ( .D(n14639), .CLK(clk), .RST(rst), .Q(ereg[738]) );
  DFF \ereg_reg[739]  ( .D(n14638), .CLK(clk), .RST(rst), .Q(ereg[739]) );
  DFF \ereg_reg[740]  ( .D(n14637), .CLK(clk), .RST(rst), .Q(ereg[740]) );
  DFF \ereg_reg[741]  ( .D(n14636), .CLK(clk), .RST(rst), .Q(ereg[741]) );
  DFF \ereg_reg[742]  ( .D(n14635), .CLK(clk), .RST(rst), .Q(ereg[742]) );
  DFF \ereg_reg[743]  ( .D(n14634), .CLK(clk), .RST(rst), .Q(ereg[743]) );
  DFF \ereg_reg[744]  ( .D(n14633), .CLK(clk), .RST(rst), .Q(ereg[744]) );
  DFF \ereg_reg[745]  ( .D(n14632), .CLK(clk), .RST(rst), .Q(ereg[745]) );
  DFF \ereg_reg[746]  ( .D(n14631), .CLK(clk), .RST(rst), .Q(ereg[746]) );
  DFF \ereg_reg[747]  ( .D(n14630), .CLK(clk), .RST(rst), .Q(ereg[747]) );
  DFF \ereg_reg[748]  ( .D(n14629), .CLK(clk), .RST(rst), .Q(ereg[748]) );
  DFF \ereg_reg[749]  ( .D(n14628), .CLK(clk), .RST(rst), .Q(ereg[749]) );
  DFF \ereg_reg[750]  ( .D(n14627), .CLK(clk), .RST(rst), .Q(ereg[750]) );
  DFF \ereg_reg[751]  ( .D(n14626), .CLK(clk), .RST(rst), .Q(ereg[751]) );
  DFF \ereg_reg[752]  ( .D(n14625), .CLK(clk), .RST(rst), .Q(ereg[752]) );
  DFF \ereg_reg[753]  ( .D(n14624), .CLK(clk), .RST(rst), .Q(ereg[753]) );
  DFF \ereg_reg[754]  ( .D(n14623), .CLK(clk), .RST(rst), .Q(ereg[754]) );
  DFF \ereg_reg[755]  ( .D(n14622), .CLK(clk), .RST(rst), .Q(ereg[755]) );
  DFF \ereg_reg[756]  ( .D(n14621), .CLK(clk), .RST(rst), .Q(ereg[756]) );
  DFF \ereg_reg[757]  ( .D(n14620), .CLK(clk), .RST(rst), .Q(ereg[757]) );
  DFF \ereg_reg[758]  ( .D(n14619), .CLK(clk), .RST(rst), .Q(ereg[758]) );
  DFF \ereg_reg[759]  ( .D(n14618), .CLK(clk), .RST(rst), .Q(ereg[759]) );
  DFF \ereg_reg[760]  ( .D(n14617), .CLK(clk), .RST(rst), .Q(ereg[760]) );
  DFF \ereg_reg[761]  ( .D(n14616), .CLK(clk), .RST(rst), .Q(ereg[761]) );
  DFF \ereg_reg[762]  ( .D(n14615), .CLK(clk), .RST(rst), .Q(ereg[762]) );
  DFF \ereg_reg[763]  ( .D(n14614), .CLK(clk), .RST(rst), .Q(ereg[763]) );
  DFF \ereg_reg[764]  ( .D(n14613), .CLK(clk), .RST(rst), .Q(ereg[764]) );
  DFF \ereg_reg[765]  ( .D(n14612), .CLK(clk), .RST(rst), .Q(ereg[765]) );
  DFF \ereg_reg[766]  ( .D(n14611), .CLK(clk), .RST(rst), .Q(ereg[766]) );
  DFF \ereg_reg[767]  ( .D(n14610), .CLK(clk), .RST(rst), .Q(ereg[767]) );
  DFF \ereg_reg[768]  ( .D(n14609), .CLK(clk), .RST(rst), .Q(ereg[768]) );
  DFF \ereg_reg[769]  ( .D(n14608), .CLK(clk), .RST(rst), .Q(ereg[769]) );
  DFF \ereg_reg[770]  ( .D(n14607), .CLK(clk), .RST(rst), .Q(ereg[770]) );
  DFF \ereg_reg[771]  ( .D(n14606), .CLK(clk), .RST(rst), .Q(ereg[771]) );
  DFF \ereg_reg[772]  ( .D(n14605), .CLK(clk), .RST(rst), .Q(ereg[772]) );
  DFF \ereg_reg[773]  ( .D(n14604), .CLK(clk), .RST(rst), .Q(ereg[773]) );
  DFF \ereg_reg[774]  ( .D(n14603), .CLK(clk), .RST(rst), .Q(ereg[774]) );
  DFF \ereg_reg[775]  ( .D(n14602), .CLK(clk), .RST(rst), .Q(ereg[775]) );
  DFF \ereg_reg[776]  ( .D(n14601), .CLK(clk), .RST(rst), .Q(ereg[776]) );
  DFF \ereg_reg[777]  ( .D(n14600), .CLK(clk), .RST(rst), .Q(ereg[777]) );
  DFF \ereg_reg[778]  ( .D(n14599), .CLK(clk), .RST(rst), .Q(ereg[778]) );
  DFF \ereg_reg[779]  ( .D(n14598), .CLK(clk), .RST(rst), .Q(ereg[779]) );
  DFF \ereg_reg[780]  ( .D(n14597), .CLK(clk), .RST(rst), .Q(ereg[780]) );
  DFF \ereg_reg[781]  ( .D(n14596), .CLK(clk), .RST(rst), .Q(ereg[781]) );
  DFF \ereg_reg[782]  ( .D(n14595), .CLK(clk), .RST(rst), .Q(ereg[782]) );
  DFF \ereg_reg[783]  ( .D(n14594), .CLK(clk), .RST(rst), .Q(ereg[783]) );
  DFF \ereg_reg[784]  ( .D(n14593), .CLK(clk), .RST(rst), .Q(ereg[784]) );
  DFF \ereg_reg[785]  ( .D(n14592), .CLK(clk), .RST(rst), .Q(ereg[785]) );
  DFF \ereg_reg[786]  ( .D(n14591), .CLK(clk), .RST(rst), .Q(ereg[786]) );
  DFF \ereg_reg[787]  ( .D(n14590), .CLK(clk), .RST(rst), .Q(ereg[787]) );
  DFF \ereg_reg[788]  ( .D(n14589), .CLK(clk), .RST(rst), .Q(ereg[788]) );
  DFF \ereg_reg[789]  ( .D(n14588), .CLK(clk), .RST(rst), .Q(ereg[789]) );
  DFF \ereg_reg[790]  ( .D(n14587), .CLK(clk), .RST(rst), .Q(ereg[790]) );
  DFF \ereg_reg[791]  ( .D(n14586), .CLK(clk), .RST(rst), .Q(ereg[791]) );
  DFF \ereg_reg[792]  ( .D(n14585), .CLK(clk), .RST(rst), .Q(ereg[792]) );
  DFF \ereg_reg[793]  ( .D(n14584), .CLK(clk), .RST(rst), .Q(ereg[793]) );
  DFF \ereg_reg[794]  ( .D(n14583), .CLK(clk), .RST(rst), .Q(ereg[794]) );
  DFF \ereg_reg[795]  ( .D(n14582), .CLK(clk), .RST(rst), .Q(ereg[795]) );
  DFF \ereg_reg[796]  ( .D(n14581), .CLK(clk), .RST(rst), .Q(ereg[796]) );
  DFF \ereg_reg[797]  ( .D(n14580), .CLK(clk), .RST(rst), .Q(ereg[797]) );
  DFF \ereg_reg[798]  ( .D(n14579), .CLK(clk), .RST(rst), .Q(ereg[798]) );
  DFF \ereg_reg[799]  ( .D(n14578), .CLK(clk), .RST(rst), .Q(ereg[799]) );
  DFF \ereg_reg[800]  ( .D(n14577), .CLK(clk), .RST(rst), .Q(ereg[800]) );
  DFF \ereg_reg[801]  ( .D(n14576), .CLK(clk), .RST(rst), .Q(ereg[801]) );
  DFF \ereg_reg[802]  ( .D(n14575), .CLK(clk), .RST(rst), .Q(ereg[802]) );
  DFF \ereg_reg[803]  ( .D(n14574), .CLK(clk), .RST(rst), .Q(ereg[803]) );
  DFF \ereg_reg[804]  ( .D(n14573), .CLK(clk), .RST(rst), .Q(ereg[804]) );
  DFF \ereg_reg[805]  ( .D(n14572), .CLK(clk), .RST(rst), .Q(ereg[805]) );
  DFF \ereg_reg[806]  ( .D(n14571), .CLK(clk), .RST(rst), .Q(ereg[806]) );
  DFF \ereg_reg[807]  ( .D(n14570), .CLK(clk), .RST(rst), .Q(ereg[807]) );
  DFF \ereg_reg[808]  ( .D(n14569), .CLK(clk), .RST(rst), .Q(ereg[808]) );
  DFF \ereg_reg[809]  ( .D(n14568), .CLK(clk), .RST(rst), .Q(ereg[809]) );
  DFF \ereg_reg[810]  ( .D(n14567), .CLK(clk), .RST(rst), .Q(ereg[810]) );
  DFF \ereg_reg[811]  ( .D(n14566), .CLK(clk), .RST(rst), .Q(ereg[811]) );
  DFF \ereg_reg[812]  ( .D(n14565), .CLK(clk), .RST(rst), .Q(ereg[812]) );
  DFF \ereg_reg[813]  ( .D(n14564), .CLK(clk), .RST(rst), .Q(ereg[813]) );
  DFF \ereg_reg[814]  ( .D(n14563), .CLK(clk), .RST(rst), .Q(ereg[814]) );
  DFF \ereg_reg[815]  ( .D(n14562), .CLK(clk), .RST(rst), .Q(ereg[815]) );
  DFF \ereg_reg[816]  ( .D(n14561), .CLK(clk), .RST(rst), .Q(ereg[816]) );
  DFF \ereg_reg[817]  ( .D(n14560), .CLK(clk), .RST(rst), .Q(ereg[817]) );
  DFF \ereg_reg[818]  ( .D(n14559), .CLK(clk), .RST(rst), .Q(ereg[818]) );
  DFF \ereg_reg[819]  ( .D(n14558), .CLK(clk), .RST(rst), .Q(ereg[819]) );
  DFF \ereg_reg[820]  ( .D(n14557), .CLK(clk), .RST(rst), .Q(ereg[820]) );
  DFF \ereg_reg[821]  ( .D(n14556), .CLK(clk), .RST(rst), .Q(ereg[821]) );
  DFF \ereg_reg[822]  ( .D(n14555), .CLK(clk), .RST(rst), .Q(ereg[822]) );
  DFF \ereg_reg[823]  ( .D(n14554), .CLK(clk), .RST(rst), .Q(ereg[823]) );
  DFF \ereg_reg[824]  ( .D(n14553), .CLK(clk), .RST(rst), .Q(ereg[824]) );
  DFF \ereg_reg[825]  ( .D(n14552), .CLK(clk), .RST(rst), .Q(ereg[825]) );
  DFF \ereg_reg[826]  ( .D(n14551), .CLK(clk), .RST(rst), .Q(ereg[826]) );
  DFF \ereg_reg[827]  ( .D(n14550), .CLK(clk), .RST(rst), .Q(ereg[827]) );
  DFF \ereg_reg[828]  ( .D(n14549), .CLK(clk), .RST(rst), .Q(ereg[828]) );
  DFF \ereg_reg[829]  ( .D(n14548), .CLK(clk), .RST(rst), .Q(ereg[829]) );
  DFF \ereg_reg[830]  ( .D(n14547), .CLK(clk), .RST(rst), .Q(ereg[830]) );
  DFF \ereg_reg[831]  ( .D(n14546), .CLK(clk), .RST(rst), .Q(ereg[831]) );
  DFF \ereg_reg[832]  ( .D(n14545), .CLK(clk), .RST(rst), .Q(ereg[832]) );
  DFF \ereg_reg[833]  ( .D(n14544), .CLK(clk), .RST(rst), .Q(ereg[833]) );
  DFF \ereg_reg[834]  ( .D(n14543), .CLK(clk), .RST(rst), .Q(ereg[834]) );
  DFF \ereg_reg[835]  ( .D(n14542), .CLK(clk), .RST(rst), .Q(ereg[835]) );
  DFF \ereg_reg[836]  ( .D(n14541), .CLK(clk), .RST(rst), .Q(ereg[836]) );
  DFF \ereg_reg[837]  ( .D(n14540), .CLK(clk), .RST(rst), .Q(ereg[837]) );
  DFF \ereg_reg[838]  ( .D(n14539), .CLK(clk), .RST(rst), .Q(ereg[838]) );
  DFF \ereg_reg[839]  ( .D(n14538), .CLK(clk), .RST(rst), .Q(ereg[839]) );
  DFF \ereg_reg[840]  ( .D(n14537), .CLK(clk), .RST(rst), .Q(ereg[840]) );
  DFF \ereg_reg[841]  ( .D(n14536), .CLK(clk), .RST(rst), .Q(ereg[841]) );
  DFF \ereg_reg[842]  ( .D(n14535), .CLK(clk), .RST(rst), .Q(ereg[842]) );
  DFF \ereg_reg[843]  ( .D(n14534), .CLK(clk), .RST(rst), .Q(ereg[843]) );
  DFF \ereg_reg[844]  ( .D(n14533), .CLK(clk), .RST(rst), .Q(ereg[844]) );
  DFF \ereg_reg[845]  ( .D(n14532), .CLK(clk), .RST(rst), .Q(ereg[845]) );
  DFF \ereg_reg[846]  ( .D(n14531), .CLK(clk), .RST(rst), .Q(ereg[846]) );
  DFF \ereg_reg[847]  ( .D(n14530), .CLK(clk), .RST(rst), .Q(ereg[847]) );
  DFF \ereg_reg[848]  ( .D(n14529), .CLK(clk), .RST(rst), .Q(ereg[848]) );
  DFF \ereg_reg[849]  ( .D(n14528), .CLK(clk), .RST(rst), .Q(ereg[849]) );
  DFF \ereg_reg[850]  ( .D(n14527), .CLK(clk), .RST(rst), .Q(ereg[850]) );
  DFF \ereg_reg[851]  ( .D(n14526), .CLK(clk), .RST(rst), .Q(ereg[851]) );
  DFF \ereg_reg[852]  ( .D(n14525), .CLK(clk), .RST(rst), .Q(ereg[852]) );
  DFF \ereg_reg[853]  ( .D(n14524), .CLK(clk), .RST(rst), .Q(ereg[853]) );
  DFF \ereg_reg[854]  ( .D(n14523), .CLK(clk), .RST(rst), .Q(ereg[854]) );
  DFF \ereg_reg[855]  ( .D(n14522), .CLK(clk), .RST(rst), .Q(ereg[855]) );
  DFF \ereg_reg[856]  ( .D(n14521), .CLK(clk), .RST(rst), .Q(ereg[856]) );
  DFF \ereg_reg[857]  ( .D(n14520), .CLK(clk), .RST(rst), .Q(ereg[857]) );
  DFF \ereg_reg[858]  ( .D(n14519), .CLK(clk), .RST(rst), .Q(ereg[858]) );
  DFF \ereg_reg[859]  ( .D(n14518), .CLK(clk), .RST(rst), .Q(ereg[859]) );
  DFF \ereg_reg[860]  ( .D(n14517), .CLK(clk), .RST(rst), .Q(ereg[860]) );
  DFF \ereg_reg[861]  ( .D(n14516), .CLK(clk), .RST(rst), .Q(ereg[861]) );
  DFF \ereg_reg[862]  ( .D(n14515), .CLK(clk), .RST(rst), .Q(ereg[862]) );
  DFF \ereg_reg[863]  ( .D(n14514), .CLK(clk), .RST(rst), .Q(ereg[863]) );
  DFF \ereg_reg[864]  ( .D(n14513), .CLK(clk), .RST(rst), .Q(ereg[864]) );
  DFF \ereg_reg[865]  ( .D(n14512), .CLK(clk), .RST(rst), .Q(ereg[865]) );
  DFF \ereg_reg[866]  ( .D(n14511), .CLK(clk), .RST(rst), .Q(ereg[866]) );
  DFF \ereg_reg[867]  ( .D(n14510), .CLK(clk), .RST(rst), .Q(ereg[867]) );
  DFF \ereg_reg[868]  ( .D(n14509), .CLK(clk), .RST(rst), .Q(ereg[868]) );
  DFF \ereg_reg[869]  ( .D(n14508), .CLK(clk), .RST(rst), .Q(ereg[869]) );
  DFF \ereg_reg[870]  ( .D(n14507), .CLK(clk), .RST(rst), .Q(ereg[870]) );
  DFF \ereg_reg[871]  ( .D(n14506), .CLK(clk), .RST(rst), .Q(ereg[871]) );
  DFF \ereg_reg[872]  ( .D(n14505), .CLK(clk), .RST(rst), .Q(ereg[872]) );
  DFF \ereg_reg[873]  ( .D(n14504), .CLK(clk), .RST(rst), .Q(ereg[873]) );
  DFF \ereg_reg[874]  ( .D(n14503), .CLK(clk), .RST(rst), .Q(ereg[874]) );
  DFF \ereg_reg[875]  ( .D(n14502), .CLK(clk), .RST(rst), .Q(ereg[875]) );
  DFF \ereg_reg[876]  ( .D(n14501), .CLK(clk), .RST(rst), .Q(ereg[876]) );
  DFF \ereg_reg[877]  ( .D(n14500), .CLK(clk), .RST(rst), .Q(ereg[877]) );
  DFF \ereg_reg[878]  ( .D(n14499), .CLK(clk), .RST(rst), .Q(ereg[878]) );
  DFF \ereg_reg[879]  ( .D(n14498), .CLK(clk), .RST(rst), .Q(ereg[879]) );
  DFF \ereg_reg[880]  ( .D(n14497), .CLK(clk), .RST(rst), .Q(ereg[880]) );
  DFF \ereg_reg[881]  ( .D(n14496), .CLK(clk), .RST(rst), .Q(ereg[881]) );
  DFF \ereg_reg[882]  ( .D(n14495), .CLK(clk), .RST(rst), .Q(ereg[882]) );
  DFF \ereg_reg[883]  ( .D(n14494), .CLK(clk), .RST(rst), .Q(ereg[883]) );
  DFF \ereg_reg[884]  ( .D(n14493), .CLK(clk), .RST(rst), .Q(ereg[884]) );
  DFF \ereg_reg[885]  ( .D(n14492), .CLK(clk), .RST(rst), .Q(ereg[885]) );
  DFF \ereg_reg[886]  ( .D(n14491), .CLK(clk), .RST(rst), .Q(ereg[886]) );
  DFF \ereg_reg[887]  ( .D(n14490), .CLK(clk), .RST(rst), .Q(ereg[887]) );
  DFF \ereg_reg[888]  ( .D(n14489), .CLK(clk), .RST(rst), .Q(ereg[888]) );
  DFF \ereg_reg[889]  ( .D(n14488), .CLK(clk), .RST(rst), .Q(ereg[889]) );
  DFF \ereg_reg[890]  ( .D(n14487), .CLK(clk), .RST(rst), .Q(ereg[890]) );
  DFF \ereg_reg[891]  ( .D(n14486), .CLK(clk), .RST(rst), .Q(ereg[891]) );
  DFF \ereg_reg[892]  ( .D(n14485), .CLK(clk), .RST(rst), .Q(ereg[892]) );
  DFF \ereg_reg[893]  ( .D(n14484), .CLK(clk), .RST(rst), .Q(ereg[893]) );
  DFF \ereg_reg[894]  ( .D(n14483), .CLK(clk), .RST(rst), .Q(ereg[894]) );
  DFF \ereg_reg[895]  ( .D(n14482), .CLK(clk), .RST(rst), .Q(ereg[895]) );
  DFF \ereg_reg[896]  ( .D(n14481), .CLK(clk), .RST(rst), .Q(ereg[896]) );
  DFF \ereg_reg[897]  ( .D(n14480), .CLK(clk), .RST(rst), .Q(ereg[897]) );
  DFF \ereg_reg[898]  ( .D(n14479), .CLK(clk), .RST(rst), .Q(ereg[898]) );
  DFF \ereg_reg[899]  ( .D(n14478), .CLK(clk), .RST(rst), .Q(ereg[899]) );
  DFF \ereg_reg[900]  ( .D(n14477), .CLK(clk), .RST(rst), .Q(ereg[900]) );
  DFF \ereg_reg[901]  ( .D(n14476), .CLK(clk), .RST(rst), .Q(ereg[901]) );
  DFF \ereg_reg[902]  ( .D(n14475), .CLK(clk), .RST(rst), .Q(ereg[902]) );
  DFF \ereg_reg[903]  ( .D(n14474), .CLK(clk), .RST(rst), .Q(ereg[903]) );
  DFF \ereg_reg[904]  ( .D(n14473), .CLK(clk), .RST(rst), .Q(ereg[904]) );
  DFF \ereg_reg[905]  ( .D(n14472), .CLK(clk), .RST(rst), .Q(ereg[905]) );
  DFF \ereg_reg[906]  ( .D(n14471), .CLK(clk), .RST(rst), .Q(ereg[906]) );
  DFF \ereg_reg[907]  ( .D(n14470), .CLK(clk), .RST(rst), .Q(ereg[907]) );
  DFF \ereg_reg[908]  ( .D(n14469), .CLK(clk), .RST(rst), .Q(ereg[908]) );
  DFF \ereg_reg[909]  ( .D(n14468), .CLK(clk), .RST(rst), .Q(ereg[909]) );
  DFF \ereg_reg[910]  ( .D(n14467), .CLK(clk), .RST(rst), .Q(ereg[910]) );
  DFF \ereg_reg[911]  ( .D(n14466), .CLK(clk), .RST(rst), .Q(ereg[911]) );
  DFF \ereg_reg[912]  ( .D(n14465), .CLK(clk), .RST(rst), .Q(ereg[912]) );
  DFF \ereg_reg[913]  ( .D(n14464), .CLK(clk), .RST(rst), .Q(ereg[913]) );
  DFF \ereg_reg[914]  ( .D(n14463), .CLK(clk), .RST(rst), .Q(ereg[914]) );
  DFF \ereg_reg[915]  ( .D(n14462), .CLK(clk), .RST(rst), .Q(ereg[915]) );
  DFF \ereg_reg[916]  ( .D(n14461), .CLK(clk), .RST(rst), .Q(ereg[916]) );
  DFF \ereg_reg[917]  ( .D(n14460), .CLK(clk), .RST(rst), .Q(ereg[917]) );
  DFF \ereg_reg[918]  ( .D(n14459), .CLK(clk), .RST(rst), .Q(ereg[918]) );
  DFF \ereg_reg[919]  ( .D(n14458), .CLK(clk), .RST(rst), .Q(ereg[919]) );
  DFF \ereg_reg[920]  ( .D(n14457), .CLK(clk), .RST(rst), .Q(ereg[920]) );
  DFF \ereg_reg[921]  ( .D(n14456), .CLK(clk), .RST(rst), .Q(ereg[921]) );
  DFF \ereg_reg[922]  ( .D(n14455), .CLK(clk), .RST(rst), .Q(ereg[922]) );
  DFF \ereg_reg[923]  ( .D(n14454), .CLK(clk), .RST(rst), .Q(ereg[923]) );
  DFF \ereg_reg[924]  ( .D(n14453), .CLK(clk), .RST(rst), .Q(ereg[924]) );
  DFF \ereg_reg[925]  ( .D(n14452), .CLK(clk), .RST(rst), .Q(ereg[925]) );
  DFF \ereg_reg[926]  ( .D(n14451), .CLK(clk), .RST(rst), .Q(ereg[926]) );
  DFF \ereg_reg[927]  ( .D(n14450), .CLK(clk), .RST(rst), .Q(ereg[927]) );
  DFF \ereg_reg[928]  ( .D(n14449), .CLK(clk), .RST(rst), .Q(ereg[928]) );
  DFF \ereg_reg[929]  ( .D(n14448), .CLK(clk), .RST(rst), .Q(ereg[929]) );
  DFF \ereg_reg[930]  ( .D(n14447), .CLK(clk), .RST(rst), .Q(ereg[930]) );
  DFF \ereg_reg[931]  ( .D(n14446), .CLK(clk), .RST(rst), .Q(ereg[931]) );
  DFF \ereg_reg[932]  ( .D(n14445), .CLK(clk), .RST(rst), .Q(ereg[932]) );
  DFF \ereg_reg[933]  ( .D(n14444), .CLK(clk), .RST(rst), .Q(ereg[933]) );
  DFF \ereg_reg[934]  ( .D(n14443), .CLK(clk), .RST(rst), .Q(ereg[934]) );
  DFF \ereg_reg[935]  ( .D(n14442), .CLK(clk), .RST(rst), .Q(ereg[935]) );
  DFF \ereg_reg[936]  ( .D(n14441), .CLK(clk), .RST(rst), .Q(ereg[936]) );
  DFF \ereg_reg[937]  ( .D(n14440), .CLK(clk), .RST(rst), .Q(ereg[937]) );
  DFF \ereg_reg[938]  ( .D(n14439), .CLK(clk), .RST(rst), .Q(ereg[938]) );
  DFF \ereg_reg[939]  ( .D(n14438), .CLK(clk), .RST(rst), .Q(ereg[939]) );
  DFF \ereg_reg[940]  ( .D(n14437), .CLK(clk), .RST(rst), .Q(ereg[940]) );
  DFF \ereg_reg[941]  ( .D(n14436), .CLK(clk), .RST(rst), .Q(ereg[941]) );
  DFF \ereg_reg[942]  ( .D(n14435), .CLK(clk), .RST(rst), .Q(ereg[942]) );
  DFF \ereg_reg[943]  ( .D(n14434), .CLK(clk), .RST(rst), .Q(ereg[943]) );
  DFF \ereg_reg[944]  ( .D(n14433), .CLK(clk), .RST(rst), .Q(ereg[944]) );
  DFF \ereg_reg[945]  ( .D(n14432), .CLK(clk), .RST(rst), .Q(ereg[945]) );
  DFF \ereg_reg[946]  ( .D(n14431), .CLK(clk), .RST(rst), .Q(ereg[946]) );
  DFF \ereg_reg[947]  ( .D(n14430), .CLK(clk), .RST(rst), .Q(ereg[947]) );
  DFF \ereg_reg[948]  ( .D(n14429), .CLK(clk), .RST(rst), .Q(ereg[948]) );
  DFF \ereg_reg[949]  ( .D(n14428), .CLK(clk), .RST(rst), .Q(ereg[949]) );
  DFF \ereg_reg[950]  ( .D(n14427), .CLK(clk), .RST(rst), .Q(ereg[950]) );
  DFF \ereg_reg[951]  ( .D(n14426), .CLK(clk), .RST(rst), .Q(ereg[951]) );
  DFF \ereg_reg[952]  ( .D(n14425), .CLK(clk), .RST(rst), .Q(ereg[952]) );
  DFF \ereg_reg[953]  ( .D(n14424), .CLK(clk), .RST(rst), .Q(ereg[953]) );
  DFF \ereg_reg[954]  ( .D(n14423), .CLK(clk), .RST(rst), .Q(ereg[954]) );
  DFF \ereg_reg[955]  ( .D(n14422), .CLK(clk), .RST(rst), .Q(ereg[955]) );
  DFF \ereg_reg[956]  ( .D(n14421), .CLK(clk), .RST(rst), .Q(ereg[956]) );
  DFF \ereg_reg[957]  ( .D(n14420), .CLK(clk), .RST(rst), .Q(ereg[957]) );
  DFF \ereg_reg[958]  ( .D(n14419), .CLK(clk), .RST(rst), .Q(ereg[958]) );
  DFF \ereg_reg[959]  ( .D(n14418), .CLK(clk), .RST(rst), .Q(ereg[959]) );
  DFF \ereg_reg[960]  ( .D(n14417), .CLK(clk), .RST(rst), .Q(ereg[960]) );
  DFF \ereg_reg[961]  ( .D(n14416), .CLK(clk), .RST(rst), .Q(ereg[961]) );
  DFF \ereg_reg[962]  ( .D(n14415), .CLK(clk), .RST(rst), .Q(ereg[962]) );
  DFF \ereg_reg[963]  ( .D(n14414), .CLK(clk), .RST(rst), .Q(ereg[963]) );
  DFF \ereg_reg[964]  ( .D(n14413), .CLK(clk), .RST(rst), .Q(ereg[964]) );
  DFF \ereg_reg[965]  ( .D(n14412), .CLK(clk), .RST(rst), .Q(ereg[965]) );
  DFF \ereg_reg[966]  ( .D(n14411), .CLK(clk), .RST(rst), .Q(ereg[966]) );
  DFF \ereg_reg[967]  ( .D(n14410), .CLK(clk), .RST(rst), .Q(ereg[967]) );
  DFF \ereg_reg[968]  ( .D(n14409), .CLK(clk), .RST(rst), .Q(ereg[968]) );
  DFF \ereg_reg[969]  ( .D(n14408), .CLK(clk), .RST(rst), .Q(ereg[969]) );
  DFF \ereg_reg[970]  ( .D(n14407), .CLK(clk), .RST(rst), .Q(ereg[970]) );
  DFF \ereg_reg[971]  ( .D(n14406), .CLK(clk), .RST(rst), .Q(ereg[971]) );
  DFF \ereg_reg[972]  ( .D(n14405), .CLK(clk), .RST(rst), .Q(ereg[972]) );
  DFF \ereg_reg[973]  ( .D(n14404), .CLK(clk), .RST(rst), .Q(ereg[973]) );
  DFF \ereg_reg[974]  ( .D(n14403), .CLK(clk), .RST(rst), .Q(ereg[974]) );
  DFF \ereg_reg[975]  ( .D(n14402), .CLK(clk), .RST(rst), .Q(ereg[975]) );
  DFF \ereg_reg[976]  ( .D(n14401), .CLK(clk), .RST(rst), .Q(ereg[976]) );
  DFF \ereg_reg[977]  ( .D(n14400), .CLK(clk), .RST(rst), .Q(ereg[977]) );
  DFF \ereg_reg[978]  ( .D(n14399), .CLK(clk), .RST(rst), .Q(ereg[978]) );
  DFF \ereg_reg[979]  ( .D(n14398), .CLK(clk), .RST(rst), .Q(ereg[979]) );
  DFF \ereg_reg[980]  ( .D(n14397), .CLK(clk), .RST(rst), .Q(ereg[980]) );
  DFF \ereg_reg[981]  ( .D(n14396), .CLK(clk), .RST(rst), .Q(ereg[981]) );
  DFF \ereg_reg[982]  ( .D(n14395), .CLK(clk), .RST(rst), .Q(ereg[982]) );
  DFF \ereg_reg[983]  ( .D(n14394), .CLK(clk), .RST(rst), .Q(ereg[983]) );
  DFF \ereg_reg[984]  ( .D(n14393), .CLK(clk), .RST(rst), .Q(ereg[984]) );
  DFF \ereg_reg[985]  ( .D(n14392), .CLK(clk), .RST(rst), .Q(ereg[985]) );
  DFF \ereg_reg[986]  ( .D(n14391), .CLK(clk), .RST(rst), .Q(ereg[986]) );
  DFF \ereg_reg[987]  ( .D(n14390), .CLK(clk), .RST(rst), .Q(ereg[987]) );
  DFF \ereg_reg[988]  ( .D(n14389), .CLK(clk), .RST(rst), .Q(ereg[988]) );
  DFF \ereg_reg[989]  ( .D(n14388), .CLK(clk), .RST(rst), .Q(ereg[989]) );
  DFF \ereg_reg[990]  ( .D(n14387), .CLK(clk), .RST(rst), .Q(ereg[990]) );
  DFF \ereg_reg[991]  ( .D(n14386), .CLK(clk), .RST(rst), .Q(ereg[991]) );
  DFF \ereg_reg[992]  ( .D(n14385), .CLK(clk), .RST(rst), .Q(ereg[992]) );
  DFF \ereg_reg[993]  ( .D(n14384), .CLK(clk), .RST(rst), .Q(ereg[993]) );
  DFF \ereg_reg[994]  ( .D(n14383), .CLK(clk), .RST(rst), .Q(ereg[994]) );
  DFF \ereg_reg[995]  ( .D(n14382), .CLK(clk), .RST(rst), .Q(ereg[995]) );
  DFF \ereg_reg[996]  ( .D(n14381), .CLK(clk), .RST(rst), .Q(ereg[996]) );
  DFF \ereg_reg[997]  ( .D(n14380), .CLK(clk), .RST(rst), .Q(ereg[997]) );
  DFF \ereg_reg[998]  ( .D(n14379), .CLK(clk), .RST(rst), .Q(ereg[998]) );
  DFF \ereg_reg[999]  ( .D(n14378), .CLK(clk), .RST(rst), .Q(ereg[999]) );
  DFF \ereg_reg[1000]  ( .D(n14377), .CLK(clk), .RST(rst), .Q(ereg[1000]) );
  DFF \ereg_reg[1001]  ( .D(n14376), .CLK(clk), .RST(rst), .Q(ereg[1001]) );
  DFF \ereg_reg[1002]  ( .D(n14375), .CLK(clk), .RST(rst), .Q(ereg[1002]) );
  DFF \ereg_reg[1003]  ( .D(n14374), .CLK(clk), .RST(rst), .Q(ereg[1003]) );
  DFF \ereg_reg[1004]  ( .D(n14373), .CLK(clk), .RST(rst), .Q(ereg[1004]) );
  DFF \ereg_reg[1005]  ( .D(n14372), .CLK(clk), .RST(rst), .Q(ereg[1005]) );
  DFF \ereg_reg[1006]  ( .D(n14371), .CLK(clk), .RST(rst), .Q(ereg[1006]) );
  DFF \ereg_reg[1007]  ( .D(n14370), .CLK(clk), .RST(rst), .Q(ereg[1007]) );
  DFF \ereg_reg[1008]  ( .D(n14369), .CLK(clk), .RST(rst), .Q(ereg[1008]) );
  DFF \ereg_reg[1009]  ( .D(n14368), .CLK(clk), .RST(rst), .Q(ereg[1009]) );
  DFF \ereg_reg[1010]  ( .D(n14367), .CLK(clk), .RST(rst), .Q(ereg[1010]) );
  DFF \ereg_reg[1011]  ( .D(n14366), .CLK(clk), .RST(rst), .Q(ereg[1011]) );
  DFF \ereg_reg[1012]  ( .D(n14365), .CLK(clk), .RST(rst), .Q(ereg[1012]) );
  DFF \ereg_reg[1013]  ( .D(n14364), .CLK(clk), .RST(rst), .Q(ereg[1013]) );
  DFF \ereg_reg[1014]  ( .D(n14363), .CLK(clk), .RST(rst), .Q(ereg[1014]) );
  DFF \ereg_reg[1015]  ( .D(n14362), .CLK(clk), .RST(rst), .Q(ereg[1015]) );
  DFF \ereg_reg[1016]  ( .D(n14361), .CLK(clk), .RST(rst), .Q(ereg[1016]) );
  DFF \ereg_reg[1017]  ( .D(n14360), .CLK(clk), .RST(rst), .Q(ereg[1017]) );
  DFF \ereg_reg[1018]  ( .D(n14359), .CLK(clk), .RST(rst), .Q(ereg[1018]) );
  DFF \ereg_reg[1019]  ( .D(n14358), .CLK(clk), .RST(rst), .Q(ereg[1019]) );
  DFF \ereg_reg[1020]  ( .D(n14357), .CLK(clk), .RST(rst), .Q(ereg[1020]) );
  DFF \ereg_reg[1021]  ( .D(n14356), .CLK(clk), .RST(rst), .Q(ereg[1021]) );
  DFF \ereg_reg[1022]  ( .D(n14355), .CLK(clk), .RST(rst), .Q(ereg[1022]) );
  DFF \ereg_reg[1023]  ( .D(n14354), .CLK(clk), .RST(rst), .Q(ereg[1023]) );
  DFF first_one_reg ( .D(n13329), .CLK(clk), .RST(rst), .Q(first_one) );
  DFF \creg_reg[0]  ( .D(n14352), .CLK(clk), .RST(rst), .Q(creg[0]) );
  DFF \creg_reg[1]  ( .D(n14351), .CLK(clk), .RST(rst), .Q(creg[1]) );
  DFF \creg_reg[2]  ( .D(n14350), .CLK(clk), .RST(rst), .Q(creg[2]) );
  DFF \creg_reg[3]  ( .D(n14349), .CLK(clk), .RST(rst), .Q(creg[3]) );
  DFF \creg_reg[4]  ( .D(n14348), .CLK(clk), .RST(rst), .Q(creg[4]) );
  DFF \creg_reg[5]  ( .D(n14347), .CLK(clk), .RST(rst), .Q(creg[5]) );
  DFF \creg_reg[6]  ( .D(n14346), .CLK(clk), .RST(rst), .Q(creg[6]) );
  DFF \creg_reg[7]  ( .D(n14345), .CLK(clk), .RST(rst), .Q(creg[7]) );
  DFF \creg_reg[8]  ( .D(n14344), .CLK(clk), .RST(rst), .Q(creg[8]) );
  DFF \creg_reg[9]  ( .D(n14343), .CLK(clk), .RST(rst), .Q(creg[9]) );
  DFF \creg_reg[10]  ( .D(n14342), .CLK(clk), .RST(rst), .Q(creg[10]) );
  DFF \creg_reg[11]  ( .D(n14341), .CLK(clk), .RST(rst), .Q(creg[11]) );
  DFF \creg_reg[12]  ( .D(n14340), .CLK(clk), .RST(rst), .Q(creg[12]) );
  DFF \creg_reg[13]  ( .D(n14339), .CLK(clk), .RST(rst), .Q(creg[13]) );
  DFF \creg_reg[14]  ( .D(n14338), .CLK(clk), .RST(rst), .Q(creg[14]) );
  DFF \creg_reg[15]  ( .D(n14337), .CLK(clk), .RST(rst), .Q(creg[15]) );
  DFF \creg_reg[16]  ( .D(n14336), .CLK(clk), .RST(rst), .Q(creg[16]) );
  DFF \creg_reg[17]  ( .D(n14335), .CLK(clk), .RST(rst), .Q(creg[17]) );
  DFF \creg_reg[18]  ( .D(n14334), .CLK(clk), .RST(rst), .Q(creg[18]) );
  DFF \creg_reg[19]  ( .D(n14333), .CLK(clk), .RST(rst), .Q(creg[19]) );
  DFF \creg_reg[20]  ( .D(n14332), .CLK(clk), .RST(rst), .Q(creg[20]) );
  DFF \creg_reg[21]  ( .D(n14331), .CLK(clk), .RST(rst), .Q(creg[21]) );
  DFF \creg_reg[22]  ( .D(n14330), .CLK(clk), .RST(rst), .Q(creg[22]) );
  DFF \creg_reg[23]  ( .D(n14329), .CLK(clk), .RST(rst), .Q(creg[23]) );
  DFF \creg_reg[24]  ( .D(n14328), .CLK(clk), .RST(rst), .Q(creg[24]) );
  DFF \creg_reg[25]  ( .D(n14327), .CLK(clk), .RST(rst), .Q(creg[25]) );
  DFF \creg_reg[26]  ( .D(n14326), .CLK(clk), .RST(rst), .Q(creg[26]) );
  DFF \creg_reg[27]  ( .D(n14325), .CLK(clk), .RST(rst), .Q(creg[27]) );
  DFF \creg_reg[28]  ( .D(n14324), .CLK(clk), .RST(rst), .Q(creg[28]) );
  DFF \creg_reg[29]  ( .D(n14323), .CLK(clk), .RST(rst), .Q(creg[29]) );
  DFF \creg_reg[30]  ( .D(n14322), .CLK(clk), .RST(rst), .Q(creg[30]) );
  DFF \creg_reg[31]  ( .D(n14321), .CLK(clk), .RST(rst), .Q(creg[31]) );
  DFF \creg_reg[32]  ( .D(n14320), .CLK(clk), .RST(rst), .Q(creg[32]) );
  DFF \creg_reg[33]  ( .D(n14319), .CLK(clk), .RST(rst), .Q(creg[33]) );
  DFF \creg_reg[34]  ( .D(n14318), .CLK(clk), .RST(rst), .Q(creg[34]) );
  DFF \creg_reg[35]  ( .D(n14317), .CLK(clk), .RST(rst), .Q(creg[35]) );
  DFF \creg_reg[36]  ( .D(n14316), .CLK(clk), .RST(rst), .Q(creg[36]) );
  DFF \creg_reg[37]  ( .D(n14315), .CLK(clk), .RST(rst), .Q(creg[37]) );
  DFF \creg_reg[38]  ( .D(n14314), .CLK(clk), .RST(rst), .Q(creg[38]) );
  DFF \creg_reg[39]  ( .D(n14313), .CLK(clk), .RST(rst), .Q(creg[39]) );
  DFF \creg_reg[40]  ( .D(n14312), .CLK(clk), .RST(rst), .Q(creg[40]) );
  DFF \creg_reg[41]  ( .D(n14311), .CLK(clk), .RST(rst), .Q(creg[41]) );
  DFF \creg_reg[42]  ( .D(n14310), .CLK(clk), .RST(rst), .Q(creg[42]) );
  DFF \creg_reg[43]  ( .D(n14309), .CLK(clk), .RST(rst), .Q(creg[43]) );
  DFF \creg_reg[44]  ( .D(n14308), .CLK(clk), .RST(rst), .Q(creg[44]) );
  DFF \creg_reg[45]  ( .D(n14307), .CLK(clk), .RST(rst), .Q(creg[45]) );
  DFF \creg_reg[46]  ( .D(n14306), .CLK(clk), .RST(rst), .Q(creg[46]) );
  DFF \creg_reg[47]  ( .D(n14305), .CLK(clk), .RST(rst), .Q(creg[47]) );
  DFF \creg_reg[48]  ( .D(n14304), .CLK(clk), .RST(rst), .Q(creg[48]) );
  DFF \creg_reg[49]  ( .D(n14303), .CLK(clk), .RST(rst), .Q(creg[49]) );
  DFF \creg_reg[50]  ( .D(n14302), .CLK(clk), .RST(rst), .Q(creg[50]) );
  DFF \creg_reg[51]  ( .D(n14301), .CLK(clk), .RST(rst), .Q(creg[51]) );
  DFF \creg_reg[52]  ( .D(n14300), .CLK(clk), .RST(rst), .Q(creg[52]) );
  DFF \creg_reg[53]  ( .D(n14299), .CLK(clk), .RST(rst), .Q(creg[53]) );
  DFF \creg_reg[54]  ( .D(n14298), .CLK(clk), .RST(rst), .Q(creg[54]) );
  DFF \creg_reg[55]  ( .D(n14297), .CLK(clk), .RST(rst), .Q(creg[55]) );
  DFF \creg_reg[56]  ( .D(n14296), .CLK(clk), .RST(rst), .Q(creg[56]) );
  DFF \creg_reg[57]  ( .D(n14295), .CLK(clk), .RST(rst), .Q(creg[57]) );
  DFF \creg_reg[58]  ( .D(n14294), .CLK(clk), .RST(rst), .Q(creg[58]) );
  DFF \creg_reg[59]  ( .D(n14293), .CLK(clk), .RST(rst), .Q(creg[59]) );
  DFF \creg_reg[60]  ( .D(n14292), .CLK(clk), .RST(rst), .Q(creg[60]) );
  DFF \creg_reg[61]  ( .D(n14291), .CLK(clk), .RST(rst), .Q(creg[61]) );
  DFF \creg_reg[62]  ( .D(n14290), .CLK(clk), .RST(rst), .Q(creg[62]) );
  DFF \creg_reg[63]  ( .D(n14289), .CLK(clk), .RST(rst), .Q(creg[63]) );
  DFF \creg_reg[64]  ( .D(n14288), .CLK(clk), .RST(rst), .Q(creg[64]) );
  DFF \creg_reg[65]  ( .D(n14287), .CLK(clk), .RST(rst), .Q(creg[65]) );
  DFF \creg_reg[66]  ( .D(n14286), .CLK(clk), .RST(rst), .Q(creg[66]) );
  DFF \creg_reg[67]  ( .D(n14285), .CLK(clk), .RST(rst), .Q(creg[67]) );
  DFF \creg_reg[68]  ( .D(n14284), .CLK(clk), .RST(rst), .Q(creg[68]) );
  DFF \creg_reg[69]  ( .D(n14283), .CLK(clk), .RST(rst), .Q(creg[69]) );
  DFF \creg_reg[70]  ( .D(n14282), .CLK(clk), .RST(rst), .Q(creg[70]) );
  DFF \creg_reg[71]  ( .D(n14281), .CLK(clk), .RST(rst), .Q(creg[71]) );
  DFF \creg_reg[72]  ( .D(n14280), .CLK(clk), .RST(rst), .Q(creg[72]) );
  DFF \creg_reg[73]  ( .D(n14279), .CLK(clk), .RST(rst), .Q(creg[73]) );
  DFF \creg_reg[74]  ( .D(n14278), .CLK(clk), .RST(rst), .Q(creg[74]) );
  DFF \creg_reg[75]  ( .D(n14277), .CLK(clk), .RST(rst), .Q(creg[75]) );
  DFF \creg_reg[76]  ( .D(n14276), .CLK(clk), .RST(rst), .Q(creg[76]) );
  DFF \creg_reg[77]  ( .D(n14275), .CLK(clk), .RST(rst), .Q(creg[77]) );
  DFF \creg_reg[78]  ( .D(n14274), .CLK(clk), .RST(rst), .Q(creg[78]) );
  DFF \creg_reg[79]  ( .D(n14273), .CLK(clk), .RST(rst), .Q(creg[79]) );
  DFF \creg_reg[80]  ( .D(n14272), .CLK(clk), .RST(rst), .Q(creg[80]) );
  DFF \creg_reg[81]  ( .D(n14271), .CLK(clk), .RST(rst), .Q(creg[81]) );
  DFF \creg_reg[82]  ( .D(n14270), .CLK(clk), .RST(rst), .Q(creg[82]) );
  DFF \creg_reg[83]  ( .D(n14269), .CLK(clk), .RST(rst), .Q(creg[83]) );
  DFF \creg_reg[84]  ( .D(n14268), .CLK(clk), .RST(rst), .Q(creg[84]) );
  DFF \creg_reg[85]  ( .D(n14267), .CLK(clk), .RST(rst), .Q(creg[85]) );
  DFF \creg_reg[86]  ( .D(n14266), .CLK(clk), .RST(rst), .Q(creg[86]) );
  DFF \creg_reg[87]  ( .D(n14265), .CLK(clk), .RST(rst), .Q(creg[87]) );
  DFF \creg_reg[88]  ( .D(n14264), .CLK(clk), .RST(rst), .Q(creg[88]) );
  DFF \creg_reg[89]  ( .D(n14263), .CLK(clk), .RST(rst), .Q(creg[89]) );
  DFF \creg_reg[90]  ( .D(n14262), .CLK(clk), .RST(rst), .Q(creg[90]) );
  DFF \creg_reg[91]  ( .D(n14261), .CLK(clk), .RST(rst), .Q(creg[91]) );
  DFF \creg_reg[92]  ( .D(n14260), .CLK(clk), .RST(rst), .Q(creg[92]) );
  DFF \creg_reg[93]  ( .D(n14259), .CLK(clk), .RST(rst), .Q(creg[93]) );
  DFF \creg_reg[94]  ( .D(n14258), .CLK(clk), .RST(rst), .Q(creg[94]) );
  DFF \creg_reg[95]  ( .D(n14257), .CLK(clk), .RST(rst), .Q(creg[95]) );
  DFF \creg_reg[96]  ( .D(n14256), .CLK(clk), .RST(rst), .Q(creg[96]) );
  DFF \creg_reg[97]  ( .D(n14255), .CLK(clk), .RST(rst), .Q(creg[97]) );
  DFF \creg_reg[98]  ( .D(n14254), .CLK(clk), .RST(rst), .Q(creg[98]) );
  DFF \creg_reg[99]  ( .D(n14253), .CLK(clk), .RST(rst), .Q(creg[99]) );
  DFF \creg_reg[100]  ( .D(n14252), .CLK(clk), .RST(rst), .Q(creg[100]) );
  DFF \creg_reg[101]  ( .D(n14251), .CLK(clk), .RST(rst), .Q(creg[101]) );
  DFF \creg_reg[102]  ( .D(n14250), .CLK(clk), .RST(rst), .Q(creg[102]) );
  DFF \creg_reg[103]  ( .D(n14249), .CLK(clk), .RST(rst), .Q(creg[103]) );
  DFF \creg_reg[104]  ( .D(n14248), .CLK(clk), .RST(rst), .Q(creg[104]) );
  DFF \creg_reg[105]  ( .D(n14247), .CLK(clk), .RST(rst), .Q(creg[105]) );
  DFF \creg_reg[106]  ( .D(n14246), .CLK(clk), .RST(rst), .Q(creg[106]) );
  DFF \creg_reg[107]  ( .D(n14245), .CLK(clk), .RST(rst), .Q(creg[107]) );
  DFF \creg_reg[108]  ( .D(n14244), .CLK(clk), .RST(rst), .Q(creg[108]) );
  DFF \creg_reg[109]  ( .D(n14243), .CLK(clk), .RST(rst), .Q(creg[109]) );
  DFF \creg_reg[110]  ( .D(n14242), .CLK(clk), .RST(rst), .Q(creg[110]) );
  DFF \creg_reg[111]  ( .D(n14241), .CLK(clk), .RST(rst), .Q(creg[111]) );
  DFF \creg_reg[112]  ( .D(n14240), .CLK(clk), .RST(rst), .Q(creg[112]) );
  DFF \creg_reg[113]  ( .D(n14239), .CLK(clk), .RST(rst), .Q(creg[113]) );
  DFF \creg_reg[114]  ( .D(n14238), .CLK(clk), .RST(rst), .Q(creg[114]) );
  DFF \creg_reg[115]  ( .D(n14237), .CLK(clk), .RST(rst), .Q(creg[115]) );
  DFF \creg_reg[116]  ( .D(n14236), .CLK(clk), .RST(rst), .Q(creg[116]) );
  DFF \creg_reg[117]  ( .D(n14235), .CLK(clk), .RST(rst), .Q(creg[117]) );
  DFF \creg_reg[118]  ( .D(n14234), .CLK(clk), .RST(rst), .Q(creg[118]) );
  DFF \creg_reg[119]  ( .D(n14233), .CLK(clk), .RST(rst), .Q(creg[119]) );
  DFF \creg_reg[120]  ( .D(n14232), .CLK(clk), .RST(rst), .Q(creg[120]) );
  DFF \creg_reg[121]  ( .D(n14231), .CLK(clk), .RST(rst), .Q(creg[121]) );
  DFF \creg_reg[122]  ( .D(n14230), .CLK(clk), .RST(rst), .Q(creg[122]) );
  DFF \creg_reg[123]  ( .D(n14229), .CLK(clk), .RST(rst), .Q(creg[123]) );
  DFF \creg_reg[124]  ( .D(n14228), .CLK(clk), .RST(rst), .Q(creg[124]) );
  DFF \creg_reg[125]  ( .D(n14227), .CLK(clk), .RST(rst), .Q(creg[125]) );
  DFF \creg_reg[126]  ( .D(n14226), .CLK(clk), .RST(rst), .Q(creg[126]) );
  DFF \creg_reg[127]  ( .D(n14225), .CLK(clk), .RST(rst), .Q(creg[127]) );
  DFF \creg_reg[128]  ( .D(n14224), .CLK(clk), .RST(rst), .Q(creg[128]) );
  DFF \creg_reg[129]  ( .D(n14223), .CLK(clk), .RST(rst), .Q(creg[129]) );
  DFF \creg_reg[130]  ( .D(n14222), .CLK(clk), .RST(rst), .Q(creg[130]) );
  DFF \creg_reg[131]  ( .D(n14221), .CLK(clk), .RST(rst), .Q(creg[131]) );
  DFF \creg_reg[132]  ( .D(n14220), .CLK(clk), .RST(rst), .Q(creg[132]) );
  DFF \creg_reg[133]  ( .D(n14219), .CLK(clk), .RST(rst), .Q(creg[133]) );
  DFF \creg_reg[134]  ( .D(n14218), .CLK(clk), .RST(rst), .Q(creg[134]) );
  DFF \creg_reg[135]  ( .D(n14217), .CLK(clk), .RST(rst), .Q(creg[135]) );
  DFF \creg_reg[136]  ( .D(n14216), .CLK(clk), .RST(rst), .Q(creg[136]) );
  DFF \creg_reg[137]  ( .D(n14215), .CLK(clk), .RST(rst), .Q(creg[137]) );
  DFF \creg_reg[138]  ( .D(n14214), .CLK(clk), .RST(rst), .Q(creg[138]) );
  DFF \creg_reg[139]  ( .D(n14213), .CLK(clk), .RST(rst), .Q(creg[139]) );
  DFF \creg_reg[140]  ( .D(n14212), .CLK(clk), .RST(rst), .Q(creg[140]) );
  DFF \creg_reg[141]  ( .D(n14211), .CLK(clk), .RST(rst), .Q(creg[141]) );
  DFF \creg_reg[142]  ( .D(n14210), .CLK(clk), .RST(rst), .Q(creg[142]) );
  DFF \creg_reg[143]  ( .D(n14209), .CLK(clk), .RST(rst), .Q(creg[143]) );
  DFF \creg_reg[144]  ( .D(n14208), .CLK(clk), .RST(rst), .Q(creg[144]) );
  DFF \creg_reg[145]  ( .D(n14207), .CLK(clk), .RST(rst), .Q(creg[145]) );
  DFF \creg_reg[146]  ( .D(n14206), .CLK(clk), .RST(rst), .Q(creg[146]) );
  DFF \creg_reg[147]  ( .D(n14205), .CLK(clk), .RST(rst), .Q(creg[147]) );
  DFF \creg_reg[148]  ( .D(n14204), .CLK(clk), .RST(rst), .Q(creg[148]) );
  DFF \creg_reg[149]  ( .D(n14203), .CLK(clk), .RST(rst), .Q(creg[149]) );
  DFF \creg_reg[150]  ( .D(n14202), .CLK(clk), .RST(rst), .Q(creg[150]) );
  DFF \creg_reg[151]  ( .D(n14201), .CLK(clk), .RST(rst), .Q(creg[151]) );
  DFF \creg_reg[152]  ( .D(n14200), .CLK(clk), .RST(rst), .Q(creg[152]) );
  DFF \creg_reg[153]  ( .D(n14199), .CLK(clk), .RST(rst), .Q(creg[153]) );
  DFF \creg_reg[154]  ( .D(n14198), .CLK(clk), .RST(rst), .Q(creg[154]) );
  DFF \creg_reg[155]  ( .D(n14197), .CLK(clk), .RST(rst), .Q(creg[155]) );
  DFF \creg_reg[156]  ( .D(n14196), .CLK(clk), .RST(rst), .Q(creg[156]) );
  DFF \creg_reg[157]  ( .D(n14195), .CLK(clk), .RST(rst), .Q(creg[157]) );
  DFF \creg_reg[158]  ( .D(n14194), .CLK(clk), .RST(rst), .Q(creg[158]) );
  DFF \creg_reg[159]  ( .D(n14193), .CLK(clk), .RST(rst), .Q(creg[159]) );
  DFF \creg_reg[160]  ( .D(n14192), .CLK(clk), .RST(rst), .Q(creg[160]) );
  DFF \creg_reg[161]  ( .D(n14191), .CLK(clk), .RST(rst), .Q(creg[161]) );
  DFF \creg_reg[162]  ( .D(n14190), .CLK(clk), .RST(rst), .Q(creg[162]) );
  DFF \creg_reg[163]  ( .D(n14189), .CLK(clk), .RST(rst), .Q(creg[163]) );
  DFF \creg_reg[164]  ( .D(n14188), .CLK(clk), .RST(rst), .Q(creg[164]) );
  DFF \creg_reg[165]  ( .D(n14187), .CLK(clk), .RST(rst), .Q(creg[165]) );
  DFF \creg_reg[166]  ( .D(n14186), .CLK(clk), .RST(rst), .Q(creg[166]) );
  DFF \creg_reg[167]  ( .D(n14185), .CLK(clk), .RST(rst), .Q(creg[167]) );
  DFF \creg_reg[168]  ( .D(n14184), .CLK(clk), .RST(rst), .Q(creg[168]) );
  DFF \creg_reg[169]  ( .D(n14183), .CLK(clk), .RST(rst), .Q(creg[169]) );
  DFF \creg_reg[170]  ( .D(n14182), .CLK(clk), .RST(rst), .Q(creg[170]) );
  DFF \creg_reg[171]  ( .D(n14181), .CLK(clk), .RST(rst), .Q(creg[171]) );
  DFF \creg_reg[172]  ( .D(n14180), .CLK(clk), .RST(rst), .Q(creg[172]) );
  DFF \creg_reg[173]  ( .D(n14179), .CLK(clk), .RST(rst), .Q(creg[173]) );
  DFF \creg_reg[174]  ( .D(n14178), .CLK(clk), .RST(rst), .Q(creg[174]) );
  DFF \creg_reg[175]  ( .D(n14177), .CLK(clk), .RST(rst), .Q(creg[175]) );
  DFF \creg_reg[176]  ( .D(n14176), .CLK(clk), .RST(rst), .Q(creg[176]) );
  DFF \creg_reg[177]  ( .D(n14175), .CLK(clk), .RST(rst), .Q(creg[177]) );
  DFF \creg_reg[178]  ( .D(n14174), .CLK(clk), .RST(rst), .Q(creg[178]) );
  DFF \creg_reg[179]  ( .D(n14173), .CLK(clk), .RST(rst), .Q(creg[179]) );
  DFF \creg_reg[180]  ( .D(n14172), .CLK(clk), .RST(rst), .Q(creg[180]) );
  DFF \creg_reg[181]  ( .D(n14171), .CLK(clk), .RST(rst), .Q(creg[181]) );
  DFF \creg_reg[182]  ( .D(n14170), .CLK(clk), .RST(rst), .Q(creg[182]) );
  DFF \creg_reg[183]  ( .D(n14169), .CLK(clk), .RST(rst), .Q(creg[183]) );
  DFF \creg_reg[184]  ( .D(n14168), .CLK(clk), .RST(rst), .Q(creg[184]) );
  DFF \creg_reg[185]  ( .D(n14167), .CLK(clk), .RST(rst), .Q(creg[185]) );
  DFF \creg_reg[186]  ( .D(n14166), .CLK(clk), .RST(rst), .Q(creg[186]) );
  DFF \creg_reg[187]  ( .D(n14165), .CLK(clk), .RST(rst), .Q(creg[187]) );
  DFF \creg_reg[188]  ( .D(n14164), .CLK(clk), .RST(rst), .Q(creg[188]) );
  DFF \creg_reg[189]  ( .D(n14163), .CLK(clk), .RST(rst), .Q(creg[189]) );
  DFF \creg_reg[190]  ( .D(n14162), .CLK(clk), .RST(rst), .Q(creg[190]) );
  DFF \creg_reg[191]  ( .D(n14161), .CLK(clk), .RST(rst), .Q(creg[191]) );
  DFF \creg_reg[192]  ( .D(n14160), .CLK(clk), .RST(rst), .Q(creg[192]) );
  DFF \creg_reg[193]  ( .D(n14159), .CLK(clk), .RST(rst), .Q(creg[193]) );
  DFF \creg_reg[194]  ( .D(n14158), .CLK(clk), .RST(rst), .Q(creg[194]) );
  DFF \creg_reg[195]  ( .D(n14157), .CLK(clk), .RST(rst), .Q(creg[195]) );
  DFF \creg_reg[196]  ( .D(n14156), .CLK(clk), .RST(rst), .Q(creg[196]) );
  DFF \creg_reg[197]  ( .D(n14155), .CLK(clk), .RST(rst), .Q(creg[197]) );
  DFF \creg_reg[198]  ( .D(n14154), .CLK(clk), .RST(rst), .Q(creg[198]) );
  DFF \creg_reg[199]  ( .D(n14153), .CLK(clk), .RST(rst), .Q(creg[199]) );
  DFF \creg_reg[200]  ( .D(n14152), .CLK(clk), .RST(rst), .Q(creg[200]) );
  DFF \creg_reg[201]  ( .D(n14151), .CLK(clk), .RST(rst), .Q(creg[201]) );
  DFF \creg_reg[202]  ( .D(n14150), .CLK(clk), .RST(rst), .Q(creg[202]) );
  DFF \creg_reg[203]  ( .D(n14149), .CLK(clk), .RST(rst), .Q(creg[203]) );
  DFF \creg_reg[204]  ( .D(n14148), .CLK(clk), .RST(rst), .Q(creg[204]) );
  DFF \creg_reg[205]  ( .D(n14147), .CLK(clk), .RST(rst), .Q(creg[205]) );
  DFF \creg_reg[206]  ( .D(n14146), .CLK(clk), .RST(rst), .Q(creg[206]) );
  DFF \creg_reg[207]  ( .D(n14145), .CLK(clk), .RST(rst), .Q(creg[207]) );
  DFF \creg_reg[208]  ( .D(n14144), .CLK(clk), .RST(rst), .Q(creg[208]) );
  DFF \creg_reg[209]  ( .D(n14143), .CLK(clk), .RST(rst), .Q(creg[209]) );
  DFF \creg_reg[210]  ( .D(n14142), .CLK(clk), .RST(rst), .Q(creg[210]) );
  DFF \creg_reg[211]  ( .D(n14141), .CLK(clk), .RST(rst), .Q(creg[211]) );
  DFF \creg_reg[212]  ( .D(n14140), .CLK(clk), .RST(rst), .Q(creg[212]) );
  DFF \creg_reg[213]  ( .D(n14139), .CLK(clk), .RST(rst), .Q(creg[213]) );
  DFF \creg_reg[214]  ( .D(n14138), .CLK(clk), .RST(rst), .Q(creg[214]) );
  DFF \creg_reg[215]  ( .D(n14137), .CLK(clk), .RST(rst), .Q(creg[215]) );
  DFF \creg_reg[216]  ( .D(n14136), .CLK(clk), .RST(rst), .Q(creg[216]) );
  DFF \creg_reg[217]  ( .D(n14135), .CLK(clk), .RST(rst), .Q(creg[217]) );
  DFF \creg_reg[218]  ( .D(n14134), .CLK(clk), .RST(rst), .Q(creg[218]) );
  DFF \creg_reg[219]  ( .D(n14133), .CLK(clk), .RST(rst), .Q(creg[219]) );
  DFF \creg_reg[220]  ( .D(n14132), .CLK(clk), .RST(rst), .Q(creg[220]) );
  DFF \creg_reg[221]  ( .D(n14131), .CLK(clk), .RST(rst), .Q(creg[221]) );
  DFF \creg_reg[222]  ( .D(n14130), .CLK(clk), .RST(rst), .Q(creg[222]) );
  DFF \creg_reg[223]  ( .D(n14129), .CLK(clk), .RST(rst), .Q(creg[223]) );
  DFF \creg_reg[224]  ( .D(n14128), .CLK(clk), .RST(rst), .Q(creg[224]) );
  DFF \creg_reg[225]  ( .D(n14127), .CLK(clk), .RST(rst), .Q(creg[225]) );
  DFF \creg_reg[226]  ( .D(n14126), .CLK(clk), .RST(rst), .Q(creg[226]) );
  DFF \creg_reg[227]  ( .D(n14125), .CLK(clk), .RST(rst), .Q(creg[227]) );
  DFF \creg_reg[228]  ( .D(n14124), .CLK(clk), .RST(rst), .Q(creg[228]) );
  DFF \creg_reg[229]  ( .D(n14123), .CLK(clk), .RST(rst), .Q(creg[229]) );
  DFF \creg_reg[230]  ( .D(n14122), .CLK(clk), .RST(rst), .Q(creg[230]) );
  DFF \creg_reg[231]  ( .D(n14121), .CLK(clk), .RST(rst), .Q(creg[231]) );
  DFF \creg_reg[232]  ( .D(n14120), .CLK(clk), .RST(rst), .Q(creg[232]) );
  DFF \creg_reg[233]  ( .D(n14119), .CLK(clk), .RST(rst), .Q(creg[233]) );
  DFF \creg_reg[234]  ( .D(n14118), .CLK(clk), .RST(rst), .Q(creg[234]) );
  DFF \creg_reg[235]  ( .D(n14117), .CLK(clk), .RST(rst), .Q(creg[235]) );
  DFF \creg_reg[236]  ( .D(n14116), .CLK(clk), .RST(rst), .Q(creg[236]) );
  DFF \creg_reg[237]  ( .D(n14115), .CLK(clk), .RST(rst), .Q(creg[237]) );
  DFF \creg_reg[238]  ( .D(n14114), .CLK(clk), .RST(rst), .Q(creg[238]) );
  DFF \creg_reg[239]  ( .D(n14113), .CLK(clk), .RST(rst), .Q(creg[239]) );
  DFF \creg_reg[240]  ( .D(n14112), .CLK(clk), .RST(rst), .Q(creg[240]) );
  DFF \creg_reg[241]  ( .D(n14111), .CLK(clk), .RST(rst), .Q(creg[241]) );
  DFF \creg_reg[242]  ( .D(n14110), .CLK(clk), .RST(rst), .Q(creg[242]) );
  DFF \creg_reg[243]  ( .D(n14109), .CLK(clk), .RST(rst), .Q(creg[243]) );
  DFF \creg_reg[244]  ( .D(n14108), .CLK(clk), .RST(rst), .Q(creg[244]) );
  DFF \creg_reg[245]  ( .D(n14107), .CLK(clk), .RST(rst), .Q(creg[245]) );
  DFF \creg_reg[246]  ( .D(n14106), .CLK(clk), .RST(rst), .Q(creg[246]) );
  DFF \creg_reg[247]  ( .D(n14105), .CLK(clk), .RST(rst), .Q(creg[247]) );
  DFF \creg_reg[248]  ( .D(n14104), .CLK(clk), .RST(rst), .Q(creg[248]) );
  DFF \creg_reg[249]  ( .D(n14103), .CLK(clk), .RST(rst), .Q(creg[249]) );
  DFF \creg_reg[250]  ( .D(n14102), .CLK(clk), .RST(rst), .Q(creg[250]) );
  DFF \creg_reg[251]  ( .D(n14101), .CLK(clk), .RST(rst), .Q(creg[251]) );
  DFF \creg_reg[252]  ( .D(n14100), .CLK(clk), .RST(rst), .Q(creg[252]) );
  DFF \creg_reg[253]  ( .D(n14099), .CLK(clk), .RST(rst), .Q(creg[253]) );
  DFF \creg_reg[254]  ( .D(n14098), .CLK(clk), .RST(rst), .Q(creg[254]) );
  DFF \creg_reg[255]  ( .D(n14097), .CLK(clk), .RST(rst), .Q(creg[255]) );
  DFF \creg_reg[256]  ( .D(n14096), .CLK(clk), .RST(rst), .Q(creg[256]) );
  DFF \creg_reg[257]  ( .D(n14095), .CLK(clk), .RST(rst), .Q(creg[257]) );
  DFF \creg_reg[258]  ( .D(n14094), .CLK(clk), .RST(rst), .Q(creg[258]) );
  DFF \creg_reg[259]  ( .D(n14093), .CLK(clk), .RST(rst), .Q(creg[259]) );
  DFF \creg_reg[260]  ( .D(n14092), .CLK(clk), .RST(rst), .Q(creg[260]) );
  DFF \creg_reg[261]  ( .D(n14091), .CLK(clk), .RST(rst), .Q(creg[261]) );
  DFF \creg_reg[262]  ( .D(n14090), .CLK(clk), .RST(rst), .Q(creg[262]) );
  DFF \creg_reg[263]  ( .D(n14089), .CLK(clk), .RST(rst), .Q(creg[263]) );
  DFF \creg_reg[264]  ( .D(n14088), .CLK(clk), .RST(rst), .Q(creg[264]) );
  DFF \creg_reg[265]  ( .D(n14087), .CLK(clk), .RST(rst), .Q(creg[265]) );
  DFF \creg_reg[266]  ( .D(n14086), .CLK(clk), .RST(rst), .Q(creg[266]) );
  DFF \creg_reg[267]  ( .D(n14085), .CLK(clk), .RST(rst), .Q(creg[267]) );
  DFF \creg_reg[268]  ( .D(n14084), .CLK(clk), .RST(rst), .Q(creg[268]) );
  DFF \creg_reg[269]  ( .D(n14083), .CLK(clk), .RST(rst), .Q(creg[269]) );
  DFF \creg_reg[270]  ( .D(n14082), .CLK(clk), .RST(rst), .Q(creg[270]) );
  DFF \creg_reg[271]  ( .D(n14081), .CLK(clk), .RST(rst), .Q(creg[271]) );
  DFF \creg_reg[272]  ( .D(n14080), .CLK(clk), .RST(rst), .Q(creg[272]) );
  DFF \creg_reg[273]  ( .D(n14079), .CLK(clk), .RST(rst), .Q(creg[273]) );
  DFF \creg_reg[274]  ( .D(n14078), .CLK(clk), .RST(rst), .Q(creg[274]) );
  DFF \creg_reg[275]  ( .D(n14077), .CLK(clk), .RST(rst), .Q(creg[275]) );
  DFF \creg_reg[276]  ( .D(n14076), .CLK(clk), .RST(rst), .Q(creg[276]) );
  DFF \creg_reg[277]  ( .D(n14075), .CLK(clk), .RST(rst), .Q(creg[277]) );
  DFF \creg_reg[278]  ( .D(n14074), .CLK(clk), .RST(rst), .Q(creg[278]) );
  DFF \creg_reg[279]  ( .D(n14073), .CLK(clk), .RST(rst), .Q(creg[279]) );
  DFF \creg_reg[280]  ( .D(n14072), .CLK(clk), .RST(rst), .Q(creg[280]) );
  DFF \creg_reg[281]  ( .D(n14071), .CLK(clk), .RST(rst), .Q(creg[281]) );
  DFF \creg_reg[282]  ( .D(n14070), .CLK(clk), .RST(rst), .Q(creg[282]) );
  DFF \creg_reg[283]  ( .D(n14069), .CLK(clk), .RST(rst), .Q(creg[283]) );
  DFF \creg_reg[284]  ( .D(n14068), .CLK(clk), .RST(rst), .Q(creg[284]) );
  DFF \creg_reg[285]  ( .D(n14067), .CLK(clk), .RST(rst), .Q(creg[285]) );
  DFF \creg_reg[286]  ( .D(n14066), .CLK(clk), .RST(rst), .Q(creg[286]) );
  DFF \creg_reg[287]  ( .D(n14065), .CLK(clk), .RST(rst), .Q(creg[287]) );
  DFF \creg_reg[288]  ( .D(n14064), .CLK(clk), .RST(rst), .Q(creg[288]) );
  DFF \creg_reg[289]  ( .D(n14063), .CLK(clk), .RST(rst), .Q(creg[289]) );
  DFF \creg_reg[290]  ( .D(n14062), .CLK(clk), .RST(rst), .Q(creg[290]) );
  DFF \creg_reg[291]  ( .D(n14061), .CLK(clk), .RST(rst), .Q(creg[291]) );
  DFF \creg_reg[292]  ( .D(n14060), .CLK(clk), .RST(rst), .Q(creg[292]) );
  DFF \creg_reg[293]  ( .D(n14059), .CLK(clk), .RST(rst), .Q(creg[293]) );
  DFF \creg_reg[294]  ( .D(n14058), .CLK(clk), .RST(rst), .Q(creg[294]) );
  DFF \creg_reg[295]  ( .D(n14057), .CLK(clk), .RST(rst), .Q(creg[295]) );
  DFF \creg_reg[296]  ( .D(n14056), .CLK(clk), .RST(rst), .Q(creg[296]) );
  DFF \creg_reg[297]  ( .D(n14055), .CLK(clk), .RST(rst), .Q(creg[297]) );
  DFF \creg_reg[298]  ( .D(n14054), .CLK(clk), .RST(rst), .Q(creg[298]) );
  DFF \creg_reg[299]  ( .D(n14053), .CLK(clk), .RST(rst), .Q(creg[299]) );
  DFF \creg_reg[300]  ( .D(n14052), .CLK(clk), .RST(rst), .Q(creg[300]) );
  DFF \creg_reg[301]  ( .D(n14051), .CLK(clk), .RST(rst), .Q(creg[301]) );
  DFF \creg_reg[302]  ( .D(n14050), .CLK(clk), .RST(rst), .Q(creg[302]) );
  DFF \creg_reg[303]  ( .D(n14049), .CLK(clk), .RST(rst), .Q(creg[303]) );
  DFF \creg_reg[304]  ( .D(n14048), .CLK(clk), .RST(rst), .Q(creg[304]) );
  DFF \creg_reg[305]  ( .D(n14047), .CLK(clk), .RST(rst), .Q(creg[305]) );
  DFF \creg_reg[306]  ( .D(n14046), .CLK(clk), .RST(rst), .Q(creg[306]) );
  DFF \creg_reg[307]  ( .D(n14045), .CLK(clk), .RST(rst), .Q(creg[307]) );
  DFF \creg_reg[308]  ( .D(n14044), .CLK(clk), .RST(rst), .Q(creg[308]) );
  DFF \creg_reg[309]  ( .D(n14043), .CLK(clk), .RST(rst), .Q(creg[309]) );
  DFF \creg_reg[310]  ( .D(n14042), .CLK(clk), .RST(rst), .Q(creg[310]) );
  DFF \creg_reg[311]  ( .D(n14041), .CLK(clk), .RST(rst), .Q(creg[311]) );
  DFF \creg_reg[312]  ( .D(n14040), .CLK(clk), .RST(rst), .Q(creg[312]) );
  DFF \creg_reg[313]  ( .D(n14039), .CLK(clk), .RST(rst), .Q(creg[313]) );
  DFF \creg_reg[314]  ( .D(n14038), .CLK(clk), .RST(rst), .Q(creg[314]) );
  DFF \creg_reg[315]  ( .D(n14037), .CLK(clk), .RST(rst), .Q(creg[315]) );
  DFF \creg_reg[316]  ( .D(n14036), .CLK(clk), .RST(rst), .Q(creg[316]) );
  DFF \creg_reg[317]  ( .D(n14035), .CLK(clk), .RST(rst), .Q(creg[317]) );
  DFF \creg_reg[318]  ( .D(n14034), .CLK(clk), .RST(rst), .Q(creg[318]) );
  DFF \creg_reg[319]  ( .D(n14033), .CLK(clk), .RST(rst), .Q(creg[319]) );
  DFF \creg_reg[320]  ( .D(n14032), .CLK(clk), .RST(rst), .Q(creg[320]) );
  DFF \creg_reg[321]  ( .D(n14031), .CLK(clk), .RST(rst), .Q(creg[321]) );
  DFF \creg_reg[322]  ( .D(n14030), .CLK(clk), .RST(rst), .Q(creg[322]) );
  DFF \creg_reg[323]  ( .D(n14029), .CLK(clk), .RST(rst), .Q(creg[323]) );
  DFF \creg_reg[324]  ( .D(n14028), .CLK(clk), .RST(rst), .Q(creg[324]) );
  DFF \creg_reg[325]  ( .D(n14027), .CLK(clk), .RST(rst), .Q(creg[325]) );
  DFF \creg_reg[326]  ( .D(n14026), .CLK(clk), .RST(rst), .Q(creg[326]) );
  DFF \creg_reg[327]  ( .D(n14025), .CLK(clk), .RST(rst), .Q(creg[327]) );
  DFF \creg_reg[328]  ( .D(n14024), .CLK(clk), .RST(rst), .Q(creg[328]) );
  DFF \creg_reg[329]  ( .D(n14023), .CLK(clk), .RST(rst), .Q(creg[329]) );
  DFF \creg_reg[330]  ( .D(n14022), .CLK(clk), .RST(rst), .Q(creg[330]) );
  DFF \creg_reg[331]  ( .D(n14021), .CLK(clk), .RST(rst), .Q(creg[331]) );
  DFF \creg_reg[332]  ( .D(n14020), .CLK(clk), .RST(rst), .Q(creg[332]) );
  DFF \creg_reg[333]  ( .D(n14019), .CLK(clk), .RST(rst), .Q(creg[333]) );
  DFF \creg_reg[334]  ( .D(n14018), .CLK(clk), .RST(rst), .Q(creg[334]) );
  DFF \creg_reg[335]  ( .D(n14017), .CLK(clk), .RST(rst), .Q(creg[335]) );
  DFF \creg_reg[336]  ( .D(n14016), .CLK(clk), .RST(rst), .Q(creg[336]) );
  DFF \creg_reg[337]  ( .D(n14015), .CLK(clk), .RST(rst), .Q(creg[337]) );
  DFF \creg_reg[338]  ( .D(n14014), .CLK(clk), .RST(rst), .Q(creg[338]) );
  DFF \creg_reg[339]  ( .D(n14013), .CLK(clk), .RST(rst), .Q(creg[339]) );
  DFF \creg_reg[340]  ( .D(n14012), .CLK(clk), .RST(rst), .Q(creg[340]) );
  DFF \creg_reg[341]  ( .D(n14011), .CLK(clk), .RST(rst), .Q(creg[341]) );
  DFF \creg_reg[342]  ( .D(n14010), .CLK(clk), .RST(rst), .Q(creg[342]) );
  DFF \creg_reg[343]  ( .D(n14009), .CLK(clk), .RST(rst), .Q(creg[343]) );
  DFF \creg_reg[344]  ( .D(n14008), .CLK(clk), .RST(rst), .Q(creg[344]) );
  DFF \creg_reg[345]  ( .D(n14007), .CLK(clk), .RST(rst), .Q(creg[345]) );
  DFF \creg_reg[346]  ( .D(n14006), .CLK(clk), .RST(rst), .Q(creg[346]) );
  DFF \creg_reg[347]  ( .D(n14005), .CLK(clk), .RST(rst), .Q(creg[347]) );
  DFF \creg_reg[348]  ( .D(n14004), .CLK(clk), .RST(rst), .Q(creg[348]) );
  DFF \creg_reg[349]  ( .D(n14003), .CLK(clk), .RST(rst), .Q(creg[349]) );
  DFF \creg_reg[350]  ( .D(n14002), .CLK(clk), .RST(rst), .Q(creg[350]) );
  DFF \creg_reg[351]  ( .D(n14001), .CLK(clk), .RST(rst), .Q(creg[351]) );
  DFF \creg_reg[352]  ( .D(n14000), .CLK(clk), .RST(rst), .Q(creg[352]) );
  DFF \creg_reg[353]  ( .D(n13999), .CLK(clk), .RST(rst), .Q(creg[353]) );
  DFF \creg_reg[354]  ( .D(n13998), .CLK(clk), .RST(rst), .Q(creg[354]) );
  DFF \creg_reg[355]  ( .D(n13997), .CLK(clk), .RST(rst), .Q(creg[355]) );
  DFF \creg_reg[356]  ( .D(n13996), .CLK(clk), .RST(rst), .Q(creg[356]) );
  DFF \creg_reg[357]  ( .D(n13995), .CLK(clk), .RST(rst), .Q(creg[357]) );
  DFF \creg_reg[358]  ( .D(n13994), .CLK(clk), .RST(rst), .Q(creg[358]) );
  DFF \creg_reg[359]  ( .D(n13993), .CLK(clk), .RST(rst), .Q(creg[359]) );
  DFF \creg_reg[360]  ( .D(n13992), .CLK(clk), .RST(rst), .Q(creg[360]) );
  DFF \creg_reg[361]  ( .D(n13991), .CLK(clk), .RST(rst), .Q(creg[361]) );
  DFF \creg_reg[362]  ( .D(n13990), .CLK(clk), .RST(rst), .Q(creg[362]) );
  DFF \creg_reg[363]  ( .D(n13989), .CLK(clk), .RST(rst), .Q(creg[363]) );
  DFF \creg_reg[364]  ( .D(n13988), .CLK(clk), .RST(rst), .Q(creg[364]) );
  DFF \creg_reg[365]  ( .D(n13987), .CLK(clk), .RST(rst), .Q(creg[365]) );
  DFF \creg_reg[366]  ( .D(n13986), .CLK(clk), .RST(rst), .Q(creg[366]) );
  DFF \creg_reg[367]  ( .D(n13985), .CLK(clk), .RST(rst), .Q(creg[367]) );
  DFF \creg_reg[368]  ( .D(n13984), .CLK(clk), .RST(rst), .Q(creg[368]) );
  DFF \creg_reg[369]  ( .D(n13983), .CLK(clk), .RST(rst), .Q(creg[369]) );
  DFF \creg_reg[370]  ( .D(n13982), .CLK(clk), .RST(rst), .Q(creg[370]) );
  DFF \creg_reg[371]  ( .D(n13981), .CLK(clk), .RST(rst), .Q(creg[371]) );
  DFF \creg_reg[372]  ( .D(n13980), .CLK(clk), .RST(rst), .Q(creg[372]) );
  DFF \creg_reg[373]  ( .D(n13979), .CLK(clk), .RST(rst), .Q(creg[373]) );
  DFF \creg_reg[374]  ( .D(n13978), .CLK(clk), .RST(rst), .Q(creg[374]) );
  DFF \creg_reg[375]  ( .D(n13977), .CLK(clk), .RST(rst), .Q(creg[375]) );
  DFF \creg_reg[376]  ( .D(n13976), .CLK(clk), .RST(rst), .Q(creg[376]) );
  DFF \creg_reg[377]  ( .D(n13975), .CLK(clk), .RST(rst), .Q(creg[377]) );
  DFF \creg_reg[378]  ( .D(n13974), .CLK(clk), .RST(rst), .Q(creg[378]) );
  DFF \creg_reg[379]  ( .D(n13973), .CLK(clk), .RST(rst), .Q(creg[379]) );
  DFF \creg_reg[380]  ( .D(n13972), .CLK(clk), .RST(rst), .Q(creg[380]) );
  DFF \creg_reg[381]  ( .D(n13971), .CLK(clk), .RST(rst), .Q(creg[381]) );
  DFF \creg_reg[382]  ( .D(n13970), .CLK(clk), .RST(rst), .Q(creg[382]) );
  DFF \creg_reg[383]  ( .D(n13969), .CLK(clk), .RST(rst), .Q(creg[383]) );
  DFF \creg_reg[384]  ( .D(n13968), .CLK(clk), .RST(rst), .Q(creg[384]) );
  DFF \creg_reg[385]  ( .D(n13967), .CLK(clk), .RST(rst), .Q(creg[385]) );
  DFF \creg_reg[386]  ( .D(n13966), .CLK(clk), .RST(rst), .Q(creg[386]) );
  DFF \creg_reg[387]  ( .D(n13965), .CLK(clk), .RST(rst), .Q(creg[387]) );
  DFF \creg_reg[388]  ( .D(n13964), .CLK(clk), .RST(rst), .Q(creg[388]) );
  DFF \creg_reg[389]  ( .D(n13963), .CLK(clk), .RST(rst), .Q(creg[389]) );
  DFF \creg_reg[390]  ( .D(n13962), .CLK(clk), .RST(rst), .Q(creg[390]) );
  DFF \creg_reg[391]  ( .D(n13961), .CLK(clk), .RST(rst), .Q(creg[391]) );
  DFF \creg_reg[392]  ( .D(n13960), .CLK(clk), .RST(rst), .Q(creg[392]) );
  DFF \creg_reg[393]  ( .D(n13959), .CLK(clk), .RST(rst), .Q(creg[393]) );
  DFF \creg_reg[394]  ( .D(n13958), .CLK(clk), .RST(rst), .Q(creg[394]) );
  DFF \creg_reg[395]  ( .D(n13957), .CLK(clk), .RST(rst), .Q(creg[395]) );
  DFF \creg_reg[396]  ( .D(n13956), .CLK(clk), .RST(rst), .Q(creg[396]) );
  DFF \creg_reg[397]  ( .D(n13955), .CLK(clk), .RST(rst), .Q(creg[397]) );
  DFF \creg_reg[398]  ( .D(n13954), .CLK(clk), .RST(rst), .Q(creg[398]) );
  DFF \creg_reg[399]  ( .D(n13953), .CLK(clk), .RST(rst), .Q(creg[399]) );
  DFF \creg_reg[400]  ( .D(n13952), .CLK(clk), .RST(rst), .Q(creg[400]) );
  DFF \creg_reg[401]  ( .D(n13951), .CLK(clk), .RST(rst), .Q(creg[401]) );
  DFF \creg_reg[402]  ( .D(n13950), .CLK(clk), .RST(rst), .Q(creg[402]) );
  DFF \creg_reg[403]  ( .D(n13949), .CLK(clk), .RST(rst), .Q(creg[403]) );
  DFF \creg_reg[404]  ( .D(n13948), .CLK(clk), .RST(rst), .Q(creg[404]) );
  DFF \creg_reg[405]  ( .D(n13947), .CLK(clk), .RST(rst), .Q(creg[405]) );
  DFF \creg_reg[406]  ( .D(n13946), .CLK(clk), .RST(rst), .Q(creg[406]) );
  DFF \creg_reg[407]  ( .D(n13945), .CLK(clk), .RST(rst), .Q(creg[407]) );
  DFF \creg_reg[408]  ( .D(n13944), .CLK(clk), .RST(rst), .Q(creg[408]) );
  DFF \creg_reg[409]  ( .D(n13943), .CLK(clk), .RST(rst), .Q(creg[409]) );
  DFF \creg_reg[410]  ( .D(n13942), .CLK(clk), .RST(rst), .Q(creg[410]) );
  DFF \creg_reg[411]  ( .D(n13941), .CLK(clk), .RST(rst), .Q(creg[411]) );
  DFF \creg_reg[412]  ( .D(n13940), .CLK(clk), .RST(rst), .Q(creg[412]) );
  DFF \creg_reg[413]  ( .D(n13939), .CLK(clk), .RST(rst), .Q(creg[413]) );
  DFF \creg_reg[414]  ( .D(n13938), .CLK(clk), .RST(rst), .Q(creg[414]) );
  DFF \creg_reg[415]  ( .D(n13937), .CLK(clk), .RST(rst), .Q(creg[415]) );
  DFF \creg_reg[416]  ( .D(n13936), .CLK(clk), .RST(rst), .Q(creg[416]) );
  DFF \creg_reg[417]  ( .D(n13935), .CLK(clk), .RST(rst), .Q(creg[417]) );
  DFF \creg_reg[418]  ( .D(n13934), .CLK(clk), .RST(rst), .Q(creg[418]) );
  DFF \creg_reg[419]  ( .D(n13933), .CLK(clk), .RST(rst), .Q(creg[419]) );
  DFF \creg_reg[420]  ( .D(n13932), .CLK(clk), .RST(rst), .Q(creg[420]) );
  DFF \creg_reg[421]  ( .D(n13931), .CLK(clk), .RST(rst), .Q(creg[421]) );
  DFF \creg_reg[422]  ( .D(n13930), .CLK(clk), .RST(rst), .Q(creg[422]) );
  DFF \creg_reg[423]  ( .D(n13929), .CLK(clk), .RST(rst), .Q(creg[423]) );
  DFF \creg_reg[424]  ( .D(n13928), .CLK(clk), .RST(rst), .Q(creg[424]) );
  DFF \creg_reg[425]  ( .D(n13927), .CLK(clk), .RST(rst), .Q(creg[425]) );
  DFF \creg_reg[426]  ( .D(n13926), .CLK(clk), .RST(rst), .Q(creg[426]) );
  DFF \creg_reg[427]  ( .D(n13925), .CLK(clk), .RST(rst), .Q(creg[427]) );
  DFF \creg_reg[428]  ( .D(n13924), .CLK(clk), .RST(rst), .Q(creg[428]) );
  DFF \creg_reg[429]  ( .D(n13923), .CLK(clk), .RST(rst), .Q(creg[429]) );
  DFF \creg_reg[430]  ( .D(n13922), .CLK(clk), .RST(rst), .Q(creg[430]) );
  DFF \creg_reg[431]  ( .D(n13921), .CLK(clk), .RST(rst), .Q(creg[431]) );
  DFF \creg_reg[432]  ( .D(n13920), .CLK(clk), .RST(rst), .Q(creg[432]) );
  DFF \creg_reg[433]  ( .D(n13919), .CLK(clk), .RST(rst), .Q(creg[433]) );
  DFF \creg_reg[434]  ( .D(n13918), .CLK(clk), .RST(rst), .Q(creg[434]) );
  DFF \creg_reg[435]  ( .D(n13917), .CLK(clk), .RST(rst), .Q(creg[435]) );
  DFF \creg_reg[436]  ( .D(n13916), .CLK(clk), .RST(rst), .Q(creg[436]) );
  DFF \creg_reg[437]  ( .D(n13915), .CLK(clk), .RST(rst), .Q(creg[437]) );
  DFF \creg_reg[438]  ( .D(n13914), .CLK(clk), .RST(rst), .Q(creg[438]) );
  DFF \creg_reg[439]  ( .D(n13913), .CLK(clk), .RST(rst), .Q(creg[439]) );
  DFF \creg_reg[440]  ( .D(n13912), .CLK(clk), .RST(rst), .Q(creg[440]) );
  DFF \creg_reg[441]  ( .D(n13911), .CLK(clk), .RST(rst), .Q(creg[441]) );
  DFF \creg_reg[442]  ( .D(n13910), .CLK(clk), .RST(rst), .Q(creg[442]) );
  DFF \creg_reg[443]  ( .D(n13909), .CLK(clk), .RST(rst), .Q(creg[443]) );
  DFF \creg_reg[444]  ( .D(n13908), .CLK(clk), .RST(rst), .Q(creg[444]) );
  DFF \creg_reg[445]  ( .D(n13907), .CLK(clk), .RST(rst), .Q(creg[445]) );
  DFF \creg_reg[446]  ( .D(n13906), .CLK(clk), .RST(rst), .Q(creg[446]) );
  DFF \creg_reg[447]  ( .D(n13905), .CLK(clk), .RST(rst), .Q(creg[447]) );
  DFF \creg_reg[448]  ( .D(n13904), .CLK(clk), .RST(rst), .Q(creg[448]) );
  DFF \creg_reg[449]  ( .D(n13903), .CLK(clk), .RST(rst), .Q(creg[449]) );
  DFF \creg_reg[450]  ( .D(n13902), .CLK(clk), .RST(rst), .Q(creg[450]) );
  DFF \creg_reg[451]  ( .D(n13901), .CLK(clk), .RST(rst), .Q(creg[451]) );
  DFF \creg_reg[452]  ( .D(n13900), .CLK(clk), .RST(rst), .Q(creg[452]) );
  DFF \creg_reg[453]  ( .D(n13899), .CLK(clk), .RST(rst), .Q(creg[453]) );
  DFF \creg_reg[454]  ( .D(n13898), .CLK(clk), .RST(rst), .Q(creg[454]) );
  DFF \creg_reg[455]  ( .D(n13897), .CLK(clk), .RST(rst), .Q(creg[455]) );
  DFF \creg_reg[456]  ( .D(n13896), .CLK(clk), .RST(rst), .Q(creg[456]) );
  DFF \creg_reg[457]  ( .D(n13895), .CLK(clk), .RST(rst), .Q(creg[457]) );
  DFF \creg_reg[458]  ( .D(n13894), .CLK(clk), .RST(rst), .Q(creg[458]) );
  DFF \creg_reg[459]  ( .D(n13893), .CLK(clk), .RST(rst), .Q(creg[459]) );
  DFF \creg_reg[460]  ( .D(n13892), .CLK(clk), .RST(rst), .Q(creg[460]) );
  DFF \creg_reg[461]  ( .D(n13891), .CLK(clk), .RST(rst), .Q(creg[461]) );
  DFF \creg_reg[462]  ( .D(n13890), .CLK(clk), .RST(rst), .Q(creg[462]) );
  DFF \creg_reg[463]  ( .D(n13889), .CLK(clk), .RST(rst), .Q(creg[463]) );
  DFF \creg_reg[464]  ( .D(n13888), .CLK(clk), .RST(rst), .Q(creg[464]) );
  DFF \creg_reg[465]  ( .D(n13887), .CLK(clk), .RST(rst), .Q(creg[465]) );
  DFF \creg_reg[466]  ( .D(n13886), .CLK(clk), .RST(rst), .Q(creg[466]) );
  DFF \creg_reg[467]  ( .D(n13885), .CLK(clk), .RST(rst), .Q(creg[467]) );
  DFF \creg_reg[468]  ( .D(n13884), .CLK(clk), .RST(rst), .Q(creg[468]) );
  DFF \creg_reg[469]  ( .D(n13883), .CLK(clk), .RST(rst), .Q(creg[469]) );
  DFF \creg_reg[470]  ( .D(n13882), .CLK(clk), .RST(rst), .Q(creg[470]) );
  DFF \creg_reg[471]  ( .D(n13881), .CLK(clk), .RST(rst), .Q(creg[471]) );
  DFF \creg_reg[472]  ( .D(n13880), .CLK(clk), .RST(rst), .Q(creg[472]) );
  DFF \creg_reg[473]  ( .D(n13879), .CLK(clk), .RST(rst), .Q(creg[473]) );
  DFF \creg_reg[474]  ( .D(n13878), .CLK(clk), .RST(rst), .Q(creg[474]) );
  DFF \creg_reg[475]  ( .D(n13877), .CLK(clk), .RST(rst), .Q(creg[475]) );
  DFF \creg_reg[476]  ( .D(n13876), .CLK(clk), .RST(rst), .Q(creg[476]) );
  DFF \creg_reg[477]  ( .D(n13875), .CLK(clk), .RST(rst), .Q(creg[477]) );
  DFF \creg_reg[478]  ( .D(n13874), .CLK(clk), .RST(rst), .Q(creg[478]) );
  DFF \creg_reg[479]  ( .D(n13873), .CLK(clk), .RST(rst), .Q(creg[479]) );
  DFF \creg_reg[480]  ( .D(n13872), .CLK(clk), .RST(rst), .Q(creg[480]) );
  DFF \creg_reg[481]  ( .D(n13871), .CLK(clk), .RST(rst), .Q(creg[481]) );
  DFF \creg_reg[482]  ( .D(n13870), .CLK(clk), .RST(rst), .Q(creg[482]) );
  DFF \creg_reg[483]  ( .D(n13869), .CLK(clk), .RST(rst), .Q(creg[483]) );
  DFF \creg_reg[484]  ( .D(n13868), .CLK(clk), .RST(rst), .Q(creg[484]) );
  DFF \creg_reg[485]  ( .D(n13867), .CLK(clk), .RST(rst), .Q(creg[485]) );
  DFF \creg_reg[486]  ( .D(n13866), .CLK(clk), .RST(rst), .Q(creg[486]) );
  DFF \creg_reg[487]  ( .D(n13865), .CLK(clk), .RST(rst), .Q(creg[487]) );
  DFF \creg_reg[488]  ( .D(n13864), .CLK(clk), .RST(rst), .Q(creg[488]) );
  DFF \creg_reg[489]  ( .D(n13863), .CLK(clk), .RST(rst), .Q(creg[489]) );
  DFF \creg_reg[490]  ( .D(n13862), .CLK(clk), .RST(rst), .Q(creg[490]) );
  DFF \creg_reg[491]  ( .D(n13861), .CLK(clk), .RST(rst), .Q(creg[491]) );
  DFF \creg_reg[492]  ( .D(n13860), .CLK(clk), .RST(rst), .Q(creg[492]) );
  DFF \creg_reg[493]  ( .D(n13859), .CLK(clk), .RST(rst), .Q(creg[493]) );
  DFF \creg_reg[494]  ( .D(n13858), .CLK(clk), .RST(rst), .Q(creg[494]) );
  DFF \creg_reg[495]  ( .D(n13857), .CLK(clk), .RST(rst), .Q(creg[495]) );
  DFF \creg_reg[496]  ( .D(n13856), .CLK(clk), .RST(rst), .Q(creg[496]) );
  DFF \creg_reg[497]  ( .D(n13855), .CLK(clk), .RST(rst), .Q(creg[497]) );
  DFF \creg_reg[498]  ( .D(n13854), .CLK(clk), .RST(rst), .Q(creg[498]) );
  DFF \creg_reg[499]  ( .D(n13853), .CLK(clk), .RST(rst), .Q(creg[499]) );
  DFF \creg_reg[500]  ( .D(n13852), .CLK(clk), .RST(rst), .Q(creg[500]) );
  DFF \creg_reg[501]  ( .D(n13851), .CLK(clk), .RST(rst), .Q(creg[501]) );
  DFF \creg_reg[502]  ( .D(n13850), .CLK(clk), .RST(rst), .Q(creg[502]) );
  DFF \creg_reg[503]  ( .D(n13849), .CLK(clk), .RST(rst), .Q(creg[503]) );
  DFF \creg_reg[504]  ( .D(n13848), .CLK(clk), .RST(rst), .Q(creg[504]) );
  DFF \creg_reg[505]  ( .D(n13847), .CLK(clk), .RST(rst), .Q(creg[505]) );
  DFF \creg_reg[506]  ( .D(n13846), .CLK(clk), .RST(rst), .Q(creg[506]) );
  DFF \creg_reg[507]  ( .D(n13845), .CLK(clk), .RST(rst), .Q(creg[507]) );
  DFF \creg_reg[508]  ( .D(n13844), .CLK(clk), .RST(rst), .Q(creg[508]) );
  DFF \creg_reg[509]  ( .D(n13843), .CLK(clk), .RST(rst), .Q(creg[509]) );
  DFF \creg_reg[510]  ( .D(n13842), .CLK(clk), .RST(rst), .Q(creg[510]) );
  DFF \creg_reg[511]  ( .D(n13841), .CLK(clk), .RST(rst), .Q(creg[511]) );
  DFF \creg_reg[512]  ( .D(n13840), .CLK(clk), .RST(rst), .Q(creg[512]) );
  DFF \creg_reg[513]  ( .D(n13839), .CLK(clk), .RST(rst), .Q(creg[513]) );
  DFF \creg_reg[514]  ( .D(n13838), .CLK(clk), .RST(rst), .Q(creg[514]) );
  DFF \creg_reg[515]  ( .D(n13837), .CLK(clk), .RST(rst), .Q(creg[515]) );
  DFF \creg_reg[516]  ( .D(n13836), .CLK(clk), .RST(rst), .Q(creg[516]) );
  DFF \creg_reg[517]  ( .D(n13835), .CLK(clk), .RST(rst), .Q(creg[517]) );
  DFF \creg_reg[518]  ( .D(n13834), .CLK(clk), .RST(rst), .Q(creg[518]) );
  DFF \creg_reg[519]  ( .D(n13833), .CLK(clk), .RST(rst), .Q(creg[519]) );
  DFF \creg_reg[520]  ( .D(n13832), .CLK(clk), .RST(rst), .Q(creg[520]) );
  DFF \creg_reg[521]  ( .D(n13831), .CLK(clk), .RST(rst), .Q(creg[521]) );
  DFF \creg_reg[522]  ( .D(n13830), .CLK(clk), .RST(rst), .Q(creg[522]) );
  DFF \creg_reg[523]  ( .D(n13829), .CLK(clk), .RST(rst), .Q(creg[523]) );
  DFF \creg_reg[524]  ( .D(n13828), .CLK(clk), .RST(rst), .Q(creg[524]) );
  DFF \creg_reg[525]  ( .D(n13827), .CLK(clk), .RST(rst), .Q(creg[525]) );
  DFF \creg_reg[526]  ( .D(n13826), .CLK(clk), .RST(rst), .Q(creg[526]) );
  DFF \creg_reg[527]  ( .D(n13825), .CLK(clk), .RST(rst), .Q(creg[527]) );
  DFF \creg_reg[528]  ( .D(n13824), .CLK(clk), .RST(rst), .Q(creg[528]) );
  DFF \creg_reg[529]  ( .D(n13823), .CLK(clk), .RST(rst), .Q(creg[529]) );
  DFF \creg_reg[530]  ( .D(n13822), .CLK(clk), .RST(rst), .Q(creg[530]) );
  DFF \creg_reg[531]  ( .D(n13821), .CLK(clk), .RST(rst), .Q(creg[531]) );
  DFF \creg_reg[532]  ( .D(n13820), .CLK(clk), .RST(rst), .Q(creg[532]) );
  DFF \creg_reg[533]  ( .D(n13819), .CLK(clk), .RST(rst), .Q(creg[533]) );
  DFF \creg_reg[534]  ( .D(n13818), .CLK(clk), .RST(rst), .Q(creg[534]) );
  DFF \creg_reg[535]  ( .D(n13817), .CLK(clk), .RST(rst), .Q(creg[535]) );
  DFF \creg_reg[536]  ( .D(n13816), .CLK(clk), .RST(rst), .Q(creg[536]) );
  DFF \creg_reg[537]  ( .D(n13815), .CLK(clk), .RST(rst), .Q(creg[537]) );
  DFF \creg_reg[538]  ( .D(n13814), .CLK(clk), .RST(rst), .Q(creg[538]) );
  DFF \creg_reg[539]  ( .D(n13813), .CLK(clk), .RST(rst), .Q(creg[539]) );
  DFF \creg_reg[540]  ( .D(n13812), .CLK(clk), .RST(rst), .Q(creg[540]) );
  DFF \creg_reg[541]  ( .D(n13811), .CLK(clk), .RST(rst), .Q(creg[541]) );
  DFF \creg_reg[542]  ( .D(n13810), .CLK(clk), .RST(rst), .Q(creg[542]) );
  DFF \creg_reg[543]  ( .D(n13809), .CLK(clk), .RST(rst), .Q(creg[543]) );
  DFF \creg_reg[544]  ( .D(n13808), .CLK(clk), .RST(rst), .Q(creg[544]) );
  DFF \creg_reg[545]  ( .D(n13807), .CLK(clk), .RST(rst), .Q(creg[545]) );
  DFF \creg_reg[546]  ( .D(n13806), .CLK(clk), .RST(rst), .Q(creg[546]) );
  DFF \creg_reg[547]  ( .D(n13805), .CLK(clk), .RST(rst), .Q(creg[547]) );
  DFF \creg_reg[548]  ( .D(n13804), .CLK(clk), .RST(rst), .Q(creg[548]) );
  DFF \creg_reg[549]  ( .D(n13803), .CLK(clk), .RST(rst), .Q(creg[549]) );
  DFF \creg_reg[550]  ( .D(n13802), .CLK(clk), .RST(rst), .Q(creg[550]) );
  DFF \creg_reg[551]  ( .D(n13801), .CLK(clk), .RST(rst), .Q(creg[551]) );
  DFF \creg_reg[552]  ( .D(n13800), .CLK(clk), .RST(rst), .Q(creg[552]) );
  DFF \creg_reg[553]  ( .D(n13799), .CLK(clk), .RST(rst), .Q(creg[553]) );
  DFF \creg_reg[554]  ( .D(n13798), .CLK(clk), .RST(rst), .Q(creg[554]) );
  DFF \creg_reg[555]  ( .D(n13797), .CLK(clk), .RST(rst), .Q(creg[555]) );
  DFF \creg_reg[556]  ( .D(n13796), .CLK(clk), .RST(rst), .Q(creg[556]) );
  DFF \creg_reg[557]  ( .D(n13795), .CLK(clk), .RST(rst), .Q(creg[557]) );
  DFF \creg_reg[558]  ( .D(n13794), .CLK(clk), .RST(rst), .Q(creg[558]) );
  DFF \creg_reg[559]  ( .D(n13793), .CLK(clk), .RST(rst), .Q(creg[559]) );
  DFF \creg_reg[560]  ( .D(n13792), .CLK(clk), .RST(rst), .Q(creg[560]) );
  DFF \creg_reg[561]  ( .D(n13791), .CLK(clk), .RST(rst), .Q(creg[561]) );
  DFF \creg_reg[562]  ( .D(n13790), .CLK(clk), .RST(rst), .Q(creg[562]) );
  DFF \creg_reg[563]  ( .D(n13789), .CLK(clk), .RST(rst), .Q(creg[563]) );
  DFF \creg_reg[564]  ( .D(n13788), .CLK(clk), .RST(rst), .Q(creg[564]) );
  DFF \creg_reg[565]  ( .D(n13787), .CLK(clk), .RST(rst), .Q(creg[565]) );
  DFF \creg_reg[566]  ( .D(n13786), .CLK(clk), .RST(rst), .Q(creg[566]) );
  DFF \creg_reg[567]  ( .D(n13785), .CLK(clk), .RST(rst), .Q(creg[567]) );
  DFF \creg_reg[568]  ( .D(n13784), .CLK(clk), .RST(rst), .Q(creg[568]) );
  DFF \creg_reg[569]  ( .D(n13783), .CLK(clk), .RST(rst), .Q(creg[569]) );
  DFF \creg_reg[570]  ( .D(n13782), .CLK(clk), .RST(rst), .Q(creg[570]) );
  DFF \creg_reg[571]  ( .D(n13781), .CLK(clk), .RST(rst), .Q(creg[571]) );
  DFF \creg_reg[572]  ( .D(n13780), .CLK(clk), .RST(rst), .Q(creg[572]) );
  DFF \creg_reg[573]  ( .D(n13779), .CLK(clk), .RST(rst), .Q(creg[573]) );
  DFF \creg_reg[574]  ( .D(n13778), .CLK(clk), .RST(rst), .Q(creg[574]) );
  DFF \creg_reg[575]  ( .D(n13777), .CLK(clk), .RST(rst), .Q(creg[575]) );
  DFF \creg_reg[576]  ( .D(n13776), .CLK(clk), .RST(rst), .Q(creg[576]) );
  DFF \creg_reg[577]  ( .D(n13775), .CLK(clk), .RST(rst), .Q(creg[577]) );
  DFF \creg_reg[578]  ( .D(n13774), .CLK(clk), .RST(rst), .Q(creg[578]) );
  DFF \creg_reg[579]  ( .D(n13773), .CLK(clk), .RST(rst), .Q(creg[579]) );
  DFF \creg_reg[580]  ( .D(n13772), .CLK(clk), .RST(rst), .Q(creg[580]) );
  DFF \creg_reg[581]  ( .D(n13771), .CLK(clk), .RST(rst), .Q(creg[581]) );
  DFF \creg_reg[582]  ( .D(n13770), .CLK(clk), .RST(rst), .Q(creg[582]) );
  DFF \creg_reg[583]  ( .D(n13769), .CLK(clk), .RST(rst), .Q(creg[583]) );
  DFF \creg_reg[584]  ( .D(n13768), .CLK(clk), .RST(rst), .Q(creg[584]) );
  DFF \creg_reg[585]  ( .D(n13767), .CLK(clk), .RST(rst), .Q(creg[585]) );
  DFF \creg_reg[586]  ( .D(n13766), .CLK(clk), .RST(rst), .Q(creg[586]) );
  DFF \creg_reg[587]  ( .D(n13765), .CLK(clk), .RST(rst), .Q(creg[587]) );
  DFF \creg_reg[588]  ( .D(n13764), .CLK(clk), .RST(rst), .Q(creg[588]) );
  DFF \creg_reg[589]  ( .D(n13763), .CLK(clk), .RST(rst), .Q(creg[589]) );
  DFF \creg_reg[590]  ( .D(n13762), .CLK(clk), .RST(rst), .Q(creg[590]) );
  DFF \creg_reg[591]  ( .D(n13761), .CLK(clk), .RST(rst), .Q(creg[591]) );
  DFF \creg_reg[592]  ( .D(n13760), .CLK(clk), .RST(rst), .Q(creg[592]) );
  DFF \creg_reg[593]  ( .D(n13759), .CLK(clk), .RST(rst), .Q(creg[593]) );
  DFF \creg_reg[594]  ( .D(n13758), .CLK(clk), .RST(rst), .Q(creg[594]) );
  DFF \creg_reg[595]  ( .D(n13757), .CLK(clk), .RST(rst), .Q(creg[595]) );
  DFF \creg_reg[596]  ( .D(n13756), .CLK(clk), .RST(rst), .Q(creg[596]) );
  DFF \creg_reg[597]  ( .D(n13755), .CLK(clk), .RST(rst), .Q(creg[597]) );
  DFF \creg_reg[598]  ( .D(n13754), .CLK(clk), .RST(rst), .Q(creg[598]) );
  DFF \creg_reg[599]  ( .D(n13753), .CLK(clk), .RST(rst), .Q(creg[599]) );
  DFF \creg_reg[600]  ( .D(n13752), .CLK(clk), .RST(rst), .Q(creg[600]) );
  DFF \creg_reg[601]  ( .D(n13751), .CLK(clk), .RST(rst), .Q(creg[601]) );
  DFF \creg_reg[602]  ( .D(n13750), .CLK(clk), .RST(rst), .Q(creg[602]) );
  DFF \creg_reg[603]  ( .D(n13749), .CLK(clk), .RST(rst), .Q(creg[603]) );
  DFF \creg_reg[604]  ( .D(n13748), .CLK(clk), .RST(rst), .Q(creg[604]) );
  DFF \creg_reg[605]  ( .D(n13747), .CLK(clk), .RST(rst), .Q(creg[605]) );
  DFF \creg_reg[606]  ( .D(n13746), .CLK(clk), .RST(rst), .Q(creg[606]) );
  DFF \creg_reg[607]  ( .D(n13745), .CLK(clk), .RST(rst), .Q(creg[607]) );
  DFF \creg_reg[608]  ( .D(n13744), .CLK(clk), .RST(rst), .Q(creg[608]) );
  DFF \creg_reg[609]  ( .D(n13743), .CLK(clk), .RST(rst), .Q(creg[609]) );
  DFF \creg_reg[610]  ( .D(n13742), .CLK(clk), .RST(rst), .Q(creg[610]) );
  DFF \creg_reg[611]  ( .D(n13741), .CLK(clk), .RST(rst), .Q(creg[611]) );
  DFF \creg_reg[612]  ( .D(n13740), .CLK(clk), .RST(rst), .Q(creg[612]) );
  DFF \creg_reg[613]  ( .D(n13739), .CLK(clk), .RST(rst), .Q(creg[613]) );
  DFF \creg_reg[614]  ( .D(n13738), .CLK(clk), .RST(rst), .Q(creg[614]) );
  DFF \creg_reg[615]  ( .D(n13737), .CLK(clk), .RST(rst), .Q(creg[615]) );
  DFF \creg_reg[616]  ( .D(n13736), .CLK(clk), .RST(rst), .Q(creg[616]) );
  DFF \creg_reg[617]  ( .D(n13735), .CLK(clk), .RST(rst), .Q(creg[617]) );
  DFF \creg_reg[618]  ( .D(n13734), .CLK(clk), .RST(rst), .Q(creg[618]) );
  DFF \creg_reg[619]  ( .D(n13733), .CLK(clk), .RST(rst), .Q(creg[619]) );
  DFF \creg_reg[620]  ( .D(n13732), .CLK(clk), .RST(rst), .Q(creg[620]) );
  DFF \creg_reg[621]  ( .D(n13731), .CLK(clk), .RST(rst), .Q(creg[621]) );
  DFF \creg_reg[622]  ( .D(n13730), .CLK(clk), .RST(rst), .Q(creg[622]) );
  DFF \creg_reg[623]  ( .D(n13729), .CLK(clk), .RST(rst), .Q(creg[623]) );
  DFF \creg_reg[624]  ( .D(n13728), .CLK(clk), .RST(rst), .Q(creg[624]) );
  DFF \creg_reg[625]  ( .D(n13727), .CLK(clk), .RST(rst), .Q(creg[625]) );
  DFF \creg_reg[626]  ( .D(n13726), .CLK(clk), .RST(rst), .Q(creg[626]) );
  DFF \creg_reg[627]  ( .D(n13725), .CLK(clk), .RST(rst), .Q(creg[627]) );
  DFF \creg_reg[628]  ( .D(n13724), .CLK(clk), .RST(rst), .Q(creg[628]) );
  DFF \creg_reg[629]  ( .D(n13723), .CLK(clk), .RST(rst), .Q(creg[629]) );
  DFF \creg_reg[630]  ( .D(n13722), .CLK(clk), .RST(rst), .Q(creg[630]) );
  DFF \creg_reg[631]  ( .D(n13721), .CLK(clk), .RST(rst), .Q(creg[631]) );
  DFF \creg_reg[632]  ( .D(n13720), .CLK(clk), .RST(rst), .Q(creg[632]) );
  DFF \creg_reg[633]  ( .D(n13719), .CLK(clk), .RST(rst), .Q(creg[633]) );
  DFF \creg_reg[634]  ( .D(n13718), .CLK(clk), .RST(rst), .Q(creg[634]) );
  DFF \creg_reg[635]  ( .D(n13717), .CLK(clk), .RST(rst), .Q(creg[635]) );
  DFF \creg_reg[636]  ( .D(n13716), .CLK(clk), .RST(rst), .Q(creg[636]) );
  DFF \creg_reg[637]  ( .D(n13715), .CLK(clk), .RST(rst), .Q(creg[637]) );
  DFF \creg_reg[638]  ( .D(n13714), .CLK(clk), .RST(rst), .Q(creg[638]) );
  DFF \creg_reg[639]  ( .D(n13713), .CLK(clk), .RST(rst), .Q(creg[639]) );
  DFF \creg_reg[640]  ( .D(n13712), .CLK(clk), .RST(rst), .Q(creg[640]) );
  DFF \creg_reg[641]  ( .D(n13711), .CLK(clk), .RST(rst), .Q(creg[641]) );
  DFF \creg_reg[642]  ( .D(n13710), .CLK(clk), .RST(rst), .Q(creg[642]) );
  DFF \creg_reg[643]  ( .D(n13709), .CLK(clk), .RST(rst), .Q(creg[643]) );
  DFF \creg_reg[644]  ( .D(n13708), .CLK(clk), .RST(rst), .Q(creg[644]) );
  DFF \creg_reg[645]  ( .D(n13707), .CLK(clk), .RST(rst), .Q(creg[645]) );
  DFF \creg_reg[646]  ( .D(n13706), .CLK(clk), .RST(rst), .Q(creg[646]) );
  DFF \creg_reg[647]  ( .D(n13705), .CLK(clk), .RST(rst), .Q(creg[647]) );
  DFF \creg_reg[648]  ( .D(n13704), .CLK(clk), .RST(rst), .Q(creg[648]) );
  DFF \creg_reg[649]  ( .D(n13703), .CLK(clk), .RST(rst), .Q(creg[649]) );
  DFF \creg_reg[650]  ( .D(n13702), .CLK(clk), .RST(rst), .Q(creg[650]) );
  DFF \creg_reg[651]  ( .D(n13701), .CLK(clk), .RST(rst), .Q(creg[651]) );
  DFF \creg_reg[652]  ( .D(n13700), .CLK(clk), .RST(rst), .Q(creg[652]) );
  DFF \creg_reg[653]  ( .D(n13699), .CLK(clk), .RST(rst), .Q(creg[653]) );
  DFF \creg_reg[654]  ( .D(n13698), .CLK(clk), .RST(rst), .Q(creg[654]) );
  DFF \creg_reg[655]  ( .D(n13697), .CLK(clk), .RST(rst), .Q(creg[655]) );
  DFF \creg_reg[656]  ( .D(n13696), .CLK(clk), .RST(rst), .Q(creg[656]) );
  DFF \creg_reg[657]  ( .D(n13695), .CLK(clk), .RST(rst), .Q(creg[657]) );
  DFF \creg_reg[658]  ( .D(n13694), .CLK(clk), .RST(rst), .Q(creg[658]) );
  DFF \creg_reg[659]  ( .D(n13693), .CLK(clk), .RST(rst), .Q(creg[659]) );
  DFF \creg_reg[660]  ( .D(n13692), .CLK(clk), .RST(rst), .Q(creg[660]) );
  DFF \creg_reg[661]  ( .D(n13691), .CLK(clk), .RST(rst), .Q(creg[661]) );
  DFF \creg_reg[662]  ( .D(n13690), .CLK(clk), .RST(rst), .Q(creg[662]) );
  DFF \creg_reg[663]  ( .D(n13689), .CLK(clk), .RST(rst), .Q(creg[663]) );
  DFF \creg_reg[664]  ( .D(n13688), .CLK(clk), .RST(rst), .Q(creg[664]) );
  DFF \creg_reg[665]  ( .D(n13687), .CLK(clk), .RST(rst), .Q(creg[665]) );
  DFF \creg_reg[666]  ( .D(n13686), .CLK(clk), .RST(rst), .Q(creg[666]) );
  DFF \creg_reg[667]  ( .D(n13685), .CLK(clk), .RST(rst), .Q(creg[667]) );
  DFF \creg_reg[668]  ( .D(n13684), .CLK(clk), .RST(rst), .Q(creg[668]) );
  DFF \creg_reg[669]  ( .D(n13683), .CLK(clk), .RST(rst), .Q(creg[669]) );
  DFF \creg_reg[670]  ( .D(n13682), .CLK(clk), .RST(rst), .Q(creg[670]) );
  DFF \creg_reg[671]  ( .D(n13681), .CLK(clk), .RST(rst), .Q(creg[671]) );
  DFF \creg_reg[672]  ( .D(n13680), .CLK(clk), .RST(rst), .Q(creg[672]) );
  DFF \creg_reg[673]  ( .D(n13679), .CLK(clk), .RST(rst), .Q(creg[673]) );
  DFF \creg_reg[674]  ( .D(n13678), .CLK(clk), .RST(rst), .Q(creg[674]) );
  DFF \creg_reg[675]  ( .D(n13677), .CLK(clk), .RST(rst), .Q(creg[675]) );
  DFF \creg_reg[676]  ( .D(n13676), .CLK(clk), .RST(rst), .Q(creg[676]) );
  DFF \creg_reg[677]  ( .D(n13675), .CLK(clk), .RST(rst), .Q(creg[677]) );
  DFF \creg_reg[678]  ( .D(n13674), .CLK(clk), .RST(rst), .Q(creg[678]) );
  DFF \creg_reg[679]  ( .D(n13673), .CLK(clk), .RST(rst), .Q(creg[679]) );
  DFF \creg_reg[680]  ( .D(n13672), .CLK(clk), .RST(rst), .Q(creg[680]) );
  DFF \creg_reg[681]  ( .D(n13671), .CLK(clk), .RST(rst), .Q(creg[681]) );
  DFF \creg_reg[682]  ( .D(n13670), .CLK(clk), .RST(rst), .Q(creg[682]) );
  DFF \creg_reg[683]  ( .D(n13669), .CLK(clk), .RST(rst), .Q(creg[683]) );
  DFF \creg_reg[684]  ( .D(n13668), .CLK(clk), .RST(rst), .Q(creg[684]) );
  DFF \creg_reg[685]  ( .D(n13667), .CLK(clk), .RST(rst), .Q(creg[685]) );
  DFF \creg_reg[686]  ( .D(n13666), .CLK(clk), .RST(rst), .Q(creg[686]) );
  DFF \creg_reg[687]  ( .D(n13665), .CLK(clk), .RST(rst), .Q(creg[687]) );
  DFF \creg_reg[688]  ( .D(n13664), .CLK(clk), .RST(rst), .Q(creg[688]) );
  DFF \creg_reg[689]  ( .D(n13663), .CLK(clk), .RST(rst), .Q(creg[689]) );
  DFF \creg_reg[690]  ( .D(n13662), .CLK(clk), .RST(rst), .Q(creg[690]) );
  DFF \creg_reg[691]  ( .D(n13661), .CLK(clk), .RST(rst), .Q(creg[691]) );
  DFF \creg_reg[692]  ( .D(n13660), .CLK(clk), .RST(rst), .Q(creg[692]) );
  DFF \creg_reg[693]  ( .D(n13659), .CLK(clk), .RST(rst), .Q(creg[693]) );
  DFF \creg_reg[694]  ( .D(n13658), .CLK(clk), .RST(rst), .Q(creg[694]) );
  DFF \creg_reg[695]  ( .D(n13657), .CLK(clk), .RST(rst), .Q(creg[695]) );
  DFF \creg_reg[696]  ( .D(n13656), .CLK(clk), .RST(rst), .Q(creg[696]) );
  DFF \creg_reg[697]  ( .D(n13655), .CLK(clk), .RST(rst), .Q(creg[697]) );
  DFF \creg_reg[698]  ( .D(n13654), .CLK(clk), .RST(rst), .Q(creg[698]) );
  DFF \creg_reg[699]  ( .D(n13653), .CLK(clk), .RST(rst), .Q(creg[699]) );
  DFF \creg_reg[700]  ( .D(n13652), .CLK(clk), .RST(rst), .Q(creg[700]) );
  DFF \creg_reg[701]  ( .D(n13651), .CLK(clk), .RST(rst), .Q(creg[701]) );
  DFF \creg_reg[702]  ( .D(n13650), .CLK(clk), .RST(rst), .Q(creg[702]) );
  DFF \creg_reg[703]  ( .D(n13649), .CLK(clk), .RST(rst), .Q(creg[703]) );
  DFF \creg_reg[704]  ( .D(n13648), .CLK(clk), .RST(rst), .Q(creg[704]) );
  DFF \creg_reg[705]  ( .D(n13647), .CLK(clk), .RST(rst), .Q(creg[705]) );
  DFF \creg_reg[706]  ( .D(n13646), .CLK(clk), .RST(rst), .Q(creg[706]) );
  DFF \creg_reg[707]  ( .D(n13645), .CLK(clk), .RST(rst), .Q(creg[707]) );
  DFF \creg_reg[708]  ( .D(n13644), .CLK(clk), .RST(rst), .Q(creg[708]) );
  DFF \creg_reg[709]  ( .D(n13643), .CLK(clk), .RST(rst), .Q(creg[709]) );
  DFF \creg_reg[710]  ( .D(n13642), .CLK(clk), .RST(rst), .Q(creg[710]) );
  DFF \creg_reg[711]  ( .D(n13641), .CLK(clk), .RST(rst), .Q(creg[711]) );
  DFF \creg_reg[712]  ( .D(n13640), .CLK(clk), .RST(rst), .Q(creg[712]) );
  DFF \creg_reg[713]  ( .D(n13639), .CLK(clk), .RST(rst), .Q(creg[713]) );
  DFF \creg_reg[714]  ( .D(n13638), .CLK(clk), .RST(rst), .Q(creg[714]) );
  DFF \creg_reg[715]  ( .D(n13637), .CLK(clk), .RST(rst), .Q(creg[715]) );
  DFF \creg_reg[716]  ( .D(n13636), .CLK(clk), .RST(rst), .Q(creg[716]) );
  DFF \creg_reg[717]  ( .D(n13635), .CLK(clk), .RST(rst), .Q(creg[717]) );
  DFF \creg_reg[718]  ( .D(n13634), .CLK(clk), .RST(rst), .Q(creg[718]) );
  DFF \creg_reg[719]  ( .D(n13633), .CLK(clk), .RST(rst), .Q(creg[719]) );
  DFF \creg_reg[720]  ( .D(n13632), .CLK(clk), .RST(rst), .Q(creg[720]) );
  DFF \creg_reg[721]  ( .D(n13631), .CLK(clk), .RST(rst), .Q(creg[721]) );
  DFF \creg_reg[722]  ( .D(n13630), .CLK(clk), .RST(rst), .Q(creg[722]) );
  DFF \creg_reg[723]  ( .D(n13629), .CLK(clk), .RST(rst), .Q(creg[723]) );
  DFF \creg_reg[724]  ( .D(n13628), .CLK(clk), .RST(rst), .Q(creg[724]) );
  DFF \creg_reg[725]  ( .D(n13627), .CLK(clk), .RST(rst), .Q(creg[725]) );
  DFF \creg_reg[726]  ( .D(n13626), .CLK(clk), .RST(rst), .Q(creg[726]) );
  DFF \creg_reg[727]  ( .D(n13625), .CLK(clk), .RST(rst), .Q(creg[727]) );
  DFF \creg_reg[728]  ( .D(n13624), .CLK(clk), .RST(rst), .Q(creg[728]) );
  DFF \creg_reg[729]  ( .D(n13623), .CLK(clk), .RST(rst), .Q(creg[729]) );
  DFF \creg_reg[730]  ( .D(n13622), .CLK(clk), .RST(rst), .Q(creg[730]) );
  DFF \creg_reg[731]  ( .D(n13621), .CLK(clk), .RST(rst), .Q(creg[731]) );
  DFF \creg_reg[732]  ( .D(n13620), .CLK(clk), .RST(rst), .Q(creg[732]) );
  DFF \creg_reg[733]  ( .D(n13619), .CLK(clk), .RST(rst), .Q(creg[733]) );
  DFF \creg_reg[734]  ( .D(n13618), .CLK(clk), .RST(rst), .Q(creg[734]) );
  DFF \creg_reg[735]  ( .D(n13617), .CLK(clk), .RST(rst), .Q(creg[735]) );
  DFF \creg_reg[736]  ( .D(n13616), .CLK(clk), .RST(rst), .Q(creg[736]) );
  DFF \creg_reg[737]  ( .D(n13615), .CLK(clk), .RST(rst), .Q(creg[737]) );
  DFF \creg_reg[738]  ( .D(n13614), .CLK(clk), .RST(rst), .Q(creg[738]) );
  DFF \creg_reg[739]  ( .D(n13613), .CLK(clk), .RST(rst), .Q(creg[739]) );
  DFF \creg_reg[740]  ( .D(n13612), .CLK(clk), .RST(rst), .Q(creg[740]) );
  DFF \creg_reg[741]  ( .D(n13611), .CLK(clk), .RST(rst), .Q(creg[741]) );
  DFF \creg_reg[742]  ( .D(n13610), .CLK(clk), .RST(rst), .Q(creg[742]) );
  DFF \creg_reg[743]  ( .D(n13609), .CLK(clk), .RST(rst), .Q(creg[743]) );
  DFF \creg_reg[744]  ( .D(n13608), .CLK(clk), .RST(rst), .Q(creg[744]) );
  DFF \creg_reg[745]  ( .D(n13607), .CLK(clk), .RST(rst), .Q(creg[745]) );
  DFF \creg_reg[746]  ( .D(n13606), .CLK(clk), .RST(rst), .Q(creg[746]) );
  DFF \creg_reg[747]  ( .D(n13605), .CLK(clk), .RST(rst), .Q(creg[747]) );
  DFF \creg_reg[748]  ( .D(n13604), .CLK(clk), .RST(rst), .Q(creg[748]) );
  DFF \creg_reg[749]  ( .D(n13603), .CLK(clk), .RST(rst), .Q(creg[749]) );
  DFF \creg_reg[750]  ( .D(n13602), .CLK(clk), .RST(rst), .Q(creg[750]) );
  DFF \creg_reg[751]  ( .D(n13601), .CLK(clk), .RST(rst), .Q(creg[751]) );
  DFF \creg_reg[752]  ( .D(n13600), .CLK(clk), .RST(rst), .Q(creg[752]) );
  DFF \creg_reg[753]  ( .D(n13599), .CLK(clk), .RST(rst), .Q(creg[753]) );
  DFF \creg_reg[754]  ( .D(n13598), .CLK(clk), .RST(rst), .Q(creg[754]) );
  DFF \creg_reg[755]  ( .D(n13597), .CLK(clk), .RST(rst), .Q(creg[755]) );
  DFF \creg_reg[756]  ( .D(n13596), .CLK(clk), .RST(rst), .Q(creg[756]) );
  DFF \creg_reg[757]  ( .D(n13595), .CLK(clk), .RST(rst), .Q(creg[757]) );
  DFF \creg_reg[758]  ( .D(n13594), .CLK(clk), .RST(rst), .Q(creg[758]) );
  DFF \creg_reg[759]  ( .D(n13593), .CLK(clk), .RST(rst), .Q(creg[759]) );
  DFF \creg_reg[760]  ( .D(n13592), .CLK(clk), .RST(rst), .Q(creg[760]) );
  DFF \creg_reg[761]  ( .D(n13591), .CLK(clk), .RST(rst), .Q(creg[761]) );
  DFF \creg_reg[762]  ( .D(n13590), .CLK(clk), .RST(rst), .Q(creg[762]) );
  DFF \creg_reg[763]  ( .D(n13589), .CLK(clk), .RST(rst), .Q(creg[763]) );
  DFF \creg_reg[764]  ( .D(n13588), .CLK(clk), .RST(rst), .Q(creg[764]) );
  DFF \creg_reg[765]  ( .D(n13587), .CLK(clk), .RST(rst), .Q(creg[765]) );
  DFF \creg_reg[766]  ( .D(n13586), .CLK(clk), .RST(rst), .Q(creg[766]) );
  DFF \creg_reg[767]  ( .D(n13585), .CLK(clk), .RST(rst), .Q(creg[767]) );
  DFF \creg_reg[768]  ( .D(n13584), .CLK(clk), .RST(rst), .Q(creg[768]) );
  DFF \creg_reg[769]  ( .D(n13583), .CLK(clk), .RST(rst), .Q(creg[769]) );
  DFF \creg_reg[770]  ( .D(n13582), .CLK(clk), .RST(rst), .Q(creg[770]) );
  DFF \creg_reg[771]  ( .D(n13581), .CLK(clk), .RST(rst), .Q(creg[771]) );
  DFF \creg_reg[772]  ( .D(n13580), .CLK(clk), .RST(rst), .Q(creg[772]) );
  DFF \creg_reg[773]  ( .D(n13579), .CLK(clk), .RST(rst), .Q(creg[773]) );
  DFF \creg_reg[774]  ( .D(n13578), .CLK(clk), .RST(rst), .Q(creg[774]) );
  DFF \creg_reg[775]  ( .D(n13577), .CLK(clk), .RST(rst), .Q(creg[775]) );
  DFF \creg_reg[776]  ( .D(n13576), .CLK(clk), .RST(rst), .Q(creg[776]) );
  DFF \creg_reg[777]  ( .D(n13575), .CLK(clk), .RST(rst), .Q(creg[777]) );
  DFF \creg_reg[778]  ( .D(n13574), .CLK(clk), .RST(rst), .Q(creg[778]) );
  DFF \creg_reg[779]  ( .D(n13573), .CLK(clk), .RST(rst), .Q(creg[779]) );
  DFF \creg_reg[780]  ( .D(n13572), .CLK(clk), .RST(rst), .Q(creg[780]) );
  DFF \creg_reg[781]  ( .D(n13571), .CLK(clk), .RST(rst), .Q(creg[781]) );
  DFF \creg_reg[782]  ( .D(n13570), .CLK(clk), .RST(rst), .Q(creg[782]) );
  DFF \creg_reg[783]  ( .D(n13569), .CLK(clk), .RST(rst), .Q(creg[783]) );
  DFF \creg_reg[784]  ( .D(n13568), .CLK(clk), .RST(rst), .Q(creg[784]) );
  DFF \creg_reg[785]  ( .D(n13567), .CLK(clk), .RST(rst), .Q(creg[785]) );
  DFF \creg_reg[786]  ( .D(n13566), .CLK(clk), .RST(rst), .Q(creg[786]) );
  DFF \creg_reg[787]  ( .D(n13565), .CLK(clk), .RST(rst), .Q(creg[787]) );
  DFF \creg_reg[788]  ( .D(n13564), .CLK(clk), .RST(rst), .Q(creg[788]) );
  DFF \creg_reg[789]  ( .D(n13563), .CLK(clk), .RST(rst), .Q(creg[789]) );
  DFF \creg_reg[790]  ( .D(n13562), .CLK(clk), .RST(rst), .Q(creg[790]) );
  DFF \creg_reg[791]  ( .D(n13561), .CLK(clk), .RST(rst), .Q(creg[791]) );
  DFF \creg_reg[792]  ( .D(n13560), .CLK(clk), .RST(rst), .Q(creg[792]) );
  DFF \creg_reg[793]  ( .D(n13559), .CLK(clk), .RST(rst), .Q(creg[793]) );
  DFF \creg_reg[794]  ( .D(n13558), .CLK(clk), .RST(rst), .Q(creg[794]) );
  DFF \creg_reg[795]  ( .D(n13557), .CLK(clk), .RST(rst), .Q(creg[795]) );
  DFF \creg_reg[796]  ( .D(n13556), .CLK(clk), .RST(rst), .Q(creg[796]) );
  DFF \creg_reg[797]  ( .D(n13555), .CLK(clk), .RST(rst), .Q(creg[797]) );
  DFF \creg_reg[798]  ( .D(n13554), .CLK(clk), .RST(rst), .Q(creg[798]) );
  DFF \creg_reg[799]  ( .D(n13553), .CLK(clk), .RST(rst), .Q(creg[799]) );
  DFF \creg_reg[800]  ( .D(n13552), .CLK(clk), .RST(rst), .Q(creg[800]) );
  DFF \creg_reg[801]  ( .D(n13551), .CLK(clk), .RST(rst), .Q(creg[801]) );
  DFF \creg_reg[802]  ( .D(n13550), .CLK(clk), .RST(rst), .Q(creg[802]) );
  DFF \creg_reg[803]  ( .D(n13549), .CLK(clk), .RST(rst), .Q(creg[803]) );
  DFF \creg_reg[804]  ( .D(n13548), .CLK(clk), .RST(rst), .Q(creg[804]) );
  DFF \creg_reg[805]  ( .D(n13547), .CLK(clk), .RST(rst), .Q(creg[805]) );
  DFF \creg_reg[806]  ( .D(n13546), .CLK(clk), .RST(rst), .Q(creg[806]) );
  DFF \creg_reg[807]  ( .D(n13545), .CLK(clk), .RST(rst), .Q(creg[807]) );
  DFF \creg_reg[808]  ( .D(n13544), .CLK(clk), .RST(rst), .Q(creg[808]) );
  DFF \creg_reg[809]  ( .D(n13543), .CLK(clk), .RST(rst), .Q(creg[809]) );
  DFF \creg_reg[810]  ( .D(n13542), .CLK(clk), .RST(rst), .Q(creg[810]) );
  DFF \creg_reg[811]  ( .D(n13541), .CLK(clk), .RST(rst), .Q(creg[811]) );
  DFF \creg_reg[812]  ( .D(n13540), .CLK(clk), .RST(rst), .Q(creg[812]) );
  DFF \creg_reg[813]  ( .D(n13539), .CLK(clk), .RST(rst), .Q(creg[813]) );
  DFF \creg_reg[814]  ( .D(n13538), .CLK(clk), .RST(rst), .Q(creg[814]) );
  DFF \creg_reg[815]  ( .D(n13537), .CLK(clk), .RST(rst), .Q(creg[815]) );
  DFF \creg_reg[816]  ( .D(n13536), .CLK(clk), .RST(rst), .Q(creg[816]) );
  DFF \creg_reg[817]  ( .D(n13535), .CLK(clk), .RST(rst), .Q(creg[817]) );
  DFF \creg_reg[818]  ( .D(n13534), .CLK(clk), .RST(rst), .Q(creg[818]) );
  DFF \creg_reg[819]  ( .D(n13533), .CLK(clk), .RST(rst), .Q(creg[819]) );
  DFF \creg_reg[820]  ( .D(n13532), .CLK(clk), .RST(rst), .Q(creg[820]) );
  DFF \creg_reg[821]  ( .D(n13531), .CLK(clk), .RST(rst), .Q(creg[821]) );
  DFF \creg_reg[822]  ( .D(n13530), .CLK(clk), .RST(rst), .Q(creg[822]) );
  DFF \creg_reg[823]  ( .D(n13529), .CLK(clk), .RST(rst), .Q(creg[823]) );
  DFF \creg_reg[824]  ( .D(n13528), .CLK(clk), .RST(rst), .Q(creg[824]) );
  DFF \creg_reg[825]  ( .D(n13527), .CLK(clk), .RST(rst), .Q(creg[825]) );
  DFF \creg_reg[826]  ( .D(n13526), .CLK(clk), .RST(rst), .Q(creg[826]) );
  DFF \creg_reg[827]  ( .D(n13525), .CLK(clk), .RST(rst), .Q(creg[827]) );
  DFF \creg_reg[828]  ( .D(n13524), .CLK(clk), .RST(rst), .Q(creg[828]) );
  DFF \creg_reg[829]  ( .D(n13523), .CLK(clk), .RST(rst), .Q(creg[829]) );
  DFF \creg_reg[830]  ( .D(n13522), .CLK(clk), .RST(rst), .Q(creg[830]) );
  DFF \creg_reg[831]  ( .D(n13521), .CLK(clk), .RST(rst), .Q(creg[831]) );
  DFF \creg_reg[832]  ( .D(n13520), .CLK(clk), .RST(rst), .Q(creg[832]) );
  DFF \creg_reg[833]  ( .D(n13519), .CLK(clk), .RST(rst), .Q(creg[833]) );
  DFF \creg_reg[834]  ( .D(n13518), .CLK(clk), .RST(rst), .Q(creg[834]) );
  DFF \creg_reg[835]  ( .D(n13517), .CLK(clk), .RST(rst), .Q(creg[835]) );
  DFF \creg_reg[836]  ( .D(n13516), .CLK(clk), .RST(rst), .Q(creg[836]) );
  DFF \creg_reg[837]  ( .D(n13515), .CLK(clk), .RST(rst), .Q(creg[837]) );
  DFF \creg_reg[838]  ( .D(n13514), .CLK(clk), .RST(rst), .Q(creg[838]) );
  DFF \creg_reg[839]  ( .D(n13513), .CLK(clk), .RST(rst), .Q(creg[839]) );
  DFF \creg_reg[840]  ( .D(n13512), .CLK(clk), .RST(rst), .Q(creg[840]) );
  DFF \creg_reg[841]  ( .D(n13511), .CLK(clk), .RST(rst), .Q(creg[841]) );
  DFF \creg_reg[842]  ( .D(n13510), .CLK(clk), .RST(rst), .Q(creg[842]) );
  DFF \creg_reg[843]  ( .D(n13509), .CLK(clk), .RST(rst), .Q(creg[843]) );
  DFF \creg_reg[844]  ( .D(n13508), .CLK(clk), .RST(rst), .Q(creg[844]) );
  DFF \creg_reg[845]  ( .D(n13507), .CLK(clk), .RST(rst), .Q(creg[845]) );
  DFF \creg_reg[846]  ( .D(n13506), .CLK(clk), .RST(rst), .Q(creg[846]) );
  DFF \creg_reg[847]  ( .D(n13505), .CLK(clk), .RST(rst), .Q(creg[847]) );
  DFF \creg_reg[848]  ( .D(n13504), .CLK(clk), .RST(rst), .Q(creg[848]) );
  DFF \creg_reg[849]  ( .D(n13503), .CLK(clk), .RST(rst), .Q(creg[849]) );
  DFF \creg_reg[850]  ( .D(n13502), .CLK(clk), .RST(rst), .Q(creg[850]) );
  DFF \creg_reg[851]  ( .D(n13501), .CLK(clk), .RST(rst), .Q(creg[851]) );
  DFF \creg_reg[852]  ( .D(n13500), .CLK(clk), .RST(rst), .Q(creg[852]) );
  DFF \creg_reg[853]  ( .D(n13499), .CLK(clk), .RST(rst), .Q(creg[853]) );
  DFF \creg_reg[854]  ( .D(n13498), .CLK(clk), .RST(rst), .Q(creg[854]) );
  DFF \creg_reg[855]  ( .D(n13497), .CLK(clk), .RST(rst), .Q(creg[855]) );
  DFF \creg_reg[856]  ( .D(n13496), .CLK(clk), .RST(rst), .Q(creg[856]) );
  DFF \creg_reg[857]  ( .D(n13495), .CLK(clk), .RST(rst), .Q(creg[857]) );
  DFF \creg_reg[858]  ( .D(n13494), .CLK(clk), .RST(rst), .Q(creg[858]) );
  DFF \creg_reg[859]  ( .D(n13493), .CLK(clk), .RST(rst), .Q(creg[859]) );
  DFF \creg_reg[860]  ( .D(n13492), .CLK(clk), .RST(rst), .Q(creg[860]) );
  DFF \creg_reg[861]  ( .D(n13491), .CLK(clk), .RST(rst), .Q(creg[861]) );
  DFF \creg_reg[862]  ( .D(n13490), .CLK(clk), .RST(rst), .Q(creg[862]) );
  DFF \creg_reg[863]  ( .D(n13489), .CLK(clk), .RST(rst), .Q(creg[863]) );
  DFF \creg_reg[864]  ( .D(n13488), .CLK(clk), .RST(rst), .Q(creg[864]) );
  DFF \creg_reg[865]  ( .D(n13487), .CLK(clk), .RST(rst), .Q(creg[865]) );
  DFF \creg_reg[866]  ( .D(n13486), .CLK(clk), .RST(rst), .Q(creg[866]) );
  DFF \creg_reg[867]  ( .D(n13485), .CLK(clk), .RST(rst), .Q(creg[867]) );
  DFF \creg_reg[868]  ( .D(n13484), .CLK(clk), .RST(rst), .Q(creg[868]) );
  DFF \creg_reg[869]  ( .D(n13483), .CLK(clk), .RST(rst), .Q(creg[869]) );
  DFF \creg_reg[870]  ( .D(n13482), .CLK(clk), .RST(rst), .Q(creg[870]) );
  DFF \creg_reg[871]  ( .D(n13481), .CLK(clk), .RST(rst), .Q(creg[871]) );
  DFF \creg_reg[872]  ( .D(n13480), .CLK(clk), .RST(rst), .Q(creg[872]) );
  DFF \creg_reg[873]  ( .D(n13479), .CLK(clk), .RST(rst), .Q(creg[873]) );
  DFF \creg_reg[874]  ( .D(n13478), .CLK(clk), .RST(rst), .Q(creg[874]) );
  DFF \creg_reg[875]  ( .D(n13477), .CLK(clk), .RST(rst), .Q(creg[875]) );
  DFF \creg_reg[876]  ( .D(n13476), .CLK(clk), .RST(rst), .Q(creg[876]) );
  DFF \creg_reg[877]  ( .D(n13475), .CLK(clk), .RST(rst), .Q(creg[877]) );
  DFF \creg_reg[878]  ( .D(n13474), .CLK(clk), .RST(rst), .Q(creg[878]) );
  DFF \creg_reg[879]  ( .D(n13473), .CLK(clk), .RST(rst), .Q(creg[879]) );
  DFF \creg_reg[880]  ( .D(n13472), .CLK(clk), .RST(rst), .Q(creg[880]) );
  DFF \creg_reg[881]  ( .D(n13471), .CLK(clk), .RST(rst), .Q(creg[881]) );
  DFF \creg_reg[882]  ( .D(n13470), .CLK(clk), .RST(rst), .Q(creg[882]) );
  DFF \creg_reg[883]  ( .D(n13469), .CLK(clk), .RST(rst), .Q(creg[883]) );
  DFF \creg_reg[884]  ( .D(n13468), .CLK(clk), .RST(rst), .Q(creg[884]) );
  DFF \creg_reg[885]  ( .D(n13467), .CLK(clk), .RST(rst), .Q(creg[885]) );
  DFF \creg_reg[886]  ( .D(n13466), .CLK(clk), .RST(rst), .Q(creg[886]) );
  DFF \creg_reg[887]  ( .D(n13465), .CLK(clk), .RST(rst), .Q(creg[887]) );
  DFF \creg_reg[888]  ( .D(n13464), .CLK(clk), .RST(rst), .Q(creg[888]) );
  DFF \creg_reg[889]  ( .D(n13463), .CLK(clk), .RST(rst), .Q(creg[889]) );
  DFF \creg_reg[890]  ( .D(n13462), .CLK(clk), .RST(rst), .Q(creg[890]) );
  DFF \creg_reg[891]  ( .D(n13461), .CLK(clk), .RST(rst), .Q(creg[891]) );
  DFF \creg_reg[892]  ( .D(n13460), .CLK(clk), .RST(rst), .Q(creg[892]) );
  DFF \creg_reg[893]  ( .D(n13459), .CLK(clk), .RST(rst), .Q(creg[893]) );
  DFF \creg_reg[894]  ( .D(n13458), .CLK(clk), .RST(rst), .Q(creg[894]) );
  DFF \creg_reg[895]  ( .D(n13457), .CLK(clk), .RST(rst), .Q(creg[895]) );
  DFF \creg_reg[896]  ( .D(n13456), .CLK(clk), .RST(rst), .Q(creg[896]) );
  DFF \creg_reg[897]  ( .D(n13455), .CLK(clk), .RST(rst), .Q(creg[897]) );
  DFF \creg_reg[898]  ( .D(n13454), .CLK(clk), .RST(rst), .Q(creg[898]) );
  DFF \creg_reg[899]  ( .D(n13453), .CLK(clk), .RST(rst), .Q(creg[899]) );
  DFF \creg_reg[900]  ( .D(n13452), .CLK(clk), .RST(rst), .Q(creg[900]) );
  DFF \creg_reg[901]  ( .D(n13451), .CLK(clk), .RST(rst), .Q(creg[901]) );
  DFF \creg_reg[902]  ( .D(n13450), .CLK(clk), .RST(rst), .Q(creg[902]) );
  DFF \creg_reg[903]  ( .D(n13449), .CLK(clk), .RST(rst), .Q(creg[903]) );
  DFF \creg_reg[904]  ( .D(n13448), .CLK(clk), .RST(rst), .Q(creg[904]) );
  DFF \creg_reg[905]  ( .D(n13447), .CLK(clk), .RST(rst), .Q(creg[905]) );
  DFF \creg_reg[906]  ( .D(n13446), .CLK(clk), .RST(rst), .Q(creg[906]) );
  DFF \creg_reg[907]  ( .D(n13445), .CLK(clk), .RST(rst), .Q(creg[907]) );
  DFF \creg_reg[908]  ( .D(n13444), .CLK(clk), .RST(rst), .Q(creg[908]) );
  DFF \creg_reg[909]  ( .D(n13443), .CLK(clk), .RST(rst), .Q(creg[909]) );
  DFF \creg_reg[910]  ( .D(n13442), .CLK(clk), .RST(rst), .Q(creg[910]) );
  DFF \creg_reg[911]  ( .D(n13441), .CLK(clk), .RST(rst), .Q(creg[911]) );
  DFF \creg_reg[912]  ( .D(n13440), .CLK(clk), .RST(rst), .Q(creg[912]) );
  DFF \creg_reg[913]  ( .D(n13439), .CLK(clk), .RST(rst), .Q(creg[913]) );
  DFF \creg_reg[914]  ( .D(n13438), .CLK(clk), .RST(rst), .Q(creg[914]) );
  DFF \creg_reg[915]  ( .D(n13437), .CLK(clk), .RST(rst), .Q(creg[915]) );
  DFF \creg_reg[916]  ( .D(n13436), .CLK(clk), .RST(rst), .Q(creg[916]) );
  DFF \creg_reg[917]  ( .D(n13435), .CLK(clk), .RST(rst), .Q(creg[917]) );
  DFF \creg_reg[918]  ( .D(n13434), .CLK(clk), .RST(rst), .Q(creg[918]) );
  DFF \creg_reg[919]  ( .D(n13433), .CLK(clk), .RST(rst), .Q(creg[919]) );
  DFF \creg_reg[920]  ( .D(n13432), .CLK(clk), .RST(rst), .Q(creg[920]) );
  DFF \creg_reg[921]  ( .D(n13431), .CLK(clk), .RST(rst), .Q(creg[921]) );
  DFF \creg_reg[922]  ( .D(n13430), .CLK(clk), .RST(rst), .Q(creg[922]) );
  DFF \creg_reg[923]  ( .D(n13429), .CLK(clk), .RST(rst), .Q(creg[923]) );
  DFF \creg_reg[924]  ( .D(n13428), .CLK(clk), .RST(rst), .Q(creg[924]) );
  DFF \creg_reg[925]  ( .D(n13427), .CLK(clk), .RST(rst), .Q(creg[925]) );
  DFF \creg_reg[926]  ( .D(n13426), .CLK(clk), .RST(rst), .Q(creg[926]) );
  DFF \creg_reg[927]  ( .D(n13425), .CLK(clk), .RST(rst), .Q(creg[927]) );
  DFF \creg_reg[928]  ( .D(n13424), .CLK(clk), .RST(rst), .Q(creg[928]) );
  DFF \creg_reg[929]  ( .D(n13423), .CLK(clk), .RST(rst), .Q(creg[929]) );
  DFF \creg_reg[930]  ( .D(n13422), .CLK(clk), .RST(rst), .Q(creg[930]) );
  DFF \creg_reg[931]  ( .D(n13421), .CLK(clk), .RST(rst), .Q(creg[931]) );
  DFF \creg_reg[932]  ( .D(n13420), .CLK(clk), .RST(rst), .Q(creg[932]) );
  DFF \creg_reg[933]  ( .D(n13419), .CLK(clk), .RST(rst), .Q(creg[933]) );
  DFF \creg_reg[934]  ( .D(n13418), .CLK(clk), .RST(rst), .Q(creg[934]) );
  DFF \creg_reg[935]  ( .D(n13417), .CLK(clk), .RST(rst), .Q(creg[935]) );
  DFF \creg_reg[936]  ( .D(n13416), .CLK(clk), .RST(rst), .Q(creg[936]) );
  DFF \creg_reg[937]  ( .D(n13415), .CLK(clk), .RST(rst), .Q(creg[937]) );
  DFF \creg_reg[938]  ( .D(n13414), .CLK(clk), .RST(rst), .Q(creg[938]) );
  DFF \creg_reg[939]  ( .D(n13413), .CLK(clk), .RST(rst), .Q(creg[939]) );
  DFF \creg_reg[940]  ( .D(n13412), .CLK(clk), .RST(rst), .Q(creg[940]) );
  DFF \creg_reg[941]  ( .D(n13411), .CLK(clk), .RST(rst), .Q(creg[941]) );
  DFF \creg_reg[942]  ( .D(n13410), .CLK(clk), .RST(rst), .Q(creg[942]) );
  DFF \creg_reg[943]  ( .D(n13409), .CLK(clk), .RST(rst), .Q(creg[943]) );
  DFF \creg_reg[944]  ( .D(n13408), .CLK(clk), .RST(rst), .Q(creg[944]) );
  DFF \creg_reg[945]  ( .D(n13407), .CLK(clk), .RST(rst), .Q(creg[945]) );
  DFF \creg_reg[946]  ( .D(n13406), .CLK(clk), .RST(rst), .Q(creg[946]) );
  DFF \creg_reg[947]  ( .D(n13405), .CLK(clk), .RST(rst), .Q(creg[947]) );
  DFF \creg_reg[948]  ( .D(n13404), .CLK(clk), .RST(rst), .Q(creg[948]) );
  DFF \creg_reg[949]  ( .D(n13403), .CLK(clk), .RST(rst), .Q(creg[949]) );
  DFF \creg_reg[950]  ( .D(n13402), .CLK(clk), .RST(rst), .Q(creg[950]) );
  DFF \creg_reg[951]  ( .D(n13401), .CLK(clk), .RST(rst), .Q(creg[951]) );
  DFF \creg_reg[952]  ( .D(n13400), .CLK(clk), .RST(rst), .Q(creg[952]) );
  DFF \creg_reg[953]  ( .D(n13399), .CLK(clk), .RST(rst), .Q(creg[953]) );
  DFF \creg_reg[954]  ( .D(n13398), .CLK(clk), .RST(rst), .Q(creg[954]) );
  DFF \creg_reg[955]  ( .D(n13397), .CLK(clk), .RST(rst), .Q(creg[955]) );
  DFF \creg_reg[956]  ( .D(n13396), .CLK(clk), .RST(rst), .Q(creg[956]) );
  DFF \creg_reg[957]  ( .D(n13395), .CLK(clk), .RST(rst), .Q(creg[957]) );
  DFF \creg_reg[958]  ( .D(n13394), .CLK(clk), .RST(rst), .Q(creg[958]) );
  DFF \creg_reg[959]  ( .D(n13393), .CLK(clk), .RST(rst), .Q(creg[959]) );
  DFF \creg_reg[960]  ( .D(n13392), .CLK(clk), .RST(rst), .Q(creg[960]) );
  DFF \creg_reg[961]  ( .D(n13391), .CLK(clk), .RST(rst), .Q(creg[961]) );
  DFF \creg_reg[962]  ( .D(n13390), .CLK(clk), .RST(rst), .Q(creg[962]) );
  DFF \creg_reg[963]  ( .D(n13389), .CLK(clk), .RST(rst), .Q(creg[963]) );
  DFF \creg_reg[964]  ( .D(n13388), .CLK(clk), .RST(rst), .Q(creg[964]) );
  DFF \creg_reg[965]  ( .D(n13387), .CLK(clk), .RST(rst), .Q(creg[965]) );
  DFF \creg_reg[966]  ( .D(n13386), .CLK(clk), .RST(rst), .Q(creg[966]) );
  DFF \creg_reg[967]  ( .D(n13385), .CLK(clk), .RST(rst), .Q(creg[967]) );
  DFF \creg_reg[968]  ( .D(n13384), .CLK(clk), .RST(rst), .Q(creg[968]) );
  DFF \creg_reg[969]  ( .D(n13383), .CLK(clk), .RST(rst), .Q(creg[969]) );
  DFF \creg_reg[970]  ( .D(n13382), .CLK(clk), .RST(rst), .Q(creg[970]) );
  DFF \creg_reg[971]  ( .D(n13381), .CLK(clk), .RST(rst), .Q(creg[971]) );
  DFF \creg_reg[972]  ( .D(n13380), .CLK(clk), .RST(rst), .Q(creg[972]) );
  DFF \creg_reg[973]  ( .D(n13379), .CLK(clk), .RST(rst), .Q(creg[973]) );
  DFF \creg_reg[974]  ( .D(n13378), .CLK(clk), .RST(rst), .Q(creg[974]) );
  DFF \creg_reg[975]  ( .D(n13377), .CLK(clk), .RST(rst), .Q(creg[975]) );
  DFF \creg_reg[976]  ( .D(n13376), .CLK(clk), .RST(rst), .Q(creg[976]) );
  DFF \creg_reg[977]  ( .D(n13375), .CLK(clk), .RST(rst), .Q(creg[977]) );
  DFF \creg_reg[978]  ( .D(n13374), .CLK(clk), .RST(rst), .Q(creg[978]) );
  DFF \creg_reg[979]  ( .D(n13373), .CLK(clk), .RST(rst), .Q(creg[979]) );
  DFF \creg_reg[980]  ( .D(n13372), .CLK(clk), .RST(rst), .Q(creg[980]) );
  DFF \creg_reg[981]  ( .D(n13371), .CLK(clk), .RST(rst), .Q(creg[981]) );
  DFF \creg_reg[982]  ( .D(n13370), .CLK(clk), .RST(rst), .Q(creg[982]) );
  DFF \creg_reg[983]  ( .D(n13369), .CLK(clk), .RST(rst), .Q(creg[983]) );
  DFF \creg_reg[984]  ( .D(n13368), .CLK(clk), .RST(rst), .Q(creg[984]) );
  DFF \creg_reg[985]  ( .D(n13367), .CLK(clk), .RST(rst), .Q(creg[985]) );
  DFF \creg_reg[986]  ( .D(n13366), .CLK(clk), .RST(rst), .Q(creg[986]) );
  DFF \creg_reg[987]  ( .D(n13365), .CLK(clk), .RST(rst), .Q(creg[987]) );
  DFF \creg_reg[988]  ( .D(n13364), .CLK(clk), .RST(rst), .Q(creg[988]) );
  DFF \creg_reg[989]  ( .D(n13363), .CLK(clk), .RST(rst), .Q(creg[989]) );
  DFF \creg_reg[990]  ( .D(n13362), .CLK(clk), .RST(rst), .Q(creg[990]) );
  DFF \creg_reg[991]  ( .D(n13361), .CLK(clk), .RST(rst), .Q(creg[991]) );
  DFF \creg_reg[992]  ( .D(n13360), .CLK(clk), .RST(rst), .Q(creg[992]) );
  DFF \creg_reg[993]  ( .D(n13359), .CLK(clk), .RST(rst), .Q(creg[993]) );
  DFF \creg_reg[994]  ( .D(n13358), .CLK(clk), .RST(rst), .Q(creg[994]) );
  DFF \creg_reg[995]  ( .D(n13357), .CLK(clk), .RST(rst), .Q(creg[995]) );
  DFF \creg_reg[996]  ( .D(n13356), .CLK(clk), .RST(rst), .Q(creg[996]) );
  DFF \creg_reg[997]  ( .D(n13355), .CLK(clk), .RST(rst), .Q(creg[997]) );
  DFF \creg_reg[998]  ( .D(n13354), .CLK(clk), .RST(rst), .Q(creg[998]) );
  DFF \creg_reg[999]  ( .D(n13353), .CLK(clk), .RST(rst), .Q(creg[999]) );
  DFF \creg_reg[1000]  ( .D(n13352), .CLK(clk), .RST(rst), .Q(creg[1000]) );
  DFF \creg_reg[1001]  ( .D(n13351), .CLK(clk), .RST(rst), .Q(creg[1001]) );
  DFF \creg_reg[1002]  ( .D(n13350), .CLK(clk), .RST(rst), .Q(creg[1002]) );
  DFF \creg_reg[1003]  ( .D(n13349), .CLK(clk), .RST(rst), .Q(creg[1003]) );
  DFF \creg_reg[1004]  ( .D(n13348), .CLK(clk), .RST(rst), .Q(creg[1004]) );
  DFF \creg_reg[1005]  ( .D(n13347), .CLK(clk), .RST(rst), .Q(creg[1005]) );
  DFF \creg_reg[1006]  ( .D(n13346), .CLK(clk), .RST(rst), .Q(creg[1006]) );
  DFF \creg_reg[1007]  ( .D(n13345), .CLK(clk), .RST(rst), .Q(creg[1007]) );
  DFF \creg_reg[1008]  ( .D(n13344), .CLK(clk), .RST(rst), .Q(creg[1008]) );
  DFF \creg_reg[1009]  ( .D(n13343), .CLK(clk), .RST(rst), .Q(creg[1009]) );
  DFF \creg_reg[1010]  ( .D(n13342), .CLK(clk), .RST(rst), .Q(creg[1010]) );
  DFF \creg_reg[1011]  ( .D(n13341), .CLK(clk), .RST(rst), .Q(creg[1011]) );
  DFF \creg_reg[1012]  ( .D(n13340), .CLK(clk), .RST(rst), .Q(creg[1012]) );
  DFF \creg_reg[1013]  ( .D(n13339), .CLK(clk), .RST(rst), .Q(creg[1013]) );
  DFF \creg_reg[1014]  ( .D(n13338), .CLK(clk), .RST(rst), .Q(creg[1014]) );
  DFF \creg_reg[1015]  ( .D(n13337), .CLK(clk), .RST(rst), .Q(creg[1015]) );
  DFF \creg_reg[1016]  ( .D(n13336), .CLK(clk), .RST(rst), .Q(creg[1016]) );
  DFF \creg_reg[1017]  ( .D(n13335), .CLK(clk), .RST(rst), .Q(creg[1017]) );
  DFF \creg_reg[1018]  ( .D(n13334), .CLK(clk), .RST(rst), .Q(creg[1018]) );
  DFF \creg_reg[1019]  ( .D(n13333), .CLK(clk), .RST(rst), .Q(creg[1019]) );
  DFF \creg_reg[1020]  ( .D(n13332), .CLK(clk), .RST(rst), .Q(creg[1020]) );
  DFF \creg_reg[1021]  ( .D(n13331), .CLK(clk), .RST(rst), .Q(creg[1021]) );
  DFF \creg_reg[1022]  ( .D(n13330), .CLK(clk), .RST(rst), .Q(creg[1022]) );
  DFF \creg_reg[1023]  ( .D(n14353), .CLK(clk), .RST(rst), .Q(creg[1023]) );
  modmult_N1024_CC1024 modmult_1 ( .clk(clk), .rst(rst), .start(start_in[0]), 
        .x(x), .y(y), .n(n), .o(o) );
  NAND U19477 ( .A(n15379), .B(n15380), .Z(y[9]) );
  NAND U19478 ( .A(n15381), .B(m[9]), .Z(n15380) );
  NAND U19479 ( .A(n15382), .B(creg[9]), .Z(n15379) );
  NAND U19480 ( .A(n15383), .B(n15384), .Z(y[99]) );
  NAND U19481 ( .A(n15381), .B(m[99]), .Z(n15384) );
  NAND U19482 ( .A(n15382), .B(creg[99]), .Z(n15383) );
  NAND U19483 ( .A(n15385), .B(n15386), .Z(y[999]) );
  NAND U19484 ( .A(n15381), .B(m[999]), .Z(n15386) );
  NAND U19485 ( .A(n15382), .B(creg[999]), .Z(n15385) );
  NAND U19486 ( .A(n15387), .B(n15388), .Z(y[998]) );
  NAND U19487 ( .A(n15381), .B(m[998]), .Z(n15388) );
  NAND U19488 ( .A(n15382), .B(creg[998]), .Z(n15387) );
  NAND U19489 ( .A(n15389), .B(n15390), .Z(y[997]) );
  NAND U19490 ( .A(n15381), .B(m[997]), .Z(n15390) );
  NAND U19491 ( .A(n15382), .B(creg[997]), .Z(n15389) );
  NAND U19492 ( .A(n15391), .B(n15392), .Z(y[996]) );
  NAND U19493 ( .A(n15381), .B(m[996]), .Z(n15392) );
  NAND U19494 ( .A(n15382), .B(creg[996]), .Z(n15391) );
  NAND U19495 ( .A(n15393), .B(n15394), .Z(y[995]) );
  NAND U19496 ( .A(n15381), .B(m[995]), .Z(n15394) );
  NAND U19497 ( .A(n15382), .B(creg[995]), .Z(n15393) );
  NAND U19498 ( .A(n15395), .B(n15396), .Z(y[994]) );
  NAND U19499 ( .A(n15381), .B(m[994]), .Z(n15396) );
  NAND U19500 ( .A(n15382), .B(creg[994]), .Z(n15395) );
  NAND U19501 ( .A(n15397), .B(n15398), .Z(y[993]) );
  NAND U19502 ( .A(n15381), .B(m[993]), .Z(n15398) );
  NAND U19503 ( .A(n15382), .B(creg[993]), .Z(n15397) );
  NAND U19504 ( .A(n15399), .B(n15400), .Z(y[992]) );
  NAND U19505 ( .A(n15381), .B(m[992]), .Z(n15400) );
  NAND U19506 ( .A(n15382), .B(creg[992]), .Z(n15399) );
  NAND U19507 ( .A(n15401), .B(n15402), .Z(y[991]) );
  NAND U19508 ( .A(n15381), .B(m[991]), .Z(n15402) );
  NAND U19509 ( .A(n15382), .B(creg[991]), .Z(n15401) );
  NAND U19510 ( .A(n15403), .B(n15404), .Z(y[990]) );
  NAND U19511 ( .A(n15381), .B(m[990]), .Z(n15404) );
  NAND U19512 ( .A(n15382), .B(creg[990]), .Z(n15403) );
  NAND U19513 ( .A(n15405), .B(n15406), .Z(y[98]) );
  NAND U19514 ( .A(n15381), .B(m[98]), .Z(n15406) );
  NAND U19515 ( .A(n15382), .B(creg[98]), .Z(n15405) );
  NAND U19516 ( .A(n15407), .B(n15408), .Z(y[989]) );
  NAND U19517 ( .A(n15381), .B(m[989]), .Z(n15408) );
  NAND U19518 ( .A(n15382), .B(creg[989]), .Z(n15407) );
  NAND U19519 ( .A(n15409), .B(n15410), .Z(y[988]) );
  NAND U19520 ( .A(n15381), .B(m[988]), .Z(n15410) );
  NAND U19521 ( .A(n15382), .B(creg[988]), .Z(n15409) );
  NAND U19522 ( .A(n15411), .B(n15412), .Z(y[987]) );
  NAND U19523 ( .A(n15381), .B(m[987]), .Z(n15412) );
  NAND U19524 ( .A(n15382), .B(creg[987]), .Z(n15411) );
  NAND U19525 ( .A(n15413), .B(n15414), .Z(y[986]) );
  NAND U19526 ( .A(n15381), .B(m[986]), .Z(n15414) );
  NAND U19527 ( .A(n15382), .B(creg[986]), .Z(n15413) );
  NAND U19528 ( .A(n15415), .B(n15416), .Z(y[985]) );
  NAND U19529 ( .A(n15381), .B(m[985]), .Z(n15416) );
  NAND U19530 ( .A(n15382), .B(creg[985]), .Z(n15415) );
  NAND U19531 ( .A(n15417), .B(n15418), .Z(y[984]) );
  NAND U19532 ( .A(n15381), .B(m[984]), .Z(n15418) );
  NAND U19533 ( .A(n15382), .B(creg[984]), .Z(n15417) );
  NAND U19534 ( .A(n15419), .B(n15420), .Z(y[983]) );
  NAND U19535 ( .A(n15381), .B(m[983]), .Z(n15420) );
  NAND U19536 ( .A(n15382), .B(creg[983]), .Z(n15419) );
  NAND U19537 ( .A(n15421), .B(n15422), .Z(y[982]) );
  NAND U19538 ( .A(n15381), .B(m[982]), .Z(n15422) );
  NAND U19539 ( .A(n15382), .B(creg[982]), .Z(n15421) );
  NAND U19540 ( .A(n15423), .B(n15424), .Z(y[981]) );
  NAND U19541 ( .A(n15381), .B(m[981]), .Z(n15424) );
  NAND U19542 ( .A(n15382), .B(creg[981]), .Z(n15423) );
  NAND U19543 ( .A(n15425), .B(n15426), .Z(y[980]) );
  NAND U19544 ( .A(n15381), .B(m[980]), .Z(n15426) );
  NAND U19545 ( .A(n15382), .B(creg[980]), .Z(n15425) );
  NAND U19546 ( .A(n15427), .B(n15428), .Z(y[97]) );
  NAND U19547 ( .A(n15381), .B(m[97]), .Z(n15428) );
  NAND U19548 ( .A(n15382), .B(creg[97]), .Z(n15427) );
  NAND U19549 ( .A(n15429), .B(n15430), .Z(y[979]) );
  NAND U19550 ( .A(n15381), .B(m[979]), .Z(n15430) );
  NAND U19551 ( .A(n15382), .B(creg[979]), .Z(n15429) );
  NAND U19552 ( .A(n15431), .B(n15432), .Z(y[978]) );
  NAND U19553 ( .A(n15381), .B(m[978]), .Z(n15432) );
  NAND U19554 ( .A(n15382), .B(creg[978]), .Z(n15431) );
  NAND U19555 ( .A(n15433), .B(n15434), .Z(y[977]) );
  NAND U19556 ( .A(n15381), .B(m[977]), .Z(n15434) );
  NAND U19557 ( .A(n15382), .B(creg[977]), .Z(n15433) );
  NAND U19558 ( .A(n15435), .B(n15436), .Z(y[976]) );
  NAND U19559 ( .A(n15381), .B(m[976]), .Z(n15436) );
  NAND U19560 ( .A(n15382), .B(creg[976]), .Z(n15435) );
  NAND U19561 ( .A(n15437), .B(n15438), .Z(y[975]) );
  NAND U19562 ( .A(n15381), .B(m[975]), .Z(n15438) );
  NAND U19563 ( .A(n15382), .B(creg[975]), .Z(n15437) );
  NAND U19564 ( .A(n15439), .B(n15440), .Z(y[974]) );
  NAND U19565 ( .A(n15381), .B(m[974]), .Z(n15440) );
  NAND U19566 ( .A(n15382), .B(creg[974]), .Z(n15439) );
  NAND U19567 ( .A(n15441), .B(n15442), .Z(y[973]) );
  NAND U19568 ( .A(n15381), .B(m[973]), .Z(n15442) );
  NAND U19569 ( .A(n15382), .B(creg[973]), .Z(n15441) );
  NAND U19570 ( .A(n15443), .B(n15444), .Z(y[972]) );
  NAND U19571 ( .A(n15381), .B(m[972]), .Z(n15444) );
  NAND U19572 ( .A(n15382), .B(creg[972]), .Z(n15443) );
  NAND U19573 ( .A(n15445), .B(n15446), .Z(y[971]) );
  NAND U19574 ( .A(n15381), .B(m[971]), .Z(n15446) );
  NAND U19575 ( .A(n15382), .B(creg[971]), .Z(n15445) );
  NAND U19576 ( .A(n15447), .B(n15448), .Z(y[970]) );
  NAND U19577 ( .A(n15381), .B(m[970]), .Z(n15448) );
  NAND U19578 ( .A(n15382), .B(creg[970]), .Z(n15447) );
  NAND U19579 ( .A(n15449), .B(n15450), .Z(y[96]) );
  NAND U19580 ( .A(n15381), .B(m[96]), .Z(n15450) );
  NAND U19581 ( .A(n15382), .B(creg[96]), .Z(n15449) );
  NAND U19582 ( .A(n15451), .B(n15452), .Z(y[969]) );
  NAND U19583 ( .A(n15381), .B(m[969]), .Z(n15452) );
  NAND U19584 ( .A(n15382), .B(creg[969]), .Z(n15451) );
  NAND U19585 ( .A(n15453), .B(n15454), .Z(y[968]) );
  NAND U19586 ( .A(n15381), .B(m[968]), .Z(n15454) );
  NAND U19587 ( .A(n15382), .B(creg[968]), .Z(n15453) );
  NAND U19588 ( .A(n15455), .B(n15456), .Z(y[967]) );
  NAND U19589 ( .A(n15381), .B(m[967]), .Z(n15456) );
  NAND U19590 ( .A(n15382), .B(creg[967]), .Z(n15455) );
  NAND U19591 ( .A(n15457), .B(n15458), .Z(y[966]) );
  NAND U19592 ( .A(n15381), .B(m[966]), .Z(n15458) );
  NAND U19593 ( .A(n15382), .B(creg[966]), .Z(n15457) );
  NAND U19594 ( .A(n15459), .B(n15460), .Z(y[965]) );
  NAND U19595 ( .A(n15381), .B(m[965]), .Z(n15460) );
  NAND U19596 ( .A(n15382), .B(creg[965]), .Z(n15459) );
  NAND U19597 ( .A(n15461), .B(n15462), .Z(y[964]) );
  NAND U19598 ( .A(n15381), .B(m[964]), .Z(n15462) );
  NAND U19599 ( .A(n15382), .B(creg[964]), .Z(n15461) );
  NAND U19600 ( .A(n15463), .B(n15464), .Z(y[963]) );
  NAND U19601 ( .A(n15381), .B(m[963]), .Z(n15464) );
  NAND U19602 ( .A(n15382), .B(creg[963]), .Z(n15463) );
  NAND U19603 ( .A(n15465), .B(n15466), .Z(y[962]) );
  NAND U19604 ( .A(n15381), .B(m[962]), .Z(n15466) );
  NAND U19605 ( .A(n15382), .B(creg[962]), .Z(n15465) );
  NAND U19606 ( .A(n15467), .B(n15468), .Z(y[961]) );
  NAND U19607 ( .A(n15381), .B(m[961]), .Z(n15468) );
  NAND U19608 ( .A(n15382), .B(creg[961]), .Z(n15467) );
  NAND U19609 ( .A(n15469), .B(n15470), .Z(y[960]) );
  NAND U19610 ( .A(n15381), .B(m[960]), .Z(n15470) );
  NAND U19611 ( .A(n15382), .B(creg[960]), .Z(n15469) );
  NAND U19612 ( .A(n15471), .B(n15472), .Z(y[95]) );
  NAND U19613 ( .A(n15381), .B(m[95]), .Z(n15472) );
  NAND U19614 ( .A(n15382), .B(creg[95]), .Z(n15471) );
  NAND U19615 ( .A(n15473), .B(n15474), .Z(y[959]) );
  NAND U19616 ( .A(n15381), .B(m[959]), .Z(n15474) );
  NAND U19617 ( .A(n15382), .B(creg[959]), .Z(n15473) );
  NAND U19618 ( .A(n15475), .B(n15476), .Z(y[958]) );
  NAND U19619 ( .A(n15381), .B(m[958]), .Z(n15476) );
  NAND U19620 ( .A(n15382), .B(creg[958]), .Z(n15475) );
  NAND U19621 ( .A(n15477), .B(n15478), .Z(y[957]) );
  NAND U19622 ( .A(n15381), .B(m[957]), .Z(n15478) );
  NAND U19623 ( .A(n15382), .B(creg[957]), .Z(n15477) );
  NAND U19624 ( .A(n15479), .B(n15480), .Z(y[956]) );
  NAND U19625 ( .A(n15381), .B(m[956]), .Z(n15480) );
  NAND U19626 ( .A(n15382), .B(creg[956]), .Z(n15479) );
  NAND U19627 ( .A(n15481), .B(n15482), .Z(y[955]) );
  NAND U19628 ( .A(n15381), .B(m[955]), .Z(n15482) );
  NAND U19629 ( .A(n15382), .B(creg[955]), .Z(n15481) );
  NAND U19630 ( .A(n15483), .B(n15484), .Z(y[954]) );
  NAND U19631 ( .A(n15381), .B(m[954]), .Z(n15484) );
  NAND U19632 ( .A(n15382), .B(creg[954]), .Z(n15483) );
  NAND U19633 ( .A(n15485), .B(n15486), .Z(y[953]) );
  NAND U19634 ( .A(n15381), .B(m[953]), .Z(n15486) );
  NAND U19635 ( .A(n15382), .B(creg[953]), .Z(n15485) );
  NAND U19636 ( .A(n15487), .B(n15488), .Z(y[952]) );
  NAND U19637 ( .A(n15381), .B(m[952]), .Z(n15488) );
  NAND U19638 ( .A(n15382), .B(creg[952]), .Z(n15487) );
  NAND U19639 ( .A(n15489), .B(n15490), .Z(y[951]) );
  NAND U19640 ( .A(n15381), .B(m[951]), .Z(n15490) );
  NAND U19641 ( .A(n15382), .B(creg[951]), .Z(n15489) );
  NAND U19642 ( .A(n15491), .B(n15492), .Z(y[950]) );
  NAND U19643 ( .A(n15381), .B(m[950]), .Z(n15492) );
  NAND U19644 ( .A(n15382), .B(creg[950]), .Z(n15491) );
  NAND U19645 ( .A(n15493), .B(n15494), .Z(y[94]) );
  NAND U19646 ( .A(n15381), .B(m[94]), .Z(n15494) );
  NAND U19647 ( .A(n15382), .B(creg[94]), .Z(n15493) );
  NAND U19648 ( .A(n15495), .B(n15496), .Z(y[949]) );
  NAND U19649 ( .A(n15381), .B(m[949]), .Z(n15496) );
  NAND U19650 ( .A(n15382), .B(creg[949]), .Z(n15495) );
  NAND U19651 ( .A(n15497), .B(n15498), .Z(y[948]) );
  NAND U19652 ( .A(n15381), .B(m[948]), .Z(n15498) );
  NAND U19653 ( .A(n15382), .B(creg[948]), .Z(n15497) );
  NAND U19654 ( .A(n15499), .B(n15500), .Z(y[947]) );
  NAND U19655 ( .A(n15381), .B(m[947]), .Z(n15500) );
  NAND U19656 ( .A(n15382), .B(creg[947]), .Z(n15499) );
  NAND U19657 ( .A(n15501), .B(n15502), .Z(y[946]) );
  NAND U19658 ( .A(n15381), .B(m[946]), .Z(n15502) );
  NAND U19659 ( .A(n15382), .B(creg[946]), .Z(n15501) );
  NAND U19660 ( .A(n15503), .B(n15504), .Z(y[945]) );
  NAND U19661 ( .A(n15381), .B(m[945]), .Z(n15504) );
  NAND U19662 ( .A(n15382), .B(creg[945]), .Z(n15503) );
  NAND U19663 ( .A(n15505), .B(n15506), .Z(y[944]) );
  NAND U19664 ( .A(n15381), .B(m[944]), .Z(n15506) );
  NAND U19665 ( .A(n15382), .B(creg[944]), .Z(n15505) );
  NAND U19666 ( .A(n15507), .B(n15508), .Z(y[943]) );
  NAND U19667 ( .A(n15381), .B(m[943]), .Z(n15508) );
  NAND U19668 ( .A(n15382), .B(creg[943]), .Z(n15507) );
  NAND U19669 ( .A(n15509), .B(n15510), .Z(y[942]) );
  NAND U19670 ( .A(n15381), .B(m[942]), .Z(n15510) );
  NAND U19671 ( .A(n15382), .B(creg[942]), .Z(n15509) );
  NAND U19672 ( .A(n15511), .B(n15512), .Z(y[941]) );
  NAND U19673 ( .A(n15381), .B(m[941]), .Z(n15512) );
  NAND U19674 ( .A(n15382), .B(creg[941]), .Z(n15511) );
  NAND U19675 ( .A(n15513), .B(n15514), .Z(y[940]) );
  NAND U19676 ( .A(n15381), .B(m[940]), .Z(n15514) );
  NAND U19677 ( .A(n15382), .B(creg[940]), .Z(n15513) );
  NAND U19678 ( .A(n15515), .B(n15516), .Z(y[93]) );
  NAND U19679 ( .A(n15381), .B(m[93]), .Z(n15516) );
  NAND U19680 ( .A(n15382), .B(creg[93]), .Z(n15515) );
  NAND U19681 ( .A(n15517), .B(n15518), .Z(y[939]) );
  NAND U19682 ( .A(n15381), .B(m[939]), .Z(n15518) );
  NAND U19683 ( .A(n15382), .B(creg[939]), .Z(n15517) );
  NAND U19684 ( .A(n15519), .B(n15520), .Z(y[938]) );
  NAND U19685 ( .A(n15381), .B(m[938]), .Z(n15520) );
  NAND U19686 ( .A(n15382), .B(creg[938]), .Z(n15519) );
  NAND U19687 ( .A(n15521), .B(n15522), .Z(y[937]) );
  NAND U19688 ( .A(n15381), .B(m[937]), .Z(n15522) );
  NAND U19689 ( .A(n15382), .B(creg[937]), .Z(n15521) );
  NAND U19690 ( .A(n15523), .B(n15524), .Z(y[936]) );
  NAND U19691 ( .A(n15381), .B(m[936]), .Z(n15524) );
  NAND U19692 ( .A(n15382), .B(creg[936]), .Z(n15523) );
  NAND U19693 ( .A(n15525), .B(n15526), .Z(y[935]) );
  NAND U19694 ( .A(n15381), .B(m[935]), .Z(n15526) );
  NAND U19695 ( .A(n15382), .B(creg[935]), .Z(n15525) );
  NAND U19696 ( .A(n15527), .B(n15528), .Z(y[934]) );
  NAND U19697 ( .A(n15381), .B(m[934]), .Z(n15528) );
  NAND U19698 ( .A(n15382), .B(creg[934]), .Z(n15527) );
  NAND U19699 ( .A(n15529), .B(n15530), .Z(y[933]) );
  NAND U19700 ( .A(n15381), .B(m[933]), .Z(n15530) );
  NAND U19701 ( .A(n15382), .B(creg[933]), .Z(n15529) );
  NAND U19702 ( .A(n15531), .B(n15532), .Z(y[932]) );
  NAND U19703 ( .A(n15381), .B(m[932]), .Z(n15532) );
  NAND U19704 ( .A(n15382), .B(creg[932]), .Z(n15531) );
  NAND U19705 ( .A(n15533), .B(n15534), .Z(y[931]) );
  NAND U19706 ( .A(n15381), .B(m[931]), .Z(n15534) );
  NAND U19707 ( .A(n15382), .B(creg[931]), .Z(n15533) );
  NAND U19708 ( .A(n15535), .B(n15536), .Z(y[930]) );
  NAND U19709 ( .A(n15381), .B(m[930]), .Z(n15536) );
  NAND U19710 ( .A(n15382), .B(creg[930]), .Z(n15535) );
  NAND U19711 ( .A(n15537), .B(n15538), .Z(y[92]) );
  NAND U19712 ( .A(n15381), .B(m[92]), .Z(n15538) );
  NAND U19713 ( .A(n15382), .B(creg[92]), .Z(n15537) );
  NAND U19714 ( .A(n15539), .B(n15540), .Z(y[929]) );
  NAND U19715 ( .A(n15381), .B(m[929]), .Z(n15540) );
  NAND U19716 ( .A(n15382), .B(creg[929]), .Z(n15539) );
  NAND U19717 ( .A(n15541), .B(n15542), .Z(y[928]) );
  NAND U19718 ( .A(n15381), .B(m[928]), .Z(n15542) );
  NAND U19719 ( .A(n15382), .B(creg[928]), .Z(n15541) );
  NAND U19720 ( .A(n15543), .B(n15544), .Z(y[927]) );
  NAND U19721 ( .A(n15381), .B(m[927]), .Z(n15544) );
  NAND U19722 ( .A(n15382), .B(creg[927]), .Z(n15543) );
  NAND U19723 ( .A(n15545), .B(n15546), .Z(y[926]) );
  NAND U19724 ( .A(n15381), .B(m[926]), .Z(n15546) );
  NAND U19725 ( .A(n15382), .B(creg[926]), .Z(n15545) );
  NAND U19726 ( .A(n15547), .B(n15548), .Z(y[925]) );
  NAND U19727 ( .A(n15381), .B(m[925]), .Z(n15548) );
  NAND U19728 ( .A(n15382), .B(creg[925]), .Z(n15547) );
  NAND U19729 ( .A(n15549), .B(n15550), .Z(y[924]) );
  NAND U19730 ( .A(n15381), .B(m[924]), .Z(n15550) );
  NAND U19731 ( .A(n15382), .B(creg[924]), .Z(n15549) );
  NAND U19732 ( .A(n15551), .B(n15552), .Z(y[923]) );
  NAND U19733 ( .A(n15381), .B(m[923]), .Z(n15552) );
  NAND U19734 ( .A(n15382), .B(creg[923]), .Z(n15551) );
  NAND U19735 ( .A(n15553), .B(n15554), .Z(y[922]) );
  NAND U19736 ( .A(n15381), .B(m[922]), .Z(n15554) );
  NAND U19737 ( .A(n15382), .B(creg[922]), .Z(n15553) );
  NAND U19738 ( .A(n15555), .B(n15556), .Z(y[921]) );
  NAND U19739 ( .A(n15381), .B(m[921]), .Z(n15556) );
  NAND U19740 ( .A(n15382), .B(creg[921]), .Z(n15555) );
  NAND U19741 ( .A(n15557), .B(n15558), .Z(y[920]) );
  NAND U19742 ( .A(n15381), .B(m[920]), .Z(n15558) );
  NAND U19743 ( .A(n15382), .B(creg[920]), .Z(n15557) );
  NAND U19744 ( .A(n15559), .B(n15560), .Z(y[91]) );
  NAND U19745 ( .A(n15381), .B(m[91]), .Z(n15560) );
  NAND U19746 ( .A(n15382), .B(creg[91]), .Z(n15559) );
  NAND U19747 ( .A(n15561), .B(n15562), .Z(y[919]) );
  NAND U19748 ( .A(n15381), .B(m[919]), .Z(n15562) );
  NAND U19749 ( .A(n15382), .B(creg[919]), .Z(n15561) );
  NAND U19750 ( .A(n15563), .B(n15564), .Z(y[918]) );
  NAND U19751 ( .A(n15381), .B(m[918]), .Z(n15564) );
  NAND U19752 ( .A(n15382), .B(creg[918]), .Z(n15563) );
  NAND U19753 ( .A(n15565), .B(n15566), .Z(y[917]) );
  NAND U19754 ( .A(n15381), .B(m[917]), .Z(n15566) );
  NAND U19755 ( .A(n15382), .B(creg[917]), .Z(n15565) );
  NAND U19756 ( .A(n15567), .B(n15568), .Z(y[916]) );
  NAND U19757 ( .A(n15381), .B(m[916]), .Z(n15568) );
  NAND U19758 ( .A(n15382), .B(creg[916]), .Z(n15567) );
  NAND U19759 ( .A(n15569), .B(n15570), .Z(y[915]) );
  NAND U19760 ( .A(n15381), .B(m[915]), .Z(n15570) );
  NAND U19761 ( .A(n15382), .B(creg[915]), .Z(n15569) );
  NAND U19762 ( .A(n15571), .B(n15572), .Z(y[914]) );
  NAND U19763 ( .A(n15381), .B(m[914]), .Z(n15572) );
  NAND U19764 ( .A(n15382), .B(creg[914]), .Z(n15571) );
  NAND U19765 ( .A(n15573), .B(n15574), .Z(y[913]) );
  NAND U19766 ( .A(n15381), .B(m[913]), .Z(n15574) );
  NAND U19767 ( .A(n15382), .B(creg[913]), .Z(n15573) );
  NAND U19768 ( .A(n15575), .B(n15576), .Z(y[912]) );
  NAND U19769 ( .A(n15381), .B(m[912]), .Z(n15576) );
  NAND U19770 ( .A(n15382), .B(creg[912]), .Z(n15575) );
  NAND U19771 ( .A(n15577), .B(n15578), .Z(y[911]) );
  NAND U19772 ( .A(n15381), .B(m[911]), .Z(n15578) );
  NAND U19773 ( .A(n15382), .B(creg[911]), .Z(n15577) );
  NAND U19774 ( .A(n15579), .B(n15580), .Z(y[910]) );
  NAND U19775 ( .A(n15381), .B(m[910]), .Z(n15580) );
  NAND U19776 ( .A(n15382), .B(creg[910]), .Z(n15579) );
  NAND U19777 ( .A(n15581), .B(n15582), .Z(y[90]) );
  NAND U19778 ( .A(n15381), .B(m[90]), .Z(n15582) );
  NAND U19779 ( .A(n15382), .B(creg[90]), .Z(n15581) );
  NAND U19780 ( .A(n15583), .B(n15584), .Z(y[909]) );
  NAND U19781 ( .A(n15381), .B(m[909]), .Z(n15584) );
  NAND U19782 ( .A(n15382), .B(creg[909]), .Z(n15583) );
  NAND U19783 ( .A(n15585), .B(n15586), .Z(y[908]) );
  NAND U19784 ( .A(n15381), .B(m[908]), .Z(n15586) );
  NAND U19785 ( .A(n15382), .B(creg[908]), .Z(n15585) );
  NAND U19786 ( .A(n15587), .B(n15588), .Z(y[907]) );
  NAND U19787 ( .A(n15381), .B(m[907]), .Z(n15588) );
  NAND U19788 ( .A(n15382), .B(creg[907]), .Z(n15587) );
  NAND U19789 ( .A(n15589), .B(n15590), .Z(y[906]) );
  NAND U19790 ( .A(n15381), .B(m[906]), .Z(n15590) );
  NAND U19791 ( .A(n15382), .B(creg[906]), .Z(n15589) );
  NAND U19792 ( .A(n15591), .B(n15592), .Z(y[905]) );
  NAND U19793 ( .A(n15381), .B(m[905]), .Z(n15592) );
  NAND U19794 ( .A(n15382), .B(creg[905]), .Z(n15591) );
  NAND U19795 ( .A(n15593), .B(n15594), .Z(y[904]) );
  NAND U19796 ( .A(n15381), .B(m[904]), .Z(n15594) );
  NAND U19797 ( .A(n15382), .B(creg[904]), .Z(n15593) );
  NAND U19798 ( .A(n15595), .B(n15596), .Z(y[903]) );
  NAND U19799 ( .A(n15381), .B(m[903]), .Z(n15596) );
  NAND U19800 ( .A(n15382), .B(creg[903]), .Z(n15595) );
  NAND U19801 ( .A(n15597), .B(n15598), .Z(y[902]) );
  NAND U19802 ( .A(n15381), .B(m[902]), .Z(n15598) );
  NAND U19803 ( .A(n15382), .B(creg[902]), .Z(n15597) );
  NAND U19804 ( .A(n15599), .B(n15600), .Z(y[901]) );
  NAND U19805 ( .A(n15381), .B(m[901]), .Z(n15600) );
  NAND U19806 ( .A(n15382), .B(creg[901]), .Z(n15599) );
  NAND U19807 ( .A(n15601), .B(n15602), .Z(y[900]) );
  NAND U19808 ( .A(n15381), .B(m[900]), .Z(n15602) );
  NAND U19809 ( .A(n15382), .B(creg[900]), .Z(n15601) );
  NAND U19810 ( .A(n15603), .B(n15604), .Z(y[8]) );
  NAND U19811 ( .A(n15381), .B(m[8]), .Z(n15604) );
  NAND U19812 ( .A(n15382), .B(creg[8]), .Z(n15603) );
  NAND U19813 ( .A(n15605), .B(n15606), .Z(y[89]) );
  NAND U19814 ( .A(n15381), .B(m[89]), .Z(n15606) );
  NAND U19815 ( .A(n15382), .B(creg[89]), .Z(n15605) );
  NAND U19816 ( .A(n15607), .B(n15608), .Z(y[899]) );
  NAND U19817 ( .A(n15381), .B(m[899]), .Z(n15608) );
  NAND U19818 ( .A(n15382), .B(creg[899]), .Z(n15607) );
  NAND U19819 ( .A(n15609), .B(n15610), .Z(y[898]) );
  NAND U19820 ( .A(n15381), .B(m[898]), .Z(n15610) );
  NAND U19821 ( .A(n15382), .B(creg[898]), .Z(n15609) );
  NAND U19822 ( .A(n15611), .B(n15612), .Z(y[897]) );
  NAND U19823 ( .A(n15381), .B(m[897]), .Z(n15612) );
  NAND U19824 ( .A(n15382), .B(creg[897]), .Z(n15611) );
  NAND U19825 ( .A(n15613), .B(n15614), .Z(y[896]) );
  NAND U19826 ( .A(n15381), .B(m[896]), .Z(n15614) );
  NAND U19827 ( .A(n15382), .B(creg[896]), .Z(n15613) );
  NAND U19828 ( .A(n15615), .B(n15616), .Z(y[895]) );
  NAND U19829 ( .A(n15381), .B(m[895]), .Z(n15616) );
  NAND U19830 ( .A(n15382), .B(creg[895]), .Z(n15615) );
  NAND U19831 ( .A(n15617), .B(n15618), .Z(y[894]) );
  NAND U19832 ( .A(n15381), .B(m[894]), .Z(n15618) );
  NAND U19833 ( .A(n15382), .B(creg[894]), .Z(n15617) );
  NAND U19834 ( .A(n15619), .B(n15620), .Z(y[893]) );
  NAND U19835 ( .A(n15381), .B(m[893]), .Z(n15620) );
  NAND U19836 ( .A(n15382), .B(creg[893]), .Z(n15619) );
  NAND U19837 ( .A(n15621), .B(n15622), .Z(y[892]) );
  NAND U19838 ( .A(n15381), .B(m[892]), .Z(n15622) );
  NAND U19839 ( .A(n15382), .B(creg[892]), .Z(n15621) );
  NAND U19840 ( .A(n15623), .B(n15624), .Z(y[891]) );
  NAND U19841 ( .A(n15381), .B(m[891]), .Z(n15624) );
  NAND U19842 ( .A(n15382), .B(creg[891]), .Z(n15623) );
  NAND U19843 ( .A(n15625), .B(n15626), .Z(y[890]) );
  NAND U19844 ( .A(n15381), .B(m[890]), .Z(n15626) );
  NAND U19845 ( .A(n15382), .B(creg[890]), .Z(n15625) );
  NAND U19846 ( .A(n15627), .B(n15628), .Z(y[88]) );
  NAND U19847 ( .A(n15381), .B(m[88]), .Z(n15628) );
  NAND U19848 ( .A(n15382), .B(creg[88]), .Z(n15627) );
  NAND U19849 ( .A(n15629), .B(n15630), .Z(y[889]) );
  NAND U19850 ( .A(n15381), .B(m[889]), .Z(n15630) );
  NAND U19851 ( .A(n15382), .B(creg[889]), .Z(n15629) );
  NAND U19852 ( .A(n15631), .B(n15632), .Z(y[888]) );
  NAND U19853 ( .A(n15381), .B(m[888]), .Z(n15632) );
  NAND U19854 ( .A(n15382), .B(creg[888]), .Z(n15631) );
  NAND U19855 ( .A(n15633), .B(n15634), .Z(y[887]) );
  NAND U19856 ( .A(n15381), .B(m[887]), .Z(n15634) );
  NAND U19857 ( .A(n15382), .B(creg[887]), .Z(n15633) );
  NAND U19858 ( .A(n15635), .B(n15636), .Z(y[886]) );
  NAND U19859 ( .A(n15381), .B(m[886]), .Z(n15636) );
  NAND U19860 ( .A(n15382), .B(creg[886]), .Z(n15635) );
  NAND U19861 ( .A(n15637), .B(n15638), .Z(y[885]) );
  NAND U19862 ( .A(n15381), .B(m[885]), .Z(n15638) );
  NAND U19863 ( .A(n15382), .B(creg[885]), .Z(n15637) );
  NAND U19864 ( .A(n15639), .B(n15640), .Z(y[884]) );
  NAND U19865 ( .A(n15381), .B(m[884]), .Z(n15640) );
  NAND U19866 ( .A(n15382), .B(creg[884]), .Z(n15639) );
  NAND U19867 ( .A(n15641), .B(n15642), .Z(y[883]) );
  NAND U19868 ( .A(n15381), .B(m[883]), .Z(n15642) );
  NAND U19869 ( .A(n15382), .B(creg[883]), .Z(n15641) );
  NAND U19870 ( .A(n15643), .B(n15644), .Z(y[882]) );
  NAND U19871 ( .A(n15381), .B(m[882]), .Z(n15644) );
  NAND U19872 ( .A(n15382), .B(creg[882]), .Z(n15643) );
  NAND U19873 ( .A(n15645), .B(n15646), .Z(y[881]) );
  NAND U19874 ( .A(n15381), .B(m[881]), .Z(n15646) );
  NAND U19875 ( .A(n15382), .B(creg[881]), .Z(n15645) );
  NAND U19876 ( .A(n15647), .B(n15648), .Z(y[880]) );
  NAND U19877 ( .A(n15381), .B(m[880]), .Z(n15648) );
  NAND U19878 ( .A(n15382), .B(creg[880]), .Z(n15647) );
  NAND U19879 ( .A(n15649), .B(n15650), .Z(y[87]) );
  NAND U19880 ( .A(n15381), .B(m[87]), .Z(n15650) );
  NAND U19881 ( .A(n15382), .B(creg[87]), .Z(n15649) );
  NAND U19882 ( .A(n15651), .B(n15652), .Z(y[879]) );
  NAND U19883 ( .A(n15381), .B(m[879]), .Z(n15652) );
  NAND U19884 ( .A(n15382), .B(creg[879]), .Z(n15651) );
  NAND U19885 ( .A(n15653), .B(n15654), .Z(y[878]) );
  NAND U19886 ( .A(n15381), .B(m[878]), .Z(n15654) );
  NAND U19887 ( .A(n15382), .B(creg[878]), .Z(n15653) );
  NAND U19888 ( .A(n15655), .B(n15656), .Z(y[877]) );
  NAND U19889 ( .A(n15381), .B(m[877]), .Z(n15656) );
  NAND U19890 ( .A(n15382), .B(creg[877]), .Z(n15655) );
  NAND U19891 ( .A(n15657), .B(n15658), .Z(y[876]) );
  NAND U19892 ( .A(n15381), .B(m[876]), .Z(n15658) );
  NAND U19893 ( .A(n15382), .B(creg[876]), .Z(n15657) );
  NAND U19894 ( .A(n15659), .B(n15660), .Z(y[875]) );
  NAND U19895 ( .A(n15381), .B(m[875]), .Z(n15660) );
  NAND U19896 ( .A(n15382), .B(creg[875]), .Z(n15659) );
  NAND U19897 ( .A(n15661), .B(n15662), .Z(y[874]) );
  NAND U19898 ( .A(n15381), .B(m[874]), .Z(n15662) );
  NAND U19899 ( .A(n15382), .B(creg[874]), .Z(n15661) );
  NAND U19900 ( .A(n15663), .B(n15664), .Z(y[873]) );
  NAND U19901 ( .A(n15381), .B(m[873]), .Z(n15664) );
  NAND U19902 ( .A(n15382), .B(creg[873]), .Z(n15663) );
  NAND U19903 ( .A(n15665), .B(n15666), .Z(y[872]) );
  NAND U19904 ( .A(n15381), .B(m[872]), .Z(n15666) );
  NAND U19905 ( .A(n15382), .B(creg[872]), .Z(n15665) );
  NAND U19906 ( .A(n15667), .B(n15668), .Z(y[871]) );
  NAND U19907 ( .A(n15381), .B(m[871]), .Z(n15668) );
  NAND U19908 ( .A(n15382), .B(creg[871]), .Z(n15667) );
  NAND U19909 ( .A(n15669), .B(n15670), .Z(y[870]) );
  NAND U19910 ( .A(n15381), .B(m[870]), .Z(n15670) );
  NAND U19911 ( .A(n15382), .B(creg[870]), .Z(n15669) );
  NAND U19912 ( .A(n15671), .B(n15672), .Z(y[86]) );
  NAND U19913 ( .A(n15381), .B(m[86]), .Z(n15672) );
  NAND U19914 ( .A(n15382), .B(creg[86]), .Z(n15671) );
  NAND U19915 ( .A(n15673), .B(n15674), .Z(y[869]) );
  NAND U19916 ( .A(n15381), .B(m[869]), .Z(n15674) );
  NAND U19917 ( .A(n15382), .B(creg[869]), .Z(n15673) );
  NAND U19918 ( .A(n15675), .B(n15676), .Z(y[868]) );
  NAND U19919 ( .A(n15381), .B(m[868]), .Z(n15676) );
  NAND U19920 ( .A(n15382), .B(creg[868]), .Z(n15675) );
  NAND U19921 ( .A(n15677), .B(n15678), .Z(y[867]) );
  NAND U19922 ( .A(n15381), .B(m[867]), .Z(n15678) );
  NAND U19923 ( .A(n15382), .B(creg[867]), .Z(n15677) );
  NAND U19924 ( .A(n15679), .B(n15680), .Z(y[866]) );
  NAND U19925 ( .A(n15381), .B(m[866]), .Z(n15680) );
  NAND U19926 ( .A(n15382), .B(creg[866]), .Z(n15679) );
  NAND U19927 ( .A(n15681), .B(n15682), .Z(y[865]) );
  NAND U19928 ( .A(n15381), .B(m[865]), .Z(n15682) );
  NAND U19929 ( .A(n15382), .B(creg[865]), .Z(n15681) );
  NAND U19930 ( .A(n15683), .B(n15684), .Z(y[864]) );
  NAND U19931 ( .A(n15381), .B(m[864]), .Z(n15684) );
  NAND U19932 ( .A(n15382), .B(creg[864]), .Z(n15683) );
  NAND U19933 ( .A(n15685), .B(n15686), .Z(y[863]) );
  NAND U19934 ( .A(n15381), .B(m[863]), .Z(n15686) );
  NAND U19935 ( .A(n15382), .B(creg[863]), .Z(n15685) );
  NAND U19936 ( .A(n15687), .B(n15688), .Z(y[862]) );
  NAND U19937 ( .A(n15381), .B(m[862]), .Z(n15688) );
  NAND U19938 ( .A(n15382), .B(creg[862]), .Z(n15687) );
  NAND U19939 ( .A(n15689), .B(n15690), .Z(y[861]) );
  NAND U19940 ( .A(n15381), .B(m[861]), .Z(n15690) );
  NAND U19941 ( .A(n15382), .B(creg[861]), .Z(n15689) );
  NAND U19942 ( .A(n15691), .B(n15692), .Z(y[860]) );
  NAND U19943 ( .A(n15381), .B(m[860]), .Z(n15692) );
  NAND U19944 ( .A(n15382), .B(creg[860]), .Z(n15691) );
  NAND U19945 ( .A(n15693), .B(n15694), .Z(y[85]) );
  NAND U19946 ( .A(n15381), .B(m[85]), .Z(n15694) );
  NAND U19947 ( .A(n15382), .B(creg[85]), .Z(n15693) );
  NAND U19948 ( .A(n15695), .B(n15696), .Z(y[859]) );
  NAND U19949 ( .A(n15381), .B(m[859]), .Z(n15696) );
  NAND U19950 ( .A(n15382), .B(creg[859]), .Z(n15695) );
  NAND U19951 ( .A(n15697), .B(n15698), .Z(y[858]) );
  NAND U19952 ( .A(n15381), .B(m[858]), .Z(n15698) );
  NAND U19953 ( .A(n15382), .B(creg[858]), .Z(n15697) );
  NAND U19954 ( .A(n15699), .B(n15700), .Z(y[857]) );
  NAND U19955 ( .A(n15381), .B(m[857]), .Z(n15700) );
  NAND U19956 ( .A(n15382), .B(creg[857]), .Z(n15699) );
  NAND U19957 ( .A(n15701), .B(n15702), .Z(y[856]) );
  NAND U19958 ( .A(n15381), .B(m[856]), .Z(n15702) );
  NAND U19959 ( .A(n15382), .B(creg[856]), .Z(n15701) );
  NAND U19960 ( .A(n15703), .B(n15704), .Z(y[855]) );
  NAND U19961 ( .A(n15381), .B(m[855]), .Z(n15704) );
  NAND U19962 ( .A(n15382), .B(creg[855]), .Z(n15703) );
  NAND U19963 ( .A(n15705), .B(n15706), .Z(y[854]) );
  NAND U19964 ( .A(n15381), .B(m[854]), .Z(n15706) );
  NAND U19965 ( .A(n15382), .B(creg[854]), .Z(n15705) );
  NAND U19966 ( .A(n15707), .B(n15708), .Z(y[853]) );
  NAND U19967 ( .A(n15381), .B(m[853]), .Z(n15708) );
  NAND U19968 ( .A(n15382), .B(creg[853]), .Z(n15707) );
  NAND U19969 ( .A(n15709), .B(n15710), .Z(y[852]) );
  NAND U19970 ( .A(n15381), .B(m[852]), .Z(n15710) );
  NAND U19971 ( .A(n15382), .B(creg[852]), .Z(n15709) );
  NAND U19972 ( .A(n15711), .B(n15712), .Z(y[851]) );
  NAND U19973 ( .A(n15381), .B(m[851]), .Z(n15712) );
  NAND U19974 ( .A(n15382), .B(creg[851]), .Z(n15711) );
  NAND U19975 ( .A(n15713), .B(n15714), .Z(y[850]) );
  NAND U19976 ( .A(n15381), .B(m[850]), .Z(n15714) );
  NAND U19977 ( .A(n15382), .B(creg[850]), .Z(n15713) );
  NAND U19978 ( .A(n15715), .B(n15716), .Z(y[84]) );
  NAND U19979 ( .A(n15381), .B(m[84]), .Z(n15716) );
  NAND U19980 ( .A(n15382), .B(creg[84]), .Z(n15715) );
  NAND U19981 ( .A(n15717), .B(n15718), .Z(y[849]) );
  NAND U19982 ( .A(n15381), .B(m[849]), .Z(n15718) );
  NAND U19983 ( .A(n15382), .B(creg[849]), .Z(n15717) );
  NAND U19984 ( .A(n15719), .B(n15720), .Z(y[848]) );
  NAND U19985 ( .A(n15381), .B(m[848]), .Z(n15720) );
  NAND U19986 ( .A(n15382), .B(creg[848]), .Z(n15719) );
  NAND U19987 ( .A(n15721), .B(n15722), .Z(y[847]) );
  NAND U19988 ( .A(n15381), .B(m[847]), .Z(n15722) );
  NAND U19989 ( .A(n15382), .B(creg[847]), .Z(n15721) );
  NAND U19990 ( .A(n15723), .B(n15724), .Z(y[846]) );
  NAND U19991 ( .A(n15381), .B(m[846]), .Z(n15724) );
  NAND U19992 ( .A(n15382), .B(creg[846]), .Z(n15723) );
  NAND U19993 ( .A(n15725), .B(n15726), .Z(y[845]) );
  NAND U19994 ( .A(n15381), .B(m[845]), .Z(n15726) );
  NAND U19995 ( .A(n15382), .B(creg[845]), .Z(n15725) );
  NAND U19996 ( .A(n15727), .B(n15728), .Z(y[844]) );
  NAND U19997 ( .A(n15381), .B(m[844]), .Z(n15728) );
  NAND U19998 ( .A(n15382), .B(creg[844]), .Z(n15727) );
  NAND U19999 ( .A(n15729), .B(n15730), .Z(y[843]) );
  NAND U20000 ( .A(n15381), .B(m[843]), .Z(n15730) );
  NAND U20001 ( .A(n15382), .B(creg[843]), .Z(n15729) );
  NAND U20002 ( .A(n15731), .B(n15732), .Z(y[842]) );
  NAND U20003 ( .A(n15381), .B(m[842]), .Z(n15732) );
  NAND U20004 ( .A(n15382), .B(creg[842]), .Z(n15731) );
  NAND U20005 ( .A(n15733), .B(n15734), .Z(y[841]) );
  NAND U20006 ( .A(n15381), .B(m[841]), .Z(n15734) );
  NAND U20007 ( .A(n15382), .B(creg[841]), .Z(n15733) );
  NAND U20008 ( .A(n15735), .B(n15736), .Z(y[840]) );
  NAND U20009 ( .A(n15381), .B(m[840]), .Z(n15736) );
  NAND U20010 ( .A(n15382), .B(creg[840]), .Z(n15735) );
  NAND U20011 ( .A(n15737), .B(n15738), .Z(y[83]) );
  NAND U20012 ( .A(n15381), .B(m[83]), .Z(n15738) );
  NAND U20013 ( .A(n15382), .B(creg[83]), .Z(n15737) );
  NAND U20014 ( .A(n15739), .B(n15740), .Z(y[839]) );
  NAND U20015 ( .A(n15381), .B(m[839]), .Z(n15740) );
  NAND U20016 ( .A(n15382), .B(creg[839]), .Z(n15739) );
  NAND U20017 ( .A(n15741), .B(n15742), .Z(y[838]) );
  NAND U20018 ( .A(n15381), .B(m[838]), .Z(n15742) );
  NAND U20019 ( .A(n15382), .B(creg[838]), .Z(n15741) );
  NAND U20020 ( .A(n15743), .B(n15744), .Z(y[837]) );
  NAND U20021 ( .A(n15381), .B(m[837]), .Z(n15744) );
  NAND U20022 ( .A(n15382), .B(creg[837]), .Z(n15743) );
  NAND U20023 ( .A(n15745), .B(n15746), .Z(y[836]) );
  NAND U20024 ( .A(n15381), .B(m[836]), .Z(n15746) );
  NAND U20025 ( .A(n15382), .B(creg[836]), .Z(n15745) );
  NAND U20026 ( .A(n15747), .B(n15748), .Z(y[835]) );
  NAND U20027 ( .A(n15381), .B(m[835]), .Z(n15748) );
  NAND U20028 ( .A(n15382), .B(creg[835]), .Z(n15747) );
  NAND U20029 ( .A(n15749), .B(n15750), .Z(y[834]) );
  NAND U20030 ( .A(n15381), .B(m[834]), .Z(n15750) );
  NAND U20031 ( .A(n15382), .B(creg[834]), .Z(n15749) );
  NAND U20032 ( .A(n15751), .B(n15752), .Z(y[833]) );
  NAND U20033 ( .A(n15381), .B(m[833]), .Z(n15752) );
  NAND U20034 ( .A(n15382), .B(creg[833]), .Z(n15751) );
  NAND U20035 ( .A(n15753), .B(n15754), .Z(y[832]) );
  NAND U20036 ( .A(n15381), .B(m[832]), .Z(n15754) );
  NAND U20037 ( .A(n15382), .B(creg[832]), .Z(n15753) );
  NAND U20038 ( .A(n15755), .B(n15756), .Z(y[831]) );
  NAND U20039 ( .A(n15381), .B(m[831]), .Z(n15756) );
  NAND U20040 ( .A(n15382), .B(creg[831]), .Z(n15755) );
  NAND U20041 ( .A(n15757), .B(n15758), .Z(y[830]) );
  NAND U20042 ( .A(n15381), .B(m[830]), .Z(n15758) );
  NAND U20043 ( .A(n15382), .B(creg[830]), .Z(n15757) );
  NAND U20044 ( .A(n15759), .B(n15760), .Z(y[82]) );
  NAND U20045 ( .A(n15381), .B(m[82]), .Z(n15760) );
  NAND U20046 ( .A(n15382), .B(creg[82]), .Z(n15759) );
  NAND U20047 ( .A(n15761), .B(n15762), .Z(y[829]) );
  NAND U20048 ( .A(n15381), .B(m[829]), .Z(n15762) );
  NAND U20049 ( .A(n15382), .B(creg[829]), .Z(n15761) );
  NAND U20050 ( .A(n15763), .B(n15764), .Z(y[828]) );
  NAND U20051 ( .A(n15381), .B(m[828]), .Z(n15764) );
  NAND U20052 ( .A(n15382), .B(creg[828]), .Z(n15763) );
  NAND U20053 ( .A(n15765), .B(n15766), .Z(y[827]) );
  NAND U20054 ( .A(n15381), .B(m[827]), .Z(n15766) );
  NAND U20055 ( .A(n15382), .B(creg[827]), .Z(n15765) );
  NAND U20056 ( .A(n15767), .B(n15768), .Z(y[826]) );
  NAND U20057 ( .A(n15381), .B(m[826]), .Z(n15768) );
  NAND U20058 ( .A(n15382), .B(creg[826]), .Z(n15767) );
  NAND U20059 ( .A(n15769), .B(n15770), .Z(y[825]) );
  NAND U20060 ( .A(n15381), .B(m[825]), .Z(n15770) );
  NAND U20061 ( .A(n15382), .B(creg[825]), .Z(n15769) );
  NAND U20062 ( .A(n15771), .B(n15772), .Z(y[824]) );
  NAND U20063 ( .A(n15381), .B(m[824]), .Z(n15772) );
  NAND U20064 ( .A(n15382), .B(creg[824]), .Z(n15771) );
  NAND U20065 ( .A(n15773), .B(n15774), .Z(y[823]) );
  NAND U20066 ( .A(n15381), .B(m[823]), .Z(n15774) );
  NAND U20067 ( .A(n15382), .B(creg[823]), .Z(n15773) );
  NAND U20068 ( .A(n15775), .B(n15776), .Z(y[822]) );
  NAND U20069 ( .A(n15381), .B(m[822]), .Z(n15776) );
  NAND U20070 ( .A(n15382), .B(creg[822]), .Z(n15775) );
  NAND U20071 ( .A(n15777), .B(n15778), .Z(y[821]) );
  NAND U20072 ( .A(n15381), .B(m[821]), .Z(n15778) );
  NAND U20073 ( .A(n15382), .B(creg[821]), .Z(n15777) );
  NAND U20074 ( .A(n15779), .B(n15780), .Z(y[820]) );
  NAND U20075 ( .A(n15381), .B(m[820]), .Z(n15780) );
  NAND U20076 ( .A(n15382), .B(creg[820]), .Z(n15779) );
  NAND U20077 ( .A(n15781), .B(n15782), .Z(y[81]) );
  NAND U20078 ( .A(n15381), .B(m[81]), .Z(n15782) );
  NAND U20079 ( .A(n15382), .B(creg[81]), .Z(n15781) );
  NAND U20080 ( .A(n15783), .B(n15784), .Z(y[819]) );
  NAND U20081 ( .A(n15381), .B(m[819]), .Z(n15784) );
  NAND U20082 ( .A(n15382), .B(creg[819]), .Z(n15783) );
  NAND U20083 ( .A(n15785), .B(n15786), .Z(y[818]) );
  NAND U20084 ( .A(n15381), .B(m[818]), .Z(n15786) );
  NAND U20085 ( .A(n15382), .B(creg[818]), .Z(n15785) );
  NAND U20086 ( .A(n15787), .B(n15788), .Z(y[817]) );
  NAND U20087 ( .A(n15381), .B(m[817]), .Z(n15788) );
  NAND U20088 ( .A(n15382), .B(creg[817]), .Z(n15787) );
  NAND U20089 ( .A(n15789), .B(n15790), .Z(y[816]) );
  NAND U20090 ( .A(n15381), .B(m[816]), .Z(n15790) );
  NAND U20091 ( .A(n15382), .B(creg[816]), .Z(n15789) );
  NAND U20092 ( .A(n15791), .B(n15792), .Z(y[815]) );
  NAND U20093 ( .A(n15381), .B(m[815]), .Z(n15792) );
  NAND U20094 ( .A(n15382), .B(creg[815]), .Z(n15791) );
  NAND U20095 ( .A(n15793), .B(n15794), .Z(y[814]) );
  NAND U20096 ( .A(n15381), .B(m[814]), .Z(n15794) );
  NAND U20097 ( .A(n15382), .B(creg[814]), .Z(n15793) );
  NAND U20098 ( .A(n15795), .B(n15796), .Z(y[813]) );
  NAND U20099 ( .A(n15381), .B(m[813]), .Z(n15796) );
  NAND U20100 ( .A(n15382), .B(creg[813]), .Z(n15795) );
  NAND U20101 ( .A(n15797), .B(n15798), .Z(y[812]) );
  NAND U20102 ( .A(n15381), .B(m[812]), .Z(n15798) );
  NAND U20103 ( .A(n15382), .B(creg[812]), .Z(n15797) );
  NAND U20104 ( .A(n15799), .B(n15800), .Z(y[811]) );
  NAND U20105 ( .A(n15381), .B(m[811]), .Z(n15800) );
  NAND U20106 ( .A(n15382), .B(creg[811]), .Z(n15799) );
  NAND U20107 ( .A(n15801), .B(n15802), .Z(y[810]) );
  NAND U20108 ( .A(n15381), .B(m[810]), .Z(n15802) );
  NAND U20109 ( .A(n15382), .B(creg[810]), .Z(n15801) );
  NAND U20110 ( .A(n15803), .B(n15804), .Z(y[80]) );
  NAND U20111 ( .A(n15381), .B(m[80]), .Z(n15804) );
  NAND U20112 ( .A(n15382), .B(creg[80]), .Z(n15803) );
  NAND U20113 ( .A(n15805), .B(n15806), .Z(y[809]) );
  NAND U20114 ( .A(n15381), .B(m[809]), .Z(n15806) );
  NAND U20115 ( .A(n15382), .B(creg[809]), .Z(n15805) );
  NAND U20116 ( .A(n15807), .B(n15808), .Z(y[808]) );
  NAND U20117 ( .A(n15381), .B(m[808]), .Z(n15808) );
  NAND U20118 ( .A(n15382), .B(creg[808]), .Z(n15807) );
  NAND U20119 ( .A(n15809), .B(n15810), .Z(y[807]) );
  NAND U20120 ( .A(n15381), .B(m[807]), .Z(n15810) );
  NAND U20121 ( .A(n15382), .B(creg[807]), .Z(n15809) );
  NAND U20122 ( .A(n15811), .B(n15812), .Z(y[806]) );
  NAND U20123 ( .A(n15381), .B(m[806]), .Z(n15812) );
  NAND U20124 ( .A(n15382), .B(creg[806]), .Z(n15811) );
  NAND U20125 ( .A(n15813), .B(n15814), .Z(y[805]) );
  NAND U20126 ( .A(n15381), .B(m[805]), .Z(n15814) );
  NAND U20127 ( .A(n15382), .B(creg[805]), .Z(n15813) );
  NAND U20128 ( .A(n15815), .B(n15816), .Z(y[804]) );
  NAND U20129 ( .A(n15381), .B(m[804]), .Z(n15816) );
  NAND U20130 ( .A(n15382), .B(creg[804]), .Z(n15815) );
  NAND U20131 ( .A(n15817), .B(n15818), .Z(y[803]) );
  NAND U20132 ( .A(n15381), .B(m[803]), .Z(n15818) );
  NAND U20133 ( .A(n15382), .B(creg[803]), .Z(n15817) );
  NAND U20134 ( .A(n15819), .B(n15820), .Z(y[802]) );
  NAND U20135 ( .A(n15381), .B(m[802]), .Z(n15820) );
  NAND U20136 ( .A(n15382), .B(creg[802]), .Z(n15819) );
  NAND U20137 ( .A(n15821), .B(n15822), .Z(y[801]) );
  NAND U20138 ( .A(n15381), .B(m[801]), .Z(n15822) );
  NAND U20139 ( .A(n15382), .B(creg[801]), .Z(n15821) );
  NAND U20140 ( .A(n15823), .B(n15824), .Z(y[800]) );
  NAND U20141 ( .A(n15381), .B(m[800]), .Z(n15824) );
  NAND U20142 ( .A(n15382), .B(creg[800]), .Z(n15823) );
  NAND U20143 ( .A(n15825), .B(n15826), .Z(y[7]) );
  NAND U20144 ( .A(n15381), .B(m[7]), .Z(n15826) );
  NAND U20145 ( .A(n15382), .B(creg[7]), .Z(n15825) );
  NAND U20146 ( .A(n15827), .B(n15828), .Z(y[79]) );
  NAND U20147 ( .A(n15381), .B(m[79]), .Z(n15828) );
  NAND U20148 ( .A(n15382), .B(creg[79]), .Z(n15827) );
  NAND U20149 ( .A(n15829), .B(n15830), .Z(y[799]) );
  NAND U20150 ( .A(n15381), .B(m[799]), .Z(n15830) );
  NAND U20151 ( .A(n15382), .B(creg[799]), .Z(n15829) );
  NAND U20152 ( .A(n15831), .B(n15832), .Z(y[798]) );
  NAND U20153 ( .A(n15381), .B(m[798]), .Z(n15832) );
  NAND U20154 ( .A(n15382), .B(creg[798]), .Z(n15831) );
  NAND U20155 ( .A(n15833), .B(n15834), .Z(y[797]) );
  NAND U20156 ( .A(n15381), .B(m[797]), .Z(n15834) );
  NAND U20157 ( .A(n15382), .B(creg[797]), .Z(n15833) );
  NAND U20158 ( .A(n15835), .B(n15836), .Z(y[796]) );
  NAND U20159 ( .A(n15381), .B(m[796]), .Z(n15836) );
  NAND U20160 ( .A(n15382), .B(creg[796]), .Z(n15835) );
  NAND U20161 ( .A(n15837), .B(n15838), .Z(y[795]) );
  NAND U20162 ( .A(n15381), .B(m[795]), .Z(n15838) );
  NAND U20163 ( .A(n15382), .B(creg[795]), .Z(n15837) );
  NAND U20164 ( .A(n15839), .B(n15840), .Z(y[794]) );
  NAND U20165 ( .A(n15381), .B(m[794]), .Z(n15840) );
  NAND U20166 ( .A(n15382), .B(creg[794]), .Z(n15839) );
  NAND U20167 ( .A(n15841), .B(n15842), .Z(y[793]) );
  NAND U20168 ( .A(n15381), .B(m[793]), .Z(n15842) );
  NAND U20169 ( .A(n15382), .B(creg[793]), .Z(n15841) );
  NAND U20170 ( .A(n15843), .B(n15844), .Z(y[792]) );
  NAND U20171 ( .A(n15381), .B(m[792]), .Z(n15844) );
  NAND U20172 ( .A(n15382), .B(creg[792]), .Z(n15843) );
  NAND U20173 ( .A(n15845), .B(n15846), .Z(y[791]) );
  NAND U20174 ( .A(n15381), .B(m[791]), .Z(n15846) );
  NAND U20175 ( .A(n15382), .B(creg[791]), .Z(n15845) );
  NAND U20176 ( .A(n15847), .B(n15848), .Z(y[790]) );
  NAND U20177 ( .A(n15381), .B(m[790]), .Z(n15848) );
  NAND U20178 ( .A(n15382), .B(creg[790]), .Z(n15847) );
  NAND U20179 ( .A(n15849), .B(n15850), .Z(y[78]) );
  NAND U20180 ( .A(n15381), .B(m[78]), .Z(n15850) );
  NAND U20181 ( .A(n15382), .B(creg[78]), .Z(n15849) );
  NAND U20182 ( .A(n15851), .B(n15852), .Z(y[789]) );
  NAND U20183 ( .A(n15381), .B(m[789]), .Z(n15852) );
  NAND U20184 ( .A(n15382), .B(creg[789]), .Z(n15851) );
  NAND U20185 ( .A(n15853), .B(n15854), .Z(y[788]) );
  NAND U20186 ( .A(n15381), .B(m[788]), .Z(n15854) );
  NAND U20187 ( .A(n15382), .B(creg[788]), .Z(n15853) );
  NAND U20188 ( .A(n15855), .B(n15856), .Z(y[787]) );
  NAND U20189 ( .A(n15381), .B(m[787]), .Z(n15856) );
  NAND U20190 ( .A(n15382), .B(creg[787]), .Z(n15855) );
  NAND U20191 ( .A(n15857), .B(n15858), .Z(y[786]) );
  NAND U20192 ( .A(n15381), .B(m[786]), .Z(n15858) );
  NAND U20193 ( .A(n15382), .B(creg[786]), .Z(n15857) );
  NAND U20194 ( .A(n15859), .B(n15860), .Z(y[785]) );
  NAND U20195 ( .A(n15381), .B(m[785]), .Z(n15860) );
  NAND U20196 ( .A(n15382), .B(creg[785]), .Z(n15859) );
  NAND U20197 ( .A(n15861), .B(n15862), .Z(y[784]) );
  NAND U20198 ( .A(n15381), .B(m[784]), .Z(n15862) );
  NAND U20199 ( .A(n15382), .B(creg[784]), .Z(n15861) );
  NAND U20200 ( .A(n15863), .B(n15864), .Z(y[783]) );
  NAND U20201 ( .A(n15381), .B(m[783]), .Z(n15864) );
  NAND U20202 ( .A(n15382), .B(creg[783]), .Z(n15863) );
  NAND U20203 ( .A(n15865), .B(n15866), .Z(y[782]) );
  NAND U20204 ( .A(n15381), .B(m[782]), .Z(n15866) );
  NAND U20205 ( .A(n15382), .B(creg[782]), .Z(n15865) );
  NAND U20206 ( .A(n15867), .B(n15868), .Z(y[781]) );
  NAND U20207 ( .A(n15381), .B(m[781]), .Z(n15868) );
  NAND U20208 ( .A(n15382), .B(creg[781]), .Z(n15867) );
  NAND U20209 ( .A(n15869), .B(n15870), .Z(y[780]) );
  NAND U20210 ( .A(n15381), .B(m[780]), .Z(n15870) );
  NAND U20211 ( .A(n15382), .B(creg[780]), .Z(n15869) );
  NAND U20212 ( .A(n15871), .B(n15872), .Z(y[77]) );
  NAND U20213 ( .A(n15381), .B(m[77]), .Z(n15872) );
  NAND U20214 ( .A(n15382), .B(creg[77]), .Z(n15871) );
  NAND U20215 ( .A(n15873), .B(n15874), .Z(y[779]) );
  NAND U20216 ( .A(n15381), .B(m[779]), .Z(n15874) );
  NAND U20217 ( .A(n15382), .B(creg[779]), .Z(n15873) );
  NAND U20218 ( .A(n15875), .B(n15876), .Z(y[778]) );
  NAND U20219 ( .A(n15381), .B(m[778]), .Z(n15876) );
  NAND U20220 ( .A(n15382), .B(creg[778]), .Z(n15875) );
  NAND U20221 ( .A(n15877), .B(n15878), .Z(y[777]) );
  NAND U20222 ( .A(n15381), .B(m[777]), .Z(n15878) );
  NAND U20223 ( .A(n15382), .B(creg[777]), .Z(n15877) );
  NAND U20224 ( .A(n15879), .B(n15880), .Z(y[776]) );
  NAND U20225 ( .A(n15381), .B(m[776]), .Z(n15880) );
  NAND U20226 ( .A(n15382), .B(creg[776]), .Z(n15879) );
  NAND U20227 ( .A(n15881), .B(n15882), .Z(y[775]) );
  NAND U20228 ( .A(n15381), .B(m[775]), .Z(n15882) );
  NAND U20229 ( .A(n15382), .B(creg[775]), .Z(n15881) );
  NAND U20230 ( .A(n15883), .B(n15884), .Z(y[774]) );
  NAND U20231 ( .A(n15381), .B(m[774]), .Z(n15884) );
  NAND U20232 ( .A(n15382), .B(creg[774]), .Z(n15883) );
  NAND U20233 ( .A(n15885), .B(n15886), .Z(y[773]) );
  NAND U20234 ( .A(n15381), .B(m[773]), .Z(n15886) );
  NAND U20235 ( .A(n15382), .B(creg[773]), .Z(n15885) );
  NAND U20236 ( .A(n15887), .B(n15888), .Z(y[772]) );
  NAND U20237 ( .A(n15381), .B(m[772]), .Z(n15888) );
  NAND U20238 ( .A(n15382), .B(creg[772]), .Z(n15887) );
  NAND U20239 ( .A(n15889), .B(n15890), .Z(y[771]) );
  NAND U20240 ( .A(n15381), .B(m[771]), .Z(n15890) );
  NAND U20241 ( .A(n15382), .B(creg[771]), .Z(n15889) );
  NAND U20242 ( .A(n15891), .B(n15892), .Z(y[770]) );
  NAND U20243 ( .A(n15381), .B(m[770]), .Z(n15892) );
  NAND U20244 ( .A(n15382), .B(creg[770]), .Z(n15891) );
  NAND U20245 ( .A(n15893), .B(n15894), .Z(y[76]) );
  NAND U20246 ( .A(n15381), .B(m[76]), .Z(n15894) );
  NAND U20247 ( .A(n15382), .B(creg[76]), .Z(n15893) );
  NAND U20248 ( .A(n15895), .B(n15896), .Z(y[769]) );
  NAND U20249 ( .A(n15381), .B(m[769]), .Z(n15896) );
  NAND U20250 ( .A(n15382), .B(creg[769]), .Z(n15895) );
  NAND U20251 ( .A(n15897), .B(n15898), .Z(y[768]) );
  NAND U20252 ( .A(n15381), .B(m[768]), .Z(n15898) );
  NAND U20253 ( .A(n15382), .B(creg[768]), .Z(n15897) );
  NAND U20254 ( .A(n15899), .B(n15900), .Z(y[767]) );
  NAND U20255 ( .A(n15381), .B(m[767]), .Z(n15900) );
  NAND U20256 ( .A(n15382), .B(creg[767]), .Z(n15899) );
  NAND U20257 ( .A(n15901), .B(n15902), .Z(y[766]) );
  NAND U20258 ( .A(n15381), .B(m[766]), .Z(n15902) );
  NAND U20259 ( .A(n15382), .B(creg[766]), .Z(n15901) );
  NAND U20260 ( .A(n15903), .B(n15904), .Z(y[765]) );
  NAND U20261 ( .A(n15381), .B(m[765]), .Z(n15904) );
  NAND U20262 ( .A(n15382), .B(creg[765]), .Z(n15903) );
  NAND U20263 ( .A(n15905), .B(n15906), .Z(y[764]) );
  NAND U20264 ( .A(n15381), .B(m[764]), .Z(n15906) );
  NAND U20265 ( .A(n15382), .B(creg[764]), .Z(n15905) );
  NAND U20266 ( .A(n15907), .B(n15908), .Z(y[763]) );
  NAND U20267 ( .A(n15381), .B(m[763]), .Z(n15908) );
  NAND U20268 ( .A(n15382), .B(creg[763]), .Z(n15907) );
  NAND U20269 ( .A(n15909), .B(n15910), .Z(y[762]) );
  NAND U20270 ( .A(n15381), .B(m[762]), .Z(n15910) );
  NAND U20271 ( .A(n15382), .B(creg[762]), .Z(n15909) );
  NAND U20272 ( .A(n15911), .B(n15912), .Z(y[761]) );
  NAND U20273 ( .A(n15381), .B(m[761]), .Z(n15912) );
  NAND U20274 ( .A(n15382), .B(creg[761]), .Z(n15911) );
  NAND U20275 ( .A(n15913), .B(n15914), .Z(y[760]) );
  NAND U20276 ( .A(n15381), .B(m[760]), .Z(n15914) );
  NAND U20277 ( .A(n15382), .B(creg[760]), .Z(n15913) );
  NAND U20278 ( .A(n15915), .B(n15916), .Z(y[75]) );
  NAND U20279 ( .A(n15381), .B(m[75]), .Z(n15916) );
  NAND U20280 ( .A(n15382), .B(creg[75]), .Z(n15915) );
  NAND U20281 ( .A(n15917), .B(n15918), .Z(y[759]) );
  NAND U20282 ( .A(n15381), .B(m[759]), .Z(n15918) );
  NAND U20283 ( .A(n15382), .B(creg[759]), .Z(n15917) );
  NAND U20284 ( .A(n15919), .B(n15920), .Z(y[758]) );
  NAND U20285 ( .A(n15381), .B(m[758]), .Z(n15920) );
  NAND U20286 ( .A(n15382), .B(creg[758]), .Z(n15919) );
  NAND U20287 ( .A(n15921), .B(n15922), .Z(y[757]) );
  NAND U20288 ( .A(n15381), .B(m[757]), .Z(n15922) );
  NAND U20289 ( .A(n15382), .B(creg[757]), .Z(n15921) );
  NAND U20290 ( .A(n15923), .B(n15924), .Z(y[756]) );
  NAND U20291 ( .A(n15381), .B(m[756]), .Z(n15924) );
  NAND U20292 ( .A(n15382), .B(creg[756]), .Z(n15923) );
  NAND U20293 ( .A(n15925), .B(n15926), .Z(y[755]) );
  NAND U20294 ( .A(n15381), .B(m[755]), .Z(n15926) );
  NAND U20295 ( .A(n15382), .B(creg[755]), .Z(n15925) );
  NAND U20296 ( .A(n15927), .B(n15928), .Z(y[754]) );
  NAND U20297 ( .A(n15381), .B(m[754]), .Z(n15928) );
  NAND U20298 ( .A(n15382), .B(creg[754]), .Z(n15927) );
  NAND U20299 ( .A(n15929), .B(n15930), .Z(y[753]) );
  NAND U20300 ( .A(n15381), .B(m[753]), .Z(n15930) );
  NAND U20301 ( .A(n15382), .B(creg[753]), .Z(n15929) );
  NAND U20302 ( .A(n15931), .B(n15932), .Z(y[752]) );
  NAND U20303 ( .A(n15381), .B(m[752]), .Z(n15932) );
  NAND U20304 ( .A(n15382), .B(creg[752]), .Z(n15931) );
  NAND U20305 ( .A(n15933), .B(n15934), .Z(y[751]) );
  NAND U20306 ( .A(n15381), .B(m[751]), .Z(n15934) );
  NAND U20307 ( .A(n15382), .B(creg[751]), .Z(n15933) );
  NAND U20308 ( .A(n15935), .B(n15936), .Z(y[750]) );
  NAND U20309 ( .A(n15381), .B(m[750]), .Z(n15936) );
  NAND U20310 ( .A(n15382), .B(creg[750]), .Z(n15935) );
  NAND U20311 ( .A(n15937), .B(n15938), .Z(y[74]) );
  NAND U20312 ( .A(n15381), .B(m[74]), .Z(n15938) );
  NAND U20313 ( .A(n15382), .B(creg[74]), .Z(n15937) );
  NAND U20314 ( .A(n15939), .B(n15940), .Z(y[749]) );
  NAND U20315 ( .A(n15381), .B(m[749]), .Z(n15940) );
  NAND U20316 ( .A(n15382), .B(creg[749]), .Z(n15939) );
  NAND U20317 ( .A(n15941), .B(n15942), .Z(y[748]) );
  NAND U20318 ( .A(n15381), .B(m[748]), .Z(n15942) );
  NAND U20319 ( .A(n15382), .B(creg[748]), .Z(n15941) );
  NAND U20320 ( .A(n15943), .B(n15944), .Z(y[747]) );
  NAND U20321 ( .A(n15381), .B(m[747]), .Z(n15944) );
  NAND U20322 ( .A(n15382), .B(creg[747]), .Z(n15943) );
  NAND U20323 ( .A(n15945), .B(n15946), .Z(y[746]) );
  NAND U20324 ( .A(n15381), .B(m[746]), .Z(n15946) );
  NAND U20325 ( .A(n15382), .B(creg[746]), .Z(n15945) );
  NAND U20326 ( .A(n15947), .B(n15948), .Z(y[745]) );
  NAND U20327 ( .A(n15381), .B(m[745]), .Z(n15948) );
  NAND U20328 ( .A(n15382), .B(creg[745]), .Z(n15947) );
  NAND U20329 ( .A(n15949), .B(n15950), .Z(y[744]) );
  NAND U20330 ( .A(n15381), .B(m[744]), .Z(n15950) );
  NAND U20331 ( .A(n15382), .B(creg[744]), .Z(n15949) );
  NAND U20332 ( .A(n15951), .B(n15952), .Z(y[743]) );
  NAND U20333 ( .A(n15381), .B(m[743]), .Z(n15952) );
  NAND U20334 ( .A(n15382), .B(creg[743]), .Z(n15951) );
  NAND U20335 ( .A(n15953), .B(n15954), .Z(y[742]) );
  NAND U20336 ( .A(n15381), .B(m[742]), .Z(n15954) );
  NAND U20337 ( .A(n15382), .B(creg[742]), .Z(n15953) );
  NAND U20338 ( .A(n15955), .B(n15956), .Z(y[741]) );
  NAND U20339 ( .A(n15381), .B(m[741]), .Z(n15956) );
  NAND U20340 ( .A(n15382), .B(creg[741]), .Z(n15955) );
  NAND U20341 ( .A(n15957), .B(n15958), .Z(y[740]) );
  NAND U20342 ( .A(n15381), .B(m[740]), .Z(n15958) );
  NAND U20343 ( .A(n15382), .B(creg[740]), .Z(n15957) );
  NAND U20344 ( .A(n15959), .B(n15960), .Z(y[73]) );
  NAND U20345 ( .A(n15381), .B(m[73]), .Z(n15960) );
  NAND U20346 ( .A(n15382), .B(creg[73]), .Z(n15959) );
  NAND U20347 ( .A(n15961), .B(n15962), .Z(y[739]) );
  NAND U20348 ( .A(n15381), .B(m[739]), .Z(n15962) );
  NAND U20349 ( .A(n15382), .B(creg[739]), .Z(n15961) );
  NAND U20350 ( .A(n15963), .B(n15964), .Z(y[738]) );
  NAND U20351 ( .A(n15381), .B(m[738]), .Z(n15964) );
  NAND U20352 ( .A(n15382), .B(creg[738]), .Z(n15963) );
  NAND U20353 ( .A(n15965), .B(n15966), .Z(y[737]) );
  NAND U20354 ( .A(n15381), .B(m[737]), .Z(n15966) );
  NAND U20355 ( .A(n15382), .B(creg[737]), .Z(n15965) );
  NAND U20356 ( .A(n15967), .B(n15968), .Z(y[736]) );
  NAND U20357 ( .A(n15381), .B(m[736]), .Z(n15968) );
  NAND U20358 ( .A(n15382), .B(creg[736]), .Z(n15967) );
  NAND U20359 ( .A(n15969), .B(n15970), .Z(y[735]) );
  NAND U20360 ( .A(n15381), .B(m[735]), .Z(n15970) );
  NAND U20361 ( .A(n15382), .B(creg[735]), .Z(n15969) );
  NAND U20362 ( .A(n15971), .B(n15972), .Z(y[734]) );
  NAND U20363 ( .A(n15381), .B(m[734]), .Z(n15972) );
  NAND U20364 ( .A(n15382), .B(creg[734]), .Z(n15971) );
  NAND U20365 ( .A(n15973), .B(n15974), .Z(y[733]) );
  NAND U20366 ( .A(n15381), .B(m[733]), .Z(n15974) );
  NAND U20367 ( .A(n15382), .B(creg[733]), .Z(n15973) );
  NAND U20368 ( .A(n15975), .B(n15976), .Z(y[732]) );
  NAND U20369 ( .A(n15381), .B(m[732]), .Z(n15976) );
  NAND U20370 ( .A(n15382), .B(creg[732]), .Z(n15975) );
  NAND U20371 ( .A(n15977), .B(n15978), .Z(y[731]) );
  NAND U20372 ( .A(n15381), .B(m[731]), .Z(n15978) );
  NAND U20373 ( .A(n15382), .B(creg[731]), .Z(n15977) );
  NAND U20374 ( .A(n15979), .B(n15980), .Z(y[730]) );
  NAND U20375 ( .A(n15381), .B(m[730]), .Z(n15980) );
  NAND U20376 ( .A(n15382), .B(creg[730]), .Z(n15979) );
  NAND U20377 ( .A(n15981), .B(n15982), .Z(y[72]) );
  NAND U20378 ( .A(n15381), .B(m[72]), .Z(n15982) );
  NAND U20379 ( .A(n15382), .B(creg[72]), .Z(n15981) );
  NAND U20380 ( .A(n15983), .B(n15984), .Z(y[729]) );
  NAND U20381 ( .A(n15381), .B(m[729]), .Z(n15984) );
  NAND U20382 ( .A(n15382), .B(creg[729]), .Z(n15983) );
  NAND U20383 ( .A(n15985), .B(n15986), .Z(y[728]) );
  NAND U20384 ( .A(n15381), .B(m[728]), .Z(n15986) );
  NAND U20385 ( .A(n15382), .B(creg[728]), .Z(n15985) );
  NAND U20386 ( .A(n15987), .B(n15988), .Z(y[727]) );
  NAND U20387 ( .A(n15381), .B(m[727]), .Z(n15988) );
  NAND U20388 ( .A(n15382), .B(creg[727]), .Z(n15987) );
  NAND U20389 ( .A(n15989), .B(n15990), .Z(y[726]) );
  NAND U20390 ( .A(n15381), .B(m[726]), .Z(n15990) );
  NAND U20391 ( .A(n15382), .B(creg[726]), .Z(n15989) );
  NAND U20392 ( .A(n15991), .B(n15992), .Z(y[725]) );
  NAND U20393 ( .A(n15381), .B(m[725]), .Z(n15992) );
  NAND U20394 ( .A(n15382), .B(creg[725]), .Z(n15991) );
  NAND U20395 ( .A(n15993), .B(n15994), .Z(y[724]) );
  NAND U20396 ( .A(n15381), .B(m[724]), .Z(n15994) );
  NAND U20397 ( .A(n15382), .B(creg[724]), .Z(n15993) );
  NAND U20398 ( .A(n15995), .B(n15996), .Z(y[723]) );
  NAND U20399 ( .A(n15381), .B(m[723]), .Z(n15996) );
  NAND U20400 ( .A(n15382), .B(creg[723]), .Z(n15995) );
  NAND U20401 ( .A(n15997), .B(n15998), .Z(y[722]) );
  NAND U20402 ( .A(n15381), .B(m[722]), .Z(n15998) );
  NAND U20403 ( .A(n15382), .B(creg[722]), .Z(n15997) );
  NAND U20404 ( .A(n15999), .B(n16000), .Z(y[721]) );
  NAND U20405 ( .A(n15381), .B(m[721]), .Z(n16000) );
  NAND U20406 ( .A(n15382), .B(creg[721]), .Z(n15999) );
  NAND U20407 ( .A(n16001), .B(n16002), .Z(y[720]) );
  NAND U20408 ( .A(n15381), .B(m[720]), .Z(n16002) );
  NAND U20409 ( .A(n15382), .B(creg[720]), .Z(n16001) );
  NAND U20410 ( .A(n16003), .B(n16004), .Z(y[71]) );
  NAND U20411 ( .A(n15381), .B(m[71]), .Z(n16004) );
  NAND U20412 ( .A(n15382), .B(creg[71]), .Z(n16003) );
  NAND U20413 ( .A(n16005), .B(n16006), .Z(y[719]) );
  NAND U20414 ( .A(n15381), .B(m[719]), .Z(n16006) );
  NAND U20415 ( .A(n15382), .B(creg[719]), .Z(n16005) );
  NAND U20416 ( .A(n16007), .B(n16008), .Z(y[718]) );
  NAND U20417 ( .A(n15381), .B(m[718]), .Z(n16008) );
  NAND U20418 ( .A(n15382), .B(creg[718]), .Z(n16007) );
  NAND U20419 ( .A(n16009), .B(n16010), .Z(y[717]) );
  NAND U20420 ( .A(n15381), .B(m[717]), .Z(n16010) );
  NAND U20421 ( .A(n15382), .B(creg[717]), .Z(n16009) );
  NAND U20422 ( .A(n16011), .B(n16012), .Z(y[716]) );
  NAND U20423 ( .A(n15381), .B(m[716]), .Z(n16012) );
  NAND U20424 ( .A(n15382), .B(creg[716]), .Z(n16011) );
  NAND U20425 ( .A(n16013), .B(n16014), .Z(y[715]) );
  NAND U20426 ( .A(n15381), .B(m[715]), .Z(n16014) );
  NAND U20427 ( .A(n15382), .B(creg[715]), .Z(n16013) );
  NAND U20428 ( .A(n16015), .B(n16016), .Z(y[714]) );
  NAND U20429 ( .A(n15381), .B(m[714]), .Z(n16016) );
  NAND U20430 ( .A(n15382), .B(creg[714]), .Z(n16015) );
  NAND U20431 ( .A(n16017), .B(n16018), .Z(y[713]) );
  NAND U20432 ( .A(n15381), .B(m[713]), .Z(n16018) );
  NAND U20433 ( .A(n15382), .B(creg[713]), .Z(n16017) );
  NAND U20434 ( .A(n16019), .B(n16020), .Z(y[712]) );
  NAND U20435 ( .A(n15381), .B(m[712]), .Z(n16020) );
  NAND U20436 ( .A(n15382), .B(creg[712]), .Z(n16019) );
  NAND U20437 ( .A(n16021), .B(n16022), .Z(y[711]) );
  NAND U20438 ( .A(n15381), .B(m[711]), .Z(n16022) );
  NAND U20439 ( .A(n15382), .B(creg[711]), .Z(n16021) );
  NAND U20440 ( .A(n16023), .B(n16024), .Z(y[710]) );
  NAND U20441 ( .A(n15381), .B(m[710]), .Z(n16024) );
  NAND U20442 ( .A(n15382), .B(creg[710]), .Z(n16023) );
  NAND U20443 ( .A(n16025), .B(n16026), .Z(y[70]) );
  NAND U20444 ( .A(n15381), .B(m[70]), .Z(n16026) );
  NAND U20445 ( .A(n15382), .B(creg[70]), .Z(n16025) );
  NAND U20446 ( .A(n16027), .B(n16028), .Z(y[709]) );
  NAND U20447 ( .A(n15381), .B(m[709]), .Z(n16028) );
  NAND U20448 ( .A(n15382), .B(creg[709]), .Z(n16027) );
  NAND U20449 ( .A(n16029), .B(n16030), .Z(y[708]) );
  NAND U20450 ( .A(n15381), .B(m[708]), .Z(n16030) );
  NAND U20451 ( .A(n15382), .B(creg[708]), .Z(n16029) );
  NAND U20452 ( .A(n16031), .B(n16032), .Z(y[707]) );
  NAND U20453 ( .A(n15381), .B(m[707]), .Z(n16032) );
  NAND U20454 ( .A(n15382), .B(creg[707]), .Z(n16031) );
  NAND U20455 ( .A(n16033), .B(n16034), .Z(y[706]) );
  NAND U20456 ( .A(n15381), .B(m[706]), .Z(n16034) );
  NAND U20457 ( .A(n15382), .B(creg[706]), .Z(n16033) );
  NAND U20458 ( .A(n16035), .B(n16036), .Z(y[705]) );
  NAND U20459 ( .A(n15381), .B(m[705]), .Z(n16036) );
  NAND U20460 ( .A(n15382), .B(creg[705]), .Z(n16035) );
  NAND U20461 ( .A(n16037), .B(n16038), .Z(y[704]) );
  NAND U20462 ( .A(n15381), .B(m[704]), .Z(n16038) );
  NAND U20463 ( .A(n15382), .B(creg[704]), .Z(n16037) );
  NAND U20464 ( .A(n16039), .B(n16040), .Z(y[703]) );
  NAND U20465 ( .A(n15381), .B(m[703]), .Z(n16040) );
  NAND U20466 ( .A(n15382), .B(creg[703]), .Z(n16039) );
  NAND U20467 ( .A(n16041), .B(n16042), .Z(y[702]) );
  NAND U20468 ( .A(n15381), .B(m[702]), .Z(n16042) );
  NAND U20469 ( .A(n15382), .B(creg[702]), .Z(n16041) );
  NAND U20470 ( .A(n16043), .B(n16044), .Z(y[701]) );
  NAND U20471 ( .A(n15381), .B(m[701]), .Z(n16044) );
  NAND U20472 ( .A(n15382), .B(creg[701]), .Z(n16043) );
  NAND U20473 ( .A(n16045), .B(n16046), .Z(y[700]) );
  NAND U20474 ( .A(n15381), .B(m[700]), .Z(n16046) );
  NAND U20475 ( .A(n15382), .B(creg[700]), .Z(n16045) );
  NAND U20476 ( .A(n16047), .B(n16048), .Z(y[6]) );
  NAND U20477 ( .A(n15381), .B(m[6]), .Z(n16048) );
  NAND U20478 ( .A(n15382), .B(creg[6]), .Z(n16047) );
  NAND U20479 ( .A(n16049), .B(n16050), .Z(y[69]) );
  NAND U20480 ( .A(n15381), .B(m[69]), .Z(n16050) );
  NAND U20481 ( .A(n15382), .B(creg[69]), .Z(n16049) );
  NAND U20482 ( .A(n16051), .B(n16052), .Z(y[699]) );
  NAND U20483 ( .A(n15381), .B(m[699]), .Z(n16052) );
  NAND U20484 ( .A(n15382), .B(creg[699]), .Z(n16051) );
  NAND U20485 ( .A(n16053), .B(n16054), .Z(y[698]) );
  NAND U20486 ( .A(n15381), .B(m[698]), .Z(n16054) );
  NAND U20487 ( .A(n15382), .B(creg[698]), .Z(n16053) );
  NAND U20488 ( .A(n16055), .B(n16056), .Z(y[697]) );
  NAND U20489 ( .A(n15381), .B(m[697]), .Z(n16056) );
  NAND U20490 ( .A(n15382), .B(creg[697]), .Z(n16055) );
  NAND U20491 ( .A(n16057), .B(n16058), .Z(y[696]) );
  NAND U20492 ( .A(n15381), .B(m[696]), .Z(n16058) );
  NAND U20493 ( .A(n15382), .B(creg[696]), .Z(n16057) );
  NAND U20494 ( .A(n16059), .B(n16060), .Z(y[695]) );
  NAND U20495 ( .A(n15381), .B(m[695]), .Z(n16060) );
  NAND U20496 ( .A(n15382), .B(creg[695]), .Z(n16059) );
  NAND U20497 ( .A(n16061), .B(n16062), .Z(y[694]) );
  NAND U20498 ( .A(n15381), .B(m[694]), .Z(n16062) );
  NAND U20499 ( .A(n15382), .B(creg[694]), .Z(n16061) );
  NAND U20500 ( .A(n16063), .B(n16064), .Z(y[693]) );
  NAND U20501 ( .A(n15381), .B(m[693]), .Z(n16064) );
  NAND U20502 ( .A(n15382), .B(creg[693]), .Z(n16063) );
  NAND U20503 ( .A(n16065), .B(n16066), .Z(y[692]) );
  NAND U20504 ( .A(n15381), .B(m[692]), .Z(n16066) );
  NAND U20505 ( .A(n15382), .B(creg[692]), .Z(n16065) );
  NAND U20506 ( .A(n16067), .B(n16068), .Z(y[691]) );
  NAND U20507 ( .A(n15381), .B(m[691]), .Z(n16068) );
  NAND U20508 ( .A(n15382), .B(creg[691]), .Z(n16067) );
  NAND U20509 ( .A(n16069), .B(n16070), .Z(y[690]) );
  NAND U20510 ( .A(n15381), .B(m[690]), .Z(n16070) );
  NAND U20511 ( .A(n15382), .B(creg[690]), .Z(n16069) );
  NAND U20512 ( .A(n16071), .B(n16072), .Z(y[68]) );
  NAND U20513 ( .A(n15381), .B(m[68]), .Z(n16072) );
  NAND U20514 ( .A(n15382), .B(creg[68]), .Z(n16071) );
  NAND U20515 ( .A(n16073), .B(n16074), .Z(y[689]) );
  NAND U20516 ( .A(n15381), .B(m[689]), .Z(n16074) );
  NAND U20517 ( .A(n15382), .B(creg[689]), .Z(n16073) );
  NAND U20518 ( .A(n16075), .B(n16076), .Z(y[688]) );
  NAND U20519 ( .A(n15381), .B(m[688]), .Z(n16076) );
  NAND U20520 ( .A(n15382), .B(creg[688]), .Z(n16075) );
  NAND U20521 ( .A(n16077), .B(n16078), .Z(y[687]) );
  NAND U20522 ( .A(n15381), .B(m[687]), .Z(n16078) );
  NAND U20523 ( .A(n15382), .B(creg[687]), .Z(n16077) );
  NAND U20524 ( .A(n16079), .B(n16080), .Z(y[686]) );
  NAND U20525 ( .A(n15381), .B(m[686]), .Z(n16080) );
  NAND U20526 ( .A(n15382), .B(creg[686]), .Z(n16079) );
  NAND U20527 ( .A(n16081), .B(n16082), .Z(y[685]) );
  NAND U20528 ( .A(n15381), .B(m[685]), .Z(n16082) );
  NAND U20529 ( .A(n15382), .B(creg[685]), .Z(n16081) );
  NAND U20530 ( .A(n16083), .B(n16084), .Z(y[684]) );
  NAND U20531 ( .A(n15381), .B(m[684]), .Z(n16084) );
  NAND U20532 ( .A(n15382), .B(creg[684]), .Z(n16083) );
  NAND U20533 ( .A(n16085), .B(n16086), .Z(y[683]) );
  NAND U20534 ( .A(n15381), .B(m[683]), .Z(n16086) );
  NAND U20535 ( .A(n15382), .B(creg[683]), .Z(n16085) );
  NAND U20536 ( .A(n16087), .B(n16088), .Z(y[682]) );
  NAND U20537 ( .A(n15381), .B(m[682]), .Z(n16088) );
  NAND U20538 ( .A(n15382), .B(creg[682]), .Z(n16087) );
  NAND U20539 ( .A(n16089), .B(n16090), .Z(y[681]) );
  NAND U20540 ( .A(n15381), .B(m[681]), .Z(n16090) );
  NAND U20541 ( .A(n15382), .B(creg[681]), .Z(n16089) );
  NAND U20542 ( .A(n16091), .B(n16092), .Z(y[680]) );
  NAND U20543 ( .A(n15381), .B(m[680]), .Z(n16092) );
  NAND U20544 ( .A(n15382), .B(creg[680]), .Z(n16091) );
  NAND U20545 ( .A(n16093), .B(n16094), .Z(y[67]) );
  NAND U20546 ( .A(n15381), .B(m[67]), .Z(n16094) );
  NAND U20547 ( .A(n15382), .B(creg[67]), .Z(n16093) );
  NAND U20548 ( .A(n16095), .B(n16096), .Z(y[679]) );
  NAND U20549 ( .A(n15381), .B(m[679]), .Z(n16096) );
  NAND U20550 ( .A(n15382), .B(creg[679]), .Z(n16095) );
  NAND U20551 ( .A(n16097), .B(n16098), .Z(y[678]) );
  NAND U20552 ( .A(n15381), .B(m[678]), .Z(n16098) );
  NAND U20553 ( .A(n15382), .B(creg[678]), .Z(n16097) );
  NAND U20554 ( .A(n16099), .B(n16100), .Z(y[677]) );
  NAND U20555 ( .A(n15381), .B(m[677]), .Z(n16100) );
  NAND U20556 ( .A(n15382), .B(creg[677]), .Z(n16099) );
  NAND U20557 ( .A(n16101), .B(n16102), .Z(y[676]) );
  NAND U20558 ( .A(n15381), .B(m[676]), .Z(n16102) );
  NAND U20559 ( .A(n15382), .B(creg[676]), .Z(n16101) );
  NAND U20560 ( .A(n16103), .B(n16104), .Z(y[675]) );
  NAND U20561 ( .A(n15381), .B(m[675]), .Z(n16104) );
  NAND U20562 ( .A(n15382), .B(creg[675]), .Z(n16103) );
  NAND U20563 ( .A(n16105), .B(n16106), .Z(y[674]) );
  NAND U20564 ( .A(n15381), .B(m[674]), .Z(n16106) );
  NAND U20565 ( .A(n15382), .B(creg[674]), .Z(n16105) );
  NAND U20566 ( .A(n16107), .B(n16108), .Z(y[673]) );
  NAND U20567 ( .A(n15381), .B(m[673]), .Z(n16108) );
  NAND U20568 ( .A(n15382), .B(creg[673]), .Z(n16107) );
  NAND U20569 ( .A(n16109), .B(n16110), .Z(y[672]) );
  NAND U20570 ( .A(n15381), .B(m[672]), .Z(n16110) );
  NAND U20571 ( .A(n15382), .B(creg[672]), .Z(n16109) );
  NAND U20572 ( .A(n16111), .B(n16112), .Z(y[671]) );
  NAND U20573 ( .A(n15381), .B(m[671]), .Z(n16112) );
  NAND U20574 ( .A(n15382), .B(creg[671]), .Z(n16111) );
  NAND U20575 ( .A(n16113), .B(n16114), .Z(y[670]) );
  NAND U20576 ( .A(n15381), .B(m[670]), .Z(n16114) );
  NAND U20577 ( .A(n15382), .B(creg[670]), .Z(n16113) );
  NAND U20578 ( .A(n16115), .B(n16116), .Z(y[66]) );
  NAND U20579 ( .A(n15381), .B(m[66]), .Z(n16116) );
  NAND U20580 ( .A(n15382), .B(creg[66]), .Z(n16115) );
  NAND U20581 ( .A(n16117), .B(n16118), .Z(y[669]) );
  NAND U20582 ( .A(n15381), .B(m[669]), .Z(n16118) );
  NAND U20583 ( .A(n15382), .B(creg[669]), .Z(n16117) );
  NAND U20584 ( .A(n16119), .B(n16120), .Z(y[668]) );
  NAND U20585 ( .A(n15381), .B(m[668]), .Z(n16120) );
  NAND U20586 ( .A(n15382), .B(creg[668]), .Z(n16119) );
  NAND U20587 ( .A(n16121), .B(n16122), .Z(y[667]) );
  NAND U20588 ( .A(n15381), .B(m[667]), .Z(n16122) );
  NAND U20589 ( .A(n15382), .B(creg[667]), .Z(n16121) );
  NAND U20590 ( .A(n16123), .B(n16124), .Z(y[666]) );
  NAND U20591 ( .A(n15381), .B(m[666]), .Z(n16124) );
  NAND U20592 ( .A(n15382), .B(creg[666]), .Z(n16123) );
  NAND U20593 ( .A(n16125), .B(n16126), .Z(y[665]) );
  NAND U20594 ( .A(n15381), .B(m[665]), .Z(n16126) );
  NAND U20595 ( .A(n15382), .B(creg[665]), .Z(n16125) );
  NAND U20596 ( .A(n16127), .B(n16128), .Z(y[664]) );
  NAND U20597 ( .A(n15381), .B(m[664]), .Z(n16128) );
  NAND U20598 ( .A(n15382), .B(creg[664]), .Z(n16127) );
  NAND U20599 ( .A(n16129), .B(n16130), .Z(y[663]) );
  NAND U20600 ( .A(n15381), .B(m[663]), .Z(n16130) );
  NAND U20601 ( .A(n15382), .B(creg[663]), .Z(n16129) );
  NAND U20602 ( .A(n16131), .B(n16132), .Z(y[662]) );
  NAND U20603 ( .A(n15381), .B(m[662]), .Z(n16132) );
  NAND U20604 ( .A(n15382), .B(creg[662]), .Z(n16131) );
  NAND U20605 ( .A(n16133), .B(n16134), .Z(y[661]) );
  NAND U20606 ( .A(n15381), .B(m[661]), .Z(n16134) );
  NAND U20607 ( .A(n15382), .B(creg[661]), .Z(n16133) );
  NAND U20608 ( .A(n16135), .B(n16136), .Z(y[660]) );
  NAND U20609 ( .A(n15381), .B(m[660]), .Z(n16136) );
  NAND U20610 ( .A(n15382), .B(creg[660]), .Z(n16135) );
  NAND U20611 ( .A(n16137), .B(n16138), .Z(y[65]) );
  NAND U20612 ( .A(n15381), .B(m[65]), .Z(n16138) );
  NAND U20613 ( .A(n15382), .B(creg[65]), .Z(n16137) );
  NAND U20614 ( .A(n16139), .B(n16140), .Z(y[659]) );
  NAND U20615 ( .A(n15381), .B(m[659]), .Z(n16140) );
  NAND U20616 ( .A(n15382), .B(creg[659]), .Z(n16139) );
  NAND U20617 ( .A(n16141), .B(n16142), .Z(y[658]) );
  NAND U20618 ( .A(n15381), .B(m[658]), .Z(n16142) );
  NAND U20619 ( .A(n15382), .B(creg[658]), .Z(n16141) );
  NAND U20620 ( .A(n16143), .B(n16144), .Z(y[657]) );
  NAND U20621 ( .A(n15381), .B(m[657]), .Z(n16144) );
  NAND U20622 ( .A(n15382), .B(creg[657]), .Z(n16143) );
  NAND U20623 ( .A(n16145), .B(n16146), .Z(y[656]) );
  NAND U20624 ( .A(n15381), .B(m[656]), .Z(n16146) );
  NAND U20625 ( .A(n15382), .B(creg[656]), .Z(n16145) );
  NAND U20626 ( .A(n16147), .B(n16148), .Z(y[655]) );
  NAND U20627 ( .A(n15381), .B(m[655]), .Z(n16148) );
  NAND U20628 ( .A(n15382), .B(creg[655]), .Z(n16147) );
  NAND U20629 ( .A(n16149), .B(n16150), .Z(y[654]) );
  NAND U20630 ( .A(n15381), .B(m[654]), .Z(n16150) );
  NAND U20631 ( .A(n15382), .B(creg[654]), .Z(n16149) );
  NAND U20632 ( .A(n16151), .B(n16152), .Z(y[653]) );
  NAND U20633 ( .A(n15381), .B(m[653]), .Z(n16152) );
  NAND U20634 ( .A(n15382), .B(creg[653]), .Z(n16151) );
  NAND U20635 ( .A(n16153), .B(n16154), .Z(y[652]) );
  NAND U20636 ( .A(n15381), .B(m[652]), .Z(n16154) );
  NAND U20637 ( .A(n15382), .B(creg[652]), .Z(n16153) );
  NAND U20638 ( .A(n16155), .B(n16156), .Z(y[651]) );
  NAND U20639 ( .A(n15381), .B(m[651]), .Z(n16156) );
  NAND U20640 ( .A(n15382), .B(creg[651]), .Z(n16155) );
  NAND U20641 ( .A(n16157), .B(n16158), .Z(y[650]) );
  NAND U20642 ( .A(n15381), .B(m[650]), .Z(n16158) );
  NAND U20643 ( .A(n15382), .B(creg[650]), .Z(n16157) );
  NAND U20644 ( .A(n16159), .B(n16160), .Z(y[64]) );
  NAND U20645 ( .A(n15381), .B(m[64]), .Z(n16160) );
  NAND U20646 ( .A(n15382), .B(creg[64]), .Z(n16159) );
  NAND U20647 ( .A(n16161), .B(n16162), .Z(y[649]) );
  NAND U20648 ( .A(n15381), .B(m[649]), .Z(n16162) );
  NAND U20649 ( .A(n15382), .B(creg[649]), .Z(n16161) );
  NAND U20650 ( .A(n16163), .B(n16164), .Z(y[648]) );
  NAND U20651 ( .A(n15381), .B(m[648]), .Z(n16164) );
  NAND U20652 ( .A(n15382), .B(creg[648]), .Z(n16163) );
  NAND U20653 ( .A(n16165), .B(n16166), .Z(y[647]) );
  NAND U20654 ( .A(n15381), .B(m[647]), .Z(n16166) );
  NAND U20655 ( .A(n15382), .B(creg[647]), .Z(n16165) );
  NAND U20656 ( .A(n16167), .B(n16168), .Z(y[646]) );
  NAND U20657 ( .A(n15381), .B(m[646]), .Z(n16168) );
  NAND U20658 ( .A(n15382), .B(creg[646]), .Z(n16167) );
  NAND U20659 ( .A(n16169), .B(n16170), .Z(y[645]) );
  NAND U20660 ( .A(n15381), .B(m[645]), .Z(n16170) );
  NAND U20661 ( .A(n15382), .B(creg[645]), .Z(n16169) );
  NAND U20662 ( .A(n16171), .B(n16172), .Z(y[644]) );
  NAND U20663 ( .A(n15381), .B(m[644]), .Z(n16172) );
  NAND U20664 ( .A(n15382), .B(creg[644]), .Z(n16171) );
  NAND U20665 ( .A(n16173), .B(n16174), .Z(y[643]) );
  NAND U20666 ( .A(n15381), .B(m[643]), .Z(n16174) );
  NAND U20667 ( .A(n15382), .B(creg[643]), .Z(n16173) );
  NAND U20668 ( .A(n16175), .B(n16176), .Z(y[642]) );
  NAND U20669 ( .A(n15381), .B(m[642]), .Z(n16176) );
  NAND U20670 ( .A(n15382), .B(creg[642]), .Z(n16175) );
  NAND U20671 ( .A(n16177), .B(n16178), .Z(y[641]) );
  NAND U20672 ( .A(n15381), .B(m[641]), .Z(n16178) );
  NAND U20673 ( .A(n15382), .B(creg[641]), .Z(n16177) );
  NAND U20674 ( .A(n16179), .B(n16180), .Z(y[640]) );
  NAND U20675 ( .A(n15381), .B(m[640]), .Z(n16180) );
  NAND U20676 ( .A(n15382), .B(creg[640]), .Z(n16179) );
  NAND U20677 ( .A(n16181), .B(n16182), .Z(y[63]) );
  NAND U20678 ( .A(n15381), .B(m[63]), .Z(n16182) );
  NAND U20679 ( .A(n15382), .B(creg[63]), .Z(n16181) );
  NAND U20680 ( .A(n16183), .B(n16184), .Z(y[639]) );
  NAND U20681 ( .A(n15381), .B(m[639]), .Z(n16184) );
  NAND U20682 ( .A(n15382), .B(creg[639]), .Z(n16183) );
  NAND U20683 ( .A(n16185), .B(n16186), .Z(y[638]) );
  NAND U20684 ( .A(n15381), .B(m[638]), .Z(n16186) );
  NAND U20685 ( .A(n15382), .B(creg[638]), .Z(n16185) );
  NAND U20686 ( .A(n16187), .B(n16188), .Z(y[637]) );
  NAND U20687 ( .A(n15381), .B(m[637]), .Z(n16188) );
  NAND U20688 ( .A(n15382), .B(creg[637]), .Z(n16187) );
  NAND U20689 ( .A(n16189), .B(n16190), .Z(y[636]) );
  NAND U20690 ( .A(n15381), .B(m[636]), .Z(n16190) );
  NAND U20691 ( .A(n15382), .B(creg[636]), .Z(n16189) );
  NAND U20692 ( .A(n16191), .B(n16192), .Z(y[635]) );
  NAND U20693 ( .A(n15381), .B(m[635]), .Z(n16192) );
  NAND U20694 ( .A(n15382), .B(creg[635]), .Z(n16191) );
  NAND U20695 ( .A(n16193), .B(n16194), .Z(y[634]) );
  NAND U20696 ( .A(n15381), .B(m[634]), .Z(n16194) );
  NAND U20697 ( .A(n15382), .B(creg[634]), .Z(n16193) );
  NAND U20698 ( .A(n16195), .B(n16196), .Z(y[633]) );
  NAND U20699 ( .A(n15381), .B(m[633]), .Z(n16196) );
  NAND U20700 ( .A(n15382), .B(creg[633]), .Z(n16195) );
  NAND U20701 ( .A(n16197), .B(n16198), .Z(y[632]) );
  NAND U20702 ( .A(n15381), .B(m[632]), .Z(n16198) );
  NAND U20703 ( .A(n15382), .B(creg[632]), .Z(n16197) );
  NAND U20704 ( .A(n16199), .B(n16200), .Z(y[631]) );
  NAND U20705 ( .A(n15381), .B(m[631]), .Z(n16200) );
  NAND U20706 ( .A(n15382), .B(creg[631]), .Z(n16199) );
  NAND U20707 ( .A(n16201), .B(n16202), .Z(y[630]) );
  NAND U20708 ( .A(n15381), .B(m[630]), .Z(n16202) );
  NAND U20709 ( .A(n15382), .B(creg[630]), .Z(n16201) );
  NAND U20710 ( .A(n16203), .B(n16204), .Z(y[62]) );
  NAND U20711 ( .A(n15381), .B(m[62]), .Z(n16204) );
  NAND U20712 ( .A(n15382), .B(creg[62]), .Z(n16203) );
  NAND U20713 ( .A(n16205), .B(n16206), .Z(y[629]) );
  NAND U20714 ( .A(n15381), .B(m[629]), .Z(n16206) );
  NAND U20715 ( .A(n15382), .B(creg[629]), .Z(n16205) );
  NAND U20716 ( .A(n16207), .B(n16208), .Z(y[628]) );
  NAND U20717 ( .A(n15381), .B(m[628]), .Z(n16208) );
  NAND U20718 ( .A(n15382), .B(creg[628]), .Z(n16207) );
  NAND U20719 ( .A(n16209), .B(n16210), .Z(y[627]) );
  NAND U20720 ( .A(n15381), .B(m[627]), .Z(n16210) );
  NAND U20721 ( .A(n15382), .B(creg[627]), .Z(n16209) );
  NAND U20722 ( .A(n16211), .B(n16212), .Z(y[626]) );
  NAND U20723 ( .A(n15381), .B(m[626]), .Z(n16212) );
  NAND U20724 ( .A(n15382), .B(creg[626]), .Z(n16211) );
  NAND U20725 ( .A(n16213), .B(n16214), .Z(y[625]) );
  NAND U20726 ( .A(n15381), .B(m[625]), .Z(n16214) );
  NAND U20727 ( .A(n15382), .B(creg[625]), .Z(n16213) );
  NAND U20728 ( .A(n16215), .B(n16216), .Z(y[624]) );
  NAND U20729 ( .A(n15381), .B(m[624]), .Z(n16216) );
  NAND U20730 ( .A(n15382), .B(creg[624]), .Z(n16215) );
  NAND U20731 ( .A(n16217), .B(n16218), .Z(y[623]) );
  NAND U20732 ( .A(n15381), .B(m[623]), .Z(n16218) );
  NAND U20733 ( .A(n15382), .B(creg[623]), .Z(n16217) );
  NAND U20734 ( .A(n16219), .B(n16220), .Z(y[622]) );
  NAND U20735 ( .A(n15381), .B(m[622]), .Z(n16220) );
  NAND U20736 ( .A(n15382), .B(creg[622]), .Z(n16219) );
  NAND U20737 ( .A(n16221), .B(n16222), .Z(y[621]) );
  NAND U20738 ( .A(n15381), .B(m[621]), .Z(n16222) );
  NAND U20739 ( .A(n15382), .B(creg[621]), .Z(n16221) );
  NAND U20740 ( .A(n16223), .B(n16224), .Z(y[620]) );
  NAND U20741 ( .A(n15381), .B(m[620]), .Z(n16224) );
  NAND U20742 ( .A(n15382), .B(creg[620]), .Z(n16223) );
  NAND U20743 ( .A(n16225), .B(n16226), .Z(y[61]) );
  NAND U20744 ( .A(n15381), .B(m[61]), .Z(n16226) );
  NAND U20745 ( .A(n15382), .B(creg[61]), .Z(n16225) );
  NAND U20746 ( .A(n16227), .B(n16228), .Z(y[619]) );
  NAND U20747 ( .A(n15381), .B(m[619]), .Z(n16228) );
  NAND U20748 ( .A(n15382), .B(creg[619]), .Z(n16227) );
  NAND U20749 ( .A(n16229), .B(n16230), .Z(y[618]) );
  NAND U20750 ( .A(n15381), .B(m[618]), .Z(n16230) );
  NAND U20751 ( .A(n15382), .B(creg[618]), .Z(n16229) );
  NAND U20752 ( .A(n16231), .B(n16232), .Z(y[617]) );
  NAND U20753 ( .A(n15381), .B(m[617]), .Z(n16232) );
  NAND U20754 ( .A(n15382), .B(creg[617]), .Z(n16231) );
  NAND U20755 ( .A(n16233), .B(n16234), .Z(y[616]) );
  NAND U20756 ( .A(n15381), .B(m[616]), .Z(n16234) );
  NAND U20757 ( .A(n15382), .B(creg[616]), .Z(n16233) );
  NAND U20758 ( .A(n16235), .B(n16236), .Z(y[615]) );
  NAND U20759 ( .A(n15381), .B(m[615]), .Z(n16236) );
  NAND U20760 ( .A(n15382), .B(creg[615]), .Z(n16235) );
  NAND U20761 ( .A(n16237), .B(n16238), .Z(y[614]) );
  NAND U20762 ( .A(n15381), .B(m[614]), .Z(n16238) );
  NAND U20763 ( .A(n15382), .B(creg[614]), .Z(n16237) );
  NAND U20764 ( .A(n16239), .B(n16240), .Z(y[613]) );
  NAND U20765 ( .A(n15381), .B(m[613]), .Z(n16240) );
  NAND U20766 ( .A(n15382), .B(creg[613]), .Z(n16239) );
  NAND U20767 ( .A(n16241), .B(n16242), .Z(y[612]) );
  NAND U20768 ( .A(n15381), .B(m[612]), .Z(n16242) );
  NAND U20769 ( .A(n15382), .B(creg[612]), .Z(n16241) );
  NAND U20770 ( .A(n16243), .B(n16244), .Z(y[611]) );
  NAND U20771 ( .A(n15381), .B(m[611]), .Z(n16244) );
  NAND U20772 ( .A(n15382), .B(creg[611]), .Z(n16243) );
  NAND U20773 ( .A(n16245), .B(n16246), .Z(y[610]) );
  NAND U20774 ( .A(n15381), .B(m[610]), .Z(n16246) );
  NAND U20775 ( .A(n15382), .B(creg[610]), .Z(n16245) );
  NAND U20776 ( .A(n16247), .B(n16248), .Z(y[60]) );
  NAND U20777 ( .A(n15381), .B(m[60]), .Z(n16248) );
  NAND U20778 ( .A(n15382), .B(creg[60]), .Z(n16247) );
  NAND U20779 ( .A(n16249), .B(n16250), .Z(y[609]) );
  NAND U20780 ( .A(n15381), .B(m[609]), .Z(n16250) );
  NAND U20781 ( .A(n15382), .B(creg[609]), .Z(n16249) );
  NAND U20782 ( .A(n16251), .B(n16252), .Z(y[608]) );
  NAND U20783 ( .A(n15381), .B(m[608]), .Z(n16252) );
  NAND U20784 ( .A(n15382), .B(creg[608]), .Z(n16251) );
  NAND U20785 ( .A(n16253), .B(n16254), .Z(y[607]) );
  NAND U20786 ( .A(n15381), .B(m[607]), .Z(n16254) );
  NAND U20787 ( .A(n15382), .B(creg[607]), .Z(n16253) );
  NAND U20788 ( .A(n16255), .B(n16256), .Z(y[606]) );
  NAND U20789 ( .A(n15381), .B(m[606]), .Z(n16256) );
  NAND U20790 ( .A(n15382), .B(creg[606]), .Z(n16255) );
  NAND U20791 ( .A(n16257), .B(n16258), .Z(y[605]) );
  NAND U20792 ( .A(n15381), .B(m[605]), .Z(n16258) );
  NAND U20793 ( .A(n15382), .B(creg[605]), .Z(n16257) );
  NAND U20794 ( .A(n16259), .B(n16260), .Z(y[604]) );
  NAND U20795 ( .A(n15381), .B(m[604]), .Z(n16260) );
  NAND U20796 ( .A(n15382), .B(creg[604]), .Z(n16259) );
  NAND U20797 ( .A(n16261), .B(n16262), .Z(y[603]) );
  NAND U20798 ( .A(n15381), .B(m[603]), .Z(n16262) );
  NAND U20799 ( .A(n15382), .B(creg[603]), .Z(n16261) );
  NAND U20800 ( .A(n16263), .B(n16264), .Z(y[602]) );
  NAND U20801 ( .A(n15381), .B(m[602]), .Z(n16264) );
  NAND U20802 ( .A(n15382), .B(creg[602]), .Z(n16263) );
  NAND U20803 ( .A(n16265), .B(n16266), .Z(y[601]) );
  NAND U20804 ( .A(n15381), .B(m[601]), .Z(n16266) );
  NAND U20805 ( .A(n15382), .B(creg[601]), .Z(n16265) );
  NAND U20806 ( .A(n16267), .B(n16268), .Z(y[600]) );
  NAND U20807 ( .A(n15381), .B(m[600]), .Z(n16268) );
  NAND U20808 ( .A(n15382), .B(creg[600]), .Z(n16267) );
  NAND U20809 ( .A(n16269), .B(n16270), .Z(y[5]) );
  NAND U20810 ( .A(n15381), .B(m[5]), .Z(n16270) );
  NAND U20811 ( .A(n15382), .B(creg[5]), .Z(n16269) );
  NAND U20812 ( .A(n16271), .B(n16272), .Z(y[59]) );
  NAND U20813 ( .A(n15381), .B(m[59]), .Z(n16272) );
  NAND U20814 ( .A(n15382), .B(creg[59]), .Z(n16271) );
  NAND U20815 ( .A(n16273), .B(n16274), .Z(y[599]) );
  NAND U20816 ( .A(n15381), .B(m[599]), .Z(n16274) );
  NAND U20817 ( .A(n15382), .B(creg[599]), .Z(n16273) );
  NAND U20818 ( .A(n16275), .B(n16276), .Z(y[598]) );
  NAND U20819 ( .A(n15381), .B(m[598]), .Z(n16276) );
  NAND U20820 ( .A(n15382), .B(creg[598]), .Z(n16275) );
  NAND U20821 ( .A(n16277), .B(n16278), .Z(y[597]) );
  NAND U20822 ( .A(n15381), .B(m[597]), .Z(n16278) );
  NAND U20823 ( .A(n15382), .B(creg[597]), .Z(n16277) );
  NAND U20824 ( .A(n16279), .B(n16280), .Z(y[596]) );
  NAND U20825 ( .A(n15381), .B(m[596]), .Z(n16280) );
  NAND U20826 ( .A(n15382), .B(creg[596]), .Z(n16279) );
  NAND U20827 ( .A(n16281), .B(n16282), .Z(y[595]) );
  NAND U20828 ( .A(n15381), .B(m[595]), .Z(n16282) );
  NAND U20829 ( .A(n15382), .B(creg[595]), .Z(n16281) );
  NAND U20830 ( .A(n16283), .B(n16284), .Z(y[594]) );
  NAND U20831 ( .A(n15381), .B(m[594]), .Z(n16284) );
  NAND U20832 ( .A(n15382), .B(creg[594]), .Z(n16283) );
  NAND U20833 ( .A(n16285), .B(n16286), .Z(y[593]) );
  NAND U20834 ( .A(n15381), .B(m[593]), .Z(n16286) );
  NAND U20835 ( .A(n15382), .B(creg[593]), .Z(n16285) );
  NAND U20836 ( .A(n16287), .B(n16288), .Z(y[592]) );
  NAND U20837 ( .A(n15381), .B(m[592]), .Z(n16288) );
  NAND U20838 ( .A(n15382), .B(creg[592]), .Z(n16287) );
  NAND U20839 ( .A(n16289), .B(n16290), .Z(y[591]) );
  NAND U20840 ( .A(n15381), .B(m[591]), .Z(n16290) );
  NAND U20841 ( .A(n15382), .B(creg[591]), .Z(n16289) );
  NAND U20842 ( .A(n16291), .B(n16292), .Z(y[590]) );
  NAND U20843 ( .A(n15381), .B(m[590]), .Z(n16292) );
  NAND U20844 ( .A(n15382), .B(creg[590]), .Z(n16291) );
  NAND U20845 ( .A(n16293), .B(n16294), .Z(y[58]) );
  NAND U20846 ( .A(n15381), .B(m[58]), .Z(n16294) );
  NAND U20847 ( .A(n15382), .B(creg[58]), .Z(n16293) );
  NAND U20848 ( .A(n16295), .B(n16296), .Z(y[589]) );
  NAND U20849 ( .A(n15381), .B(m[589]), .Z(n16296) );
  NAND U20850 ( .A(n15382), .B(creg[589]), .Z(n16295) );
  NAND U20851 ( .A(n16297), .B(n16298), .Z(y[588]) );
  NAND U20852 ( .A(n15381), .B(m[588]), .Z(n16298) );
  NAND U20853 ( .A(n15382), .B(creg[588]), .Z(n16297) );
  NAND U20854 ( .A(n16299), .B(n16300), .Z(y[587]) );
  NAND U20855 ( .A(n15381), .B(m[587]), .Z(n16300) );
  NAND U20856 ( .A(n15382), .B(creg[587]), .Z(n16299) );
  NAND U20857 ( .A(n16301), .B(n16302), .Z(y[586]) );
  NAND U20858 ( .A(n15381), .B(m[586]), .Z(n16302) );
  NAND U20859 ( .A(n15382), .B(creg[586]), .Z(n16301) );
  NAND U20860 ( .A(n16303), .B(n16304), .Z(y[585]) );
  NAND U20861 ( .A(n15381), .B(m[585]), .Z(n16304) );
  NAND U20862 ( .A(n15382), .B(creg[585]), .Z(n16303) );
  NAND U20863 ( .A(n16305), .B(n16306), .Z(y[584]) );
  NAND U20864 ( .A(n15381), .B(m[584]), .Z(n16306) );
  NAND U20865 ( .A(n15382), .B(creg[584]), .Z(n16305) );
  NAND U20866 ( .A(n16307), .B(n16308), .Z(y[583]) );
  NAND U20867 ( .A(n15381), .B(m[583]), .Z(n16308) );
  NAND U20868 ( .A(n15382), .B(creg[583]), .Z(n16307) );
  NAND U20869 ( .A(n16309), .B(n16310), .Z(y[582]) );
  NAND U20870 ( .A(n15381), .B(m[582]), .Z(n16310) );
  NAND U20871 ( .A(n15382), .B(creg[582]), .Z(n16309) );
  NAND U20872 ( .A(n16311), .B(n16312), .Z(y[581]) );
  NAND U20873 ( .A(n15381), .B(m[581]), .Z(n16312) );
  NAND U20874 ( .A(n15382), .B(creg[581]), .Z(n16311) );
  NAND U20875 ( .A(n16313), .B(n16314), .Z(y[580]) );
  NAND U20876 ( .A(n15381), .B(m[580]), .Z(n16314) );
  NAND U20877 ( .A(n15382), .B(creg[580]), .Z(n16313) );
  NAND U20878 ( .A(n16315), .B(n16316), .Z(y[57]) );
  NAND U20879 ( .A(n15381), .B(m[57]), .Z(n16316) );
  NAND U20880 ( .A(n15382), .B(creg[57]), .Z(n16315) );
  NAND U20881 ( .A(n16317), .B(n16318), .Z(y[579]) );
  NAND U20882 ( .A(n15381), .B(m[579]), .Z(n16318) );
  NAND U20883 ( .A(n15382), .B(creg[579]), .Z(n16317) );
  NAND U20884 ( .A(n16319), .B(n16320), .Z(y[578]) );
  NAND U20885 ( .A(n15381), .B(m[578]), .Z(n16320) );
  NAND U20886 ( .A(n15382), .B(creg[578]), .Z(n16319) );
  NAND U20887 ( .A(n16321), .B(n16322), .Z(y[577]) );
  NAND U20888 ( .A(n15381), .B(m[577]), .Z(n16322) );
  NAND U20889 ( .A(n15382), .B(creg[577]), .Z(n16321) );
  NAND U20890 ( .A(n16323), .B(n16324), .Z(y[576]) );
  NAND U20891 ( .A(n15381), .B(m[576]), .Z(n16324) );
  NAND U20892 ( .A(n15382), .B(creg[576]), .Z(n16323) );
  NAND U20893 ( .A(n16325), .B(n16326), .Z(y[575]) );
  NAND U20894 ( .A(n15381), .B(m[575]), .Z(n16326) );
  NAND U20895 ( .A(n15382), .B(creg[575]), .Z(n16325) );
  NAND U20896 ( .A(n16327), .B(n16328), .Z(y[574]) );
  NAND U20897 ( .A(n15381), .B(m[574]), .Z(n16328) );
  NAND U20898 ( .A(n15382), .B(creg[574]), .Z(n16327) );
  NAND U20899 ( .A(n16329), .B(n16330), .Z(y[573]) );
  NAND U20900 ( .A(n15381), .B(m[573]), .Z(n16330) );
  NAND U20901 ( .A(n15382), .B(creg[573]), .Z(n16329) );
  NAND U20902 ( .A(n16331), .B(n16332), .Z(y[572]) );
  NAND U20903 ( .A(n15381), .B(m[572]), .Z(n16332) );
  NAND U20904 ( .A(n15382), .B(creg[572]), .Z(n16331) );
  NAND U20905 ( .A(n16333), .B(n16334), .Z(y[571]) );
  NAND U20906 ( .A(n15381), .B(m[571]), .Z(n16334) );
  NAND U20907 ( .A(n15382), .B(creg[571]), .Z(n16333) );
  NAND U20908 ( .A(n16335), .B(n16336), .Z(y[570]) );
  NAND U20909 ( .A(n15381), .B(m[570]), .Z(n16336) );
  NAND U20910 ( .A(n15382), .B(creg[570]), .Z(n16335) );
  NAND U20911 ( .A(n16337), .B(n16338), .Z(y[56]) );
  NAND U20912 ( .A(n15381), .B(m[56]), .Z(n16338) );
  NAND U20913 ( .A(n15382), .B(creg[56]), .Z(n16337) );
  NAND U20914 ( .A(n16339), .B(n16340), .Z(y[569]) );
  NAND U20915 ( .A(n15381), .B(m[569]), .Z(n16340) );
  NAND U20916 ( .A(n15382), .B(creg[569]), .Z(n16339) );
  NAND U20917 ( .A(n16341), .B(n16342), .Z(y[568]) );
  NAND U20918 ( .A(n15381), .B(m[568]), .Z(n16342) );
  NAND U20919 ( .A(n15382), .B(creg[568]), .Z(n16341) );
  NAND U20920 ( .A(n16343), .B(n16344), .Z(y[567]) );
  NAND U20921 ( .A(n15381), .B(m[567]), .Z(n16344) );
  NAND U20922 ( .A(n15382), .B(creg[567]), .Z(n16343) );
  NAND U20923 ( .A(n16345), .B(n16346), .Z(y[566]) );
  NAND U20924 ( .A(n15381), .B(m[566]), .Z(n16346) );
  NAND U20925 ( .A(n15382), .B(creg[566]), .Z(n16345) );
  NAND U20926 ( .A(n16347), .B(n16348), .Z(y[565]) );
  NAND U20927 ( .A(n15381), .B(m[565]), .Z(n16348) );
  NAND U20928 ( .A(n15382), .B(creg[565]), .Z(n16347) );
  NAND U20929 ( .A(n16349), .B(n16350), .Z(y[564]) );
  NAND U20930 ( .A(n15381), .B(m[564]), .Z(n16350) );
  NAND U20931 ( .A(n15382), .B(creg[564]), .Z(n16349) );
  NAND U20932 ( .A(n16351), .B(n16352), .Z(y[563]) );
  NAND U20933 ( .A(n15381), .B(m[563]), .Z(n16352) );
  NAND U20934 ( .A(n15382), .B(creg[563]), .Z(n16351) );
  NAND U20935 ( .A(n16353), .B(n16354), .Z(y[562]) );
  NAND U20936 ( .A(n15381), .B(m[562]), .Z(n16354) );
  NAND U20937 ( .A(n15382), .B(creg[562]), .Z(n16353) );
  NAND U20938 ( .A(n16355), .B(n16356), .Z(y[561]) );
  NAND U20939 ( .A(n15381), .B(m[561]), .Z(n16356) );
  NAND U20940 ( .A(n15382), .B(creg[561]), .Z(n16355) );
  NAND U20941 ( .A(n16357), .B(n16358), .Z(y[560]) );
  NAND U20942 ( .A(n15381), .B(m[560]), .Z(n16358) );
  NAND U20943 ( .A(n15382), .B(creg[560]), .Z(n16357) );
  NAND U20944 ( .A(n16359), .B(n16360), .Z(y[55]) );
  NAND U20945 ( .A(n15381), .B(m[55]), .Z(n16360) );
  NAND U20946 ( .A(n15382), .B(creg[55]), .Z(n16359) );
  NAND U20947 ( .A(n16361), .B(n16362), .Z(y[559]) );
  NAND U20948 ( .A(n15381), .B(m[559]), .Z(n16362) );
  NAND U20949 ( .A(n15382), .B(creg[559]), .Z(n16361) );
  NAND U20950 ( .A(n16363), .B(n16364), .Z(y[558]) );
  NAND U20951 ( .A(n15381), .B(m[558]), .Z(n16364) );
  NAND U20952 ( .A(n15382), .B(creg[558]), .Z(n16363) );
  NAND U20953 ( .A(n16365), .B(n16366), .Z(y[557]) );
  NAND U20954 ( .A(n15381), .B(m[557]), .Z(n16366) );
  NAND U20955 ( .A(n15382), .B(creg[557]), .Z(n16365) );
  NAND U20956 ( .A(n16367), .B(n16368), .Z(y[556]) );
  NAND U20957 ( .A(n15381), .B(m[556]), .Z(n16368) );
  NAND U20958 ( .A(n15382), .B(creg[556]), .Z(n16367) );
  NAND U20959 ( .A(n16369), .B(n16370), .Z(y[555]) );
  NAND U20960 ( .A(n15381), .B(m[555]), .Z(n16370) );
  NAND U20961 ( .A(n15382), .B(creg[555]), .Z(n16369) );
  NAND U20962 ( .A(n16371), .B(n16372), .Z(y[554]) );
  NAND U20963 ( .A(n15381), .B(m[554]), .Z(n16372) );
  NAND U20964 ( .A(n15382), .B(creg[554]), .Z(n16371) );
  NAND U20965 ( .A(n16373), .B(n16374), .Z(y[553]) );
  NAND U20966 ( .A(n15381), .B(m[553]), .Z(n16374) );
  NAND U20967 ( .A(n15382), .B(creg[553]), .Z(n16373) );
  NAND U20968 ( .A(n16375), .B(n16376), .Z(y[552]) );
  NAND U20969 ( .A(n15381), .B(m[552]), .Z(n16376) );
  NAND U20970 ( .A(n15382), .B(creg[552]), .Z(n16375) );
  NAND U20971 ( .A(n16377), .B(n16378), .Z(y[551]) );
  NAND U20972 ( .A(n15381), .B(m[551]), .Z(n16378) );
  NAND U20973 ( .A(n15382), .B(creg[551]), .Z(n16377) );
  NAND U20974 ( .A(n16379), .B(n16380), .Z(y[550]) );
  NAND U20975 ( .A(n15381), .B(m[550]), .Z(n16380) );
  NAND U20976 ( .A(n15382), .B(creg[550]), .Z(n16379) );
  NAND U20977 ( .A(n16381), .B(n16382), .Z(y[54]) );
  NAND U20978 ( .A(n15381), .B(m[54]), .Z(n16382) );
  NAND U20979 ( .A(n15382), .B(creg[54]), .Z(n16381) );
  NAND U20980 ( .A(n16383), .B(n16384), .Z(y[549]) );
  NAND U20981 ( .A(n15381), .B(m[549]), .Z(n16384) );
  NAND U20982 ( .A(n15382), .B(creg[549]), .Z(n16383) );
  NAND U20983 ( .A(n16385), .B(n16386), .Z(y[548]) );
  NAND U20984 ( .A(n15381), .B(m[548]), .Z(n16386) );
  NAND U20985 ( .A(n15382), .B(creg[548]), .Z(n16385) );
  NAND U20986 ( .A(n16387), .B(n16388), .Z(y[547]) );
  NAND U20987 ( .A(n15381), .B(m[547]), .Z(n16388) );
  NAND U20988 ( .A(n15382), .B(creg[547]), .Z(n16387) );
  NAND U20989 ( .A(n16389), .B(n16390), .Z(y[546]) );
  NAND U20990 ( .A(n15381), .B(m[546]), .Z(n16390) );
  NAND U20991 ( .A(n15382), .B(creg[546]), .Z(n16389) );
  NAND U20992 ( .A(n16391), .B(n16392), .Z(y[545]) );
  NAND U20993 ( .A(n15381), .B(m[545]), .Z(n16392) );
  NAND U20994 ( .A(n15382), .B(creg[545]), .Z(n16391) );
  NAND U20995 ( .A(n16393), .B(n16394), .Z(y[544]) );
  NAND U20996 ( .A(n15381), .B(m[544]), .Z(n16394) );
  NAND U20997 ( .A(n15382), .B(creg[544]), .Z(n16393) );
  NAND U20998 ( .A(n16395), .B(n16396), .Z(y[543]) );
  NAND U20999 ( .A(n15381), .B(m[543]), .Z(n16396) );
  NAND U21000 ( .A(n15382), .B(creg[543]), .Z(n16395) );
  NAND U21001 ( .A(n16397), .B(n16398), .Z(y[542]) );
  NAND U21002 ( .A(n15381), .B(m[542]), .Z(n16398) );
  NAND U21003 ( .A(n15382), .B(creg[542]), .Z(n16397) );
  NAND U21004 ( .A(n16399), .B(n16400), .Z(y[541]) );
  NAND U21005 ( .A(n15381), .B(m[541]), .Z(n16400) );
  NAND U21006 ( .A(n15382), .B(creg[541]), .Z(n16399) );
  NAND U21007 ( .A(n16401), .B(n16402), .Z(y[540]) );
  NAND U21008 ( .A(n15381), .B(m[540]), .Z(n16402) );
  NAND U21009 ( .A(n15382), .B(creg[540]), .Z(n16401) );
  NAND U21010 ( .A(n16403), .B(n16404), .Z(y[53]) );
  NAND U21011 ( .A(n15381), .B(m[53]), .Z(n16404) );
  NAND U21012 ( .A(n15382), .B(creg[53]), .Z(n16403) );
  NAND U21013 ( .A(n16405), .B(n16406), .Z(y[539]) );
  NAND U21014 ( .A(n15381), .B(m[539]), .Z(n16406) );
  NAND U21015 ( .A(n15382), .B(creg[539]), .Z(n16405) );
  NAND U21016 ( .A(n16407), .B(n16408), .Z(y[538]) );
  NAND U21017 ( .A(n15381), .B(m[538]), .Z(n16408) );
  NAND U21018 ( .A(n15382), .B(creg[538]), .Z(n16407) );
  NAND U21019 ( .A(n16409), .B(n16410), .Z(y[537]) );
  NAND U21020 ( .A(n15381), .B(m[537]), .Z(n16410) );
  NAND U21021 ( .A(n15382), .B(creg[537]), .Z(n16409) );
  NAND U21022 ( .A(n16411), .B(n16412), .Z(y[536]) );
  NAND U21023 ( .A(n15381), .B(m[536]), .Z(n16412) );
  NAND U21024 ( .A(n15382), .B(creg[536]), .Z(n16411) );
  NAND U21025 ( .A(n16413), .B(n16414), .Z(y[535]) );
  NAND U21026 ( .A(n15381), .B(m[535]), .Z(n16414) );
  NAND U21027 ( .A(n15382), .B(creg[535]), .Z(n16413) );
  NAND U21028 ( .A(n16415), .B(n16416), .Z(y[534]) );
  NAND U21029 ( .A(n15381), .B(m[534]), .Z(n16416) );
  NAND U21030 ( .A(n15382), .B(creg[534]), .Z(n16415) );
  NAND U21031 ( .A(n16417), .B(n16418), .Z(y[533]) );
  NAND U21032 ( .A(n15381), .B(m[533]), .Z(n16418) );
  NAND U21033 ( .A(n15382), .B(creg[533]), .Z(n16417) );
  NAND U21034 ( .A(n16419), .B(n16420), .Z(y[532]) );
  NAND U21035 ( .A(n15381), .B(m[532]), .Z(n16420) );
  NAND U21036 ( .A(n15382), .B(creg[532]), .Z(n16419) );
  NAND U21037 ( .A(n16421), .B(n16422), .Z(y[531]) );
  NAND U21038 ( .A(n15381), .B(m[531]), .Z(n16422) );
  NAND U21039 ( .A(n15382), .B(creg[531]), .Z(n16421) );
  NAND U21040 ( .A(n16423), .B(n16424), .Z(y[530]) );
  NAND U21041 ( .A(n15381), .B(m[530]), .Z(n16424) );
  NAND U21042 ( .A(n15382), .B(creg[530]), .Z(n16423) );
  NAND U21043 ( .A(n16425), .B(n16426), .Z(y[52]) );
  NAND U21044 ( .A(n15381), .B(m[52]), .Z(n16426) );
  NAND U21045 ( .A(n15382), .B(creg[52]), .Z(n16425) );
  NAND U21046 ( .A(n16427), .B(n16428), .Z(y[529]) );
  NAND U21047 ( .A(n15381), .B(m[529]), .Z(n16428) );
  NAND U21048 ( .A(n15382), .B(creg[529]), .Z(n16427) );
  NAND U21049 ( .A(n16429), .B(n16430), .Z(y[528]) );
  NAND U21050 ( .A(n15381), .B(m[528]), .Z(n16430) );
  NAND U21051 ( .A(n15382), .B(creg[528]), .Z(n16429) );
  NAND U21052 ( .A(n16431), .B(n16432), .Z(y[527]) );
  NAND U21053 ( .A(n15381), .B(m[527]), .Z(n16432) );
  NAND U21054 ( .A(n15382), .B(creg[527]), .Z(n16431) );
  NAND U21055 ( .A(n16433), .B(n16434), .Z(y[526]) );
  NAND U21056 ( .A(n15381), .B(m[526]), .Z(n16434) );
  NAND U21057 ( .A(n15382), .B(creg[526]), .Z(n16433) );
  NAND U21058 ( .A(n16435), .B(n16436), .Z(y[525]) );
  NAND U21059 ( .A(n15381), .B(m[525]), .Z(n16436) );
  NAND U21060 ( .A(n15382), .B(creg[525]), .Z(n16435) );
  NAND U21061 ( .A(n16437), .B(n16438), .Z(y[524]) );
  NAND U21062 ( .A(n15381), .B(m[524]), .Z(n16438) );
  NAND U21063 ( .A(n15382), .B(creg[524]), .Z(n16437) );
  NAND U21064 ( .A(n16439), .B(n16440), .Z(y[523]) );
  NAND U21065 ( .A(n15381), .B(m[523]), .Z(n16440) );
  NAND U21066 ( .A(n15382), .B(creg[523]), .Z(n16439) );
  NAND U21067 ( .A(n16441), .B(n16442), .Z(y[522]) );
  NAND U21068 ( .A(n15381), .B(m[522]), .Z(n16442) );
  NAND U21069 ( .A(n15382), .B(creg[522]), .Z(n16441) );
  NAND U21070 ( .A(n16443), .B(n16444), .Z(y[521]) );
  NAND U21071 ( .A(n15381), .B(m[521]), .Z(n16444) );
  NAND U21072 ( .A(n15382), .B(creg[521]), .Z(n16443) );
  NAND U21073 ( .A(n16445), .B(n16446), .Z(y[520]) );
  NAND U21074 ( .A(n15381), .B(m[520]), .Z(n16446) );
  NAND U21075 ( .A(n15382), .B(creg[520]), .Z(n16445) );
  NAND U21076 ( .A(n16447), .B(n16448), .Z(y[51]) );
  NAND U21077 ( .A(n15381), .B(m[51]), .Z(n16448) );
  NAND U21078 ( .A(n15382), .B(creg[51]), .Z(n16447) );
  NAND U21079 ( .A(n16449), .B(n16450), .Z(y[519]) );
  NAND U21080 ( .A(n15381), .B(m[519]), .Z(n16450) );
  NAND U21081 ( .A(n15382), .B(creg[519]), .Z(n16449) );
  NAND U21082 ( .A(n16451), .B(n16452), .Z(y[518]) );
  NAND U21083 ( .A(n15381), .B(m[518]), .Z(n16452) );
  NAND U21084 ( .A(n15382), .B(creg[518]), .Z(n16451) );
  NAND U21085 ( .A(n16453), .B(n16454), .Z(y[517]) );
  NAND U21086 ( .A(n15381), .B(m[517]), .Z(n16454) );
  NAND U21087 ( .A(n15382), .B(creg[517]), .Z(n16453) );
  NAND U21088 ( .A(n16455), .B(n16456), .Z(y[516]) );
  NAND U21089 ( .A(n15381), .B(m[516]), .Z(n16456) );
  NAND U21090 ( .A(n15382), .B(creg[516]), .Z(n16455) );
  NAND U21091 ( .A(n16457), .B(n16458), .Z(y[515]) );
  NAND U21092 ( .A(n15381), .B(m[515]), .Z(n16458) );
  NAND U21093 ( .A(n15382), .B(creg[515]), .Z(n16457) );
  NAND U21094 ( .A(n16459), .B(n16460), .Z(y[514]) );
  NAND U21095 ( .A(n15381), .B(m[514]), .Z(n16460) );
  NAND U21096 ( .A(n15382), .B(creg[514]), .Z(n16459) );
  NAND U21097 ( .A(n16461), .B(n16462), .Z(y[513]) );
  NAND U21098 ( .A(n15381), .B(m[513]), .Z(n16462) );
  NAND U21099 ( .A(n15382), .B(creg[513]), .Z(n16461) );
  NAND U21100 ( .A(n16463), .B(n16464), .Z(y[512]) );
  NAND U21101 ( .A(n15381), .B(m[512]), .Z(n16464) );
  NAND U21102 ( .A(n15382), .B(creg[512]), .Z(n16463) );
  NAND U21103 ( .A(n16465), .B(n16466), .Z(y[511]) );
  NAND U21104 ( .A(n15381), .B(m[511]), .Z(n16466) );
  NAND U21105 ( .A(n15382), .B(creg[511]), .Z(n16465) );
  NAND U21106 ( .A(n16467), .B(n16468), .Z(y[510]) );
  NAND U21107 ( .A(n15381), .B(m[510]), .Z(n16468) );
  NAND U21108 ( .A(n15382), .B(creg[510]), .Z(n16467) );
  NAND U21109 ( .A(n16469), .B(n16470), .Z(y[50]) );
  NAND U21110 ( .A(n15381), .B(m[50]), .Z(n16470) );
  NAND U21111 ( .A(n15382), .B(creg[50]), .Z(n16469) );
  NAND U21112 ( .A(n16471), .B(n16472), .Z(y[509]) );
  NAND U21113 ( .A(n15381), .B(m[509]), .Z(n16472) );
  NAND U21114 ( .A(n15382), .B(creg[509]), .Z(n16471) );
  NAND U21115 ( .A(n16473), .B(n16474), .Z(y[508]) );
  NAND U21116 ( .A(n15381), .B(m[508]), .Z(n16474) );
  NAND U21117 ( .A(n15382), .B(creg[508]), .Z(n16473) );
  NAND U21118 ( .A(n16475), .B(n16476), .Z(y[507]) );
  NAND U21119 ( .A(n15381), .B(m[507]), .Z(n16476) );
  NAND U21120 ( .A(n15382), .B(creg[507]), .Z(n16475) );
  NAND U21121 ( .A(n16477), .B(n16478), .Z(y[506]) );
  NAND U21122 ( .A(n15381), .B(m[506]), .Z(n16478) );
  NAND U21123 ( .A(n15382), .B(creg[506]), .Z(n16477) );
  NAND U21124 ( .A(n16479), .B(n16480), .Z(y[505]) );
  NAND U21125 ( .A(n15381), .B(m[505]), .Z(n16480) );
  NAND U21126 ( .A(n15382), .B(creg[505]), .Z(n16479) );
  NAND U21127 ( .A(n16481), .B(n16482), .Z(y[504]) );
  NAND U21128 ( .A(n15381), .B(m[504]), .Z(n16482) );
  NAND U21129 ( .A(n15382), .B(creg[504]), .Z(n16481) );
  NAND U21130 ( .A(n16483), .B(n16484), .Z(y[503]) );
  NAND U21131 ( .A(n15381), .B(m[503]), .Z(n16484) );
  NAND U21132 ( .A(n15382), .B(creg[503]), .Z(n16483) );
  NAND U21133 ( .A(n16485), .B(n16486), .Z(y[502]) );
  NAND U21134 ( .A(n15381), .B(m[502]), .Z(n16486) );
  NAND U21135 ( .A(n15382), .B(creg[502]), .Z(n16485) );
  NAND U21136 ( .A(n16487), .B(n16488), .Z(y[501]) );
  NAND U21137 ( .A(n15381), .B(m[501]), .Z(n16488) );
  NAND U21138 ( .A(n15382), .B(creg[501]), .Z(n16487) );
  NAND U21139 ( .A(n16489), .B(n16490), .Z(y[500]) );
  NAND U21140 ( .A(n15381), .B(m[500]), .Z(n16490) );
  NAND U21141 ( .A(n15382), .B(creg[500]), .Z(n16489) );
  NAND U21142 ( .A(n16491), .B(n16492), .Z(y[4]) );
  NAND U21143 ( .A(n15381), .B(m[4]), .Z(n16492) );
  NAND U21144 ( .A(n15382), .B(creg[4]), .Z(n16491) );
  NAND U21145 ( .A(n16493), .B(n16494), .Z(y[49]) );
  NAND U21146 ( .A(n15381), .B(m[49]), .Z(n16494) );
  NAND U21147 ( .A(n15382), .B(creg[49]), .Z(n16493) );
  NAND U21148 ( .A(n16495), .B(n16496), .Z(y[499]) );
  NAND U21149 ( .A(n15381), .B(m[499]), .Z(n16496) );
  NAND U21150 ( .A(n15382), .B(creg[499]), .Z(n16495) );
  NAND U21151 ( .A(n16497), .B(n16498), .Z(y[498]) );
  NAND U21152 ( .A(n15381), .B(m[498]), .Z(n16498) );
  NAND U21153 ( .A(n15382), .B(creg[498]), .Z(n16497) );
  NAND U21154 ( .A(n16499), .B(n16500), .Z(y[497]) );
  NAND U21155 ( .A(n15381), .B(m[497]), .Z(n16500) );
  NAND U21156 ( .A(n15382), .B(creg[497]), .Z(n16499) );
  NAND U21157 ( .A(n16501), .B(n16502), .Z(y[496]) );
  NAND U21158 ( .A(n15381), .B(m[496]), .Z(n16502) );
  NAND U21159 ( .A(n15382), .B(creg[496]), .Z(n16501) );
  NAND U21160 ( .A(n16503), .B(n16504), .Z(y[495]) );
  NAND U21161 ( .A(n15381), .B(m[495]), .Z(n16504) );
  NAND U21162 ( .A(n15382), .B(creg[495]), .Z(n16503) );
  NAND U21163 ( .A(n16505), .B(n16506), .Z(y[494]) );
  NAND U21164 ( .A(n15381), .B(m[494]), .Z(n16506) );
  NAND U21165 ( .A(n15382), .B(creg[494]), .Z(n16505) );
  NAND U21166 ( .A(n16507), .B(n16508), .Z(y[493]) );
  NAND U21167 ( .A(n15381), .B(m[493]), .Z(n16508) );
  NAND U21168 ( .A(n15382), .B(creg[493]), .Z(n16507) );
  NAND U21169 ( .A(n16509), .B(n16510), .Z(y[492]) );
  NAND U21170 ( .A(n15381), .B(m[492]), .Z(n16510) );
  NAND U21171 ( .A(n15382), .B(creg[492]), .Z(n16509) );
  NAND U21172 ( .A(n16511), .B(n16512), .Z(y[491]) );
  NAND U21173 ( .A(n15381), .B(m[491]), .Z(n16512) );
  NAND U21174 ( .A(n15382), .B(creg[491]), .Z(n16511) );
  NAND U21175 ( .A(n16513), .B(n16514), .Z(y[490]) );
  NAND U21176 ( .A(n15381), .B(m[490]), .Z(n16514) );
  NAND U21177 ( .A(n15382), .B(creg[490]), .Z(n16513) );
  NAND U21178 ( .A(n16515), .B(n16516), .Z(y[48]) );
  NAND U21179 ( .A(n15381), .B(m[48]), .Z(n16516) );
  NAND U21180 ( .A(n15382), .B(creg[48]), .Z(n16515) );
  NAND U21181 ( .A(n16517), .B(n16518), .Z(y[489]) );
  NAND U21182 ( .A(n15381), .B(m[489]), .Z(n16518) );
  NAND U21183 ( .A(n15382), .B(creg[489]), .Z(n16517) );
  NAND U21184 ( .A(n16519), .B(n16520), .Z(y[488]) );
  NAND U21185 ( .A(n15381), .B(m[488]), .Z(n16520) );
  NAND U21186 ( .A(n15382), .B(creg[488]), .Z(n16519) );
  NAND U21187 ( .A(n16521), .B(n16522), .Z(y[487]) );
  NAND U21188 ( .A(n15381), .B(m[487]), .Z(n16522) );
  NAND U21189 ( .A(n15382), .B(creg[487]), .Z(n16521) );
  NAND U21190 ( .A(n16523), .B(n16524), .Z(y[486]) );
  NAND U21191 ( .A(n15381), .B(m[486]), .Z(n16524) );
  NAND U21192 ( .A(n15382), .B(creg[486]), .Z(n16523) );
  NAND U21193 ( .A(n16525), .B(n16526), .Z(y[485]) );
  NAND U21194 ( .A(n15381), .B(m[485]), .Z(n16526) );
  NAND U21195 ( .A(n15382), .B(creg[485]), .Z(n16525) );
  NAND U21196 ( .A(n16527), .B(n16528), .Z(y[484]) );
  NAND U21197 ( .A(n15381), .B(m[484]), .Z(n16528) );
  NAND U21198 ( .A(n15382), .B(creg[484]), .Z(n16527) );
  NAND U21199 ( .A(n16529), .B(n16530), .Z(y[483]) );
  NAND U21200 ( .A(n15381), .B(m[483]), .Z(n16530) );
  NAND U21201 ( .A(n15382), .B(creg[483]), .Z(n16529) );
  NAND U21202 ( .A(n16531), .B(n16532), .Z(y[482]) );
  NAND U21203 ( .A(n15381), .B(m[482]), .Z(n16532) );
  NAND U21204 ( .A(n15382), .B(creg[482]), .Z(n16531) );
  NAND U21205 ( .A(n16533), .B(n16534), .Z(y[481]) );
  NAND U21206 ( .A(n15381), .B(m[481]), .Z(n16534) );
  NAND U21207 ( .A(n15382), .B(creg[481]), .Z(n16533) );
  NAND U21208 ( .A(n16535), .B(n16536), .Z(y[480]) );
  NAND U21209 ( .A(n15381), .B(m[480]), .Z(n16536) );
  NAND U21210 ( .A(n15382), .B(creg[480]), .Z(n16535) );
  NAND U21211 ( .A(n16537), .B(n16538), .Z(y[47]) );
  NAND U21212 ( .A(n15381), .B(m[47]), .Z(n16538) );
  NAND U21213 ( .A(n15382), .B(creg[47]), .Z(n16537) );
  NAND U21214 ( .A(n16539), .B(n16540), .Z(y[479]) );
  NAND U21215 ( .A(n15381), .B(m[479]), .Z(n16540) );
  NAND U21216 ( .A(n15382), .B(creg[479]), .Z(n16539) );
  NAND U21217 ( .A(n16541), .B(n16542), .Z(y[478]) );
  NAND U21218 ( .A(n15381), .B(m[478]), .Z(n16542) );
  NAND U21219 ( .A(n15382), .B(creg[478]), .Z(n16541) );
  NAND U21220 ( .A(n16543), .B(n16544), .Z(y[477]) );
  NAND U21221 ( .A(n15381), .B(m[477]), .Z(n16544) );
  NAND U21222 ( .A(n15382), .B(creg[477]), .Z(n16543) );
  NAND U21223 ( .A(n16545), .B(n16546), .Z(y[476]) );
  NAND U21224 ( .A(n15381), .B(m[476]), .Z(n16546) );
  NAND U21225 ( .A(n15382), .B(creg[476]), .Z(n16545) );
  NAND U21226 ( .A(n16547), .B(n16548), .Z(y[475]) );
  NAND U21227 ( .A(n15381), .B(m[475]), .Z(n16548) );
  NAND U21228 ( .A(n15382), .B(creg[475]), .Z(n16547) );
  NAND U21229 ( .A(n16549), .B(n16550), .Z(y[474]) );
  NAND U21230 ( .A(n15381), .B(m[474]), .Z(n16550) );
  NAND U21231 ( .A(n15382), .B(creg[474]), .Z(n16549) );
  NAND U21232 ( .A(n16551), .B(n16552), .Z(y[473]) );
  NAND U21233 ( .A(n15381), .B(m[473]), .Z(n16552) );
  NAND U21234 ( .A(n15382), .B(creg[473]), .Z(n16551) );
  NAND U21235 ( .A(n16553), .B(n16554), .Z(y[472]) );
  NAND U21236 ( .A(n15381), .B(m[472]), .Z(n16554) );
  NAND U21237 ( .A(n15382), .B(creg[472]), .Z(n16553) );
  NAND U21238 ( .A(n16555), .B(n16556), .Z(y[471]) );
  NAND U21239 ( .A(n15381), .B(m[471]), .Z(n16556) );
  NAND U21240 ( .A(n15382), .B(creg[471]), .Z(n16555) );
  NAND U21241 ( .A(n16557), .B(n16558), .Z(y[470]) );
  NAND U21242 ( .A(n15381), .B(m[470]), .Z(n16558) );
  NAND U21243 ( .A(n15382), .B(creg[470]), .Z(n16557) );
  NAND U21244 ( .A(n16559), .B(n16560), .Z(y[46]) );
  NAND U21245 ( .A(n15381), .B(m[46]), .Z(n16560) );
  NAND U21246 ( .A(n15382), .B(creg[46]), .Z(n16559) );
  NAND U21247 ( .A(n16561), .B(n16562), .Z(y[469]) );
  NAND U21248 ( .A(n15381), .B(m[469]), .Z(n16562) );
  NAND U21249 ( .A(n15382), .B(creg[469]), .Z(n16561) );
  NAND U21250 ( .A(n16563), .B(n16564), .Z(y[468]) );
  NAND U21251 ( .A(n15381), .B(m[468]), .Z(n16564) );
  NAND U21252 ( .A(n15382), .B(creg[468]), .Z(n16563) );
  NAND U21253 ( .A(n16565), .B(n16566), .Z(y[467]) );
  NAND U21254 ( .A(n15381), .B(m[467]), .Z(n16566) );
  NAND U21255 ( .A(n15382), .B(creg[467]), .Z(n16565) );
  NAND U21256 ( .A(n16567), .B(n16568), .Z(y[466]) );
  NAND U21257 ( .A(n15381), .B(m[466]), .Z(n16568) );
  NAND U21258 ( .A(n15382), .B(creg[466]), .Z(n16567) );
  NAND U21259 ( .A(n16569), .B(n16570), .Z(y[465]) );
  NAND U21260 ( .A(n15381), .B(m[465]), .Z(n16570) );
  NAND U21261 ( .A(n15382), .B(creg[465]), .Z(n16569) );
  NAND U21262 ( .A(n16571), .B(n16572), .Z(y[464]) );
  NAND U21263 ( .A(n15381), .B(m[464]), .Z(n16572) );
  NAND U21264 ( .A(n15382), .B(creg[464]), .Z(n16571) );
  NAND U21265 ( .A(n16573), .B(n16574), .Z(y[463]) );
  NAND U21266 ( .A(n15381), .B(m[463]), .Z(n16574) );
  NAND U21267 ( .A(n15382), .B(creg[463]), .Z(n16573) );
  NAND U21268 ( .A(n16575), .B(n16576), .Z(y[462]) );
  NAND U21269 ( .A(n15381), .B(m[462]), .Z(n16576) );
  NAND U21270 ( .A(n15382), .B(creg[462]), .Z(n16575) );
  NAND U21271 ( .A(n16577), .B(n16578), .Z(y[461]) );
  NAND U21272 ( .A(n15381), .B(m[461]), .Z(n16578) );
  NAND U21273 ( .A(n15382), .B(creg[461]), .Z(n16577) );
  NAND U21274 ( .A(n16579), .B(n16580), .Z(y[460]) );
  NAND U21275 ( .A(n15381), .B(m[460]), .Z(n16580) );
  NAND U21276 ( .A(n15382), .B(creg[460]), .Z(n16579) );
  NAND U21277 ( .A(n16581), .B(n16582), .Z(y[45]) );
  NAND U21278 ( .A(n15381), .B(m[45]), .Z(n16582) );
  NAND U21279 ( .A(n15382), .B(creg[45]), .Z(n16581) );
  NAND U21280 ( .A(n16583), .B(n16584), .Z(y[459]) );
  NAND U21281 ( .A(n15381), .B(m[459]), .Z(n16584) );
  NAND U21282 ( .A(n15382), .B(creg[459]), .Z(n16583) );
  NAND U21283 ( .A(n16585), .B(n16586), .Z(y[458]) );
  NAND U21284 ( .A(n15381), .B(m[458]), .Z(n16586) );
  NAND U21285 ( .A(n15382), .B(creg[458]), .Z(n16585) );
  NAND U21286 ( .A(n16587), .B(n16588), .Z(y[457]) );
  NAND U21287 ( .A(n15381), .B(m[457]), .Z(n16588) );
  NAND U21288 ( .A(n15382), .B(creg[457]), .Z(n16587) );
  NAND U21289 ( .A(n16589), .B(n16590), .Z(y[456]) );
  NAND U21290 ( .A(n15381), .B(m[456]), .Z(n16590) );
  NAND U21291 ( .A(n15382), .B(creg[456]), .Z(n16589) );
  NAND U21292 ( .A(n16591), .B(n16592), .Z(y[455]) );
  NAND U21293 ( .A(n15381), .B(m[455]), .Z(n16592) );
  NAND U21294 ( .A(n15382), .B(creg[455]), .Z(n16591) );
  NAND U21295 ( .A(n16593), .B(n16594), .Z(y[454]) );
  NAND U21296 ( .A(n15381), .B(m[454]), .Z(n16594) );
  NAND U21297 ( .A(n15382), .B(creg[454]), .Z(n16593) );
  NAND U21298 ( .A(n16595), .B(n16596), .Z(y[453]) );
  NAND U21299 ( .A(n15381), .B(m[453]), .Z(n16596) );
  NAND U21300 ( .A(n15382), .B(creg[453]), .Z(n16595) );
  NAND U21301 ( .A(n16597), .B(n16598), .Z(y[452]) );
  NAND U21302 ( .A(n15381), .B(m[452]), .Z(n16598) );
  NAND U21303 ( .A(n15382), .B(creg[452]), .Z(n16597) );
  NAND U21304 ( .A(n16599), .B(n16600), .Z(y[451]) );
  NAND U21305 ( .A(n15381), .B(m[451]), .Z(n16600) );
  NAND U21306 ( .A(n15382), .B(creg[451]), .Z(n16599) );
  NAND U21307 ( .A(n16601), .B(n16602), .Z(y[450]) );
  NAND U21308 ( .A(n15381), .B(m[450]), .Z(n16602) );
  NAND U21309 ( .A(n15382), .B(creg[450]), .Z(n16601) );
  NAND U21310 ( .A(n16603), .B(n16604), .Z(y[44]) );
  NAND U21311 ( .A(n15381), .B(m[44]), .Z(n16604) );
  NAND U21312 ( .A(n15382), .B(creg[44]), .Z(n16603) );
  NAND U21313 ( .A(n16605), .B(n16606), .Z(y[449]) );
  NAND U21314 ( .A(n15381), .B(m[449]), .Z(n16606) );
  NAND U21315 ( .A(n15382), .B(creg[449]), .Z(n16605) );
  NAND U21316 ( .A(n16607), .B(n16608), .Z(y[448]) );
  NAND U21317 ( .A(n15381), .B(m[448]), .Z(n16608) );
  NAND U21318 ( .A(n15382), .B(creg[448]), .Z(n16607) );
  NAND U21319 ( .A(n16609), .B(n16610), .Z(y[447]) );
  NAND U21320 ( .A(n15381), .B(m[447]), .Z(n16610) );
  NAND U21321 ( .A(n15382), .B(creg[447]), .Z(n16609) );
  NAND U21322 ( .A(n16611), .B(n16612), .Z(y[446]) );
  NAND U21323 ( .A(n15381), .B(m[446]), .Z(n16612) );
  NAND U21324 ( .A(n15382), .B(creg[446]), .Z(n16611) );
  NAND U21325 ( .A(n16613), .B(n16614), .Z(y[445]) );
  NAND U21326 ( .A(n15381), .B(m[445]), .Z(n16614) );
  NAND U21327 ( .A(n15382), .B(creg[445]), .Z(n16613) );
  NAND U21328 ( .A(n16615), .B(n16616), .Z(y[444]) );
  NAND U21329 ( .A(n15381), .B(m[444]), .Z(n16616) );
  NAND U21330 ( .A(n15382), .B(creg[444]), .Z(n16615) );
  NAND U21331 ( .A(n16617), .B(n16618), .Z(y[443]) );
  NAND U21332 ( .A(n15381), .B(m[443]), .Z(n16618) );
  NAND U21333 ( .A(n15382), .B(creg[443]), .Z(n16617) );
  NAND U21334 ( .A(n16619), .B(n16620), .Z(y[442]) );
  NAND U21335 ( .A(n15381), .B(m[442]), .Z(n16620) );
  NAND U21336 ( .A(n15382), .B(creg[442]), .Z(n16619) );
  NAND U21337 ( .A(n16621), .B(n16622), .Z(y[441]) );
  NAND U21338 ( .A(n15381), .B(m[441]), .Z(n16622) );
  NAND U21339 ( .A(n15382), .B(creg[441]), .Z(n16621) );
  NAND U21340 ( .A(n16623), .B(n16624), .Z(y[440]) );
  NAND U21341 ( .A(n15381), .B(m[440]), .Z(n16624) );
  NAND U21342 ( .A(n15382), .B(creg[440]), .Z(n16623) );
  NAND U21343 ( .A(n16625), .B(n16626), .Z(y[43]) );
  NAND U21344 ( .A(n15381), .B(m[43]), .Z(n16626) );
  NAND U21345 ( .A(n15382), .B(creg[43]), .Z(n16625) );
  NAND U21346 ( .A(n16627), .B(n16628), .Z(y[439]) );
  NAND U21347 ( .A(n15381), .B(m[439]), .Z(n16628) );
  NAND U21348 ( .A(n15382), .B(creg[439]), .Z(n16627) );
  NAND U21349 ( .A(n16629), .B(n16630), .Z(y[438]) );
  NAND U21350 ( .A(n15381), .B(m[438]), .Z(n16630) );
  NAND U21351 ( .A(n15382), .B(creg[438]), .Z(n16629) );
  NAND U21352 ( .A(n16631), .B(n16632), .Z(y[437]) );
  NAND U21353 ( .A(n15381), .B(m[437]), .Z(n16632) );
  NAND U21354 ( .A(n15382), .B(creg[437]), .Z(n16631) );
  NAND U21355 ( .A(n16633), .B(n16634), .Z(y[436]) );
  NAND U21356 ( .A(n15381), .B(m[436]), .Z(n16634) );
  NAND U21357 ( .A(n15382), .B(creg[436]), .Z(n16633) );
  NAND U21358 ( .A(n16635), .B(n16636), .Z(y[435]) );
  NAND U21359 ( .A(n15381), .B(m[435]), .Z(n16636) );
  NAND U21360 ( .A(n15382), .B(creg[435]), .Z(n16635) );
  NAND U21361 ( .A(n16637), .B(n16638), .Z(y[434]) );
  NAND U21362 ( .A(n15381), .B(m[434]), .Z(n16638) );
  NAND U21363 ( .A(n15382), .B(creg[434]), .Z(n16637) );
  NAND U21364 ( .A(n16639), .B(n16640), .Z(y[433]) );
  NAND U21365 ( .A(n15381), .B(m[433]), .Z(n16640) );
  NAND U21366 ( .A(n15382), .B(creg[433]), .Z(n16639) );
  NAND U21367 ( .A(n16641), .B(n16642), .Z(y[432]) );
  NAND U21368 ( .A(n15381), .B(m[432]), .Z(n16642) );
  NAND U21369 ( .A(n15382), .B(creg[432]), .Z(n16641) );
  NAND U21370 ( .A(n16643), .B(n16644), .Z(y[431]) );
  NAND U21371 ( .A(n15381), .B(m[431]), .Z(n16644) );
  NAND U21372 ( .A(n15382), .B(creg[431]), .Z(n16643) );
  NAND U21373 ( .A(n16645), .B(n16646), .Z(y[430]) );
  NAND U21374 ( .A(n15381), .B(m[430]), .Z(n16646) );
  NAND U21375 ( .A(n15382), .B(creg[430]), .Z(n16645) );
  NAND U21376 ( .A(n16647), .B(n16648), .Z(y[42]) );
  NAND U21377 ( .A(n15381), .B(m[42]), .Z(n16648) );
  NAND U21378 ( .A(n15382), .B(creg[42]), .Z(n16647) );
  NAND U21379 ( .A(n16649), .B(n16650), .Z(y[429]) );
  NAND U21380 ( .A(n15381), .B(m[429]), .Z(n16650) );
  NAND U21381 ( .A(n15382), .B(creg[429]), .Z(n16649) );
  NAND U21382 ( .A(n16651), .B(n16652), .Z(y[428]) );
  NAND U21383 ( .A(n15381), .B(m[428]), .Z(n16652) );
  NAND U21384 ( .A(n15382), .B(creg[428]), .Z(n16651) );
  NAND U21385 ( .A(n16653), .B(n16654), .Z(y[427]) );
  NAND U21386 ( .A(n15381), .B(m[427]), .Z(n16654) );
  NAND U21387 ( .A(n15382), .B(creg[427]), .Z(n16653) );
  NAND U21388 ( .A(n16655), .B(n16656), .Z(y[426]) );
  NAND U21389 ( .A(n15381), .B(m[426]), .Z(n16656) );
  NAND U21390 ( .A(n15382), .B(creg[426]), .Z(n16655) );
  NAND U21391 ( .A(n16657), .B(n16658), .Z(y[425]) );
  NAND U21392 ( .A(n15381), .B(m[425]), .Z(n16658) );
  NAND U21393 ( .A(n15382), .B(creg[425]), .Z(n16657) );
  NAND U21394 ( .A(n16659), .B(n16660), .Z(y[424]) );
  NAND U21395 ( .A(n15381), .B(m[424]), .Z(n16660) );
  NAND U21396 ( .A(n15382), .B(creg[424]), .Z(n16659) );
  NAND U21397 ( .A(n16661), .B(n16662), .Z(y[423]) );
  NAND U21398 ( .A(n15381), .B(m[423]), .Z(n16662) );
  NAND U21399 ( .A(n15382), .B(creg[423]), .Z(n16661) );
  NAND U21400 ( .A(n16663), .B(n16664), .Z(y[422]) );
  NAND U21401 ( .A(n15381), .B(m[422]), .Z(n16664) );
  NAND U21402 ( .A(n15382), .B(creg[422]), .Z(n16663) );
  NAND U21403 ( .A(n16665), .B(n16666), .Z(y[421]) );
  NAND U21404 ( .A(n15381), .B(m[421]), .Z(n16666) );
  NAND U21405 ( .A(n15382), .B(creg[421]), .Z(n16665) );
  NAND U21406 ( .A(n16667), .B(n16668), .Z(y[420]) );
  NAND U21407 ( .A(n15381), .B(m[420]), .Z(n16668) );
  NAND U21408 ( .A(n15382), .B(creg[420]), .Z(n16667) );
  NAND U21409 ( .A(n16669), .B(n16670), .Z(y[41]) );
  NAND U21410 ( .A(n15381), .B(m[41]), .Z(n16670) );
  NAND U21411 ( .A(n15382), .B(creg[41]), .Z(n16669) );
  NAND U21412 ( .A(n16671), .B(n16672), .Z(y[419]) );
  NAND U21413 ( .A(n15381), .B(m[419]), .Z(n16672) );
  NAND U21414 ( .A(n15382), .B(creg[419]), .Z(n16671) );
  NAND U21415 ( .A(n16673), .B(n16674), .Z(y[418]) );
  NAND U21416 ( .A(n15381), .B(m[418]), .Z(n16674) );
  NAND U21417 ( .A(n15382), .B(creg[418]), .Z(n16673) );
  NAND U21418 ( .A(n16675), .B(n16676), .Z(y[417]) );
  NAND U21419 ( .A(n15381), .B(m[417]), .Z(n16676) );
  NAND U21420 ( .A(n15382), .B(creg[417]), .Z(n16675) );
  NAND U21421 ( .A(n16677), .B(n16678), .Z(y[416]) );
  NAND U21422 ( .A(n15381), .B(m[416]), .Z(n16678) );
  NAND U21423 ( .A(n15382), .B(creg[416]), .Z(n16677) );
  NAND U21424 ( .A(n16679), .B(n16680), .Z(y[415]) );
  NAND U21425 ( .A(n15381), .B(m[415]), .Z(n16680) );
  NAND U21426 ( .A(n15382), .B(creg[415]), .Z(n16679) );
  NAND U21427 ( .A(n16681), .B(n16682), .Z(y[414]) );
  NAND U21428 ( .A(n15381), .B(m[414]), .Z(n16682) );
  NAND U21429 ( .A(n15382), .B(creg[414]), .Z(n16681) );
  NAND U21430 ( .A(n16683), .B(n16684), .Z(y[413]) );
  NAND U21431 ( .A(n15381), .B(m[413]), .Z(n16684) );
  NAND U21432 ( .A(n15382), .B(creg[413]), .Z(n16683) );
  NAND U21433 ( .A(n16685), .B(n16686), .Z(y[412]) );
  NAND U21434 ( .A(n15381), .B(m[412]), .Z(n16686) );
  NAND U21435 ( .A(n15382), .B(creg[412]), .Z(n16685) );
  NAND U21436 ( .A(n16687), .B(n16688), .Z(y[411]) );
  NAND U21437 ( .A(n15381), .B(m[411]), .Z(n16688) );
  NAND U21438 ( .A(n15382), .B(creg[411]), .Z(n16687) );
  NAND U21439 ( .A(n16689), .B(n16690), .Z(y[410]) );
  NAND U21440 ( .A(n15381), .B(m[410]), .Z(n16690) );
  NAND U21441 ( .A(n15382), .B(creg[410]), .Z(n16689) );
  NAND U21442 ( .A(n16691), .B(n16692), .Z(y[40]) );
  NAND U21443 ( .A(n15381), .B(m[40]), .Z(n16692) );
  NAND U21444 ( .A(n15382), .B(creg[40]), .Z(n16691) );
  NAND U21445 ( .A(n16693), .B(n16694), .Z(y[409]) );
  NAND U21446 ( .A(n15381), .B(m[409]), .Z(n16694) );
  NAND U21447 ( .A(n15382), .B(creg[409]), .Z(n16693) );
  NAND U21448 ( .A(n16695), .B(n16696), .Z(y[408]) );
  NAND U21449 ( .A(n15381), .B(m[408]), .Z(n16696) );
  NAND U21450 ( .A(n15382), .B(creg[408]), .Z(n16695) );
  NAND U21451 ( .A(n16697), .B(n16698), .Z(y[407]) );
  NAND U21452 ( .A(n15381), .B(m[407]), .Z(n16698) );
  NAND U21453 ( .A(n15382), .B(creg[407]), .Z(n16697) );
  NAND U21454 ( .A(n16699), .B(n16700), .Z(y[406]) );
  NAND U21455 ( .A(n15381), .B(m[406]), .Z(n16700) );
  NAND U21456 ( .A(n15382), .B(creg[406]), .Z(n16699) );
  NAND U21457 ( .A(n16701), .B(n16702), .Z(y[405]) );
  NAND U21458 ( .A(n15381), .B(m[405]), .Z(n16702) );
  NAND U21459 ( .A(n15382), .B(creg[405]), .Z(n16701) );
  NAND U21460 ( .A(n16703), .B(n16704), .Z(y[404]) );
  NAND U21461 ( .A(n15381), .B(m[404]), .Z(n16704) );
  NAND U21462 ( .A(n15382), .B(creg[404]), .Z(n16703) );
  NAND U21463 ( .A(n16705), .B(n16706), .Z(y[403]) );
  NAND U21464 ( .A(n15381), .B(m[403]), .Z(n16706) );
  NAND U21465 ( .A(n15382), .B(creg[403]), .Z(n16705) );
  NAND U21466 ( .A(n16707), .B(n16708), .Z(y[402]) );
  NAND U21467 ( .A(n15381), .B(m[402]), .Z(n16708) );
  NAND U21468 ( .A(n15382), .B(creg[402]), .Z(n16707) );
  NAND U21469 ( .A(n16709), .B(n16710), .Z(y[401]) );
  NAND U21470 ( .A(n15381), .B(m[401]), .Z(n16710) );
  NAND U21471 ( .A(n15382), .B(creg[401]), .Z(n16709) );
  NAND U21472 ( .A(n16711), .B(n16712), .Z(y[400]) );
  NAND U21473 ( .A(n15381), .B(m[400]), .Z(n16712) );
  NAND U21474 ( .A(n15382), .B(creg[400]), .Z(n16711) );
  NAND U21475 ( .A(n16713), .B(n16714), .Z(y[3]) );
  NAND U21476 ( .A(n15381), .B(m[3]), .Z(n16714) );
  NAND U21477 ( .A(n15382), .B(creg[3]), .Z(n16713) );
  NAND U21478 ( .A(n16715), .B(n16716), .Z(y[39]) );
  NAND U21479 ( .A(n15381), .B(m[39]), .Z(n16716) );
  NAND U21480 ( .A(n15382), .B(creg[39]), .Z(n16715) );
  NAND U21481 ( .A(n16717), .B(n16718), .Z(y[399]) );
  NAND U21482 ( .A(n15381), .B(m[399]), .Z(n16718) );
  NAND U21483 ( .A(n15382), .B(creg[399]), .Z(n16717) );
  NAND U21484 ( .A(n16719), .B(n16720), .Z(y[398]) );
  NAND U21485 ( .A(n15381), .B(m[398]), .Z(n16720) );
  NAND U21486 ( .A(n15382), .B(creg[398]), .Z(n16719) );
  NAND U21487 ( .A(n16721), .B(n16722), .Z(y[397]) );
  NAND U21488 ( .A(n15381), .B(m[397]), .Z(n16722) );
  NAND U21489 ( .A(n15382), .B(creg[397]), .Z(n16721) );
  NAND U21490 ( .A(n16723), .B(n16724), .Z(y[396]) );
  NAND U21491 ( .A(n15381), .B(m[396]), .Z(n16724) );
  NAND U21492 ( .A(n15382), .B(creg[396]), .Z(n16723) );
  NAND U21493 ( .A(n16725), .B(n16726), .Z(y[395]) );
  NAND U21494 ( .A(n15381), .B(m[395]), .Z(n16726) );
  NAND U21495 ( .A(n15382), .B(creg[395]), .Z(n16725) );
  NAND U21496 ( .A(n16727), .B(n16728), .Z(y[394]) );
  NAND U21497 ( .A(n15381), .B(m[394]), .Z(n16728) );
  NAND U21498 ( .A(n15382), .B(creg[394]), .Z(n16727) );
  NAND U21499 ( .A(n16729), .B(n16730), .Z(y[393]) );
  NAND U21500 ( .A(n15381), .B(m[393]), .Z(n16730) );
  NAND U21501 ( .A(n15382), .B(creg[393]), .Z(n16729) );
  NAND U21502 ( .A(n16731), .B(n16732), .Z(y[392]) );
  NAND U21503 ( .A(n15381), .B(m[392]), .Z(n16732) );
  NAND U21504 ( .A(n15382), .B(creg[392]), .Z(n16731) );
  NAND U21505 ( .A(n16733), .B(n16734), .Z(y[391]) );
  NAND U21506 ( .A(n15381), .B(m[391]), .Z(n16734) );
  NAND U21507 ( .A(n15382), .B(creg[391]), .Z(n16733) );
  NAND U21508 ( .A(n16735), .B(n16736), .Z(y[390]) );
  NAND U21509 ( .A(n15381), .B(m[390]), .Z(n16736) );
  NAND U21510 ( .A(n15382), .B(creg[390]), .Z(n16735) );
  NAND U21511 ( .A(n16737), .B(n16738), .Z(y[38]) );
  NAND U21512 ( .A(n15381), .B(m[38]), .Z(n16738) );
  NAND U21513 ( .A(n15382), .B(creg[38]), .Z(n16737) );
  NAND U21514 ( .A(n16739), .B(n16740), .Z(y[389]) );
  NAND U21515 ( .A(n15381), .B(m[389]), .Z(n16740) );
  NAND U21516 ( .A(n15382), .B(creg[389]), .Z(n16739) );
  NAND U21517 ( .A(n16741), .B(n16742), .Z(y[388]) );
  NAND U21518 ( .A(n15381), .B(m[388]), .Z(n16742) );
  NAND U21519 ( .A(n15382), .B(creg[388]), .Z(n16741) );
  NAND U21520 ( .A(n16743), .B(n16744), .Z(y[387]) );
  NAND U21521 ( .A(n15381), .B(m[387]), .Z(n16744) );
  NAND U21522 ( .A(n15382), .B(creg[387]), .Z(n16743) );
  NAND U21523 ( .A(n16745), .B(n16746), .Z(y[386]) );
  NAND U21524 ( .A(n15381), .B(m[386]), .Z(n16746) );
  NAND U21525 ( .A(n15382), .B(creg[386]), .Z(n16745) );
  NAND U21526 ( .A(n16747), .B(n16748), .Z(y[385]) );
  NAND U21527 ( .A(n15381), .B(m[385]), .Z(n16748) );
  NAND U21528 ( .A(n15382), .B(creg[385]), .Z(n16747) );
  NAND U21529 ( .A(n16749), .B(n16750), .Z(y[384]) );
  NAND U21530 ( .A(n15381), .B(m[384]), .Z(n16750) );
  NAND U21531 ( .A(n15382), .B(creg[384]), .Z(n16749) );
  NAND U21532 ( .A(n16751), .B(n16752), .Z(y[383]) );
  NAND U21533 ( .A(n15381), .B(m[383]), .Z(n16752) );
  NAND U21534 ( .A(n15382), .B(creg[383]), .Z(n16751) );
  NAND U21535 ( .A(n16753), .B(n16754), .Z(y[382]) );
  NAND U21536 ( .A(n15381), .B(m[382]), .Z(n16754) );
  NAND U21537 ( .A(n15382), .B(creg[382]), .Z(n16753) );
  NAND U21538 ( .A(n16755), .B(n16756), .Z(y[381]) );
  NAND U21539 ( .A(n15381), .B(m[381]), .Z(n16756) );
  NAND U21540 ( .A(n15382), .B(creg[381]), .Z(n16755) );
  NAND U21541 ( .A(n16757), .B(n16758), .Z(y[380]) );
  NAND U21542 ( .A(n15381), .B(m[380]), .Z(n16758) );
  NAND U21543 ( .A(n15382), .B(creg[380]), .Z(n16757) );
  NAND U21544 ( .A(n16759), .B(n16760), .Z(y[37]) );
  NAND U21545 ( .A(n15381), .B(m[37]), .Z(n16760) );
  NAND U21546 ( .A(n15382), .B(creg[37]), .Z(n16759) );
  NAND U21547 ( .A(n16761), .B(n16762), .Z(y[379]) );
  NAND U21548 ( .A(n15381), .B(m[379]), .Z(n16762) );
  NAND U21549 ( .A(n15382), .B(creg[379]), .Z(n16761) );
  NAND U21550 ( .A(n16763), .B(n16764), .Z(y[378]) );
  NAND U21551 ( .A(n15381), .B(m[378]), .Z(n16764) );
  NAND U21552 ( .A(n15382), .B(creg[378]), .Z(n16763) );
  NAND U21553 ( .A(n16765), .B(n16766), .Z(y[377]) );
  NAND U21554 ( .A(n15381), .B(m[377]), .Z(n16766) );
  NAND U21555 ( .A(n15382), .B(creg[377]), .Z(n16765) );
  NAND U21556 ( .A(n16767), .B(n16768), .Z(y[376]) );
  NAND U21557 ( .A(n15381), .B(m[376]), .Z(n16768) );
  NAND U21558 ( .A(n15382), .B(creg[376]), .Z(n16767) );
  NAND U21559 ( .A(n16769), .B(n16770), .Z(y[375]) );
  NAND U21560 ( .A(n15381), .B(m[375]), .Z(n16770) );
  NAND U21561 ( .A(n15382), .B(creg[375]), .Z(n16769) );
  NAND U21562 ( .A(n16771), .B(n16772), .Z(y[374]) );
  NAND U21563 ( .A(n15381), .B(m[374]), .Z(n16772) );
  NAND U21564 ( .A(n15382), .B(creg[374]), .Z(n16771) );
  NAND U21565 ( .A(n16773), .B(n16774), .Z(y[373]) );
  NAND U21566 ( .A(n15381), .B(m[373]), .Z(n16774) );
  NAND U21567 ( .A(n15382), .B(creg[373]), .Z(n16773) );
  NAND U21568 ( .A(n16775), .B(n16776), .Z(y[372]) );
  NAND U21569 ( .A(n15381), .B(m[372]), .Z(n16776) );
  NAND U21570 ( .A(n15382), .B(creg[372]), .Z(n16775) );
  NAND U21571 ( .A(n16777), .B(n16778), .Z(y[371]) );
  NAND U21572 ( .A(n15381), .B(m[371]), .Z(n16778) );
  NAND U21573 ( .A(n15382), .B(creg[371]), .Z(n16777) );
  NAND U21574 ( .A(n16779), .B(n16780), .Z(y[370]) );
  NAND U21575 ( .A(n15381), .B(m[370]), .Z(n16780) );
  NAND U21576 ( .A(n15382), .B(creg[370]), .Z(n16779) );
  NAND U21577 ( .A(n16781), .B(n16782), .Z(y[36]) );
  NAND U21578 ( .A(n15381), .B(m[36]), .Z(n16782) );
  NAND U21579 ( .A(n15382), .B(creg[36]), .Z(n16781) );
  NAND U21580 ( .A(n16783), .B(n16784), .Z(y[369]) );
  NAND U21581 ( .A(n15381), .B(m[369]), .Z(n16784) );
  NAND U21582 ( .A(n15382), .B(creg[369]), .Z(n16783) );
  NAND U21583 ( .A(n16785), .B(n16786), .Z(y[368]) );
  NAND U21584 ( .A(n15381), .B(m[368]), .Z(n16786) );
  NAND U21585 ( .A(n15382), .B(creg[368]), .Z(n16785) );
  NAND U21586 ( .A(n16787), .B(n16788), .Z(y[367]) );
  NAND U21587 ( .A(n15381), .B(m[367]), .Z(n16788) );
  NAND U21588 ( .A(n15382), .B(creg[367]), .Z(n16787) );
  NAND U21589 ( .A(n16789), .B(n16790), .Z(y[366]) );
  NAND U21590 ( .A(n15381), .B(m[366]), .Z(n16790) );
  NAND U21591 ( .A(n15382), .B(creg[366]), .Z(n16789) );
  NAND U21592 ( .A(n16791), .B(n16792), .Z(y[365]) );
  NAND U21593 ( .A(n15381), .B(m[365]), .Z(n16792) );
  NAND U21594 ( .A(n15382), .B(creg[365]), .Z(n16791) );
  NAND U21595 ( .A(n16793), .B(n16794), .Z(y[364]) );
  NAND U21596 ( .A(n15381), .B(m[364]), .Z(n16794) );
  NAND U21597 ( .A(n15382), .B(creg[364]), .Z(n16793) );
  NAND U21598 ( .A(n16795), .B(n16796), .Z(y[363]) );
  NAND U21599 ( .A(n15381), .B(m[363]), .Z(n16796) );
  NAND U21600 ( .A(n15382), .B(creg[363]), .Z(n16795) );
  NAND U21601 ( .A(n16797), .B(n16798), .Z(y[362]) );
  NAND U21602 ( .A(n15381), .B(m[362]), .Z(n16798) );
  NAND U21603 ( .A(n15382), .B(creg[362]), .Z(n16797) );
  NAND U21604 ( .A(n16799), .B(n16800), .Z(y[361]) );
  NAND U21605 ( .A(n15381), .B(m[361]), .Z(n16800) );
  NAND U21606 ( .A(n15382), .B(creg[361]), .Z(n16799) );
  NAND U21607 ( .A(n16801), .B(n16802), .Z(y[360]) );
  NAND U21608 ( .A(n15381), .B(m[360]), .Z(n16802) );
  NAND U21609 ( .A(n15382), .B(creg[360]), .Z(n16801) );
  NAND U21610 ( .A(n16803), .B(n16804), .Z(y[35]) );
  NAND U21611 ( .A(n15381), .B(m[35]), .Z(n16804) );
  NAND U21612 ( .A(n15382), .B(creg[35]), .Z(n16803) );
  NAND U21613 ( .A(n16805), .B(n16806), .Z(y[359]) );
  NAND U21614 ( .A(n15381), .B(m[359]), .Z(n16806) );
  NAND U21615 ( .A(n15382), .B(creg[359]), .Z(n16805) );
  NAND U21616 ( .A(n16807), .B(n16808), .Z(y[358]) );
  NAND U21617 ( .A(n15381), .B(m[358]), .Z(n16808) );
  NAND U21618 ( .A(n15382), .B(creg[358]), .Z(n16807) );
  NAND U21619 ( .A(n16809), .B(n16810), .Z(y[357]) );
  NAND U21620 ( .A(n15381), .B(m[357]), .Z(n16810) );
  NAND U21621 ( .A(n15382), .B(creg[357]), .Z(n16809) );
  NAND U21622 ( .A(n16811), .B(n16812), .Z(y[356]) );
  NAND U21623 ( .A(n15381), .B(m[356]), .Z(n16812) );
  NAND U21624 ( .A(n15382), .B(creg[356]), .Z(n16811) );
  NAND U21625 ( .A(n16813), .B(n16814), .Z(y[355]) );
  NAND U21626 ( .A(n15381), .B(m[355]), .Z(n16814) );
  NAND U21627 ( .A(n15382), .B(creg[355]), .Z(n16813) );
  NAND U21628 ( .A(n16815), .B(n16816), .Z(y[354]) );
  NAND U21629 ( .A(n15381), .B(m[354]), .Z(n16816) );
  NAND U21630 ( .A(n15382), .B(creg[354]), .Z(n16815) );
  NAND U21631 ( .A(n16817), .B(n16818), .Z(y[353]) );
  NAND U21632 ( .A(n15381), .B(m[353]), .Z(n16818) );
  NAND U21633 ( .A(n15382), .B(creg[353]), .Z(n16817) );
  NAND U21634 ( .A(n16819), .B(n16820), .Z(y[352]) );
  NAND U21635 ( .A(n15381), .B(m[352]), .Z(n16820) );
  NAND U21636 ( .A(n15382), .B(creg[352]), .Z(n16819) );
  NAND U21637 ( .A(n16821), .B(n16822), .Z(y[351]) );
  NAND U21638 ( .A(n15381), .B(m[351]), .Z(n16822) );
  NAND U21639 ( .A(n15382), .B(creg[351]), .Z(n16821) );
  NAND U21640 ( .A(n16823), .B(n16824), .Z(y[350]) );
  NAND U21641 ( .A(n15381), .B(m[350]), .Z(n16824) );
  NAND U21642 ( .A(n15382), .B(creg[350]), .Z(n16823) );
  NAND U21643 ( .A(n16825), .B(n16826), .Z(y[34]) );
  NAND U21644 ( .A(n15381), .B(m[34]), .Z(n16826) );
  NAND U21645 ( .A(n15382), .B(creg[34]), .Z(n16825) );
  NAND U21646 ( .A(n16827), .B(n16828), .Z(y[349]) );
  NAND U21647 ( .A(n15381), .B(m[349]), .Z(n16828) );
  NAND U21648 ( .A(n15382), .B(creg[349]), .Z(n16827) );
  NAND U21649 ( .A(n16829), .B(n16830), .Z(y[348]) );
  NAND U21650 ( .A(n15381), .B(m[348]), .Z(n16830) );
  NAND U21651 ( .A(n15382), .B(creg[348]), .Z(n16829) );
  NAND U21652 ( .A(n16831), .B(n16832), .Z(y[347]) );
  NAND U21653 ( .A(n15381), .B(m[347]), .Z(n16832) );
  NAND U21654 ( .A(n15382), .B(creg[347]), .Z(n16831) );
  NAND U21655 ( .A(n16833), .B(n16834), .Z(y[346]) );
  NAND U21656 ( .A(n15381), .B(m[346]), .Z(n16834) );
  NAND U21657 ( .A(n15382), .B(creg[346]), .Z(n16833) );
  NAND U21658 ( .A(n16835), .B(n16836), .Z(y[345]) );
  NAND U21659 ( .A(n15381), .B(m[345]), .Z(n16836) );
  NAND U21660 ( .A(n15382), .B(creg[345]), .Z(n16835) );
  NAND U21661 ( .A(n16837), .B(n16838), .Z(y[344]) );
  NAND U21662 ( .A(n15381), .B(m[344]), .Z(n16838) );
  NAND U21663 ( .A(n15382), .B(creg[344]), .Z(n16837) );
  NAND U21664 ( .A(n16839), .B(n16840), .Z(y[343]) );
  NAND U21665 ( .A(n15381), .B(m[343]), .Z(n16840) );
  NAND U21666 ( .A(n15382), .B(creg[343]), .Z(n16839) );
  NAND U21667 ( .A(n16841), .B(n16842), .Z(y[342]) );
  NAND U21668 ( .A(n15381), .B(m[342]), .Z(n16842) );
  NAND U21669 ( .A(n15382), .B(creg[342]), .Z(n16841) );
  NAND U21670 ( .A(n16843), .B(n16844), .Z(y[341]) );
  NAND U21671 ( .A(n15381), .B(m[341]), .Z(n16844) );
  NAND U21672 ( .A(n15382), .B(creg[341]), .Z(n16843) );
  NAND U21673 ( .A(n16845), .B(n16846), .Z(y[340]) );
  NAND U21674 ( .A(n15381), .B(m[340]), .Z(n16846) );
  NAND U21675 ( .A(n15382), .B(creg[340]), .Z(n16845) );
  NAND U21676 ( .A(n16847), .B(n16848), .Z(y[33]) );
  NAND U21677 ( .A(n15381), .B(m[33]), .Z(n16848) );
  NAND U21678 ( .A(n15382), .B(creg[33]), .Z(n16847) );
  NAND U21679 ( .A(n16849), .B(n16850), .Z(y[339]) );
  NAND U21680 ( .A(n15381), .B(m[339]), .Z(n16850) );
  NAND U21681 ( .A(n15382), .B(creg[339]), .Z(n16849) );
  NAND U21682 ( .A(n16851), .B(n16852), .Z(y[338]) );
  NAND U21683 ( .A(n15381), .B(m[338]), .Z(n16852) );
  NAND U21684 ( .A(n15382), .B(creg[338]), .Z(n16851) );
  NAND U21685 ( .A(n16853), .B(n16854), .Z(y[337]) );
  NAND U21686 ( .A(n15381), .B(m[337]), .Z(n16854) );
  NAND U21687 ( .A(n15382), .B(creg[337]), .Z(n16853) );
  NAND U21688 ( .A(n16855), .B(n16856), .Z(y[336]) );
  NAND U21689 ( .A(n15381), .B(m[336]), .Z(n16856) );
  NAND U21690 ( .A(n15382), .B(creg[336]), .Z(n16855) );
  NAND U21691 ( .A(n16857), .B(n16858), .Z(y[335]) );
  NAND U21692 ( .A(n15381), .B(m[335]), .Z(n16858) );
  NAND U21693 ( .A(n15382), .B(creg[335]), .Z(n16857) );
  NAND U21694 ( .A(n16859), .B(n16860), .Z(y[334]) );
  NAND U21695 ( .A(n15381), .B(m[334]), .Z(n16860) );
  NAND U21696 ( .A(n15382), .B(creg[334]), .Z(n16859) );
  NAND U21697 ( .A(n16861), .B(n16862), .Z(y[333]) );
  NAND U21698 ( .A(n15381), .B(m[333]), .Z(n16862) );
  NAND U21699 ( .A(n15382), .B(creg[333]), .Z(n16861) );
  NAND U21700 ( .A(n16863), .B(n16864), .Z(y[332]) );
  NAND U21701 ( .A(n15381), .B(m[332]), .Z(n16864) );
  NAND U21702 ( .A(n15382), .B(creg[332]), .Z(n16863) );
  NAND U21703 ( .A(n16865), .B(n16866), .Z(y[331]) );
  NAND U21704 ( .A(n15381), .B(m[331]), .Z(n16866) );
  NAND U21705 ( .A(n15382), .B(creg[331]), .Z(n16865) );
  NAND U21706 ( .A(n16867), .B(n16868), .Z(y[330]) );
  NAND U21707 ( .A(n15381), .B(m[330]), .Z(n16868) );
  NAND U21708 ( .A(n15382), .B(creg[330]), .Z(n16867) );
  NAND U21709 ( .A(n16869), .B(n16870), .Z(y[32]) );
  NAND U21710 ( .A(n15381), .B(m[32]), .Z(n16870) );
  NAND U21711 ( .A(n15382), .B(creg[32]), .Z(n16869) );
  NAND U21712 ( .A(n16871), .B(n16872), .Z(y[329]) );
  NAND U21713 ( .A(n15381), .B(m[329]), .Z(n16872) );
  NAND U21714 ( .A(n15382), .B(creg[329]), .Z(n16871) );
  NAND U21715 ( .A(n16873), .B(n16874), .Z(y[328]) );
  NAND U21716 ( .A(n15381), .B(m[328]), .Z(n16874) );
  NAND U21717 ( .A(n15382), .B(creg[328]), .Z(n16873) );
  NAND U21718 ( .A(n16875), .B(n16876), .Z(y[327]) );
  NAND U21719 ( .A(n15381), .B(m[327]), .Z(n16876) );
  NAND U21720 ( .A(n15382), .B(creg[327]), .Z(n16875) );
  NAND U21721 ( .A(n16877), .B(n16878), .Z(y[326]) );
  NAND U21722 ( .A(n15381), .B(m[326]), .Z(n16878) );
  NAND U21723 ( .A(n15382), .B(creg[326]), .Z(n16877) );
  NAND U21724 ( .A(n16879), .B(n16880), .Z(y[325]) );
  NAND U21725 ( .A(n15381), .B(m[325]), .Z(n16880) );
  NAND U21726 ( .A(n15382), .B(creg[325]), .Z(n16879) );
  NAND U21727 ( .A(n16881), .B(n16882), .Z(y[324]) );
  NAND U21728 ( .A(n15381), .B(m[324]), .Z(n16882) );
  NAND U21729 ( .A(n15382), .B(creg[324]), .Z(n16881) );
  NAND U21730 ( .A(n16883), .B(n16884), .Z(y[323]) );
  NAND U21731 ( .A(n15381), .B(m[323]), .Z(n16884) );
  NAND U21732 ( .A(n15382), .B(creg[323]), .Z(n16883) );
  NAND U21733 ( .A(n16885), .B(n16886), .Z(y[322]) );
  NAND U21734 ( .A(n15381), .B(m[322]), .Z(n16886) );
  NAND U21735 ( .A(n15382), .B(creg[322]), .Z(n16885) );
  NAND U21736 ( .A(n16887), .B(n16888), .Z(y[321]) );
  NAND U21737 ( .A(n15381), .B(m[321]), .Z(n16888) );
  NAND U21738 ( .A(n15382), .B(creg[321]), .Z(n16887) );
  NAND U21739 ( .A(n16889), .B(n16890), .Z(y[320]) );
  NAND U21740 ( .A(n15381), .B(m[320]), .Z(n16890) );
  NAND U21741 ( .A(n15382), .B(creg[320]), .Z(n16889) );
  NAND U21742 ( .A(n16891), .B(n16892), .Z(y[31]) );
  NAND U21743 ( .A(n15381), .B(m[31]), .Z(n16892) );
  NAND U21744 ( .A(n15382), .B(creg[31]), .Z(n16891) );
  NAND U21745 ( .A(n16893), .B(n16894), .Z(y[319]) );
  NAND U21746 ( .A(n15381), .B(m[319]), .Z(n16894) );
  NAND U21747 ( .A(n15382), .B(creg[319]), .Z(n16893) );
  NAND U21748 ( .A(n16895), .B(n16896), .Z(y[318]) );
  NAND U21749 ( .A(n15381), .B(m[318]), .Z(n16896) );
  NAND U21750 ( .A(n15382), .B(creg[318]), .Z(n16895) );
  NAND U21751 ( .A(n16897), .B(n16898), .Z(y[317]) );
  NAND U21752 ( .A(n15381), .B(m[317]), .Z(n16898) );
  NAND U21753 ( .A(n15382), .B(creg[317]), .Z(n16897) );
  NAND U21754 ( .A(n16899), .B(n16900), .Z(y[316]) );
  NAND U21755 ( .A(n15381), .B(m[316]), .Z(n16900) );
  NAND U21756 ( .A(n15382), .B(creg[316]), .Z(n16899) );
  NAND U21757 ( .A(n16901), .B(n16902), .Z(y[315]) );
  NAND U21758 ( .A(n15381), .B(m[315]), .Z(n16902) );
  NAND U21759 ( .A(n15382), .B(creg[315]), .Z(n16901) );
  NAND U21760 ( .A(n16903), .B(n16904), .Z(y[314]) );
  NAND U21761 ( .A(n15381), .B(m[314]), .Z(n16904) );
  NAND U21762 ( .A(n15382), .B(creg[314]), .Z(n16903) );
  NAND U21763 ( .A(n16905), .B(n16906), .Z(y[313]) );
  NAND U21764 ( .A(n15381), .B(m[313]), .Z(n16906) );
  NAND U21765 ( .A(n15382), .B(creg[313]), .Z(n16905) );
  NAND U21766 ( .A(n16907), .B(n16908), .Z(y[312]) );
  NAND U21767 ( .A(n15381), .B(m[312]), .Z(n16908) );
  NAND U21768 ( .A(n15382), .B(creg[312]), .Z(n16907) );
  NAND U21769 ( .A(n16909), .B(n16910), .Z(y[311]) );
  NAND U21770 ( .A(n15381), .B(m[311]), .Z(n16910) );
  NAND U21771 ( .A(n15382), .B(creg[311]), .Z(n16909) );
  NAND U21772 ( .A(n16911), .B(n16912), .Z(y[310]) );
  NAND U21773 ( .A(n15381), .B(m[310]), .Z(n16912) );
  NAND U21774 ( .A(n15382), .B(creg[310]), .Z(n16911) );
  NAND U21775 ( .A(n16913), .B(n16914), .Z(y[30]) );
  NAND U21776 ( .A(n15381), .B(m[30]), .Z(n16914) );
  NAND U21777 ( .A(n15382), .B(creg[30]), .Z(n16913) );
  NAND U21778 ( .A(n16915), .B(n16916), .Z(y[309]) );
  NAND U21779 ( .A(n15381), .B(m[309]), .Z(n16916) );
  NAND U21780 ( .A(n15382), .B(creg[309]), .Z(n16915) );
  NAND U21781 ( .A(n16917), .B(n16918), .Z(y[308]) );
  NAND U21782 ( .A(n15381), .B(m[308]), .Z(n16918) );
  NAND U21783 ( .A(n15382), .B(creg[308]), .Z(n16917) );
  NAND U21784 ( .A(n16919), .B(n16920), .Z(y[307]) );
  NAND U21785 ( .A(n15381), .B(m[307]), .Z(n16920) );
  NAND U21786 ( .A(n15382), .B(creg[307]), .Z(n16919) );
  NAND U21787 ( .A(n16921), .B(n16922), .Z(y[306]) );
  NAND U21788 ( .A(n15381), .B(m[306]), .Z(n16922) );
  NAND U21789 ( .A(n15382), .B(creg[306]), .Z(n16921) );
  NAND U21790 ( .A(n16923), .B(n16924), .Z(y[305]) );
  NAND U21791 ( .A(n15381), .B(m[305]), .Z(n16924) );
  NAND U21792 ( .A(n15382), .B(creg[305]), .Z(n16923) );
  NAND U21793 ( .A(n16925), .B(n16926), .Z(y[304]) );
  NAND U21794 ( .A(n15381), .B(m[304]), .Z(n16926) );
  NAND U21795 ( .A(n15382), .B(creg[304]), .Z(n16925) );
  NAND U21796 ( .A(n16927), .B(n16928), .Z(y[303]) );
  NAND U21797 ( .A(n15381), .B(m[303]), .Z(n16928) );
  NAND U21798 ( .A(n15382), .B(creg[303]), .Z(n16927) );
  NAND U21799 ( .A(n16929), .B(n16930), .Z(y[302]) );
  NAND U21800 ( .A(n15381), .B(m[302]), .Z(n16930) );
  NAND U21801 ( .A(n15382), .B(creg[302]), .Z(n16929) );
  NAND U21802 ( .A(n16931), .B(n16932), .Z(y[301]) );
  NAND U21803 ( .A(n15381), .B(m[301]), .Z(n16932) );
  NAND U21804 ( .A(n15382), .B(creg[301]), .Z(n16931) );
  NAND U21805 ( .A(n16933), .B(n16934), .Z(y[300]) );
  NAND U21806 ( .A(n15381), .B(m[300]), .Z(n16934) );
  NAND U21807 ( .A(n15382), .B(creg[300]), .Z(n16933) );
  NAND U21808 ( .A(n16935), .B(n16936), .Z(y[2]) );
  NAND U21809 ( .A(n15381), .B(m[2]), .Z(n16936) );
  NAND U21810 ( .A(n15382), .B(creg[2]), .Z(n16935) );
  NAND U21811 ( .A(n16937), .B(n16938), .Z(y[29]) );
  NAND U21812 ( .A(n15381), .B(m[29]), .Z(n16938) );
  NAND U21813 ( .A(n15382), .B(creg[29]), .Z(n16937) );
  NAND U21814 ( .A(n16939), .B(n16940), .Z(y[299]) );
  NAND U21815 ( .A(n15381), .B(m[299]), .Z(n16940) );
  NAND U21816 ( .A(n15382), .B(creg[299]), .Z(n16939) );
  NAND U21817 ( .A(n16941), .B(n16942), .Z(y[298]) );
  NAND U21818 ( .A(n15381), .B(m[298]), .Z(n16942) );
  NAND U21819 ( .A(n15382), .B(creg[298]), .Z(n16941) );
  NAND U21820 ( .A(n16943), .B(n16944), .Z(y[297]) );
  NAND U21821 ( .A(n15381), .B(m[297]), .Z(n16944) );
  NAND U21822 ( .A(n15382), .B(creg[297]), .Z(n16943) );
  NAND U21823 ( .A(n16945), .B(n16946), .Z(y[296]) );
  NAND U21824 ( .A(n15381), .B(m[296]), .Z(n16946) );
  NAND U21825 ( .A(n15382), .B(creg[296]), .Z(n16945) );
  NAND U21826 ( .A(n16947), .B(n16948), .Z(y[295]) );
  NAND U21827 ( .A(n15381), .B(m[295]), .Z(n16948) );
  NAND U21828 ( .A(n15382), .B(creg[295]), .Z(n16947) );
  NAND U21829 ( .A(n16949), .B(n16950), .Z(y[294]) );
  NAND U21830 ( .A(n15381), .B(m[294]), .Z(n16950) );
  NAND U21831 ( .A(n15382), .B(creg[294]), .Z(n16949) );
  NAND U21832 ( .A(n16951), .B(n16952), .Z(y[293]) );
  NAND U21833 ( .A(n15381), .B(m[293]), .Z(n16952) );
  NAND U21834 ( .A(n15382), .B(creg[293]), .Z(n16951) );
  NAND U21835 ( .A(n16953), .B(n16954), .Z(y[292]) );
  NAND U21836 ( .A(n15381), .B(m[292]), .Z(n16954) );
  NAND U21837 ( .A(n15382), .B(creg[292]), .Z(n16953) );
  NAND U21838 ( .A(n16955), .B(n16956), .Z(y[291]) );
  NAND U21839 ( .A(n15381), .B(m[291]), .Z(n16956) );
  NAND U21840 ( .A(n15382), .B(creg[291]), .Z(n16955) );
  NAND U21841 ( .A(n16957), .B(n16958), .Z(y[290]) );
  NAND U21842 ( .A(n15381), .B(m[290]), .Z(n16958) );
  NAND U21843 ( .A(n15382), .B(creg[290]), .Z(n16957) );
  NAND U21844 ( .A(n16959), .B(n16960), .Z(y[28]) );
  NAND U21845 ( .A(n15381), .B(m[28]), .Z(n16960) );
  NAND U21846 ( .A(n15382), .B(creg[28]), .Z(n16959) );
  NAND U21847 ( .A(n16961), .B(n16962), .Z(y[289]) );
  NAND U21848 ( .A(n15381), .B(m[289]), .Z(n16962) );
  NAND U21849 ( .A(n15382), .B(creg[289]), .Z(n16961) );
  NAND U21850 ( .A(n16963), .B(n16964), .Z(y[288]) );
  NAND U21851 ( .A(n15381), .B(m[288]), .Z(n16964) );
  NAND U21852 ( .A(n15382), .B(creg[288]), .Z(n16963) );
  NAND U21853 ( .A(n16965), .B(n16966), .Z(y[287]) );
  NAND U21854 ( .A(n15381), .B(m[287]), .Z(n16966) );
  NAND U21855 ( .A(n15382), .B(creg[287]), .Z(n16965) );
  NAND U21856 ( .A(n16967), .B(n16968), .Z(y[286]) );
  NAND U21857 ( .A(n15381), .B(m[286]), .Z(n16968) );
  NAND U21858 ( .A(n15382), .B(creg[286]), .Z(n16967) );
  NAND U21859 ( .A(n16969), .B(n16970), .Z(y[285]) );
  NAND U21860 ( .A(n15381), .B(m[285]), .Z(n16970) );
  NAND U21861 ( .A(n15382), .B(creg[285]), .Z(n16969) );
  NAND U21862 ( .A(n16971), .B(n16972), .Z(y[284]) );
  NAND U21863 ( .A(n15381), .B(m[284]), .Z(n16972) );
  NAND U21864 ( .A(n15382), .B(creg[284]), .Z(n16971) );
  NAND U21865 ( .A(n16973), .B(n16974), .Z(y[283]) );
  NAND U21866 ( .A(n15381), .B(m[283]), .Z(n16974) );
  NAND U21867 ( .A(n15382), .B(creg[283]), .Z(n16973) );
  NAND U21868 ( .A(n16975), .B(n16976), .Z(y[282]) );
  NAND U21869 ( .A(n15381), .B(m[282]), .Z(n16976) );
  NAND U21870 ( .A(n15382), .B(creg[282]), .Z(n16975) );
  NAND U21871 ( .A(n16977), .B(n16978), .Z(y[281]) );
  NAND U21872 ( .A(n15381), .B(m[281]), .Z(n16978) );
  NAND U21873 ( .A(n15382), .B(creg[281]), .Z(n16977) );
  NAND U21874 ( .A(n16979), .B(n16980), .Z(y[280]) );
  NAND U21875 ( .A(n15381), .B(m[280]), .Z(n16980) );
  NAND U21876 ( .A(n15382), .B(creg[280]), .Z(n16979) );
  NAND U21877 ( .A(n16981), .B(n16982), .Z(y[27]) );
  NAND U21878 ( .A(n15381), .B(m[27]), .Z(n16982) );
  NAND U21879 ( .A(n15382), .B(creg[27]), .Z(n16981) );
  NAND U21880 ( .A(n16983), .B(n16984), .Z(y[279]) );
  NAND U21881 ( .A(n15381), .B(m[279]), .Z(n16984) );
  NAND U21882 ( .A(n15382), .B(creg[279]), .Z(n16983) );
  NAND U21883 ( .A(n16985), .B(n16986), .Z(y[278]) );
  NAND U21884 ( .A(n15381), .B(m[278]), .Z(n16986) );
  NAND U21885 ( .A(n15382), .B(creg[278]), .Z(n16985) );
  NAND U21886 ( .A(n16987), .B(n16988), .Z(y[277]) );
  NAND U21887 ( .A(n15381), .B(m[277]), .Z(n16988) );
  NAND U21888 ( .A(n15382), .B(creg[277]), .Z(n16987) );
  NAND U21889 ( .A(n16989), .B(n16990), .Z(y[276]) );
  NAND U21890 ( .A(n15381), .B(m[276]), .Z(n16990) );
  NAND U21891 ( .A(n15382), .B(creg[276]), .Z(n16989) );
  NAND U21892 ( .A(n16991), .B(n16992), .Z(y[275]) );
  NAND U21893 ( .A(n15381), .B(m[275]), .Z(n16992) );
  NAND U21894 ( .A(n15382), .B(creg[275]), .Z(n16991) );
  NAND U21895 ( .A(n16993), .B(n16994), .Z(y[274]) );
  NAND U21896 ( .A(n15381), .B(m[274]), .Z(n16994) );
  NAND U21897 ( .A(n15382), .B(creg[274]), .Z(n16993) );
  NAND U21898 ( .A(n16995), .B(n16996), .Z(y[273]) );
  NAND U21899 ( .A(n15381), .B(m[273]), .Z(n16996) );
  NAND U21900 ( .A(n15382), .B(creg[273]), .Z(n16995) );
  NAND U21901 ( .A(n16997), .B(n16998), .Z(y[272]) );
  NAND U21902 ( .A(n15381), .B(m[272]), .Z(n16998) );
  NAND U21903 ( .A(n15382), .B(creg[272]), .Z(n16997) );
  NAND U21904 ( .A(n16999), .B(n17000), .Z(y[271]) );
  NAND U21905 ( .A(n15381), .B(m[271]), .Z(n17000) );
  NAND U21906 ( .A(n15382), .B(creg[271]), .Z(n16999) );
  NAND U21907 ( .A(n17001), .B(n17002), .Z(y[270]) );
  NAND U21908 ( .A(n15381), .B(m[270]), .Z(n17002) );
  NAND U21909 ( .A(n15382), .B(creg[270]), .Z(n17001) );
  NAND U21910 ( .A(n17003), .B(n17004), .Z(y[26]) );
  NAND U21911 ( .A(n15381), .B(m[26]), .Z(n17004) );
  NAND U21912 ( .A(n15382), .B(creg[26]), .Z(n17003) );
  NAND U21913 ( .A(n17005), .B(n17006), .Z(y[269]) );
  NAND U21914 ( .A(n15381), .B(m[269]), .Z(n17006) );
  NAND U21915 ( .A(n15382), .B(creg[269]), .Z(n17005) );
  NAND U21916 ( .A(n17007), .B(n17008), .Z(y[268]) );
  NAND U21917 ( .A(n15381), .B(m[268]), .Z(n17008) );
  NAND U21918 ( .A(n15382), .B(creg[268]), .Z(n17007) );
  NAND U21919 ( .A(n17009), .B(n17010), .Z(y[267]) );
  NAND U21920 ( .A(n15381), .B(m[267]), .Z(n17010) );
  NAND U21921 ( .A(n15382), .B(creg[267]), .Z(n17009) );
  NAND U21922 ( .A(n17011), .B(n17012), .Z(y[266]) );
  NAND U21923 ( .A(n15381), .B(m[266]), .Z(n17012) );
  NAND U21924 ( .A(n15382), .B(creg[266]), .Z(n17011) );
  NAND U21925 ( .A(n17013), .B(n17014), .Z(y[265]) );
  NAND U21926 ( .A(n15381), .B(m[265]), .Z(n17014) );
  NAND U21927 ( .A(n15382), .B(creg[265]), .Z(n17013) );
  NAND U21928 ( .A(n17015), .B(n17016), .Z(y[264]) );
  NAND U21929 ( .A(n15381), .B(m[264]), .Z(n17016) );
  NAND U21930 ( .A(n15382), .B(creg[264]), .Z(n17015) );
  NAND U21931 ( .A(n17017), .B(n17018), .Z(y[263]) );
  NAND U21932 ( .A(n15381), .B(m[263]), .Z(n17018) );
  NAND U21933 ( .A(n15382), .B(creg[263]), .Z(n17017) );
  NAND U21934 ( .A(n17019), .B(n17020), .Z(y[262]) );
  NAND U21935 ( .A(n15381), .B(m[262]), .Z(n17020) );
  NAND U21936 ( .A(n15382), .B(creg[262]), .Z(n17019) );
  NAND U21937 ( .A(n17021), .B(n17022), .Z(y[261]) );
  NAND U21938 ( .A(n15381), .B(m[261]), .Z(n17022) );
  NAND U21939 ( .A(n15382), .B(creg[261]), .Z(n17021) );
  NAND U21940 ( .A(n17023), .B(n17024), .Z(y[260]) );
  NAND U21941 ( .A(n15381), .B(m[260]), .Z(n17024) );
  NAND U21942 ( .A(n15382), .B(creg[260]), .Z(n17023) );
  NAND U21943 ( .A(n17025), .B(n17026), .Z(y[25]) );
  NAND U21944 ( .A(n15381), .B(m[25]), .Z(n17026) );
  NAND U21945 ( .A(n15382), .B(creg[25]), .Z(n17025) );
  NAND U21946 ( .A(n17027), .B(n17028), .Z(y[259]) );
  NAND U21947 ( .A(n15381), .B(m[259]), .Z(n17028) );
  NAND U21948 ( .A(n15382), .B(creg[259]), .Z(n17027) );
  NAND U21949 ( .A(n17029), .B(n17030), .Z(y[258]) );
  NAND U21950 ( .A(n15381), .B(m[258]), .Z(n17030) );
  NAND U21951 ( .A(n15382), .B(creg[258]), .Z(n17029) );
  NAND U21952 ( .A(n17031), .B(n17032), .Z(y[257]) );
  NAND U21953 ( .A(n15381), .B(m[257]), .Z(n17032) );
  NAND U21954 ( .A(n15382), .B(creg[257]), .Z(n17031) );
  NAND U21955 ( .A(n17033), .B(n17034), .Z(y[256]) );
  NAND U21956 ( .A(n15381), .B(m[256]), .Z(n17034) );
  NAND U21957 ( .A(n15382), .B(creg[256]), .Z(n17033) );
  NAND U21958 ( .A(n17035), .B(n17036), .Z(y[255]) );
  NAND U21959 ( .A(n15381), .B(m[255]), .Z(n17036) );
  NAND U21960 ( .A(n15382), .B(creg[255]), .Z(n17035) );
  NAND U21961 ( .A(n17037), .B(n17038), .Z(y[254]) );
  NAND U21962 ( .A(n15381), .B(m[254]), .Z(n17038) );
  NAND U21963 ( .A(n15382), .B(creg[254]), .Z(n17037) );
  NAND U21964 ( .A(n17039), .B(n17040), .Z(y[253]) );
  NAND U21965 ( .A(n15381), .B(m[253]), .Z(n17040) );
  NAND U21966 ( .A(n15382), .B(creg[253]), .Z(n17039) );
  NAND U21967 ( .A(n17041), .B(n17042), .Z(y[252]) );
  NAND U21968 ( .A(n15381), .B(m[252]), .Z(n17042) );
  NAND U21969 ( .A(n15382), .B(creg[252]), .Z(n17041) );
  NAND U21970 ( .A(n17043), .B(n17044), .Z(y[251]) );
  NAND U21971 ( .A(n15381), .B(m[251]), .Z(n17044) );
  NAND U21972 ( .A(n15382), .B(creg[251]), .Z(n17043) );
  NAND U21973 ( .A(n17045), .B(n17046), .Z(y[250]) );
  NAND U21974 ( .A(n15381), .B(m[250]), .Z(n17046) );
  NAND U21975 ( .A(n15382), .B(creg[250]), .Z(n17045) );
  NAND U21976 ( .A(n17047), .B(n17048), .Z(y[24]) );
  NAND U21977 ( .A(n15381), .B(m[24]), .Z(n17048) );
  NAND U21978 ( .A(n15382), .B(creg[24]), .Z(n17047) );
  NAND U21979 ( .A(n17049), .B(n17050), .Z(y[249]) );
  NAND U21980 ( .A(n15381), .B(m[249]), .Z(n17050) );
  NAND U21981 ( .A(n15382), .B(creg[249]), .Z(n17049) );
  NAND U21982 ( .A(n17051), .B(n17052), .Z(y[248]) );
  NAND U21983 ( .A(n15381), .B(m[248]), .Z(n17052) );
  NAND U21984 ( .A(n15382), .B(creg[248]), .Z(n17051) );
  NAND U21985 ( .A(n17053), .B(n17054), .Z(y[247]) );
  NAND U21986 ( .A(n15381), .B(m[247]), .Z(n17054) );
  NAND U21987 ( .A(n15382), .B(creg[247]), .Z(n17053) );
  NAND U21988 ( .A(n17055), .B(n17056), .Z(y[246]) );
  NAND U21989 ( .A(n15381), .B(m[246]), .Z(n17056) );
  NAND U21990 ( .A(n15382), .B(creg[246]), .Z(n17055) );
  NAND U21991 ( .A(n17057), .B(n17058), .Z(y[245]) );
  NAND U21992 ( .A(n15381), .B(m[245]), .Z(n17058) );
  NAND U21993 ( .A(n15382), .B(creg[245]), .Z(n17057) );
  NAND U21994 ( .A(n17059), .B(n17060), .Z(y[244]) );
  NAND U21995 ( .A(n15381), .B(m[244]), .Z(n17060) );
  NAND U21996 ( .A(n15382), .B(creg[244]), .Z(n17059) );
  NAND U21997 ( .A(n17061), .B(n17062), .Z(y[243]) );
  NAND U21998 ( .A(n15381), .B(m[243]), .Z(n17062) );
  NAND U21999 ( .A(n15382), .B(creg[243]), .Z(n17061) );
  NAND U22000 ( .A(n17063), .B(n17064), .Z(y[242]) );
  NAND U22001 ( .A(n15381), .B(m[242]), .Z(n17064) );
  NAND U22002 ( .A(n15382), .B(creg[242]), .Z(n17063) );
  NAND U22003 ( .A(n17065), .B(n17066), .Z(y[241]) );
  NAND U22004 ( .A(n15381), .B(m[241]), .Z(n17066) );
  NAND U22005 ( .A(n15382), .B(creg[241]), .Z(n17065) );
  NAND U22006 ( .A(n17067), .B(n17068), .Z(y[240]) );
  NAND U22007 ( .A(n15381), .B(m[240]), .Z(n17068) );
  NAND U22008 ( .A(n15382), .B(creg[240]), .Z(n17067) );
  NAND U22009 ( .A(n17069), .B(n17070), .Z(y[23]) );
  NAND U22010 ( .A(n15381), .B(m[23]), .Z(n17070) );
  NAND U22011 ( .A(n15382), .B(creg[23]), .Z(n17069) );
  NAND U22012 ( .A(n17071), .B(n17072), .Z(y[239]) );
  NAND U22013 ( .A(n15381), .B(m[239]), .Z(n17072) );
  NAND U22014 ( .A(n15382), .B(creg[239]), .Z(n17071) );
  NAND U22015 ( .A(n17073), .B(n17074), .Z(y[238]) );
  NAND U22016 ( .A(n15381), .B(m[238]), .Z(n17074) );
  NAND U22017 ( .A(n15382), .B(creg[238]), .Z(n17073) );
  NAND U22018 ( .A(n17075), .B(n17076), .Z(y[237]) );
  NAND U22019 ( .A(n15381), .B(m[237]), .Z(n17076) );
  NAND U22020 ( .A(n15382), .B(creg[237]), .Z(n17075) );
  NAND U22021 ( .A(n17077), .B(n17078), .Z(y[236]) );
  NAND U22022 ( .A(n15381), .B(m[236]), .Z(n17078) );
  NAND U22023 ( .A(n15382), .B(creg[236]), .Z(n17077) );
  NAND U22024 ( .A(n17079), .B(n17080), .Z(y[235]) );
  NAND U22025 ( .A(n15381), .B(m[235]), .Z(n17080) );
  NAND U22026 ( .A(n15382), .B(creg[235]), .Z(n17079) );
  NAND U22027 ( .A(n17081), .B(n17082), .Z(y[234]) );
  NAND U22028 ( .A(n15381), .B(m[234]), .Z(n17082) );
  NAND U22029 ( .A(n15382), .B(creg[234]), .Z(n17081) );
  NAND U22030 ( .A(n17083), .B(n17084), .Z(y[233]) );
  NAND U22031 ( .A(n15381), .B(m[233]), .Z(n17084) );
  NAND U22032 ( .A(n15382), .B(creg[233]), .Z(n17083) );
  NAND U22033 ( .A(n17085), .B(n17086), .Z(y[232]) );
  NAND U22034 ( .A(n15381), .B(m[232]), .Z(n17086) );
  NAND U22035 ( .A(n15382), .B(creg[232]), .Z(n17085) );
  NAND U22036 ( .A(n17087), .B(n17088), .Z(y[231]) );
  NAND U22037 ( .A(n15381), .B(m[231]), .Z(n17088) );
  NAND U22038 ( .A(n15382), .B(creg[231]), .Z(n17087) );
  NAND U22039 ( .A(n17089), .B(n17090), .Z(y[230]) );
  NAND U22040 ( .A(n15381), .B(m[230]), .Z(n17090) );
  NAND U22041 ( .A(n15382), .B(creg[230]), .Z(n17089) );
  NAND U22042 ( .A(n17091), .B(n17092), .Z(y[22]) );
  NAND U22043 ( .A(n15381), .B(m[22]), .Z(n17092) );
  NAND U22044 ( .A(n15382), .B(creg[22]), .Z(n17091) );
  NAND U22045 ( .A(n17093), .B(n17094), .Z(y[229]) );
  NAND U22046 ( .A(n15381), .B(m[229]), .Z(n17094) );
  NAND U22047 ( .A(n15382), .B(creg[229]), .Z(n17093) );
  NAND U22048 ( .A(n17095), .B(n17096), .Z(y[228]) );
  NAND U22049 ( .A(n15381), .B(m[228]), .Z(n17096) );
  NAND U22050 ( .A(n15382), .B(creg[228]), .Z(n17095) );
  NAND U22051 ( .A(n17097), .B(n17098), .Z(y[227]) );
  NAND U22052 ( .A(n15381), .B(m[227]), .Z(n17098) );
  NAND U22053 ( .A(n15382), .B(creg[227]), .Z(n17097) );
  NAND U22054 ( .A(n17099), .B(n17100), .Z(y[226]) );
  NAND U22055 ( .A(n15381), .B(m[226]), .Z(n17100) );
  NAND U22056 ( .A(n15382), .B(creg[226]), .Z(n17099) );
  NAND U22057 ( .A(n17101), .B(n17102), .Z(y[225]) );
  NAND U22058 ( .A(n15381), .B(m[225]), .Z(n17102) );
  NAND U22059 ( .A(n15382), .B(creg[225]), .Z(n17101) );
  NAND U22060 ( .A(n17103), .B(n17104), .Z(y[224]) );
  NAND U22061 ( .A(n15381), .B(m[224]), .Z(n17104) );
  NAND U22062 ( .A(n15382), .B(creg[224]), .Z(n17103) );
  NAND U22063 ( .A(n17105), .B(n17106), .Z(y[223]) );
  NAND U22064 ( .A(n15381), .B(m[223]), .Z(n17106) );
  NAND U22065 ( .A(n15382), .B(creg[223]), .Z(n17105) );
  NAND U22066 ( .A(n17107), .B(n17108), .Z(y[222]) );
  NAND U22067 ( .A(n15381), .B(m[222]), .Z(n17108) );
  NAND U22068 ( .A(n15382), .B(creg[222]), .Z(n17107) );
  NAND U22069 ( .A(n17109), .B(n17110), .Z(y[221]) );
  NAND U22070 ( .A(n15381), .B(m[221]), .Z(n17110) );
  NAND U22071 ( .A(n15382), .B(creg[221]), .Z(n17109) );
  NAND U22072 ( .A(n17111), .B(n17112), .Z(y[220]) );
  NAND U22073 ( .A(n15381), .B(m[220]), .Z(n17112) );
  NAND U22074 ( .A(n15382), .B(creg[220]), .Z(n17111) );
  NAND U22075 ( .A(n17113), .B(n17114), .Z(y[21]) );
  NAND U22076 ( .A(n15381), .B(m[21]), .Z(n17114) );
  NAND U22077 ( .A(n15382), .B(creg[21]), .Z(n17113) );
  NAND U22078 ( .A(n17115), .B(n17116), .Z(y[219]) );
  NAND U22079 ( .A(n15381), .B(m[219]), .Z(n17116) );
  NAND U22080 ( .A(n15382), .B(creg[219]), .Z(n17115) );
  NAND U22081 ( .A(n17117), .B(n17118), .Z(y[218]) );
  NAND U22082 ( .A(n15381), .B(m[218]), .Z(n17118) );
  NAND U22083 ( .A(n15382), .B(creg[218]), .Z(n17117) );
  NAND U22084 ( .A(n17119), .B(n17120), .Z(y[217]) );
  NAND U22085 ( .A(n15381), .B(m[217]), .Z(n17120) );
  NAND U22086 ( .A(n15382), .B(creg[217]), .Z(n17119) );
  NAND U22087 ( .A(n17121), .B(n17122), .Z(y[216]) );
  NAND U22088 ( .A(n15381), .B(m[216]), .Z(n17122) );
  NAND U22089 ( .A(n15382), .B(creg[216]), .Z(n17121) );
  NAND U22090 ( .A(n17123), .B(n17124), .Z(y[215]) );
  NAND U22091 ( .A(n15381), .B(m[215]), .Z(n17124) );
  NAND U22092 ( .A(n15382), .B(creg[215]), .Z(n17123) );
  NAND U22093 ( .A(n17125), .B(n17126), .Z(y[214]) );
  NAND U22094 ( .A(n15381), .B(m[214]), .Z(n17126) );
  NAND U22095 ( .A(n15382), .B(creg[214]), .Z(n17125) );
  NAND U22096 ( .A(n17127), .B(n17128), .Z(y[213]) );
  NAND U22097 ( .A(n15381), .B(m[213]), .Z(n17128) );
  NAND U22098 ( .A(n15382), .B(creg[213]), .Z(n17127) );
  NAND U22099 ( .A(n17129), .B(n17130), .Z(y[212]) );
  NAND U22100 ( .A(n15381), .B(m[212]), .Z(n17130) );
  NAND U22101 ( .A(n15382), .B(creg[212]), .Z(n17129) );
  NAND U22102 ( .A(n17131), .B(n17132), .Z(y[211]) );
  NAND U22103 ( .A(n15381), .B(m[211]), .Z(n17132) );
  NAND U22104 ( .A(n15382), .B(creg[211]), .Z(n17131) );
  NAND U22105 ( .A(n17133), .B(n17134), .Z(y[210]) );
  NAND U22106 ( .A(n15381), .B(m[210]), .Z(n17134) );
  NAND U22107 ( .A(n15382), .B(creg[210]), .Z(n17133) );
  NAND U22108 ( .A(n17135), .B(n17136), .Z(y[20]) );
  NAND U22109 ( .A(n15381), .B(m[20]), .Z(n17136) );
  NAND U22110 ( .A(n15382), .B(creg[20]), .Z(n17135) );
  NAND U22111 ( .A(n17137), .B(n17138), .Z(y[209]) );
  NAND U22112 ( .A(n15381), .B(m[209]), .Z(n17138) );
  NAND U22113 ( .A(n15382), .B(creg[209]), .Z(n17137) );
  NAND U22114 ( .A(n17139), .B(n17140), .Z(y[208]) );
  NAND U22115 ( .A(n15381), .B(m[208]), .Z(n17140) );
  NAND U22116 ( .A(n15382), .B(creg[208]), .Z(n17139) );
  NAND U22117 ( .A(n17141), .B(n17142), .Z(y[207]) );
  NAND U22118 ( .A(n15381), .B(m[207]), .Z(n17142) );
  NAND U22119 ( .A(n15382), .B(creg[207]), .Z(n17141) );
  NAND U22120 ( .A(n17143), .B(n17144), .Z(y[206]) );
  NAND U22121 ( .A(n15381), .B(m[206]), .Z(n17144) );
  NAND U22122 ( .A(n15382), .B(creg[206]), .Z(n17143) );
  NAND U22123 ( .A(n17145), .B(n17146), .Z(y[205]) );
  NAND U22124 ( .A(n15381), .B(m[205]), .Z(n17146) );
  NAND U22125 ( .A(n15382), .B(creg[205]), .Z(n17145) );
  NAND U22126 ( .A(n17147), .B(n17148), .Z(y[204]) );
  NAND U22127 ( .A(n15381), .B(m[204]), .Z(n17148) );
  NAND U22128 ( .A(n15382), .B(creg[204]), .Z(n17147) );
  NAND U22129 ( .A(n17149), .B(n17150), .Z(y[203]) );
  NAND U22130 ( .A(n15381), .B(m[203]), .Z(n17150) );
  NAND U22131 ( .A(n15382), .B(creg[203]), .Z(n17149) );
  NAND U22132 ( .A(n17151), .B(n17152), .Z(y[202]) );
  NAND U22133 ( .A(n15381), .B(m[202]), .Z(n17152) );
  NAND U22134 ( .A(n15382), .B(creg[202]), .Z(n17151) );
  NAND U22135 ( .A(n17153), .B(n17154), .Z(y[201]) );
  NAND U22136 ( .A(n15381), .B(m[201]), .Z(n17154) );
  NAND U22137 ( .A(n15382), .B(creg[201]), .Z(n17153) );
  NAND U22138 ( .A(n17155), .B(n17156), .Z(y[200]) );
  NAND U22139 ( .A(n15381), .B(m[200]), .Z(n17156) );
  NAND U22140 ( .A(n15382), .B(creg[200]), .Z(n17155) );
  NAND U22141 ( .A(n17157), .B(n17158), .Z(y[1]) );
  NAND U22142 ( .A(n15381), .B(m[1]), .Z(n17158) );
  NAND U22143 ( .A(n15382), .B(creg[1]), .Z(n17157) );
  NAND U22144 ( .A(n17159), .B(n17160), .Z(y[19]) );
  NAND U22145 ( .A(n15381), .B(m[19]), .Z(n17160) );
  NAND U22146 ( .A(n15382), .B(creg[19]), .Z(n17159) );
  NAND U22147 ( .A(n17161), .B(n17162), .Z(y[199]) );
  NAND U22148 ( .A(n15381), .B(m[199]), .Z(n17162) );
  NAND U22149 ( .A(n15382), .B(creg[199]), .Z(n17161) );
  NAND U22150 ( .A(n17163), .B(n17164), .Z(y[198]) );
  NAND U22151 ( .A(n15381), .B(m[198]), .Z(n17164) );
  NAND U22152 ( .A(n15382), .B(creg[198]), .Z(n17163) );
  NAND U22153 ( .A(n17165), .B(n17166), .Z(y[197]) );
  NAND U22154 ( .A(n15381), .B(m[197]), .Z(n17166) );
  NAND U22155 ( .A(n15382), .B(creg[197]), .Z(n17165) );
  NAND U22156 ( .A(n17167), .B(n17168), .Z(y[196]) );
  NAND U22157 ( .A(n15381), .B(m[196]), .Z(n17168) );
  NAND U22158 ( .A(n15382), .B(creg[196]), .Z(n17167) );
  NAND U22159 ( .A(n17169), .B(n17170), .Z(y[195]) );
  NAND U22160 ( .A(n15381), .B(m[195]), .Z(n17170) );
  NAND U22161 ( .A(n15382), .B(creg[195]), .Z(n17169) );
  NAND U22162 ( .A(n17171), .B(n17172), .Z(y[194]) );
  NAND U22163 ( .A(n15381), .B(m[194]), .Z(n17172) );
  NAND U22164 ( .A(n15382), .B(creg[194]), .Z(n17171) );
  NAND U22165 ( .A(n17173), .B(n17174), .Z(y[193]) );
  NAND U22166 ( .A(n15381), .B(m[193]), .Z(n17174) );
  NAND U22167 ( .A(n15382), .B(creg[193]), .Z(n17173) );
  NAND U22168 ( .A(n17175), .B(n17176), .Z(y[192]) );
  NAND U22169 ( .A(n15381), .B(m[192]), .Z(n17176) );
  NAND U22170 ( .A(n15382), .B(creg[192]), .Z(n17175) );
  NAND U22171 ( .A(n17177), .B(n17178), .Z(y[191]) );
  NAND U22172 ( .A(n15381), .B(m[191]), .Z(n17178) );
  NAND U22173 ( .A(n15382), .B(creg[191]), .Z(n17177) );
  NAND U22174 ( .A(n17179), .B(n17180), .Z(y[190]) );
  NAND U22175 ( .A(n15381), .B(m[190]), .Z(n17180) );
  NAND U22176 ( .A(n15382), .B(creg[190]), .Z(n17179) );
  NAND U22177 ( .A(n17181), .B(n17182), .Z(y[18]) );
  NAND U22178 ( .A(n15381), .B(m[18]), .Z(n17182) );
  NAND U22179 ( .A(n15382), .B(creg[18]), .Z(n17181) );
  NAND U22180 ( .A(n17183), .B(n17184), .Z(y[189]) );
  NAND U22181 ( .A(n15381), .B(m[189]), .Z(n17184) );
  NAND U22182 ( .A(n15382), .B(creg[189]), .Z(n17183) );
  NAND U22183 ( .A(n17185), .B(n17186), .Z(y[188]) );
  NAND U22184 ( .A(n15381), .B(m[188]), .Z(n17186) );
  NAND U22185 ( .A(n15382), .B(creg[188]), .Z(n17185) );
  NAND U22186 ( .A(n17187), .B(n17188), .Z(y[187]) );
  NAND U22187 ( .A(n15381), .B(m[187]), .Z(n17188) );
  NAND U22188 ( .A(n15382), .B(creg[187]), .Z(n17187) );
  NAND U22189 ( .A(n17189), .B(n17190), .Z(y[186]) );
  NAND U22190 ( .A(n15381), .B(m[186]), .Z(n17190) );
  NAND U22191 ( .A(n15382), .B(creg[186]), .Z(n17189) );
  NAND U22192 ( .A(n17191), .B(n17192), .Z(y[185]) );
  NAND U22193 ( .A(n15381), .B(m[185]), .Z(n17192) );
  NAND U22194 ( .A(n15382), .B(creg[185]), .Z(n17191) );
  NAND U22195 ( .A(n17193), .B(n17194), .Z(y[184]) );
  NAND U22196 ( .A(n15381), .B(m[184]), .Z(n17194) );
  NAND U22197 ( .A(n15382), .B(creg[184]), .Z(n17193) );
  NAND U22198 ( .A(n17195), .B(n17196), .Z(y[183]) );
  NAND U22199 ( .A(n15381), .B(m[183]), .Z(n17196) );
  NAND U22200 ( .A(n15382), .B(creg[183]), .Z(n17195) );
  NAND U22201 ( .A(n17197), .B(n17198), .Z(y[182]) );
  NAND U22202 ( .A(n15381), .B(m[182]), .Z(n17198) );
  NAND U22203 ( .A(n15382), .B(creg[182]), .Z(n17197) );
  NAND U22204 ( .A(n17199), .B(n17200), .Z(y[181]) );
  NAND U22205 ( .A(n15381), .B(m[181]), .Z(n17200) );
  NAND U22206 ( .A(n15382), .B(creg[181]), .Z(n17199) );
  NAND U22207 ( .A(n17201), .B(n17202), .Z(y[180]) );
  NAND U22208 ( .A(n15381), .B(m[180]), .Z(n17202) );
  NAND U22209 ( .A(n15382), .B(creg[180]), .Z(n17201) );
  NAND U22210 ( .A(n17203), .B(n17204), .Z(y[17]) );
  NAND U22211 ( .A(n15381), .B(m[17]), .Z(n17204) );
  NAND U22212 ( .A(n15382), .B(creg[17]), .Z(n17203) );
  NAND U22213 ( .A(n17205), .B(n17206), .Z(y[179]) );
  NAND U22214 ( .A(n15381), .B(m[179]), .Z(n17206) );
  NAND U22215 ( .A(n15382), .B(creg[179]), .Z(n17205) );
  NAND U22216 ( .A(n17207), .B(n17208), .Z(y[178]) );
  NAND U22217 ( .A(n15381), .B(m[178]), .Z(n17208) );
  NAND U22218 ( .A(n15382), .B(creg[178]), .Z(n17207) );
  NAND U22219 ( .A(n17209), .B(n17210), .Z(y[177]) );
  NAND U22220 ( .A(n15381), .B(m[177]), .Z(n17210) );
  NAND U22221 ( .A(n15382), .B(creg[177]), .Z(n17209) );
  NAND U22222 ( .A(n17211), .B(n17212), .Z(y[176]) );
  NAND U22223 ( .A(n15381), .B(m[176]), .Z(n17212) );
  NAND U22224 ( .A(n15382), .B(creg[176]), .Z(n17211) );
  NAND U22225 ( .A(n17213), .B(n17214), .Z(y[175]) );
  NAND U22226 ( .A(n15381), .B(m[175]), .Z(n17214) );
  NAND U22227 ( .A(n15382), .B(creg[175]), .Z(n17213) );
  NAND U22228 ( .A(n17215), .B(n17216), .Z(y[174]) );
  NAND U22229 ( .A(n15381), .B(m[174]), .Z(n17216) );
  NAND U22230 ( .A(n15382), .B(creg[174]), .Z(n17215) );
  NAND U22231 ( .A(n17217), .B(n17218), .Z(y[173]) );
  NAND U22232 ( .A(n15381), .B(m[173]), .Z(n17218) );
  NAND U22233 ( .A(n15382), .B(creg[173]), .Z(n17217) );
  NAND U22234 ( .A(n17219), .B(n17220), .Z(y[172]) );
  NAND U22235 ( .A(n15381), .B(m[172]), .Z(n17220) );
  NAND U22236 ( .A(n15382), .B(creg[172]), .Z(n17219) );
  NAND U22237 ( .A(n17221), .B(n17222), .Z(y[171]) );
  NAND U22238 ( .A(n15381), .B(m[171]), .Z(n17222) );
  NAND U22239 ( .A(n15382), .B(creg[171]), .Z(n17221) );
  NAND U22240 ( .A(n17223), .B(n17224), .Z(y[170]) );
  NAND U22241 ( .A(n15381), .B(m[170]), .Z(n17224) );
  NAND U22242 ( .A(n15382), .B(creg[170]), .Z(n17223) );
  NAND U22243 ( .A(n17225), .B(n17226), .Z(y[16]) );
  NAND U22244 ( .A(n15381), .B(m[16]), .Z(n17226) );
  NAND U22245 ( .A(n15382), .B(creg[16]), .Z(n17225) );
  NAND U22246 ( .A(n17227), .B(n17228), .Z(y[169]) );
  NAND U22247 ( .A(n15381), .B(m[169]), .Z(n17228) );
  NAND U22248 ( .A(n15382), .B(creg[169]), .Z(n17227) );
  NAND U22249 ( .A(n17229), .B(n17230), .Z(y[168]) );
  NAND U22250 ( .A(n15381), .B(m[168]), .Z(n17230) );
  NAND U22251 ( .A(n15382), .B(creg[168]), .Z(n17229) );
  NAND U22252 ( .A(n17231), .B(n17232), .Z(y[167]) );
  NAND U22253 ( .A(n15381), .B(m[167]), .Z(n17232) );
  NAND U22254 ( .A(n15382), .B(creg[167]), .Z(n17231) );
  NAND U22255 ( .A(n17233), .B(n17234), .Z(y[166]) );
  NAND U22256 ( .A(n15381), .B(m[166]), .Z(n17234) );
  NAND U22257 ( .A(n15382), .B(creg[166]), .Z(n17233) );
  NAND U22258 ( .A(n17235), .B(n17236), .Z(y[165]) );
  NAND U22259 ( .A(n15381), .B(m[165]), .Z(n17236) );
  NAND U22260 ( .A(n15382), .B(creg[165]), .Z(n17235) );
  NAND U22261 ( .A(n17237), .B(n17238), .Z(y[164]) );
  NAND U22262 ( .A(n15381), .B(m[164]), .Z(n17238) );
  NAND U22263 ( .A(n15382), .B(creg[164]), .Z(n17237) );
  NAND U22264 ( .A(n17239), .B(n17240), .Z(y[163]) );
  NAND U22265 ( .A(n15381), .B(m[163]), .Z(n17240) );
  NAND U22266 ( .A(n15382), .B(creg[163]), .Z(n17239) );
  NAND U22267 ( .A(n17241), .B(n17242), .Z(y[162]) );
  NAND U22268 ( .A(n15381), .B(m[162]), .Z(n17242) );
  NAND U22269 ( .A(n15382), .B(creg[162]), .Z(n17241) );
  NAND U22270 ( .A(n17243), .B(n17244), .Z(y[161]) );
  NAND U22271 ( .A(n15381), .B(m[161]), .Z(n17244) );
  NAND U22272 ( .A(n15382), .B(creg[161]), .Z(n17243) );
  NAND U22273 ( .A(n17245), .B(n17246), .Z(y[160]) );
  NAND U22274 ( .A(n15381), .B(m[160]), .Z(n17246) );
  NAND U22275 ( .A(n15382), .B(creg[160]), .Z(n17245) );
  NAND U22276 ( .A(n17247), .B(n17248), .Z(y[15]) );
  NAND U22277 ( .A(n15381), .B(m[15]), .Z(n17248) );
  NAND U22278 ( .A(n15382), .B(creg[15]), .Z(n17247) );
  NAND U22279 ( .A(n17249), .B(n17250), .Z(y[159]) );
  NAND U22280 ( .A(n15381), .B(m[159]), .Z(n17250) );
  NAND U22281 ( .A(n15382), .B(creg[159]), .Z(n17249) );
  NAND U22282 ( .A(n17251), .B(n17252), .Z(y[158]) );
  NAND U22283 ( .A(n15381), .B(m[158]), .Z(n17252) );
  NAND U22284 ( .A(n15382), .B(creg[158]), .Z(n17251) );
  NAND U22285 ( .A(n17253), .B(n17254), .Z(y[157]) );
  NAND U22286 ( .A(n15381), .B(m[157]), .Z(n17254) );
  NAND U22287 ( .A(n15382), .B(creg[157]), .Z(n17253) );
  NAND U22288 ( .A(n17255), .B(n17256), .Z(y[156]) );
  NAND U22289 ( .A(n15381), .B(m[156]), .Z(n17256) );
  NAND U22290 ( .A(n15382), .B(creg[156]), .Z(n17255) );
  NAND U22291 ( .A(n17257), .B(n17258), .Z(y[155]) );
  NAND U22292 ( .A(n15381), .B(m[155]), .Z(n17258) );
  NAND U22293 ( .A(n15382), .B(creg[155]), .Z(n17257) );
  NAND U22294 ( .A(n17259), .B(n17260), .Z(y[154]) );
  NAND U22295 ( .A(n15381), .B(m[154]), .Z(n17260) );
  NAND U22296 ( .A(n15382), .B(creg[154]), .Z(n17259) );
  NAND U22297 ( .A(n17261), .B(n17262), .Z(y[153]) );
  NAND U22298 ( .A(n15381), .B(m[153]), .Z(n17262) );
  NAND U22299 ( .A(n15382), .B(creg[153]), .Z(n17261) );
  NAND U22300 ( .A(n17263), .B(n17264), .Z(y[152]) );
  NAND U22301 ( .A(n15381), .B(m[152]), .Z(n17264) );
  NAND U22302 ( .A(n15382), .B(creg[152]), .Z(n17263) );
  NAND U22303 ( .A(n17265), .B(n17266), .Z(y[151]) );
  NAND U22304 ( .A(n15381), .B(m[151]), .Z(n17266) );
  NAND U22305 ( .A(n15382), .B(creg[151]), .Z(n17265) );
  NAND U22306 ( .A(n17267), .B(n17268), .Z(y[150]) );
  NAND U22307 ( .A(n15381), .B(m[150]), .Z(n17268) );
  NAND U22308 ( .A(n15382), .B(creg[150]), .Z(n17267) );
  NAND U22309 ( .A(n17269), .B(n17270), .Z(y[14]) );
  NAND U22310 ( .A(n15381), .B(m[14]), .Z(n17270) );
  NAND U22311 ( .A(n15382), .B(creg[14]), .Z(n17269) );
  NAND U22312 ( .A(n17271), .B(n17272), .Z(y[149]) );
  NAND U22313 ( .A(n15381), .B(m[149]), .Z(n17272) );
  NAND U22314 ( .A(n15382), .B(creg[149]), .Z(n17271) );
  NAND U22315 ( .A(n17273), .B(n17274), .Z(y[148]) );
  NAND U22316 ( .A(n15381), .B(m[148]), .Z(n17274) );
  NAND U22317 ( .A(n15382), .B(creg[148]), .Z(n17273) );
  NAND U22318 ( .A(n17275), .B(n17276), .Z(y[147]) );
  NAND U22319 ( .A(n15381), .B(m[147]), .Z(n17276) );
  NAND U22320 ( .A(n15382), .B(creg[147]), .Z(n17275) );
  NAND U22321 ( .A(n17277), .B(n17278), .Z(y[146]) );
  NAND U22322 ( .A(n15381), .B(m[146]), .Z(n17278) );
  NAND U22323 ( .A(n15382), .B(creg[146]), .Z(n17277) );
  NAND U22324 ( .A(n17279), .B(n17280), .Z(y[145]) );
  NAND U22325 ( .A(n15381), .B(m[145]), .Z(n17280) );
  NAND U22326 ( .A(n15382), .B(creg[145]), .Z(n17279) );
  NAND U22327 ( .A(n17281), .B(n17282), .Z(y[144]) );
  NAND U22328 ( .A(n15381), .B(m[144]), .Z(n17282) );
  NAND U22329 ( .A(n15382), .B(creg[144]), .Z(n17281) );
  NAND U22330 ( .A(n17283), .B(n17284), .Z(y[143]) );
  NAND U22331 ( .A(n15381), .B(m[143]), .Z(n17284) );
  NAND U22332 ( .A(n15382), .B(creg[143]), .Z(n17283) );
  NAND U22333 ( .A(n17285), .B(n17286), .Z(y[142]) );
  NAND U22334 ( .A(n15381), .B(m[142]), .Z(n17286) );
  NAND U22335 ( .A(n15382), .B(creg[142]), .Z(n17285) );
  NAND U22336 ( .A(n17287), .B(n17288), .Z(y[141]) );
  NAND U22337 ( .A(n15381), .B(m[141]), .Z(n17288) );
  NAND U22338 ( .A(n15382), .B(creg[141]), .Z(n17287) );
  NAND U22339 ( .A(n17289), .B(n17290), .Z(y[140]) );
  NAND U22340 ( .A(n15381), .B(m[140]), .Z(n17290) );
  NAND U22341 ( .A(n15382), .B(creg[140]), .Z(n17289) );
  NAND U22342 ( .A(n17291), .B(n17292), .Z(y[13]) );
  NAND U22343 ( .A(n15381), .B(m[13]), .Z(n17292) );
  NAND U22344 ( .A(n15382), .B(creg[13]), .Z(n17291) );
  NAND U22345 ( .A(n17293), .B(n17294), .Z(y[139]) );
  NAND U22346 ( .A(n15381), .B(m[139]), .Z(n17294) );
  NAND U22347 ( .A(n15382), .B(creg[139]), .Z(n17293) );
  NAND U22348 ( .A(n17295), .B(n17296), .Z(y[138]) );
  NAND U22349 ( .A(n15381), .B(m[138]), .Z(n17296) );
  NAND U22350 ( .A(n15382), .B(creg[138]), .Z(n17295) );
  NAND U22351 ( .A(n17297), .B(n17298), .Z(y[137]) );
  NAND U22352 ( .A(n15381), .B(m[137]), .Z(n17298) );
  NAND U22353 ( .A(n15382), .B(creg[137]), .Z(n17297) );
  NAND U22354 ( .A(n17299), .B(n17300), .Z(y[136]) );
  NAND U22355 ( .A(n15381), .B(m[136]), .Z(n17300) );
  NAND U22356 ( .A(n15382), .B(creg[136]), .Z(n17299) );
  NAND U22357 ( .A(n17301), .B(n17302), .Z(y[135]) );
  NAND U22358 ( .A(n15381), .B(m[135]), .Z(n17302) );
  NAND U22359 ( .A(n15382), .B(creg[135]), .Z(n17301) );
  NAND U22360 ( .A(n17303), .B(n17304), .Z(y[134]) );
  NAND U22361 ( .A(n15381), .B(m[134]), .Z(n17304) );
  NAND U22362 ( .A(n15382), .B(creg[134]), .Z(n17303) );
  NAND U22363 ( .A(n17305), .B(n17306), .Z(y[133]) );
  NAND U22364 ( .A(n15381), .B(m[133]), .Z(n17306) );
  NAND U22365 ( .A(n15382), .B(creg[133]), .Z(n17305) );
  NAND U22366 ( .A(n17307), .B(n17308), .Z(y[132]) );
  NAND U22367 ( .A(n15381), .B(m[132]), .Z(n17308) );
  NAND U22368 ( .A(n15382), .B(creg[132]), .Z(n17307) );
  NAND U22369 ( .A(n17309), .B(n17310), .Z(y[131]) );
  NAND U22370 ( .A(n15381), .B(m[131]), .Z(n17310) );
  NAND U22371 ( .A(n15382), .B(creg[131]), .Z(n17309) );
  NAND U22372 ( .A(n17311), .B(n17312), .Z(y[130]) );
  NAND U22373 ( .A(n15381), .B(m[130]), .Z(n17312) );
  NAND U22374 ( .A(n15382), .B(creg[130]), .Z(n17311) );
  NAND U22375 ( .A(n17313), .B(n17314), .Z(y[12]) );
  NAND U22376 ( .A(n15381), .B(m[12]), .Z(n17314) );
  NAND U22377 ( .A(n15382), .B(creg[12]), .Z(n17313) );
  NAND U22378 ( .A(n17315), .B(n17316), .Z(y[129]) );
  NAND U22379 ( .A(n15381), .B(m[129]), .Z(n17316) );
  NAND U22380 ( .A(n15382), .B(creg[129]), .Z(n17315) );
  NAND U22381 ( .A(n17317), .B(n17318), .Z(y[128]) );
  NAND U22382 ( .A(n15381), .B(m[128]), .Z(n17318) );
  NAND U22383 ( .A(n15382), .B(creg[128]), .Z(n17317) );
  NAND U22384 ( .A(n17319), .B(n17320), .Z(y[127]) );
  NAND U22385 ( .A(n15381), .B(m[127]), .Z(n17320) );
  NAND U22386 ( .A(n15382), .B(creg[127]), .Z(n17319) );
  NAND U22387 ( .A(n17321), .B(n17322), .Z(y[126]) );
  NAND U22388 ( .A(n15381), .B(m[126]), .Z(n17322) );
  NAND U22389 ( .A(n15382), .B(creg[126]), .Z(n17321) );
  NAND U22390 ( .A(n17323), .B(n17324), .Z(y[125]) );
  NAND U22391 ( .A(n15381), .B(m[125]), .Z(n17324) );
  NAND U22392 ( .A(n15382), .B(creg[125]), .Z(n17323) );
  NAND U22393 ( .A(n17325), .B(n17326), .Z(y[124]) );
  NAND U22394 ( .A(n15381), .B(m[124]), .Z(n17326) );
  NAND U22395 ( .A(n15382), .B(creg[124]), .Z(n17325) );
  NAND U22396 ( .A(n17327), .B(n17328), .Z(y[123]) );
  NAND U22397 ( .A(n15381), .B(m[123]), .Z(n17328) );
  NAND U22398 ( .A(n15382), .B(creg[123]), .Z(n17327) );
  NAND U22399 ( .A(n17329), .B(n17330), .Z(y[122]) );
  NAND U22400 ( .A(n15381), .B(m[122]), .Z(n17330) );
  NAND U22401 ( .A(n15382), .B(creg[122]), .Z(n17329) );
  NAND U22402 ( .A(n17331), .B(n17332), .Z(y[121]) );
  NAND U22403 ( .A(n15381), .B(m[121]), .Z(n17332) );
  NAND U22404 ( .A(n15382), .B(creg[121]), .Z(n17331) );
  NAND U22405 ( .A(n17333), .B(n17334), .Z(y[120]) );
  NAND U22406 ( .A(n15381), .B(m[120]), .Z(n17334) );
  NAND U22407 ( .A(n15382), .B(creg[120]), .Z(n17333) );
  NAND U22408 ( .A(n17335), .B(n17336), .Z(y[11]) );
  NAND U22409 ( .A(n15381), .B(m[11]), .Z(n17336) );
  NAND U22410 ( .A(n15382), .B(creg[11]), .Z(n17335) );
  NAND U22411 ( .A(n17337), .B(n17338), .Z(y[119]) );
  NAND U22412 ( .A(n15381), .B(m[119]), .Z(n17338) );
  NAND U22413 ( .A(n15382), .B(creg[119]), .Z(n17337) );
  NAND U22414 ( .A(n17339), .B(n17340), .Z(y[118]) );
  NAND U22415 ( .A(n15381), .B(m[118]), .Z(n17340) );
  NAND U22416 ( .A(n15382), .B(creg[118]), .Z(n17339) );
  NAND U22417 ( .A(n17341), .B(n17342), .Z(y[117]) );
  NAND U22418 ( .A(n15381), .B(m[117]), .Z(n17342) );
  NAND U22419 ( .A(n15382), .B(creg[117]), .Z(n17341) );
  NAND U22420 ( .A(n17343), .B(n17344), .Z(y[116]) );
  NAND U22421 ( .A(n15381), .B(m[116]), .Z(n17344) );
  NAND U22422 ( .A(n15382), .B(creg[116]), .Z(n17343) );
  NAND U22423 ( .A(n17345), .B(n17346), .Z(y[115]) );
  NAND U22424 ( .A(n15381), .B(m[115]), .Z(n17346) );
  NAND U22425 ( .A(n15382), .B(creg[115]), .Z(n17345) );
  NAND U22426 ( .A(n17347), .B(n17348), .Z(y[114]) );
  NAND U22427 ( .A(n15381), .B(m[114]), .Z(n17348) );
  NAND U22428 ( .A(n15382), .B(creg[114]), .Z(n17347) );
  NAND U22429 ( .A(n17349), .B(n17350), .Z(y[113]) );
  NAND U22430 ( .A(n15381), .B(m[113]), .Z(n17350) );
  NAND U22431 ( .A(n15382), .B(creg[113]), .Z(n17349) );
  NAND U22432 ( .A(n17351), .B(n17352), .Z(y[112]) );
  NAND U22433 ( .A(n15381), .B(m[112]), .Z(n17352) );
  NAND U22434 ( .A(n15382), .B(creg[112]), .Z(n17351) );
  NAND U22435 ( .A(n17353), .B(n17354), .Z(y[111]) );
  NAND U22436 ( .A(n15381), .B(m[111]), .Z(n17354) );
  NAND U22437 ( .A(n15382), .B(creg[111]), .Z(n17353) );
  NAND U22438 ( .A(n17355), .B(n17356), .Z(y[110]) );
  NAND U22439 ( .A(n15381), .B(m[110]), .Z(n17356) );
  NAND U22440 ( .A(n15382), .B(creg[110]), .Z(n17355) );
  NAND U22441 ( .A(n17357), .B(n17358), .Z(y[10]) );
  NAND U22442 ( .A(n15381), .B(m[10]), .Z(n17358) );
  NAND U22443 ( .A(n15382), .B(creg[10]), .Z(n17357) );
  NAND U22444 ( .A(n17359), .B(n17360), .Z(y[109]) );
  NAND U22445 ( .A(n15381), .B(m[109]), .Z(n17360) );
  NAND U22446 ( .A(n15382), .B(creg[109]), .Z(n17359) );
  NAND U22447 ( .A(n17361), .B(n17362), .Z(y[108]) );
  NAND U22448 ( .A(n15381), .B(m[108]), .Z(n17362) );
  NAND U22449 ( .A(n15382), .B(creg[108]), .Z(n17361) );
  NAND U22450 ( .A(n17363), .B(n17364), .Z(y[107]) );
  NAND U22451 ( .A(n15381), .B(m[107]), .Z(n17364) );
  NAND U22452 ( .A(n15382), .B(creg[107]), .Z(n17363) );
  NAND U22453 ( .A(n17365), .B(n17366), .Z(y[106]) );
  NAND U22454 ( .A(n15381), .B(m[106]), .Z(n17366) );
  NAND U22455 ( .A(n15382), .B(creg[106]), .Z(n17365) );
  NAND U22456 ( .A(n17367), .B(n17368), .Z(y[105]) );
  NAND U22457 ( .A(n15381), .B(m[105]), .Z(n17368) );
  NAND U22458 ( .A(n15382), .B(creg[105]), .Z(n17367) );
  NAND U22459 ( .A(n17369), .B(n17370), .Z(y[104]) );
  NAND U22460 ( .A(n15381), .B(m[104]), .Z(n17370) );
  NAND U22461 ( .A(n15382), .B(creg[104]), .Z(n17369) );
  NAND U22462 ( .A(n17371), .B(n17372), .Z(y[103]) );
  NAND U22463 ( .A(n15381), .B(m[103]), .Z(n17372) );
  NAND U22464 ( .A(n15382), .B(creg[103]), .Z(n17371) );
  NAND U22465 ( .A(n17373), .B(n17374), .Z(y[102]) );
  NAND U22466 ( .A(n15381), .B(m[102]), .Z(n17374) );
  NAND U22467 ( .A(n15382), .B(creg[102]), .Z(n17373) );
  NAND U22468 ( .A(n17375), .B(n17376), .Z(y[1023]) );
  NAND U22469 ( .A(n15381), .B(m[1023]), .Z(n17376) );
  NAND U22470 ( .A(n15382), .B(creg[1023]), .Z(n17375) );
  NAND U22471 ( .A(n17377), .B(n17378), .Z(y[1022]) );
  NAND U22472 ( .A(n15381), .B(m[1022]), .Z(n17378) );
  NAND U22473 ( .A(n15382), .B(creg[1022]), .Z(n17377) );
  NAND U22474 ( .A(n17379), .B(n17380), .Z(y[1021]) );
  NAND U22475 ( .A(n15381), .B(m[1021]), .Z(n17380) );
  NAND U22476 ( .A(n15382), .B(creg[1021]), .Z(n17379) );
  NAND U22477 ( .A(n17381), .B(n17382), .Z(y[1020]) );
  NAND U22478 ( .A(n15381), .B(m[1020]), .Z(n17382) );
  NAND U22479 ( .A(n15382), .B(creg[1020]), .Z(n17381) );
  NAND U22480 ( .A(n17383), .B(n17384), .Z(y[101]) );
  NAND U22481 ( .A(n15381), .B(m[101]), .Z(n17384) );
  NAND U22482 ( .A(n15382), .B(creg[101]), .Z(n17383) );
  NAND U22483 ( .A(n17385), .B(n17386), .Z(y[1019]) );
  NAND U22484 ( .A(n15381), .B(m[1019]), .Z(n17386) );
  NAND U22485 ( .A(n15382), .B(creg[1019]), .Z(n17385) );
  NAND U22486 ( .A(n17387), .B(n17388), .Z(y[1018]) );
  NAND U22487 ( .A(n15381), .B(m[1018]), .Z(n17388) );
  NAND U22488 ( .A(n15382), .B(creg[1018]), .Z(n17387) );
  NAND U22489 ( .A(n17389), .B(n17390), .Z(y[1017]) );
  NAND U22490 ( .A(n15381), .B(m[1017]), .Z(n17390) );
  NAND U22491 ( .A(n15382), .B(creg[1017]), .Z(n17389) );
  NAND U22492 ( .A(n17391), .B(n17392), .Z(y[1016]) );
  NAND U22493 ( .A(n15381), .B(m[1016]), .Z(n17392) );
  NAND U22494 ( .A(n15382), .B(creg[1016]), .Z(n17391) );
  NAND U22495 ( .A(n17393), .B(n17394), .Z(y[1015]) );
  NAND U22496 ( .A(n15381), .B(m[1015]), .Z(n17394) );
  NAND U22497 ( .A(n15382), .B(creg[1015]), .Z(n17393) );
  NAND U22498 ( .A(n17395), .B(n17396), .Z(y[1014]) );
  NAND U22499 ( .A(n15381), .B(m[1014]), .Z(n17396) );
  NAND U22500 ( .A(n15382), .B(creg[1014]), .Z(n17395) );
  NAND U22501 ( .A(n17397), .B(n17398), .Z(y[1013]) );
  NAND U22502 ( .A(n15381), .B(m[1013]), .Z(n17398) );
  NAND U22503 ( .A(n15382), .B(creg[1013]), .Z(n17397) );
  NAND U22504 ( .A(n17399), .B(n17400), .Z(y[1012]) );
  NAND U22505 ( .A(n15381), .B(m[1012]), .Z(n17400) );
  NAND U22506 ( .A(n15382), .B(creg[1012]), .Z(n17399) );
  NAND U22507 ( .A(n17401), .B(n17402), .Z(y[1011]) );
  NAND U22508 ( .A(n15381), .B(m[1011]), .Z(n17402) );
  NAND U22509 ( .A(n15382), .B(creg[1011]), .Z(n17401) );
  NAND U22510 ( .A(n17403), .B(n17404), .Z(y[1010]) );
  NAND U22511 ( .A(n15381), .B(m[1010]), .Z(n17404) );
  NAND U22512 ( .A(n15382), .B(creg[1010]), .Z(n17403) );
  NAND U22513 ( .A(n17405), .B(n17406), .Z(y[100]) );
  NAND U22514 ( .A(n15381), .B(m[100]), .Z(n17406) );
  NAND U22515 ( .A(n15382), .B(creg[100]), .Z(n17405) );
  NAND U22516 ( .A(n17407), .B(n17408), .Z(y[1009]) );
  NAND U22517 ( .A(n15381), .B(m[1009]), .Z(n17408) );
  NAND U22518 ( .A(n15382), .B(creg[1009]), .Z(n17407) );
  NAND U22519 ( .A(n17409), .B(n17410), .Z(y[1008]) );
  NAND U22520 ( .A(n15381), .B(m[1008]), .Z(n17410) );
  NAND U22521 ( .A(n15382), .B(creg[1008]), .Z(n17409) );
  NAND U22522 ( .A(n17411), .B(n17412), .Z(y[1007]) );
  NAND U22523 ( .A(n15381), .B(m[1007]), .Z(n17412) );
  NAND U22524 ( .A(n15382), .B(creg[1007]), .Z(n17411) );
  NAND U22525 ( .A(n17413), .B(n17414), .Z(y[1006]) );
  NAND U22526 ( .A(n15381), .B(m[1006]), .Z(n17414) );
  NAND U22527 ( .A(n15382), .B(creg[1006]), .Z(n17413) );
  NAND U22528 ( .A(n17415), .B(n17416), .Z(y[1005]) );
  NAND U22529 ( .A(n15381), .B(m[1005]), .Z(n17416) );
  NAND U22530 ( .A(n15382), .B(creg[1005]), .Z(n17415) );
  NAND U22531 ( .A(n17417), .B(n17418), .Z(y[1004]) );
  NAND U22532 ( .A(n15381), .B(m[1004]), .Z(n17418) );
  NAND U22533 ( .A(n15382), .B(creg[1004]), .Z(n17417) );
  NAND U22534 ( .A(n17419), .B(n17420), .Z(y[1003]) );
  NAND U22535 ( .A(n15381), .B(m[1003]), .Z(n17420) );
  NAND U22536 ( .A(n15382), .B(creg[1003]), .Z(n17419) );
  NAND U22537 ( .A(n17421), .B(n17422), .Z(y[1002]) );
  NAND U22538 ( .A(n15381), .B(m[1002]), .Z(n17422) );
  NAND U22539 ( .A(n15382), .B(creg[1002]), .Z(n17421) );
  NAND U22540 ( .A(n17423), .B(n17424), .Z(y[1001]) );
  NAND U22541 ( .A(n15381), .B(m[1001]), .Z(n17424) );
  NAND U22542 ( .A(n15382), .B(creg[1001]), .Z(n17423) );
  NAND U22543 ( .A(n17425), .B(n17426), .Z(y[1000]) );
  NAND U22544 ( .A(n15381), .B(m[1000]), .Z(n17426) );
  NAND U22545 ( .A(n15382), .B(creg[1000]), .Z(n17425) );
  NAND U22546 ( .A(n17427), .B(n17428), .Z(y[0]) );
  NAND U22547 ( .A(n15381), .B(m[0]), .Z(n17428) );
  NAND U22548 ( .A(n15382), .B(creg[0]), .Z(n17427) );
  NAND U22549 ( .A(n17429), .B(n17430), .Z(x[9]) );
  NAND U22550 ( .A(creg[9]), .B(init), .Z(n17429) );
  NAND U22551 ( .A(n17431), .B(n17432), .Z(x[99]) );
  NAND U22552 ( .A(creg[99]), .B(init), .Z(n17431) );
  NAND U22553 ( .A(n17433), .B(n17434), .Z(x[999]) );
  NAND U22554 ( .A(creg[999]), .B(init), .Z(n17433) );
  NAND U22555 ( .A(n17435), .B(n17436), .Z(x[998]) );
  NAND U22556 ( .A(creg[998]), .B(init), .Z(n17435) );
  NAND U22557 ( .A(n17437), .B(n17438), .Z(x[997]) );
  NAND U22558 ( .A(creg[997]), .B(init), .Z(n17437) );
  NAND U22559 ( .A(n17439), .B(n17440), .Z(x[996]) );
  NAND U22560 ( .A(creg[996]), .B(init), .Z(n17439) );
  NAND U22561 ( .A(n17441), .B(n17442), .Z(x[995]) );
  NAND U22562 ( .A(creg[995]), .B(init), .Z(n17441) );
  NAND U22563 ( .A(n17443), .B(n17444), .Z(x[994]) );
  NAND U22564 ( .A(creg[994]), .B(init), .Z(n17443) );
  NAND U22565 ( .A(n17445), .B(n17446), .Z(x[993]) );
  NAND U22566 ( .A(creg[993]), .B(init), .Z(n17445) );
  NAND U22567 ( .A(n17447), .B(n17448), .Z(x[992]) );
  NAND U22568 ( .A(creg[992]), .B(init), .Z(n17447) );
  NAND U22569 ( .A(n17449), .B(n17450), .Z(x[991]) );
  NAND U22570 ( .A(creg[991]), .B(init), .Z(n17449) );
  NAND U22571 ( .A(n17451), .B(n17452), .Z(x[990]) );
  NAND U22572 ( .A(creg[990]), .B(init), .Z(n17451) );
  NAND U22573 ( .A(n17453), .B(n17454), .Z(x[98]) );
  NAND U22574 ( .A(creg[98]), .B(init), .Z(n17453) );
  NAND U22575 ( .A(n17455), .B(n17456), .Z(x[989]) );
  NAND U22576 ( .A(creg[989]), .B(init), .Z(n17455) );
  NAND U22577 ( .A(n17457), .B(n17458), .Z(x[988]) );
  NAND U22578 ( .A(creg[988]), .B(init), .Z(n17457) );
  NAND U22579 ( .A(n17459), .B(n17460), .Z(x[987]) );
  NAND U22580 ( .A(creg[987]), .B(init), .Z(n17459) );
  NAND U22581 ( .A(n17461), .B(n17462), .Z(x[986]) );
  NAND U22582 ( .A(creg[986]), .B(init), .Z(n17461) );
  NAND U22583 ( .A(n17463), .B(n17464), .Z(x[985]) );
  NAND U22584 ( .A(creg[985]), .B(init), .Z(n17463) );
  NAND U22585 ( .A(n17465), .B(n17466), .Z(x[984]) );
  NAND U22586 ( .A(creg[984]), .B(init), .Z(n17465) );
  NAND U22587 ( .A(n17467), .B(n17468), .Z(x[983]) );
  NAND U22588 ( .A(creg[983]), .B(init), .Z(n17467) );
  NAND U22589 ( .A(n17469), .B(n17470), .Z(x[982]) );
  NAND U22590 ( .A(creg[982]), .B(init), .Z(n17469) );
  NAND U22591 ( .A(n17471), .B(n17472), .Z(x[981]) );
  NAND U22592 ( .A(creg[981]), .B(init), .Z(n17471) );
  NAND U22593 ( .A(n17473), .B(n17474), .Z(x[980]) );
  NAND U22594 ( .A(creg[980]), .B(init), .Z(n17473) );
  NAND U22595 ( .A(n17475), .B(n17476), .Z(x[97]) );
  NAND U22596 ( .A(creg[97]), .B(init), .Z(n17475) );
  NAND U22597 ( .A(n17477), .B(n17478), .Z(x[979]) );
  NAND U22598 ( .A(creg[979]), .B(init), .Z(n17477) );
  NAND U22599 ( .A(n17479), .B(n17480), .Z(x[978]) );
  NAND U22600 ( .A(creg[978]), .B(init), .Z(n17479) );
  NAND U22601 ( .A(n17481), .B(n17482), .Z(x[977]) );
  NAND U22602 ( .A(creg[977]), .B(init), .Z(n17481) );
  NAND U22603 ( .A(n17483), .B(n17484), .Z(x[976]) );
  NAND U22604 ( .A(creg[976]), .B(init), .Z(n17483) );
  NAND U22605 ( .A(n17485), .B(n17486), .Z(x[975]) );
  NAND U22606 ( .A(creg[975]), .B(init), .Z(n17485) );
  NAND U22607 ( .A(n17487), .B(n17488), .Z(x[974]) );
  NAND U22608 ( .A(creg[974]), .B(init), .Z(n17487) );
  NAND U22609 ( .A(n17489), .B(n17490), .Z(x[973]) );
  NAND U22610 ( .A(creg[973]), .B(init), .Z(n17489) );
  NAND U22611 ( .A(n17491), .B(n17492), .Z(x[972]) );
  NAND U22612 ( .A(creg[972]), .B(init), .Z(n17491) );
  NAND U22613 ( .A(n17493), .B(n17494), .Z(x[971]) );
  NAND U22614 ( .A(creg[971]), .B(init), .Z(n17493) );
  NAND U22615 ( .A(n17495), .B(n17496), .Z(x[970]) );
  NAND U22616 ( .A(creg[970]), .B(init), .Z(n17495) );
  NAND U22617 ( .A(n17497), .B(n17498), .Z(x[96]) );
  NAND U22618 ( .A(creg[96]), .B(init), .Z(n17497) );
  NAND U22619 ( .A(n17499), .B(n17500), .Z(x[969]) );
  NAND U22620 ( .A(creg[969]), .B(init), .Z(n17499) );
  NAND U22621 ( .A(n17501), .B(n17502), .Z(x[968]) );
  NAND U22622 ( .A(creg[968]), .B(init), .Z(n17501) );
  NAND U22623 ( .A(n17503), .B(n17504), .Z(x[967]) );
  NAND U22624 ( .A(creg[967]), .B(init), .Z(n17503) );
  NAND U22625 ( .A(n17505), .B(n17506), .Z(x[966]) );
  NAND U22626 ( .A(creg[966]), .B(init), .Z(n17505) );
  NAND U22627 ( .A(n17507), .B(n17508), .Z(x[965]) );
  NAND U22628 ( .A(creg[965]), .B(init), .Z(n17507) );
  NAND U22629 ( .A(n17509), .B(n17510), .Z(x[964]) );
  NAND U22630 ( .A(creg[964]), .B(init), .Z(n17509) );
  NAND U22631 ( .A(n17511), .B(n17512), .Z(x[963]) );
  NAND U22632 ( .A(creg[963]), .B(init), .Z(n17511) );
  NAND U22633 ( .A(n17513), .B(n17514), .Z(x[962]) );
  NAND U22634 ( .A(creg[962]), .B(init), .Z(n17513) );
  NAND U22635 ( .A(n17515), .B(n17516), .Z(x[961]) );
  NAND U22636 ( .A(creg[961]), .B(init), .Z(n17515) );
  NAND U22637 ( .A(n17517), .B(n17518), .Z(x[960]) );
  NAND U22638 ( .A(creg[960]), .B(init), .Z(n17517) );
  NAND U22639 ( .A(n17519), .B(n17520), .Z(x[95]) );
  NAND U22640 ( .A(creg[95]), .B(init), .Z(n17519) );
  NAND U22641 ( .A(n17521), .B(n17522), .Z(x[959]) );
  NAND U22642 ( .A(creg[959]), .B(init), .Z(n17521) );
  NAND U22643 ( .A(n17523), .B(n17524), .Z(x[958]) );
  NAND U22644 ( .A(creg[958]), .B(init), .Z(n17523) );
  NAND U22645 ( .A(n17525), .B(n17526), .Z(x[957]) );
  NAND U22646 ( .A(creg[957]), .B(init), .Z(n17525) );
  NAND U22647 ( .A(n17527), .B(n17528), .Z(x[956]) );
  NAND U22648 ( .A(creg[956]), .B(init), .Z(n17527) );
  NAND U22649 ( .A(n17529), .B(n17530), .Z(x[955]) );
  NAND U22650 ( .A(creg[955]), .B(init), .Z(n17529) );
  NAND U22651 ( .A(n17531), .B(n17532), .Z(x[954]) );
  NAND U22652 ( .A(creg[954]), .B(init), .Z(n17531) );
  NAND U22653 ( .A(n17533), .B(n17534), .Z(x[953]) );
  NAND U22654 ( .A(creg[953]), .B(init), .Z(n17533) );
  NAND U22655 ( .A(n17535), .B(n17536), .Z(x[952]) );
  NAND U22656 ( .A(creg[952]), .B(init), .Z(n17535) );
  NAND U22657 ( .A(n17537), .B(n17538), .Z(x[951]) );
  NAND U22658 ( .A(creg[951]), .B(init), .Z(n17537) );
  NAND U22659 ( .A(n17539), .B(n17540), .Z(x[950]) );
  NAND U22660 ( .A(creg[950]), .B(init), .Z(n17539) );
  NAND U22661 ( .A(n17541), .B(n17542), .Z(x[94]) );
  NAND U22662 ( .A(creg[94]), .B(init), .Z(n17541) );
  NAND U22663 ( .A(n17543), .B(n17544), .Z(x[949]) );
  NAND U22664 ( .A(creg[949]), .B(init), .Z(n17543) );
  NAND U22665 ( .A(n17545), .B(n17546), .Z(x[948]) );
  NAND U22666 ( .A(creg[948]), .B(init), .Z(n17545) );
  NAND U22667 ( .A(n17547), .B(n17548), .Z(x[947]) );
  NAND U22668 ( .A(creg[947]), .B(init), .Z(n17547) );
  NAND U22669 ( .A(n17549), .B(n17550), .Z(x[946]) );
  NAND U22670 ( .A(creg[946]), .B(init), .Z(n17549) );
  NAND U22671 ( .A(n17551), .B(n17552), .Z(x[945]) );
  NAND U22672 ( .A(creg[945]), .B(init), .Z(n17551) );
  NAND U22673 ( .A(n17553), .B(n17554), .Z(x[944]) );
  NAND U22674 ( .A(creg[944]), .B(init), .Z(n17553) );
  NAND U22675 ( .A(n17555), .B(n17556), .Z(x[943]) );
  NAND U22676 ( .A(creg[943]), .B(init), .Z(n17555) );
  NAND U22677 ( .A(n17557), .B(n17558), .Z(x[942]) );
  NAND U22678 ( .A(creg[942]), .B(init), .Z(n17557) );
  NAND U22679 ( .A(n17559), .B(n17560), .Z(x[941]) );
  NAND U22680 ( .A(creg[941]), .B(init), .Z(n17559) );
  NAND U22681 ( .A(n17561), .B(n17562), .Z(x[940]) );
  NAND U22682 ( .A(creg[940]), .B(init), .Z(n17561) );
  NAND U22683 ( .A(n17563), .B(n17564), .Z(x[93]) );
  NAND U22684 ( .A(creg[93]), .B(init), .Z(n17563) );
  NAND U22685 ( .A(n17565), .B(n17566), .Z(x[939]) );
  NAND U22686 ( .A(creg[939]), .B(init), .Z(n17565) );
  NAND U22687 ( .A(n17567), .B(n17568), .Z(x[938]) );
  NAND U22688 ( .A(creg[938]), .B(init), .Z(n17567) );
  NAND U22689 ( .A(n17569), .B(n17570), .Z(x[937]) );
  NAND U22690 ( .A(creg[937]), .B(init), .Z(n17569) );
  NAND U22691 ( .A(n17571), .B(n17572), .Z(x[936]) );
  NAND U22692 ( .A(creg[936]), .B(init), .Z(n17571) );
  NAND U22693 ( .A(n17573), .B(n17574), .Z(x[935]) );
  NAND U22694 ( .A(creg[935]), .B(init), .Z(n17573) );
  NAND U22695 ( .A(n17575), .B(n17576), .Z(x[934]) );
  NAND U22696 ( .A(creg[934]), .B(init), .Z(n17575) );
  NAND U22697 ( .A(n17577), .B(n17578), .Z(x[933]) );
  NAND U22698 ( .A(creg[933]), .B(init), .Z(n17577) );
  NAND U22699 ( .A(n17579), .B(n17580), .Z(x[932]) );
  NAND U22700 ( .A(creg[932]), .B(init), .Z(n17579) );
  NAND U22701 ( .A(n17581), .B(n17582), .Z(x[931]) );
  NAND U22702 ( .A(creg[931]), .B(init), .Z(n17581) );
  NAND U22703 ( .A(n17583), .B(n17584), .Z(x[930]) );
  NAND U22704 ( .A(creg[930]), .B(init), .Z(n17583) );
  NAND U22705 ( .A(n17585), .B(n17586), .Z(x[92]) );
  NAND U22706 ( .A(creg[92]), .B(init), .Z(n17585) );
  NAND U22707 ( .A(n17587), .B(n17588), .Z(x[929]) );
  NAND U22708 ( .A(creg[929]), .B(init), .Z(n17587) );
  NAND U22709 ( .A(n17589), .B(n17590), .Z(x[928]) );
  NAND U22710 ( .A(creg[928]), .B(init), .Z(n17589) );
  NAND U22711 ( .A(n17591), .B(n17592), .Z(x[927]) );
  NAND U22712 ( .A(creg[927]), .B(init), .Z(n17591) );
  NAND U22713 ( .A(n17593), .B(n17594), .Z(x[926]) );
  NAND U22714 ( .A(creg[926]), .B(init), .Z(n17593) );
  NAND U22715 ( .A(n17595), .B(n17596), .Z(x[925]) );
  NAND U22716 ( .A(creg[925]), .B(init), .Z(n17595) );
  NAND U22717 ( .A(n17597), .B(n17598), .Z(x[924]) );
  NAND U22718 ( .A(creg[924]), .B(init), .Z(n17597) );
  NAND U22719 ( .A(n17599), .B(n17600), .Z(x[923]) );
  NAND U22720 ( .A(creg[923]), .B(init), .Z(n17599) );
  NAND U22721 ( .A(n17601), .B(n17602), .Z(x[922]) );
  NAND U22722 ( .A(creg[922]), .B(init), .Z(n17601) );
  NAND U22723 ( .A(n17603), .B(n17604), .Z(x[921]) );
  NAND U22724 ( .A(creg[921]), .B(init), .Z(n17603) );
  NAND U22725 ( .A(n17605), .B(n17606), .Z(x[920]) );
  NAND U22726 ( .A(creg[920]), .B(init), .Z(n17605) );
  NAND U22727 ( .A(n17607), .B(n17608), .Z(x[91]) );
  NAND U22728 ( .A(creg[91]), .B(init), .Z(n17607) );
  NAND U22729 ( .A(n17609), .B(n17610), .Z(x[919]) );
  NAND U22730 ( .A(creg[919]), .B(init), .Z(n17609) );
  NAND U22731 ( .A(n17611), .B(n17612), .Z(x[918]) );
  NAND U22732 ( .A(creg[918]), .B(init), .Z(n17611) );
  NAND U22733 ( .A(n17613), .B(n17614), .Z(x[917]) );
  NAND U22734 ( .A(creg[917]), .B(init), .Z(n17613) );
  NAND U22735 ( .A(n17615), .B(n17616), .Z(x[916]) );
  NAND U22736 ( .A(creg[916]), .B(init), .Z(n17615) );
  NAND U22737 ( .A(n17617), .B(n17618), .Z(x[915]) );
  NAND U22738 ( .A(creg[915]), .B(init), .Z(n17617) );
  NAND U22739 ( .A(n17619), .B(n17620), .Z(x[914]) );
  NAND U22740 ( .A(creg[914]), .B(init), .Z(n17619) );
  NAND U22741 ( .A(n17621), .B(n17622), .Z(x[913]) );
  NAND U22742 ( .A(creg[913]), .B(init), .Z(n17621) );
  NAND U22743 ( .A(n17623), .B(n17624), .Z(x[912]) );
  NAND U22744 ( .A(creg[912]), .B(init), .Z(n17623) );
  NAND U22745 ( .A(n17625), .B(n17626), .Z(x[911]) );
  NAND U22746 ( .A(creg[911]), .B(init), .Z(n17625) );
  NAND U22747 ( .A(n17627), .B(n17628), .Z(x[910]) );
  NAND U22748 ( .A(creg[910]), .B(init), .Z(n17627) );
  NAND U22749 ( .A(n17629), .B(n17630), .Z(x[90]) );
  NAND U22750 ( .A(creg[90]), .B(init), .Z(n17629) );
  NAND U22751 ( .A(n17631), .B(n17632), .Z(x[909]) );
  NAND U22752 ( .A(creg[909]), .B(init), .Z(n17631) );
  NAND U22753 ( .A(n17633), .B(n17634), .Z(x[908]) );
  NAND U22754 ( .A(creg[908]), .B(init), .Z(n17633) );
  NAND U22755 ( .A(n17635), .B(n17636), .Z(x[907]) );
  NAND U22756 ( .A(creg[907]), .B(init), .Z(n17635) );
  NAND U22757 ( .A(n17637), .B(n17638), .Z(x[906]) );
  NAND U22758 ( .A(creg[906]), .B(init), .Z(n17637) );
  NAND U22759 ( .A(n17639), .B(n17640), .Z(x[905]) );
  NAND U22760 ( .A(creg[905]), .B(init), .Z(n17639) );
  NAND U22761 ( .A(n17641), .B(n17642), .Z(x[904]) );
  NAND U22762 ( .A(creg[904]), .B(init), .Z(n17641) );
  NAND U22763 ( .A(n17643), .B(n17644), .Z(x[903]) );
  NAND U22764 ( .A(creg[903]), .B(init), .Z(n17643) );
  NAND U22765 ( .A(n17645), .B(n17646), .Z(x[902]) );
  NAND U22766 ( .A(creg[902]), .B(init), .Z(n17645) );
  NAND U22767 ( .A(n17647), .B(n17648), .Z(x[901]) );
  NAND U22768 ( .A(creg[901]), .B(init), .Z(n17647) );
  NAND U22769 ( .A(n17649), .B(n17650), .Z(x[900]) );
  NAND U22770 ( .A(creg[900]), .B(init), .Z(n17649) );
  NAND U22771 ( .A(n17651), .B(n17652), .Z(x[8]) );
  NAND U22772 ( .A(creg[8]), .B(init), .Z(n17651) );
  NAND U22773 ( .A(n17653), .B(n17654), .Z(x[89]) );
  NAND U22774 ( .A(creg[89]), .B(init), .Z(n17653) );
  NAND U22775 ( .A(n17655), .B(n17656), .Z(x[899]) );
  NAND U22776 ( .A(creg[899]), .B(init), .Z(n17655) );
  NAND U22777 ( .A(n17657), .B(n17658), .Z(x[898]) );
  NAND U22778 ( .A(creg[898]), .B(init), .Z(n17657) );
  NAND U22779 ( .A(n17659), .B(n17660), .Z(x[897]) );
  NAND U22780 ( .A(creg[897]), .B(init), .Z(n17659) );
  NAND U22781 ( .A(n17661), .B(n17662), .Z(x[896]) );
  NAND U22782 ( .A(creg[896]), .B(init), .Z(n17661) );
  NAND U22783 ( .A(n17663), .B(n17664), .Z(x[895]) );
  NAND U22784 ( .A(creg[895]), .B(init), .Z(n17663) );
  NAND U22785 ( .A(n17665), .B(n17666), .Z(x[894]) );
  NAND U22786 ( .A(creg[894]), .B(init), .Z(n17665) );
  NAND U22787 ( .A(n17667), .B(n17668), .Z(x[893]) );
  NAND U22788 ( .A(creg[893]), .B(init), .Z(n17667) );
  NAND U22789 ( .A(n17669), .B(n17670), .Z(x[892]) );
  NAND U22790 ( .A(creg[892]), .B(init), .Z(n17669) );
  NAND U22791 ( .A(n17671), .B(n17672), .Z(x[891]) );
  NAND U22792 ( .A(creg[891]), .B(init), .Z(n17671) );
  NAND U22793 ( .A(n17673), .B(n17674), .Z(x[890]) );
  NAND U22794 ( .A(creg[890]), .B(init), .Z(n17673) );
  NAND U22795 ( .A(n17675), .B(n17676), .Z(x[88]) );
  NAND U22796 ( .A(creg[88]), .B(init), .Z(n17675) );
  NAND U22797 ( .A(n17677), .B(n17678), .Z(x[889]) );
  NAND U22798 ( .A(creg[889]), .B(init), .Z(n17677) );
  NAND U22799 ( .A(n17679), .B(n17680), .Z(x[888]) );
  NAND U22800 ( .A(creg[888]), .B(init), .Z(n17679) );
  NAND U22801 ( .A(n17681), .B(n17682), .Z(x[887]) );
  NAND U22802 ( .A(creg[887]), .B(init), .Z(n17681) );
  NAND U22803 ( .A(n17683), .B(n17684), .Z(x[886]) );
  NAND U22804 ( .A(creg[886]), .B(init), .Z(n17683) );
  NAND U22805 ( .A(n17685), .B(n17686), .Z(x[885]) );
  NAND U22806 ( .A(creg[885]), .B(init), .Z(n17685) );
  NAND U22807 ( .A(n17687), .B(n17688), .Z(x[884]) );
  NAND U22808 ( .A(creg[884]), .B(init), .Z(n17687) );
  NAND U22809 ( .A(n17689), .B(n17690), .Z(x[883]) );
  NAND U22810 ( .A(creg[883]), .B(init), .Z(n17689) );
  NAND U22811 ( .A(n17691), .B(n17692), .Z(x[882]) );
  NAND U22812 ( .A(creg[882]), .B(init), .Z(n17691) );
  NAND U22813 ( .A(n17693), .B(n17694), .Z(x[881]) );
  NAND U22814 ( .A(creg[881]), .B(init), .Z(n17693) );
  NAND U22815 ( .A(n17695), .B(n17696), .Z(x[880]) );
  NAND U22816 ( .A(creg[880]), .B(init), .Z(n17695) );
  NAND U22817 ( .A(n17697), .B(n17698), .Z(x[87]) );
  NAND U22818 ( .A(creg[87]), .B(init), .Z(n17697) );
  NAND U22819 ( .A(n17699), .B(n17700), .Z(x[879]) );
  NAND U22820 ( .A(creg[879]), .B(init), .Z(n17699) );
  NAND U22821 ( .A(n17701), .B(n17702), .Z(x[878]) );
  NAND U22822 ( .A(creg[878]), .B(init), .Z(n17701) );
  NAND U22823 ( .A(n17703), .B(n17704), .Z(x[877]) );
  NAND U22824 ( .A(creg[877]), .B(init), .Z(n17703) );
  NAND U22825 ( .A(n17705), .B(n17706), .Z(x[876]) );
  NAND U22826 ( .A(creg[876]), .B(init), .Z(n17705) );
  NAND U22827 ( .A(n17707), .B(n17708), .Z(x[875]) );
  NAND U22828 ( .A(creg[875]), .B(init), .Z(n17707) );
  NAND U22829 ( .A(n17709), .B(n17710), .Z(x[874]) );
  NAND U22830 ( .A(creg[874]), .B(init), .Z(n17709) );
  NAND U22831 ( .A(n17711), .B(n17712), .Z(x[873]) );
  NAND U22832 ( .A(creg[873]), .B(init), .Z(n17711) );
  NAND U22833 ( .A(n17713), .B(n17714), .Z(x[872]) );
  NAND U22834 ( .A(creg[872]), .B(init), .Z(n17713) );
  NAND U22835 ( .A(n17715), .B(n17716), .Z(x[871]) );
  NAND U22836 ( .A(creg[871]), .B(init), .Z(n17715) );
  NAND U22837 ( .A(n17717), .B(n17718), .Z(x[870]) );
  NAND U22838 ( .A(creg[870]), .B(init), .Z(n17717) );
  NAND U22839 ( .A(n17719), .B(n17720), .Z(x[86]) );
  NAND U22840 ( .A(creg[86]), .B(init), .Z(n17719) );
  NAND U22841 ( .A(n17721), .B(n17722), .Z(x[869]) );
  NAND U22842 ( .A(creg[869]), .B(init), .Z(n17721) );
  NAND U22843 ( .A(n17723), .B(n17724), .Z(x[868]) );
  NAND U22844 ( .A(creg[868]), .B(init), .Z(n17723) );
  NAND U22845 ( .A(n17725), .B(n17726), .Z(x[867]) );
  NAND U22846 ( .A(creg[867]), .B(init), .Z(n17725) );
  NAND U22847 ( .A(n17727), .B(n17728), .Z(x[866]) );
  NAND U22848 ( .A(creg[866]), .B(init), .Z(n17727) );
  NAND U22849 ( .A(n17729), .B(n17730), .Z(x[865]) );
  NAND U22850 ( .A(creg[865]), .B(init), .Z(n17729) );
  NAND U22851 ( .A(n17731), .B(n17732), .Z(x[864]) );
  NAND U22852 ( .A(creg[864]), .B(init), .Z(n17731) );
  NAND U22853 ( .A(n17733), .B(n17734), .Z(x[863]) );
  NAND U22854 ( .A(creg[863]), .B(init), .Z(n17733) );
  NAND U22855 ( .A(n17735), .B(n17736), .Z(x[862]) );
  NAND U22856 ( .A(creg[862]), .B(init), .Z(n17735) );
  NAND U22857 ( .A(n17737), .B(n17738), .Z(x[861]) );
  NAND U22858 ( .A(creg[861]), .B(init), .Z(n17737) );
  NAND U22859 ( .A(n17739), .B(n17740), .Z(x[860]) );
  NAND U22860 ( .A(creg[860]), .B(init), .Z(n17739) );
  NAND U22861 ( .A(n17741), .B(n17742), .Z(x[85]) );
  NAND U22862 ( .A(creg[85]), .B(init), .Z(n17741) );
  NAND U22863 ( .A(n17743), .B(n17744), .Z(x[859]) );
  NAND U22864 ( .A(creg[859]), .B(init), .Z(n17743) );
  NAND U22865 ( .A(n17745), .B(n17746), .Z(x[858]) );
  NAND U22866 ( .A(creg[858]), .B(init), .Z(n17745) );
  NAND U22867 ( .A(n17747), .B(n17748), .Z(x[857]) );
  NAND U22868 ( .A(creg[857]), .B(init), .Z(n17747) );
  NAND U22869 ( .A(n17749), .B(n17750), .Z(x[856]) );
  NAND U22870 ( .A(creg[856]), .B(init), .Z(n17749) );
  NAND U22871 ( .A(n17751), .B(n17752), .Z(x[855]) );
  NAND U22872 ( .A(creg[855]), .B(init), .Z(n17751) );
  NAND U22873 ( .A(n17753), .B(n17754), .Z(x[854]) );
  NAND U22874 ( .A(creg[854]), .B(init), .Z(n17753) );
  NAND U22875 ( .A(n17755), .B(n17756), .Z(x[853]) );
  NAND U22876 ( .A(creg[853]), .B(init), .Z(n17755) );
  NAND U22877 ( .A(n17757), .B(n17758), .Z(x[852]) );
  NAND U22878 ( .A(creg[852]), .B(init), .Z(n17757) );
  NAND U22879 ( .A(n17759), .B(n17760), .Z(x[851]) );
  NAND U22880 ( .A(creg[851]), .B(init), .Z(n17759) );
  NAND U22881 ( .A(n17761), .B(n17762), .Z(x[850]) );
  NAND U22882 ( .A(creg[850]), .B(init), .Z(n17761) );
  NAND U22883 ( .A(n17763), .B(n17764), .Z(x[84]) );
  NAND U22884 ( .A(creg[84]), .B(init), .Z(n17763) );
  NAND U22885 ( .A(n17765), .B(n17766), .Z(x[849]) );
  NAND U22886 ( .A(creg[849]), .B(init), .Z(n17765) );
  NAND U22887 ( .A(n17767), .B(n17768), .Z(x[848]) );
  NAND U22888 ( .A(creg[848]), .B(init), .Z(n17767) );
  NAND U22889 ( .A(n17769), .B(n17770), .Z(x[847]) );
  NAND U22890 ( .A(creg[847]), .B(init), .Z(n17769) );
  NAND U22891 ( .A(n17771), .B(n17772), .Z(x[846]) );
  NAND U22892 ( .A(creg[846]), .B(init), .Z(n17771) );
  NAND U22893 ( .A(n17773), .B(n17774), .Z(x[845]) );
  NAND U22894 ( .A(creg[845]), .B(init), .Z(n17773) );
  NAND U22895 ( .A(n17775), .B(n17776), .Z(x[844]) );
  NAND U22896 ( .A(creg[844]), .B(init), .Z(n17775) );
  NAND U22897 ( .A(n17777), .B(n17778), .Z(x[843]) );
  NAND U22898 ( .A(creg[843]), .B(init), .Z(n17777) );
  NAND U22899 ( .A(n17779), .B(n17780), .Z(x[842]) );
  NAND U22900 ( .A(creg[842]), .B(init), .Z(n17779) );
  NAND U22901 ( .A(n17781), .B(n17782), .Z(x[841]) );
  NAND U22902 ( .A(creg[841]), .B(init), .Z(n17781) );
  NAND U22903 ( .A(n17783), .B(n17784), .Z(x[840]) );
  NAND U22904 ( .A(creg[840]), .B(init), .Z(n17783) );
  NAND U22905 ( .A(n17785), .B(n17786), .Z(x[83]) );
  NAND U22906 ( .A(creg[83]), .B(init), .Z(n17785) );
  NAND U22907 ( .A(n17787), .B(n17788), .Z(x[839]) );
  NAND U22908 ( .A(creg[839]), .B(init), .Z(n17787) );
  NAND U22909 ( .A(n17789), .B(n17790), .Z(x[838]) );
  NAND U22910 ( .A(creg[838]), .B(init), .Z(n17789) );
  NAND U22911 ( .A(n17791), .B(n17792), .Z(x[837]) );
  NAND U22912 ( .A(creg[837]), .B(init), .Z(n17791) );
  NAND U22913 ( .A(n17793), .B(n17794), .Z(x[836]) );
  NAND U22914 ( .A(creg[836]), .B(init), .Z(n17793) );
  NAND U22915 ( .A(n17795), .B(n17796), .Z(x[835]) );
  NAND U22916 ( .A(creg[835]), .B(init), .Z(n17795) );
  NAND U22917 ( .A(n17797), .B(n17798), .Z(x[834]) );
  NAND U22918 ( .A(creg[834]), .B(init), .Z(n17797) );
  NAND U22919 ( .A(n17799), .B(n17800), .Z(x[833]) );
  NAND U22920 ( .A(creg[833]), .B(init), .Z(n17799) );
  NAND U22921 ( .A(n17801), .B(n17802), .Z(x[832]) );
  NAND U22922 ( .A(creg[832]), .B(init), .Z(n17801) );
  NAND U22923 ( .A(n17803), .B(n17804), .Z(x[831]) );
  NAND U22924 ( .A(creg[831]), .B(init), .Z(n17803) );
  NAND U22925 ( .A(n17805), .B(n17806), .Z(x[830]) );
  NAND U22926 ( .A(creg[830]), .B(init), .Z(n17805) );
  NAND U22927 ( .A(n17807), .B(n17808), .Z(x[82]) );
  NAND U22928 ( .A(creg[82]), .B(init), .Z(n17807) );
  NAND U22929 ( .A(n17809), .B(n17810), .Z(x[829]) );
  NAND U22930 ( .A(creg[829]), .B(init), .Z(n17809) );
  NAND U22931 ( .A(n17811), .B(n17812), .Z(x[828]) );
  NAND U22932 ( .A(creg[828]), .B(init), .Z(n17811) );
  NAND U22933 ( .A(n17813), .B(n17814), .Z(x[827]) );
  NAND U22934 ( .A(creg[827]), .B(init), .Z(n17813) );
  NAND U22935 ( .A(n17815), .B(n17816), .Z(x[826]) );
  NAND U22936 ( .A(creg[826]), .B(init), .Z(n17815) );
  NAND U22937 ( .A(n17817), .B(n17818), .Z(x[825]) );
  NAND U22938 ( .A(creg[825]), .B(init), .Z(n17817) );
  NAND U22939 ( .A(n17819), .B(n17820), .Z(x[824]) );
  NAND U22940 ( .A(creg[824]), .B(init), .Z(n17819) );
  NAND U22941 ( .A(n17821), .B(n17822), .Z(x[823]) );
  NAND U22942 ( .A(creg[823]), .B(init), .Z(n17821) );
  NAND U22943 ( .A(n17823), .B(n17824), .Z(x[822]) );
  NAND U22944 ( .A(creg[822]), .B(init), .Z(n17823) );
  NAND U22945 ( .A(n17825), .B(n17826), .Z(x[821]) );
  NAND U22946 ( .A(creg[821]), .B(init), .Z(n17825) );
  NAND U22947 ( .A(n17827), .B(n17828), .Z(x[820]) );
  NAND U22948 ( .A(creg[820]), .B(init), .Z(n17827) );
  NAND U22949 ( .A(n17829), .B(n17830), .Z(x[81]) );
  NAND U22950 ( .A(creg[81]), .B(init), .Z(n17829) );
  NAND U22951 ( .A(n17831), .B(n17832), .Z(x[819]) );
  NAND U22952 ( .A(creg[819]), .B(init), .Z(n17831) );
  NAND U22953 ( .A(n17833), .B(n17834), .Z(x[818]) );
  NAND U22954 ( .A(creg[818]), .B(init), .Z(n17833) );
  NAND U22955 ( .A(n17835), .B(n17836), .Z(x[817]) );
  NAND U22956 ( .A(creg[817]), .B(init), .Z(n17835) );
  NAND U22957 ( .A(n17837), .B(n17838), .Z(x[816]) );
  NAND U22958 ( .A(creg[816]), .B(init), .Z(n17837) );
  NAND U22959 ( .A(n17839), .B(n17840), .Z(x[815]) );
  NAND U22960 ( .A(creg[815]), .B(init), .Z(n17839) );
  NAND U22961 ( .A(n17841), .B(n17842), .Z(x[814]) );
  NAND U22962 ( .A(creg[814]), .B(init), .Z(n17841) );
  NAND U22963 ( .A(n17843), .B(n17844), .Z(x[813]) );
  NAND U22964 ( .A(creg[813]), .B(init), .Z(n17843) );
  NAND U22965 ( .A(n17845), .B(n17846), .Z(x[812]) );
  NAND U22966 ( .A(creg[812]), .B(init), .Z(n17845) );
  NAND U22967 ( .A(n17847), .B(n17848), .Z(x[811]) );
  NAND U22968 ( .A(creg[811]), .B(init), .Z(n17847) );
  NAND U22969 ( .A(n17849), .B(n17850), .Z(x[810]) );
  NAND U22970 ( .A(creg[810]), .B(init), .Z(n17849) );
  NAND U22971 ( .A(n17851), .B(n17852), .Z(x[80]) );
  NAND U22972 ( .A(creg[80]), .B(init), .Z(n17851) );
  NAND U22973 ( .A(n17853), .B(n17854), .Z(x[809]) );
  NAND U22974 ( .A(creg[809]), .B(init), .Z(n17853) );
  NAND U22975 ( .A(n17855), .B(n17856), .Z(x[808]) );
  NAND U22976 ( .A(creg[808]), .B(init), .Z(n17855) );
  NAND U22977 ( .A(n17857), .B(n17858), .Z(x[807]) );
  NAND U22978 ( .A(creg[807]), .B(init), .Z(n17857) );
  NAND U22979 ( .A(n17859), .B(n17860), .Z(x[806]) );
  NAND U22980 ( .A(creg[806]), .B(init), .Z(n17859) );
  NAND U22981 ( .A(n17861), .B(n17862), .Z(x[805]) );
  NAND U22982 ( .A(creg[805]), .B(init), .Z(n17861) );
  NAND U22983 ( .A(n17863), .B(n17864), .Z(x[804]) );
  NAND U22984 ( .A(creg[804]), .B(init), .Z(n17863) );
  NAND U22985 ( .A(n17865), .B(n17866), .Z(x[803]) );
  NAND U22986 ( .A(creg[803]), .B(init), .Z(n17865) );
  NAND U22987 ( .A(n17867), .B(n17868), .Z(x[802]) );
  NAND U22988 ( .A(creg[802]), .B(init), .Z(n17867) );
  NAND U22989 ( .A(n17869), .B(n17870), .Z(x[801]) );
  NAND U22990 ( .A(creg[801]), .B(init), .Z(n17869) );
  NAND U22991 ( .A(n17871), .B(n17872), .Z(x[800]) );
  NAND U22992 ( .A(creg[800]), .B(init), .Z(n17871) );
  NAND U22993 ( .A(n17873), .B(n17874), .Z(x[7]) );
  NAND U22994 ( .A(creg[7]), .B(init), .Z(n17873) );
  NAND U22995 ( .A(n17875), .B(n17876), .Z(x[79]) );
  NAND U22996 ( .A(creg[79]), .B(init), .Z(n17875) );
  NAND U22997 ( .A(n17877), .B(n17878), .Z(x[799]) );
  NAND U22998 ( .A(creg[799]), .B(init), .Z(n17877) );
  NAND U22999 ( .A(n17879), .B(n17880), .Z(x[798]) );
  NAND U23000 ( .A(creg[798]), .B(init), .Z(n17879) );
  NAND U23001 ( .A(n17881), .B(n17882), .Z(x[797]) );
  NAND U23002 ( .A(creg[797]), .B(init), .Z(n17881) );
  NAND U23003 ( .A(n17883), .B(n17884), .Z(x[796]) );
  NAND U23004 ( .A(creg[796]), .B(init), .Z(n17883) );
  NAND U23005 ( .A(n17885), .B(n17886), .Z(x[795]) );
  NAND U23006 ( .A(creg[795]), .B(init), .Z(n17885) );
  NAND U23007 ( .A(n17887), .B(n17888), .Z(x[794]) );
  NAND U23008 ( .A(creg[794]), .B(init), .Z(n17887) );
  NAND U23009 ( .A(n17889), .B(n17890), .Z(x[793]) );
  NAND U23010 ( .A(creg[793]), .B(init), .Z(n17889) );
  NAND U23011 ( .A(n17891), .B(n17892), .Z(x[792]) );
  NAND U23012 ( .A(creg[792]), .B(init), .Z(n17891) );
  NAND U23013 ( .A(n17893), .B(n17894), .Z(x[791]) );
  NAND U23014 ( .A(creg[791]), .B(init), .Z(n17893) );
  NAND U23015 ( .A(n17895), .B(n17896), .Z(x[790]) );
  NAND U23016 ( .A(creg[790]), .B(init), .Z(n17895) );
  NAND U23017 ( .A(n17897), .B(n17898), .Z(x[78]) );
  NAND U23018 ( .A(creg[78]), .B(init), .Z(n17897) );
  NAND U23019 ( .A(n17899), .B(n17900), .Z(x[789]) );
  NAND U23020 ( .A(creg[789]), .B(init), .Z(n17899) );
  NAND U23021 ( .A(n17901), .B(n17902), .Z(x[788]) );
  NAND U23022 ( .A(creg[788]), .B(init), .Z(n17901) );
  NAND U23023 ( .A(n17903), .B(n17904), .Z(x[787]) );
  NAND U23024 ( .A(creg[787]), .B(init), .Z(n17903) );
  NAND U23025 ( .A(n17905), .B(n17906), .Z(x[786]) );
  NAND U23026 ( .A(creg[786]), .B(init), .Z(n17905) );
  NAND U23027 ( .A(n17907), .B(n17908), .Z(x[785]) );
  NAND U23028 ( .A(creg[785]), .B(init), .Z(n17907) );
  NAND U23029 ( .A(n17909), .B(n17910), .Z(x[784]) );
  NAND U23030 ( .A(creg[784]), .B(init), .Z(n17909) );
  NAND U23031 ( .A(n17911), .B(n17912), .Z(x[783]) );
  NAND U23032 ( .A(creg[783]), .B(init), .Z(n17911) );
  NAND U23033 ( .A(n17913), .B(n17914), .Z(x[782]) );
  NAND U23034 ( .A(creg[782]), .B(init), .Z(n17913) );
  NAND U23035 ( .A(n17915), .B(n17916), .Z(x[781]) );
  NAND U23036 ( .A(creg[781]), .B(init), .Z(n17915) );
  NAND U23037 ( .A(n17917), .B(n17918), .Z(x[780]) );
  NAND U23038 ( .A(creg[780]), .B(init), .Z(n17917) );
  NAND U23039 ( .A(n17919), .B(n17920), .Z(x[77]) );
  NAND U23040 ( .A(creg[77]), .B(init), .Z(n17919) );
  NAND U23041 ( .A(n17921), .B(n17922), .Z(x[779]) );
  NAND U23042 ( .A(creg[779]), .B(init), .Z(n17921) );
  NAND U23043 ( .A(n17923), .B(n17924), .Z(x[778]) );
  NAND U23044 ( .A(creg[778]), .B(init), .Z(n17923) );
  NAND U23045 ( .A(n17925), .B(n17926), .Z(x[777]) );
  NAND U23046 ( .A(creg[777]), .B(init), .Z(n17925) );
  NAND U23047 ( .A(n17927), .B(n17928), .Z(x[776]) );
  NAND U23048 ( .A(creg[776]), .B(init), .Z(n17927) );
  NAND U23049 ( .A(n17929), .B(n17930), .Z(x[775]) );
  NAND U23050 ( .A(creg[775]), .B(init), .Z(n17929) );
  NAND U23051 ( .A(n17931), .B(n17932), .Z(x[774]) );
  NAND U23052 ( .A(creg[774]), .B(init), .Z(n17931) );
  NAND U23053 ( .A(n17933), .B(n17934), .Z(x[773]) );
  NAND U23054 ( .A(creg[773]), .B(init), .Z(n17933) );
  NAND U23055 ( .A(n17935), .B(n17936), .Z(x[772]) );
  NAND U23056 ( .A(creg[772]), .B(init), .Z(n17935) );
  NAND U23057 ( .A(n17937), .B(n17938), .Z(x[771]) );
  NAND U23058 ( .A(creg[771]), .B(init), .Z(n17937) );
  NAND U23059 ( .A(n17939), .B(n17940), .Z(x[770]) );
  NAND U23060 ( .A(creg[770]), .B(init), .Z(n17939) );
  NAND U23061 ( .A(n17941), .B(n17942), .Z(x[76]) );
  NAND U23062 ( .A(creg[76]), .B(init), .Z(n17941) );
  NAND U23063 ( .A(n17943), .B(n17944), .Z(x[769]) );
  NAND U23064 ( .A(creg[769]), .B(init), .Z(n17943) );
  NAND U23065 ( .A(n17945), .B(n17946), .Z(x[768]) );
  NAND U23066 ( .A(creg[768]), .B(init), .Z(n17945) );
  NAND U23067 ( .A(n17947), .B(n17948), .Z(x[767]) );
  NAND U23068 ( .A(creg[767]), .B(init), .Z(n17947) );
  NAND U23069 ( .A(n17949), .B(n17950), .Z(x[766]) );
  NAND U23070 ( .A(creg[766]), .B(init), .Z(n17949) );
  NAND U23071 ( .A(n17951), .B(n17952), .Z(x[765]) );
  NAND U23072 ( .A(creg[765]), .B(init), .Z(n17951) );
  NAND U23073 ( .A(n17953), .B(n17954), .Z(x[764]) );
  NAND U23074 ( .A(creg[764]), .B(init), .Z(n17953) );
  NAND U23075 ( .A(n17955), .B(n17956), .Z(x[763]) );
  NAND U23076 ( .A(creg[763]), .B(init), .Z(n17955) );
  NAND U23077 ( .A(n17957), .B(n17958), .Z(x[762]) );
  NAND U23078 ( .A(creg[762]), .B(init), .Z(n17957) );
  NAND U23079 ( .A(n17959), .B(n17960), .Z(x[761]) );
  NAND U23080 ( .A(creg[761]), .B(init), .Z(n17959) );
  NAND U23081 ( .A(n17961), .B(n17962), .Z(x[760]) );
  NAND U23082 ( .A(creg[760]), .B(init), .Z(n17961) );
  NAND U23083 ( .A(n17963), .B(n17964), .Z(x[75]) );
  NAND U23084 ( .A(creg[75]), .B(init), .Z(n17963) );
  NAND U23085 ( .A(n17965), .B(n17966), .Z(x[759]) );
  NAND U23086 ( .A(creg[759]), .B(init), .Z(n17965) );
  NAND U23087 ( .A(n17967), .B(n17968), .Z(x[758]) );
  NAND U23088 ( .A(creg[758]), .B(init), .Z(n17967) );
  NAND U23089 ( .A(n17969), .B(n17970), .Z(x[757]) );
  NAND U23090 ( .A(creg[757]), .B(init), .Z(n17969) );
  NAND U23091 ( .A(n17971), .B(n17972), .Z(x[756]) );
  NAND U23092 ( .A(creg[756]), .B(init), .Z(n17971) );
  NAND U23093 ( .A(n17973), .B(n17974), .Z(x[755]) );
  NAND U23094 ( .A(creg[755]), .B(init), .Z(n17973) );
  NAND U23095 ( .A(n17975), .B(n17976), .Z(x[754]) );
  NAND U23096 ( .A(creg[754]), .B(init), .Z(n17975) );
  NAND U23097 ( .A(n17977), .B(n17978), .Z(x[753]) );
  NAND U23098 ( .A(creg[753]), .B(init), .Z(n17977) );
  NAND U23099 ( .A(n17979), .B(n17980), .Z(x[752]) );
  NAND U23100 ( .A(creg[752]), .B(init), .Z(n17979) );
  NAND U23101 ( .A(n17981), .B(n17982), .Z(x[751]) );
  NAND U23102 ( .A(creg[751]), .B(init), .Z(n17981) );
  NAND U23103 ( .A(n17983), .B(n17984), .Z(x[750]) );
  NAND U23104 ( .A(creg[750]), .B(init), .Z(n17983) );
  NAND U23105 ( .A(n17985), .B(n17986), .Z(x[74]) );
  NAND U23106 ( .A(creg[74]), .B(init), .Z(n17985) );
  NAND U23107 ( .A(n17987), .B(n17988), .Z(x[749]) );
  NAND U23108 ( .A(creg[749]), .B(init), .Z(n17987) );
  NAND U23109 ( .A(n17989), .B(n17990), .Z(x[748]) );
  NAND U23110 ( .A(creg[748]), .B(init), .Z(n17989) );
  NAND U23111 ( .A(n17991), .B(n17992), .Z(x[747]) );
  NAND U23112 ( .A(creg[747]), .B(init), .Z(n17991) );
  NAND U23113 ( .A(n17993), .B(n17994), .Z(x[746]) );
  NAND U23114 ( .A(creg[746]), .B(init), .Z(n17993) );
  NAND U23115 ( .A(n17995), .B(n17996), .Z(x[745]) );
  NAND U23116 ( .A(creg[745]), .B(init), .Z(n17995) );
  NAND U23117 ( .A(n17997), .B(n17998), .Z(x[744]) );
  NAND U23118 ( .A(creg[744]), .B(init), .Z(n17997) );
  NAND U23119 ( .A(n17999), .B(n18000), .Z(x[743]) );
  NAND U23120 ( .A(creg[743]), .B(init), .Z(n17999) );
  NAND U23121 ( .A(n18001), .B(n18002), .Z(x[742]) );
  NAND U23122 ( .A(creg[742]), .B(init), .Z(n18001) );
  NAND U23123 ( .A(n18003), .B(n18004), .Z(x[741]) );
  NAND U23124 ( .A(creg[741]), .B(init), .Z(n18003) );
  NAND U23125 ( .A(n18005), .B(n18006), .Z(x[740]) );
  NAND U23126 ( .A(creg[740]), .B(init), .Z(n18005) );
  NAND U23127 ( .A(n18007), .B(n18008), .Z(x[73]) );
  NAND U23128 ( .A(creg[73]), .B(init), .Z(n18007) );
  NAND U23129 ( .A(n18009), .B(n18010), .Z(x[739]) );
  NAND U23130 ( .A(creg[739]), .B(init), .Z(n18009) );
  NAND U23131 ( .A(n18011), .B(n18012), .Z(x[738]) );
  NAND U23132 ( .A(creg[738]), .B(init), .Z(n18011) );
  NAND U23133 ( .A(n18013), .B(n18014), .Z(x[737]) );
  NAND U23134 ( .A(creg[737]), .B(init), .Z(n18013) );
  NAND U23135 ( .A(n18015), .B(n18016), .Z(x[736]) );
  NAND U23136 ( .A(creg[736]), .B(init), .Z(n18015) );
  NAND U23137 ( .A(n18017), .B(n18018), .Z(x[735]) );
  NAND U23138 ( .A(creg[735]), .B(init), .Z(n18017) );
  NAND U23139 ( .A(n18019), .B(n18020), .Z(x[734]) );
  NAND U23140 ( .A(creg[734]), .B(init), .Z(n18019) );
  NAND U23141 ( .A(n18021), .B(n18022), .Z(x[733]) );
  NAND U23142 ( .A(creg[733]), .B(init), .Z(n18021) );
  NAND U23143 ( .A(n18023), .B(n18024), .Z(x[732]) );
  NAND U23144 ( .A(creg[732]), .B(init), .Z(n18023) );
  NAND U23145 ( .A(n18025), .B(n18026), .Z(x[731]) );
  NAND U23146 ( .A(creg[731]), .B(init), .Z(n18025) );
  NAND U23147 ( .A(n18027), .B(n18028), .Z(x[730]) );
  NAND U23148 ( .A(creg[730]), .B(init), .Z(n18027) );
  NAND U23149 ( .A(n18029), .B(n18030), .Z(x[72]) );
  NAND U23150 ( .A(creg[72]), .B(init), .Z(n18029) );
  NAND U23151 ( .A(n18031), .B(n18032), .Z(x[729]) );
  NAND U23152 ( .A(creg[729]), .B(init), .Z(n18031) );
  NAND U23153 ( .A(n18033), .B(n18034), .Z(x[728]) );
  NAND U23154 ( .A(creg[728]), .B(init), .Z(n18033) );
  NAND U23155 ( .A(n18035), .B(n18036), .Z(x[727]) );
  NAND U23156 ( .A(creg[727]), .B(init), .Z(n18035) );
  NAND U23157 ( .A(n18037), .B(n18038), .Z(x[726]) );
  NAND U23158 ( .A(creg[726]), .B(init), .Z(n18037) );
  NAND U23159 ( .A(n18039), .B(n18040), .Z(x[725]) );
  NAND U23160 ( .A(creg[725]), .B(init), .Z(n18039) );
  NAND U23161 ( .A(n18041), .B(n18042), .Z(x[724]) );
  NAND U23162 ( .A(creg[724]), .B(init), .Z(n18041) );
  NAND U23163 ( .A(n18043), .B(n18044), .Z(x[723]) );
  NAND U23164 ( .A(creg[723]), .B(init), .Z(n18043) );
  NAND U23165 ( .A(n18045), .B(n18046), .Z(x[722]) );
  NAND U23166 ( .A(creg[722]), .B(init), .Z(n18045) );
  NAND U23167 ( .A(n18047), .B(n18048), .Z(x[721]) );
  NAND U23168 ( .A(creg[721]), .B(init), .Z(n18047) );
  NAND U23169 ( .A(n18049), .B(n18050), .Z(x[720]) );
  NAND U23170 ( .A(creg[720]), .B(init), .Z(n18049) );
  NAND U23171 ( .A(n18051), .B(n18052), .Z(x[71]) );
  NAND U23172 ( .A(creg[71]), .B(init), .Z(n18051) );
  NAND U23173 ( .A(n18053), .B(n18054), .Z(x[719]) );
  NAND U23174 ( .A(creg[719]), .B(init), .Z(n18053) );
  NAND U23175 ( .A(n18055), .B(n18056), .Z(x[718]) );
  NAND U23176 ( .A(creg[718]), .B(init), .Z(n18055) );
  NAND U23177 ( .A(n18057), .B(n18058), .Z(x[717]) );
  NAND U23178 ( .A(creg[717]), .B(init), .Z(n18057) );
  NAND U23179 ( .A(n18059), .B(n18060), .Z(x[716]) );
  NAND U23180 ( .A(creg[716]), .B(init), .Z(n18059) );
  NAND U23181 ( .A(n18061), .B(n18062), .Z(x[715]) );
  NAND U23182 ( .A(creg[715]), .B(init), .Z(n18061) );
  NAND U23183 ( .A(n18063), .B(n18064), .Z(x[714]) );
  NAND U23184 ( .A(creg[714]), .B(init), .Z(n18063) );
  NAND U23185 ( .A(n18065), .B(n18066), .Z(x[713]) );
  NAND U23186 ( .A(creg[713]), .B(init), .Z(n18065) );
  NAND U23187 ( .A(n18067), .B(n18068), .Z(x[712]) );
  NAND U23188 ( .A(creg[712]), .B(init), .Z(n18067) );
  NAND U23189 ( .A(n18069), .B(n18070), .Z(x[711]) );
  NAND U23190 ( .A(creg[711]), .B(init), .Z(n18069) );
  NAND U23191 ( .A(n18071), .B(n18072), .Z(x[710]) );
  NAND U23192 ( .A(creg[710]), .B(init), .Z(n18071) );
  NAND U23193 ( .A(n18073), .B(n18074), .Z(x[70]) );
  NAND U23194 ( .A(creg[70]), .B(init), .Z(n18073) );
  NAND U23195 ( .A(n18075), .B(n18076), .Z(x[709]) );
  NAND U23196 ( .A(creg[709]), .B(init), .Z(n18075) );
  NAND U23197 ( .A(n18077), .B(n18078), .Z(x[708]) );
  NAND U23198 ( .A(creg[708]), .B(init), .Z(n18077) );
  NAND U23199 ( .A(n18079), .B(n18080), .Z(x[707]) );
  NAND U23200 ( .A(creg[707]), .B(init), .Z(n18079) );
  NAND U23201 ( .A(n18081), .B(n18082), .Z(x[706]) );
  NAND U23202 ( .A(creg[706]), .B(init), .Z(n18081) );
  NAND U23203 ( .A(n18083), .B(n18084), .Z(x[705]) );
  NAND U23204 ( .A(creg[705]), .B(init), .Z(n18083) );
  NAND U23205 ( .A(n18085), .B(n18086), .Z(x[704]) );
  NAND U23206 ( .A(creg[704]), .B(init), .Z(n18085) );
  NAND U23207 ( .A(n18087), .B(n18088), .Z(x[703]) );
  NAND U23208 ( .A(creg[703]), .B(init), .Z(n18087) );
  NAND U23209 ( .A(n18089), .B(n18090), .Z(x[702]) );
  NAND U23210 ( .A(creg[702]), .B(init), .Z(n18089) );
  NAND U23211 ( .A(n18091), .B(n18092), .Z(x[701]) );
  NAND U23212 ( .A(creg[701]), .B(init), .Z(n18091) );
  NAND U23213 ( .A(n18093), .B(n18094), .Z(x[700]) );
  NAND U23214 ( .A(creg[700]), .B(init), .Z(n18093) );
  NAND U23215 ( .A(n18095), .B(n18096), .Z(x[6]) );
  NAND U23216 ( .A(creg[6]), .B(init), .Z(n18095) );
  NAND U23217 ( .A(n18097), .B(n18098), .Z(x[69]) );
  NAND U23218 ( .A(creg[69]), .B(init), .Z(n18097) );
  NAND U23219 ( .A(n18099), .B(n18100), .Z(x[699]) );
  NAND U23220 ( .A(creg[699]), .B(init), .Z(n18099) );
  NAND U23221 ( .A(n18101), .B(n18102), .Z(x[698]) );
  NAND U23222 ( .A(creg[698]), .B(init), .Z(n18101) );
  NAND U23223 ( .A(n18103), .B(n18104), .Z(x[697]) );
  NAND U23224 ( .A(creg[697]), .B(init), .Z(n18103) );
  NAND U23225 ( .A(n18105), .B(n18106), .Z(x[696]) );
  NAND U23226 ( .A(creg[696]), .B(init), .Z(n18105) );
  NAND U23227 ( .A(n18107), .B(n18108), .Z(x[695]) );
  NAND U23228 ( .A(creg[695]), .B(init), .Z(n18107) );
  NAND U23229 ( .A(n18109), .B(n18110), .Z(x[694]) );
  NAND U23230 ( .A(creg[694]), .B(init), .Z(n18109) );
  NAND U23231 ( .A(n18111), .B(n18112), .Z(x[693]) );
  NAND U23232 ( .A(creg[693]), .B(init), .Z(n18111) );
  NAND U23233 ( .A(n18113), .B(n18114), .Z(x[692]) );
  NAND U23234 ( .A(creg[692]), .B(init), .Z(n18113) );
  NAND U23235 ( .A(n18115), .B(n18116), .Z(x[691]) );
  NAND U23236 ( .A(creg[691]), .B(init), .Z(n18115) );
  NAND U23237 ( .A(n18117), .B(n18118), .Z(x[690]) );
  NAND U23238 ( .A(creg[690]), .B(init), .Z(n18117) );
  NAND U23239 ( .A(n18119), .B(n18120), .Z(x[68]) );
  NAND U23240 ( .A(creg[68]), .B(init), .Z(n18119) );
  NAND U23241 ( .A(n18121), .B(n18122), .Z(x[689]) );
  NAND U23242 ( .A(creg[689]), .B(init), .Z(n18121) );
  NAND U23243 ( .A(n18123), .B(n18124), .Z(x[688]) );
  NAND U23244 ( .A(creg[688]), .B(init), .Z(n18123) );
  NAND U23245 ( .A(n18125), .B(n18126), .Z(x[687]) );
  NAND U23246 ( .A(creg[687]), .B(init), .Z(n18125) );
  NAND U23247 ( .A(n18127), .B(n18128), .Z(x[686]) );
  NAND U23248 ( .A(creg[686]), .B(init), .Z(n18127) );
  NAND U23249 ( .A(n18129), .B(n18130), .Z(x[685]) );
  NAND U23250 ( .A(creg[685]), .B(init), .Z(n18129) );
  NAND U23251 ( .A(n18131), .B(n18132), .Z(x[684]) );
  NAND U23252 ( .A(creg[684]), .B(init), .Z(n18131) );
  NAND U23253 ( .A(n18133), .B(n18134), .Z(x[683]) );
  NAND U23254 ( .A(creg[683]), .B(init), .Z(n18133) );
  NAND U23255 ( .A(n18135), .B(n18136), .Z(x[682]) );
  NAND U23256 ( .A(creg[682]), .B(init), .Z(n18135) );
  NAND U23257 ( .A(n18137), .B(n18138), .Z(x[681]) );
  NAND U23258 ( .A(creg[681]), .B(init), .Z(n18137) );
  NAND U23259 ( .A(n18139), .B(n18140), .Z(x[680]) );
  NAND U23260 ( .A(creg[680]), .B(init), .Z(n18139) );
  NAND U23261 ( .A(n18141), .B(n18142), .Z(x[67]) );
  NAND U23262 ( .A(creg[67]), .B(init), .Z(n18141) );
  NAND U23263 ( .A(n18143), .B(n18144), .Z(x[679]) );
  NAND U23264 ( .A(creg[679]), .B(init), .Z(n18143) );
  NAND U23265 ( .A(n18145), .B(n18146), .Z(x[678]) );
  NAND U23266 ( .A(creg[678]), .B(init), .Z(n18145) );
  NAND U23267 ( .A(n18147), .B(n18148), .Z(x[677]) );
  NAND U23268 ( .A(creg[677]), .B(init), .Z(n18147) );
  NAND U23269 ( .A(n18149), .B(n18150), .Z(x[676]) );
  NAND U23270 ( .A(creg[676]), .B(init), .Z(n18149) );
  NAND U23271 ( .A(n18151), .B(n18152), .Z(x[675]) );
  NAND U23272 ( .A(creg[675]), .B(init), .Z(n18151) );
  NAND U23273 ( .A(n18153), .B(n18154), .Z(x[674]) );
  NAND U23274 ( .A(creg[674]), .B(init), .Z(n18153) );
  NAND U23275 ( .A(n18155), .B(n18156), .Z(x[673]) );
  NAND U23276 ( .A(creg[673]), .B(init), .Z(n18155) );
  NAND U23277 ( .A(n18157), .B(n18158), .Z(x[672]) );
  NAND U23278 ( .A(creg[672]), .B(init), .Z(n18157) );
  NAND U23279 ( .A(n18159), .B(n18160), .Z(x[671]) );
  NAND U23280 ( .A(creg[671]), .B(init), .Z(n18159) );
  NAND U23281 ( .A(n18161), .B(n18162), .Z(x[670]) );
  NAND U23282 ( .A(creg[670]), .B(init), .Z(n18161) );
  NAND U23283 ( .A(n18163), .B(n18164), .Z(x[66]) );
  NAND U23284 ( .A(creg[66]), .B(init), .Z(n18163) );
  NAND U23285 ( .A(n18165), .B(n18166), .Z(x[669]) );
  NAND U23286 ( .A(creg[669]), .B(init), .Z(n18165) );
  NAND U23287 ( .A(n18167), .B(n18168), .Z(x[668]) );
  NAND U23288 ( .A(creg[668]), .B(init), .Z(n18167) );
  NAND U23289 ( .A(n18169), .B(n18170), .Z(x[667]) );
  NAND U23290 ( .A(creg[667]), .B(init), .Z(n18169) );
  NAND U23291 ( .A(n18171), .B(n18172), .Z(x[666]) );
  NAND U23292 ( .A(creg[666]), .B(init), .Z(n18171) );
  NAND U23293 ( .A(n18173), .B(n18174), .Z(x[665]) );
  NAND U23294 ( .A(creg[665]), .B(init), .Z(n18173) );
  NAND U23295 ( .A(n18175), .B(n18176), .Z(x[664]) );
  NAND U23296 ( .A(creg[664]), .B(init), .Z(n18175) );
  NAND U23297 ( .A(n18177), .B(n18178), .Z(x[663]) );
  NAND U23298 ( .A(creg[663]), .B(init), .Z(n18177) );
  NAND U23299 ( .A(n18179), .B(n18180), .Z(x[662]) );
  NAND U23300 ( .A(creg[662]), .B(init), .Z(n18179) );
  NAND U23301 ( .A(n18181), .B(n18182), .Z(x[661]) );
  NAND U23302 ( .A(creg[661]), .B(init), .Z(n18181) );
  NAND U23303 ( .A(n18183), .B(n18184), .Z(x[660]) );
  NAND U23304 ( .A(creg[660]), .B(init), .Z(n18183) );
  NAND U23305 ( .A(n18185), .B(n18186), .Z(x[65]) );
  NAND U23306 ( .A(creg[65]), .B(init), .Z(n18185) );
  NAND U23307 ( .A(n18187), .B(n18188), .Z(x[659]) );
  NAND U23308 ( .A(creg[659]), .B(init), .Z(n18187) );
  NAND U23309 ( .A(n18189), .B(n18190), .Z(x[658]) );
  NAND U23310 ( .A(creg[658]), .B(init), .Z(n18189) );
  NAND U23311 ( .A(n18191), .B(n18192), .Z(x[657]) );
  NAND U23312 ( .A(creg[657]), .B(init), .Z(n18191) );
  NAND U23313 ( .A(n18193), .B(n18194), .Z(x[656]) );
  NAND U23314 ( .A(creg[656]), .B(init), .Z(n18193) );
  NAND U23315 ( .A(n18195), .B(n18196), .Z(x[655]) );
  NAND U23316 ( .A(creg[655]), .B(init), .Z(n18195) );
  NAND U23317 ( .A(n18197), .B(n18198), .Z(x[654]) );
  NAND U23318 ( .A(creg[654]), .B(init), .Z(n18197) );
  NAND U23319 ( .A(n18199), .B(n18200), .Z(x[653]) );
  NAND U23320 ( .A(creg[653]), .B(init), .Z(n18199) );
  NAND U23321 ( .A(n18201), .B(n18202), .Z(x[652]) );
  NAND U23322 ( .A(creg[652]), .B(init), .Z(n18201) );
  NAND U23323 ( .A(n18203), .B(n18204), .Z(x[651]) );
  NAND U23324 ( .A(creg[651]), .B(init), .Z(n18203) );
  NAND U23325 ( .A(n18205), .B(n18206), .Z(x[650]) );
  NAND U23326 ( .A(creg[650]), .B(init), .Z(n18205) );
  NAND U23327 ( .A(n18207), .B(n18208), .Z(x[64]) );
  NAND U23328 ( .A(creg[64]), .B(init), .Z(n18207) );
  NAND U23329 ( .A(n18209), .B(n18210), .Z(x[649]) );
  NAND U23330 ( .A(creg[649]), .B(init), .Z(n18209) );
  NAND U23331 ( .A(n18211), .B(n18212), .Z(x[648]) );
  NAND U23332 ( .A(creg[648]), .B(init), .Z(n18211) );
  NAND U23333 ( .A(n18213), .B(n18214), .Z(x[647]) );
  NAND U23334 ( .A(creg[647]), .B(init), .Z(n18213) );
  NAND U23335 ( .A(n18215), .B(n18216), .Z(x[646]) );
  NAND U23336 ( .A(creg[646]), .B(init), .Z(n18215) );
  NAND U23337 ( .A(n18217), .B(n18218), .Z(x[645]) );
  NAND U23338 ( .A(creg[645]), .B(init), .Z(n18217) );
  NAND U23339 ( .A(n18219), .B(n18220), .Z(x[644]) );
  NAND U23340 ( .A(creg[644]), .B(init), .Z(n18219) );
  NAND U23341 ( .A(n18221), .B(n18222), .Z(x[643]) );
  NAND U23342 ( .A(creg[643]), .B(init), .Z(n18221) );
  NAND U23343 ( .A(n18223), .B(n18224), .Z(x[642]) );
  NAND U23344 ( .A(creg[642]), .B(init), .Z(n18223) );
  NAND U23345 ( .A(n18225), .B(n18226), .Z(x[641]) );
  NAND U23346 ( .A(creg[641]), .B(init), .Z(n18225) );
  NAND U23347 ( .A(n18227), .B(n18228), .Z(x[640]) );
  NAND U23348 ( .A(creg[640]), .B(init), .Z(n18227) );
  NAND U23349 ( .A(n18229), .B(n18230), .Z(x[63]) );
  NAND U23350 ( .A(creg[63]), .B(init), .Z(n18229) );
  NAND U23351 ( .A(n18231), .B(n18232), .Z(x[639]) );
  NAND U23352 ( .A(creg[639]), .B(init), .Z(n18231) );
  NAND U23353 ( .A(n18233), .B(n18234), .Z(x[638]) );
  NAND U23354 ( .A(creg[638]), .B(init), .Z(n18233) );
  NAND U23355 ( .A(n18235), .B(n18236), .Z(x[637]) );
  NAND U23356 ( .A(creg[637]), .B(init), .Z(n18235) );
  NAND U23357 ( .A(n18237), .B(n18238), .Z(x[636]) );
  NAND U23358 ( .A(creg[636]), .B(init), .Z(n18237) );
  NAND U23359 ( .A(n18239), .B(n18240), .Z(x[635]) );
  NAND U23360 ( .A(creg[635]), .B(init), .Z(n18239) );
  NAND U23361 ( .A(n18241), .B(n18242), .Z(x[634]) );
  NAND U23362 ( .A(creg[634]), .B(init), .Z(n18241) );
  NAND U23363 ( .A(n18243), .B(n18244), .Z(x[633]) );
  NAND U23364 ( .A(creg[633]), .B(init), .Z(n18243) );
  NAND U23365 ( .A(n18245), .B(n18246), .Z(x[632]) );
  NAND U23366 ( .A(creg[632]), .B(init), .Z(n18245) );
  NAND U23367 ( .A(n18247), .B(n18248), .Z(x[631]) );
  NAND U23368 ( .A(creg[631]), .B(init), .Z(n18247) );
  NAND U23369 ( .A(n18249), .B(n18250), .Z(x[630]) );
  NAND U23370 ( .A(creg[630]), .B(init), .Z(n18249) );
  NAND U23371 ( .A(n18251), .B(n18252), .Z(x[62]) );
  NAND U23372 ( .A(creg[62]), .B(init), .Z(n18251) );
  NAND U23373 ( .A(n18253), .B(n18254), .Z(x[629]) );
  NAND U23374 ( .A(creg[629]), .B(init), .Z(n18253) );
  NAND U23375 ( .A(n18255), .B(n18256), .Z(x[628]) );
  NAND U23376 ( .A(creg[628]), .B(init), .Z(n18255) );
  NAND U23377 ( .A(n18257), .B(n18258), .Z(x[627]) );
  NAND U23378 ( .A(creg[627]), .B(init), .Z(n18257) );
  NAND U23379 ( .A(n18259), .B(n18260), .Z(x[626]) );
  NAND U23380 ( .A(creg[626]), .B(init), .Z(n18259) );
  NAND U23381 ( .A(n18261), .B(n18262), .Z(x[625]) );
  NAND U23382 ( .A(creg[625]), .B(init), .Z(n18261) );
  NAND U23383 ( .A(n18263), .B(n18264), .Z(x[624]) );
  NAND U23384 ( .A(creg[624]), .B(init), .Z(n18263) );
  NAND U23385 ( .A(n18265), .B(n18266), .Z(x[623]) );
  NAND U23386 ( .A(creg[623]), .B(init), .Z(n18265) );
  NAND U23387 ( .A(n18267), .B(n18268), .Z(x[622]) );
  NAND U23388 ( .A(creg[622]), .B(init), .Z(n18267) );
  NAND U23389 ( .A(n18269), .B(n18270), .Z(x[621]) );
  NAND U23390 ( .A(creg[621]), .B(init), .Z(n18269) );
  NAND U23391 ( .A(n18271), .B(n18272), .Z(x[620]) );
  NAND U23392 ( .A(creg[620]), .B(init), .Z(n18271) );
  NAND U23393 ( .A(n18273), .B(n18274), .Z(x[61]) );
  NAND U23394 ( .A(creg[61]), .B(init), .Z(n18273) );
  NAND U23395 ( .A(n18275), .B(n18276), .Z(x[619]) );
  NAND U23396 ( .A(creg[619]), .B(init), .Z(n18275) );
  NAND U23397 ( .A(n18277), .B(n18278), .Z(x[618]) );
  NAND U23398 ( .A(creg[618]), .B(init), .Z(n18277) );
  NAND U23399 ( .A(n18279), .B(n18280), .Z(x[617]) );
  NAND U23400 ( .A(creg[617]), .B(init), .Z(n18279) );
  NAND U23401 ( .A(n18281), .B(n18282), .Z(x[616]) );
  NAND U23402 ( .A(creg[616]), .B(init), .Z(n18281) );
  NAND U23403 ( .A(n18283), .B(n18284), .Z(x[615]) );
  NAND U23404 ( .A(creg[615]), .B(init), .Z(n18283) );
  NAND U23405 ( .A(n18285), .B(n18286), .Z(x[614]) );
  NAND U23406 ( .A(creg[614]), .B(init), .Z(n18285) );
  NAND U23407 ( .A(n18287), .B(n18288), .Z(x[613]) );
  NAND U23408 ( .A(creg[613]), .B(init), .Z(n18287) );
  NAND U23409 ( .A(n18289), .B(n18290), .Z(x[612]) );
  NAND U23410 ( .A(creg[612]), .B(init), .Z(n18289) );
  NAND U23411 ( .A(n18291), .B(n18292), .Z(x[611]) );
  NAND U23412 ( .A(creg[611]), .B(init), .Z(n18291) );
  NAND U23413 ( .A(n18293), .B(n18294), .Z(x[610]) );
  NAND U23414 ( .A(creg[610]), .B(init), .Z(n18293) );
  NAND U23415 ( .A(n18295), .B(n18296), .Z(x[60]) );
  NAND U23416 ( .A(creg[60]), .B(init), .Z(n18295) );
  NAND U23417 ( .A(n18297), .B(n18298), .Z(x[609]) );
  NAND U23418 ( .A(creg[609]), .B(init), .Z(n18297) );
  NAND U23419 ( .A(n18299), .B(n18300), .Z(x[608]) );
  NAND U23420 ( .A(creg[608]), .B(init), .Z(n18299) );
  NAND U23421 ( .A(n18301), .B(n18302), .Z(x[607]) );
  NAND U23422 ( .A(creg[607]), .B(init), .Z(n18301) );
  NAND U23423 ( .A(n18303), .B(n18304), .Z(x[606]) );
  NAND U23424 ( .A(creg[606]), .B(init), .Z(n18303) );
  NAND U23425 ( .A(n18305), .B(n18306), .Z(x[605]) );
  NAND U23426 ( .A(creg[605]), .B(init), .Z(n18305) );
  NAND U23427 ( .A(n18307), .B(n18308), .Z(x[604]) );
  NAND U23428 ( .A(creg[604]), .B(init), .Z(n18307) );
  NAND U23429 ( .A(n18309), .B(n18310), .Z(x[603]) );
  NAND U23430 ( .A(creg[603]), .B(init), .Z(n18309) );
  NAND U23431 ( .A(n18311), .B(n18312), .Z(x[602]) );
  NAND U23432 ( .A(creg[602]), .B(init), .Z(n18311) );
  NAND U23433 ( .A(n18313), .B(n18314), .Z(x[601]) );
  NAND U23434 ( .A(creg[601]), .B(init), .Z(n18313) );
  NAND U23435 ( .A(n18315), .B(n18316), .Z(x[600]) );
  NAND U23436 ( .A(creg[600]), .B(init), .Z(n18315) );
  NAND U23437 ( .A(n18317), .B(n18318), .Z(x[5]) );
  NAND U23438 ( .A(creg[5]), .B(init), .Z(n18317) );
  NAND U23439 ( .A(n18319), .B(n18320), .Z(x[59]) );
  NAND U23440 ( .A(creg[59]), .B(init), .Z(n18319) );
  NAND U23441 ( .A(n18321), .B(n18322), .Z(x[599]) );
  NAND U23442 ( .A(creg[599]), .B(init), .Z(n18321) );
  NAND U23443 ( .A(n18323), .B(n18324), .Z(x[598]) );
  NAND U23444 ( .A(creg[598]), .B(init), .Z(n18323) );
  NAND U23445 ( .A(n18325), .B(n18326), .Z(x[597]) );
  NAND U23446 ( .A(creg[597]), .B(init), .Z(n18325) );
  NAND U23447 ( .A(n18327), .B(n18328), .Z(x[596]) );
  NAND U23448 ( .A(creg[596]), .B(init), .Z(n18327) );
  NAND U23449 ( .A(n18329), .B(n18330), .Z(x[595]) );
  NAND U23450 ( .A(creg[595]), .B(init), .Z(n18329) );
  NAND U23451 ( .A(n18331), .B(n18332), .Z(x[594]) );
  NAND U23452 ( .A(creg[594]), .B(init), .Z(n18331) );
  NAND U23453 ( .A(n18333), .B(n18334), .Z(x[593]) );
  NAND U23454 ( .A(creg[593]), .B(init), .Z(n18333) );
  NAND U23455 ( .A(n18335), .B(n18336), .Z(x[592]) );
  NAND U23456 ( .A(creg[592]), .B(init), .Z(n18335) );
  NAND U23457 ( .A(n18337), .B(n18338), .Z(x[591]) );
  NAND U23458 ( .A(creg[591]), .B(init), .Z(n18337) );
  NAND U23459 ( .A(n18339), .B(n18340), .Z(x[590]) );
  NAND U23460 ( .A(creg[590]), .B(init), .Z(n18339) );
  NAND U23461 ( .A(n18341), .B(n18342), .Z(x[58]) );
  NAND U23462 ( .A(creg[58]), .B(init), .Z(n18341) );
  NAND U23463 ( .A(n18343), .B(n18344), .Z(x[589]) );
  NAND U23464 ( .A(creg[589]), .B(init), .Z(n18343) );
  NAND U23465 ( .A(n18345), .B(n18346), .Z(x[588]) );
  NAND U23466 ( .A(creg[588]), .B(init), .Z(n18345) );
  NAND U23467 ( .A(n18347), .B(n18348), .Z(x[587]) );
  NAND U23468 ( .A(creg[587]), .B(init), .Z(n18347) );
  NAND U23469 ( .A(n18349), .B(n18350), .Z(x[586]) );
  NAND U23470 ( .A(creg[586]), .B(init), .Z(n18349) );
  NAND U23471 ( .A(n18351), .B(n18352), .Z(x[585]) );
  NAND U23472 ( .A(creg[585]), .B(init), .Z(n18351) );
  NAND U23473 ( .A(n18353), .B(n18354), .Z(x[584]) );
  NAND U23474 ( .A(creg[584]), .B(init), .Z(n18353) );
  NAND U23475 ( .A(n18355), .B(n18356), .Z(x[583]) );
  NAND U23476 ( .A(creg[583]), .B(init), .Z(n18355) );
  NAND U23477 ( .A(n18357), .B(n18358), .Z(x[582]) );
  NAND U23478 ( .A(creg[582]), .B(init), .Z(n18357) );
  NAND U23479 ( .A(n18359), .B(n18360), .Z(x[581]) );
  NAND U23480 ( .A(creg[581]), .B(init), .Z(n18359) );
  NAND U23481 ( .A(n18361), .B(n18362), .Z(x[580]) );
  NAND U23482 ( .A(creg[580]), .B(init), .Z(n18361) );
  NAND U23483 ( .A(n18363), .B(n18364), .Z(x[57]) );
  NAND U23484 ( .A(creg[57]), .B(init), .Z(n18363) );
  NAND U23485 ( .A(n18365), .B(n18366), .Z(x[579]) );
  NAND U23486 ( .A(creg[579]), .B(init), .Z(n18365) );
  NAND U23487 ( .A(n18367), .B(n18368), .Z(x[578]) );
  NAND U23488 ( .A(creg[578]), .B(init), .Z(n18367) );
  NAND U23489 ( .A(n18369), .B(n18370), .Z(x[577]) );
  NAND U23490 ( .A(creg[577]), .B(init), .Z(n18369) );
  NAND U23491 ( .A(n18371), .B(n18372), .Z(x[576]) );
  NAND U23492 ( .A(creg[576]), .B(init), .Z(n18371) );
  NAND U23493 ( .A(n18373), .B(n18374), .Z(x[575]) );
  NAND U23494 ( .A(creg[575]), .B(init), .Z(n18373) );
  NAND U23495 ( .A(n18375), .B(n18376), .Z(x[574]) );
  NAND U23496 ( .A(creg[574]), .B(init), .Z(n18375) );
  NAND U23497 ( .A(n18377), .B(n18378), .Z(x[573]) );
  NAND U23498 ( .A(creg[573]), .B(init), .Z(n18377) );
  NAND U23499 ( .A(n18379), .B(n18380), .Z(x[572]) );
  NAND U23500 ( .A(creg[572]), .B(init), .Z(n18379) );
  NAND U23501 ( .A(n18381), .B(n18382), .Z(x[571]) );
  NAND U23502 ( .A(creg[571]), .B(init), .Z(n18381) );
  NAND U23503 ( .A(n18383), .B(n18384), .Z(x[570]) );
  NAND U23504 ( .A(creg[570]), .B(init), .Z(n18383) );
  NAND U23505 ( .A(n18385), .B(n18386), .Z(x[56]) );
  NAND U23506 ( .A(creg[56]), .B(init), .Z(n18385) );
  NAND U23507 ( .A(n18387), .B(n18388), .Z(x[569]) );
  NAND U23508 ( .A(creg[569]), .B(init), .Z(n18387) );
  NAND U23509 ( .A(n18389), .B(n18390), .Z(x[568]) );
  NAND U23510 ( .A(creg[568]), .B(init), .Z(n18389) );
  NAND U23511 ( .A(n18391), .B(n18392), .Z(x[567]) );
  NAND U23512 ( .A(creg[567]), .B(init), .Z(n18391) );
  NAND U23513 ( .A(n18393), .B(n18394), .Z(x[566]) );
  NAND U23514 ( .A(creg[566]), .B(init), .Z(n18393) );
  NAND U23515 ( .A(n18395), .B(n18396), .Z(x[565]) );
  NAND U23516 ( .A(creg[565]), .B(init), .Z(n18395) );
  NAND U23517 ( .A(n18397), .B(n18398), .Z(x[564]) );
  NAND U23518 ( .A(creg[564]), .B(init), .Z(n18397) );
  NAND U23519 ( .A(n18399), .B(n18400), .Z(x[563]) );
  NAND U23520 ( .A(creg[563]), .B(init), .Z(n18399) );
  NAND U23521 ( .A(n18401), .B(n18402), .Z(x[562]) );
  NAND U23522 ( .A(creg[562]), .B(init), .Z(n18401) );
  NAND U23523 ( .A(n18403), .B(n18404), .Z(x[561]) );
  NAND U23524 ( .A(creg[561]), .B(init), .Z(n18403) );
  NAND U23525 ( .A(n18405), .B(n18406), .Z(x[560]) );
  NAND U23526 ( .A(creg[560]), .B(init), .Z(n18405) );
  NAND U23527 ( .A(n18407), .B(n18408), .Z(x[55]) );
  NAND U23528 ( .A(creg[55]), .B(init), .Z(n18407) );
  NAND U23529 ( .A(n18409), .B(n18410), .Z(x[559]) );
  NAND U23530 ( .A(creg[559]), .B(init), .Z(n18409) );
  NAND U23531 ( .A(n18411), .B(n18412), .Z(x[558]) );
  NAND U23532 ( .A(creg[558]), .B(init), .Z(n18411) );
  NAND U23533 ( .A(n18413), .B(n18414), .Z(x[557]) );
  NAND U23534 ( .A(creg[557]), .B(init), .Z(n18413) );
  NAND U23535 ( .A(n18415), .B(n18416), .Z(x[556]) );
  NAND U23536 ( .A(creg[556]), .B(init), .Z(n18415) );
  NAND U23537 ( .A(n18417), .B(n18418), .Z(x[555]) );
  NAND U23538 ( .A(creg[555]), .B(init), .Z(n18417) );
  NAND U23539 ( .A(n18419), .B(n18420), .Z(x[554]) );
  NAND U23540 ( .A(creg[554]), .B(init), .Z(n18419) );
  NAND U23541 ( .A(n18421), .B(n18422), .Z(x[553]) );
  NAND U23542 ( .A(creg[553]), .B(init), .Z(n18421) );
  NAND U23543 ( .A(n18423), .B(n18424), .Z(x[552]) );
  NAND U23544 ( .A(creg[552]), .B(init), .Z(n18423) );
  NAND U23545 ( .A(n18425), .B(n18426), .Z(x[551]) );
  NAND U23546 ( .A(creg[551]), .B(init), .Z(n18425) );
  NAND U23547 ( .A(n18427), .B(n18428), .Z(x[550]) );
  NAND U23548 ( .A(creg[550]), .B(init), .Z(n18427) );
  NAND U23549 ( .A(n18429), .B(n18430), .Z(x[54]) );
  NAND U23550 ( .A(creg[54]), .B(init), .Z(n18429) );
  NAND U23551 ( .A(n18431), .B(n18432), .Z(x[549]) );
  NAND U23552 ( .A(creg[549]), .B(init), .Z(n18431) );
  NAND U23553 ( .A(n18433), .B(n18434), .Z(x[548]) );
  NAND U23554 ( .A(creg[548]), .B(init), .Z(n18433) );
  NAND U23555 ( .A(n18435), .B(n18436), .Z(x[547]) );
  NAND U23556 ( .A(creg[547]), .B(init), .Z(n18435) );
  NAND U23557 ( .A(n18437), .B(n18438), .Z(x[546]) );
  NAND U23558 ( .A(creg[546]), .B(init), .Z(n18437) );
  NAND U23559 ( .A(n18439), .B(n18440), .Z(x[545]) );
  NAND U23560 ( .A(creg[545]), .B(init), .Z(n18439) );
  NAND U23561 ( .A(n18441), .B(n18442), .Z(x[544]) );
  NAND U23562 ( .A(creg[544]), .B(init), .Z(n18441) );
  NAND U23563 ( .A(n18443), .B(n18444), .Z(x[543]) );
  NAND U23564 ( .A(creg[543]), .B(init), .Z(n18443) );
  NAND U23565 ( .A(n18445), .B(n18446), .Z(x[542]) );
  NAND U23566 ( .A(creg[542]), .B(init), .Z(n18445) );
  NAND U23567 ( .A(n18447), .B(n18448), .Z(x[541]) );
  NAND U23568 ( .A(creg[541]), .B(init), .Z(n18447) );
  NAND U23569 ( .A(n18449), .B(n18450), .Z(x[540]) );
  NAND U23570 ( .A(creg[540]), .B(init), .Z(n18449) );
  NAND U23571 ( .A(n18451), .B(n18452), .Z(x[53]) );
  NAND U23572 ( .A(creg[53]), .B(init), .Z(n18451) );
  NAND U23573 ( .A(n18453), .B(n18454), .Z(x[539]) );
  NAND U23574 ( .A(creg[539]), .B(init), .Z(n18453) );
  NAND U23575 ( .A(n18455), .B(n18456), .Z(x[538]) );
  NAND U23576 ( .A(creg[538]), .B(init), .Z(n18455) );
  NAND U23577 ( .A(n18457), .B(n18458), .Z(x[537]) );
  NAND U23578 ( .A(creg[537]), .B(init), .Z(n18457) );
  NAND U23579 ( .A(n18459), .B(n18460), .Z(x[536]) );
  NAND U23580 ( .A(creg[536]), .B(init), .Z(n18459) );
  NAND U23581 ( .A(n18461), .B(n18462), .Z(x[535]) );
  NAND U23582 ( .A(creg[535]), .B(init), .Z(n18461) );
  NAND U23583 ( .A(n18463), .B(n18464), .Z(x[534]) );
  NAND U23584 ( .A(creg[534]), .B(init), .Z(n18463) );
  NAND U23585 ( .A(n18465), .B(n18466), .Z(x[533]) );
  NAND U23586 ( .A(creg[533]), .B(init), .Z(n18465) );
  NAND U23587 ( .A(n18467), .B(n18468), .Z(x[532]) );
  NAND U23588 ( .A(creg[532]), .B(init), .Z(n18467) );
  NAND U23589 ( .A(n18469), .B(n18470), .Z(x[531]) );
  NAND U23590 ( .A(creg[531]), .B(init), .Z(n18469) );
  NAND U23591 ( .A(n18471), .B(n18472), .Z(x[530]) );
  NAND U23592 ( .A(creg[530]), .B(init), .Z(n18471) );
  NAND U23593 ( .A(n18473), .B(n18474), .Z(x[52]) );
  NAND U23594 ( .A(creg[52]), .B(init), .Z(n18473) );
  NAND U23595 ( .A(n18475), .B(n18476), .Z(x[529]) );
  NAND U23596 ( .A(creg[529]), .B(init), .Z(n18475) );
  NAND U23597 ( .A(n18477), .B(n18478), .Z(x[528]) );
  NAND U23598 ( .A(creg[528]), .B(init), .Z(n18477) );
  NAND U23599 ( .A(n18479), .B(n18480), .Z(x[527]) );
  NAND U23600 ( .A(creg[527]), .B(init), .Z(n18479) );
  NAND U23601 ( .A(n18481), .B(n18482), .Z(x[526]) );
  NAND U23602 ( .A(creg[526]), .B(init), .Z(n18481) );
  NAND U23603 ( .A(n18483), .B(n18484), .Z(x[525]) );
  NAND U23604 ( .A(creg[525]), .B(init), .Z(n18483) );
  NAND U23605 ( .A(n18485), .B(n18486), .Z(x[524]) );
  NAND U23606 ( .A(creg[524]), .B(init), .Z(n18485) );
  NAND U23607 ( .A(n18487), .B(n18488), .Z(x[523]) );
  NAND U23608 ( .A(creg[523]), .B(init), .Z(n18487) );
  NAND U23609 ( .A(n18489), .B(n18490), .Z(x[522]) );
  NAND U23610 ( .A(creg[522]), .B(init), .Z(n18489) );
  NAND U23611 ( .A(n18491), .B(n18492), .Z(x[521]) );
  NAND U23612 ( .A(creg[521]), .B(init), .Z(n18491) );
  NAND U23613 ( .A(n18493), .B(n18494), .Z(x[520]) );
  NAND U23614 ( .A(creg[520]), .B(init), .Z(n18493) );
  NAND U23615 ( .A(n18495), .B(n18496), .Z(x[51]) );
  NAND U23616 ( .A(creg[51]), .B(init), .Z(n18495) );
  NAND U23617 ( .A(n18497), .B(n18498), .Z(x[519]) );
  NAND U23618 ( .A(creg[519]), .B(init), .Z(n18497) );
  NAND U23619 ( .A(n18499), .B(n18500), .Z(x[518]) );
  NAND U23620 ( .A(creg[518]), .B(init), .Z(n18499) );
  NAND U23621 ( .A(n18501), .B(n18502), .Z(x[517]) );
  NAND U23622 ( .A(creg[517]), .B(init), .Z(n18501) );
  NAND U23623 ( .A(n18503), .B(n18504), .Z(x[516]) );
  NAND U23624 ( .A(creg[516]), .B(init), .Z(n18503) );
  NAND U23625 ( .A(n18505), .B(n18506), .Z(x[515]) );
  NAND U23626 ( .A(creg[515]), .B(init), .Z(n18505) );
  NAND U23627 ( .A(n18507), .B(n18508), .Z(x[514]) );
  NAND U23628 ( .A(creg[514]), .B(init), .Z(n18507) );
  NAND U23629 ( .A(n18509), .B(n18510), .Z(x[513]) );
  NAND U23630 ( .A(creg[513]), .B(init), .Z(n18509) );
  NAND U23631 ( .A(n18511), .B(n18512), .Z(x[512]) );
  NAND U23632 ( .A(creg[512]), .B(init), .Z(n18511) );
  NAND U23633 ( .A(n18513), .B(n18514), .Z(x[511]) );
  NAND U23634 ( .A(creg[511]), .B(init), .Z(n18513) );
  NAND U23635 ( .A(n18515), .B(n18516), .Z(x[510]) );
  NAND U23636 ( .A(creg[510]), .B(init), .Z(n18515) );
  NAND U23637 ( .A(n18517), .B(n18518), .Z(x[50]) );
  NAND U23638 ( .A(creg[50]), .B(init), .Z(n18517) );
  NAND U23639 ( .A(n18519), .B(n18520), .Z(x[509]) );
  NAND U23640 ( .A(creg[509]), .B(init), .Z(n18519) );
  NAND U23641 ( .A(n18521), .B(n18522), .Z(x[508]) );
  NAND U23642 ( .A(creg[508]), .B(init), .Z(n18521) );
  NAND U23643 ( .A(n18523), .B(n18524), .Z(x[507]) );
  NAND U23644 ( .A(creg[507]), .B(init), .Z(n18523) );
  NAND U23645 ( .A(n18525), .B(n18526), .Z(x[506]) );
  NAND U23646 ( .A(creg[506]), .B(init), .Z(n18525) );
  NAND U23647 ( .A(n18527), .B(n18528), .Z(x[505]) );
  NAND U23648 ( .A(creg[505]), .B(init), .Z(n18527) );
  NAND U23649 ( .A(n18529), .B(n18530), .Z(x[504]) );
  NAND U23650 ( .A(creg[504]), .B(init), .Z(n18529) );
  NAND U23651 ( .A(n18531), .B(n18532), .Z(x[503]) );
  NAND U23652 ( .A(creg[503]), .B(init), .Z(n18531) );
  NAND U23653 ( .A(n18533), .B(n18534), .Z(x[502]) );
  NAND U23654 ( .A(creg[502]), .B(init), .Z(n18533) );
  NAND U23655 ( .A(n18535), .B(n18536), .Z(x[501]) );
  NAND U23656 ( .A(creg[501]), .B(init), .Z(n18535) );
  NAND U23657 ( .A(n18537), .B(n18538), .Z(x[500]) );
  NAND U23658 ( .A(creg[500]), .B(init), .Z(n18537) );
  NAND U23659 ( .A(n18539), .B(n18540), .Z(x[4]) );
  NAND U23660 ( .A(creg[4]), .B(init), .Z(n18539) );
  NAND U23661 ( .A(n18541), .B(n18542), .Z(x[49]) );
  NAND U23662 ( .A(creg[49]), .B(init), .Z(n18541) );
  NAND U23663 ( .A(n18543), .B(n18544), .Z(x[499]) );
  NAND U23664 ( .A(creg[499]), .B(init), .Z(n18543) );
  NAND U23665 ( .A(n18545), .B(n18546), .Z(x[498]) );
  NAND U23666 ( .A(creg[498]), .B(init), .Z(n18545) );
  NAND U23667 ( .A(n18547), .B(n18548), .Z(x[497]) );
  NAND U23668 ( .A(creg[497]), .B(init), .Z(n18547) );
  NAND U23669 ( .A(n18549), .B(n18550), .Z(x[496]) );
  NAND U23670 ( .A(creg[496]), .B(init), .Z(n18549) );
  NAND U23671 ( .A(n18551), .B(n18552), .Z(x[495]) );
  NAND U23672 ( .A(creg[495]), .B(init), .Z(n18551) );
  NAND U23673 ( .A(n18553), .B(n18554), .Z(x[494]) );
  NAND U23674 ( .A(creg[494]), .B(init), .Z(n18553) );
  NAND U23675 ( .A(n18555), .B(n18556), .Z(x[493]) );
  NAND U23676 ( .A(creg[493]), .B(init), .Z(n18555) );
  NAND U23677 ( .A(n18557), .B(n18558), .Z(x[492]) );
  NAND U23678 ( .A(creg[492]), .B(init), .Z(n18557) );
  NAND U23679 ( .A(n18559), .B(n18560), .Z(x[491]) );
  NAND U23680 ( .A(creg[491]), .B(init), .Z(n18559) );
  NAND U23681 ( .A(n18561), .B(n18562), .Z(x[490]) );
  NAND U23682 ( .A(creg[490]), .B(init), .Z(n18561) );
  NAND U23683 ( .A(n18563), .B(n18564), .Z(x[48]) );
  NAND U23684 ( .A(creg[48]), .B(init), .Z(n18563) );
  NAND U23685 ( .A(n18565), .B(n18566), .Z(x[489]) );
  NAND U23686 ( .A(creg[489]), .B(init), .Z(n18565) );
  NAND U23687 ( .A(n18567), .B(n18568), .Z(x[488]) );
  NAND U23688 ( .A(creg[488]), .B(init), .Z(n18567) );
  NAND U23689 ( .A(n18569), .B(n18570), .Z(x[487]) );
  NAND U23690 ( .A(creg[487]), .B(init), .Z(n18569) );
  NAND U23691 ( .A(n18571), .B(n18572), .Z(x[486]) );
  NAND U23692 ( .A(creg[486]), .B(init), .Z(n18571) );
  NAND U23693 ( .A(n18573), .B(n18574), .Z(x[485]) );
  NAND U23694 ( .A(creg[485]), .B(init), .Z(n18573) );
  NAND U23695 ( .A(n18575), .B(n18576), .Z(x[484]) );
  NAND U23696 ( .A(creg[484]), .B(init), .Z(n18575) );
  NAND U23697 ( .A(n18577), .B(n18578), .Z(x[483]) );
  NAND U23698 ( .A(creg[483]), .B(init), .Z(n18577) );
  NAND U23699 ( .A(n18579), .B(n18580), .Z(x[482]) );
  NAND U23700 ( .A(creg[482]), .B(init), .Z(n18579) );
  NAND U23701 ( .A(n18581), .B(n18582), .Z(x[481]) );
  NAND U23702 ( .A(creg[481]), .B(init), .Z(n18581) );
  NAND U23703 ( .A(n18583), .B(n18584), .Z(x[480]) );
  NAND U23704 ( .A(creg[480]), .B(init), .Z(n18583) );
  NAND U23705 ( .A(n18585), .B(n18586), .Z(x[47]) );
  NAND U23706 ( .A(creg[47]), .B(init), .Z(n18585) );
  NAND U23707 ( .A(n18587), .B(n18588), .Z(x[479]) );
  NAND U23708 ( .A(creg[479]), .B(init), .Z(n18587) );
  NAND U23709 ( .A(n18589), .B(n18590), .Z(x[478]) );
  NAND U23710 ( .A(creg[478]), .B(init), .Z(n18589) );
  NAND U23711 ( .A(n18591), .B(n18592), .Z(x[477]) );
  NAND U23712 ( .A(creg[477]), .B(init), .Z(n18591) );
  NAND U23713 ( .A(n18593), .B(n18594), .Z(x[476]) );
  NAND U23714 ( .A(creg[476]), .B(init), .Z(n18593) );
  NAND U23715 ( .A(n18595), .B(n18596), .Z(x[475]) );
  NAND U23716 ( .A(creg[475]), .B(init), .Z(n18595) );
  NAND U23717 ( .A(n18597), .B(n18598), .Z(x[474]) );
  NAND U23718 ( .A(creg[474]), .B(init), .Z(n18597) );
  NAND U23719 ( .A(n18599), .B(n18600), .Z(x[473]) );
  NAND U23720 ( .A(creg[473]), .B(init), .Z(n18599) );
  NAND U23721 ( .A(n18601), .B(n18602), .Z(x[472]) );
  NAND U23722 ( .A(creg[472]), .B(init), .Z(n18601) );
  NAND U23723 ( .A(n18603), .B(n18604), .Z(x[471]) );
  NAND U23724 ( .A(creg[471]), .B(init), .Z(n18603) );
  NAND U23725 ( .A(n18605), .B(n18606), .Z(x[470]) );
  NAND U23726 ( .A(creg[470]), .B(init), .Z(n18605) );
  NAND U23727 ( .A(n18607), .B(n18608), .Z(x[46]) );
  NAND U23728 ( .A(creg[46]), .B(init), .Z(n18607) );
  NAND U23729 ( .A(n18609), .B(n18610), .Z(x[469]) );
  NAND U23730 ( .A(creg[469]), .B(init), .Z(n18609) );
  NAND U23731 ( .A(n18611), .B(n18612), .Z(x[468]) );
  NAND U23732 ( .A(creg[468]), .B(init), .Z(n18611) );
  NAND U23733 ( .A(n18613), .B(n18614), .Z(x[467]) );
  NAND U23734 ( .A(creg[467]), .B(init), .Z(n18613) );
  NAND U23735 ( .A(n18615), .B(n18616), .Z(x[466]) );
  NAND U23736 ( .A(creg[466]), .B(init), .Z(n18615) );
  NAND U23737 ( .A(n18617), .B(n18618), .Z(x[465]) );
  NAND U23738 ( .A(creg[465]), .B(init), .Z(n18617) );
  NAND U23739 ( .A(n18619), .B(n18620), .Z(x[464]) );
  NAND U23740 ( .A(creg[464]), .B(init), .Z(n18619) );
  NAND U23741 ( .A(n18621), .B(n18622), .Z(x[463]) );
  NAND U23742 ( .A(creg[463]), .B(init), .Z(n18621) );
  NAND U23743 ( .A(n18623), .B(n18624), .Z(x[462]) );
  NAND U23744 ( .A(creg[462]), .B(init), .Z(n18623) );
  NAND U23745 ( .A(n18625), .B(n18626), .Z(x[461]) );
  NAND U23746 ( .A(creg[461]), .B(init), .Z(n18625) );
  NAND U23747 ( .A(n18627), .B(n18628), .Z(x[460]) );
  NAND U23748 ( .A(creg[460]), .B(init), .Z(n18627) );
  NAND U23749 ( .A(n18629), .B(n18630), .Z(x[45]) );
  NAND U23750 ( .A(creg[45]), .B(init), .Z(n18629) );
  NAND U23751 ( .A(n18631), .B(n18632), .Z(x[459]) );
  NAND U23752 ( .A(creg[459]), .B(init), .Z(n18631) );
  NAND U23753 ( .A(n18633), .B(n18634), .Z(x[458]) );
  NAND U23754 ( .A(creg[458]), .B(init), .Z(n18633) );
  NAND U23755 ( .A(n18635), .B(n18636), .Z(x[457]) );
  NAND U23756 ( .A(creg[457]), .B(init), .Z(n18635) );
  NAND U23757 ( .A(n18637), .B(n18638), .Z(x[456]) );
  NAND U23758 ( .A(creg[456]), .B(init), .Z(n18637) );
  NAND U23759 ( .A(n18639), .B(n18640), .Z(x[455]) );
  NAND U23760 ( .A(creg[455]), .B(init), .Z(n18639) );
  NAND U23761 ( .A(n18641), .B(n18642), .Z(x[454]) );
  NAND U23762 ( .A(creg[454]), .B(init), .Z(n18641) );
  NAND U23763 ( .A(n18643), .B(n18644), .Z(x[453]) );
  NAND U23764 ( .A(creg[453]), .B(init), .Z(n18643) );
  NAND U23765 ( .A(n18645), .B(n18646), .Z(x[452]) );
  NAND U23766 ( .A(creg[452]), .B(init), .Z(n18645) );
  NAND U23767 ( .A(n18647), .B(n18648), .Z(x[451]) );
  NAND U23768 ( .A(creg[451]), .B(init), .Z(n18647) );
  NAND U23769 ( .A(n18649), .B(n18650), .Z(x[450]) );
  NAND U23770 ( .A(creg[450]), .B(init), .Z(n18649) );
  NAND U23771 ( .A(n18651), .B(n18652), .Z(x[44]) );
  NAND U23772 ( .A(creg[44]), .B(init), .Z(n18651) );
  NAND U23773 ( .A(n18653), .B(n18654), .Z(x[449]) );
  NAND U23774 ( .A(creg[449]), .B(init), .Z(n18653) );
  NAND U23775 ( .A(n18655), .B(n18656), .Z(x[448]) );
  NAND U23776 ( .A(creg[448]), .B(init), .Z(n18655) );
  NAND U23777 ( .A(n18657), .B(n18658), .Z(x[447]) );
  NAND U23778 ( .A(creg[447]), .B(init), .Z(n18657) );
  NAND U23779 ( .A(n18659), .B(n18660), .Z(x[446]) );
  NAND U23780 ( .A(creg[446]), .B(init), .Z(n18659) );
  NAND U23781 ( .A(n18661), .B(n18662), .Z(x[445]) );
  NAND U23782 ( .A(creg[445]), .B(init), .Z(n18661) );
  NAND U23783 ( .A(n18663), .B(n18664), .Z(x[444]) );
  NAND U23784 ( .A(creg[444]), .B(init), .Z(n18663) );
  NAND U23785 ( .A(n18665), .B(n18666), .Z(x[443]) );
  NAND U23786 ( .A(creg[443]), .B(init), .Z(n18665) );
  NAND U23787 ( .A(n18667), .B(n18668), .Z(x[442]) );
  NAND U23788 ( .A(creg[442]), .B(init), .Z(n18667) );
  NAND U23789 ( .A(n18669), .B(n18670), .Z(x[441]) );
  NAND U23790 ( .A(creg[441]), .B(init), .Z(n18669) );
  NAND U23791 ( .A(n18671), .B(n18672), .Z(x[440]) );
  NAND U23792 ( .A(creg[440]), .B(init), .Z(n18671) );
  NAND U23793 ( .A(n18673), .B(n18674), .Z(x[43]) );
  NAND U23794 ( .A(creg[43]), .B(init), .Z(n18673) );
  NAND U23795 ( .A(n18675), .B(n18676), .Z(x[439]) );
  NAND U23796 ( .A(creg[439]), .B(init), .Z(n18675) );
  NAND U23797 ( .A(n18677), .B(n18678), .Z(x[438]) );
  NAND U23798 ( .A(creg[438]), .B(init), .Z(n18677) );
  NAND U23799 ( .A(n18679), .B(n18680), .Z(x[437]) );
  NAND U23800 ( .A(creg[437]), .B(init), .Z(n18679) );
  NAND U23801 ( .A(n18681), .B(n18682), .Z(x[436]) );
  NAND U23802 ( .A(creg[436]), .B(init), .Z(n18681) );
  NAND U23803 ( .A(n18683), .B(n18684), .Z(x[435]) );
  NAND U23804 ( .A(creg[435]), .B(init), .Z(n18683) );
  NAND U23805 ( .A(n18685), .B(n18686), .Z(x[434]) );
  NAND U23806 ( .A(creg[434]), .B(init), .Z(n18685) );
  NAND U23807 ( .A(n18687), .B(n18688), .Z(x[433]) );
  NAND U23808 ( .A(creg[433]), .B(init), .Z(n18687) );
  NAND U23809 ( .A(n18689), .B(n18690), .Z(x[432]) );
  NAND U23810 ( .A(creg[432]), .B(init), .Z(n18689) );
  NAND U23811 ( .A(n18691), .B(n18692), .Z(x[431]) );
  NAND U23812 ( .A(creg[431]), .B(init), .Z(n18691) );
  NAND U23813 ( .A(n18693), .B(n18694), .Z(x[430]) );
  NAND U23814 ( .A(creg[430]), .B(init), .Z(n18693) );
  NAND U23815 ( .A(n18695), .B(n18696), .Z(x[42]) );
  NAND U23816 ( .A(creg[42]), .B(init), .Z(n18695) );
  NAND U23817 ( .A(n18697), .B(n18698), .Z(x[429]) );
  NAND U23818 ( .A(creg[429]), .B(init), .Z(n18697) );
  NAND U23819 ( .A(n18699), .B(n18700), .Z(x[428]) );
  NAND U23820 ( .A(creg[428]), .B(init), .Z(n18699) );
  NAND U23821 ( .A(n18701), .B(n18702), .Z(x[427]) );
  NAND U23822 ( .A(creg[427]), .B(init), .Z(n18701) );
  NAND U23823 ( .A(n18703), .B(n18704), .Z(x[426]) );
  NAND U23824 ( .A(creg[426]), .B(init), .Z(n18703) );
  NAND U23825 ( .A(n18705), .B(n18706), .Z(x[425]) );
  NAND U23826 ( .A(creg[425]), .B(init), .Z(n18705) );
  NAND U23827 ( .A(n18707), .B(n18708), .Z(x[424]) );
  NAND U23828 ( .A(creg[424]), .B(init), .Z(n18707) );
  NAND U23829 ( .A(n18709), .B(n18710), .Z(x[423]) );
  NAND U23830 ( .A(creg[423]), .B(init), .Z(n18709) );
  NAND U23831 ( .A(n18711), .B(n18712), .Z(x[422]) );
  NAND U23832 ( .A(creg[422]), .B(init), .Z(n18711) );
  NAND U23833 ( .A(n18713), .B(n18714), .Z(x[421]) );
  NAND U23834 ( .A(creg[421]), .B(init), .Z(n18713) );
  NAND U23835 ( .A(n18715), .B(n18716), .Z(x[420]) );
  NAND U23836 ( .A(creg[420]), .B(init), .Z(n18715) );
  NAND U23837 ( .A(n18717), .B(n18718), .Z(x[41]) );
  NAND U23838 ( .A(creg[41]), .B(init), .Z(n18717) );
  NAND U23839 ( .A(n18719), .B(n18720), .Z(x[419]) );
  NAND U23840 ( .A(creg[419]), .B(init), .Z(n18719) );
  NAND U23841 ( .A(n18721), .B(n18722), .Z(x[418]) );
  NAND U23842 ( .A(creg[418]), .B(init), .Z(n18721) );
  NAND U23843 ( .A(n18723), .B(n18724), .Z(x[417]) );
  NAND U23844 ( .A(creg[417]), .B(init), .Z(n18723) );
  NAND U23845 ( .A(n18725), .B(n18726), .Z(x[416]) );
  NAND U23846 ( .A(creg[416]), .B(init), .Z(n18725) );
  NAND U23847 ( .A(n18727), .B(n18728), .Z(x[415]) );
  NAND U23848 ( .A(creg[415]), .B(init), .Z(n18727) );
  NAND U23849 ( .A(n18729), .B(n18730), .Z(x[414]) );
  NAND U23850 ( .A(creg[414]), .B(init), .Z(n18729) );
  NAND U23851 ( .A(n18731), .B(n18732), .Z(x[413]) );
  NAND U23852 ( .A(creg[413]), .B(init), .Z(n18731) );
  NAND U23853 ( .A(n18733), .B(n18734), .Z(x[412]) );
  NAND U23854 ( .A(creg[412]), .B(init), .Z(n18733) );
  NAND U23855 ( .A(n18735), .B(n18736), .Z(x[411]) );
  NAND U23856 ( .A(creg[411]), .B(init), .Z(n18735) );
  NAND U23857 ( .A(n18737), .B(n18738), .Z(x[410]) );
  NAND U23858 ( .A(creg[410]), .B(init), .Z(n18737) );
  NAND U23859 ( .A(n18739), .B(n18740), .Z(x[40]) );
  NAND U23860 ( .A(creg[40]), .B(init), .Z(n18739) );
  NAND U23861 ( .A(n18741), .B(n18742), .Z(x[409]) );
  NAND U23862 ( .A(creg[409]), .B(init), .Z(n18741) );
  NAND U23863 ( .A(n18743), .B(n18744), .Z(x[408]) );
  NAND U23864 ( .A(creg[408]), .B(init), .Z(n18743) );
  NAND U23865 ( .A(n18745), .B(n18746), .Z(x[407]) );
  NAND U23866 ( .A(creg[407]), .B(init), .Z(n18745) );
  NAND U23867 ( .A(n18747), .B(n18748), .Z(x[406]) );
  NAND U23868 ( .A(creg[406]), .B(init), .Z(n18747) );
  NAND U23869 ( .A(n18749), .B(n18750), .Z(x[405]) );
  NAND U23870 ( .A(creg[405]), .B(init), .Z(n18749) );
  NAND U23871 ( .A(n18751), .B(n18752), .Z(x[404]) );
  NAND U23872 ( .A(creg[404]), .B(init), .Z(n18751) );
  NAND U23873 ( .A(n18753), .B(n18754), .Z(x[403]) );
  NAND U23874 ( .A(creg[403]), .B(init), .Z(n18753) );
  NAND U23875 ( .A(n18755), .B(n18756), .Z(x[402]) );
  NAND U23876 ( .A(creg[402]), .B(init), .Z(n18755) );
  NAND U23877 ( .A(n18757), .B(n18758), .Z(x[401]) );
  NAND U23878 ( .A(creg[401]), .B(init), .Z(n18757) );
  NAND U23879 ( .A(n18759), .B(n18760), .Z(x[400]) );
  NAND U23880 ( .A(creg[400]), .B(init), .Z(n18759) );
  NAND U23881 ( .A(n18761), .B(n18762), .Z(x[3]) );
  NAND U23882 ( .A(creg[3]), .B(init), .Z(n18761) );
  NAND U23883 ( .A(n18763), .B(n18764), .Z(x[39]) );
  NAND U23884 ( .A(creg[39]), .B(init), .Z(n18763) );
  NAND U23885 ( .A(n18765), .B(n18766), .Z(x[399]) );
  NAND U23886 ( .A(creg[399]), .B(init), .Z(n18765) );
  NAND U23887 ( .A(n18767), .B(n18768), .Z(x[398]) );
  NAND U23888 ( .A(creg[398]), .B(init), .Z(n18767) );
  NAND U23889 ( .A(n18769), .B(n18770), .Z(x[397]) );
  NAND U23890 ( .A(creg[397]), .B(init), .Z(n18769) );
  NAND U23891 ( .A(n18771), .B(n18772), .Z(x[396]) );
  NAND U23892 ( .A(creg[396]), .B(init), .Z(n18771) );
  NAND U23893 ( .A(n18773), .B(n18774), .Z(x[395]) );
  NAND U23894 ( .A(creg[395]), .B(init), .Z(n18773) );
  NAND U23895 ( .A(n18775), .B(n18776), .Z(x[394]) );
  NAND U23896 ( .A(creg[394]), .B(init), .Z(n18775) );
  NAND U23897 ( .A(n18777), .B(n18778), .Z(x[393]) );
  NAND U23898 ( .A(creg[393]), .B(init), .Z(n18777) );
  NAND U23899 ( .A(n18779), .B(n18780), .Z(x[392]) );
  NAND U23900 ( .A(creg[392]), .B(init), .Z(n18779) );
  NAND U23901 ( .A(n18781), .B(n18782), .Z(x[391]) );
  NAND U23902 ( .A(creg[391]), .B(init), .Z(n18781) );
  NAND U23903 ( .A(n18783), .B(n18784), .Z(x[390]) );
  NAND U23904 ( .A(creg[390]), .B(init), .Z(n18783) );
  NAND U23905 ( .A(n18785), .B(n18786), .Z(x[38]) );
  NAND U23906 ( .A(creg[38]), .B(init), .Z(n18785) );
  NAND U23907 ( .A(n18787), .B(n18788), .Z(x[389]) );
  NAND U23908 ( .A(creg[389]), .B(init), .Z(n18787) );
  NAND U23909 ( .A(n18789), .B(n18790), .Z(x[388]) );
  NAND U23910 ( .A(creg[388]), .B(init), .Z(n18789) );
  NAND U23911 ( .A(n18791), .B(n18792), .Z(x[387]) );
  NAND U23912 ( .A(creg[387]), .B(init), .Z(n18791) );
  NAND U23913 ( .A(n18793), .B(n18794), .Z(x[386]) );
  NAND U23914 ( .A(creg[386]), .B(init), .Z(n18793) );
  NAND U23915 ( .A(n18795), .B(n18796), .Z(x[385]) );
  NAND U23916 ( .A(creg[385]), .B(init), .Z(n18795) );
  NAND U23917 ( .A(n18797), .B(n18798), .Z(x[384]) );
  NAND U23918 ( .A(creg[384]), .B(init), .Z(n18797) );
  NAND U23919 ( .A(n18799), .B(n18800), .Z(x[383]) );
  NAND U23920 ( .A(creg[383]), .B(init), .Z(n18799) );
  NAND U23921 ( .A(n18801), .B(n18802), .Z(x[382]) );
  NAND U23922 ( .A(creg[382]), .B(init), .Z(n18801) );
  NAND U23923 ( .A(n18803), .B(n18804), .Z(x[381]) );
  NAND U23924 ( .A(creg[381]), .B(init), .Z(n18803) );
  NAND U23925 ( .A(n18805), .B(n18806), .Z(x[380]) );
  NAND U23926 ( .A(creg[380]), .B(init), .Z(n18805) );
  NAND U23927 ( .A(n18807), .B(n18808), .Z(x[37]) );
  NAND U23928 ( .A(creg[37]), .B(init), .Z(n18807) );
  NAND U23929 ( .A(n18809), .B(n18810), .Z(x[379]) );
  NAND U23930 ( .A(creg[379]), .B(init), .Z(n18809) );
  NAND U23931 ( .A(n18811), .B(n18812), .Z(x[378]) );
  NAND U23932 ( .A(creg[378]), .B(init), .Z(n18811) );
  NAND U23933 ( .A(n18813), .B(n18814), .Z(x[377]) );
  NAND U23934 ( .A(creg[377]), .B(init), .Z(n18813) );
  NAND U23935 ( .A(n18815), .B(n18816), .Z(x[376]) );
  NAND U23936 ( .A(creg[376]), .B(init), .Z(n18815) );
  NAND U23937 ( .A(n18817), .B(n18818), .Z(x[375]) );
  NAND U23938 ( .A(creg[375]), .B(init), .Z(n18817) );
  NAND U23939 ( .A(n18819), .B(n18820), .Z(x[374]) );
  NAND U23940 ( .A(creg[374]), .B(init), .Z(n18819) );
  NAND U23941 ( .A(n18821), .B(n18822), .Z(x[373]) );
  NAND U23942 ( .A(creg[373]), .B(init), .Z(n18821) );
  NAND U23943 ( .A(n18823), .B(n18824), .Z(x[372]) );
  NAND U23944 ( .A(creg[372]), .B(init), .Z(n18823) );
  NAND U23945 ( .A(n18825), .B(n18826), .Z(x[371]) );
  NAND U23946 ( .A(creg[371]), .B(init), .Z(n18825) );
  NAND U23947 ( .A(n18827), .B(n18828), .Z(x[370]) );
  NAND U23948 ( .A(creg[370]), .B(init), .Z(n18827) );
  NAND U23949 ( .A(n18829), .B(n18830), .Z(x[36]) );
  NAND U23950 ( .A(creg[36]), .B(init), .Z(n18829) );
  NAND U23951 ( .A(n18831), .B(n18832), .Z(x[369]) );
  NAND U23952 ( .A(creg[369]), .B(init), .Z(n18831) );
  NAND U23953 ( .A(n18833), .B(n18834), .Z(x[368]) );
  NAND U23954 ( .A(creg[368]), .B(init), .Z(n18833) );
  NAND U23955 ( .A(n18835), .B(n18836), .Z(x[367]) );
  NAND U23956 ( .A(creg[367]), .B(init), .Z(n18835) );
  NAND U23957 ( .A(n18837), .B(n18838), .Z(x[366]) );
  NAND U23958 ( .A(creg[366]), .B(init), .Z(n18837) );
  NAND U23959 ( .A(n18839), .B(n18840), .Z(x[365]) );
  NAND U23960 ( .A(creg[365]), .B(init), .Z(n18839) );
  NAND U23961 ( .A(n18841), .B(n18842), .Z(x[364]) );
  NAND U23962 ( .A(creg[364]), .B(init), .Z(n18841) );
  NAND U23963 ( .A(n18843), .B(n18844), .Z(x[363]) );
  NAND U23964 ( .A(creg[363]), .B(init), .Z(n18843) );
  NAND U23965 ( .A(n18845), .B(n18846), .Z(x[362]) );
  NAND U23966 ( .A(creg[362]), .B(init), .Z(n18845) );
  NAND U23967 ( .A(n18847), .B(n18848), .Z(x[361]) );
  NAND U23968 ( .A(creg[361]), .B(init), .Z(n18847) );
  NAND U23969 ( .A(n18849), .B(n18850), .Z(x[360]) );
  NAND U23970 ( .A(creg[360]), .B(init), .Z(n18849) );
  NAND U23971 ( .A(n18851), .B(n18852), .Z(x[35]) );
  NAND U23972 ( .A(creg[35]), .B(init), .Z(n18851) );
  NAND U23973 ( .A(n18853), .B(n18854), .Z(x[359]) );
  NAND U23974 ( .A(creg[359]), .B(init), .Z(n18853) );
  NAND U23975 ( .A(n18855), .B(n18856), .Z(x[358]) );
  NAND U23976 ( .A(creg[358]), .B(init), .Z(n18855) );
  NAND U23977 ( .A(n18857), .B(n18858), .Z(x[357]) );
  NAND U23978 ( .A(creg[357]), .B(init), .Z(n18857) );
  NAND U23979 ( .A(n18859), .B(n18860), .Z(x[356]) );
  NAND U23980 ( .A(creg[356]), .B(init), .Z(n18859) );
  NAND U23981 ( .A(n18861), .B(n18862), .Z(x[355]) );
  NAND U23982 ( .A(creg[355]), .B(init), .Z(n18861) );
  NAND U23983 ( .A(n18863), .B(n18864), .Z(x[354]) );
  NAND U23984 ( .A(creg[354]), .B(init), .Z(n18863) );
  NAND U23985 ( .A(n18865), .B(n18866), .Z(x[353]) );
  NAND U23986 ( .A(creg[353]), .B(init), .Z(n18865) );
  NAND U23987 ( .A(n18867), .B(n18868), .Z(x[352]) );
  NAND U23988 ( .A(creg[352]), .B(init), .Z(n18867) );
  NAND U23989 ( .A(n18869), .B(n18870), .Z(x[351]) );
  NAND U23990 ( .A(creg[351]), .B(init), .Z(n18869) );
  NAND U23991 ( .A(n18871), .B(n18872), .Z(x[350]) );
  NAND U23992 ( .A(creg[350]), .B(init), .Z(n18871) );
  NAND U23993 ( .A(n18873), .B(n18874), .Z(x[34]) );
  NAND U23994 ( .A(creg[34]), .B(init), .Z(n18873) );
  NAND U23995 ( .A(n18875), .B(n18876), .Z(x[349]) );
  NAND U23996 ( .A(creg[349]), .B(init), .Z(n18875) );
  NAND U23997 ( .A(n18877), .B(n18878), .Z(x[348]) );
  NAND U23998 ( .A(creg[348]), .B(init), .Z(n18877) );
  NAND U23999 ( .A(n18879), .B(n18880), .Z(x[347]) );
  NAND U24000 ( .A(creg[347]), .B(init), .Z(n18879) );
  NAND U24001 ( .A(n18881), .B(n18882), .Z(x[346]) );
  NAND U24002 ( .A(creg[346]), .B(init), .Z(n18881) );
  NAND U24003 ( .A(n18883), .B(n18884), .Z(x[345]) );
  NAND U24004 ( .A(creg[345]), .B(init), .Z(n18883) );
  NAND U24005 ( .A(n18885), .B(n18886), .Z(x[344]) );
  NAND U24006 ( .A(creg[344]), .B(init), .Z(n18885) );
  NAND U24007 ( .A(n18887), .B(n18888), .Z(x[343]) );
  NAND U24008 ( .A(creg[343]), .B(init), .Z(n18887) );
  NAND U24009 ( .A(n18889), .B(n18890), .Z(x[342]) );
  NAND U24010 ( .A(creg[342]), .B(init), .Z(n18889) );
  NAND U24011 ( .A(n18891), .B(n18892), .Z(x[341]) );
  NAND U24012 ( .A(creg[341]), .B(init), .Z(n18891) );
  NAND U24013 ( .A(n18893), .B(n18894), .Z(x[340]) );
  NAND U24014 ( .A(creg[340]), .B(init), .Z(n18893) );
  NAND U24015 ( .A(n18895), .B(n18896), .Z(x[33]) );
  NAND U24016 ( .A(creg[33]), .B(init), .Z(n18895) );
  NAND U24017 ( .A(n18897), .B(n18898), .Z(x[339]) );
  NAND U24018 ( .A(creg[339]), .B(init), .Z(n18897) );
  NAND U24019 ( .A(n18899), .B(n18900), .Z(x[338]) );
  NAND U24020 ( .A(creg[338]), .B(init), .Z(n18899) );
  NAND U24021 ( .A(n18901), .B(n18902), .Z(x[337]) );
  NAND U24022 ( .A(creg[337]), .B(init), .Z(n18901) );
  NAND U24023 ( .A(n18903), .B(n18904), .Z(x[336]) );
  NAND U24024 ( .A(creg[336]), .B(init), .Z(n18903) );
  NAND U24025 ( .A(n18905), .B(n18906), .Z(x[335]) );
  NAND U24026 ( .A(creg[335]), .B(init), .Z(n18905) );
  NAND U24027 ( .A(n18907), .B(n18908), .Z(x[334]) );
  NAND U24028 ( .A(creg[334]), .B(init), .Z(n18907) );
  NAND U24029 ( .A(n18909), .B(n18910), .Z(x[333]) );
  NAND U24030 ( .A(creg[333]), .B(init), .Z(n18909) );
  NAND U24031 ( .A(n18911), .B(n18912), .Z(x[332]) );
  NAND U24032 ( .A(creg[332]), .B(init), .Z(n18911) );
  NAND U24033 ( .A(n18913), .B(n18914), .Z(x[331]) );
  NAND U24034 ( .A(creg[331]), .B(init), .Z(n18913) );
  NAND U24035 ( .A(n18915), .B(n18916), .Z(x[330]) );
  NAND U24036 ( .A(creg[330]), .B(init), .Z(n18915) );
  NAND U24037 ( .A(n18917), .B(n18918), .Z(x[32]) );
  NAND U24038 ( .A(creg[32]), .B(init), .Z(n18917) );
  NAND U24039 ( .A(n18919), .B(n18920), .Z(x[329]) );
  NAND U24040 ( .A(creg[329]), .B(init), .Z(n18919) );
  NAND U24041 ( .A(n18921), .B(n18922), .Z(x[328]) );
  NAND U24042 ( .A(creg[328]), .B(init), .Z(n18921) );
  NAND U24043 ( .A(n18923), .B(n18924), .Z(x[327]) );
  NAND U24044 ( .A(creg[327]), .B(init), .Z(n18923) );
  NAND U24045 ( .A(n18925), .B(n18926), .Z(x[326]) );
  NAND U24046 ( .A(creg[326]), .B(init), .Z(n18925) );
  NAND U24047 ( .A(n18927), .B(n18928), .Z(x[325]) );
  NAND U24048 ( .A(creg[325]), .B(init), .Z(n18927) );
  NAND U24049 ( .A(n18929), .B(n18930), .Z(x[324]) );
  NAND U24050 ( .A(creg[324]), .B(init), .Z(n18929) );
  NAND U24051 ( .A(n18931), .B(n18932), .Z(x[323]) );
  NAND U24052 ( .A(creg[323]), .B(init), .Z(n18931) );
  NAND U24053 ( .A(n18933), .B(n18934), .Z(x[322]) );
  NAND U24054 ( .A(creg[322]), .B(init), .Z(n18933) );
  NAND U24055 ( .A(n18935), .B(n18936), .Z(x[321]) );
  NAND U24056 ( .A(creg[321]), .B(init), .Z(n18935) );
  NAND U24057 ( .A(n18937), .B(n18938), .Z(x[320]) );
  NAND U24058 ( .A(creg[320]), .B(init), .Z(n18937) );
  NAND U24059 ( .A(n18939), .B(n18940), .Z(x[31]) );
  NAND U24060 ( .A(creg[31]), .B(init), .Z(n18939) );
  NAND U24061 ( .A(n18941), .B(n18942), .Z(x[319]) );
  NAND U24062 ( .A(creg[319]), .B(init), .Z(n18941) );
  NAND U24063 ( .A(n18943), .B(n18944), .Z(x[318]) );
  NAND U24064 ( .A(creg[318]), .B(init), .Z(n18943) );
  NAND U24065 ( .A(n18945), .B(n18946), .Z(x[317]) );
  NAND U24066 ( .A(creg[317]), .B(init), .Z(n18945) );
  NAND U24067 ( .A(n18947), .B(n18948), .Z(x[316]) );
  NAND U24068 ( .A(creg[316]), .B(init), .Z(n18947) );
  NAND U24069 ( .A(n18949), .B(n18950), .Z(x[315]) );
  NAND U24070 ( .A(creg[315]), .B(init), .Z(n18949) );
  NAND U24071 ( .A(n18951), .B(n18952), .Z(x[314]) );
  NAND U24072 ( .A(creg[314]), .B(init), .Z(n18951) );
  NAND U24073 ( .A(n18953), .B(n18954), .Z(x[313]) );
  NAND U24074 ( .A(creg[313]), .B(init), .Z(n18953) );
  NAND U24075 ( .A(n18955), .B(n18956), .Z(x[312]) );
  NAND U24076 ( .A(creg[312]), .B(init), .Z(n18955) );
  NAND U24077 ( .A(n18957), .B(n18958), .Z(x[311]) );
  NAND U24078 ( .A(creg[311]), .B(init), .Z(n18957) );
  NAND U24079 ( .A(n18959), .B(n18960), .Z(x[310]) );
  NAND U24080 ( .A(creg[310]), .B(init), .Z(n18959) );
  NAND U24081 ( .A(n18961), .B(n18962), .Z(x[30]) );
  NAND U24082 ( .A(creg[30]), .B(init), .Z(n18961) );
  NAND U24083 ( .A(n18963), .B(n18964), .Z(x[309]) );
  NAND U24084 ( .A(creg[309]), .B(init), .Z(n18963) );
  NAND U24085 ( .A(n18965), .B(n18966), .Z(x[308]) );
  NAND U24086 ( .A(creg[308]), .B(init), .Z(n18965) );
  NAND U24087 ( .A(n18967), .B(n18968), .Z(x[307]) );
  NAND U24088 ( .A(creg[307]), .B(init), .Z(n18967) );
  NAND U24089 ( .A(n18969), .B(n18970), .Z(x[306]) );
  NAND U24090 ( .A(creg[306]), .B(init), .Z(n18969) );
  NAND U24091 ( .A(n18971), .B(n18972), .Z(x[305]) );
  NAND U24092 ( .A(creg[305]), .B(init), .Z(n18971) );
  NAND U24093 ( .A(n18973), .B(n18974), .Z(x[304]) );
  NAND U24094 ( .A(creg[304]), .B(init), .Z(n18973) );
  NAND U24095 ( .A(n18975), .B(n18976), .Z(x[303]) );
  NAND U24096 ( .A(creg[303]), .B(init), .Z(n18975) );
  NAND U24097 ( .A(n18977), .B(n18978), .Z(x[302]) );
  NAND U24098 ( .A(creg[302]), .B(init), .Z(n18977) );
  NAND U24099 ( .A(n18979), .B(n18980), .Z(x[301]) );
  NAND U24100 ( .A(creg[301]), .B(init), .Z(n18979) );
  NAND U24101 ( .A(n18981), .B(n18982), .Z(x[300]) );
  NAND U24102 ( .A(creg[300]), .B(init), .Z(n18981) );
  NAND U24103 ( .A(n18983), .B(n18984), .Z(x[2]) );
  NAND U24104 ( .A(creg[2]), .B(init), .Z(n18983) );
  NAND U24105 ( .A(n18985), .B(n18986), .Z(x[29]) );
  NAND U24106 ( .A(creg[29]), .B(init), .Z(n18985) );
  NAND U24107 ( .A(n18987), .B(n18988), .Z(x[299]) );
  NAND U24108 ( .A(creg[299]), .B(init), .Z(n18987) );
  NAND U24109 ( .A(n18989), .B(n18990), .Z(x[298]) );
  NAND U24110 ( .A(creg[298]), .B(init), .Z(n18989) );
  NAND U24111 ( .A(n18991), .B(n18992), .Z(x[297]) );
  NAND U24112 ( .A(creg[297]), .B(init), .Z(n18991) );
  NAND U24113 ( .A(n18993), .B(n18994), .Z(x[296]) );
  NAND U24114 ( .A(creg[296]), .B(init), .Z(n18993) );
  NAND U24115 ( .A(n18995), .B(n18996), .Z(x[295]) );
  NAND U24116 ( .A(creg[295]), .B(init), .Z(n18995) );
  NAND U24117 ( .A(n18997), .B(n18998), .Z(x[294]) );
  NAND U24118 ( .A(creg[294]), .B(init), .Z(n18997) );
  NAND U24119 ( .A(n18999), .B(n19000), .Z(x[293]) );
  NAND U24120 ( .A(creg[293]), .B(init), .Z(n18999) );
  NAND U24121 ( .A(n19001), .B(n19002), .Z(x[292]) );
  NAND U24122 ( .A(creg[292]), .B(init), .Z(n19001) );
  NAND U24123 ( .A(n19003), .B(n19004), .Z(x[291]) );
  NAND U24124 ( .A(creg[291]), .B(init), .Z(n19003) );
  NAND U24125 ( .A(n19005), .B(n19006), .Z(x[290]) );
  NAND U24126 ( .A(creg[290]), .B(init), .Z(n19005) );
  NAND U24127 ( .A(n19007), .B(n19008), .Z(x[28]) );
  NAND U24128 ( .A(creg[28]), .B(init), .Z(n19007) );
  NAND U24129 ( .A(n19009), .B(n19010), .Z(x[289]) );
  NAND U24130 ( .A(creg[289]), .B(init), .Z(n19009) );
  NAND U24131 ( .A(n19011), .B(n19012), .Z(x[288]) );
  NAND U24132 ( .A(creg[288]), .B(init), .Z(n19011) );
  NAND U24133 ( .A(n19013), .B(n19014), .Z(x[287]) );
  NAND U24134 ( .A(creg[287]), .B(init), .Z(n19013) );
  NAND U24135 ( .A(n19015), .B(n19016), .Z(x[286]) );
  NAND U24136 ( .A(creg[286]), .B(init), .Z(n19015) );
  NAND U24137 ( .A(n19017), .B(n19018), .Z(x[285]) );
  NAND U24138 ( .A(creg[285]), .B(init), .Z(n19017) );
  NAND U24139 ( .A(n19019), .B(n19020), .Z(x[284]) );
  NAND U24140 ( .A(creg[284]), .B(init), .Z(n19019) );
  NAND U24141 ( .A(n19021), .B(n19022), .Z(x[283]) );
  NAND U24142 ( .A(creg[283]), .B(init), .Z(n19021) );
  NAND U24143 ( .A(n19023), .B(n19024), .Z(x[282]) );
  NAND U24144 ( .A(creg[282]), .B(init), .Z(n19023) );
  NAND U24145 ( .A(n19025), .B(n19026), .Z(x[281]) );
  NAND U24146 ( .A(creg[281]), .B(init), .Z(n19025) );
  NAND U24147 ( .A(n19027), .B(n19028), .Z(x[280]) );
  NAND U24148 ( .A(creg[280]), .B(init), .Z(n19027) );
  NAND U24149 ( .A(n19029), .B(n19030), .Z(x[27]) );
  NAND U24150 ( .A(creg[27]), .B(init), .Z(n19029) );
  NAND U24151 ( .A(n19031), .B(n19032), .Z(x[279]) );
  NAND U24152 ( .A(creg[279]), .B(init), .Z(n19031) );
  NAND U24153 ( .A(n19033), .B(n19034), .Z(x[278]) );
  NAND U24154 ( .A(creg[278]), .B(init), .Z(n19033) );
  NAND U24155 ( .A(n19035), .B(n19036), .Z(x[277]) );
  NAND U24156 ( .A(creg[277]), .B(init), .Z(n19035) );
  NAND U24157 ( .A(n19037), .B(n19038), .Z(x[276]) );
  NAND U24158 ( .A(creg[276]), .B(init), .Z(n19037) );
  NAND U24159 ( .A(n19039), .B(n19040), .Z(x[275]) );
  NAND U24160 ( .A(creg[275]), .B(init), .Z(n19039) );
  NAND U24161 ( .A(n19041), .B(n19042), .Z(x[274]) );
  NAND U24162 ( .A(creg[274]), .B(init), .Z(n19041) );
  NAND U24163 ( .A(n19043), .B(n19044), .Z(x[273]) );
  NAND U24164 ( .A(creg[273]), .B(init), .Z(n19043) );
  NAND U24165 ( .A(n19045), .B(n19046), .Z(x[272]) );
  NAND U24166 ( .A(creg[272]), .B(init), .Z(n19045) );
  NAND U24167 ( .A(n19047), .B(n19048), .Z(x[271]) );
  NAND U24168 ( .A(creg[271]), .B(init), .Z(n19047) );
  NAND U24169 ( .A(n19049), .B(n19050), .Z(x[270]) );
  NAND U24170 ( .A(creg[270]), .B(init), .Z(n19049) );
  NAND U24171 ( .A(n19051), .B(n19052), .Z(x[26]) );
  NAND U24172 ( .A(creg[26]), .B(init), .Z(n19051) );
  NAND U24173 ( .A(n19053), .B(n19054), .Z(x[269]) );
  NAND U24174 ( .A(creg[269]), .B(init), .Z(n19053) );
  NAND U24175 ( .A(n19055), .B(n19056), .Z(x[268]) );
  NAND U24176 ( .A(creg[268]), .B(init), .Z(n19055) );
  NAND U24177 ( .A(n19057), .B(n19058), .Z(x[267]) );
  NAND U24178 ( .A(creg[267]), .B(init), .Z(n19057) );
  NAND U24179 ( .A(n19059), .B(n19060), .Z(x[266]) );
  NAND U24180 ( .A(creg[266]), .B(init), .Z(n19059) );
  NAND U24181 ( .A(n19061), .B(n19062), .Z(x[265]) );
  NAND U24182 ( .A(creg[265]), .B(init), .Z(n19061) );
  NAND U24183 ( .A(n19063), .B(n19064), .Z(x[264]) );
  NAND U24184 ( .A(creg[264]), .B(init), .Z(n19063) );
  NAND U24185 ( .A(n19065), .B(n19066), .Z(x[263]) );
  NAND U24186 ( .A(creg[263]), .B(init), .Z(n19065) );
  NAND U24187 ( .A(n19067), .B(n19068), .Z(x[262]) );
  NAND U24188 ( .A(creg[262]), .B(init), .Z(n19067) );
  NAND U24189 ( .A(n19069), .B(n19070), .Z(x[261]) );
  NAND U24190 ( .A(creg[261]), .B(init), .Z(n19069) );
  NAND U24191 ( .A(n19071), .B(n19072), .Z(x[260]) );
  NAND U24192 ( .A(creg[260]), .B(init), .Z(n19071) );
  NAND U24193 ( .A(n19073), .B(n19074), .Z(x[25]) );
  NAND U24194 ( .A(creg[25]), .B(init), .Z(n19073) );
  NAND U24195 ( .A(n19075), .B(n19076), .Z(x[259]) );
  NAND U24196 ( .A(creg[259]), .B(init), .Z(n19075) );
  NAND U24197 ( .A(n19077), .B(n19078), .Z(x[258]) );
  NAND U24198 ( .A(creg[258]), .B(init), .Z(n19077) );
  NAND U24199 ( .A(n19079), .B(n19080), .Z(x[257]) );
  NAND U24200 ( .A(creg[257]), .B(init), .Z(n19079) );
  NAND U24201 ( .A(n19081), .B(n19082), .Z(x[256]) );
  NAND U24202 ( .A(creg[256]), .B(init), .Z(n19081) );
  NAND U24203 ( .A(n19083), .B(n19084), .Z(x[255]) );
  NAND U24204 ( .A(creg[255]), .B(init), .Z(n19083) );
  NAND U24205 ( .A(n19085), .B(n19086), .Z(x[254]) );
  NAND U24206 ( .A(creg[254]), .B(init), .Z(n19085) );
  NAND U24207 ( .A(n19087), .B(n19088), .Z(x[253]) );
  NAND U24208 ( .A(creg[253]), .B(init), .Z(n19087) );
  NAND U24209 ( .A(n19089), .B(n19090), .Z(x[252]) );
  NAND U24210 ( .A(creg[252]), .B(init), .Z(n19089) );
  NAND U24211 ( .A(n19091), .B(n19092), .Z(x[251]) );
  NAND U24212 ( .A(creg[251]), .B(init), .Z(n19091) );
  NAND U24213 ( .A(n19093), .B(n19094), .Z(x[250]) );
  NAND U24214 ( .A(creg[250]), .B(init), .Z(n19093) );
  NAND U24215 ( .A(n19095), .B(n19096), .Z(x[24]) );
  NAND U24216 ( .A(creg[24]), .B(init), .Z(n19095) );
  NAND U24217 ( .A(n19097), .B(n19098), .Z(x[249]) );
  NAND U24218 ( .A(creg[249]), .B(init), .Z(n19097) );
  NAND U24219 ( .A(n19099), .B(n19100), .Z(x[248]) );
  NAND U24220 ( .A(creg[248]), .B(init), .Z(n19099) );
  NAND U24221 ( .A(n19101), .B(n19102), .Z(x[247]) );
  NAND U24222 ( .A(creg[247]), .B(init), .Z(n19101) );
  NAND U24223 ( .A(n19103), .B(n19104), .Z(x[246]) );
  NAND U24224 ( .A(creg[246]), .B(init), .Z(n19103) );
  NAND U24225 ( .A(n19105), .B(n19106), .Z(x[245]) );
  NAND U24226 ( .A(creg[245]), .B(init), .Z(n19105) );
  NAND U24227 ( .A(n19107), .B(n19108), .Z(x[244]) );
  NAND U24228 ( .A(creg[244]), .B(init), .Z(n19107) );
  NAND U24229 ( .A(n19109), .B(n19110), .Z(x[243]) );
  NAND U24230 ( .A(creg[243]), .B(init), .Z(n19109) );
  NAND U24231 ( .A(n19111), .B(n19112), .Z(x[242]) );
  NAND U24232 ( .A(creg[242]), .B(init), .Z(n19111) );
  NAND U24233 ( .A(n19113), .B(n19114), .Z(x[241]) );
  NAND U24234 ( .A(creg[241]), .B(init), .Z(n19113) );
  NAND U24235 ( .A(n19115), .B(n19116), .Z(x[240]) );
  NAND U24236 ( .A(creg[240]), .B(init), .Z(n19115) );
  NAND U24237 ( .A(n19117), .B(n19118), .Z(x[23]) );
  NAND U24238 ( .A(creg[23]), .B(init), .Z(n19117) );
  NAND U24239 ( .A(n19119), .B(n19120), .Z(x[239]) );
  NAND U24240 ( .A(creg[239]), .B(init), .Z(n19119) );
  NAND U24241 ( .A(n19121), .B(n19122), .Z(x[238]) );
  NAND U24242 ( .A(creg[238]), .B(init), .Z(n19121) );
  NAND U24243 ( .A(n19123), .B(n19124), .Z(x[237]) );
  NAND U24244 ( .A(creg[237]), .B(init), .Z(n19123) );
  NAND U24245 ( .A(n19125), .B(n19126), .Z(x[236]) );
  NAND U24246 ( .A(creg[236]), .B(init), .Z(n19125) );
  NAND U24247 ( .A(n19127), .B(n19128), .Z(x[235]) );
  NAND U24248 ( .A(creg[235]), .B(init), .Z(n19127) );
  NAND U24249 ( .A(n19129), .B(n19130), .Z(x[234]) );
  NAND U24250 ( .A(creg[234]), .B(init), .Z(n19129) );
  NAND U24251 ( .A(n19131), .B(n19132), .Z(x[233]) );
  NAND U24252 ( .A(creg[233]), .B(init), .Z(n19131) );
  NAND U24253 ( .A(n19133), .B(n19134), .Z(x[232]) );
  NAND U24254 ( .A(creg[232]), .B(init), .Z(n19133) );
  NAND U24255 ( .A(n19135), .B(n19136), .Z(x[231]) );
  NAND U24256 ( .A(creg[231]), .B(init), .Z(n19135) );
  NAND U24257 ( .A(n19137), .B(n19138), .Z(x[230]) );
  NAND U24258 ( .A(creg[230]), .B(init), .Z(n19137) );
  NAND U24259 ( .A(n19139), .B(n19140), .Z(x[22]) );
  NAND U24260 ( .A(creg[22]), .B(init), .Z(n19139) );
  NAND U24261 ( .A(n19141), .B(n19142), .Z(x[229]) );
  NAND U24262 ( .A(creg[229]), .B(init), .Z(n19141) );
  NAND U24263 ( .A(n19143), .B(n19144), .Z(x[228]) );
  NAND U24264 ( .A(creg[228]), .B(init), .Z(n19143) );
  NAND U24265 ( .A(n19145), .B(n19146), .Z(x[227]) );
  NAND U24266 ( .A(creg[227]), .B(init), .Z(n19145) );
  NAND U24267 ( .A(n19147), .B(n19148), .Z(x[226]) );
  NAND U24268 ( .A(creg[226]), .B(init), .Z(n19147) );
  NAND U24269 ( .A(n19149), .B(n19150), .Z(x[225]) );
  NAND U24270 ( .A(creg[225]), .B(init), .Z(n19149) );
  NAND U24271 ( .A(n19151), .B(n19152), .Z(x[224]) );
  NAND U24272 ( .A(creg[224]), .B(init), .Z(n19151) );
  NAND U24273 ( .A(n19153), .B(n19154), .Z(x[223]) );
  NAND U24274 ( .A(creg[223]), .B(init), .Z(n19153) );
  NAND U24275 ( .A(n19155), .B(n19156), .Z(x[222]) );
  NAND U24276 ( .A(creg[222]), .B(init), .Z(n19155) );
  NAND U24277 ( .A(n19157), .B(n19158), .Z(x[221]) );
  NAND U24278 ( .A(creg[221]), .B(init), .Z(n19157) );
  NAND U24279 ( .A(n19159), .B(n19160), .Z(x[220]) );
  NAND U24280 ( .A(creg[220]), .B(init), .Z(n19159) );
  NAND U24281 ( .A(n19161), .B(n19162), .Z(x[21]) );
  NAND U24282 ( .A(creg[21]), .B(init), .Z(n19161) );
  NAND U24283 ( .A(n19163), .B(n19164), .Z(x[219]) );
  NAND U24284 ( .A(creg[219]), .B(init), .Z(n19163) );
  NAND U24285 ( .A(n19165), .B(n19166), .Z(x[218]) );
  NAND U24286 ( .A(creg[218]), .B(init), .Z(n19165) );
  NAND U24287 ( .A(n19167), .B(n19168), .Z(x[217]) );
  NAND U24288 ( .A(creg[217]), .B(init), .Z(n19167) );
  NAND U24289 ( .A(n19169), .B(n19170), .Z(x[216]) );
  NAND U24290 ( .A(creg[216]), .B(init), .Z(n19169) );
  NAND U24291 ( .A(n19171), .B(n19172), .Z(x[215]) );
  NAND U24292 ( .A(creg[215]), .B(init), .Z(n19171) );
  NAND U24293 ( .A(n19173), .B(n19174), .Z(x[214]) );
  NAND U24294 ( .A(creg[214]), .B(init), .Z(n19173) );
  NAND U24295 ( .A(n19175), .B(n19176), .Z(x[213]) );
  NAND U24296 ( .A(creg[213]), .B(init), .Z(n19175) );
  NAND U24297 ( .A(n19177), .B(n19178), .Z(x[212]) );
  NAND U24298 ( .A(creg[212]), .B(init), .Z(n19177) );
  NAND U24299 ( .A(n19179), .B(n19180), .Z(x[211]) );
  NAND U24300 ( .A(creg[211]), .B(init), .Z(n19179) );
  NAND U24301 ( .A(n19181), .B(n19182), .Z(x[210]) );
  NAND U24302 ( .A(creg[210]), .B(init), .Z(n19181) );
  NAND U24303 ( .A(n19183), .B(n19184), .Z(x[20]) );
  NAND U24304 ( .A(creg[20]), .B(init), .Z(n19183) );
  NAND U24305 ( .A(n19185), .B(n19186), .Z(x[209]) );
  NAND U24306 ( .A(creg[209]), .B(init), .Z(n19185) );
  NAND U24307 ( .A(n19187), .B(n19188), .Z(x[208]) );
  NAND U24308 ( .A(creg[208]), .B(init), .Z(n19187) );
  NAND U24309 ( .A(n19189), .B(n19190), .Z(x[207]) );
  NAND U24310 ( .A(creg[207]), .B(init), .Z(n19189) );
  NAND U24311 ( .A(n19191), .B(n19192), .Z(x[206]) );
  NAND U24312 ( .A(creg[206]), .B(init), .Z(n19191) );
  NAND U24313 ( .A(n19193), .B(n19194), .Z(x[205]) );
  NAND U24314 ( .A(creg[205]), .B(init), .Z(n19193) );
  NAND U24315 ( .A(n19195), .B(n19196), .Z(x[204]) );
  NAND U24316 ( .A(creg[204]), .B(init), .Z(n19195) );
  NAND U24317 ( .A(n19197), .B(n19198), .Z(x[203]) );
  NAND U24318 ( .A(creg[203]), .B(init), .Z(n19197) );
  NAND U24319 ( .A(n19199), .B(n19200), .Z(x[202]) );
  NAND U24320 ( .A(creg[202]), .B(init), .Z(n19199) );
  NAND U24321 ( .A(n19201), .B(n19202), .Z(x[201]) );
  NAND U24322 ( .A(creg[201]), .B(init), .Z(n19201) );
  NAND U24323 ( .A(n19203), .B(n19204), .Z(x[200]) );
  NAND U24324 ( .A(creg[200]), .B(init), .Z(n19203) );
  NAND U24325 ( .A(n19205), .B(n19206), .Z(x[1]) );
  NAND U24326 ( .A(creg[1]), .B(init), .Z(n19205) );
  NAND U24327 ( .A(n19207), .B(n19208), .Z(x[19]) );
  NAND U24328 ( .A(creg[19]), .B(init), .Z(n19207) );
  NAND U24329 ( .A(n19209), .B(n19210), .Z(x[199]) );
  NAND U24330 ( .A(creg[199]), .B(init), .Z(n19209) );
  NAND U24331 ( .A(n19211), .B(n19212), .Z(x[198]) );
  NAND U24332 ( .A(creg[198]), .B(init), .Z(n19211) );
  NAND U24333 ( .A(n19213), .B(n19214), .Z(x[197]) );
  NAND U24334 ( .A(creg[197]), .B(init), .Z(n19213) );
  NAND U24335 ( .A(n19215), .B(n19216), .Z(x[196]) );
  NAND U24336 ( .A(creg[196]), .B(init), .Z(n19215) );
  NAND U24337 ( .A(n19217), .B(n19218), .Z(x[195]) );
  NAND U24338 ( .A(creg[195]), .B(init), .Z(n19217) );
  NAND U24339 ( .A(n19219), .B(n19220), .Z(x[194]) );
  NAND U24340 ( .A(creg[194]), .B(init), .Z(n19219) );
  NAND U24341 ( .A(n19221), .B(n19222), .Z(x[193]) );
  NAND U24342 ( .A(creg[193]), .B(init), .Z(n19221) );
  NAND U24343 ( .A(n19223), .B(n19224), .Z(x[192]) );
  NAND U24344 ( .A(creg[192]), .B(init), .Z(n19223) );
  NAND U24345 ( .A(n19225), .B(n19226), .Z(x[191]) );
  NAND U24346 ( .A(creg[191]), .B(init), .Z(n19225) );
  NAND U24347 ( .A(n19227), .B(n19228), .Z(x[190]) );
  NAND U24348 ( .A(creg[190]), .B(init), .Z(n19227) );
  NAND U24349 ( .A(n19229), .B(n19230), .Z(x[18]) );
  NAND U24350 ( .A(creg[18]), .B(init), .Z(n19229) );
  NAND U24351 ( .A(n19231), .B(n19232), .Z(x[189]) );
  NAND U24352 ( .A(creg[189]), .B(init), .Z(n19231) );
  NAND U24353 ( .A(n19233), .B(n19234), .Z(x[188]) );
  NAND U24354 ( .A(creg[188]), .B(init), .Z(n19233) );
  NAND U24355 ( .A(n19235), .B(n19236), .Z(x[187]) );
  NAND U24356 ( .A(creg[187]), .B(init), .Z(n19235) );
  NAND U24357 ( .A(n19237), .B(n19238), .Z(x[186]) );
  NAND U24358 ( .A(creg[186]), .B(init), .Z(n19237) );
  NAND U24359 ( .A(n19239), .B(n19240), .Z(x[185]) );
  NAND U24360 ( .A(creg[185]), .B(init), .Z(n19239) );
  NAND U24361 ( .A(n19241), .B(n19242), .Z(x[184]) );
  NAND U24362 ( .A(creg[184]), .B(init), .Z(n19241) );
  NAND U24363 ( .A(n19243), .B(n19244), .Z(x[183]) );
  NAND U24364 ( .A(creg[183]), .B(init), .Z(n19243) );
  NAND U24365 ( .A(n19245), .B(n19246), .Z(x[182]) );
  NAND U24366 ( .A(creg[182]), .B(init), .Z(n19245) );
  NAND U24367 ( .A(n19247), .B(n19248), .Z(x[181]) );
  NAND U24368 ( .A(creg[181]), .B(init), .Z(n19247) );
  NAND U24369 ( .A(n19249), .B(n19250), .Z(x[180]) );
  NAND U24370 ( .A(creg[180]), .B(init), .Z(n19249) );
  NAND U24371 ( .A(n19251), .B(n19252), .Z(x[17]) );
  NAND U24372 ( .A(creg[17]), .B(init), .Z(n19251) );
  NAND U24373 ( .A(n19253), .B(n19254), .Z(x[179]) );
  NAND U24374 ( .A(creg[179]), .B(init), .Z(n19253) );
  NAND U24375 ( .A(n19255), .B(n19256), .Z(x[178]) );
  NAND U24376 ( .A(creg[178]), .B(init), .Z(n19255) );
  NAND U24377 ( .A(n19257), .B(n19258), .Z(x[177]) );
  NAND U24378 ( .A(creg[177]), .B(init), .Z(n19257) );
  NAND U24379 ( .A(n19259), .B(n19260), .Z(x[176]) );
  NAND U24380 ( .A(creg[176]), .B(init), .Z(n19259) );
  NAND U24381 ( .A(n19261), .B(n19262), .Z(x[175]) );
  NAND U24382 ( .A(creg[175]), .B(init), .Z(n19261) );
  NAND U24383 ( .A(n19263), .B(n19264), .Z(x[174]) );
  NAND U24384 ( .A(creg[174]), .B(init), .Z(n19263) );
  NAND U24385 ( .A(n19265), .B(n19266), .Z(x[173]) );
  NAND U24386 ( .A(creg[173]), .B(init), .Z(n19265) );
  NAND U24387 ( .A(n19267), .B(n19268), .Z(x[172]) );
  NAND U24388 ( .A(creg[172]), .B(init), .Z(n19267) );
  NAND U24389 ( .A(n19269), .B(n19270), .Z(x[171]) );
  NAND U24390 ( .A(creg[171]), .B(init), .Z(n19269) );
  NAND U24391 ( .A(n19271), .B(n19272), .Z(x[170]) );
  NAND U24392 ( .A(creg[170]), .B(init), .Z(n19271) );
  NAND U24393 ( .A(n19273), .B(n19274), .Z(x[16]) );
  NAND U24394 ( .A(creg[16]), .B(init), .Z(n19273) );
  NAND U24395 ( .A(n19275), .B(n19276), .Z(x[169]) );
  NAND U24396 ( .A(creg[169]), .B(init), .Z(n19275) );
  NAND U24397 ( .A(n19277), .B(n19278), .Z(x[168]) );
  NAND U24398 ( .A(creg[168]), .B(init), .Z(n19277) );
  NAND U24399 ( .A(n19279), .B(n19280), .Z(x[167]) );
  NAND U24400 ( .A(creg[167]), .B(init), .Z(n19279) );
  NAND U24401 ( .A(n19281), .B(n19282), .Z(x[166]) );
  NAND U24402 ( .A(creg[166]), .B(init), .Z(n19281) );
  NAND U24403 ( .A(n19283), .B(n19284), .Z(x[165]) );
  NAND U24404 ( .A(creg[165]), .B(init), .Z(n19283) );
  NAND U24405 ( .A(n19285), .B(n19286), .Z(x[164]) );
  NAND U24406 ( .A(creg[164]), .B(init), .Z(n19285) );
  NAND U24407 ( .A(n19287), .B(n19288), .Z(x[163]) );
  NAND U24408 ( .A(creg[163]), .B(init), .Z(n19287) );
  NAND U24409 ( .A(n19289), .B(n19290), .Z(x[162]) );
  NAND U24410 ( .A(creg[162]), .B(init), .Z(n19289) );
  NAND U24411 ( .A(n19291), .B(n19292), .Z(x[161]) );
  NAND U24412 ( .A(creg[161]), .B(init), .Z(n19291) );
  NAND U24413 ( .A(n19293), .B(n19294), .Z(x[160]) );
  NAND U24414 ( .A(creg[160]), .B(init), .Z(n19293) );
  NAND U24415 ( .A(n19295), .B(n19296), .Z(x[15]) );
  NAND U24416 ( .A(creg[15]), .B(init), .Z(n19295) );
  NAND U24417 ( .A(n19297), .B(n19298), .Z(x[159]) );
  NAND U24418 ( .A(creg[159]), .B(init), .Z(n19297) );
  NAND U24419 ( .A(n19299), .B(n19300), .Z(x[158]) );
  NAND U24420 ( .A(creg[158]), .B(init), .Z(n19299) );
  NAND U24421 ( .A(n19301), .B(n19302), .Z(x[157]) );
  NAND U24422 ( .A(creg[157]), .B(init), .Z(n19301) );
  NAND U24423 ( .A(n19303), .B(n19304), .Z(x[156]) );
  NAND U24424 ( .A(creg[156]), .B(init), .Z(n19303) );
  NAND U24425 ( .A(n19305), .B(n19306), .Z(x[155]) );
  NAND U24426 ( .A(creg[155]), .B(init), .Z(n19305) );
  NAND U24427 ( .A(n19307), .B(n19308), .Z(x[154]) );
  NAND U24428 ( .A(creg[154]), .B(init), .Z(n19307) );
  NAND U24429 ( .A(n19309), .B(n19310), .Z(x[153]) );
  NAND U24430 ( .A(creg[153]), .B(init), .Z(n19309) );
  NAND U24431 ( .A(n19311), .B(n19312), .Z(x[152]) );
  NAND U24432 ( .A(creg[152]), .B(init), .Z(n19311) );
  NAND U24433 ( .A(n19313), .B(n19314), .Z(x[151]) );
  NAND U24434 ( .A(creg[151]), .B(init), .Z(n19313) );
  NAND U24435 ( .A(n19315), .B(n19316), .Z(x[150]) );
  NAND U24436 ( .A(creg[150]), .B(init), .Z(n19315) );
  NAND U24437 ( .A(n19317), .B(n19318), .Z(x[14]) );
  NAND U24438 ( .A(creg[14]), .B(init), .Z(n19317) );
  NAND U24439 ( .A(n19319), .B(n19320), .Z(x[149]) );
  NAND U24440 ( .A(creg[149]), .B(init), .Z(n19319) );
  NAND U24441 ( .A(n19321), .B(n19322), .Z(x[148]) );
  NAND U24442 ( .A(creg[148]), .B(init), .Z(n19321) );
  NAND U24443 ( .A(n19323), .B(n19324), .Z(x[147]) );
  NAND U24444 ( .A(creg[147]), .B(init), .Z(n19323) );
  NAND U24445 ( .A(n19325), .B(n19326), .Z(x[146]) );
  NAND U24446 ( .A(creg[146]), .B(init), .Z(n19325) );
  NAND U24447 ( .A(n19327), .B(n19328), .Z(x[145]) );
  NAND U24448 ( .A(creg[145]), .B(init), .Z(n19327) );
  NAND U24449 ( .A(n19329), .B(n19330), .Z(x[144]) );
  NAND U24450 ( .A(creg[144]), .B(init), .Z(n19329) );
  NAND U24451 ( .A(n19331), .B(n19332), .Z(x[143]) );
  NAND U24452 ( .A(creg[143]), .B(init), .Z(n19331) );
  NAND U24453 ( .A(n19333), .B(n19334), .Z(x[142]) );
  NAND U24454 ( .A(creg[142]), .B(init), .Z(n19333) );
  NAND U24455 ( .A(n19335), .B(n19336), .Z(x[141]) );
  NAND U24456 ( .A(creg[141]), .B(init), .Z(n19335) );
  NAND U24457 ( .A(n19337), .B(n19338), .Z(x[140]) );
  NAND U24458 ( .A(creg[140]), .B(init), .Z(n19337) );
  NAND U24459 ( .A(n19339), .B(n19340), .Z(x[13]) );
  NAND U24460 ( .A(creg[13]), .B(init), .Z(n19339) );
  NAND U24461 ( .A(n19341), .B(n19342), .Z(x[139]) );
  NAND U24462 ( .A(creg[139]), .B(init), .Z(n19341) );
  NAND U24463 ( .A(n19343), .B(n19344), .Z(x[138]) );
  NAND U24464 ( .A(creg[138]), .B(init), .Z(n19343) );
  NAND U24465 ( .A(n19345), .B(n19346), .Z(x[137]) );
  NAND U24466 ( .A(creg[137]), .B(init), .Z(n19345) );
  NAND U24467 ( .A(n19347), .B(n19348), .Z(x[136]) );
  NAND U24468 ( .A(creg[136]), .B(init), .Z(n19347) );
  NAND U24469 ( .A(n19349), .B(n19350), .Z(x[135]) );
  NAND U24470 ( .A(creg[135]), .B(init), .Z(n19349) );
  NAND U24471 ( .A(n19351), .B(n19352), .Z(x[134]) );
  NAND U24472 ( .A(creg[134]), .B(init), .Z(n19351) );
  NAND U24473 ( .A(n19353), .B(n19354), .Z(x[133]) );
  NAND U24474 ( .A(creg[133]), .B(init), .Z(n19353) );
  NAND U24475 ( .A(n19355), .B(n19356), .Z(x[132]) );
  NAND U24476 ( .A(creg[132]), .B(init), .Z(n19355) );
  NAND U24477 ( .A(n19357), .B(n19358), .Z(x[131]) );
  NAND U24478 ( .A(creg[131]), .B(init), .Z(n19357) );
  NAND U24479 ( .A(n19359), .B(n19360), .Z(x[130]) );
  NAND U24480 ( .A(creg[130]), .B(init), .Z(n19359) );
  NAND U24481 ( .A(n19361), .B(n19362), .Z(x[12]) );
  NAND U24482 ( .A(creg[12]), .B(init), .Z(n19361) );
  NAND U24483 ( .A(n19363), .B(n19364), .Z(x[129]) );
  NAND U24484 ( .A(creg[129]), .B(init), .Z(n19363) );
  NAND U24485 ( .A(n19365), .B(n19366), .Z(x[128]) );
  NAND U24486 ( .A(creg[128]), .B(init), .Z(n19365) );
  NAND U24487 ( .A(n19367), .B(n19368), .Z(x[127]) );
  NAND U24488 ( .A(creg[127]), .B(init), .Z(n19367) );
  NAND U24489 ( .A(n19369), .B(n19370), .Z(x[126]) );
  NAND U24490 ( .A(creg[126]), .B(init), .Z(n19369) );
  NAND U24491 ( .A(n19371), .B(n19372), .Z(x[125]) );
  NAND U24492 ( .A(creg[125]), .B(init), .Z(n19371) );
  NAND U24493 ( .A(n19373), .B(n19374), .Z(x[124]) );
  NAND U24494 ( .A(creg[124]), .B(init), .Z(n19373) );
  NAND U24495 ( .A(n19375), .B(n19376), .Z(x[123]) );
  NAND U24496 ( .A(creg[123]), .B(init), .Z(n19375) );
  NAND U24497 ( .A(n19377), .B(n19378), .Z(x[122]) );
  NAND U24498 ( .A(creg[122]), .B(init), .Z(n19377) );
  NAND U24499 ( .A(n19379), .B(n19380), .Z(x[121]) );
  NAND U24500 ( .A(creg[121]), .B(init), .Z(n19379) );
  NAND U24501 ( .A(n19381), .B(n19382), .Z(x[120]) );
  NAND U24502 ( .A(creg[120]), .B(init), .Z(n19381) );
  NAND U24503 ( .A(n19383), .B(n19384), .Z(x[11]) );
  NAND U24504 ( .A(creg[11]), .B(init), .Z(n19383) );
  NAND U24505 ( .A(n19385), .B(n19386), .Z(x[119]) );
  NAND U24506 ( .A(creg[119]), .B(init), .Z(n19385) );
  NAND U24507 ( .A(n19387), .B(n19388), .Z(x[118]) );
  NAND U24508 ( .A(creg[118]), .B(init), .Z(n19387) );
  NAND U24509 ( .A(n19389), .B(n19390), .Z(x[117]) );
  NAND U24510 ( .A(creg[117]), .B(init), .Z(n19389) );
  NAND U24511 ( .A(n19391), .B(n19392), .Z(x[116]) );
  NAND U24512 ( .A(creg[116]), .B(init), .Z(n19391) );
  NAND U24513 ( .A(n19393), .B(n19394), .Z(x[115]) );
  NAND U24514 ( .A(creg[115]), .B(init), .Z(n19393) );
  NAND U24515 ( .A(n19395), .B(n19396), .Z(x[114]) );
  NAND U24516 ( .A(creg[114]), .B(init), .Z(n19395) );
  NAND U24517 ( .A(n19397), .B(n19398), .Z(x[113]) );
  NAND U24518 ( .A(creg[113]), .B(init), .Z(n19397) );
  NAND U24519 ( .A(n19399), .B(n19400), .Z(x[112]) );
  NAND U24520 ( .A(creg[112]), .B(init), .Z(n19399) );
  NAND U24521 ( .A(n19401), .B(n19402), .Z(x[111]) );
  NAND U24522 ( .A(creg[111]), .B(init), .Z(n19401) );
  NAND U24523 ( .A(n19403), .B(n19404), .Z(x[110]) );
  NAND U24524 ( .A(creg[110]), .B(init), .Z(n19403) );
  NAND U24525 ( .A(n19405), .B(n19406), .Z(x[10]) );
  NAND U24526 ( .A(creg[10]), .B(init), .Z(n19405) );
  NAND U24527 ( .A(n19407), .B(n19408), .Z(x[109]) );
  NAND U24528 ( .A(creg[109]), .B(init), .Z(n19407) );
  NAND U24529 ( .A(n19409), .B(n19410), .Z(x[108]) );
  NAND U24530 ( .A(creg[108]), .B(init), .Z(n19409) );
  NAND U24531 ( .A(n19411), .B(n19412), .Z(x[107]) );
  NAND U24532 ( .A(creg[107]), .B(init), .Z(n19411) );
  NAND U24533 ( .A(n19413), .B(n19414), .Z(x[106]) );
  NAND U24534 ( .A(creg[106]), .B(init), .Z(n19413) );
  NAND U24535 ( .A(n19415), .B(n19416), .Z(x[105]) );
  NAND U24536 ( .A(creg[105]), .B(init), .Z(n19415) );
  NAND U24537 ( .A(n19417), .B(n19418), .Z(x[104]) );
  NAND U24538 ( .A(creg[104]), .B(init), .Z(n19417) );
  NAND U24539 ( .A(n19419), .B(n19420), .Z(x[103]) );
  NAND U24540 ( .A(creg[103]), .B(init), .Z(n19419) );
  NAND U24541 ( .A(n19421), .B(n19422), .Z(x[102]) );
  NAND U24542 ( .A(creg[102]), .B(init), .Z(n19421) );
  NAND U24543 ( .A(n19423), .B(n19424), .Z(x[1023]) );
  NAND U24544 ( .A(creg[1023]), .B(init), .Z(n19423) );
  NAND U24545 ( .A(n19425), .B(n19426), .Z(x[1022]) );
  NAND U24546 ( .A(creg[1022]), .B(init), .Z(n19425) );
  NAND U24547 ( .A(n19427), .B(n19428), .Z(x[1021]) );
  NAND U24548 ( .A(creg[1021]), .B(init), .Z(n19427) );
  NAND U24549 ( .A(n19429), .B(n19430), .Z(x[1020]) );
  NAND U24550 ( .A(creg[1020]), .B(init), .Z(n19429) );
  NAND U24551 ( .A(n19431), .B(n19432), .Z(x[101]) );
  NAND U24552 ( .A(creg[101]), .B(init), .Z(n19431) );
  NAND U24553 ( .A(n19433), .B(n19434), .Z(x[1019]) );
  NAND U24554 ( .A(creg[1019]), .B(init), .Z(n19433) );
  NAND U24555 ( .A(n19435), .B(n19436), .Z(x[1018]) );
  NAND U24556 ( .A(creg[1018]), .B(init), .Z(n19435) );
  NAND U24557 ( .A(n19437), .B(n19438), .Z(x[1017]) );
  NAND U24558 ( .A(creg[1017]), .B(init), .Z(n19437) );
  NAND U24559 ( .A(n19439), .B(n19440), .Z(x[1016]) );
  NAND U24560 ( .A(creg[1016]), .B(init), .Z(n19439) );
  NAND U24561 ( .A(n19441), .B(n19442), .Z(x[1015]) );
  NAND U24562 ( .A(creg[1015]), .B(init), .Z(n19441) );
  NAND U24563 ( .A(n19443), .B(n19444), .Z(x[1014]) );
  NAND U24564 ( .A(creg[1014]), .B(init), .Z(n19443) );
  NAND U24565 ( .A(n19445), .B(n19446), .Z(x[1013]) );
  NAND U24566 ( .A(creg[1013]), .B(init), .Z(n19445) );
  NAND U24567 ( .A(n19447), .B(n19448), .Z(x[1012]) );
  NAND U24568 ( .A(creg[1012]), .B(init), .Z(n19447) );
  NAND U24569 ( .A(n19449), .B(n19450), .Z(x[1011]) );
  NAND U24570 ( .A(creg[1011]), .B(init), .Z(n19449) );
  NAND U24571 ( .A(n19451), .B(n19452), .Z(x[1010]) );
  NAND U24572 ( .A(creg[1010]), .B(init), .Z(n19451) );
  NAND U24573 ( .A(n19453), .B(n19454), .Z(x[100]) );
  NAND U24574 ( .A(creg[100]), .B(init), .Z(n19453) );
  NAND U24575 ( .A(n19455), .B(n19456), .Z(x[1009]) );
  NAND U24576 ( .A(creg[1009]), .B(init), .Z(n19455) );
  NAND U24577 ( .A(n19457), .B(n19458), .Z(x[1008]) );
  NAND U24578 ( .A(creg[1008]), .B(init), .Z(n19457) );
  NAND U24579 ( .A(n19459), .B(n19460), .Z(x[1007]) );
  NAND U24580 ( .A(creg[1007]), .B(init), .Z(n19459) );
  NAND U24581 ( .A(n19461), .B(n19462), .Z(x[1006]) );
  NAND U24582 ( .A(creg[1006]), .B(init), .Z(n19461) );
  NAND U24583 ( .A(n19463), .B(n19464), .Z(x[1005]) );
  NAND U24584 ( .A(creg[1005]), .B(init), .Z(n19463) );
  NAND U24585 ( .A(n19465), .B(n19466), .Z(x[1004]) );
  NAND U24586 ( .A(creg[1004]), .B(init), .Z(n19465) );
  NAND U24587 ( .A(n19467), .B(n19468), .Z(x[1003]) );
  NAND U24588 ( .A(creg[1003]), .B(init), .Z(n19467) );
  NAND U24589 ( .A(n19469), .B(n19470), .Z(x[1002]) );
  NAND U24590 ( .A(creg[1002]), .B(init), .Z(n19469) );
  NAND U24591 ( .A(n19471), .B(n19472), .Z(x[1001]) );
  NAND U24592 ( .A(creg[1001]), .B(init), .Z(n19471) );
  NAND U24593 ( .A(n19473), .B(n19474), .Z(x[1000]) );
  NAND U24594 ( .A(creg[1000]), .B(init), .Z(n19473) );
  NAND U24595 ( .A(n19475), .B(n19476), .Z(x[0]) );
  NAND U24596 ( .A(creg[0]), .B(init), .Z(n19475) );
  AND U24597 ( .A(start_reg[9]), .B(init), .Z(start_in[9]) );
  AND U24598 ( .A(start_reg[99]), .B(init), .Z(start_in[99]) );
  AND U24599 ( .A(start_reg[999]), .B(init), .Z(start_in[999]) );
  AND U24600 ( .A(start_reg[998]), .B(init), .Z(start_in[998]) );
  AND U24601 ( .A(start_reg[997]), .B(init), .Z(start_in[997]) );
  AND U24602 ( .A(start_reg[996]), .B(init), .Z(start_in[996]) );
  AND U24603 ( .A(start_reg[995]), .B(init), .Z(start_in[995]) );
  AND U24604 ( .A(start_reg[994]), .B(init), .Z(start_in[994]) );
  AND U24605 ( .A(start_reg[993]), .B(init), .Z(start_in[993]) );
  AND U24606 ( .A(start_reg[992]), .B(init), .Z(start_in[992]) );
  AND U24607 ( .A(start_reg[991]), .B(init), .Z(start_in[991]) );
  AND U24608 ( .A(start_reg[990]), .B(init), .Z(start_in[990]) );
  AND U24609 ( .A(start_reg[98]), .B(init), .Z(start_in[98]) );
  AND U24610 ( .A(start_reg[989]), .B(init), .Z(start_in[989]) );
  AND U24611 ( .A(start_reg[988]), .B(init), .Z(start_in[988]) );
  AND U24612 ( .A(start_reg[987]), .B(init), .Z(start_in[987]) );
  AND U24613 ( .A(start_reg[986]), .B(init), .Z(start_in[986]) );
  AND U24614 ( .A(start_reg[985]), .B(init), .Z(start_in[985]) );
  AND U24615 ( .A(start_reg[984]), .B(init), .Z(start_in[984]) );
  AND U24616 ( .A(start_reg[983]), .B(init), .Z(start_in[983]) );
  AND U24617 ( .A(start_reg[982]), .B(init), .Z(start_in[982]) );
  AND U24618 ( .A(start_reg[981]), .B(init), .Z(start_in[981]) );
  AND U24619 ( .A(start_reg[980]), .B(init), .Z(start_in[980]) );
  AND U24620 ( .A(start_reg[97]), .B(init), .Z(start_in[97]) );
  AND U24621 ( .A(start_reg[979]), .B(init), .Z(start_in[979]) );
  AND U24622 ( .A(start_reg[978]), .B(init), .Z(start_in[978]) );
  AND U24623 ( .A(start_reg[977]), .B(init), .Z(start_in[977]) );
  AND U24624 ( .A(start_reg[976]), .B(init), .Z(start_in[976]) );
  AND U24625 ( .A(start_reg[975]), .B(init), .Z(start_in[975]) );
  AND U24626 ( .A(start_reg[974]), .B(init), .Z(start_in[974]) );
  AND U24627 ( .A(start_reg[973]), .B(init), .Z(start_in[973]) );
  AND U24628 ( .A(start_reg[972]), .B(init), .Z(start_in[972]) );
  AND U24629 ( .A(start_reg[971]), .B(init), .Z(start_in[971]) );
  AND U24630 ( .A(start_reg[970]), .B(init), .Z(start_in[970]) );
  AND U24631 ( .A(start_reg[96]), .B(init), .Z(start_in[96]) );
  AND U24632 ( .A(start_reg[969]), .B(init), .Z(start_in[969]) );
  AND U24633 ( .A(start_reg[968]), .B(init), .Z(start_in[968]) );
  AND U24634 ( .A(start_reg[967]), .B(init), .Z(start_in[967]) );
  AND U24635 ( .A(start_reg[966]), .B(init), .Z(start_in[966]) );
  AND U24636 ( .A(start_reg[965]), .B(init), .Z(start_in[965]) );
  AND U24637 ( .A(start_reg[964]), .B(init), .Z(start_in[964]) );
  AND U24638 ( .A(start_reg[963]), .B(init), .Z(start_in[963]) );
  AND U24639 ( .A(start_reg[962]), .B(init), .Z(start_in[962]) );
  AND U24640 ( .A(start_reg[961]), .B(init), .Z(start_in[961]) );
  AND U24641 ( .A(start_reg[960]), .B(init), .Z(start_in[960]) );
  AND U24642 ( .A(start_reg[95]), .B(init), .Z(start_in[95]) );
  AND U24643 ( .A(start_reg[959]), .B(init), .Z(start_in[959]) );
  AND U24644 ( .A(start_reg[958]), .B(init), .Z(start_in[958]) );
  AND U24645 ( .A(start_reg[957]), .B(init), .Z(start_in[957]) );
  AND U24646 ( .A(start_reg[956]), .B(init), .Z(start_in[956]) );
  AND U24647 ( .A(start_reg[955]), .B(init), .Z(start_in[955]) );
  AND U24648 ( .A(start_reg[954]), .B(init), .Z(start_in[954]) );
  AND U24649 ( .A(start_reg[953]), .B(init), .Z(start_in[953]) );
  AND U24650 ( .A(start_reg[952]), .B(init), .Z(start_in[952]) );
  AND U24651 ( .A(start_reg[951]), .B(init), .Z(start_in[951]) );
  AND U24652 ( .A(start_reg[950]), .B(init), .Z(start_in[950]) );
  AND U24653 ( .A(start_reg[94]), .B(init), .Z(start_in[94]) );
  AND U24654 ( .A(start_reg[949]), .B(init), .Z(start_in[949]) );
  AND U24655 ( .A(start_reg[948]), .B(init), .Z(start_in[948]) );
  AND U24656 ( .A(start_reg[947]), .B(init), .Z(start_in[947]) );
  AND U24657 ( .A(start_reg[946]), .B(init), .Z(start_in[946]) );
  AND U24658 ( .A(start_reg[945]), .B(init), .Z(start_in[945]) );
  AND U24659 ( .A(start_reg[944]), .B(init), .Z(start_in[944]) );
  AND U24660 ( .A(start_reg[943]), .B(init), .Z(start_in[943]) );
  AND U24661 ( .A(start_reg[942]), .B(init), .Z(start_in[942]) );
  AND U24662 ( .A(start_reg[941]), .B(init), .Z(start_in[941]) );
  AND U24663 ( .A(start_reg[940]), .B(init), .Z(start_in[940]) );
  AND U24664 ( .A(start_reg[93]), .B(init), .Z(start_in[93]) );
  AND U24665 ( .A(start_reg[939]), .B(init), .Z(start_in[939]) );
  AND U24666 ( .A(start_reg[938]), .B(init), .Z(start_in[938]) );
  AND U24667 ( .A(start_reg[937]), .B(init), .Z(start_in[937]) );
  AND U24668 ( .A(start_reg[936]), .B(init), .Z(start_in[936]) );
  AND U24669 ( .A(start_reg[935]), .B(init), .Z(start_in[935]) );
  AND U24670 ( .A(start_reg[934]), .B(init), .Z(start_in[934]) );
  AND U24671 ( .A(start_reg[933]), .B(init), .Z(start_in[933]) );
  AND U24672 ( .A(start_reg[932]), .B(init), .Z(start_in[932]) );
  AND U24673 ( .A(start_reg[931]), .B(init), .Z(start_in[931]) );
  AND U24674 ( .A(start_reg[930]), .B(init), .Z(start_in[930]) );
  AND U24675 ( .A(start_reg[92]), .B(init), .Z(start_in[92]) );
  AND U24676 ( .A(start_reg[929]), .B(init), .Z(start_in[929]) );
  AND U24677 ( .A(start_reg[928]), .B(init), .Z(start_in[928]) );
  AND U24678 ( .A(start_reg[927]), .B(init), .Z(start_in[927]) );
  AND U24679 ( .A(start_reg[926]), .B(init), .Z(start_in[926]) );
  AND U24680 ( .A(start_reg[925]), .B(init), .Z(start_in[925]) );
  AND U24681 ( .A(start_reg[924]), .B(init), .Z(start_in[924]) );
  AND U24682 ( .A(start_reg[923]), .B(init), .Z(start_in[923]) );
  AND U24683 ( .A(start_reg[922]), .B(init), .Z(start_in[922]) );
  AND U24684 ( .A(start_reg[921]), .B(init), .Z(start_in[921]) );
  AND U24685 ( .A(start_reg[920]), .B(init), .Z(start_in[920]) );
  AND U24686 ( .A(start_reg[91]), .B(init), .Z(start_in[91]) );
  AND U24687 ( .A(start_reg[919]), .B(init), .Z(start_in[919]) );
  AND U24688 ( .A(start_reg[918]), .B(init), .Z(start_in[918]) );
  AND U24689 ( .A(start_reg[917]), .B(init), .Z(start_in[917]) );
  AND U24690 ( .A(start_reg[916]), .B(init), .Z(start_in[916]) );
  AND U24691 ( .A(start_reg[915]), .B(init), .Z(start_in[915]) );
  AND U24692 ( .A(start_reg[914]), .B(init), .Z(start_in[914]) );
  AND U24693 ( .A(start_reg[913]), .B(init), .Z(start_in[913]) );
  AND U24694 ( .A(start_reg[912]), .B(init), .Z(start_in[912]) );
  AND U24695 ( .A(start_reg[911]), .B(init), .Z(start_in[911]) );
  AND U24696 ( .A(start_reg[910]), .B(init), .Z(start_in[910]) );
  AND U24697 ( .A(start_reg[90]), .B(init), .Z(start_in[90]) );
  AND U24698 ( .A(start_reg[909]), .B(init), .Z(start_in[909]) );
  AND U24699 ( .A(start_reg[908]), .B(init), .Z(start_in[908]) );
  AND U24700 ( .A(start_reg[907]), .B(init), .Z(start_in[907]) );
  AND U24701 ( .A(start_reg[906]), .B(init), .Z(start_in[906]) );
  AND U24702 ( .A(start_reg[905]), .B(init), .Z(start_in[905]) );
  AND U24703 ( .A(start_reg[904]), .B(init), .Z(start_in[904]) );
  AND U24704 ( .A(start_reg[903]), .B(init), .Z(start_in[903]) );
  AND U24705 ( .A(start_reg[902]), .B(init), .Z(start_in[902]) );
  AND U24706 ( .A(start_reg[901]), .B(init), .Z(start_in[901]) );
  AND U24707 ( .A(start_reg[900]), .B(init), .Z(start_in[900]) );
  AND U24708 ( .A(start_reg[8]), .B(init), .Z(start_in[8]) );
  AND U24709 ( .A(start_reg[89]), .B(init), .Z(start_in[89]) );
  AND U24710 ( .A(start_reg[899]), .B(init), .Z(start_in[899]) );
  AND U24711 ( .A(start_reg[898]), .B(init), .Z(start_in[898]) );
  AND U24712 ( .A(start_reg[897]), .B(init), .Z(start_in[897]) );
  AND U24713 ( .A(start_reg[896]), .B(init), .Z(start_in[896]) );
  AND U24714 ( .A(start_reg[895]), .B(init), .Z(start_in[895]) );
  AND U24715 ( .A(start_reg[894]), .B(init), .Z(start_in[894]) );
  AND U24716 ( .A(start_reg[893]), .B(init), .Z(start_in[893]) );
  AND U24717 ( .A(start_reg[892]), .B(init), .Z(start_in[892]) );
  AND U24718 ( .A(start_reg[891]), .B(init), .Z(start_in[891]) );
  AND U24719 ( .A(start_reg[890]), .B(init), .Z(start_in[890]) );
  AND U24720 ( .A(start_reg[88]), .B(init), .Z(start_in[88]) );
  AND U24721 ( .A(start_reg[889]), .B(init), .Z(start_in[889]) );
  AND U24722 ( .A(start_reg[888]), .B(init), .Z(start_in[888]) );
  AND U24723 ( .A(start_reg[887]), .B(init), .Z(start_in[887]) );
  AND U24724 ( .A(start_reg[886]), .B(init), .Z(start_in[886]) );
  AND U24725 ( .A(start_reg[885]), .B(init), .Z(start_in[885]) );
  AND U24726 ( .A(start_reg[884]), .B(init), .Z(start_in[884]) );
  AND U24727 ( .A(start_reg[883]), .B(init), .Z(start_in[883]) );
  AND U24728 ( .A(start_reg[882]), .B(init), .Z(start_in[882]) );
  AND U24729 ( .A(start_reg[881]), .B(init), .Z(start_in[881]) );
  AND U24730 ( .A(start_reg[880]), .B(init), .Z(start_in[880]) );
  AND U24731 ( .A(start_reg[87]), .B(init), .Z(start_in[87]) );
  AND U24732 ( .A(start_reg[879]), .B(init), .Z(start_in[879]) );
  AND U24733 ( .A(start_reg[878]), .B(init), .Z(start_in[878]) );
  AND U24734 ( .A(start_reg[877]), .B(init), .Z(start_in[877]) );
  AND U24735 ( .A(start_reg[876]), .B(init), .Z(start_in[876]) );
  AND U24736 ( .A(start_reg[875]), .B(init), .Z(start_in[875]) );
  AND U24737 ( .A(start_reg[874]), .B(init), .Z(start_in[874]) );
  AND U24738 ( .A(start_reg[873]), .B(init), .Z(start_in[873]) );
  AND U24739 ( .A(start_reg[872]), .B(init), .Z(start_in[872]) );
  AND U24740 ( .A(start_reg[871]), .B(init), .Z(start_in[871]) );
  AND U24741 ( .A(start_reg[870]), .B(init), .Z(start_in[870]) );
  AND U24742 ( .A(start_reg[86]), .B(init), .Z(start_in[86]) );
  AND U24743 ( .A(start_reg[869]), .B(init), .Z(start_in[869]) );
  AND U24744 ( .A(start_reg[868]), .B(init), .Z(start_in[868]) );
  AND U24745 ( .A(start_reg[867]), .B(init), .Z(start_in[867]) );
  AND U24746 ( .A(start_reg[866]), .B(init), .Z(start_in[866]) );
  AND U24747 ( .A(start_reg[865]), .B(init), .Z(start_in[865]) );
  AND U24748 ( .A(start_reg[864]), .B(init), .Z(start_in[864]) );
  AND U24749 ( .A(start_reg[863]), .B(init), .Z(start_in[863]) );
  AND U24750 ( .A(start_reg[862]), .B(init), .Z(start_in[862]) );
  AND U24751 ( .A(start_reg[861]), .B(init), .Z(start_in[861]) );
  AND U24752 ( .A(start_reg[860]), .B(init), .Z(start_in[860]) );
  AND U24753 ( .A(start_reg[85]), .B(init), .Z(start_in[85]) );
  AND U24754 ( .A(start_reg[859]), .B(init), .Z(start_in[859]) );
  AND U24755 ( .A(start_reg[858]), .B(init), .Z(start_in[858]) );
  AND U24756 ( .A(start_reg[857]), .B(init), .Z(start_in[857]) );
  AND U24757 ( .A(start_reg[856]), .B(init), .Z(start_in[856]) );
  AND U24758 ( .A(start_reg[855]), .B(init), .Z(start_in[855]) );
  AND U24759 ( .A(start_reg[854]), .B(init), .Z(start_in[854]) );
  AND U24760 ( .A(start_reg[853]), .B(init), .Z(start_in[853]) );
  AND U24761 ( .A(start_reg[852]), .B(init), .Z(start_in[852]) );
  AND U24762 ( .A(start_reg[851]), .B(init), .Z(start_in[851]) );
  AND U24763 ( .A(start_reg[850]), .B(init), .Z(start_in[850]) );
  AND U24764 ( .A(start_reg[84]), .B(init), .Z(start_in[84]) );
  AND U24765 ( .A(start_reg[849]), .B(init), .Z(start_in[849]) );
  AND U24766 ( .A(start_reg[848]), .B(init), .Z(start_in[848]) );
  AND U24767 ( .A(start_reg[847]), .B(init), .Z(start_in[847]) );
  AND U24768 ( .A(start_reg[846]), .B(init), .Z(start_in[846]) );
  AND U24769 ( .A(start_reg[845]), .B(init), .Z(start_in[845]) );
  AND U24770 ( .A(start_reg[844]), .B(init), .Z(start_in[844]) );
  AND U24771 ( .A(start_reg[843]), .B(init), .Z(start_in[843]) );
  AND U24772 ( .A(start_reg[842]), .B(init), .Z(start_in[842]) );
  AND U24773 ( .A(start_reg[841]), .B(init), .Z(start_in[841]) );
  AND U24774 ( .A(start_reg[840]), .B(init), .Z(start_in[840]) );
  AND U24775 ( .A(start_reg[83]), .B(init), .Z(start_in[83]) );
  AND U24776 ( .A(start_reg[839]), .B(init), .Z(start_in[839]) );
  AND U24777 ( .A(start_reg[838]), .B(init), .Z(start_in[838]) );
  AND U24778 ( .A(start_reg[837]), .B(init), .Z(start_in[837]) );
  AND U24779 ( .A(start_reg[836]), .B(init), .Z(start_in[836]) );
  AND U24780 ( .A(start_reg[835]), .B(init), .Z(start_in[835]) );
  AND U24781 ( .A(start_reg[834]), .B(init), .Z(start_in[834]) );
  AND U24782 ( .A(start_reg[833]), .B(init), .Z(start_in[833]) );
  AND U24783 ( .A(start_reg[832]), .B(init), .Z(start_in[832]) );
  AND U24784 ( .A(start_reg[831]), .B(init), .Z(start_in[831]) );
  AND U24785 ( .A(start_reg[830]), .B(init), .Z(start_in[830]) );
  AND U24786 ( .A(start_reg[82]), .B(init), .Z(start_in[82]) );
  AND U24787 ( .A(start_reg[829]), .B(init), .Z(start_in[829]) );
  AND U24788 ( .A(start_reg[828]), .B(init), .Z(start_in[828]) );
  AND U24789 ( .A(start_reg[827]), .B(init), .Z(start_in[827]) );
  AND U24790 ( .A(start_reg[826]), .B(init), .Z(start_in[826]) );
  AND U24791 ( .A(start_reg[825]), .B(init), .Z(start_in[825]) );
  AND U24792 ( .A(start_reg[824]), .B(init), .Z(start_in[824]) );
  AND U24793 ( .A(start_reg[823]), .B(init), .Z(start_in[823]) );
  AND U24794 ( .A(start_reg[822]), .B(init), .Z(start_in[822]) );
  AND U24795 ( .A(start_reg[821]), .B(init), .Z(start_in[821]) );
  AND U24796 ( .A(start_reg[820]), .B(init), .Z(start_in[820]) );
  AND U24797 ( .A(start_reg[81]), .B(init), .Z(start_in[81]) );
  AND U24798 ( .A(start_reg[819]), .B(init), .Z(start_in[819]) );
  AND U24799 ( .A(start_reg[818]), .B(init), .Z(start_in[818]) );
  AND U24800 ( .A(start_reg[817]), .B(init), .Z(start_in[817]) );
  AND U24801 ( .A(start_reg[816]), .B(init), .Z(start_in[816]) );
  AND U24802 ( .A(start_reg[815]), .B(init), .Z(start_in[815]) );
  AND U24803 ( .A(start_reg[814]), .B(init), .Z(start_in[814]) );
  AND U24804 ( .A(start_reg[813]), .B(init), .Z(start_in[813]) );
  AND U24805 ( .A(start_reg[812]), .B(init), .Z(start_in[812]) );
  AND U24806 ( .A(start_reg[811]), .B(init), .Z(start_in[811]) );
  AND U24807 ( .A(start_reg[810]), .B(init), .Z(start_in[810]) );
  AND U24808 ( .A(start_reg[80]), .B(init), .Z(start_in[80]) );
  AND U24809 ( .A(start_reg[809]), .B(init), .Z(start_in[809]) );
  AND U24810 ( .A(start_reg[808]), .B(init), .Z(start_in[808]) );
  AND U24811 ( .A(start_reg[807]), .B(init), .Z(start_in[807]) );
  AND U24812 ( .A(start_reg[806]), .B(init), .Z(start_in[806]) );
  AND U24813 ( .A(start_reg[805]), .B(init), .Z(start_in[805]) );
  AND U24814 ( .A(start_reg[804]), .B(init), .Z(start_in[804]) );
  AND U24815 ( .A(start_reg[803]), .B(init), .Z(start_in[803]) );
  AND U24816 ( .A(start_reg[802]), .B(init), .Z(start_in[802]) );
  AND U24817 ( .A(start_reg[801]), .B(init), .Z(start_in[801]) );
  AND U24818 ( .A(start_reg[800]), .B(init), .Z(start_in[800]) );
  AND U24819 ( .A(start_reg[7]), .B(init), .Z(start_in[7]) );
  AND U24820 ( .A(start_reg[79]), .B(init), .Z(start_in[79]) );
  AND U24821 ( .A(start_reg[799]), .B(init), .Z(start_in[799]) );
  AND U24822 ( .A(start_reg[798]), .B(init), .Z(start_in[798]) );
  AND U24823 ( .A(start_reg[797]), .B(init), .Z(start_in[797]) );
  AND U24824 ( .A(start_reg[796]), .B(init), .Z(start_in[796]) );
  AND U24825 ( .A(start_reg[795]), .B(init), .Z(start_in[795]) );
  AND U24826 ( .A(start_reg[794]), .B(init), .Z(start_in[794]) );
  AND U24827 ( .A(start_reg[793]), .B(init), .Z(start_in[793]) );
  AND U24828 ( .A(start_reg[792]), .B(init), .Z(start_in[792]) );
  AND U24829 ( .A(start_reg[791]), .B(init), .Z(start_in[791]) );
  AND U24830 ( .A(start_reg[790]), .B(init), .Z(start_in[790]) );
  AND U24831 ( .A(start_reg[78]), .B(init), .Z(start_in[78]) );
  AND U24832 ( .A(start_reg[789]), .B(init), .Z(start_in[789]) );
  AND U24833 ( .A(start_reg[788]), .B(init), .Z(start_in[788]) );
  AND U24834 ( .A(start_reg[787]), .B(init), .Z(start_in[787]) );
  AND U24835 ( .A(start_reg[786]), .B(init), .Z(start_in[786]) );
  AND U24836 ( .A(start_reg[785]), .B(init), .Z(start_in[785]) );
  AND U24837 ( .A(start_reg[784]), .B(init), .Z(start_in[784]) );
  AND U24838 ( .A(start_reg[783]), .B(init), .Z(start_in[783]) );
  AND U24839 ( .A(start_reg[782]), .B(init), .Z(start_in[782]) );
  AND U24840 ( .A(start_reg[781]), .B(init), .Z(start_in[781]) );
  AND U24841 ( .A(start_reg[780]), .B(init), .Z(start_in[780]) );
  AND U24842 ( .A(start_reg[77]), .B(init), .Z(start_in[77]) );
  AND U24843 ( .A(start_reg[779]), .B(init), .Z(start_in[779]) );
  AND U24844 ( .A(start_reg[778]), .B(init), .Z(start_in[778]) );
  AND U24845 ( .A(start_reg[777]), .B(init), .Z(start_in[777]) );
  AND U24846 ( .A(start_reg[776]), .B(init), .Z(start_in[776]) );
  AND U24847 ( .A(start_reg[775]), .B(init), .Z(start_in[775]) );
  AND U24848 ( .A(start_reg[774]), .B(init), .Z(start_in[774]) );
  AND U24849 ( .A(start_reg[773]), .B(init), .Z(start_in[773]) );
  AND U24850 ( .A(start_reg[772]), .B(init), .Z(start_in[772]) );
  AND U24851 ( .A(start_reg[771]), .B(init), .Z(start_in[771]) );
  AND U24852 ( .A(start_reg[770]), .B(init), .Z(start_in[770]) );
  AND U24853 ( .A(start_reg[76]), .B(init), .Z(start_in[76]) );
  AND U24854 ( .A(start_reg[769]), .B(init), .Z(start_in[769]) );
  AND U24855 ( .A(start_reg[768]), .B(init), .Z(start_in[768]) );
  AND U24856 ( .A(start_reg[767]), .B(init), .Z(start_in[767]) );
  AND U24857 ( .A(start_reg[766]), .B(init), .Z(start_in[766]) );
  AND U24858 ( .A(start_reg[765]), .B(init), .Z(start_in[765]) );
  AND U24859 ( .A(start_reg[764]), .B(init), .Z(start_in[764]) );
  AND U24860 ( .A(start_reg[763]), .B(init), .Z(start_in[763]) );
  AND U24861 ( .A(start_reg[762]), .B(init), .Z(start_in[762]) );
  AND U24862 ( .A(start_reg[761]), .B(init), .Z(start_in[761]) );
  AND U24863 ( .A(start_reg[760]), .B(init), .Z(start_in[760]) );
  AND U24864 ( .A(start_reg[75]), .B(init), .Z(start_in[75]) );
  AND U24865 ( .A(start_reg[759]), .B(init), .Z(start_in[759]) );
  AND U24866 ( .A(start_reg[758]), .B(init), .Z(start_in[758]) );
  AND U24867 ( .A(start_reg[757]), .B(init), .Z(start_in[757]) );
  AND U24868 ( .A(start_reg[756]), .B(init), .Z(start_in[756]) );
  AND U24869 ( .A(start_reg[755]), .B(init), .Z(start_in[755]) );
  AND U24870 ( .A(start_reg[754]), .B(init), .Z(start_in[754]) );
  AND U24871 ( .A(start_reg[753]), .B(init), .Z(start_in[753]) );
  AND U24872 ( .A(start_reg[752]), .B(init), .Z(start_in[752]) );
  AND U24873 ( .A(start_reg[751]), .B(init), .Z(start_in[751]) );
  AND U24874 ( .A(start_reg[750]), .B(init), .Z(start_in[750]) );
  AND U24875 ( .A(start_reg[74]), .B(init), .Z(start_in[74]) );
  AND U24876 ( .A(start_reg[749]), .B(init), .Z(start_in[749]) );
  AND U24877 ( .A(start_reg[748]), .B(init), .Z(start_in[748]) );
  AND U24878 ( .A(start_reg[747]), .B(init), .Z(start_in[747]) );
  AND U24879 ( .A(start_reg[746]), .B(init), .Z(start_in[746]) );
  AND U24880 ( .A(start_reg[745]), .B(init), .Z(start_in[745]) );
  AND U24881 ( .A(start_reg[744]), .B(init), .Z(start_in[744]) );
  AND U24882 ( .A(start_reg[743]), .B(init), .Z(start_in[743]) );
  AND U24883 ( .A(start_reg[742]), .B(init), .Z(start_in[742]) );
  AND U24884 ( .A(start_reg[741]), .B(init), .Z(start_in[741]) );
  AND U24885 ( .A(start_reg[740]), .B(init), .Z(start_in[740]) );
  AND U24886 ( .A(start_reg[73]), .B(init), .Z(start_in[73]) );
  AND U24887 ( .A(start_reg[739]), .B(init), .Z(start_in[739]) );
  AND U24888 ( .A(start_reg[738]), .B(init), .Z(start_in[738]) );
  AND U24889 ( .A(start_reg[737]), .B(init), .Z(start_in[737]) );
  AND U24890 ( .A(start_reg[736]), .B(init), .Z(start_in[736]) );
  AND U24891 ( .A(start_reg[735]), .B(init), .Z(start_in[735]) );
  AND U24892 ( .A(start_reg[734]), .B(init), .Z(start_in[734]) );
  AND U24893 ( .A(start_reg[733]), .B(init), .Z(start_in[733]) );
  AND U24894 ( .A(start_reg[732]), .B(init), .Z(start_in[732]) );
  AND U24895 ( .A(start_reg[731]), .B(init), .Z(start_in[731]) );
  AND U24896 ( .A(start_reg[730]), .B(init), .Z(start_in[730]) );
  AND U24897 ( .A(start_reg[72]), .B(init), .Z(start_in[72]) );
  AND U24898 ( .A(start_reg[729]), .B(init), .Z(start_in[729]) );
  AND U24899 ( .A(start_reg[728]), .B(init), .Z(start_in[728]) );
  AND U24900 ( .A(start_reg[727]), .B(init), .Z(start_in[727]) );
  AND U24901 ( .A(start_reg[726]), .B(init), .Z(start_in[726]) );
  AND U24902 ( .A(start_reg[725]), .B(init), .Z(start_in[725]) );
  AND U24903 ( .A(start_reg[724]), .B(init), .Z(start_in[724]) );
  AND U24904 ( .A(start_reg[723]), .B(init), .Z(start_in[723]) );
  AND U24905 ( .A(start_reg[722]), .B(init), .Z(start_in[722]) );
  AND U24906 ( .A(start_reg[721]), .B(init), .Z(start_in[721]) );
  AND U24907 ( .A(start_reg[720]), .B(init), .Z(start_in[720]) );
  AND U24908 ( .A(start_reg[71]), .B(init), .Z(start_in[71]) );
  AND U24909 ( .A(start_reg[719]), .B(init), .Z(start_in[719]) );
  AND U24910 ( .A(start_reg[718]), .B(init), .Z(start_in[718]) );
  AND U24911 ( .A(start_reg[717]), .B(init), .Z(start_in[717]) );
  AND U24912 ( .A(start_reg[716]), .B(init), .Z(start_in[716]) );
  AND U24913 ( .A(start_reg[715]), .B(init), .Z(start_in[715]) );
  AND U24914 ( .A(start_reg[714]), .B(init), .Z(start_in[714]) );
  AND U24915 ( .A(start_reg[713]), .B(init), .Z(start_in[713]) );
  AND U24916 ( .A(start_reg[712]), .B(init), .Z(start_in[712]) );
  AND U24917 ( .A(start_reg[711]), .B(init), .Z(start_in[711]) );
  AND U24918 ( .A(start_reg[710]), .B(init), .Z(start_in[710]) );
  AND U24919 ( .A(start_reg[70]), .B(init), .Z(start_in[70]) );
  AND U24920 ( .A(start_reg[709]), .B(init), .Z(start_in[709]) );
  AND U24921 ( .A(start_reg[708]), .B(init), .Z(start_in[708]) );
  AND U24922 ( .A(start_reg[707]), .B(init), .Z(start_in[707]) );
  AND U24923 ( .A(start_reg[706]), .B(init), .Z(start_in[706]) );
  AND U24924 ( .A(start_reg[705]), .B(init), .Z(start_in[705]) );
  AND U24925 ( .A(start_reg[704]), .B(init), .Z(start_in[704]) );
  AND U24926 ( .A(start_reg[703]), .B(init), .Z(start_in[703]) );
  AND U24927 ( .A(start_reg[702]), .B(init), .Z(start_in[702]) );
  AND U24928 ( .A(start_reg[701]), .B(init), .Z(start_in[701]) );
  AND U24929 ( .A(start_reg[700]), .B(init), .Z(start_in[700]) );
  AND U24930 ( .A(start_reg[6]), .B(init), .Z(start_in[6]) );
  AND U24931 ( .A(start_reg[69]), .B(init), .Z(start_in[69]) );
  AND U24932 ( .A(start_reg[699]), .B(init), .Z(start_in[699]) );
  AND U24933 ( .A(start_reg[698]), .B(init), .Z(start_in[698]) );
  AND U24934 ( .A(start_reg[697]), .B(init), .Z(start_in[697]) );
  AND U24935 ( .A(start_reg[696]), .B(init), .Z(start_in[696]) );
  AND U24936 ( .A(start_reg[695]), .B(init), .Z(start_in[695]) );
  AND U24937 ( .A(start_reg[694]), .B(init), .Z(start_in[694]) );
  AND U24938 ( .A(start_reg[693]), .B(init), .Z(start_in[693]) );
  AND U24939 ( .A(start_reg[692]), .B(init), .Z(start_in[692]) );
  AND U24940 ( .A(start_reg[691]), .B(init), .Z(start_in[691]) );
  AND U24941 ( .A(start_reg[690]), .B(init), .Z(start_in[690]) );
  AND U24942 ( .A(start_reg[68]), .B(init), .Z(start_in[68]) );
  AND U24943 ( .A(start_reg[689]), .B(init), .Z(start_in[689]) );
  AND U24944 ( .A(start_reg[688]), .B(init), .Z(start_in[688]) );
  AND U24945 ( .A(start_reg[687]), .B(init), .Z(start_in[687]) );
  AND U24946 ( .A(start_reg[686]), .B(init), .Z(start_in[686]) );
  AND U24947 ( .A(start_reg[685]), .B(init), .Z(start_in[685]) );
  AND U24948 ( .A(start_reg[684]), .B(init), .Z(start_in[684]) );
  AND U24949 ( .A(start_reg[683]), .B(init), .Z(start_in[683]) );
  AND U24950 ( .A(start_reg[682]), .B(init), .Z(start_in[682]) );
  AND U24951 ( .A(start_reg[681]), .B(init), .Z(start_in[681]) );
  AND U24952 ( .A(start_reg[680]), .B(init), .Z(start_in[680]) );
  AND U24953 ( .A(start_reg[67]), .B(init), .Z(start_in[67]) );
  AND U24954 ( .A(start_reg[679]), .B(init), .Z(start_in[679]) );
  AND U24955 ( .A(start_reg[678]), .B(init), .Z(start_in[678]) );
  AND U24956 ( .A(start_reg[677]), .B(init), .Z(start_in[677]) );
  AND U24957 ( .A(start_reg[676]), .B(init), .Z(start_in[676]) );
  AND U24958 ( .A(start_reg[675]), .B(init), .Z(start_in[675]) );
  AND U24959 ( .A(start_reg[674]), .B(init), .Z(start_in[674]) );
  AND U24960 ( .A(start_reg[673]), .B(init), .Z(start_in[673]) );
  AND U24961 ( .A(start_reg[672]), .B(init), .Z(start_in[672]) );
  AND U24962 ( .A(start_reg[671]), .B(init), .Z(start_in[671]) );
  AND U24963 ( .A(start_reg[670]), .B(init), .Z(start_in[670]) );
  AND U24964 ( .A(start_reg[66]), .B(init), .Z(start_in[66]) );
  AND U24965 ( .A(start_reg[669]), .B(init), .Z(start_in[669]) );
  AND U24966 ( .A(start_reg[668]), .B(init), .Z(start_in[668]) );
  AND U24967 ( .A(start_reg[667]), .B(init), .Z(start_in[667]) );
  AND U24968 ( .A(start_reg[666]), .B(init), .Z(start_in[666]) );
  AND U24969 ( .A(start_reg[665]), .B(init), .Z(start_in[665]) );
  AND U24970 ( .A(start_reg[664]), .B(init), .Z(start_in[664]) );
  AND U24971 ( .A(start_reg[663]), .B(init), .Z(start_in[663]) );
  AND U24972 ( .A(start_reg[662]), .B(init), .Z(start_in[662]) );
  AND U24973 ( .A(start_reg[661]), .B(init), .Z(start_in[661]) );
  AND U24974 ( .A(start_reg[660]), .B(init), .Z(start_in[660]) );
  AND U24975 ( .A(start_reg[65]), .B(init), .Z(start_in[65]) );
  AND U24976 ( .A(start_reg[659]), .B(init), .Z(start_in[659]) );
  AND U24977 ( .A(start_reg[658]), .B(init), .Z(start_in[658]) );
  AND U24978 ( .A(start_reg[657]), .B(init), .Z(start_in[657]) );
  AND U24979 ( .A(start_reg[656]), .B(init), .Z(start_in[656]) );
  AND U24980 ( .A(start_reg[655]), .B(init), .Z(start_in[655]) );
  AND U24981 ( .A(start_reg[654]), .B(init), .Z(start_in[654]) );
  AND U24982 ( .A(start_reg[653]), .B(init), .Z(start_in[653]) );
  AND U24983 ( .A(start_reg[652]), .B(init), .Z(start_in[652]) );
  AND U24984 ( .A(start_reg[651]), .B(init), .Z(start_in[651]) );
  AND U24985 ( .A(start_reg[650]), .B(init), .Z(start_in[650]) );
  AND U24986 ( .A(start_reg[64]), .B(init), .Z(start_in[64]) );
  AND U24987 ( .A(start_reg[649]), .B(init), .Z(start_in[649]) );
  AND U24988 ( .A(start_reg[648]), .B(init), .Z(start_in[648]) );
  AND U24989 ( .A(start_reg[647]), .B(init), .Z(start_in[647]) );
  AND U24990 ( .A(start_reg[646]), .B(init), .Z(start_in[646]) );
  AND U24991 ( .A(start_reg[645]), .B(init), .Z(start_in[645]) );
  AND U24992 ( .A(start_reg[644]), .B(init), .Z(start_in[644]) );
  AND U24993 ( .A(start_reg[643]), .B(init), .Z(start_in[643]) );
  AND U24994 ( .A(start_reg[642]), .B(init), .Z(start_in[642]) );
  AND U24995 ( .A(start_reg[641]), .B(init), .Z(start_in[641]) );
  AND U24996 ( .A(start_reg[640]), .B(init), .Z(start_in[640]) );
  AND U24997 ( .A(start_reg[63]), .B(init), .Z(start_in[63]) );
  AND U24998 ( .A(start_reg[639]), .B(init), .Z(start_in[639]) );
  AND U24999 ( .A(start_reg[638]), .B(init), .Z(start_in[638]) );
  AND U25000 ( .A(start_reg[637]), .B(init), .Z(start_in[637]) );
  AND U25001 ( .A(start_reg[636]), .B(init), .Z(start_in[636]) );
  AND U25002 ( .A(start_reg[635]), .B(init), .Z(start_in[635]) );
  AND U25003 ( .A(start_reg[634]), .B(init), .Z(start_in[634]) );
  AND U25004 ( .A(start_reg[633]), .B(init), .Z(start_in[633]) );
  AND U25005 ( .A(start_reg[632]), .B(init), .Z(start_in[632]) );
  AND U25006 ( .A(start_reg[631]), .B(init), .Z(start_in[631]) );
  AND U25007 ( .A(start_reg[630]), .B(init), .Z(start_in[630]) );
  AND U25008 ( .A(start_reg[62]), .B(init), .Z(start_in[62]) );
  AND U25009 ( .A(start_reg[629]), .B(init), .Z(start_in[629]) );
  AND U25010 ( .A(start_reg[628]), .B(init), .Z(start_in[628]) );
  AND U25011 ( .A(start_reg[627]), .B(init), .Z(start_in[627]) );
  AND U25012 ( .A(start_reg[626]), .B(init), .Z(start_in[626]) );
  AND U25013 ( .A(start_reg[625]), .B(init), .Z(start_in[625]) );
  AND U25014 ( .A(start_reg[624]), .B(init), .Z(start_in[624]) );
  AND U25015 ( .A(start_reg[623]), .B(init), .Z(start_in[623]) );
  AND U25016 ( .A(start_reg[622]), .B(init), .Z(start_in[622]) );
  AND U25017 ( .A(start_reg[621]), .B(init), .Z(start_in[621]) );
  AND U25018 ( .A(start_reg[620]), .B(init), .Z(start_in[620]) );
  AND U25019 ( .A(start_reg[61]), .B(init), .Z(start_in[61]) );
  AND U25020 ( .A(start_reg[619]), .B(init), .Z(start_in[619]) );
  AND U25021 ( .A(start_reg[618]), .B(init), .Z(start_in[618]) );
  AND U25022 ( .A(start_reg[617]), .B(init), .Z(start_in[617]) );
  AND U25023 ( .A(start_reg[616]), .B(init), .Z(start_in[616]) );
  AND U25024 ( .A(start_reg[615]), .B(init), .Z(start_in[615]) );
  AND U25025 ( .A(start_reg[614]), .B(init), .Z(start_in[614]) );
  AND U25026 ( .A(start_reg[613]), .B(init), .Z(start_in[613]) );
  AND U25027 ( .A(start_reg[612]), .B(init), .Z(start_in[612]) );
  AND U25028 ( .A(start_reg[611]), .B(init), .Z(start_in[611]) );
  AND U25029 ( .A(start_reg[610]), .B(init), .Z(start_in[610]) );
  AND U25030 ( .A(start_reg[60]), .B(init), .Z(start_in[60]) );
  AND U25031 ( .A(start_reg[609]), .B(init), .Z(start_in[609]) );
  AND U25032 ( .A(start_reg[608]), .B(init), .Z(start_in[608]) );
  AND U25033 ( .A(start_reg[607]), .B(init), .Z(start_in[607]) );
  AND U25034 ( .A(start_reg[606]), .B(init), .Z(start_in[606]) );
  AND U25035 ( .A(start_reg[605]), .B(init), .Z(start_in[605]) );
  AND U25036 ( .A(start_reg[604]), .B(init), .Z(start_in[604]) );
  AND U25037 ( .A(start_reg[603]), .B(init), .Z(start_in[603]) );
  AND U25038 ( .A(start_reg[602]), .B(init), .Z(start_in[602]) );
  AND U25039 ( .A(start_reg[601]), .B(init), .Z(start_in[601]) );
  AND U25040 ( .A(start_reg[600]), .B(init), .Z(start_in[600]) );
  AND U25041 ( .A(start_reg[5]), .B(init), .Z(start_in[5]) );
  AND U25042 ( .A(start_reg[59]), .B(init), .Z(start_in[59]) );
  AND U25043 ( .A(start_reg[599]), .B(init), .Z(start_in[599]) );
  AND U25044 ( .A(start_reg[598]), .B(init), .Z(start_in[598]) );
  AND U25045 ( .A(start_reg[597]), .B(init), .Z(start_in[597]) );
  AND U25046 ( .A(start_reg[596]), .B(init), .Z(start_in[596]) );
  AND U25047 ( .A(start_reg[595]), .B(init), .Z(start_in[595]) );
  AND U25048 ( .A(start_reg[594]), .B(init), .Z(start_in[594]) );
  AND U25049 ( .A(start_reg[593]), .B(init), .Z(start_in[593]) );
  AND U25050 ( .A(start_reg[592]), .B(init), .Z(start_in[592]) );
  AND U25051 ( .A(start_reg[591]), .B(init), .Z(start_in[591]) );
  AND U25052 ( .A(start_reg[590]), .B(init), .Z(start_in[590]) );
  AND U25053 ( .A(start_reg[58]), .B(init), .Z(start_in[58]) );
  AND U25054 ( .A(start_reg[589]), .B(init), .Z(start_in[589]) );
  AND U25055 ( .A(start_reg[588]), .B(init), .Z(start_in[588]) );
  AND U25056 ( .A(start_reg[587]), .B(init), .Z(start_in[587]) );
  AND U25057 ( .A(start_reg[586]), .B(init), .Z(start_in[586]) );
  AND U25058 ( .A(start_reg[585]), .B(init), .Z(start_in[585]) );
  AND U25059 ( .A(start_reg[584]), .B(init), .Z(start_in[584]) );
  AND U25060 ( .A(start_reg[583]), .B(init), .Z(start_in[583]) );
  AND U25061 ( .A(start_reg[582]), .B(init), .Z(start_in[582]) );
  AND U25062 ( .A(start_reg[581]), .B(init), .Z(start_in[581]) );
  AND U25063 ( .A(start_reg[580]), .B(init), .Z(start_in[580]) );
  AND U25064 ( .A(start_reg[57]), .B(init), .Z(start_in[57]) );
  AND U25065 ( .A(start_reg[579]), .B(init), .Z(start_in[579]) );
  AND U25066 ( .A(start_reg[578]), .B(init), .Z(start_in[578]) );
  AND U25067 ( .A(start_reg[577]), .B(init), .Z(start_in[577]) );
  AND U25068 ( .A(start_reg[576]), .B(init), .Z(start_in[576]) );
  AND U25069 ( .A(start_reg[575]), .B(init), .Z(start_in[575]) );
  AND U25070 ( .A(start_reg[574]), .B(init), .Z(start_in[574]) );
  AND U25071 ( .A(start_reg[573]), .B(init), .Z(start_in[573]) );
  AND U25072 ( .A(start_reg[572]), .B(init), .Z(start_in[572]) );
  AND U25073 ( .A(start_reg[571]), .B(init), .Z(start_in[571]) );
  AND U25074 ( .A(start_reg[570]), .B(init), .Z(start_in[570]) );
  AND U25075 ( .A(start_reg[56]), .B(init), .Z(start_in[56]) );
  AND U25076 ( .A(start_reg[569]), .B(init), .Z(start_in[569]) );
  AND U25077 ( .A(start_reg[568]), .B(init), .Z(start_in[568]) );
  AND U25078 ( .A(start_reg[567]), .B(init), .Z(start_in[567]) );
  AND U25079 ( .A(start_reg[566]), .B(init), .Z(start_in[566]) );
  AND U25080 ( .A(start_reg[565]), .B(init), .Z(start_in[565]) );
  AND U25081 ( .A(start_reg[564]), .B(init), .Z(start_in[564]) );
  AND U25082 ( .A(start_reg[563]), .B(init), .Z(start_in[563]) );
  AND U25083 ( .A(start_reg[562]), .B(init), .Z(start_in[562]) );
  AND U25084 ( .A(start_reg[561]), .B(init), .Z(start_in[561]) );
  AND U25085 ( .A(start_reg[560]), .B(init), .Z(start_in[560]) );
  AND U25086 ( .A(start_reg[55]), .B(init), .Z(start_in[55]) );
  AND U25087 ( .A(start_reg[559]), .B(init), .Z(start_in[559]) );
  AND U25088 ( .A(start_reg[558]), .B(init), .Z(start_in[558]) );
  AND U25089 ( .A(start_reg[557]), .B(init), .Z(start_in[557]) );
  AND U25090 ( .A(start_reg[556]), .B(init), .Z(start_in[556]) );
  AND U25091 ( .A(start_reg[555]), .B(init), .Z(start_in[555]) );
  AND U25092 ( .A(start_reg[554]), .B(init), .Z(start_in[554]) );
  AND U25093 ( .A(start_reg[553]), .B(init), .Z(start_in[553]) );
  AND U25094 ( .A(start_reg[552]), .B(init), .Z(start_in[552]) );
  AND U25095 ( .A(start_reg[551]), .B(init), .Z(start_in[551]) );
  AND U25096 ( .A(start_reg[550]), .B(init), .Z(start_in[550]) );
  AND U25097 ( .A(start_reg[54]), .B(init), .Z(start_in[54]) );
  AND U25098 ( .A(start_reg[549]), .B(init), .Z(start_in[549]) );
  AND U25099 ( .A(start_reg[548]), .B(init), .Z(start_in[548]) );
  AND U25100 ( .A(start_reg[547]), .B(init), .Z(start_in[547]) );
  AND U25101 ( .A(start_reg[546]), .B(init), .Z(start_in[546]) );
  AND U25102 ( .A(start_reg[545]), .B(init), .Z(start_in[545]) );
  AND U25103 ( .A(start_reg[544]), .B(init), .Z(start_in[544]) );
  AND U25104 ( .A(start_reg[543]), .B(init), .Z(start_in[543]) );
  AND U25105 ( .A(start_reg[542]), .B(init), .Z(start_in[542]) );
  AND U25106 ( .A(start_reg[541]), .B(init), .Z(start_in[541]) );
  AND U25107 ( .A(start_reg[540]), .B(init), .Z(start_in[540]) );
  AND U25108 ( .A(start_reg[53]), .B(init), .Z(start_in[53]) );
  AND U25109 ( .A(start_reg[539]), .B(init), .Z(start_in[539]) );
  AND U25110 ( .A(start_reg[538]), .B(init), .Z(start_in[538]) );
  AND U25111 ( .A(start_reg[537]), .B(init), .Z(start_in[537]) );
  AND U25112 ( .A(start_reg[536]), .B(init), .Z(start_in[536]) );
  AND U25113 ( .A(start_reg[535]), .B(init), .Z(start_in[535]) );
  AND U25114 ( .A(start_reg[534]), .B(init), .Z(start_in[534]) );
  AND U25115 ( .A(start_reg[533]), .B(init), .Z(start_in[533]) );
  AND U25116 ( .A(start_reg[532]), .B(init), .Z(start_in[532]) );
  AND U25117 ( .A(start_reg[531]), .B(init), .Z(start_in[531]) );
  AND U25118 ( .A(start_reg[530]), .B(init), .Z(start_in[530]) );
  AND U25119 ( .A(start_reg[52]), .B(init), .Z(start_in[52]) );
  AND U25120 ( .A(start_reg[529]), .B(init), .Z(start_in[529]) );
  AND U25121 ( .A(start_reg[528]), .B(init), .Z(start_in[528]) );
  AND U25122 ( .A(start_reg[527]), .B(init), .Z(start_in[527]) );
  AND U25123 ( .A(start_reg[526]), .B(init), .Z(start_in[526]) );
  AND U25124 ( .A(start_reg[525]), .B(init), .Z(start_in[525]) );
  AND U25125 ( .A(start_reg[524]), .B(init), .Z(start_in[524]) );
  AND U25126 ( .A(start_reg[523]), .B(init), .Z(start_in[523]) );
  AND U25127 ( .A(start_reg[522]), .B(init), .Z(start_in[522]) );
  AND U25128 ( .A(start_reg[521]), .B(init), .Z(start_in[521]) );
  AND U25129 ( .A(start_reg[520]), .B(init), .Z(start_in[520]) );
  AND U25130 ( .A(start_reg[51]), .B(init), .Z(start_in[51]) );
  AND U25131 ( .A(start_reg[519]), .B(init), .Z(start_in[519]) );
  AND U25132 ( .A(start_reg[518]), .B(init), .Z(start_in[518]) );
  AND U25133 ( .A(start_reg[517]), .B(init), .Z(start_in[517]) );
  AND U25134 ( .A(start_reg[516]), .B(init), .Z(start_in[516]) );
  AND U25135 ( .A(start_reg[515]), .B(init), .Z(start_in[515]) );
  AND U25136 ( .A(start_reg[514]), .B(init), .Z(start_in[514]) );
  AND U25137 ( .A(start_reg[513]), .B(init), .Z(start_in[513]) );
  AND U25138 ( .A(start_reg[512]), .B(init), .Z(start_in[512]) );
  AND U25139 ( .A(start_reg[511]), .B(init), .Z(start_in[511]) );
  AND U25140 ( .A(start_reg[510]), .B(init), .Z(start_in[510]) );
  AND U25141 ( .A(start_reg[50]), .B(init), .Z(start_in[50]) );
  AND U25142 ( .A(start_reg[509]), .B(init), .Z(start_in[509]) );
  AND U25143 ( .A(start_reg[508]), .B(init), .Z(start_in[508]) );
  AND U25144 ( .A(start_reg[507]), .B(init), .Z(start_in[507]) );
  AND U25145 ( .A(start_reg[506]), .B(init), .Z(start_in[506]) );
  AND U25146 ( .A(start_reg[505]), .B(init), .Z(start_in[505]) );
  AND U25147 ( .A(start_reg[504]), .B(init), .Z(start_in[504]) );
  AND U25148 ( .A(start_reg[503]), .B(init), .Z(start_in[503]) );
  AND U25149 ( .A(start_reg[502]), .B(init), .Z(start_in[502]) );
  AND U25150 ( .A(start_reg[501]), .B(init), .Z(start_in[501]) );
  AND U25151 ( .A(start_reg[500]), .B(init), .Z(start_in[500]) );
  AND U25152 ( .A(start_reg[4]), .B(init), .Z(start_in[4]) );
  AND U25153 ( .A(start_reg[49]), .B(init), .Z(start_in[49]) );
  AND U25154 ( .A(start_reg[499]), .B(init), .Z(start_in[499]) );
  AND U25155 ( .A(start_reg[498]), .B(init), .Z(start_in[498]) );
  AND U25156 ( .A(start_reg[497]), .B(init), .Z(start_in[497]) );
  AND U25157 ( .A(start_reg[496]), .B(init), .Z(start_in[496]) );
  AND U25158 ( .A(start_reg[495]), .B(init), .Z(start_in[495]) );
  AND U25159 ( .A(start_reg[494]), .B(init), .Z(start_in[494]) );
  AND U25160 ( .A(start_reg[493]), .B(init), .Z(start_in[493]) );
  AND U25161 ( .A(start_reg[492]), .B(init), .Z(start_in[492]) );
  AND U25162 ( .A(start_reg[491]), .B(init), .Z(start_in[491]) );
  AND U25163 ( .A(start_reg[490]), .B(init), .Z(start_in[490]) );
  AND U25164 ( .A(start_reg[48]), .B(init), .Z(start_in[48]) );
  AND U25165 ( .A(start_reg[489]), .B(init), .Z(start_in[489]) );
  AND U25166 ( .A(start_reg[488]), .B(init), .Z(start_in[488]) );
  AND U25167 ( .A(start_reg[487]), .B(init), .Z(start_in[487]) );
  AND U25168 ( .A(start_reg[486]), .B(init), .Z(start_in[486]) );
  AND U25169 ( .A(start_reg[485]), .B(init), .Z(start_in[485]) );
  AND U25170 ( .A(start_reg[484]), .B(init), .Z(start_in[484]) );
  AND U25171 ( .A(start_reg[483]), .B(init), .Z(start_in[483]) );
  AND U25172 ( .A(start_reg[482]), .B(init), .Z(start_in[482]) );
  AND U25173 ( .A(start_reg[481]), .B(init), .Z(start_in[481]) );
  AND U25174 ( .A(start_reg[480]), .B(init), .Z(start_in[480]) );
  AND U25175 ( .A(start_reg[47]), .B(init), .Z(start_in[47]) );
  AND U25176 ( .A(start_reg[479]), .B(init), .Z(start_in[479]) );
  AND U25177 ( .A(start_reg[478]), .B(init), .Z(start_in[478]) );
  AND U25178 ( .A(start_reg[477]), .B(init), .Z(start_in[477]) );
  AND U25179 ( .A(start_reg[476]), .B(init), .Z(start_in[476]) );
  AND U25180 ( .A(start_reg[475]), .B(init), .Z(start_in[475]) );
  AND U25181 ( .A(start_reg[474]), .B(init), .Z(start_in[474]) );
  AND U25182 ( .A(start_reg[473]), .B(init), .Z(start_in[473]) );
  AND U25183 ( .A(start_reg[472]), .B(init), .Z(start_in[472]) );
  AND U25184 ( .A(start_reg[471]), .B(init), .Z(start_in[471]) );
  AND U25185 ( .A(start_reg[470]), .B(init), .Z(start_in[470]) );
  AND U25186 ( .A(start_reg[46]), .B(init), .Z(start_in[46]) );
  AND U25187 ( .A(start_reg[469]), .B(init), .Z(start_in[469]) );
  AND U25188 ( .A(start_reg[468]), .B(init), .Z(start_in[468]) );
  AND U25189 ( .A(start_reg[467]), .B(init), .Z(start_in[467]) );
  AND U25190 ( .A(start_reg[466]), .B(init), .Z(start_in[466]) );
  AND U25191 ( .A(start_reg[465]), .B(init), .Z(start_in[465]) );
  AND U25192 ( .A(start_reg[464]), .B(init), .Z(start_in[464]) );
  AND U25193 ( .A(start_reg[463]), .B(init), .Z(start_in[463]) );
  AND U25194 ( .A(start_reg[462]), .B(init), .Z(start_in[462]) );
  AND U25195 ( .A(start_reg[461]), .B(init), .Z(start_in[461]) );
  AND U25196 ( .A(start_reg[460]), .B(init), .Z(start_in[460]) );
  AND U25197 ( .A(start_reg[45]), .B(init), .Z(start_in[45]) );
  AND U25198 ( .A(start_reg[459]), .B(init), .Z(start_in[459]) );
  AND U25199 ( .A(start_reg[458]), .B(init), .Z(start_in[458]) );
  AND U25200 ( .A(start_reg[457]), .B(init), .Z(start_in[457]) );
  AND U25201 ( .A(start_reg[456]), .B(init), .Z(start_in[456]) );
  AND U25202 ( .A(start_reg[455]), .B(init), .Z(start_in[455]) );
  AND U25203 ( .A(start_reg[454]), .B(init), .Z(start_in[454]) );
  AND U25204 ( .A(start_reg[453]), .B(init), .Z(start_in[453]) );
  AND U25205 ( .A(start_reg[452]), .B(init), .Z(start_in[452]) );
  AND U25206 ( .A(start_reg[451]), .B(init), .Z(start_in[451]) );
  AND U25207 ( .A(start_reg[450]), .B(init), .Z(start_in[450]) );
  AND U25208 ( .A(start_reg[44]), .B(init), .Z(start_in[44]) );
  AND U25209 ( .A(start_reg[449]), .B(init), .Z(start_in[449]) );
  AND U25210 ( .A(start_reg[448]), .B(init), .Z(start_in[448]) );
  AND U25211 ( .A(start_reg[447]), .B(init), .Z(start_in[447]) );
  AND U25212 ( .A(start_reg[446]), .B(init), .Z(start_in[446]) );
  AND U25213 ( .A(start_reg[445]), .B(init), .Z(start_in[445]) );
  AND U25214 ( .A(start_reg[444]), .B(init), .Z(start_in[444]) );
  AND U25215 ( .A(start_reg[443]), .B(init), .Z(start_in[443]) );
  AND U25216 ( .A(start_reg[442]), .B(init), .Z(start_in[442]) );
  AND U25217 ( .A(start_reg[441]), .B(init), .Z(start_in[441]) );
  AND U25218 ( .A(start_reg[440]), .B(init), .Z(start_in[440]) );
  AND U25219 ( .A(start_reg[43]), .B(init), .Z(start_in[43]) );
  AND U25220 ( .A(start_reg[439]), .B(init), .Z(start_in[439]) );
  AND U25221 ( .A(start_reg[438]), .B(init), .Z(start_in[438]) );
  AND U25222 ( .A(start_reg[437]), .B(init), .Z(start_in[437]) );
  AND U25223 ( .A(start_reg[436]), .B(init), .Z(start_in[436]) );
  AND U25224 ( .A(start_reg[435]), .B(init), .Z(start_in[435]) );
  AND U25225 ( .A(start_reg[434]), .B(init), .Z(start_in[434]) );
  AND U25226 ( .A(start_reg[433]), .B(init), .Z(start_in[433]) );
  AND U25227 ( .A(start_reg[432]), .B(init), .Z(start_in[432]) );
  AND U25228 ( .A(start_reg[431]), .B(init), .Z(start_in[431]) );
  AND U25229 ( .A(start_reg[430]), .B(init), .Z(start_in[430]) );
  AND U25230 ( .A(start_reg[42]), .B(init), .Z(start_in[42]) );
  AND U25231 ( .A(start_reg[429]), .B(init), .Z(start_in[429]) );
  AND U25232 ( .A(start_reg[428]), .B(init), .Z(start_in[428]) );
  AND U25233 ( .A(start_reg[427]), .B(init), .Z(start_in[427]) );
  AND U25234 ( .A(start_reg[426]), .B(init), .Z(start_in[426]) );
  AND U25235 ( .A(start_reg[425]), .B(init), .Z(start_in[425]) );
  AND U25236 ( .A(start_reg[424]), .B(init), .Z(start_in[424]) );
  AND U25237 ( .A(start_reg[423]), .B(init), .Z(start_in[423]) );
  AND U25238 ( .A(start_reg[422]), .B(init), .Z(start_in[422]) );
  AND U25239 ( .A(start_reg[421]), .B(init), .Z(start_in[421]) );
  AND U25240 ( .A(start_reg[420]), .B(init), .Z(start_in[420]) );
  AND U25241 ( .A(start_reg[41]), .B(init), .Z(start_in[41]) );
  AND U25242 ( .A(start_reg[419]), .B(init), .Z(start_in[419]) );
  AND U25243 ( .A(start_reg[418]), .B(init), .Z(start_in[418]) );
  AND U25244 ( .A(start_reg[417]), .B(init), .Z(start_in[417]) );
  AND U25245 ( .A(start_reg[416]), .B(init), .Z(start_in[416]) );
  AND U25246 ( .A(start_reg[415]), .B(init), .Z(start_in[415]) );
  AND U25247 ( .A(start_reg[414]), .B(init), .Z(start_in[414]) );
  AND U25248 ( .A(start_reg[413]), .B(init), .Z(start_in[413]) );
  AND U25249 ( .A(start_reg[412]), .B(init), .Z(start_in[412]) );
  AND U25250 ( .A(start_reg[411]), .B(init), .Z(start_in[411]) );
  AND U25251 ( .A(start_reg[410]), .B(init), .Z(start_in[410]) );
  AND U25252 ( .A(start_reg[40]), .B(init), .Z(start_in[40]) );
  AND U25253 ( .A(start_reg[409]), .B(init), .Z(start_in[409]) );
  AND U25254 ( .A(start_reg[408]), .B(init), .Z(start_in[408]) );
  AND U25255 ( .A(start_reg[407]), .B(init), .Z(start_in[407]) );
  AND U25256 ( .A(start_reg[406]), .B(init), .Z(start_in[406]) );
  AND U25257 ( .A(start_reg[405]), .B(init), .Z(start_in[405]) );
  AND U25258 ( .A(start_reg[404]), .B(init), .Z(start_in[404]) );
  AND U25259 ( .A(start_reg[403]), .B(init), .Z(start_in[403]) );
  AND U25260 ( .A(start_reg[402]), .B(init), .Z(start_in[402]) );
  AND U25261 ( .A(start_reg[401]), .B(init), .Z(start_in[401]) );
  AND U25262 ( .A(start_reg[400]), .B(init), .Z(start_in[400]) );
  AND U25263 ( .A(start_reg[3]), .B(init), .Z(start_in[3]) );
  AND U25264 ( .A(start_reg[39]), .B(init), .Z(start_in[39]) );
  AND U25265 ( .A(start_reg[399]), .B(init), .Z(start_in[399]) );
  AND U25266 ( .A(start_reg[398]), .B(init), .Z(start_in[398]) );
  AND U25267 ( .A(start_reg[397]), .B(init), .Z(start_in[397]) );
  AND U25268 ( .A(start_reg[396]), .B(init), .Z(start_in[396]) );
  AND U25269 ( .A(start_reg[395]), .B(init), .Z(start_in[395]) );
  AND U25270 ( .A(start_reg[394]), .B(init), .Z(start_in[394]) );
  AND U25271 ( .A(start_reg[393]), .B(init), .Z(start_in[393]) );
  AND U25272 ( .A(start_reg[392]), .B(init), .Z(start_in[392]) );
  AND U25273 ( .A(start_reg[391]), .B(init), .Z(start_in[391]) );
  AND U25274 ( .A(start_reg[390]), .B(init), .Z(start_in[390]) );
  AND U25275 ( .A(start_reg[38]), .B(init), .Z(start_in[38]) );
  AND U25276 ( .A(start_reg[389]), .B(init), .Z(start_in[389]) );
  AND U25277 ( .A(start_reg[388]), .B(init), .Z(start_in[388]) );
  AND U25278 ( .A(start_reg[387]), .B(init), .Z(start_in[387]) );
  AND U25279 ( .A(start_reg[386]), .B(init), .Z(start_in[386]) );
  AND U25280 ( .A(start_reg[385]), .B(init), .Z(start_in[385]) );
  AND U25281 ( .A(start_reg[384]), .B(init), .Z(start_in[384]) );
  AND U25282 ( .A(start_reg[383]), .B(init), .Z(start_in[383]) );
  AND U25283 ( .A(start_reg[382]), .B(init), .Z(start_in[382]) );
  AND U25284 ( .A(start_reg[381]), .B(init), .Z(start_in[381]) );
  AND U25285 ( .A(start_reg[380]), .B(init), .Z(start_in[380]) );
  AND U25286 ( .A(start_reg[37]), .B(init), .Z(start_in[37]) );
  AND U25287 ( .A(start_reg[379]), .B(init), .Z(start_in[379]) );
  AND U25288 ( .A(start_reg[378]), .B(init), .Z(start_in[378]) );
  AND U25289 ( .A(start_reg[377]), .B(init), .Z(start_in[377]) );
  AND U25290 ( .A(start_reg[376]), .B(init), .Z(start_in[376]) );
  AND U25291 ( .A(start_reg[375]), .B(init), .Z(start_in[375]) );
  AND U25292 ( .A(start_reg[374]), .B(init), .Z(start_in[374]) );
  AND U25293 ( .A(start_reg[373]), .B(init), .Z(start_in[373]) );
  AND U25294 ( .A(start_reg[372]), .B(init), .Z(start_in[372]) );
  AND U25295 ( .A(start_reg[371]), .B(init), .Z(start_in[371]) );
  AND U25296 ( .A(start_reg[370]), .B(init), .Z(start_in[370]) );
  AND U25297 ( .A(start_reg[36]), .B(init), .Z(start_in[36]) );
  AND U25298 ( .A(start_reg[369]), .B(init), .Z(start_in[369]) );
  AND U25299 ( .A(start_reg[368]), .B(init), .Z(start_in[368]) );
  AND U25300 ( .A(start_reg[367]), .B(init), .Z(start_in[367]) );
  AND U25301 ( .A(start_reg[366]), .B(init), .Z(start_in[366]) );
  AND U25302 ( .A(start_reg[365]), .B(init), .Z(start_in[365]) );
  AND U25303 ( .A(start_reg[364]), .B(init), .Z(start_in[364]) );
  AND U25304 ( .A(start_reg[363]), .B(init), .Z(start_in[363]) );
  AND U25305 ( .A(start_reg[362]), .B(init), .Z(start_in[362]) );
  AND U25306 ( .A(start_reg[361]), .B(init), .Z(start_in[361]) );
  AND U25307 ( .A(start_reg[360]), .B(init), .Z(start_in[360]) );
  AND U25308 ( .A(start_reg[35]), .B(init), .Z(start_in[35]) );
  AND U25309 ( .A(start_reg[359]), .B(init), .Z(start_in[359]) );
  AND U25310 ( .A(start_reg[358]), .B(init), .Z(start_in[358]) );
  AND U25311 ( .A(start_reg[357]), .B(init), .Z(start_in[357]) );
  AND U25312 ( .A(start_reg[356]), .B(init), .Z(start_in[356]) );
  AND U25313 ( .A(start_reg[355]), .B(init), .Z(start_in[355]) );
  AND U25314 ( .A(start_reg[354]), .B(init), .Z(start_in[354]) );
  AND U25315 ( .A(start_reg[353]), .B(init), .Z(start_in[353]) );
  AND U25316 ( .A(start_reg[352]), .B(init), .Z(start_in[352]) );
  AND U25317 ( .A(start_reg[351]), .B(init), .Z(start_in[351]) );
  AND U25318 ( .A(start_reg[350]), .B(init), .Z(start_in[350]) );
  AND U25319 ( .A(start_reg[34]), .B(init), .Z(start_in[34]) );
  AND U25320 ( .A(start_reg[349]), .B(init), .Z(start_in[349]) );
  AND U25321 ( .A(start_reg[348]), .B(init), .Z(start_in[348]) );
  AND U25322 ( .A(start_reg[347]), .B(init), .Z(start_in[347]) );
  AND U25323 ( .A(start_reg[346]), .B(init), .Z(start_in[346]) );
  AND U25324 ( .A(start_reg[345]), .B(init), .Z(start_in[345]) );
  AND U25325 ( .A(start_reg[344]), .B(init), .Z(start_in[344]) );
  AND U25326 ( .A(start_reg[343]), .B(init), .Z(start_in[343]) );
  AND U25327 ( .A(start_reg[342]), .B(init), .Z(start_in[342]) );
  AND U25328 ( .A(start_reg[341]), .B(init), .Z(start_in[341]) );
  AND U25329 ( .A(start_reg[340]), .B(init), .Z(start_in[340]) );
  AND U25330 ( .A(start_reg[33]), .B(init), .Z(start_in[33]) );
  AND U25331 ( .A(start_reg[339]), .B(init), .Z(start_in[339]) );
  AND U25332 ( .A(start_reg[338]), .B(init), .Z(start_in[338]) );
  AND U25333 ( .A(start_reg[337]), .B(init), .Z(start_in[337]) );
  AND U25334 ( .A(start_reg[336]), .B(init), .Z(start_in[336]) );
  AND U25335 ( .A(start_reg[335]), .B(init), .Z(start_in[335]) );
  AND U25336 ( .A(start_reg[334]), .B(init), .Z(start_in[334]) );
  AND U25337 ( .A(start_reg[333]), .B(init), .Z(start_in[333]) );
  AND U25338 ( .A(start_reg[332]), .B(init), .Z(start_in[332]) );
  AND U25339 ( .A(start_reg[331]), .B(init), .Z(start_in[331]) );
  AND U25340 ( .A(start_reg[330]), .B(init), .Z(start_in[330]) );
  AND U25341 ( .A(start_reg[32]), .B(init), .Z(start_in[32]) );
  AND U25342 ( .A(start_reg[329]), .B(init), .Z(start_in[329]) );
  AND U25343 ( .A(start_reg[328]), .B(init), .Z(start_in[328]) );
  AND U25344 ( .A(start_reg[327]), .B(init), .Z(start_in[327]) );
  AND U25345 ( .A(start_reg[326]), .B(init), .Z(start_in[326]) );
  AND U25346 ( .A(start_reg[325]), .B(init), .Z(start_in[325]) );
  AND U25347 ( .A(start_reg[324]), .B(init), .Z(start_in[324]) );
  AND U25348 ( .A(start_reg[323]), .B(init), .Z(start_in[323]) );
  AND U25349 ( .A(start_reg[322]), .B(init), .Z(start_in[322]) );
  AND U25350 ( .A(start_reg[321]), .B(init), .Z(start_in[321]) );
  AND U25351 ( .A(start_reg[320]), .B(init), .Z(start_in[320]) );
  AND U25352 ( .A(start_reg[31]), .B(init), .Z(start_in[31]) );
  AND U25353 ( .A(start_reg[319]), .B(init), .Z(start_in[319]) );
  AND U25354 ( .A(start_reg[318]), .B(init), .Z(start_in[318]) );
  AND U25355 ( .A(start_reg[317]), .B(init), .Z(start_in[317]) );
  AND U25356 ( .A(start_reg[316]), .B(init), .Z(start_in[316]) );
  AND U25357 ( .A(start_reg[315]), .B(init), .Z(start_in[315]) );
  AND U25358 ( .A(start_reg[314]), .B(init), .Z(start_in[314]) );
  AND U25359 ( .A(start_reg[313]), .B(init), .Z(start_in[313]) );
  AND U25360 ( .A(start_reg[312]), .B(init), .Z(start_in[312]) );
  AND U25361 ( .A(start_reg[311]), .B(init), .Z(start_in[311]) );
  AND U25362 ( .A(start_reg[310]), .B(init), .Z(start_in[310]) );
  AND U25363 ( .A(start_reg[30]), .B(init), .Z(start_in[30]) );
  AND U25364 ( .A(start_reg[309]), .B(init), .Z(start_in[309]) );
  AND U25365 ( .A(start_reg[308]), .B(init), .Z(start_in[308]) );
  AND U25366 ( .A(start_reg[307]), .B(init), .Z(start_in[307]) );
  AND U25367 ( .A(start_reg[306]), .B(init), .Z(start_in[306]) );
  AND U25368 ( .A(start_reg[305]), .B(init), .Z(start_in[305]) );
  AND U25369 ( .A(start_reg[304]), .B(init), .Z(start_in[304]) );
  AND U25370 ( .A(start_reg[303]), .B(init), .Z(start_in[303]) );
  AND U25371 ( .A(start_reg[302]), .B(init), .Z(start_in[302]) );
  AND U25372 ( .A(start_reg[301]), .B(init), .Z(start_in[301]) );
  AND U25373 ( .A(start_reg[300]), .B(init), .Z(start_in[300]) );
  AND U25374 ( .A(start_reg[2]), .B(init), .Z(start_in[2]) );
  AND U25375 ( .A(start_reg[29]), .B(init), .Z(start_in[29]) );
  AND U25376 ( .A(start_reg[299]), .B(init), .Z(start_in[299]) );
  AND U25377 ( .A(start_reg[298]), .B(init), .Z(start_in[298]) );
  AND U25378 ( .A(start_reg[297]), .B(init), .Z(start_in[297]) );
  AND U25379 ( .A(start_reg[296]), .B(init), .Z(start_in[296]) );
  AND U25380 ( .A(start_reg[295]), .B(init), .Z(start_in[295]) );
  AND U25381 ( .A(start_reg[294]), .B(init), .Z(start_in[294]) );
  AND U25382 ( .A(start_reg[293]), .B(init), .Z(start_in[293]) );
  AND U25383 ( .A(start_reg[292]), .B(init), .Z(start_in[292]) );
  AND U25384 ( .A(start_reg[291]), .B(init), .Z(start_in[291]) );
  AND U25385 ( .A(start_reg[290]), .B(init), .Z(start_in[290]) );
  AND U25386 ( .A(start_reg[28]), .B(init), .Z(start_in[28]) );
  AND U25387 ( .A(start_reg[289]), .B(init), .Z(start_in[289]) );
  AND U25388 ( .A(start_reg[288]), .B(init), .Z(start_in[288]) );
  AND U25389 ( .A(start_reg[287]), .B(init), .Z(start_in[287]) );
  AND U25390 ( .A(start_reg[286]), .B(init), .Z(start_in[286]) );
  AND U25391 ( .A(start_reg[285]), .B(init), .Z(start_in[285]) );
  AND U25392 ( .A(start_reg[284]), .B(init), .Z(start_in[284]) );
  AND U25393 ( .A(start_reg[283]), .B(init), .Z(start_in[283]) );
  AND U25394 ( .A(start_reg[282]), .B(init), .Z(start_in[282]) );
  AND U25395 ( .A(start_reg[281]), .B(init), .Z(start_in[281]) );
  AND U25396 ( .A(start_reg[280]), .B(init), .Z(start_in[280]) );
  AND U25397 ( .A(start_reg[27]), .B(init), .Z(start_in[27]) );
  AND U25398 ( .A(start_reg[279]), .B(init), .Z(start_in[279]) );
  AND U25399 ( .A(start_reg[278]), .B(init), .Z(start_in[278]) );
  AND U25400 ( .A(start_reg[277]), .B(init), .Z(start_in[277]) );
  AND U25401 ( .A(start_reg[276]), .B(init), .Z(start_in[276]) );
  AND U25402 ( .A(start_reg[275]), .B(init), .Z(start_in[275]) );
  AND U25403 ( .A(start_reg[274]), .B(init), .Z(start_in[274]) );
  AND U25404 ( .A(start_reg[273]), .B(init), .Z(start_in[273]) );
  AND U25405 ( .A(start_reg[272]), .B(init), .Z(start_in[272]) );
  AND U25406 ( .A(start_reg[271]), .B(init), .Z(start_in[271]) );
  AND U25407 ( .A(start_reg[270]), .B(init), .Z(start_in[270]) );
  AND U25408 ( .A(start_reg[26]), .B(init), .Z(start_in[26]) );
  AND U25409 ( .A(start_reg[269]), .B(init), .Z(start_in[269]) );
  AND U25410 ( .A(start_reg[268]), .B(init), .Z(start_in[268]) );
  AND U25411 ( .A(start_reg[267]), .B(init), .Z(start_in[267]) );
  AND U25412 ( .A(start_reg[266]), .B(init), .Z(start_in[266]) );
  AND U25413 ( .A(start_reg[265]), .B(init), .Z(start_in[265]) );
  AND U25414 ( .A(start_reg[264]), .B(init), .Z(start_in[264]) );
  AND U25415 ( .A(start_reg[263]), .B(init), .Z(start_in[263]) );
  AND U25416 ( .A(start_reg[262]), .B(init), .Z(start_in[262]) );
  AND U25417 ( .A(start_reg[261]), .B(init), .Z(start_in[261]) );
  AND U25418 ( .A(start_reg[260]), .B(init), .Z(start_in[260]) );
  AND U25419 ( .A(start_reg[25]), .B(init), .Z(start_in[25]) );
  AND U25420 ( .A(start_reg[259]), .B(init), .Z(start_in[259]) );
  AND U25421 ( .A(start_reg[258]), .B(init), .Z(start_in[258]) );
  AND U25422 ( .A(start_reg[257]), .B(init), .Z(start_in[257]) );
  AND U25423 ( .A(start_reg[256]), .B(init), .Z(start_in[256]) );
  AND U25424 ( .A(start_reg[255]), .B(init), .Z(start_in[255]) );
  AND U25425 ( .A(start_reg[254]), .B(init), .Z(start_in[254]) );
  AND U25426 ( .A(start_reg[253]), .B(init), .Z(start_in[253]) );
  AND U25427 ( .A(start_reg[252]), .B(init), .Z(start_in[252]) );
  AND U25428 ( .A(start_reg[251]), .B(init), .Z(start_in[251]) );
  AND U25429 ( .A(start_reg[250]), .B(init), .Z(start_in[250]) );
  AND U25430 ( .A(start_reg[24]), .B(init), .Z(start_in[24]) );
  AND U25431 ( .A(start_reg[249]), .B(init), .Z(start_in[249]) );
  AND U25432 ( .A(start_reg[248]), .B(init), .Z(start_in[248]) );
  AND U25433 ( .A(start_reg[247]), .B(init), .Z(start_in[247]) );
  AND U25434 ( .A(start_reg[246]), .B(init), .Z(start_in[246]) );
  AND U25435 ( .A(start_reg[245]), .B(init), .Z(start_in[245]) );
  AND U25436 ( .A(start_reg[244]), .B(init), .Z(start_in[244]) );
  AND U25437 ( .A(start_reg[243]), .B(init), .Z(start_in[243]) );
  AND U25438 ( .A(start_reg[242]), .B(init), .Z(start_in[242]) );
  AND U25439 ( .A(start_reg[241]), .B(init), .Z(start_in[241]) );
  AND U25440 ( .A(start_reg[240]), .B(init), .Z(start_in[240]) );
  AND U25441 ( .A(start_reg[23]), .B(init), .Z(start_in[23]) );
  AND U25442 ( .A(start_reg[239]), .B(init), .Z(start_in[239]) );
  AND U25443 ( .A(start_reg[238]), .B(init), .Z(start_in[238]) );
  AND U25444 ( .A(start_reg[237]), .B(init), .Z(start_in[237]) );
  AND U25445 ( .A(start_reg[236]), .B(init), .Z(start_in[236]) );
  AND U25446 ( .A(start_reg[235]), .B(init), .Z(start_in[235]) );
  AND U25447 ( .A(start_reg[234]), .B(init), .Z(start_in[234]) );
  AND U25448 ( .A(start_reg[233]), .B(init), .Z(start_in[233]) );
  AND U25449 ( .A(start_reg[232]), .B(init), .Z(start_in[232]) );
  AND U25450 ( .A(start_reg[231]), .B(init), .Z(start_in[231]) );
  AND U25451 ( .A(start_reg[230]), .B(init), .Z(start_in[230]) );
  AND U25452 ( .A(start_reg[22]), .B(init), .Z(start_in[22]) );
  AND U25453 ( .A(start_reg[229]), .B(init), .Z(start_in[229]) );
  AND U25454 ( .A(start_reg[228]), .B(init), .Z(start_in[228]) );
  AND U25455 ( .A(start_reg[227]), .B(init), .Z(start_in[227]) );
  AND U25456 ( .A(start_reg[226]), .B(init), .Z(start_in[226]) );
  AND U25457 ( .A(start_reg[225]), .B(init), .Z(start_in[225]) );
  AND U25458 ( .A(start_reg[224]), .B(init), .Z(start_in[224]) );
  AND U25459 ( .A(start_reg[223]), .B(init), .Z(start_in[223]) );
  AND U25460 ( .A(start_reg[222]), .B(init), .Z(start_in[222]) );
  AND U25461 ( .A(start_reg[221]), .B(init), .Z(start_in[221]) );
  AND U25462 ( .A(start_reg[220]), .B(init), .Z(start_in[220]) );
  AND U25463 ( .A(start_reg[21]), .B(init), .Z(start_in[21]) );
  AND U25464 ( .A(start_reg[219]), .B(init), .Z(start_in[219]) );
  AND U25465 ( .A(start_reg[218]), .B(init), .Z(start_in[218]) );
  AND U25466 ( .A(start_reg[217]), .B(init), .Z(start_in[217]) );
  AND U25467 ( .A(start_reg[216]), .B(init), .Z(start_in[216]) );
  AND U25468 ( .A(start_reg[215]), .B(init), .Z(start_in[215]) );
  AND U25469 ( .A(start_reg[214]), .B(init), .Z(start_in[214]) );
  AND U25470 ( .A(start_reg[213]), .B(init), .Z(start_in[213]) );
  AND U25471 ( .A(start_reg[212]), .B(init), .Z(start_in[212]) );
  AND U25472 ( .A(start_reg[211]), .B(init), .Z(start_in[211]) );
  AND U25473 ( .A(start_reg[210]), .B(init), .Z(start_in[210]) );
  AND U25474 ( .A(start_reg[20]), .B(init), .Z(start_in[20]) );
  AND U25475 ( .A(start_reg[209]), .B(init), .Z(start_in[209]) );
  AND U25476 ( .A(start_reg[208]), .B(init), .Z(start_in[208]) );
  AND U25477 ( .A(start_reg[207]), .B(init), .Z(start_in[207]) );
  AND U25478 ( .A(start_reg[206]), .B(init), .Z(start_in[206]) );
  AND U25479 ( .A(start_reg[205]), .B(init), .Z(start_in[205]) );
  AND U25480 ( .A(start_reg[204]), .B(init), .Z(start_in[204]) );
  AND U25481 ( .A(start_reg[203]), .B(init), .Z(start_in[203]) );
  AND U25482 ( .A(start_reg[202]), .B(init), .Z(start_in[202]) );
  AND U25483 ( .A(start_reg[201]), .B(init), .Z(start_in[201]) );
  AND U25484 ( .A(start_reg[200]), .B(init), .Z(start_in[200]) );
  AND U25485 ( .A(start_reg[1]), .B(init), .Z(start_in[1]) );
  AND U25486 ( .A(start_reg[19]), .B(init), .Z(start_in[19]) );
  AND U25487 ( .A(start_reg[199]), .B(init), .Z(start_in[199]) );
  AND U25488 ( .A(start_reg[198]), .B(init), .Z(start_in[198]) );
  AND U25489 ( .A(start_reg[197]), .B(init), .Z(start_in[197]) );
  AND U25490 ( .A(start_reg[196]), .B(init), .Z(start_in[196]) );
  AND U25491 ( .A(start_reg[195]), .B(init), .Z(start_in[195]) );
  AND U25492 ( .A(start_reg[194]), .B(init), .Z(start_in[194]) );
  AND U25493 ( .A(start_reg[193]), .B(init), .Z(start_in[193]) );
  AND U25494 ( .A(start_reg[192]), .B(init), .Z(start_in[192]) );
  AND U25495 ( .A(start_reg[191]), .B(init), .Z(start_in[191]) );
  AND U25496 ( .A(start_reg[190]), .B(init), .Z(start_in[190]) );
  AND U25497 ( .A(start_reg[18]), .B(init), .Z(start_in[18]) );
  AND U25498 ( .A(start_reg[189]), .B(init), .Z(start_in[189]) );
  AND U25499 ( .A(start_reg[188]), .B(init), .Z(start_in[188]) );
  AND U25500 ( .A(start_reg[187]), .B(init), .Z(start_in[187]) );
  AND U25501 ( .A(start_reg[186]), .B(init), .Z(start_in[186]) );
  AND U25502 ( .A(start_reg[185]), .B(init), .Z(start_in[185]) );
  AND U25503 ( .A(start_reg[184]), .B(init), .Z(start_in[184]) );
  AND U25504 ( .A(start_reg[183]), .B(init), .Z(start_in[183]) );
  AND U25505 ( .A(start_reg[182]), .B(init), .Z(start_in[182]) );
  AND U25506 ( .A(start_reg[181]), .B(init), .Z(start_in[181]) );
  AND U25507 ( .A(start_reg[180]), .B(init), .Z(start_in[180]) );
  AND U25508 ( .A(start_reg[17]), .B(init), .Z(start_in[17]) );
  AND U25509 ( .A(start_reg[179]), .B(init), .Z(start_in[179]) );
  AND U25510 ( .A(start_reg[178]), .B(init), .Z(start_in[178]) );
  AND U25511 ( .A(start_reg[177]), .B(init), .Z(start_in[177]) );
  AND U25512 ( .A(start_reg[176]), .B(init), .Z(start_in[176]) );
  AND U25513 ( .A(start_reg[175]), .B(init), .Z(start_in[175]) );
  AND U25514 ( .A(start_reg[174]), .B(init), .Z(start_in[174]) );
  AND U25515 ( .A(start_reg[173]), .B(init), .Z(start_in[173]) );
  AND U25516 ( .A(start_reg[172]), .B(init), .Z(start_in[172]) );
  AND U25517 ( .A(start_reg[171]), .B(init), .Z(start_in[171]) );
  AND U25518 ( .A(start_reg[170]), .B(init), .Z(start_in[170]) );
  AND U25519 ( .A(start_reg[16]), .B(init), .Z(start_in[16]) );
  AND U25520 ( .A(start_reg[169]), .B(init), .Z(start_in[169]) );
  AND U25521 ( .A(start_reg[168]), .B(init), .Z(start_in[168]) );
  AND U25522 ( .A(start_reg[167]), .B(init), .Z(start_in[167]) );
  AND U25523 ( .A(start_reg[166]), .B(init), .Z(start_in[166]) );
  AND U25524 ( .A(start_reg[165]), .B(init), .Z(start_in[165]) );
  AND U25525 ( .A(start_reg[164]), .B(init), .Z(start_in[164]) );
  AND U25526 ( .A(start_reg[163]), .B(init), .Z(start_in[163]) );
  AND U25527 ( .A(start_reg[162]), .B(init), .Z(start_in[162]) );
  AND U25528 ( .A(start_reg[161]), .B(init), .Z(start_in[161]) );
  AND U25529 ( .A(start_reg[160]), .B(init), .Z(start_in[160]) );
  AND U25530 ( .A(start_reg[15]), .B(init), .Z(start_in[15]) );
  AND U25531 ( .A(start_reg[159]), .B(init), .Z(start_in[159]) );
  AND U25532 ( .A(start_reg[158]), .B(init), .Z(start_in[158]) );
  AND U25533 ( .A(start_reg[157]), .B(init), .Z(start_in[157]) );
  AND U25534 ( .A(start_reg[156]), .B(init), .Z(start_in[156]) );
  AND U25535 ( .A(start_reg[155]), .B(init), .Z(start_in[155]) );
  AND U25536 ( .A(start_reg[154]), .B(init), .Z(start_in[154]) );
  AND U25537 ( .A(start_reg[153]), .B(init), .Z(start_in[153]) );
  AND U25538 ( .A(start_reg[152]), .B(init), .Z(start_in[152]) );
  AND U25539 ( .A(start_reg[151]), .B(init), .Z(start_in[151]) );
  AND U25540 ( .A(start_reg[150]), .B(init), .Z(start_in[150]) );
  AND U25541 ( .A(start_reg[14]), .B(init), .Z(start_in[14]) );
  AND U25542 ( .A(start_reg[149]), .B(init), .Z(start_in[149]) );
  AND U25543 ( .A(start_reg[148]), .B(init), .Z(start_in[148]) );
  AND U25544 ( .A(start_reg[147]), .B(init), .Z(start_in[147]) );
  AND U25545 ( .A(start_reg[146]), .B(init), .Z(start_in[146]) );
  AND U25546 ( .A(start_reg[145]), .B(init), .Z(start_in[145]) );
  AND U25547 ( .A(start_reg[144]), .B(init), .Z(start_in[144]) );
  AND U25548 ( .A(start_reg[143]), .B(init), .Z(start_in[143]) );
  AND U25549 ( .A(start_reg[142]), .B(init), .Z(start_in[142]) );
  AND U25550 ( .A(start_reg[141]), .B(init), .Z(start_in[141]) );
  AND U25551 ( .A(start_reg[140]), .B(init), .Z(start_in[140]) );
  AND U25552 ( .A(start_reg[13]), .B(init), .Z(start_in[13]) );
  AND U25553 ( .A(start_reg[139]), .B(init), .Z(start_in[139]) );
  AND U25554 ( .A(start_reg[138]), .B(init), .Z(start_in[138]) );
  AND U25555 ( .A(start_reg[137]), .B(init), .Z(start_in[137]) );
  AND U25556 ( .A(start_reg[136]), .B(init), .Z(start_in[136]) );
  AND U25557 ( .A(start_reg[135]), .B(init), .Z(start_in[135]) );
  AND U25558 ( .A(start_reg[134]), .B(init), .Z(start_in[134]) );
  AND U25559 ( .A(start_reg[133]), .B(init), .Z(start_in[133]) );
  AND U25560 ( .A(start_reg[132]), .B(init), .Z(start_in[132]) );
  AND U25561 ( .A(start_reg[131]), .B(init), .Z(start_in[131]) );
  AND U25562 ( .A(start_reg[130]), .B(init), .Z(start_in[130]) );
  AND U25563 ( .A(start_reg[12]), .B(init), .Z(start_in[12]) );
  AND U25564 ( .A(start_reg[129]), .B(init), .Z(start_in[129]) );
  AND U25565 ( .A(start_reg[128]), .B(init), .Z(start_in[128]) );
  AND U25566 ( .A(start_reg[127]), .B(init), .Z(start_in[127]) );
  AND U25567 ( .A(start_reg[126]), .B(init), .Z(start_in[126]) );
  AND U25568 ( .A(start_reg[125]), .B(init), .Z(start_in[125]) );
  AND U25569 ( .A(start_reg[124]), .B(init), .Z(start_in[124]) );
  AND U25570 ( .A(start_reg[123]), .B(init), .Z(start_in[123]) );
  AND U25571 ( .A(start_reg[122]), .B(init), .Z(start_in[122]) );
  AND U25572 ( .A(start_reg[121]), .B(init), .Z(start_in[121]) );
  AND U25573 ( .A(start_reg[120]), .B(init), .Z(start_in[120]) );
  AND U25574 ( .A(start_reg[11]), .B(init), .Z(start_in[11]) );
  AND U25575 ( .A(start_reg[119]), .B(init), .Z(start_in[119]) );
  AND U25576 ( .A(start_reg[118]), .B(init), .Z(start_in[118]) );
  AND U25577 ( .A(start_reg[117]), .B(init), .Z(start_in[117]) );
  AND U25578 ( .A(start_reg[116]), .B(init), .Z(start_in[116]) );
  AND U25579 ( .A(start_reg[115]), .B(init), .Z(start_in[115]) );
  AND U25580 ( .A(start_reg[114]), .B(init), .Z(start_in[114]) );
  AND U25581 ( .A(start_reg[113]), .B(init), .Z(start_in[113]) );
  AND U25582 ( .A(start_reg[112]), .B(init), .Z(start_in[112]) );
  AND U25583 ( .A(start_reg[111]), .B(init), .Z(start_in[111]) );
  AND U25584 ( .A(start_reg[110]), .B(init), .Z(start_in[110]) );
  AND U25585 ( .A(start_reg[10]), .B(init), .Z(start_in[10]) );
  AND U25586 ( .A(start_reg[109]), .B(init), .Z(start_in[109]) );
  AND U25587 ( .A(start_reg[108]), .B(init), .Z(start_in[108]) );
  AND U25588 ( .A(start_reg[107]), .B(init), .Z(start_in[107]) );
  AND U25589 ( .A(start_reg[106]), .B(init), .Z(start_in[106]) );
  AND U25590 ( .A(start_reg[105]), .B(init), .Z(start_in[105]) );
  AND U25591 ( .A(start_reg[104]), .B(init), .Z(start_in[104]) );
  AND U25592 ( .A(start_reg[103]), .B(init), .Z(start_in[103]) );
  AND U25593 ( .A(start_reg[102]), .B(init), .Z(start_in[102]) );
  AND U25594 ( .A(start_reg[1022]), .B(init), .Z(start_in[1022]) );
  AND U25595 ( .A(start_reg[1021]), .B(init), .Z(start_in[1021]) );
  AND U25596 ( .A(start_reg[1020]), .B(init), .Z(start_in[1020]) );
  AND U25597 ( .A(start_reg[101]), .B(init), .Z(start_in[101]) );
  AND U25598 ( .A(start_reg[1019]), .B(init), .Z(start_in[1019]) );
  AND U25599 ( .A(start_reg[1018]), .B(init), .Z(start_in[1018]) );
  AND U25600 ( .A(start_reg[1017]), .B(init), .Z(start_in[1017]) );
  AND U25601 ( .A(start_reg[1016]), .B(init), .Z(start_in[1016]) );
  AND U25602 ( .A(start_reg[1015]), .B(init), .Z(start_in[1015]) );
  AND U25603 ( .A(start_reg[1014]), .B(init), .Z(start_in[1014]) );
  AND U25604 ( .A(start_reg[1013]), .B(init), .Z(start_in[1013]) );
  AND U25605 ( .A(start_reg[1012]), .B(init), .Z(start_in[1012]) );
  AND U25606 ( .A(start_reg[1011]), .B(init), .Z(start_in[1011]) );
  AND U25607 ( .A(start_reg[1010]), .B(init), .Z(start_in[1010]) );
  AND U25608 ( .A(start_reg[100]), .B(init), .Z(start_in[100]) );
  AND U25609 ( .A(start_reg[1009]), .B(init), .Z(start_in[1009]) );
  AND U25610 ( .A(start_reg[1008]), .B(init), .Z(start_in[1008]) );
  AND U25611 ( .A(start_reg[1007]), .B(init), .Z(start_in[1007]) );
  AND U25612 ( .A(start_reg[1006]), .B(init), .Z(start_in[1006]) );
  AND U25613 ( .A(start_reg[1005]), .B(init), .Z(start_in[1005]) );
  AND U25614 ( .A(start_reg[1004]), .B(init), .Z(start_in[1004]) );
  AND U25615 ( .A(start_reg[1003]), .B(init), .Z(start_in[1003]) );
  AND U25616 ( .A(start_reg[1002]), .B(init), .Z(start_in[1002]) );
  AND U25617 ( .A(start_reg[1001]), .B(init), .Z(start_in[1001]) );
  AND U25618 ( .A(start_reg[1000]), .B(init), .Z(start_in[1000]) );
  NANDN U25619 ( .A(start_reg[0]), .B(init), .Z(start_in[0]) );
  NAND U25620 ( .A(n19477), .B(n19478), .Z(n15378) );
  NAND U25621 ( .A(n15382), .B(start_reg[1023]), .Z(n19478) );
  IV U25622 ( .A(n15381), .Z(n15382) );
  NANDN U25623 ( .A(start_in[1023]), .B(mul_pow), .Z(n19477) );
  NAND U25624 ( .A(n19479), .B(n19480), .Z(n15377) );
  NANDN U25625 ( .A(n19481), .B(ereg[0]), .Z(n19480) );
  NANDN U25626 ( .A(init), .B(e[0]), .Z(n19479) );
  NAND U25627 ( .A(n19482), .B(n19483), .Z(n15376) );
  NANDN U25628 ( .A(init), .B(e[1]), .Z(n19483) );
  AND U25629 ( .A(n19484), .B(n19485), .Z(n19482) );
  NAND U25630 ( .A(n19486), .B(ereg[0]), .Z(n19485) );
  NANDN U25631 ( .A(n19481), .B(ereg[1]), .Z(n19484) );
  NAND U25632 ( .A(n19487), .B(n19488), .Z(n15375) );
  NANDN U25633 ( .A(init), .B(e[2]), .Z(n19488) );
  AND U25634 ( .A(n19489), .B(n19490), .Z(n19487) );
  NAND U25635 ( .A(ereg[1]), .B(n19486), .Z(n19490) );
  NANDN U25636 ( .A(n19481), .B(ereg[2]), .Z(n19489) );
  NAND U25637 ( .A(n19491), .B(n19492), .Z(n15374) );
  NANDN U25638 ( .A(init), .B(e[3]), .Z(n19492) );
  AND U25639 ( .A(n19493), .B(n19494), .Z(n19491) );
  NAND U25640 ( .A(ereg[2]), .B(n19486), .Z(n19494) );
  NANDN U25641 ( .A(n19481), .B(ereg[3]), .Z(n19493) );
  NAND U25642 ( .A(n19495), .B(n19496), .Z(n15373) );
  NANDN U25643 ( .A(init), .B(e[4]), .Z(n19496) );
  AND U25644 ( .A(n19497), .B(n19498), .Z(n19495) );
  NAND U25645 ( .A(ereg[3]), .B(n19486), .Z(n19498) );
  NANDN U25646 ( .A(n19481), .B(ereg[4]), .Z(n19497) );
  NAND U25647 ( .A(n19499), .B(n19500), .Z(n15372) );
  NANDN U25648 ( .A(init), .B(e[5]), .Z(n19500) );
  AND U25649 ( .A(n19501), .B(n19502), .Z(n19499) );
  NAND U25650 ( .A(ereg[4]), .B(n19486), .Z(n19502) );
  NANDN U25651 ( .A(n19481), .B(ereg[5]), .Z(n19501) );
  NAND U25652 ( .A(n19503), .B(n19504), .Z(n15371) );
  NANDN U25653 ( .A(init), .B(e[6]), .Z(n19504) );
  AND U25654 ( .A(n19505), .B(n19506), .Z(n19503) );
  NAND U25655 ( .A(ereg[5]), .B(n19486), .Z(n19506) );
  NANDN U25656 ( .A(n19481), .B(ereg[6]), .Z(n19505) );
  NAND U25657 ( .A(n19507), .B(n19508), .Z(n15370) );
  NANDN U25658 ( .A(init), .B(e[7]), .Z(n19508) );
  AND U25659 ( .A(n19509), .B(n19510), .Z(n19507) );
  NAND U25660 ( .A(ereg[6]), .B(n19486), .Z(n19510) );
  NANDN U25661 ( .A(n19481), .B(ereg[7]), .Z(n19509) );
  NAND U25662 ( .A(n19511), .B(n19512), .Z(n15369) );
  NANDN U25663 ( .A(init), .B(e[8]), .Z(n19512) );
  AND U25664 ( .A(n19513), .B(n19514), .Z(n19511) );
  NAND U25665 ( .A(ereg[7]), .B(n19486), .Z(n19514) );
  NANDN U25666 ( .A(n19481), .B(ereg[8]), .Z(n19513) );
  NAND U25667 ( .A(n19515), .B(n19516), .Z(n15368) );
  NANDN U25668 ( .A(init), .B(e[9]), .Z(n19516) );
  AND U25669 ( .A(n19517), .B(n19518), .Z(n19515) );
  NAND U25670 ( .A(ereg[8]), .B(n19486), .Z(n19518) );
  NANDN U25671 ( .A(n19481), .B(ereg[9]), .Z(n19517) );
  NAND U25672 ( .A(n19519), .B(n19520), .Z(n15367) );
  NANDN U25673 ( .A(init), .B(e[10]), .Z(n19520) );
  AND U25674 ( .A(n19521), .B(n19522), .Z(n19519) );
  NAND U25675 ( .A(ereg[9]), .B(n19486), .Z(n19522) );
  NANDN U25676 ( .A(n19481), .B(ereg[10]), .Z(n19521) );
  NAND U25677 ( .A(n19523), .B(n19524), .Z(n15366) );
  NANDN U25678 ( .A(init), .B(e[11]), .Z(n19524) );
  AND U25679 ( .A(n19525), .B(n19526), .Z(n19523) );
  NAND U25680 ( .A(ereg[10]), .B(n19486), .Z(n19526) );
  NANDN U25681 ( .A(n19481), .B(ereg[11]), .Z(n19525) );
  NAND U25682 ( .A(n19527), .B(n19528), .Z(n15365) );
  NANDN U25683 ( .A(init), .B(e[12]), .Z(n19528) );
  AND U25684 ( .A(n19529), .B(n19530), .Z(n19527) );
  NAND U25685 ( .A(ereg[11]), .B(n19486), .Z(n19530) );
  NANDN U25686 ( .A(n19481), .B(ereg[12]), .Z(n19529) );
  NAND U25687 ( .A(n19531), .B(n19532), .Z(n15364) );
  NANDN U25688 ( .A(init), .B(e[13]), .Z(n19532) );
  AND U25689 ( .A(n19533), .B(n19534), .Z(n19531) );
  NAND U25690 ( .A(ereg[12]), .B(n19486), .Z(n19534) );
  NANDN U25691 ( .A(n19481), .B(ereg[13]), .Z(n19533) );
  NAND U25692 ( .A(n19535), .B(n19536), .Z(n15363) );
  NANDN U25693 ( .A(init), .B(e[14]), .Z(n19536) );
  AND U25694 ( .A(n19537), .B(n19538), .Z(n19535) );
  NAND U25695 ( .A(ereg[13]), .B(n19486), .Z(n19538) );
  NANDN U25696 ( .A(n19481), .B(ereg[14]), .Z(n19537) );
  NAND U25697 ( .A(n19539), .B(n19540), .Z(n15362) );
  NANDN U25698 ( .A(init), .B(e[15]), .Z(n19540) );
  AND U25699 ( .A(n19541), .B(n19542), .Z(n19539) );
  NAND U25700 ( .A(ereg[14]), .B(n19486), .Z(n19542) );
  NANDN U25701 ( .A(n19481), .B(ereg[15]), .Z(n19541) );
  NAND U25702 ( .A(n19543), .B(n19544), .Z(n15361) );
  NANDN U25703 ( .A(init), .B(e[16]), .Z(n19544) );
  AND U25704 ( .A(n19545), .B(n19546), .Z(n19543) );
  NAND U25705 ( .A(ereg[15]), .B(n19486), .Z(n19546) );
  NANDN U25706 ( .A(n19481), .B(ereg[16]), .Z(n19545) );
  NAND U25707 ( .A(n19547), .B(n19548), .Z(n15360) );
  NANDN U25708 ( .A(init), .B(e[17]), .Z(n19548) );
  AND U25709 ( .A(n19549), .B(n19550), .Z(n19547) );
  NAND U25710 ( .A(ereg[16]), .B(n19486), .Z(n19550) );
  NANDN U25711 ( .A(n19481), .B(ereg[17]), .Z(n19549) );
  NAND U25712 ( .A(n19551), .B(n19552), .Z(n15359) );
  NANDN U25713 ( .A(init), .B(e[18]), .Z(n19552) );
  AND U25714 ( .A(n19553), .B(n19554), .Z(n19551) );
  NAND U25715 ( .A(ereg[17]), .B(n19486), .Z(n19554) );
  NANDN U25716 ( .A(n19481), .B(ereg[18]), .Z(n19553) );
  NAND U25717 ( .A(n19555), .B(n19556), .Z(n15358) );
  NANDN U25718 ( .A(init), .B(e[19]), .Z(n19556) );
  AND U25719 ( .A(n19557), .B(n19558), .Z(n19555) );
  NAND U25720 ( .A(ereg[18]), .B(n19486), .Z(n19558) );
  NANDN U25721 ( .A(n19481), .B(ereg[19]), .Z(n19557) );
  NAND U25722 ( .A(n19559), .B(n19560), .Z(n15357) );
  NANDN U25723 ( .A(init), .B(e[20]), .Z(n19560) );
  AND U25724 ( .A(n19561), .B(n19562), .Z(n19559) );
  NAND U25725 ( .A(ereg[19]), .B(n19486), .Z(n19562) );
  NANDN U25726 ( .A(n19481), .B(ereg[20]), .Z(n19561) );
  NAND U25727 ( .A(n19563), .B(n19564), .Z(n15356) );
  NANDN U25728 ( .A(init), .B(e[21]), .Z(n19564) );
  AND U25729 ( .A(n19565), .B(n19566), .Z(n19563) );
  NAND U25730 ( .A(ereg[20]), .B(n19486), .Z(n19566) );
  NANDN U25731 ( .A(n19481), .B(ereg[21]), .Z(n19565) );
  NAND U25732 ( .A(n19567), .B(n19568), .Z(n15355) );
  NANDN U25733 ( .A(init), .B(e[22]), .Z(n19568) );
  AND U25734 ( .A(n19569), .B(n19570), .Z(n19567) );
  NAND U25735 ( .A(ereg[21]), .B(n19486), .Z(n19570) );
  NANDN U25736 ( .A(n19481), .B(ereg[22]), .Z(n19569) );
  NAND U25737 ( .A(n19571), .B(n19572), .Z(n15354) );
  NANDN U25738 ( .A(init), .B(e[23]), .Z(n19572) );
  AND U25739 ( .A(n19573), .B(n19574), .Z(n19571) );
  NAND U25740 ( .A(ereg[22]), .B(n19486), .Z(n19574) );
  NANDN U25741 ( .A(n19481), .B(ereg[23]), .Z(n19573) );
  NAND U25742 ( .A(n19575), .B(n19576), .Z(n15353) );
  NANDN U25743 ( .A(init), .B(e[24]), .Z(n19576) );
  AND U25744 ( .A(n19577), .B(n19578), .Z(n19575) );
  NAND U25745 ( .A(ereg[23]), .B(n19486), .Z(n19578) );
  NANDN U25746 ( .A(n19481), .B(ereg[24]), .Z(n19577) );
  NAND U25747 ( .A(n19579), .B(n19580), .Z(n15352) );
  NANDN U25748 ( .A(init), .B(e[25]), .Z(n19580) );
  AND U25749 ( .A(n19581), .B(n19582), .Z(n19579) );
  NAND U25750 ( .A(ereg[24]), .B(n19486), .Z(n19582) );
  NANDN U25751 ( .A(n19481), .B(ereg[25]), .Z(n19581) );
  NAND U25752 ( .A(n19583), .B(n19584), .Z(n15351) );
  NANDN U25753 ( .A(init), .B(e[26]), .Z(n19584) );
  AND U25754 ( .A(n19585), .B(n19586), .Z(n19583) );
  NAND U25755 ( .A(ereg[25]), .B(n19486), .Z(n19586) );
  NANDN U25756 ( .A(n19481), .B(ereg[26]), .Z(n19585) );
  NAND U25757 ( .A(n19587), .B(n19588), .Z(n15350) );
  NANDN U25758 ( .A(init), .B(e[27]), .Z(n19588) );
  AND U25759 ( .A(n19589), .B(n19590), .Z(n19587) );
  NAND U25760 ( .A(ereg[26]), .B(n19486), .Z(n19590) );
  NANDN U25761 ( .A(n19481), .B(ereg[27]), .Z(n19589) );
  NAND U25762 ( .A(n19591), .B(n19592), .Z(n15349) );
  NANDN U25763 ( .A(init), .B(e[28]), .Z(n19592) );
  AND U25764 ( .A(n19593), .B(n19594), .Z(n19591) );
  NAND U25765 ( .A(ereg[27]), .B(n19486), .Z(n19594) );
  NANDN U25766 ( .A(n19481), .B(ereg[28]), .Z(n19593) );
  NAND U25767 ( .A(n19595), .B(n19596), .Z(n15348) );
  NANDN U25768 ( .A(init), .B(e[29]), .Z(n19596) );
  AND U25769 ( .A(n19597), .B(n19598), .Z(n19595) );
  NAND U25770 ( .A(ereg[28]), .B(n19486), .Z(n19598) );
  NANDN U25771 ( .A(n19481), .B(ereg[29]), .Z(n19597) );
  NAND U25772 ( .A(n19599), .B(n19600), .Z(n15347) );
  NANDN U25773 ( .A(init), .B(e[30]), .Z(n19600) );
  AND U25774 ( .A(n19601), .B(n19602), .Z(n19599) );
  NAND U25775 ( .A(ereg[29]), .B(n19486), .Z(n19602) );
  NANDN U25776 ( .A(n19481), .B(ereg[30]), .Z(n19601) );
  NAND U25777 ( .A(n19603), .B(n19604), .Z(n15346) );
  NANDN U25778 ( .A(init), .B(e[31]), .Z(n19604) );
  AND U25779 ( .A(n19605), .B(n19606), .Z(n19603) );
  NAND U25780 ( .A(ereg[30]), .B(n19486), .Z(n19606) );
  NANDN U25781 ( .A(n19481), .B(ereg[31]), .Z(n19605) );
  NAND U25782 ( .A(n19607), .B(n19608), .Z(n15345) );
  NANDN U25783 ( .A(init), .B(e[32]), .Z(n19608) );
  AND U25784 ( .A(n19609), .B(n19610), .Z(n19607) );
  NAND U25785 ( .A(ereg[31]), .B(n19486), .Z(n19610) );
  NANDN U25786 ( .A(n19481), .B(ereg[32]), .Z(n19609) );
  NAND U25787 ( .A(n19611), .B(n19612), .Z(n15344) );
  NANDN U25788 ( .A(init), .B(e[33]), .Z(n19612) );
  AND U25789 ( .A(n19613), .B(n19614), .Z(n19611) );
  NAND U25790 ( .A(ereg[32]), .B(n19486), .Z(n19614) );
  NANDN U25791 ( .A(n19481), .B(ereg[33]), .Z(n19613) );
  NAND U25792 ( .A(n19615), .B(n19616), .Z(n15343) );
  NANDN U25793 ( .A(init), .B(e[34]), .Z(n19616) );
  AND U25794 ( .A(n19617), .B(n19618), .Z(n19615) );
  NAND U25795 ( .A(ereg[33]), .B(n19486), .Z(n19618) );
  NANDN U25796 ( .A(n19481), .B(ereg[34]), .Z(n19617) );
  NAND U25797 ( .A(n19619), .B(n19620), .Z(n15342) );
  NANDN U25798 ( .A(init), .B(e[35]), .Z(n19620) );
  AND U25799 ( .A(n19621), .B(n19622), .Z(n19619) );
  NAND U25800 ( .A(ereg[34]), .B(n19486), .Z(n19622) );
  NANDN U25801 ( .A(n19481), .B(ereg[35]), .Z(n19621) );
  NAND U25802 ( .A(n19623), .B(n19624), .Z(n15341) );
  NANDN U25803 ( .A(init), .B(e[36]), .Z(n19624) );
  AND U25804 ( .A(n19625), .B(n19626), .Z(n19623) );
  NAND U25805 ( .A(ereg[35]), .B(n19486), .Z(n19626) );
  NANDN U25806 ( .A(n19481), .B(ereg[36]), .Z(n19625) );
  NAND U25807 ( .A(n19627), .B(n19628), .Z(n15340) );
  NANDN U25808 ( .A(init), .B(e[37]), .Z(n19628) );
  AND U25809 ( .A(n19629), .B(n19630), .Z(n19627) );
  NAND U25810 ( .A(ereg[36]), .B(n19486), .Z(n19630) );
  NANDN U25811 ( .A(n19481), .B(ereg[37]), .Z(n19629) );
  NAND U25812 ( .A(n19631), .B(n19632), .Z(n15339) );
  NANDN U25813 ( .A(init), .B(e[38]), .Z(n19632) );
  AND U25814 ( .A(n19633), .B(n19634), .Z(n19631) );
  NAND U25815 ( .A(ereg[37]), .B(n19486), .Z(n19634) );
  NANDN U25816 ( .A(n19481), .B(ereg[38]), .Z(n19633) );
  NAND U25817 ( .A(n19635), .B(n19636), .Z(n15338) );
  NANDN U25818 ( .A(init), .B(e[39]), .Z(n19636) );
  AND U25819 ( .A(n19637), .B(n19638), .Z(n19635) );
  NAND U25820 ( .A(ereg[38]), .B(n19486), .Z(n19638) );
  NANDN U25821 ( .A(n19481), .B(ereg[39]), .Z(n19637) );
  NAND U25822 ( .A(n19639), .B(n19640), .Z(n15337) );
  NANDN U25823 ( .A(init), .B(e[40]), .Z(n19640) );
  AND U25824 ( .A(n19641), .B(n19642), .Z(n19639) );
  NAND U25825 ( .A(ereg[39]), .B(n19486), .Z(n19642) );
  NANDN U25826 ( .A(n19481), .B(ereg[40]), .Z(n19641) );
  NAND U25827 ( .A(n19643), .B(n19644), .Z(n15336) );
  NANDN U25828 ( .A(init), .B(e[41]), .Z(n19644) );
  AND U25829 ( .A(n19645), .B(n19646), .Z(n19643) );
  NAND U25830 ( .A(ereg[40]), .B(n19486), .Z(n19646) );
  NANDN U25831 ( .A(n19481), .B(ereg[41]), .Z(n19645) );
  NAND U25832 ( .A(n19647), .B(n19648), .Z(n15335) );
  NANDN U25833 ( .A(init), .B(e[42]), .Z(n19648) );
  AND U25834 ( .A(n19649), .B(n19650), .Z(n19647) );
  NAND U25835 ( .A(ereg[41]), .B(n19486), .Z(n19650) );
  NANDN U25836 ( .A(n19481), .B(ereg[42]), .Z(n19649) );
  NAND U25837 ( .A(n19651), .B(n19652), .Z(n15334) );
  NANDN U25838 ( .A(init), .B(e[43]), .Z(n19652) );
  AND U25839 ( .A(n19653), .B(n19654), .Z(n19651) );
  NAND U25840 ( .A(ereg[42]), .B(n19486), .Z(n19654) );
  NANDN U25841 ( .A(n19481), .B(ereg[43]), .Z(n19653) );
  NAND U25842 ( .A(n19655), .B(n19656), .Z(n15333) );
  NANDN U25843 ( .A(init), .B(e[44]), .Z(n19656) );
  AND U25844 ( .A(n19657), .B(n19658), .Z(n19655) );
  NAND U25845 ( .A(ereg[43]), .B(n19486), .Z(n19658) );
  NANDN U25846 ( .A(n19481), .B(ereg[44]), .Z(n19657) );
  NAND U25847 ( .A(n19659), .B(n19660), .Z(n15332) );
  NANDN U25848 ( .A(init), .B(e[45]), .Z(n19660) );
  AND U25849 ( .A(n19661), .B(n19662), .Z(n19659) );
  NAND U25850 ( .A(ereg[44]), .B(n19486), .Z(n19662) );
  NANDN U25851 ( .A(n19481), .B(ereg[45]), .Z(n19661) );
  NAND U25852 ( .A(n19663), .B(n19664), .Z(n15331) );
  NANDN U25853 ( .A(init), .B(e[46]), .Z(n19664) );
  AND U25854 ( .A(n19665), .B(n19666), .Z(n19663) );
  NAND U25855 ( .A(ereg[45]), .B(n19486), .Z(n19666) );
  NANDN U25856 ( .A(n19481), .B(ereg[46]), .Z(n19665) );
  NAND U25857 ( .A(n19667), .B(n19668), .Z(n15330) );
  NANDN U25858 ( .A(init), .B(e[47]), .Z(n19668) );
  AND U25859 ( .A(n19669), .B(n19670), .Z(n19667) );
  NAND U25860 ( .A(ereg[46]), .B(n19486), .Z(n19670) );
  NANDN U25861 ( .A(n19481), .B(ereg[47]), .Z(n19669) );
  NAND U25862 ( .A(n19671), .B(n19672), .Z(n15329) );
  NANDN U25863 ( .A(init), .B(e[48]), .Z(n19672) );
  AND U25864 ( .A(n19673), .B(n19674), .Z(n19671) );
  NAND U25865 ( .A(ereg[47]), .B(n19486), .Z(n19674) );
  NANDN U25866 ( .A(n19481), .B(ereg[48]), .Z(n19673) );
  NAND U25867 ( .A(n19675), .B(n19676), .Z(n15328) );
  NANDN U25868 ( .A(init), .B(e[49]), .Z(n19676) );
  AND U25869 ( .A(n19677), .B(n19678), .Z(n19675) );
  NAND U25870 ( .A(ereg[48]), .B(n19486), .Z(n19678) );
  NANDN U25871 ( .A(n19481), .B(ereg[49]), .Z(n19677) );
  NAND U25872 ( .A(n19679), .B(n19680), .Z(n15327) );
  NANDN U25873 ( .A(init), .B(e[50]), .Z(n19680) );
  AND U25874 ( .A(n19681), .B(n19682), .Z(n19679) );
  NAND U25875 ( .A(ereg[49]), .B(n19486), .Z(n19682) );
  NANDN U25876 ( .A(n19481), .B(ereg[50]), .Z(n19681) );
  NAND U25877 ( .A(n19683), .B(n19684), .Z(n15326) );
  NANDN U25878 ( .A(init), .B(e[51]), .Z(n19684) );
  AND U25879 ( .A(n19685), .B(n19686), .Z(n19683) );
  NAND U25880 ( .A(ereg[50]), .B(n19486), .Z(n19686) );
  NANDN U25881 ( .A(n19481), .B(ereg[51]), .Z(n19685) );
  NAND U25882 ( .A(n19687), .B(n19688), .Z(n15325) );
  NANDN U25883 ( .A(init), .B(e[52]), .Z(n19688) );
  AND U25884 ( .A(n19689), .B(n19690), .Z(n19687) );
  NAND U25885 ( .A(ereg[51]), .B(n19486), .Z(n19690) );
  NANDN U25886 ( .A(n19481), .B(ereg[52]), .Z(n19689) );
  NAND U25887 ( .A(n19691), .B(n19692), .Z(n15324) );
  NANDN U25888 ( .A(init), .B(e[53]), .Z(n19692) );
  AND U25889 ( .A(n19693), .B(n19694), .Z(n19691) );
  NAND U25890 ( .A(ereg[52]), .B(n19486), .Z(n19694) );
  NANDN U25891 ( .A(n19481), .B(ereg[53]), .Z(n19693) );
  NAND U25892 ( .A(n19695), .B(n19696), .Z(n15323) );
  NANDN U25893 ( .A(init), .B(e[54]), .Z(n19696) );
  AND U25894 ( .A(n19697), .B(n19698), .Z(n19695) );
  NAND U25895 ( .A(ereg[53]), .B(n19486), .Z(n19698) );
  NANDN U25896 ( .A(n19481), .B(ereg[54]), .Z(n19697) );
  NAND U25897 ( .A(n19699), .B(n19700), .Z(n15322) );
  NANDN U25898 ( .A(init), .B(e[55]), .Z(n19700) );
  AND U25899 ( .A(n19701), .B(n19702), .Z(n19699) );
  NAND U25900 ( .A(ereg[54]), .B(n19486), .Z(n19702) );
  NANDN U25901 ( .A(n19481), .B(ereg[55]), .Z(n19701) );
  NAND U25902 ( .A(n19703), .B(n19704), .Z(n15321) );
  NANDN U25903 ( .A(init), .B(e[56]), .Z(n19704) );
  AND U25904 ( .A(n19705), .B(n19706), .Z(n19703) );
  NAND U25905 ( .A(ereg[55]), .B(n19486), .Z(n19706) );
  NANDN U25906 ( .A(n19481), .B(ereg[56]), .Z(n19705) );
  NAND U25907 ( .A(n19707), .B(n19708), .Z(n15320) );
  NANDN U25908 ( .A(init), .B(e[57]), .Z(n19708) );
  AND U25909 ( .A(n19709), .B(n19710), .Z(n19707) );
  NAND U25910 ( .A(ereg[56]), .B(n19486), .Z(n19710) );
  NANDN U25911 ( .A(n19481), .B(ereg[57]), .Z(n19709) );
  NAND U25912 ( .A(n19711), .B(n19712), .Z(n15319) );
  NANDN U25913 ( .A(init), .B(e[58]), .Z(n19712) );
  AND U25914 ( .A(n19713), .B(n19714), .Z(n19711) );
  NAND U25915 ( .A(ereg[57]), .B(n19486), .Z(n19714) );
  NANDN U25916 ( .A(n19481), .B(ereg[58]), .Z(n19713) );
  NAND U25917 ( .A(n19715), .B(n19716), .Z(n15318) );
  NANDN U25918 ( .A(init), .B(e[59]), .Z(n19716) );
  AND U25919 ( .A(n19717), .B(n19718), .Z(n19715) );
  NAND U25920 ( .A(ereg[58]), .B(n19486), .Z(n19718) );
  NANDN U25921 ( .A(n19481), .B(ereg[59]), .Z(n19717) );
  NAND U25922 ( .A(n19719), .B(n19720), .Z(n15317) );
  NANDN U25923 ( .A(init), .B(e[60]), .Z(n19720) );
  AND U25924 ( .A(n19721), .B(n19722), .Z(n19719) );
  NAND U25925 ( .A(ereg[59]), .B(n19486), .Z(n19722) );
  NANDN U25926 ( .A(n19481), .B(ereg[60]), .Z(n19721) );
  NAND U25927 ( .A(n19723), .B(n19724), .Z(n15316) );
  NANDN U25928 ( .A(init), .B(e[61]), .Z(n19724) );
  AND U25929 ( .A(n19725), .B(n19726), .Z(n19723) );
  NAND U25930 ( .A(ereg[60]), .B(n19486), .Z(n19726) );
  NANDN U25931 ( .A(n19481), .B(ereg[61]), .Z(n19725) );
  NAND U25932 ( .A(n19727), .B(n19728), .Z(n15315) );
  NANDN U25933 ( .A(init), .B(e[62]), .Z(n19728) );
  AND U25934 ( .A(n19729), .B(n19730), .Z(n19727) );
  NAND U25935 ( .A(ereg[61]), .B(n19486), .Z(n19730) );
  NANDN U25936 ( .A(n19481), .B(ereg[62]), .Z(n19729) );
  NAND U25937 ( .A(n19731), .B(n19732), .Z(n15314) );
  NANDN U25938 ( .A(init), .B(e[63]), .Z(n19732) );
  AND U25939 ( .A(n19733), .B(n19734), .Z(n19731) );
  NAND U25940 ( .A(ereg[62]), .B(n19486), .Z(n19734) );
  NANDN U25941 ( .A(n19481), .B(ereg[63]), .Z(n19733) );
  NAND U25942 ( .A(n19735), .B(n19736), .Z(n15313) );
  NANDN U25943 ( .A(init), .B(e[64]), .Z(n19736) );
  AND U25944 ( .A(n19737), .B(n19738), .Z(n19735) );
  NAND U25945 ( .A(ereg[63]), .B(n19486), .Z(n19738) );
  NANDN U25946 ( .A(n19481), .B(ereg[64]), .Z(n19737) );
  NAND U25947 ( .A(n19739), .B(n19740), .Z(n15312) );
  NANDN U25948 ( .A(init), .B(e[65]), .Z(n19740) );
  AND U25949 ( .A(n19741), .B(n19742), .Z(n19739) );
  NAND U25950 ( .A(ereg[64]), .B(n19486), .Z(n19742) );
  NANDN U25951 ( .A(n19481), .B(ereg[65]), .Z(n19741) );
  NAND U25952 ( .A(n19743), .B(n19744), .Z(n15311) );
  NANDN U25953 ( .A(init), .B(e[66]), .Z(n19744) );
  AND U25954 ( .A(n19745), .B(n19746), .Z(n19743) );
  NAND U25955 ( .A(ereg[65]), .B(n19486), .Z(n19746) );
  NANDN U25956 ( .A(n19481), .B(ereg[66]), .Z(n19745) );
  NAND U25957 ( .A(n19747), .B(n19748), .Z(n15310) );
  NANDN U25958 ( .A(init), .B(e[67]), .Z(n19748) );
  AND U25959 ( .A(n19749), .B(n19750), .Z(n19747) );
  NAND U25960 ( .A(ereg[66]), .B(n19486), .Z(n19750) );
  NANDN U25961 ( .A(n19481), .B(ereg[67]), .Z(n19749) );
  NAND U25962 ( .A(n19751), .B(n19752), .Z(n15309) );
  NANDN U25963 ( .A(init), .B(e[68]), .Z(n19752) );
  AND U25964 ( .A(n19753), .B(n19754), .Z(n19751) );
  NAND U25965 ( .A(ereg[67]), .B(n19486), .Z(n19754) );
  NANDN U25966 ( .A(n19481), .B(ereg[68]), .Z(n19753) );
  NAND U25967 ( .A(n19755), .B(n19756), .Z(n15308) );
  NANDN U25968 ( .A(init), .B(e[69]), .Z(n19756) );
  AND U25969 ( .A(n19757), .B(n19758), .Z(n19755) );
  NAND U25970 ( .A(ereg[68]), .B(n19486), .Z(n19758) );
  NANDN U25971 ( .A(n19481), .B(ereg[69]), .Z(n19757) );
  NAND U25972 ( .A(n19759), .B(n19760), .Z(n15307) );
  NANDN U25973 ( .A(init), .B(e[70]), .Z(n19760) );
  AND U25974 ( .A(n19761), .B(n19762), .Z(n19759) );
  NAND U25975 ( .A(ereg[69]), .B(n19486), .Z(n19762) );
  NANDN U25976 ( .A(n19481), .B(ereg[70]), .Z(n19761) );
  NAND U25977 ( .A(n19763), .B(n19764), .Z(n15306) );
  NANDN U25978 ( .A(init), .B(e[71]), .Z(n19764) );
  AND U25979 ( .A(n19765), .B(n19766), .Z(n19763) );
  NAND U25980 ( .A(ereg[70]), .B(n19486), .Z(n19766) );
  NANDN U25981 ( .A(n19481), .B(ereg[71]), .Z(n19765) );
  NAND U25982 ( .A(n19767), .B(n19768), .Z(n15305) );
  NANDN U25983 ( .A(init), .B(e[72]), .Z(n19768) );
  AND U25984 ( .A(n19769), .B(n19770), .Z(n19767) );
  NAND U25985 ( .A(ereg[71]), .B(n19486), .Z(n19770) );
  NANDN U25986 ( .A(n19481), .B(ereg[72]), .Z(n19769) );
  NAND U25987 ( .A(n19771), .B(n19772), .Z(n15304) );
  NANDN U25988 ( .A(init), .B(e[73]), .Z(n19772) );
  AND U25989 ( .A(n19773), .B(n19774), .Z(n19771) );
  NAND U25990 ( .A(ereg[72]), .B(n19486), .Z(n19774) );
  NANDN U25991 ( .A(n19481), .B(ereg[73]), .Z(n19773) );
  NAND U25992 ( .A(n19775), .B(n19776), .Z(n15303) );
  NANDN U25993 ( .A(init), .B(e[74]), .Z(n19776) );
  AND U25994 ( .A(n19777), .B(n19778), .Z(n19775) );
  NAND U25995 ( .A(ereg[73]), .B(n19486), .Z(n19778) );
  NANDN U25996 ( .A(n19481), .B(ereg[74]), .Z(n19777) );
  NAND U25997 ( .A(n19779), .B(n19780), .Z(n15302) );
  NANDN U25998 ( .A(init), .B(e[75]), .Z(n19780) );
  AND U25999 ( .A(n19781), .B(n19782), .Z(n19779) );
  NAND U26000 ( .A(ereg[74]), .B(n19486), .Z(n19782) );
  NANDN U26001 ( .A(n19481), .B(ereg[75]), .Z(n19781) );
  NAND U26002 ( .A(n19783), .B(n19784), .Z(n15301) );
  NANDN U26003 ( .A(init), .B(e[76]), .Z(n19784) );
  AND U26004 ( .A(n19785), .B(n19786), .Z(n19783) );
  NAND U26005 ( .A(ereg[75]), .B(n19486), .Z(n19786) );
  NANDN U26006 ( .A(n19481), .B(ereg[76]), .Z(n19785) );
  NAND U26007 ( .A(n19787), .B(n19788), .Z(n15300) );
  NANDN U26008 ( .A(init), .B(e[77]), .Z(n19788) );
  AND U26009 ( .A(n19789), .B(n19790), .Z(n19787) );
  NAND U26010 ( .A(ereg[76]), .B(n19486), .Z(n19790) );
  NANDN U26011 ( .A(n19481), .B(ereg[77]), .Z(n19789) );
  NAND U26012 ( .A(n19791), .B(n19792), .Z(n15299) );
  NANDN U26013 ( .A(init), .B(e[78]), .Z(n19792) );
  AND U26014 ( .A(n19793), .B(n19794), .Z(n19791) );
  NAND U26015 ( .A(ereg[77]), .B(n19486), .Z(n19794) );
  NANDN U26016 ( .A(n19481), .B(ereg[78]), .Z(n19793) );
  NAND U26017 ( .A(n19795), .B(n19796), .Z(n15298) );
  NANDN U26018 ( .A(init), .B(e[79]), .Z(n19796) );
  AND U26019 ( .A(n19797), .B(n19798), .Z(n19795) );
  NAND U26020 ( .A(ereg[78]), .B(n19486), .Z(n19798) );
  NANDN U26021 ( .A(n19481), .B(ereg[79]), .Z(n19797) );
  NAND U26022 ( .A(n19799), .B(n19800), .Z(n15297) );
  NANDN U26023 ( .A(init), .B(e[80]), .Z(n19800) );
  AND U26024 ( .A(n19801), .B(n19802), .Z(n19799) );
  NAND U26025 ( .A(ereg[79]), .B(n19486), .Z(n19802) );
  NANDN U26026 ( .A(n19481), .B(ereg[80]), .Z(n19801) );
  NAND U26027 ( .A(n19803), .B(n19804), .Z(n15296) );
  NANDN U26028 ( .A(init), .B(e[81]), .Z(n19804) );
  AND U26029 ( .A(n19805), .B(n19806), .Z(n19803) );
  NAND U26030 ( .A(ereg[80]), .B(n19486), .Z(n19806) );
  NANDN U26031 ( .A(n19481), .B(ereg[81]), .Z(n19805) );
  NAND U26032 ( .A(n19807), .B(n19808), .Z(n15295) );
  NANDN U26033 ( .A(init), .B(e[82]), .Z(n19808) );
  AND U26034 ( .A(n19809), .B(n19810), .Z(n19807) );
  NAND U26035 ( .A(ereg[81]), .B(n19486), .Z(n19810) );
  NANDN U26036 ( .A(n19481), .B(ereg[82]), .Z(n19809) );
  NAND U26037 ( .A(n19811), .B(n19812), .Z(n15294) );
  NANDN U26038 ( .A(init), .B(e[83]), .Z(n19812) );
  AND U26039 ( .A(n19813), .B(n19814), .Z(n19811) );
  NAND U26040 ( .A(ereg[82]), .B(n19486), .Z(n19814) );
  NANDN U26041 ( .A(n19481), .B(ereg[83]), .Z(n19813) );
  NAND U26042 ( .A(n19815), .B(n19816), .Z(n15293) );
  NANDN U26043 ( .A(init), .B(e[84]), .Z(n19816) );
  AND U26044 ( .A(n19817), .B(n19818), .Z(n19815) );
  NAND U26045 ( .A(ereg[83]), .B(n19486), .Z(n19818) );
  NANDN U26046 ( .A(n19481), .B(ereg[84]), .Z(n19817) );
  NAND U26047 ( .A(n19819), .B(n19820), .Z(n15292) );
  NANDN U26048 ( .A(init), .B(e[85]), .Z(n19820) );
  AND U26049 ( .A(n19821), .B(n19822), .Z(n19819) );
  NAND U26050 ( .A(ereg[84]), .B(n19486), .Z(n19822) );
  NANDN U26051 ( .A(n19481), .B(ereg[85]), .Z(n19821) );
  NAND U26052 ( .A(n19823), .B(n19824), .Z(n15291) );
  NANDN U26053 ( .A(init), .B(e[86]), .Z(n19824) );
  AND U26054 ( .A(n19825), .B(n19826), .Z(n19823) );
  NAND U26055 ( .A(ereg[85]), .B(n19486), .Z(n19826) );
  NANDN U26056 ( .A(n19481), .B(ereg[86]), .Z(n19825) );
  NAND U26057 ( .A(n19827), .B(n19828), .Z(n15290) );
  NANDN U26058 ( .A(init), .B(e[87]), .Z(n19828) );
  AND U26059 ( .A(n19829), .B(n19830), .Z(n19827) );
  NAND U26060 ( .A(ereg[86]), .B(n19486), .Z(n19830) );
  NANDN U26061 ( .A(n19481), .B(ereg[87]), .Z(n19829) );
  NAND U26062 ( .A(n19831), .B(n19832), .Z(n15289) );
  NANDN U26063 ( .A(init), .B(e[88]), .Z(n19832) );
  AND U26064 ( .A(n19833), .B(n19834), .Z(n19831) );
  NAND U26065 ( .A(ereg[87]), .B(n19486), .Z(n19834) );
  NANDN U26066 ( .A(n19481), .B(ereg[88]), .Z(n19833) );
  NAND U26067 ( .A(n19835), .B(n19836), .Z(n15288) );
  NANDN U26068 ( .A(init), .B(e[89]), .Z(n19836) );
  AND U26069 ( .A(n19837), .B(n19838), .Z(n19835) );
  NAND U26070 ( .A(ereg[88]), .B(n19486), .Z(n19838) );
  NANDN U26071 ( .A(n19481), .B(ereg[89]), .Z(n19837) );
  NAND U26072 ( .A(n19839), .B(n19840), .Z(n15287) );
  NANDN U26073 ( .A(init), .B(e[90]), .Z(n19840) );
  AND U26074 ( .A(n19841), .B(n19842), .Z(n19839) );
  NAND U26075 ( .A(ereg[89]), .B(n19486), .Z(n19842) );
  NANDN U26076 ( .A(n19481), .B(ereg[90]), .Z(n19841) );
  NAND U26077 ( .A(n19843), .B(n19844), .Z(n15286) );
  NANDN U26078 ( .A(init), .B(e[91]), .Z(n19844) );
  AND U26079 ( .A(n19845), .B(n19846), .Z(n19843) );
  NAND U26080 ( .A(ereg[90]), .B(n19486), .Z(n19846) );
  NANDN U26081 ( .A(n19481), .B(ereg[91]), .Z(n19845) );
  NAND U26082 ( .A(n19847), .B(n19848), .Z(n15285) );
  NANDN U26083 ( .A(init), .B(e[92]), .Z(n19848) );
  AND U26084 ( .A(n19849), .B(n19850), .Z(n19847) );
  NAND U26085 ( .A(ereg[91]), .B(n19486), .Z(n19850) );
  NANDN U26086 ( .A(n19481), .B(ereg[92]), .Z(n19849) );
  NAND U26087 ( .A(n19851), .B(n19852), .Z(n15284) );
  NANDN U26088 ( .A(init), .B(e[93]), .Z(n19852) );
  AND U26089 ( .A(n19853), .B(n19854), .Z(n19851) );
  NAND U26090 ( .A(ereg[92]), .B(n19486), .Z(n19854) );
  NANDN U26091 ( .A(n19481), .B(ereg[93]), .Z(n19853) );
  NAND U26092 ( .A(n19855), .B(n19856), .Z(n15283) );
  NANDN U26093 ( .A(init), .B(e[94]), .Z(n19856) );
  AND U26094 ( .A(n19857), .B(n19858), .Z(n19855) );
  NAND U26095 ( .A(ereg[93]), .B(n19486), .Z(n19858) );
  NANDN U26096 ( .A(n19481), .B(ereg[94]), .Z(n19857) );
  NAND U26097 ( .A(n19859), .B(n19860), .Z(n15282) );
  NANDN U26098 ( .A(init), .B(e[95]), .Z(n19860) );
  AND U26099 ( .A(n19861), .B(n19862), .Z(n19859) );
  NAND U26100 ( .A(ereg[94]), .B(n19486), .Z(n19862) );
  NANDN U26101 ( .A(n19481), .B(ereg[95]), .Z(n19861) );
  NAND U26102 ( .A(n19863), .B(n19864), .Z(n15281) );
  NANDN U26103 ( .A(init), .B(e[96]), .Z(n19864) );
  AND U26104 ( .A(n19865), .B(n19866), .Z(n19863) );
  NAND U26105 ( .A(ereg[95]), .B(n19486), .Z(n19866) );
  NANDN U26106 ( .A(n19481), .B(ereg[96]), .Z(n19865) );
  NAND U26107 ( .A(n19867), .B(n19868), .Z(n15280) );
  NANDN U26108 ( .A(init), .B(e[97]), .Z(n19868) );
  AND U26109 ( .A(n19869), .B(n19870), .Z(n19867) );
  NAND U26110 ( .A(ereg[96]), .B(n19486), .Z(n19870) );
  NANDN U26111 ( .A(n19481), .B(ereg[97]), .Z(n19869) );
  NAND U26112 ( .A(n19871), .B(n19872), .Z(n15279) );
  NANDN U26113 ( .A(init), .B(e[98]), .Z(n19872) );
  AND U26114 ( .A(n19873), .B(n19874), .Z(n19871) );
  NAND U26115 ( .A(ereg[97]), .B(n19486), .Z(n19874) );
  NANDN U26116 ( .A(n19481), .B(ereg[98]), .Z(n19873) );
  NAND U26117 ( .A(n19875), .B(n19876), .Z(n15278) );
  NANDN U26118 ( .A(init), .B(e[99]), .Z(n19876) );
  AND U26119 ( .A(n19877), .B(n19878), .Z(n19875) );
  NAND U26120 ( .A(ereg[98]), .B(n19486), .Z(n19878) );
  NANDN U26121 ( .A(n19481), .B(ereg[99]), .Z(n19877) );
  NAND U26122 ( .A(n19879), .B(n19880), .Z(n15277) );
  NANDN U26123 ( .A(init), .B(e[100]), .Z(n19880) );
  AND U26124 ( .A(n19881), .B(n19882), .Z(n19879) );
  NAND U26125 ( .A(ereg[99]), .B(n19486), .Z(n19882) );
  NANDN U26126 ( .A(n19481), .B(ereg[100]), .Z(n19881) );
  NAND U26127 ( .A(n19883), .B(n19884), .Z(n15276) );
  NANDN U26128 ( .A(init), .B(e[101]), .Z(n19884) );
  AND U26129 ( .A(n19885), .B(n19886), .Z(n19883) );
  NAND U26130 ( .A(ereg[100]), .B(n19486), .Z(n19886) );
  NANDN U26131 ( .A(n19481), .B(ereg[101]), .Z(n19885) );
  NAND U26132 ( .A(n19887), .B(n19888), .Z(n15275) );
  NANDN U26133 ( .A(init), .B(e[102]), .Z(n19888) );
  AND U26134 ( .A(n19889), .B(n19890), .Z(n19887) );
  NAND U26135 ( .A(ereg[101]), .B(n19486), .Z(n19890) );
  NANDN U26136 ( .A(n19481), .B(ereg[102]), .Z(n19889) );
  NAND U26137 ( .A(n19891), .B(n19892), .Z(n15274) );
  NANDN U26138 ( .A(init), .B(e[103]), .Z(n19892) );
  AND U26139 ( .A(n19893), .B(n19894), .Z(n19891) );
  NAND U26140 ( .A(ereg[102]), .B(n19486), .Z(n19894) );
  NANDN U26141 ( .A(n19481), .B(ereg[103]), .Z(n19893) );
  NAND U26142 ( .A(n19895), .B(n19896), .Z(n15273) );
  NANDN U26143 ( .A(init), .B(e[104]), .Z(n19896) );
  AND U26144 ( .A(n19897), .B(n19898), .Z(n19895) );
  NAND U26145 ( .A(ereg[103]), .B(n19486), .Z(n19898) );
  NANDN U26146 ( .A(n19481), .B(ereg[104]), .Z(n19897) );
  NAND U26147 ( .A(n19899), .B(n19900), .Z(n15272) );
  NANDN U26148 ( .A(init), .B(e[105]), .Z(n19900) );
  AND U26149 ( .A(n19901), .B(n19902), .Z(n19899) );
  NAND U26150 ( .A(ereg[104]), .B(n19486), .Z(n19902) );
  NANDN U26151 ( .A(n19481), .B(ereg[105]), .Z(n19901) );
  NAND U26152 ( .A(n19903), .B(n19904), .Z(n15271) );
  NANDN U26153 ( .A(init), .B(e[106]), .Z(n19904) );
  AND U26154 ( .A(n19905), .B(n19906), .Z(n19903) );
  NAND U26155 ( .A(ereg[105]), .B(n19486), .Z(n19906) );
  NANDN U26156 ( .A(n19481), .B(ereg[106]), .Z(n19905) );
  NAND U26157 ( .A(n19907), .B(n19908), .Z(n15270) );
  NANDN U26158 ( .A(init), .B(e[107]), .Z(n19908) );
  AND U26159 ( .A(n19909), .B(n19910), .Z(n19907) );
  NAND U26160 ( .A(ereg[106]), .B(n19486), .Z(n19910) );
  NANDN U26161 ( .A(n19481), .B(ereg[107]), .Z(n19909) );
  NAND U26162 ( .A(n19911), .B(n19912), .Z(n15269) );
  NANDN U26163 ( .A(init), .B(e[108]), .Z(n19912) );
  AND U26164 ( .A(n19913), .B(n19914), .Z(n19911) );
  NAND U26165 ( .A(ereg[107]), .B(n19486), .Z(n19914) );
  NANDN U26166 ( .A(n19481), .B(ereg[108]), .Z(n19913) );
  NAND U26167 ( .A(n19915), .B(n19916), .Z(n15268) );
  NANDN U26168 ( .A(init), .B(e[109]), .Z(n19916) );
  AND U26169 ( .A(n19917), .B(n19918), .Z(n19915) );
  NAND U26170 ( .A(ereg[108]), .B(n19486), .Z(n19918) );
  NANDN U26171 ( .A(n19481), .B(ereg[109]), .Z(n19917) );
  NAND U26172 ( .A(n19919), .B(n19920), .Z(n15267) );
  NANDN U26173 ( .A(init), .B(e[110]), .Z(n19920) );
  AND U26174 ( .A(n19921), .B(n19922), .Z(n19919) );
  NAND U26175 ( .A(ereg[109]), .B(n19486), .Z(n19922) );
  NANDN U26176 ( .A(n19481), .B(ereg[110]), .Z(n19921) );
  NAND U26177 ( .A(n19923), .B(n19924), .Z(n15266) );
  NANDN U26178 ( .A(init), .B(e[111]), .Z(n19924) );
  AND U26179 ( .A(n19925), .B(n19926), .Z(n19923) );
  NAND U26180 ( .A(ereg[110]), .B(n19486), .Z(n19926) );
  NANDN U26181 ( .A(n19481), .B(ereg[111]), .Z(n19925) );
  NAND U26182 ( .A(n19927), .B(n19928), .Z(n15265) );
  NANDN U26183 ( .A(init), .B(e[112]), .Z(n19928) );
  AND U26184 ( .A(n19929), .B(n19930), .Z(n19927) );
  NAND U26185 ( .A(ereg[111]), .B(n19486), .Z(n19930) );
  NANDN U26186 ( .A(n19481), .B(ereg[112]), .Z(n19929) );
  NAND U26187 ( .A(n19931), .B(n19932), .Z(n15264) );
  NANDN U26188 ( .A(init), .B(e[113]), .Z(n19932) );
  AND U26189 ( .A(n19933), .B(n19934), .Z(n19931) );
  NAND U26190 ( .A(ereg[112]), .B(n19486), .Z(n19934) );
  NANDN U26191 ( .A(n19481), .B(ereg[113]), .Z(n19933) );
  NAND U26192 ( .A(n19935), .B(n19936), .Z(n15263) );
  NANDN U26193 ( .A(init), .B(e[114]), .Z(n19936) );
  AND U26194 ( .A(n19937), .B(n19938), .Z(n19935) );
  NAND U26195 ( .A(ereg[113]), .B(n19486), .Z(n19938) );
  NANDN U26196 ( .A(n19481), .B(ereg[114]), .Z(n19937) );
  NAND U26197 ( .A(n19939), .B(n19940), .Z(n15262) );
  NANDN U26198 ( .A(init), .B(e[115]), .Z(n19940) );
  AND U26199 ( .A(n19941), .B(n19942), .Z(n19939) );
  NAND U26200 ( .A(ereg[114]), .B(n19486), .Z(n19942) );
  NANDN U26201 ( .A(n19481), .B(ereg[115]), .Z(n19941) );
  NAND U26202 ( .A(n19943), .B(n19944), .Z(n15261) );
  NANDN U26203 ( .A(init), .B(e[116]), .Z(n19944) );
  AND U26204 ( .A(n19945), .B(n19946), .Z(n19943) );
  NAND U26205 ( .A(ereg[115]), .B(n19486), .Z(n19946) );
  NANDN U26206 ( .A(n19481), .B(ereg[116]), .Z(n19945) );
  NAND U26207 ( .A(n19947), .B(n19948), .Z(n15260) );
  NANDN U26208 ( .A(init), .B(e[117]), .Z(n19948) );
  AND U26209 ( .A(n19949), .B(n19950), .Z(n19947) );
  NAND U26210 ( .A(ereg[116]), .B(n19486), .Z(n19950) );
  NANDN U26211 ( .A(n19481), .B(ereg[117]), .Z(n19949) );
  NAND U26212 ( .A(n19951), .B(n19952), .Z(n15259) );
  NANDN U26213 ( .A(init), .B(e[118]), .Z(n19952) );
  AND U26214 ( .A(n19953), .B(n19954), .Z(n19951) );
  NAND U26215 ( .A(ereg[117]), .B(n19486), .Z(n19954) );
  NANDN U26216 ( .A(n19481), .B(ereg[118]), .Z(n19953) );
  NAND U26217 ( .A(n19955), .B(n19956), .Z(n15258) );
  NANDN U26218 ( .A(init), .B(e[119]), .Z(n19956) );
  AND U26219 ( .A(n19957), .B(n19958), .Z(n19955) );
  NAND U26220 ( .A(ereg[118]), .B(n19486), .Z(n19958) );
  NANDN U26221 ( .A(n19481), .B(ereg[119]), .Z(n19957) );
  NAND U26222 ( .A(n19959), .B(n19960), .Z(n15257) );
  NANDN U26223 ( .A(init), .B(e[120]), .Z(n19960) );
  AND U26224 ( .A(n19961), .B(n19962), .Z(n19959) );
  NAND U26225 ( .A(ereg[119]), .B(n19486), .Z(n19962) );
  NANDN U26226 ( .A(n19481), .B(ereg[120]), .Z(n19961) );
  NAND U26227 ( .A(n19963), .B(n19964), .Z(n15256) );
  NANDN U26228 ( .A(init), .B(e[121]), .Z(n19964) );
  AND U26229 ( .A(n19965), .B(n19966), .Z(n19963) );
  NAND U26230 ( .A(ereg[120]), .B(n19486), .Z(n19966) );
  NANDN U26231 ( .A(n19481), .B(ereg[121]), .Z(n19965) );
  NAND U26232 ( .A(n19967), .B(n19968), .Z(n15255) );
  NANDN U26233 ( .A(init), .B(e[122]), .Z(n19968) );
  AND U26234 ( .A(n19969), .B(n19970), .Z(n19967) );
  NAND U26235 ( .A(ereg[121]), .B(n19486), .Z(n19970) );
  NANDN U26236 ( .A(n19481), .B(ereg[122]), .Z(n19969) );
  NAND U26237 ( .A(n19971), .B(n19972), .Z(n15254) );
  NANDN U26238 ( .A(init), .B(e[123]), .Z(n19972) );
  AND U26239 ( .A(n19973), .B(n19974), .Z(n19971) );
  NAND U26240 ( .A(ereg[122]), .B(n19486), .Z(n19974) );
  NANDN U26241 ( .A(n19481), .B(ereg[123]), .Z(n19973) );
  NAND U26242 ( .A(n19975), .B(n19976), .Z(n15253) );
  NANDN U26243 ( .A(init), .B(e[124]), .Z(n19976) );
  AND U26244 ( .A(n19977), .B(n19978), .Z(n19975) );
  NAND U26245 ( .A(ereg[123]), .B(n19486), .Z(n19978) );
  NANDN U26246 ( .A(n19481), .B(ereg[124]), .Z(n19977) );
  NAND U26247 ( .A(n19979), .B(n19980), .Z(n15252) );
  NANDN U26248 ( .A(init), .B(e[125]), .Z(n19980) );
  AND U26249 ( .A(n19981), .B(n19982), .Z(n19979) );
  NAND U26250 ( .A(ereg[124]), .B(n19486), .Z(n19982) );
  NANDN U26251 ( .A(n19481), .B(ereg[125]), .Z(n19981) );
  NAND U26252 ( .A(n19983), .B(n19984), .Z(n15251) );
  NANDN U26253 ( .A(init), .B(e[126]), .Z(n19984) );
  AND U26254 ( .A(n19985), .B(n19986), .Z(n19983) );
  NAND U26255 ( .A(ereg[125]), .B(n19486), .Z(n19986) );
  NANDN U26256 ( .A(n19481), .B(ereg[126]), .Z(n19985) );
  NAND U26257 ( .A(n19987), .B(n19988), .Z(n15250) );
  NANDN U26258 ( .A(init), .B(e[127]), .Z(n19988) );
  AND U26259 ( .A(n19989), .B(n19990), .Z(n19987) );
  NAND U26260 ( .A(ereg[126]), .B(n19486), .Z(n19990) );
  NANDN U26261 ( .A(n19481), .B(ereg[127]), .Z(n19989) );
  NAND U26262 ( .A(n19991), .B(n19992), .Z(n15249) );
  NANDN U26263 ( .A(init), .B(e[128]), .Z(n19992) );
  AND U26264 ( .A(n19993), .B(n19994), .Z(n19991) );
  NAND U26265 ( .A(ereg[127]), .B(n19486), .Z(n19994) );
  NANDN U26266 ( .A(n19481), .B(ereg[128]), .Z(n19993) );
  NAND U26267 ( .A(n19995), .B(n19996), .Z(n15248) );
  NANDN U26268 ( .A(init), .B(e[129]), .Z(n19996) );
  AND U26269 ( .A(n19997), .B(n19998), .Z(n19995) );
  NAND U26270 ( .A(ereg[128]), .B(n19486), .Z(n19998) );
  NANDN U26271 ( .A(n19481), .B(ereg[129]), .Z(n19997) );
  NAND U26272 ( .A(n19999), .B(n20000), .Z(n15247) );
  NANDN U26273 ( .A(init), .B(e[130]), .Z(n20000) );
  AND U26274 ( .A(n20001), .B(n20002), .Z(n19999) );
  NAND U26275 ( .A(ereg[129]), .B(n19486), .Z(n20002) );
  NANDN U26276 ( .A(n19481), .B(ereg[130]), .Z(n20001) );
  NAND U26277 ( .A(n20003), .B(n20004), .Z(n15246) );
  NANDN U26278 ( .A(init), .B(e[131]), .Z(n20004) );
  AND U26279 ( .A(n20005), .B(n20006), .Z(n20003) );
  NAND U26280 ( .A(ereg[130]), .B(n19486), .Z(n20006) );
  NANDN U26281 ( .A(n19481), .B(ereg[131]), .Z(n20005) );
  NAND U26282 ( .A(n20007), .B(n20008), .Z(n15245) );
  NANDN U26283 ( .A(init), .B(e[132]), .Z(n20008) );
  AND U26284 ( .A(n20009), .B(n20010), .Z(n20007) );
  NAND U26285 ( .A(ereg[131]), .B(n19486), .Z(n20010) );
  NANDN U26286 ( .A(n19481), .B(ereg[132]), .Z(n20009) );
  NAND U26287 ( .A(n20011), .B(n20012), .Z(n15244) );
  NANDN U26288 ( .A(init), .B(e[133]), .Z(n20012) );
  AND U26289 ( .A(n20013), .B(n20014), .Z(n20011) );
  NAND U26290 ( .A(ereg[132]), .B(n19486), .Z(n20014) );
  NANDN U26291 ( .A(n19481), .B(ereg[133]), .Z(n20013) );
  NAND U26292 ( .A(n20015), .B(n20016), .Z(n15243) );
  NANDN U26293 ( .A(init), .B(e[134]), .Z(n20016) );
  AND U26294 ( .A(n20017), .B(n20018), .Z(n20015) );
  NAND U26295 ( .A(ereg[133]), .B(n19486), .Z(n20018) );
  NANDN U26296 ( .A(n19481), .B(ereg[134]), .Z(n20017) );
  NAND U26297 ( .A(n20019), .B(n20020), .Z(n15242) );
  NANDN U26298 ( .A(init), .B(e[135]), .Z(n20020) );
  AND U26299 ( .A(n20021), .B(n20022), .Z(n20019) );
  NAND U26300 ( .A(ereg[134]), .B(n19486), .Z(n20022) );
  NANDN U26301 ( .A(n19481), .B(ereg[135]), .Z(n20021) );
  NAND U26302 ( .A(n20023), .B(n20024), .Z(n15241) );
  NANDN U26303 ( .A(init), .B(e[136]), .Z(n20024) );
  AND U26304 ( .A(n20025), .B(n20026), .Z(n20023) );
  NAND U26305 ( .A(ereg[135]), .B(n19486), .Z(n20026) );
  NANDN U26306 ( .A(n19481), .B(ereg[136]), .Z(n20025) );
  NAND U26307 ( .A(n20027), .B(n20028), .Z(n15240) );
  NANDN U26308 ( .A(init), .B(e[137]), .Z(n20028) );
  AND U26309 ( .A(n20029), .B(n20030), .Z(n20027) );
  NAND U26310 ( .A(ereg[136]), .B(n19486), .Z(n20030) );
  NANDN U26311 ( .A(n19481), .B(ereg[137]), .Z(n20029) );
  NAND U26312 ( .A(n20031), .B(n20032), .Z(n15239) );
  NANDN U26313 ( .A(init), .B(e[138]), .Z(n20032) );
  AND U26314 ( .A(n20033), .B(n20034), .Z(n20031) );
  NAND U26315 ( .A(ereg[137]), .B(n19486), .Z(n20034) );
  NANDN U26316 ( .A(n19481), .B(ereg[138]), .Z(n20033) );
  NAND U26317 ( .A(n20035), .B(n20036), .Z(n15238) );
  NANDN U26318 ( .A(init), .B(e[139]), .Z(n20036) );
  AND U26319 ( .A(n20037), .B(n20038), .Z(n20035) );
  NAND U26320 ( .A(ereg[138]), .B(n19486), .Z(n20038) );
  NANDN U26321 ( .A(n19481), .B(ereg[139]), .Z(n20037) );
  NAND U26322 ( .A(n20039), .B(n20040), .Z(n15237) );
  NANDN U26323 ( .A(init), .B(e[140]), .Z(n20040) );
  AND U26324 ( .A(n20041), .B(n20042), .Z(n20039) );
  NAND U26325 ( .A(ereg[139]), .B(n19486), .Z(n20042) );
  NANDN U26326 ( .A(n19481), .B(ereg[140]), .Z(n20041) );
  NAND U26327 ( .A(n20043), .B(n20044), .Z(n15236) );
  NANDN U26328 ( .A(init), .B(e[141]), .Z(n20044) );
  AND U26329 ( .A(n20045), .B(n20046), .Z(n20043) );
  NAND U26330 ( .A(ereg[140]), .B(n19486), .Z(n20046) );
  NANDN U26331 ( .A(n19481), .B(ereg[141]), .Z(n20045) );
  NAND U26332 ( .A(n20047), .B(n20048), .Z(n15235) );
  NANDN U26333 ( .A(init), .B(e[142]), .Z(n20048) );
  AND U26334 ( .A(n20049), .B(n20050), .Z(n20047) );
  NAND U26335 ( .A(ereg[141]), .B(n19486), .Z(n20050) );
  NANDN U26336 ( .A(n19481), .B(ereg[142]), .Z(n20049) );
  NAND U26337 ( .A(n20051), .B(n20052), .Z(n15234) );
  NANDN U26338 ( .A(init), .B(e[143]), .Z(n20052) );
  AND U26339 ( .A(n20053), .B(n20054), .Z(n20051) );
  NAND U26340 ( .A(ereg[142]), .B(n19486), .Z(n20054) );
  NANDN U26341 ( .A(n19481), .B(ereg[143]), .Z(n20053) );
  NAND U26342 ( .A(n20055), .B(n20056), .Z(n15233) );
  NANDN U26343 ( .A(init), .B(e[144]), .Z(n20056) );
  AND U26344 ( .A(n20057), .B(n20058), .Z(n20055) );
  NAND U26345 ( .A(ereg[143]), .B(n19486), .Z(n20058) );
  NANDN U26346 ( .A(n19481), .B(ereg[144]), .Z(n20057) );
  NAND U26347 ( .A(n20059), .B(n20060), .Z(n15232) );
  NANDN U26348 ( .A(init), .B(e[145]), .Z(n20060) );
  AND U26349 ( .A(n20061), .B(n20062), .Z(n20059) );
  NAND U26350 ( .A(ereg[144]), .B(n19486), .Z(n20062) );
  NANDN U26351 ( .A(n19481), .B(ereg[145]), .Z(n20061) );
  NAND U26352 ( .A(n20063), .B(n20064), .Z(n15231) );
  NANDN U26353 ( .A(init), .B(e[146]), .Z(n20064) );
  AND U26354 ( .A(n20065), .B(n20066), .Z(n20063) );
  NAND U26355 ( .A(ereg[145]), .B(n19486), .Z(n20066) );
  NANDN U26356 ( .A(n19481), .B(ereg[146]), .Z(n20065) );
  NAND U26357 ( .A(n20067), .B(n20068), .Z(n15230) );
  NANDN U26358 ( .A(init), .B(e[147]), .Z(n20068) );
  AND U26359 ( .A(n20069), .B(n20070), .Z(n20067) );
  NAND U26360 ( .A(ereg[146]), .B(n19486), .Z(n20070) );
  NANDN U26361 ( .A(n19481), .B(ereg[147]), .Z(n20069) );
  NAND U26362 ( .A(n20071), .B(n20072), .Z(n15229) );
  NANDN U26363 ( .A(init), .B(e[148]), .Z(n20072) );
  AND U26364 ( .A(n20073), .B(n20074), .Z(n20071) );
  NAND U26365 ( .A(ereg[147]), .B(n19486), .Z(n20074) );
  NANDN U26366 ( .A(n19481), .B(ereg[148]), .Z(n20073) );
  NAND U26367 ( .A(n20075), .B(n20076), .Z(n15228) );
  NANDN U26368 ( .A(init), .B(e[149]), .Z(n20076) );
  AND U26369 ( .A(n20077), .B(n20078), .Z(n20075) );
  NAND U26370 ( .A(ereg[148]), .B(n19486), .Z(n20078) );
  NANDN U26371 ( .A(n19481), .B(ereg[149]), .Z(n20077) );
  NAND U26372 ( .A(n20079), .B(n20080), .Z(n15227) );
  NANDN U26373 ( .A(init), .B(e[150]), .Z(n20080) );
  AND U26374 ( .A(n20081), .B(n20082), .Z(n20079) );
  NAND U26375 ( .A(ereg[149]), .B(n19486), .Z(n20082) );
  NANDN U26376 ( .A(n19481), .B(ereg[150]), .Z(n20081) );
  NAND U26377 ( .A(n20083), .B(n20084), .Z(n15226) );
  NANDN U26378 ( .A(init), .B(e[151]), .Z(n20084) );
  AND U26379 ( .A(n20085), .B(n20086), .Z(n20083) );
  NAND U26380 ( .A(ereg[150]), .B(n19486), .Z(n20086) );
  NANDN U26381 ( .A(n19481), .B(ereg[151]), .Z(n20085) );
  NAND U26382 ( .A(n20087), .B(n20088), .Z(n15225) );
  NANDN U26383 ( .A(init), .B(e[152]), .Z(n20088) );
  AND U26384 ( .A(n20089), .B(n20090), .Z(n20087) );
  NAND U26385 ( .A(ereg[151]), .B(n19486), .Z(n20090) );
  NANDN U26386 ( .A(n19481), .B(ereg[152]), .Z(n20089) );
  NAND U26387 ( .A(n20091), .B(n20092), .Z(n15224) );
  NANDN U26388 ( .A(init), .B(e[153]), .Z(n20092) );
  AND U26389 ( .A(n20093), .B(n20094), .Z(n20091) );
  NAND U26390 ( .A(ereg[152]), .B(n19486), .Z(n20094) );
  NANDN U26391 ( .A(n19481), .B(ereg[153]), .Z(n20093) );
  NAND U26392 ( .A(n20095), .B(n20096), .Z(n15223) );
  NANDN U26393 ( .A(init), .B(e[154]), .Z(n20096) );
  AND U26394 ( .A(n20097), .B(n20098), .Z(n20095) );
  NAND U26395 ( .A(ereg[153]), .B(n19486), .Z(n20098) );
  NANDN U26396 ( .A(n19481), .B(ereg[154]), .Z(n20097) );
  NAND U26397 ( .A(n20099), .B(n20100), .Z(n15222) );
  NANDN U26398 ( .A(init), .B(e[155]), .Z(n20100) );
  AND U26399 ( .A(n20101), .B(n20102), .Z(n20099) );
  NAND U26400 ( .A(ereg[154]), .B(n19486), .Z(n20102) );
  NANDN U26401 ( .A(n19481), .B(ereg[155]), .Z(n20101) );
  NAND U26402 ( .A(n20103), .B(n20104), .Z(n15221) );
  NANDN U26403 ( .A(init), .B(e[156]), .Z(n20104) );
  AND U26404 ( .A(n20105), .B(n20106), .Z(n20103) );
  NAND U26405 ( .A(ereg[155]), .B(n19486), .Z(n20106) );
  NANDN U26406 ( .A(n19481), .B(ereg[156]), .Z(n20105) );
  NAND U26407 ( .A(n20107), .B(n20108), .Z(n15220) );
  NANDN U26408 ( .A(init), .B(e[157]), .Z(n20108) );
  AND U26409 ( .A(n20109), .B(n20110), .Z(n20107) );
  NAND U26410 ( .A(ereg[156]), .B(n19486), .Z(n20110) );
  NANDN U26411 ( .A(n19481), .B(ereg[157]), .Z(n20109) );
  NAND U26412 ( .A(n20111), .B(n20112), .Z(n15219) );
  NANDN U26413 ( .A(init), .B(e[158]), .Z(n20112) );
  AND U26414 ( .A(n20113), .B(n20114), .Z(n20111) );
  NAND U26415 ( .A(ereg[157]), .B(n19486), .Z(n20114) );
  NANDN U26416 ( .A(n19481), .B(ereg[158]), .Z(n20113) );
  NAND U26417 ( .A(n20115), .B(n20116), .Z(n15218) );
  NANDN U26418 ( .A(init), .B(e[159]), .Z(n20116) );
  AND U26419 ( .A(n20117), .B(n20118), .Z(n20115) );
  NAND U26420 ( .A(ereg[158]), .B(n19486), .Z(n20118) );
  NANDN U26421 ( .A(n19481), .B(ereg[159]), .Z(n20117) );
  NAND U26422 ( .A(n20119), .B(n20120), .Z(n15217) );
  NANDN U26423 ( .A(init), .B(e[160]), .Z(n20120) );
  AND U26424 ( .A(n20121), .B(n20122), .Z(n20119) );
  NAND U26425 ( .A(ereg[159]), .B(n19486), .Z(n20122) );
  NANDN U26426 ( .A(n19481), .B(ereg[160]), .Z(n20121) );
  NAND U26427 ( .A(n20123), .B(n20124), .Z(n15216) );
  NANDN U26428 ( .A(init), .B(e[161]), .Z(n20124) );
  AND U26429 ( .A(n20125), .B(n20126), .Z(n20123) );
  NAND U26430 ( .A(ereg[160]), .B(n19486), .Z(n20126) );
  NANDN U26431 ( .A(n19481), .B(ereg[161]), .Z(n20125) );
  NAND U26432 ( .A(n20127), .B(n20128), .Z(n15215) );
  NANDN U26433 ( .A(init), .B(e[162]), .Z(n20128) );
  AND U26434 ( .A(n20129), .B(n20130), .Z(n20127) );
  NAND U26435 ( .A(ereg[161]), .B(n19486), .Z(n20130) );
  NANDN U26436 ( .A(n19481), .B(ereg[162]), .Z(n20129) );
  NAND U26437 ( .A(n20131), .B(n20132), .Z(n15214) );
  NANDN U26438 ( .A(init), .B(e[163]), .Z(n20132) );
  AND U26439 ( .A(n20133), .B(n20134), .Z(n20131) );
  NAND U26440 ( .A(ereg[162]), .B(n19486), .Z(n20134) );
  NANDN U26441 ( .A(n19481), .B(ereg[163]), .Z(n20133) );
  NAND U26442 ( .A(n20135), .B(n20136), .Z(n15213) );
  NANDN U26443 ( .A(init), .B(e[164]), .Z(n20136) );
  AND U26444 ( .A(n20137), .B(n20138), .Z(n20135) );
  NAND U26445 ( .A(ereg[163]), .B(n19486), .Z(n20138) );
  NANDN U26446 ( .A(n19481), .B(ereg[164]), .Z(n20137) );
  NAND U26447 ( .A(n20139), .B(n20140), .Z(n15212) );
  NANDN U26448 ( .A(init), .B(e[165]), .Z(n20140) );
  AND U26449 ( .A(n20141), .B(n20142), .Z(n20139) );
  NAND U26450 ( .A(ereg[164]), .B(n19486), .Z(n20142) );
  NANDN U26451 ( .A(n19481), .B(ereg[165]), .Z(n20141) );
  NAND U26452 ( .A(n20143), .B(n20144), .Z(n15211) );
  NANDN U26453 ( .A(init), .B(e[166]), .Z(n20144) );
  AND U26454 ( .A(n20145), .B(n20146), .Z(n20143) );
  NAND U26455 ( .A(ereg[165]), .B(n19486), .Z(n20146) );
  NANDN U26456 ( .A(n19481), .B(ereg[166]), .Z(n20145) );
  NAND U26457 ( .A(n20147), .B(n20148), .Z(n15210) );
  NANDN U26458 ( .A(init), .B(e[167]), .Z(n20148) );
  AND U26459 ( .A(n20149), .B(n20150), .Z(n20147) );
  NAND U26460 ( .A(ereg[166]), .B(n19486), .Z(n20150) );
  NANDN U26461 ( .A(n19481), .B(ereg[167]), .Z(n20149) );
  NAND U26462 ( .A(n20151), .B(n20152), .Z(n15209) );
  NANDN U26463 ( .A(init), .B(e[168]), .Z(n20152) );
  AND U26464 ( .A(n20153), .B(n20154), .Z(n20151) );
  NAND U26465 ( .A(ereg[167]), .B(n19486), .Z(n20154) );
  NANDN U26466 ( .A(n19481), .B(ereg[168]), .Z(n20153) );
  NAND U26467 ( .A(n20155), .B(n20156), .Z(n15208) );
  NANDN U26468 ( .A(init), .B(e[169]), .Z(n20156) );
  AND U26469 ( .A(n20157), .B(n20158), .Z(n20155) );
  NAND U26470 ( .A(ereg[168]), .B(n19486), .Z(n20158) );
  NANDN U26471 ( .A(n19481), .B(ereg[169]), .Z(n20157) );
  NAND U26472 ( .A(n20159), .B(n20160), .Z(n15207) );
  NANDN U26473 ( .A(init), .B(e[170]), .Z(n20160) );
  AND U26474 ( .A(n20161), .B(n20162), .Z(n20159) );
  NAND U26475 ( .A(ereg[169]), .B(n19486), .Z(n20162) );
  NANDN U26476 ( .A(n19481), .B(ereg[170]), .Z(n20161) );
  NAND U26477 ( .A(n20163), .B(n20164), .Z(n15206) );
  NANDN U26478 ( .A(init), .B(e[171]), .Z(n20164) );
  AND U26479 ( .A(n20165), .B(n20166), .Z(n20163) );
  NAND U26480 ( .A(ereg[170]), .B(n19486), .Z(n20166) );
  NANDN U26481 ( .A(n19481), .B(ereg[171]), .Z(n20165) );
  NAND U26482 ( .A(n20167), .B(n20168), .Z(n15205) );
  NANDN U26483 ( .A(init), .B(e[172]), .Z(n20168) );
  AND U26484 ( .A(n20169), .B(n20170), .Z(n20167) );
  NAND U26485 ( .A(ereg[171]), .B(n19486), .Z(n20170) );
  NANDN U26486 ( .A(n19481), .B(ereg[172]), .Z(n20169) );
  NAND U26487 ( .A(n20171), .B(n20172), .Z(n15204) );
  NANDN U26488 ( .A(init), .B(e[173]), .Z(n20172) );
  AND U26489 ( .A(n20173), .B(n20174), .Z(n20171) );
  NAND U26490 ( .A(ereg[172]), .B(n19486), .Z(n20174) );
  NANDN U26491 ( .A(n19481), .B(ereg[173]), .Z(n20173) );
  NAND U26492 ( .A(n20175), .B(n20176), .Z(n15203) );
  NANDN U26493 ( .A(init), .B(e[174]), .Z(n20176) );
  AND U26494 ( .A(n20177), .B(n20178), .Z(n20175) );
  NAND U26495 ( .A(ereg[173]), .B(n19486), .Z(n20178) );
  NANDN U26496 ( .A(n19481), .B(ereg[174]), .Z(n20177) );
  NAND U26497 ( .A(n20179), .B(n20180), .Z(n15202) );
  NANDN U26498 ( .A(init), .B(e[175]), .Z(n20180) );
  AND U26499 ( .A(n20181), .B(n20182), .Z(n20179) );
  NAND U26500 ( .A(ereg[174]), .B(n19486), .Z(n20182) );
  NANDN U26501 ( .A(n19481), .B(ereg[175]), .Z(n20181) );
  NAND U26502 ( .A(n20183), .B(n20184), .Z(n15201) );
  NANDN U26503 ( .A(init), .B(e[176]), .Z(n20184) );
  AND U26504 ( .A(n20185), .B(n20186), .Z(n20183) );
  NAND U26505 ( .A(ereg[175]), .B(n19486), .Z(n20186) );
  NANDN U26506 ( .A(n19481), .B(ereg[176]), .Z(n20185) );
  NAND U26507 ( .A(n20187), .B(n20188), .Z(n15200) );
  NANDN U26508 ( .A(init), .B(e[177]), .Z(n20188) );
  AND U26509 ( .A(n20189), .B(n20190), .Z(n20187) );
  NAND U26510 ( .A(ereg[176]), .B(n19486), .Z(n20190) );
  NANDN U26511 ( .A(n19481), .B(ereg[177]), .Z(n20189) );
  NAND U26512 ( .A(n20191), .B(n20192), .Z(n15199) );
  NANDN U26513 ( .A(init), .B(e[178]), .Z(n20192) );
  AND U26514 ( .A(n20193), .B(n20194), .Z(n20191) );
  NAND U26515 ( .A(ereg[177]), .B(n19486), .Z(n20194) );
  NANDN U26516 ( .A(n19481), .B(ereg[178]), .Z(n20193) );
  NAND U26517 ( .A(n20195), .B(n20196), .Z(n15198) );
  NANDN U26518 ( .A(init), .B(e[179]), .Z(n20196) );
  AND U26519 ( .A(n20197), .B(n20198), .Z(n20195) );
  NAND U26520 ( .A(ereg[178]), .B(n19486), .Z(n20198) );
  NANDN U26521 ( .A(n19481), .B(ereg[179]), .Z(n20197) );
  NAND U26522 ( .A(n20199), .B(n20200), .Z(n15197) );
  NANDN U26523 ( .A(init), .B(e[180]), .Z(n20200) );
  AND U26524 ( .A(n20201), .B(n20202), .Z(n20199) );
  NAND U26525 ( .A(ereg[179]), .B(n19486), .Z(n20202) );
  NANDN U26526 ( .A(n19481), .B(ereg[180]), .Z(n20201) );
  NAND U26527 ( .A(n20203), .B(n20204), .Z(n15196) );
  NANDN U26528 ( .A(init), .B(e[181]), .Z(n20204) );
  AND U26529 ( .A(n20205), .B(n20206), .Z(n20203) );
  NAND U26530 ( .A(ereg[180]), .B(n19486), .Z(n20206) );
  NANDN U26531 ( .A(n19481), .B(ereg[181]), .Z(n20205) );
  NAND U26532 ( .A(n20207), .B(n20208), .Z(n15195) );
  NANDN U26533 ( .A(init), .B(e[182]), .Z(n20208) );
  AND U26534 ( .A(n20209), .B(n20210), .Z(n20207) );
  NAND U26535 ( .A(ereg[181]), .B(n19486), .Z(n20210) );
  NANDN U26536 ( .A(n19481), .B(ereg[182]), .Z(n20209) );
  NAND U26537 ( .A(n20211), .B(n20212), .Z(n15194) );
  NANDN U26538 ( .A(init), .B(e[183]), .Z(n20212) );
  AND U26539 ( .A(n20213), .B(n20214), .Z(n20211) );
  NAND U26540 ( .A(ereg[182]), .B(n19486), .Z(n20214) );
  NANDN U26541 ( .A(n19481), .B(ereg[183]), .Z(n20213) );
  NAND U26542 ( .A(n20215), .B(n20216), .Z(n15193) );
  NANDN U26543 ( .A(init), .B(e[184]), .Z(n20216) );
  AND U26544 ( .A(n20217), .B(n20218), .Z(n20215) );
  NAND U26545 ( .A(ereg[183]), .B(n19486), .Z(n20218) );
  NANDN U26546 ( .A(n19481), .B(ereg[184]), .Z(n20217) );
  NAND U26547 ( .A(n20219), .B(n20220), .Z(n15192) );
  NANDN U26548 ( .A(init), .B(e[185]), .Z(n20220) );
  AND U26549 ( .A(n20221), .B(n20222), .Z(n20219) );
  NAND U26550 ( .A(ereg[184]), .B(n19486), .Z(n20222) );
  NANDN U26551 ( .A(n19481), .B(ereg[185]), .Z(n20221) );
  NAND U26552 ( .A(n20223), .B(n20224), .Z(n15191) );
  NANDN U26553 ( .A(init), .B(e[186]), .Z(n20224) );
  AND U26554 ( .A(n20225), .B(n20226), .Z(n20223) );
  NAND U26555 ( .A(ereg[185]), .B(n19486), .Z(n20226) );
  NANDN U26556 ( .A(n19481), .B(ereg[186]), .Z(n20225) );
  NAND U26557 ( .A(n20227), .B(n20228), .Z(n15190) );
  NANDN U26558 ( .A(init), .B(e[187]), .Z(n20228) );
  AND U26559 ( .A(n20229), .B(n20230), .Z(n20227) );
  NAND U26560 ( .A(ereg[186]), .B(n19486), .Z(n20230) );
  NANDN U26561 ( .A(n19481), .B(ereg[187]), .Z(n20229) );
  NAND U26562 ( .A(n20231), .B(n20232), .Z(n15189) );
  NANDN U26563 ( .A(init), .B(e[188]), .Z(n20232) );
  AND U26564 ( .A(n20233), .B(n20234), .Z(n20231) );
  NAND U26565 ( .A(ereg[187]), .B(n19486), .Z(n20234) );
  NANDN U26566 ( .A(n19481), .B(ereg[188]), .Z(n20233) );
  NAND U26567 ( .A(n20235), .B(n20236), .Z(n15188) );
  NANDN U26568 ( .A(init), .B(e[189]), .Z(n20236) );
  AND U26569 ( .A(n20237), .B(n20238), .Z(n20235) );
  NAND U26570 ( .A(ereg[188]), .B(n19486), .Z(n20238) );
  NANDN U26571 ( .A(n19481), .B(ereg[189]), .Z(n20237) );
  NAND U26572 ( .A(n20239), .B(n20240), .Z(n15187) );
  NANDN U26573 ( .A(init), .B(e[190]), .Z(n20240) );
  AND U26574 ( .A(n20241), .B(n20242), .Z(n20239) );
  NAND U26575 ( .A(ereg[189]), .B(n19486), .Z(n20242) );
  NANDN U26576 ( .A(n19481), .B(ereg[190]), .Z(n20241) );
  NAND U26577 ( .A(n20243), .B(n20244), .Z(n15186) );
  NANDN U26578 ( .A(init), .B(e[191]), .Z(n20244) );
  AND U26579 ( .A(n20245), .B(n20246), .Z(n20243) );
  NAND U26580 ( .A(ereg[190]), .B(n19486), .Z(n20246) );
  NANDN U26581 ( .A(n19481), .B(ereg[191]), .Z(n20245) );
  NAND U26582 ( .A(n20247), .B(n20248), .Z(n15185) );
  NANDN U26583 ( .A(init), .B(e[192]), .Z(n20248) );
  AND U26584 ( .A(n20249), .B(n20250), .Z(n20247) );
  NAND U26585 ( .A(ereg[191]), .B(n19486), .Z(n20250) );
  NANDN U26586 ( .A(n19481), .B(ereg[192]), .Z(n20249) );
  NAND U26587 ( .A(n20251), .B(n20252), .Z(n15184) );
  NANDN U26588 ( .A(init), .B(e[193]), .Z(n20252) );
  AND U26589 ( .A(n20253), .B(n20254), .Z(n20251) );
  NAND U26590 ( .A(ereg[192]), .B(n19486), .Z(n20254) );
  NANDN U26591 ( .A(n19481), .B(ereg[193]), .Z(n20253) );
  NAND U26592 ( .A(n20255), .B(n20256), .Z(n15183) );
  NANDN U26593 ( .A(init), .B(e[194]), .Z(n20256) );
  AND U26594 ( .A(n20257), .B(n20258), .Z(n20255) );
  NAND U26595 ( .A(ereg[193]), .B(n19486), .Z(n20258) );
  NANDN U26596 ( .A(n19481), .B(ereg[194]), .Z(n20257) );
  NAND U26597 ( .A(n20259), .B(n20260), .Z(n15182) );
  NANDN U26598 ( .A(init), .B(e[195]), .Z(n20260) );
  AND U26599 ( .A(n20261), .B(n20262), .Z(n20259) );
  NAND U26600 ( .A(ereg[194]), .B(n19486), .Z(n20262) );
  NANDN U26601 ( .A(n19481), .B(ereg[195]), .Z(n20261) );
  NAND U26602 ( .A(n20263), .B(n20264), .Z(n15181) );
  NANDN U26603 ( .A(init), .B(e[196]), .Z(n20264) );
  AND U26604 ( .A(n20265), .B(n20266), .Z(n20263) );
  NAND U26605 ( .A(ereg[195]), .B(n19486), .Z(n20266) );
  NANDN U26606 ( .A(n19481), .B(ereg[196]), .Z(n20265) );
  NAND U26607 ( .A(n20267), .B(n20268), .Z(n15180) );
  NANDN U26608 ( .A(init), .B(e[197]), .Z(n20268) );
  AND U26609 ( .A(n20269), .B(n20270), .Z(n20267) );
  NAND U26610 ( .A(ereg[196]), .B(n19486), .Z(n20270) );
  NANDN U26611 ( .A(n19481), .B(ereg[197]), .Z(n20269) );
  NAND U26612 ( .A(n20271), .B(n20272), .Z(n15179) );
  NANDN U26613 ( .A(init), .B(e[198]), .Z(n20272) );
  AND U26614 ( .A(n20273), .B(n20274), .Z(n20271) );
  NAND U26615 ( .A(ereg[197]), .B(n19486), .Z(n20274) );
  NANDN U26616 ( .A(n19481), .B(ereg[198]), .Z(n20273) );
  NAND U26617 ( .A(n20275), .B(n20276), .Z(n15178) );
  NANDN U26618 ( .A(init), .B(e[199]), .Z(n20276) );
  AND U26619 ( .A(n20277), .B(n20278), .Z(n20275) );
  NAND U26620 ( .A(ereg[198]), .B(n19486), .Z(n20278) );
  NANDN U26621 ( .A(n19481), .B(ereg[199]), .Z(n20277) );
  NAND U26622 ( .A(n20279), .B(n20280), .Z(n15177) );
  NANDN U26623 ( .A(init), .B(e[200]), .Z(n20280) );
  AND U26624 ( .A(n20281), .B(n20282), .Z(n20279) );
  NAND U26625 ( .A(ereg[199]), .B(n19486), .Z(n20282) );
  NANDN U26626 ( .A(n19481), .B(ereg[200]), .Z(n20281) );
  NAND U26627 ( .A(n20283), .B(n20284), .Z(n15176) );
  NANDN U26628 ( .A(init), .B(e[201]), .Z(n20284) );
  AND U26629 ( .A(n20285), .B(n20286), .Z(n20283) );
  NAND U26630 ( .A(ereg[200]), .B(n19486), .Z(n20286) );
  NANDN U26631 ( .A(n19481), .B(ereg[201]), .Z(n20285) );
  NAND U26632 ( .A(n20287), .B(n20288), .Z(n15175) );
  NANDN U26633 ( .A(init), .B(e[202]), .Z(n20288) );
  AND U26634 ( .A(n20289), .B(n20290), .Z(n20287) );
  NAND U26635 ( .A(ereg[201]), .B(n19486), .Z(n20290) );
  NANDN U26636 ( .A(n19481), .B(ereg[202]), .Z(n20289) );
  NAND U26637 ( .A(n20291), .B(n20292), .Z(n15174) );
  NANDN U26638 ( .A(init), .B(e[203]), .Z(n20292) );
  AND U26639 ( .A(n20293), .B(n20294), .Z(n20291) );
  NAND U26640 ( .A(ereg[202]), .B(n19486), .Z(n20294) );
  NANDN U26641 ( .A(n19481), .B(ereg[203]), .Z(n20293) );
  NAND U26642 ( .A(n20295), .B(n20296), .Z(n15173) );
  NANDN U26643 ( .A(init), .B(e[204]), .Z(n20296) );
  AND U26644 ( .A(n20297), .B(n20298), .Z(n20295) );
  NAND U26645 ( .A(ereg[203]), .B(n19486), .Z(n20298) );
  NANDN U26646 ( .A(n19481), .B(ereg[204]), .Z(n20297) );
  NAND U26647 ( .A(n20299), .B(n20300), .Z(n15172) );
  NANDN U26648 ( .A(init), .B(e[205]), .Z(n20300) );
  AND U26649 ( .A(n20301), .B(n20302), .Z(n20299) );
  NAND U26650 ( .A(ereg[204]), .B(n19486), .Z(n20302) );
  NANDN U26651 ( .A(n19481), .B(ereg[205]), .Z(n20301) );
  NAND U26652 ( .A(n20303), .B(n20304), .Z(n15171) );
  NANDN U26653 ( .A(init), .B(e[206]), .Z(n20304) );
  AND U26654 ( .A(n20305), .B(n20306), .Z(n20303) );
  NAND U26655 ( .A(ereg[205]), .B(n19486), .Z(n20306) );
  NANDN U26656 ( .A(n19481), .B(ereg[206]), .Z(n20305) );
  NAND U26657 ( .A(n20307), .B(n20308), .Z(n15170) );
  NANDN U26658 ( .A(init), .B(e[207]), .Z(n20308) );
  AND U26659 ( .A(n20309), .B(n20310), .Z(n20307) );
  NAND U26660 ( .A(ereg[206]), .B(n19486), .Z(n20310) );
  NANDN U26661 ( .A(n19481), .B(ereg[207]), .Z(n20309) );
  NAND U26662 ( .A(n20311), .B(n20312), .Z(n15169) );
  NANDN U26663 ( .A(init), .B(e[208]), .Z(n20312) );
  AND U26664 ( .A(n20313), .B(n20314), .Z(n20311) );
  NAND U26665 ( .A(ereg[207]), .B(n19486), .Z(n20314) );
  NANDN U26666 ( .A(n19481), .B(ereg[208]), .Z(n20313) );
  NAND U26667 ( .A(n20315), .B(n20316), .Z(n15168) );
  NANDN U26668 ( .A(init), .B(e[209]), .Z(n20316) );
  AND U26669 ( .A(n20317), .B(n20318), .Z(n20315) );
  NAND U26670 ( .A(ereg[208]), .B(n19486), .Z(n20318) );
  NANDN U26671 ( .A(n19481), .B(ereg[209]), .Z(n20317) );
  NAND U26672 ( .A(n20319), .B(n20320), .Z(n15167) );
  NANDN U26673 ( .A(init), .B(e[210]), .Z(n20320) );
  AND U26674 ( .A(n20321), .B(n20322), .Z(n20319) );
  NAND U26675 ( .A(ereg[209]), .B(n19486), .Z(n20322) );
  NANDN U26676 ( .A(n19481), .B(ereg[210]), .Z(n20321) );
  NAND U26677 ( .A(n20323), .B(n20324), .Z(n15166) );
  NANDN U26678 ( .A(init), .B(e[211]), .Z(n20324) );
  AND U26679 ( .A(n20325), .B(n20326), .Z(n20323) );
  NAND U26680 ( .A(ereg[210]), .B(n19486), .Z(n20326) );
  NANDN U26681 ( .A(n19481), .B(ereg[211]), .Z(n20325) );
  NAND U26682 ( .A(n20327), .B(n20328), .Z(n15165) );
  NANDN U26683 ( .A(init), .B(e[212]), .Z(n20328) );
  AND U26684 ( .A(n20329), .B(n20330), .Z(n20327) );
  NAND U26685 ( .A(ereg[211]), .B(n19486), .Z(n20330) );
  NANDN U26686 ( .A(n19481), .B(ereg[212]), .Z(n20329) );
  NAND U26687 ( .A(n20331), .B(n20332), .Z(n15164) );
  NANDN U26688 ( .A(init), .B(e[213]), .Z(n20332) );
  AND U26689 ( .A(n20333), .B(n20334), .Z(n20331) );
  NAND U26690 ( .A(ereg[212]), .B(n19486), .Z(n20334) );
  NANDN U26691 ( .A(n19481), .B(ereg[213]), .Z(n20333) );
  NAND U26692 ( .A(n20335), .B(n20336), .Z(n15163) );
  NANDN U26693 ( .A(init), .B(e[214]), .Z(n20336) );
  AND U26694 ( .A(n20337), .B(n20338), .Z(n20335) );
  NAND U26695 ( .A(ereg[213]), .B(n19486), .Z(n20338) );
  NANDN U26696 ( .A(n19481), .B(ereg[214]), .Z(n20337) );
  NAND U26697 ( .A(n20339), .B(n20340), .Z(n15162) );
  NANDN U26698 ( .A(init), .B(e[215]), .Z(n20340) );
  AND U26699 ( .A(n20341), .B(n20342), .Z(n20339) );
  NAND U26700 ( .A(ereg[214]), .B(n19486), .Z(n20342) );
  NANDN U26701 ( .A(n19481), .B(ereg[215]), .Z(n20341) );
  NAND U26702 ( .A(n20343), .B(n20344), .Z(n15161) );
  NANDN U26703 ( .A(init), .B(e[216]), .Z(n20344) );
  AND U26704 ( .A(n20345), .B(n20346), .Z(n20343) );
  NAND U26705 ( .A(ereg[215]), .B(n19486), .Z(n20346) );
  NANDN U26706 ( .A(n19481), .B(ereg[216]), .Z(n20345) );
  NAND U26707 ( .A(n20347), .B(n20348), .Z(n15160) );
  NANDN U26708 ( .A(init), .B(e[217]), .Z(n20348) );
  AND U26709 ( .A(n20349), .B(n20350), .Z(n20347) );
  NAND U26710 ( .A(ereg[216]), .B(n19486), .Z(n20350) );
  NANDN U26711 ( .A(n19481), .B(ereg[217]), .Z(n20349) );
  NAND U26712 ( .A(n20351), .B(n20352), .Z(n15159) );
  NANDN U26713 ( .A(init), .B(e[218]), .Z(n20352) );
  AND U26714 ( .A(n20353), .B(n20354), .Z(n20351) );
  NAND U26715 ( .A(ereg[217]), .B(n19486), .Z(n20354) );
  NANDN U26716 ( .A(n19481), .B(ereg[218]), .Z(n20353) );
  NAND U26717 ( .A(n20355), .B(n20356), .Z(n15158) );
  NANDN U26718 ( .A(init), .B(e[219]), .Z(n20356) );
  AND U26719 ( .A(n20357), .B(n20358), .Z(n20355) );
  NAND U26720 ( .A(ereg[218]), .B(n19486), .Z(n20358) );
  NANDN U26721 ( .A(n19481), .B(ereg[219]), .Z(n20357) );
  NAND U26722 ( .A(n20359), .B(n20360), .Z(n15157) );
  NANDN U26723 ( .A(init), .B(e[220]), .Z(n20360) );
  AND U26724 ( .A(n20361), .B(n20362), .Z(n20359) );
  NAND U26725 ( .A(ereg[219]), .B(n19486), .Z(n20362) );
  NANDN U26726 ( .A(n19481), .B(ereg[220]), .Z(n20361) );
  NAND U26727 ( .A(n20363), .B(n20364), .Z(n15156) );
  NANDN U26728 ( .A(init), .B(e[221]), .Z(n20364) );
  AND U26729 ( .A(n20365), .B(n20366), .Z(n20363) );
  NAND U26730 ( .A(ereg[220]), .B(n19486), .Z(n20366) );
  NANDN U26731 ( .A(n19481), .B(ereg[221]), .Z(n20365) );
  NAND U26732 ( .A(n20367), .B(n20368), .Z(n15155) );
  NANDN U26733 ( .A(init), .B(e[222]), .Z(n20368) );
  AND U26734 ( .A(n20369), .B(n20370), .Z(n20367) );
  NAND U26735 ( .A(ereg[221]), .B(n19486), .Z(n20370) );
  NANDN U26736 ( .A(n19481), .B(ereg[222]), .Z(n20369) );
  NAND U26737 ( .A(n20371), .B(n20372), .Z(n15154) );
  NANDN U26738 ( .A(init), .B(e[223]), .Z(n20372) );
  AND U26739 ( .A(n20373), .B(n20374), .Z(n20371) );
  NAND U26740 ( .A(ereg[222]), .B(n19486), .Z(n20374) );
  NANDN U26741 ( .A(n19481), .B(ereg[223]), .Z(n20373) );
  NAND U26742 ( .A(n20375), .B(n20376), .Z(n15153) );
  NANDN U26743 ( .A(init), .B(e[224]), .Z(n20376) );
  AND U26744 ( .A(n20377), .B(n20378), .Z(n20375) );
  NAND U26745 ( .A(ereg[223]), .B(n19486), .Z(n20378) );
  NANDN U26746 ( .A(n19481), .B(ereg[224]), .Z(n20377) );
  NAND U26747 ( .A(n20379), .B(n20380), .Z(n15152) );
  NANDN U26748 ( .A(init), .B(e[225]), .Z(n20380) );
  AND U26749 ( .A(n20381), .B(n20382), .Z(n20379) );
  NAND U26750 ( .A(ereg[224]), .B(n19486), .Z(n20382) );
  NANDN U26751 ( .A(n19481), .B(ereg[225]), .Z(n20381) );
  NAND U26752 ( .A(n20383), .B(n20384), .Z(n15151) );
  NANDN U26753 ( .A(init), .B(e[226]), .Z(n20384) );
  AND U26754 ( .A(n20385), .B(n20386), .Z(n20383) );
  NAND U26755 ( .A(ereg[225]), .B(n19486), .Z(n20386) );
  NANDN U26756 ( .A(n19481), .B(ereg[226]), .Z(n20385) );
  NAND U26757 ( .A(n20387), .B(n20388), .Z(n15150) );
  NANDN U26758 ( .A(init), .B(e[227]), .Z(n20388) );
  AND U26759 ( .A(n20389), .B(n20390), .Z(n20387) );
  NAND U26760 ( .A(ereg[226]), .B(n19486), .Z(n20390) );
  NANDN U26761 ( .A(n19481), .B(ereg[227]), .Z(n20389) );
  NAND U26762 ( .A(n20391), .B(n20392), .Z(n15149) );
  NANDN U26763 ( .A(init), .B(e[228]), .Z(n20392) );
  AND U26764 ( .A(n20393), .B(n20394), .Z(n20391) );
  NAND U26765 ( .A(ereg[227]), .B(n19486), .Z(n20394) );
  NANDN U26766 ( .A(n19481), .B(ereg[228]), .Z(n20393) );
  NAND U26767 ( .A(n20395), .B(n20396), .Z(n15148) );
  NANDN U26768 ( .A(init), .B(e[229]), .Z(n20396) );
  AND U26769 ( .A(n20397), .B(n20398), .Z(n20395) );
  NAND U26770 ( .A(ereg[228]), .B(n19486), .Z(n20398) );
  NANDN U26771 ( .A(n19481), .B(ereg[229]), .Z(n20397) );
  NAND U26772 ( .A(n20399), .B(n20400), .Z(n15147) );
  NANDN U26773 ( .A(init), .B(e[230]), .Z(n20400) );
  AND U26774 ( .A(n20401), .B(n20402), .Z(n20399) );
  NAND U26775 ( .A(ereg[229]), .B(n19486), .Z(n20402) );
  NANDN U26776 ( .A(n19481), .B(ereg[230]), .Z(n20401) );
  NAND U26777 ( .A(n20403), .B(n20404), .Z(n15146) );
  NANDN U26778 ( .A(init), .B(e[231]), .Z(n20404) );
  AND U26779 ( .A(n20405), .B(n20406), .Z(n20403) );
  NAND U26780 ( .A(ereg[230]), .B(n19486), .Z(n20406) );
  NANDN U26781 ( .A(n19481), .B(ereg[231]), .Z(n20405) );
  NAND U26782 ( .A(n20407), .B(n20408), .Z(n15145) );
  NANDN U26783 ( .A(init), .B(e[232]), .Z(n20408) );
  AND U26784 ( .A(n20409), .B(n20410), .Z(n20407) );
  NAND U26785 ( .A(ereg[231]), .B(n19486), .Z(n20410) );
  NANDN U26786 ( .A(n19481), .B(ereg[232]), .Z(n20409) );
  NAND U26787 ( .A(n20411), .B(n20412), .Z(n15144) );
  NANDN U26788 ( .A(init), .B(e[233]), .Z(n20412) );
  AND U26789 ( .A(n20413), .B(n20414), .Z(n20411) );
  NAND U26790 ( .A(ereg[232]), .B(n19486), .Z(n20414) );
  NANDN U26791 ( .A(n19481), .B(ereg[233]), .Z(n20413) );
  NAND U26792 ( .A(n20415), .B(n20416), .Z(n15143) );
  NANDN U26793 ( .A(init), .B(e[234]), .Z(n20416) );
  AND U26794 ( .A(n20417), .B(n20418), .Z(n20415) );
  NAND U26795 ( .A(ereg[233]), .B(n19486), .Z(n20418) );
  NANDN U26796 ( .A(n19481), .B(ereg[234]), .Z(n20417) );
  NAND U26797 ( .A(n20419), .B(n20420), .Z(n15142) );
  NANDN U26798 ( .A(init), .B(e[235]), .Z(n20420) );
  AND U26799 ( .A(n20421), .B(n20422), .Z(n20419) );
  NAND U26800 ( .A(ereg[234]), .B(n19486), .Z(n20422) );
  NANDN U26801 ( .A(n19481), .B(ereg[235]), .Z(n20421) );
  NAND U26802 ( .A(n20423), .B(n20424), .Z(n15141) );
  NANDN U26803 ( .A(init), .B(e[236]), .Z(n20424) );
  AND U26804 ( .A(n20425), .B(n20426), .Z(n20423) );
  NAND U26805 ( .A(ereg[235]), .B(n19486), .Z(n20426) );
  NANDN U26806 ( .A(n19481), .B(ereg[236]), .Z(n20425) );
  NAND U26807 ( .A(n20427), .B(n20428), .Z(n15140) );
  NANDN U26808 ( .A(init), .B(e[237]), .Z(n20428) );
  AND U26809 ( .A(n20429), .B(n20430), .Z(n20427) );
  NAND U26810 ( .A(ereg[236]), .B(n19486), .Z(n20430) );
  NANDN U26811 ( .A(n19481), .B(ereg[237]), .Z(n20429) );
  NAND U26812 ( .A(n20431), .B(n20432), .Z(n15139) );
  NANDN U26813 ( .A(init), .B(e[238]), .Z(n20432) );
  AND U26814 ( .A(n20433), .B(n20434), .Z(n20431) );
  NAND U26815 ( .A(ereg[237]), .B(n19486), .Z(n20434) );
  NANDN U26816 ( .A(n19481), .B(ereg[238]), .Z(n20433) );
  NAND U26817 ( .A(n20435), .B(n20436), .Z(n15138) );
  NANDN U26818 ( .A(init), .B(e[239]), .Z(n20436) );
  AND U26819 ( .A(n20437), .B(n20438), .Z(n20435) );
  NAND U26820 ( .A(ereg[238]), .B(n19486), .Z(n20438) );
  NANDN U26821 ( .A(n19481), .B(ereg[239]), .Z(n20437) );
  NAND U26822 ( .A(n20439), .B(n20440), .Z(n15137) );
  NANDN U26823 ( .A(init), .B(e[240]), .Z(n20440) );
  AND U26824 ( .A(n20441), .B(n20442), .Z(n20439) );
  NAND U26825 ( .A(ereg[239]), .B(n19486), .Z(n20442) );
  NANDN U26826 ( .A(n19481), .B(ereg[240]), .Z(n20441) );
  NAND U26827 ( .A(n20443), .B(n20444), .Z(n15136) );
  NANDN U26828 ( .A(init), .B(e[241]), .Z(n20444) );
  AND U26829 ( .A(n20445), .B(n20446), .Z(n20443) );
  NAND U26830 ( .A(ereg[240]), .B(n19486), .Z(n20446) );
  NANDN U26831 ( .A(n19481), .B(ereg[241]), .Z(n20445) );
  NAND U26832 ( .A(n20447), .B(n20448), .Z(n15135) );
  NANDN U26833 ( .A(init), .B(e[242]), .Z(n20448) );
  AND U26834 ( .A(n20449), .B(n20450), .Z(n20447) );
  NAND U26835 ( .A(ereg[241]), .B(n19486), .Z(n20450) );
  NANDN U26836 ( .A(n19481), .B(ereg[242]), .Z(n20449) );
  NAND U26837 ( .A(n20451), .B(n20452), .Z(n15134) );
  NANDN U26838 ( .A(init), .B(e[243]), .Z(n20452) );
  AND U26839 ( .A(n20453), .B(n20454), .Z(n20451) );
  NAND U26840 ( .A(ereg[242]), .B(n19486), .Z(n20454) );
  NANDN U26841 ( .A(n19481), .B(ereg[243]), .Z(n20453) );
  NAND U26842 ( .A(n20455), .B(n20456), .Z(n15133) );
  NANDN U26843 ( .A(init), .B(e[244]), .Z(n20456) );
  AND U26844 ( .A(n20457), .B(n20458), .Z(n20455) );
  NAND U26845 ( .A(ereg[243]), .B(n19486), .Z(n20458) );
  NANDN U26846 ( .A(n19481), .B(ereg[244]), .Z(n20457) );
  NAND U26847 ( .A(n20459), .B(n20460), .Z(n15132) );
  NANDN U26848 ( .A(init), .B(e[245]), .Z(n20460) );
  AND U26849 ( .A(n20461), .B(n20462), .Z(n20459) );
  NAND U26850 ( .A(ereg[244]), .B(n19486), .Z(n20462) );
  NANDN U26851 ( .A(n19481), .B(ereg[245]), .Z(n20461) );
  NAND U26852 ( .A(n20463), .B(n20464), .Z(n15131) );
  NANDN U26853 ( .A(init), .B(e[246]), .Z(n20464) );
  AND U26854 ( .A(n20465), .B(n20466), .Z(n20463) );
  NAND U26855 ( .A(ereg[245]), .B(n19486), .Z(n20466) );
  NANDN U26856 ( .A(n19481), .B(ereg[246]), .Z(n20465) );
  NAND U26857 ( .A(n20467), .B(n20468), .Z(n15130) );
  NANDN U26858 ( .A(init), .B(e[247]), .Z(n20468) );
  AND U26859 ( .A(n20469), .B(n20470), .Z(n20467) );
  NAND U26860 ( .A(ereg[246]), .B(n19486), .Z(n20470) );
  NANDN U26861 ( .A(n19481), .B(ereg[247]), .Z(n20469) );
  NAND U26862 ( .A(n20471), .B(n20472), .Z(n15129) );
  NANDN U26863 ( .A(init), .B(e[248]), .Z(n20472) );
  AND U26864 ( .A(n20473), .B(n20474), .Z(n20471) );
  NAND U26865 ( .A(ereg[247]), .B(n19486), .Z(n20474) );
  NANDN U26866 ( .A(n19481), .B(ereg[248]), .Z(n20473) );
  NAND U26867 ( .A(n20475), .B(n20476), .Z(n15128) );
  NANDN U26868 ( .A(init), .B(e[249]), .Z(n20476) );
  AND U26869 ( .A(n20477), .B(n20478), .Z(n20475) );
  NAND U26870 ( .A(ereg[248]), .B(n19486), .Z(n20478) );
  NANDN U26871 ( .A(n19481), .B(ereg[249]), .Z(n20477) );
  NAND U26872 ( .A(n20479), .B(n20480), .Z(n15127) );
  NANDN U26873 ( .A(init), .B(e[250]), .Z(n20480) );
  AND U26874 ( .A(n20481), .B(n20482), .Z(n20479) );
  NAND U26875 ( .A(ereg[249]), .B(n19486), .Z(n20482) );
  NANDN U26876 ( .A(n19481), .B(ereg[250]), .Z(n20481) );
  NAND U26877 ( .A(n20483), .B(n20484), .Z(n15126) );
  NANDN U26878 ( .A(init), .B(e[251]), .Z(n20484) );
  AND U26879 ( .A(n20485), .B(n20486), .Z(n20483) );
  NAND U26880 ( .A(ereg[250]), .B(n19486), .Z(n20486) );
  NANDN U26881 ( .A(n19481), .B(ereg[251]), .Z(n20485) );
  NAND U26882 ( .A(n20487), .B(n20488), .Z(n15125) );
  NANDN U26883 ( .A(init), .B(e[252]), .Z(n20488) );
  AND U26884 ( .A(n20489), .B(n20490), .Z(n20487) );
  NAND U26885 ( .A(ereg[251]), .B(n19486), .Z(n20490) );
  NANDN U26886 ( .A(n19481), .B(ereg[252]), .Z(n20489) );
  NAND U26887 ( .A(n20491), .B(n20492), .Z(n15124) );
  NANDN U26888 ( .A(init), .B(e[253]), .Z(n20492) );
  AND U26889 ( .A(n20493), .B(n20494), .Z(n20491) );
  NAND U26890 ( .A(ereg[252]), .B(n19486), .Z(n20494) );
  NANDN U26891 ( .A(n19481), .B(ereg[253]), .Z(n20493) );
  NAND U26892 ( .A(n20495), .B(n20496), .Z(n15123) );
  NANDN U26893 ( .A(init), .B(e[254]), .Z(n20496) );
  AND U26894 ( .A(n20497), .B(n20498), .Z(n20495) );
  NAND U26895 ( .A(ereg[253]), .B(n19486), .Z(n20498) );
  NANDN U26896 ( .A(n19481), .B(ereg[254]), .Z(n20497) );
  NAND U26897 ( .A(n20499), .B(n20500), .Z(n15122) );
  NANDN U26898 ( .A(init), .B(e[255]), .Z(n20500) );
  AND U26899 ( .A(n20501), .B(n20502), .Z(n20499) );
  NAND U26900 ( .A(ereg[254]), .B(n19486), .Z(n20502) );
  NANDN U26901 ( .A(n19481), .B(ereg[255]), .Z(n20501) );
  NAND U26902 ( .A(n20503), .B(n20504), .Z(n15121) );
  NANDN U26903 ( .A(init), .B(e[256]), .Z(n20504) );
  AND U26904 ( .A(n20505), .B(n20506), .Z(n20503) );
  NAND U26905 ( .A(ereg[255]), .B(n19486), .Z(n20506) );
  NANDN U26906 ( .A(n19481), .B(ereg[256]), .Z(n20505) );
  NAND U26907 ( .A(n20507), .B(n20508), .Z(n15120) );
  NANDN U26908 ( .A(init), .B(e[257]), .Z(n20508) );
  AND U26909 ( .A(n20509), .B(n20510), .Z(n20507) );
  NAND U26910 ( .A(ereg[256]), .B(n19486), .Z(n20510) );
  NANDN U26911 ( .A(n19481), .B(ereg[257]), .Z(n20509) );
  NAND U26912 ( .A(n20511), .B(n20512), .Z(n15119) );
  NANDN U26913 ( .A(init), .B(e[258]), .Z(n20512) );
  AND U26914 ( .A(n20513), .B(n20514), .Z(n20511) );
  NAND U26915 ( .A(ereg[257]), .B(n19486), .Z(n20514) );
  NANDN U26916 ( .A(n19481), .B(ereg[258]), .Z(n20513) );
  NAND U26917 ( .A(n20515), .B(n20516), .Z(n15118) );
  NANDN U26918 ( .A(init), .B(e[259]), .Z(n20516) );
  AND U26919 ( .A(n20517), .B(n20518), .Z(n20515) );
  NAND U26920 ( .A(ereg[258]), .B(n19486), .Z(n20518) );
  NANDN U26921 ( .A(n19481), .B(ereg[259]), .Z(n20517) );
  NAND U26922 ( .A(n20519), .B(n20520), .Z(n15117) );
  NANDN U26923 ( .A(init), .B(e[260]), .Z(n20520) );
  AND U26924 ( .A(n20521), .B(n20522), .Z(n20519) );
  NAND U26925 ( .A(ereg[259]), .B(n19486), .Z(n20522) );
  NANDN U26926 ( .A(n19481), .B(ereg[260]), .Z(n20521) );
  NAND U26927 ( .A(n20523), .B(n20524), .Z(n15116) );
  NANDN U26928 ( .A(init), .B(e[261]), .Z(n20524) );
  AND U26929 ( .A(n20525), .B(n20526), .Z(n20523) );
  NAND U26930 ( .A(ereg[260]), .B(n19486), .Z(n20526) );
  NANDN U26931 ( .A(n19481), .B(ereg[261]), .Z(n20525) );
  NAND U26932 ( .A(n20527), .B(n20528), .Z(n15115) );
  NANDN U26933 ( .A(init), .B(e[262]), .Z(n20528) );
  AND U26934 ( .A(n20529), .B(n20530), .Z(n20527) );
  NAND U26935 ( .A(ereg[261]), .B(n19486), .Z(n20530) );
  NANDN U26936 ( .A(n19481), .B(ereg[262]), .Z(n20529) );
  NAND U26937 ( .A(n20531), .B(n20532), .Z(n15114) );
  NANDN U26938 ( .A(init), .B(e[263]), .Z(n20532) );
  AND U26939 ( .A(n20533), .B(n20534), .Z(n20531) );
  NAND U26940 ( .A(ereg[262]), .B(n19486), .Z(n20534) );
  NANDN U26941 ( .A(n19481), .B(ereg[263]), .Z(n20533) );
  NAND U26942 ( .A(n20535), .B(n20536), .Z(n15113) );
  NANDN U26943 ( .A(init), .B(e[264]), .Z(n20536) );
  AND U26944 ( .A(n20537), .B(n20538), .Z(n20535) );
  NAND U26945 ( .A(ereg[263]), .B(n19486), .Z(n20538) );
  NANDN U26946 ( .A(n19481), .B(ereg[264]), .Z(n20537) );
  NAND U26947 ( .A(n20539), .B(n20540), .Z(n15112) );
  NANDN U26948 ( .A(init), .B(e[265]), .Z(n20540) );
  AND U26949 ( .A(n20541), .B(n20542), .Z(n20539) );
  NAND U26950 ( .A(ereg[264]), .B(n19486), .Z(n20542) );
  NANDN U26951 ( .A(n19481), .B(ereg[265]), .Z(n20541) );
  NAND U26952 ( .A(n20543), .B(n20544), .Z(n15111) );
  NANDN U26953 ( .A(init), .B(e[266]), .Z(n20544) );
  AND U26954 ( .A(n20545), .B(n20546), .Z(n20543) );
  NAND U26955 ( .A(ereg[265]), .B(n19486), .Z(n20546) );
  NANDN U26956 ( .A(n19481), .B(ereg[266]), .Z(n20545) );
  NAND U26957 ( .A(n20547), .B(n20548), .Z(n15110) );
  NANDN U26958 ( .A(init), .B(e[267]), .Z(n20548) );
  AND U26959 ( .A(n20549), .B(n20550), .Z(n20547) );
  NAND U26960 ( .A(ereg[266]), .B(n19486), .Z(n20550) );
  NANDN U26961 ( .A(n19481), .B(ereg[267]), .Z(n20549) );
  NAND U26962 ( .A(n20551), .B(n20552), .Z(n15109) );
  NANDN U26963 ( .A(init), .B(e[268]), .Z(n20552) );
  AND U26964 ( .A(n20553), .B(n20554), .Z(n20551) );
  NAND U26965 ( .A(ereg[267]), .B(n19486), .Z(n20554) );
  NANDN U26966 ( .A(n19481), .B(ereg[268]), .Z(n20553) );
  NAND U26967 ( .A(n20555), .B(n20556), .Z(n15108) );
  NANDN U26968 ( .A(init), .B(e[269]), .Z(n20556) );
  AND U26969 ( .A(n20557), .B(n20558), .Z(n20555) );
  NAND U26970 ( .A(ereg[268]), .B(n19486), .Z(n20558) );
  NANDN U26971 ( .A(n19481), .B(ereg[269]), .Z(n20557) );
  NAND U26972 ( .A(n20559), .B(n20560), .Z(n15107) );
  NANDN U26973 ( .A(init), .B(e[270]), .Z(n20560) );
  AND U26974 ( .A(n20561), .B(n20562), .Z(n20559) );
  NAND U26975 ( .A(ereg[269]), .B(n19486), .Z(n20562) );
  NANDN U26976 ( .A(n19481), .B(ereg[270]), .Z(n20561) );
  NAND U26977 ( .A(n20563), .B(n20564), .Z(n15106) );
  NANDN U26978 ( .A(init), .B(e[271]), .Z(n20564) );
  AND U26979 ( .A(n20565), .B(n20566), .Z(n20563) );
  NAND U26980 ( .A(ereg[270]), .B(n19486), .Z(n20566) );
  NANDN U26981 ( .A(n19481), .B(ereg[271]), .Z(n20565) );
  NAND U26982 ( .A(n20567), .B(n20568), .Z(n15105) );
  NANDN U26983 ( .A(init), .B(e[272]), .Z(n20568) );
  AND U26984 ( .A(n20569), .B(n20570), .Z(n20567) );
  NAND U26985 ( .A(ereg[271]), .B(n19486), .Z(n20570) );
  NANDN U26986 ( .A(n19481), .B(ereg[272]), .Z(n20569) );
  NAND U26987 ( .A(n20571), .B(n20572), .Z(n15104) );
  NANDN U26988 ( .A(init), .B(e[273]), .Z(n20572) );
  AND U26989 ( .A(n20573), .B(n20574), .Z(n20571) );
  NAND U26990 ( .A(ereg[272]), .B(n19486), .Z(n20574) );
  NANDN U26991 ( .A(n19481), .B(ereg[273]), .Z(n20573) );
  NAND U26992 ( .A(n20575), .B(n20576), .Z(n15103) );
  NANDN U26993 ( .A(init), .B(e[274]), .Z(n20576) );
  AND U26994 ( .A(n20577), .B(n20578), .Z(n20575) );
  NAND U26995 ( .A(ereg[273]), .B(n19486), .Z(n20578) );
  NANDN U26996 ( .A(n19481), .B(ereg[274]), .Z(n20577) );
  NAND U26997 ( .A(n20579), .B(n20580), .Z(n15102) );
  NANDN U26998 ( .A(init), .B(e[275]), .Z(n20580) );
  AND U26999 ( .A(n20581), .B(n20582), .Z(n20579) );
  NAND U27000 ( .A(ereg[274]), .B(n19486), .Z(n20582) );
  NANDN U27001 ( .A(n19481), .B(ereg[275]), .Z(n20581) );
  NAND U27002 ( .A(n20583), .B(n20584), .Z(n15101) );
  NANDN U27003 ( .A(init), .B(e[276]), .Z(n20584) );
  AND U27004 ( .A(n20585), .B(n20586), .Z(n20583) );
  NAND U27005 ( .A(ereg[275]), .B(n19486), .Z(n20586) );
  NANDN U27006 ( .A(n19481), .B(ereg[276]), .Z(n20585) );
  NAND U27007 ( .A(n20587), .B(n20588), .Z(n15100) );
  NANDN U27008 ( .A(init), .B(e[277]), .Z(n20588) );
  AND U27009 ( .A(n20589), .B(n20590), .Z(n20587) );
  NAND U27010 ( .A(ereg[276]), .B(n19486), .Z(n20590) );
  NANDN U27011 ( .A(n19481), .B(ereg[277]), .Z(n20589) );
  NAND U27012 ( .A(n20591), .B(n20592), .Z(n15099) );
  NANDN U27013 ( .A(init), .B(e[278]), .Z(n20592) );
  AND U27014 ( .A(n20593), .B(n20594), .Z(n20591) );
  NAND U27015 ( .A(ereg[277]), .B(n19486), .Z(n20594) );
  NANDN U27016 ( .A(n19481), .B(ereg[278]), .Z(n20593) );
  NAND U27017 ( .A(n20595), .B(n20596), .Z(n15098) );
  NANDN U27018 ( .A(init), .B(e[279]), .Z(n20596) );
  AND U27019 ( .A(n20597), .B(n20598), .Z(n20595) );
  NAND U27020 ( .A(ereg[278]), .B(n19486), .Z(n20598) );
  NANDN U27021 ( .A(n19481), .B(ereg[279]), .Z(n20597) );
  NAND U27022 ( .A(n20599), .B(n20600), .Z(n15097) );
  NANDN U27023 ( .A(init), .B(e[280]), .Z(n20600) );
  AND U27024 ( .A(n20601), .B(n20602), .Z(n20599) );
  NAND U27025 ( .A(ereg[279]), .B(n19486), .Z(n20602) );
  NANDN U27026 ( .A(n19481), .B(ereg[280]), .Z(n20601) );
  NAND U27027 ( .A(n20603), .B(n20604), .Z(n15096) );
  NANDN U27028 ( .A(init), .B(e[281]), .Z(n20604) );
  AND U27029 ( .A(n20605), .B(n20606), .Z(n20603) );
  NAND U27030 ( .A(ereg[280]), .B(n19486), .Z(n20606) );
  NANDN U27031 ( .A(n19481), .B(ereg[281]), .Z(n20605) );
  NAND U27032 ( .A(n20607), .B(n20608), .Z(n15095) );
  NANDN U27033 ( .A(init), .B(e[282]), .Z(n20608) );
  AND U27034 ( .A(n20609), .B(n20610), .Z(n20607) );
  NAND U27035 ( .A(ereg[281]), .B(n19486), .Z(n20610) );
  NANDN U27036 ( .A(n19481), .B(ereg[282]), .Z(n20609) );
  NAND U27037 ( .A(n20611), .B(n20612), .Z(n15094) );
  NANDN U27038 ( .A(init), .B(e[283]), .Z(n20612) );
  AND U27039 ( .A(n20613), .B(n20614), .Z(n20611) );
  NAND U27040 ( .A(ereg[282]), .B(n19486), .Z(n20614) );
  NANDN U27041 ( .A(n19481), .B(ereg[283]), .Z(n20613) );
  NAND U27042 ( .A(n20615), .B(n20616), .Z(n15093) );
  NANDN U27043 ( .A(init), .B(e[284]), .Z(n20616) );
  AND U27044 ( .A(n20617), .B(n20618), .Z(n20615) );
  NAND U27045 ( .A(ereg[283]), .B(n19486), .Z(n20618) );
  NANDN U27046 ( .A(n19481), .B(ereg[284]), .Z(n20617) );
  NAND U27047 ( .A(n20619), .B(n20620), .Z(n15092) );
  NANDN U27048 ( .A(init), .B(e[285]), .Z(n20620) );
  AND U27049 ( .A(n20621), .B(n20622), .Z(n20619) );
  NAND U27050 ( .A(ereg[284]), .B(n19486), .Z(n20622) );
  NANDN U27051 ( .A(n19481), .B(ereg[285]), .Z(n20621) );
  NAND U27052 ( .A(n20623), .B(n20624), .Z(n15091) );
  NANDN U27053 ( .A(init), .B(e[286]), .Z(n20624) );
  AND U27054 ( .A(n20625), .B(n20626), .Z(n20623) );
  NAND U27055 ( .A(ereg[285]), .B(n19486), .Z(n20626) );
  NANDN U27056 ( .A(n19481), .B(ereg[286]), .Z(n20625) );
  NAND U27057 ( .A(n20627), .B(n20628), .Z(n15090) );
  NANDN U27058 ( .A(init), .B(e[287]), .Z(n20628) );
  AND U27059 ( .A(n20629), .B(n20630), .Z(n20627) );
  NAND U27060 ( .A(ereg[286]), .B(n19486), .Z(n20630) );
  NANDN U27061 ( .A(n19481), .B(ereg[287]), .Z(n20629) );
  NAND U27062 ( .A(n20631), .B(n20632), .Z(n15089) );
  NANDN U27063 ( .A(init), .B(e[288]), .Z(n20632) );
  AND U27064 ( .A(n20633), .B(n20634), .Z(n20631) );
  NAND U27065 ( .A(ereg[287]), .B(n19486), .Z(n20634) );
  NANDN U27066 ( .A(n19481), .B(ereg[288]), .Z(n20633) );
  NAND U27067 ( .A(n20635), .B(n20636), .Z(n15088) );
  NANDN U27068 ( .A(init), .B(e[289]), .Z(n20636) );
  AND U27069 ( .A(n20637), .B(n20638), .Z(n20635) );
  NAND U27070 ( .A(ereg[288]), .B(n19486), .Z(n20638) );
  NANDN U27071 ( .A(n19481), .B(ereg[289]), .Z(n20637) );
  NAND U27072 ( .A(n20639), .B(n20640), .Z(n15087) );
  NANDN U27073 ( .A(init), .B(e[290]), .Z(n20640) );
  AND U27074 ( .A(n20641), .B(n20642), .Z(n20639) );
  NAND U27075 ( .A(ereg[289]), .B(n19486), .Z(n20642) );
  NANDN U27076 ( .A(n19481), .B(ereg[290]), .Z(n20641) );
  NAND U27077 ( .A(n20643), .B(n20644), .Z(n15086) );
  NANDN U27078 ( .A(init), .B(e[291]), .Z(n20644) );
  AND U27079 ( .A(n20645), .B(n20646), .Z(n20643) );
  NAND U27080 ( .A(ereg[290]), .B(n19486), .Z(n20646) );
  NANDN U27081 ( .A(n19481), .B(ereg[291]), .Z(n20645) );
  NAND U27082 ( .A(n20647), .B(n20648), .Z(n15085) );
  NANDN U27083 ( .A(init), .B(e[292]), .Z(n20648) );
  AND U27084 ( .A(n20649), .B(n20650), .Z(n20647) );
  NAND U27085 ( .A(ereg[291]), .B(n19486), .Z(n20650) );
  NANDN U27086 ( .A(n19481), .B(ereg[292]), .Z(n20649) );
  NAND U27087 ( .A(n20651), .B(n20652), .Z(n15084) );
  NANDN U27088 ( .A(init), .B(e[293]), .Z(n20652) );
  AND U27089 ( .A(n20653), .B(n20654), .Z(n20651) );
  NAND U27090 ( .A(ereg[292]), .B(n19486), .Z(n20654) );
  NANDN U27091 ( .A(n19481), .B(ereg[293]), .Z(n20653) );
  NAND U27092 ( .A(n20655), .B(n20656), .Z(n15083) );
  NANDN U27093 ( .A(init), .B(e[294]), .Z(n20656) );
  AND U27094 ( .A(n20657), .B(n20658), .Z(n20655) );
  NAND U27095 ( .A(ereg[293]), .B(n19486), .Z(n20658) );
  NANDN U27096 ( .A(n19481), .B(ereg[294]), .Z(n20657) );
  NAND U27097 ( .A(n20659), .B(n20660), .Z(n15082) );
  NANDN U27098 ( .A(init), .B(e[295]), .Z(n20660) );
  AND U27099 ( .A(n20661), .B(n20662), .Z(n20659) );
  NAND U27100 ( .A(ereg[294]), .B(n19486), .Z(n20662) );
  NANDN U27101 ( .A(n19481), .B(ereg[295]), .Z(n20661) );
  NAND U27102 ( .A(n20663), .B(n20664), .Z(n15081) );
  NANDN U27103 ( .A(init), .B(e[296]), .Z(n20664) );
  AND U27104 ( .A(n20665), .B(n20666), .Z(n20663) );
  NAND U27105 ( .A(ereg[295]), .B(n19486), .Z(n20666) );
  NANDN U27106 ( .A(n19481), .B(ereg[296]), .Z(n20665) );
  NAND U27107 ( .A(n20667), .B(n20668), .Z(n15080) );
  NANDN U27108 ( .A(init), .B(e[297]), .Z(n20668) );
  AND U27109 ( .A(n20669), .B(n20670), .Z(n20667) );
  NAND U27110 ( .A(ereg[296]), .B(n19486), .Z(n20670) );
  NANDN U27111 ( .A(n19481), .B(ereg[297]), .Z(n20669) );
  NAND U27112 ( .A(n20671), .B(n20672), .Z(n15079) );
  NANDN U27113 ( .A(init), .B(e[298]), .Z(n20672) );
  AND U27114 ( .A(n20673), .B(n20674), .Z(n20671) );
  NAND U27115 ( .A(ereg[297]), .B(n19486), .Z(n20674) );
  NANDN U27116 ( .A(n19481), .B(ereg[298]), .Z(n20673) );
  NAND U27117 ( .A(n20675), .B(n20676), .Z(n15078) );
  NANDN U27118 ( .A(init), .B(e[299]), .Z(n20676) );
  AND U27119 ( .A(n20677), .B(n20678), .Z(n20675) );
  NAND U27120 ( .A(ereg[298]), .B(n19486), .Z(n20678) );
  NANDN U27121 ( .A(n19481), .B(ereg[299]), .Z(n20677) );
  NAND U27122 ( .A(n20679), .B(n20680), .Z(n15077) );
  NANDN U27123 ( .A(init), .B(e[300]), .Z(n20680) );
  AND U27124 ( .A(n20681), .B(n20682), .Z(n20679) );
  NAND U27125 ( .A(ereg[299]), .B(n19486), .Z(n20682) );
  NANDN U27126 ( .A(n19481), .B(ereg[300]), .Z(n20681) );
  NAND U27127 ( .A(n20683), .B(n20684), .Z(n15076) );
  NANDN U27128 ( .A(init), .B(e[301]), .Z(n20684) );
  AND U27129 ( .A(n20685), .B(n20686), .Z(n20683) );
  NAND U27130 ( .A(ereg[300]), .B(n19486), .Z(n20686) );
  NANDN U27131 ( .A(n19481), .B(ereg[301]), .Z(n20685) );
  NAND U27132 ( .A(n20687), .B(n20688), .Z(n15075) );
  NANDN U27133 ( .A(init), .B(e[302]), .Z(n20688) );
  AND U27134 ( .A(n20689), .B(n20690), .Z(n20687) );
  NAND U27135 ( .A(ereg[301]), .B(n19486), .Z(n20690) );
  NANDN U27136 ( .A(n19481), .B(ereg[302]), .Z(n20689) );
  NAND U27137 ( .A(n20691), .B(n20692), .Z(n15074) );
  NANDN U27138 ( .A(init), .B(e[303]), .Z(n20692) );
  AND U27139 ( .A(n20693), .B(n20694), .Z(n20691) );
  NAND U27140 ( .A(ereg[302]), .B(n19486), .Z(n20694) );
  NANDN U27141 ( .A(n19481), .B(ereg[303]), .Z(n20693) );
  NAND U27142 ( .A(n20695), .B(n20696), .Z(n15073) );
  NANDN U27143 ( .A(init), .B(e[304]), .Z(n20696) );
  AND U27144 ( .A(n20697), .B(n20698), .Z(n20695) );
  NAND U27145 ( .A(ereg[303]), .B(n19486), .Z(n20698) );
  NANDN U27146 ( .A(n19481), .B(ereg[304]), .Z(n20697) );
  NAND U27147 ( .A(n20699), .B(n20700), .Z(n15072) );
  NANDN U27148 ( .A(init), .B(e[305]), .Z(n20700) );
  AND U27149 ( .A(n20701), .B(n20702), .Z(n20699) );
  NAND U27150 ( .A(ereg[304]), .B(n19486), .Z(n20702) );
  NANDN U27151 ( .A(n19481), .B(ereg[305]), .Z(n20701) );
  NAND U27152 ( .A(n20703), .B(n20704), .Z(n15071) );
  NANDN U27153 ( .A(init), .B(e[306]), .Z(n20704) );
  AND U27154 ( .A(n20705), .B(n20706), .Z(n20703) );
  NAND U27155 ( .A(ereg[305]), .B(n19486), .Z(n20706) );
  NANDN U27156 ( .A(n19481), .B(ereg[306]), .Z(n20705) );
  NAND U27157 ( .A(n20707), .B(n20708), .Z(n15070) );
  NANDN U27158 ( .A(init), .B(e[307]), .Z(n20708) );
  AND U27159 ( .A(n20709), .B(n20710), .Z(n20707) );
  NAND U27160 ( .A(ereg[306]), .B(n19486), .Z(n20710) );
  NANDN U27161 ( .A(n19481), .B(ereg[307]), .Z(n20709) );
  NAND U27162 ( .A(n20711), .B(n20712), .Z(n15069) );
  NANDN U27163 ( .A(init), .B(e[308]), .Z(n20712) );
  AND U27164 ( .A(n20713), .B(n20714), .Z(n20711) );
  NAND U27165 ( .A(ereg[307]), .B(n19486), .Z(n20714) );
  NANDN U27166 ( .A(n19481), .B(ereg[308]), .Z(n20713) );
  NAND U27167 ( .A(n20715), .B(n20716), .Z(n15068) );
  NANDN U27168 ( .A(init), .B(e[309]), .Z(n20716) );
  AND U27169 ( .A(n20717), .B(n20718), .Z(n20715) );
  NAND U27170 ( .A(ereg[308]), .B(n19486), .Z(n20718) );
  NANDN U27171 ( .A(n19481), .B(ereg[309]), .Z(n20717) );
  NAND U27172 ( .A(n20719), .B(n20720), .Z(n15067) );
  NANDN U27173 ( .A(init), .B(e[310]), .Z(n20720) );
  AND U27174 ( .A(n20721), .B(n20722), .Z(n20719) );
  NAND U27175 ( .A(ereg[309]), .B(n19486), .Z(n20722) );
  NANDN U27176 ( .A(n19481), .B(ereg[310]), .Z(n20721) );
  NAND U27177 ( .A(n20723), .B(n20724), .Z(n15066) );
  NANDN U27178 ( .A(init), .B(e[311]), .Z(n20724) );
  AND U27179 ( .A(n20725), .B(n20726), .Z(n20723) );
  NAND U27180 ( .A(ereg[310]), .B(n19486), .Z(n20726) );
  NANDN U27181 ( .A(n19481), .B(ereg[311]), .Z(n20725) );
  NAND U27182 ( .A(n20727), .B(n20728), .Z(n15065) );
  NANDN U27183 ( .A(init), .B(e[312]), .Z(n20728) );
  AND U27184 ( .A(n20729), .B(n20730), .Z(n20727) );
  NAND U27185 ( .A(ereg[311]), .B(n19486), .Z(n20730) );
  NANDN U27186 ( .A(n19481), .B(ereg[312]), .Z(n20729) );
  NAND U27187 ( .A(n20731), .B(n20732), .Z(n15064) );
  NANDN U27188 ( .A(init), .B(e[313]), .Z(n20732) );
  AND U27189 ( .A(n20733), .B(n20734), .Z(n20731) );
  NAND U27190 ( .A(ereg[312]), .B(n19486), .Z(n20734) );
  NANDN U27191 ( .A(n19481), .B(ereg[313]), .Z(n20733) );
  NAND U27192 ( .A(n20735), .B(n20736), .Z(n15063) );
  NANDN U27193 ( .A(init), .B(e[314]), .Z(n20736) );
  AND U27194 ( .A(n20737), .B(n20738), .Z(n20735) );
  NAND U27195 ( .A(ereg[313]), .B(n19486), .Z(n20738) );
  NANDN U27196 ( .A(n19481), .B(ereg[314]), .Z(n20737) );
  NAND U27197 ( .A(n20739), .B(n20740), .Z(n15062) );
  NANDN U27198 ( .A(init), .B(e[315]), .Z(n20740) );
  AND U27199 ( .A(n20741), .B(n20742), .Z(n20739) );
  NAND U27200 ( .A(ereg[314]), .B(n19486), .Z(n20742) );
  NANDN U27201 ( .A(n19481), .B(ereg[315]), .Z(n20741) );
  NAND U27202 ( .A(n20743), .B(n20744), .Z(n15061) );
  NANDN U27203 ( .A(init), .B(e[316]), .Z(n20744) );
  AND U27204 ( .A(n20745), .B(n20746), .Z(n20743) );
  NAND U27205 ( .A(ereg[315]), .B(n19486), .Z(n20746) );
  NANDN U27206 ( .A(n19481), .B(ereg[316]), .Z(n20745) );
  NAND U27207 ( .A(n20747), .B(n20748), .Z(n15060) );
  NANDN U27208 ( .A(init), .B(e[317]), .Z(n20748) );
  AND U27209 ( .A(n20749), .B(n20750), .Z(n20747) );
  NAND U27210 ( .A(ereg[316]), .B(n19486), .Z(n20750) );
  NANDN U27211 ( .A(n19481), .B(ereg[317]), .Z(n20749) );
  NAND U27212 ( .A(n20751), .B(n20752), .Z(n15059) );
  NANDN U27213 ( .A(init), .B(e[318]), .Z(n20752) );
  AND U27214 ( .A(n20753), .B(n20754), .Z(n20751) );
  NAND U27215 ( .A(ereg[317]), .B(n19486), .Z(n20754) );
  NANDN U27216 ( .A(n19481), .B(ereg[318]), .Z(n20753) );
  NAND U27217 ( .A(n20755), .B(n20756), .Z(n15058) );
  NANDN U27218 ( .A(init), .B(e[319]), .Z(n20756) );
  AND U27219 ( .A(n20757), .B(n20758), .Z(n20755) );
  NAND U27220 ( .A(ereg[318]), .B(n19486), .Z(n20758) );
  NANDN U27221 ( .A(n19481), .B(ereg[319]), .Z(n20757) );
  NAND U27222 ( .A(n20759), .B(n20760), .Z(n15057) );
  NANDN U27223 ( .A(init), .B(e[320]), .Z(n20760) );
  AND U27224 ( .A(n20761), .B(n20762), .Z(n20759) );
  NAND U27225 ( .A(ereg[319]), .B(n19486), .Z(n20762) );
  NANDN U27226 ( .A(n19481), .B(ereg[320]), .Z(n20761) );
  NAND U27227 ( .A(n20763), .B(n20764), .Z(n15056) );
  NANDN U27228 ( .A(init), .B(e[321]), .Z(n20764) );
  AND U27229 ( .A(n20765), .B(n20766), .Z(n20763) );
  NAND U27230 ( .A(ereg[320]), .B(n19486), .Z(n20766) );
  NANDN U27231 ( .A(n19481), .B(ereg[321]), .Z(n20765) );
  NAND U27232 ( .A(n20767), .B(n20768), .Z(n15055) );
  NANDN U27233 ( .A(init), .B(e[322]), .Z(n20768) );
  AND U27234 ( .A(n20769), .B(n20770), .Z(n20767) );
  NAND U27235 ( .A(ereg[321]), .B(n19486), .Z(n20770) );
  NANDN U27236 ( .A(n19481), .B(ereg[322]), .Z(n20769) );
  NAND U27237 ( .A(n20771), .B(n20772), .Z(n15054) );
  NANDN U27238 ( .A(init), .B(e[323]), .Z(n20772) );
  AND U27239 ( .A(n20773), .B(n20774), .Z(n20771) );
  NAND U27240 ( .A(ereg[322]), .B(n19486), .Z(n20774) );
  NANDN U27241 ( .A(n19481), .B(ereg[323]), .Z(n20773) );
  NAND U27242 ( .A(n20775), .B(n20776), .Z(n15053) );
  NANDN U27243 ( .A(init), .B(e[324]), .Z(n20776) );
  AND U27244 ( .A(n20777), .B(n20778), .Z(n20775) );
  NAND U27245 ( .A(ereg[323]), .B(n19486), .Z(n20778) );
  NANDN U27246 ( .A(n19481), .B(ereg[324]), .Z(n20777) );
  NAND U27247 ( .A(n20779), .B(n20780), .Z(n15052) );
  NANDN U27248 ( .A(init), .B(e[325]), .Z(n20780) );
  AND U27249 ( .A(n20781), .B(n20782), .Z(n20779) );
  NAND U27250 ( .A(ereg[324]), .B(n19486), .Z(n20782) );
  NANDN U27251 ( .A(n19481), .B(ereg[325]), .Z(n20781) );
  NAND U27252 ( .A(n20783), .B(n20784), .Z(n15051) );
  NANDN U27253 ( .A(init), .B(e[326]), .Z(n20784) );
  AND U27254 ( .A(n20785), .B(n20786), .Z(n20783) );
  NAND U27255 ( .A(ereg[325]), .B(n19486), .Z(n20786) );
  NANDN U27256 ( .A(n19481), .B(ereg[326]), .Z(n20785) );
  NAND U27257 ( .A(n20787), .B(n20788), .Z(n15050) );
  NANDN U27258 ( .A(init), .B(e[327]), .Z(n20788) );
  AND U27259 ( .A(n20789), .B(n20790), .Z(n20787) );
  NAND U27260 ( .A(ereg[326]), .B(n19486), .Z(n20790) );
  NANDN U27261 ( .A(n19481), .B(ereg[327]), .Z(n20789) );
  NAND U27262 ( .A(n20791), .B(n20792), .Z(n15049) );
  NANDN U27263 ( .A(init), .B(e[328]), .Z(n20792) );
  AND U27264 ( .A(n20793), .B(n20794), .Z(n20791) );
  NAND U27265 ( .A(ereg[327]), .B(n19486), .Z(n20794) );
  NANDN U27266 ( .A(n19481), .B(ereg[328]), .Z(n20793) );
  NAND U27267 ( .A(n20795), .B(n20796), .Z(n15048) );
  NANDN U27268 ( .A(init), .B(e[329]), .Z(n20796) );
  AND U27269 ( .A(n20797), .B(n20798), .Z(n20795) );
  NAND U27270 ( .A(ereg[328]), .B(n19486), .Z(n20798) );
  NANDN U27271 ( .A(n19481), .B(ereg[329]), .Z(n20797) );
  NAND U27272 ( .A(n20799), .B(n20800), .Z(n15047) );
  NANDN U27273 ( .A(init), .B(e[330]), .Z(n20800) );
  AND U27274 ( .A(n20801), .B(n20802), .Z(n20799) );
  NAND U27275 ( .A(ereg[329]), .B(n19486), .Z(n20802) );
  NANDN U27276 ( .A(n19481), .B(ereg[330]), .Z(n20801) );
  NAND U27277 ( .A(n20803), .B(n20804), .Z(n15046) );
  NANDN U27278 ( .A(init), .B(e[331]), .Z(n20804) );
  AND U27279 ( .A(n20805), .B(n20806), .Z(n20803) );
  NAND U27280 ( .A(ereg[330]), .B(n19486), .Z(n20806) );
  NANDN U27281 ( .A(n19481), .B(ereg[331]), .Z(n20805) );
  NAND U27282 ( .A(n20807), .B(n20808), .Z(n15045) );
  NANDN U27283 ( .A(init), .B(e[332]), .Z(n20808) );
  AND U27284 ( .A(n20809), .B(n20810), .Z(n20807) );
  NAND U27285 ( .A(ereg[331]), .B(n19486), .Z(n20810) );
  NANDN U27286 ( .A(n19481), .B(ereg[332]), .Z(n20809) );
  NAND U27287 ( .A(n20811), .B(n20812), .Z(n15044) );
  NANDN U27288 ( .A(init), .B(e[333]), .Z(n20812) );
  AND U27289 ( .A(n20813), .B(n20814), .Z(n20811) );
  NAND U27290 ( .A(ereg[332]), .B(n19486), .Z(n20814) );
  NANDN U27291 ( .A(n19481), .B(ereg[333]), .Z(n20813) );
  NAND U27292 ( .A(n20815), .B(n20816), .Z(n15043) );
  NANDN U27293 ( .A(init), .B(e[334]), .Z(n20816) );
  AND U27294 ( .A(n20817), .B(n20818), .Z(n20815) );
  NAND U27295 ( .A(ereg[333]), .B(n19486), .Z(n20818) );
  NANDN U27296 ( .A(n19481), .B(ereg[334]), .Z(n20817) );
  NAND U27297 ( .A(n20819), .B(n20820), .Z(n15042) );
  NANDN U27298 ( .A(init), .B(e[335]), .Z(n20820) );
  AND U27299 ( .A(n20821), .B(n20822), .Z(n20819) );
  NAND U27300 ( .A(ereg[334]), .B(n19486), .Z(n20822) );
  NANDN U27301 ( .A(n19481), .B(ereg[335]), .Z(n20821) );
  NAND U27302 ( .A(n20823), .B(n20824), .Z(n15041) );
  NANDN U27303 ( .A(init), .B(e[336]), .Z(n20824) );
  AND U27304 ( .A(n20825), .B(n20826), .Z(n20823) );
  NAND U27305 ( .A(ereg[335]), .B(n19486), .Z(n20826) );
  NANDN U27306 ( .A(n19481), .B(ereg[336]), .Z(n20825) );
  NAND U27307 ( .A(n20827), .B(n20828), .Z(n15040) );
  NANDN U27308 ( .A(init), .B(e[337]), .Z(n20828) );
  AND U27309 ( .A(n20829), .B(n20830), .Z(n20827) );
  NAND U27310 ( .A(ereg[336]), .B(n19486), .Z(n20830) );
  NANDN U27311 ( .A(n19481), .B(ereg[337]), .Z(n20829) );
  NAND U27312 ( .A(n20831), .B(n20832), .Z(n15039) );
  NANDN U27313 ( .A(init), .B(e[338]), .Z(n20832) );
  AND U27314 ( .A(n20833), .B(n20834), .Z(n20831) );
  NAND U27315 ( .A(ereg[337]), .B(n19486), .Z(n20834) );
  NANDN U27316 ( .A(n19481), .B(ereg[338]), .Z(n20833) );
  NAND U27317 ( .A(n20835), .B(n20836), .Z(n15038) );
  NANDN U27318 ( .A(init), .B(e[339]), .Z(n20836) );
  AND U27319 ( .A(n20837), .B(n20838), .Z(n20835) );
  NAND U27320 ( .A(ereg[338]), .B(n19486), .Z(n20838) );
  NANDN U27321 ( .A(n19481), .B(ereg[339]), .Z(n20837) );
  NAND U27322 ( .A(n20839), .B(n20840), .Z(n15037) );
  NANDN U27323 ( .A(init), .B(e[340]), .Z(n20840) );
  AND U27324 ( .A(n20841), .B(n20842), .Z(n20839) );
  NAND U27325 ( .A(ereg[339]), .B(n19486), .Z(n20842) );
  NANDN U27326 ( .A(n19481), .B(ereg[340]), .Z(n20841) );
  NAND U27327 ( .A(n20843), .B(n20844), .Z(n15036) );
  NANDN U27328 ( .A(init), .B(e[341]), .Z(n20844) );
  AND U27329 ( .A(n20845), .B(n20846), .Z(n20843) );
  NAND U27330 ( .A(ereg[340]), .B(n19486), .Z(n20846) );
  NANDN U27331 ( .A(n19481), .B(ereg[341]), .Z(n20845) );
  NAND U27332 ( .A(n20847), .B(n20848), .Z(n15035) );
  NANDN U27333 ( .A(init), .B(e[342]), .Z(n20848) );
  AND U27334 ( .A(n20849), .B(n20850), .Z(n20847) );
  NAND U27335 ( .A(ereg[341]), .B(n19486), .Z(n20850) );
  NANDN U27336 ( .A(n19481), .B(ereg[342]), .Z(n20849) );
  NAND U27337 ( .A(n20851), .B(n20852), .Z(n15034) );
  NANDN U27338 ( .A(init), .B(e[343]), .Z(n20852) );
  AND U27339 ( .A(n20853), .B(n20854), .Z(n20851) );
  NAND U27340 ( .A(ereg[342]), .B(n19486), .Z(n20854) );
  NANDN U27341 ( .A(n19481), .B(ereg[343]), .Z(n20853) );
  NAND U27342 ( .A(n20855), .B(n20856), .Z(n15033) );
  NANDN U27343 ( .A(init), .B(e[344]), .Z(n20856) );
  AND U27344 ( .A(n20857), .B(n20858), .Z(n20855) );
  NAND U27345 ( .A(ereg[343]), .B(n19486), .Z(n20858) );
  NANDN U27346 ( .A(n19481), .B(ereg[344]), .Z(n20857) );
  NAND U27347 ( .A(n20859), .B(n20860), .Z(n15032) );
  NANDN U27348 ( .A(init), .B(e[345]), .Z(n20860) );
  AND U27349 ( .A(n20861), .B(n20862), .Z(n20859) );
  NAND U27350 ( .A(ereg[344]), .B(n19486), .Z(n20862) );
  NANDN U27351 ( .A(n19481), .B(ereg[345]), .Z(n20861) );
  NAND U27352 ( .A(n20863), .B(n20864), .Z(n15031) );
  NANDN U27353 ( .A(init), .B(e[346]), .Z(n20864) );
  AND U27354 ( .A(n20865), .B(n20866), .Z(n20863) );
  NAND U27355 ( .A(ereg[345]), .B(n19486), .Z(n20866) );
  NANDN U27356 ( .A(n19481), .B(ereg[346]), .Z(n20865) );
  NAND U27357 ( .A(n20867), .B(n20868), .Z(n15030) );
  NANDN U27358 ( .A(init), .B(e[347]), .Z(n20868) );
  AND U27359 ( .A(n20869), .B(n20870), .Z(n20867) );
  NAND U27360 ( .A(ereg[346]), .B(n19486), .Z(n20870) );
  NANDN U27361 ( .A(n19481), .B(ereg[347]), .Z(n20869) );
  NAND U27362 ( .A(n20871), .B(n20872), .Z(n15029) );
  NANDN U27363 ( .A(init), .B(e[348]), .Z(n20872) );
  AND U27364 ( .A(n20873), .B(n20874), .Z(n20871) );
  NAND U27365 ( .A(ereg[347]), .B(n19486), .Z(n20874) );
  NANDN U27366 ( .A(n19481), .B(ereg[348]), .Z(n20873) );
  NAND U27367 ( .A(n20875), .B(n20876), .Z(n15028) );
  NANDN U27368 ( .A(init), .B(e[349]), .Z(n20876) );
  AND U27369 ( .A(n20877), .B(n20878), .Z(n20875) );
  NAND U27370 ( .A(ereg[348]), .B(n19486), .Z(n20878) );
  NANDN U27371 ( .A(n19481), .B(ereg[349]), .Z(n20877) );
  NAND U27372 ( .A(n20879), .B(n20880), .Z(n15027) );
  NANDN U27373 ( .A(init), .B(e[350]), .Z(n20880) );
  AND U27374 ( .A(n20881), .B(n20882), .Z(n20879) );
  NAND U27375 ( .A(ereg[349]), .B(n19486), .Z(n20882) );
  NANDN U27376 ( .A(n19481), .B(ereg[350]), .Z(n20881) );
  NAND U27377 ( .A(n20883), .B(n20884), .Z(n15026) );
  NANDN U27378 ( .A(init), .B(e[351]), .Z(n20884) );
  AND U27379 ( .A(n20885), .B(n20886), .Z(n20883) );
  NAND U27380 ( .A(ereg[350]), .B(n19486), .Z(n20886) );
  NANDN U27381 ( .A(n19481), .B(ereg[351]), .Z(n20885) );
  NAND U27382 ( .A(n20887), .B(n20888), .Z(n15025) );
  NANDN U27383 ( .A(init), .B(e[352]), .Z(n20888) );
  AND U27384 ( .A(n20889), .B(n20890), .Z(n20887) );
  NAND U27385 ( .A(ereg[351]), .B(n19486), .Z(n20890) );
  NANDN U27386 ( .A(n19481), .B(ereg[352]), .Z(n20889) );
  NAND U27387 ( .A(n20891), .B(n20892), .Z(n15024) );
  NANDN U27388 ( .A(init), .B(e[353]), .Z(n20892) );
  AND U27389 ( .A(n20893), .B(n20894), .Z(n20891) );
  NAND U27390 ( .A(ereg[352]), .B(n19486), .Z(n20894) );
  NANDN U27391 ( .A(n19481), .B(ereg[353]), .Z(n20893) );
  NAND U27392 ( .A(n20895), .B(n20896), .Z(n15023) );
  NANDN U27393 ( .A(init), .B(e[354]), .Z(n20896) );
  AND U27394 ( .A(n20897), .B(n20898), .Z(n20895) );
  NAND U27395 ( .A(ereg[353]), .B(n19486), .Z(n20898) );
  NANDN U27396 ( .A(n19481), .B(ereg[354]), .Z(n20897) );
  NAND U27397 ( .A(n20899), .B(n20900), .Z(n15022) );
  NANDN U27398 ( .A(init), .B(e[355]), .Z(n20900) );
  AND U27399 ( .A(n20901), .B(n20902), .Z(n20899) );
  NAND U27400 ( .A(ereg[354]), .B(n19486), .Z(n20902) );
  NANDN U27401 ( .A(n19481), .B(ereg[355]), .Z(n20901) );
  NAND U27402 ( .A(n20903), .B(n20904), .Z(n15021) );
  NANDN U27403 ( .A(init), .B(e[356]), .Z(n20904) );
  AND U27404 ( .A(n20905), .B(n20906), .Z(n20903) );
  NAND U27405 ( .A(ereg[355]), .B(n19486), .Z(n20906) );
  NANDN U27406 ( .A(n19481), .B(ereg[356]), .Z(n20905) );
  NAND U27407 ( .A(n20907), .B(n20908), .Z(n15020) );
  NANDN U27408 ( .A(init), .B(e[357]), .Z(n20908) );
  AND U27409 ( .A(n20909), .B(n20910), .Z(n20907) );
  NAND U27410 ( .A(ereg[356]), .B(n19486), .Z(n20910) );
  NANDN U27411 ( .A(n19481), .B(ereg[357]), .Z(n20909) );
  NAND U27412 ( .A(n20911), .B(n20912), .Z(n15019) );
  NANDN U27413 ( .A(init), .B(e[358]), .Z(n20912) );
  AND U27414 ( .A(n20913), .B(n20914), .Z(n20911) );
  NAND U27415 ( .A(ereg[357]), .B(n19486), .Z(n20914) );
  NANDN U27416 ( .A(n19481), .B(ereg[358]), .Z(n20913) );
  NAND U27417 ( .A(n20915), .B(n20916), .Z(n15018) );
  NANDN U27418 ( .A(init), .B(e[359]), .Z(n20916) );
  AND U27419 ( .A(n20917), .B(n20918), .Z(n20915) );
  NAND U27420 ( .A(ereg[358]), .B(n19486), .Z(n20918) );
  NANDN U27421 ( .A(n19481), .B(ereg[359]), .Z(n20917) );
  NAND U27422 ( .A(n20919), .B(n20920), .Z(n15017) );
  NANDN U27423 ( .A(init), .B(e[360]), .Z(n20920) );
  AND U27424 ( .A(n20921), .B(n20922), .Z(n20919) );
  NAND U27425 ( .A(ereg[359]), .B(n19486), .Z(n20922) );
  NANDN U27426 ( .A(n19481), .B(ereg[360]), .Z(n20921) );
  NAND U27427 ( .A(n20923), .B(n20924), .Z(n15016) );
  NANDN U27428 ( .A(init), .B(e[361]), .Z(n20924) );
  AND U27429 ( .A(n20925), .B(n20926), .Z(n20923) );
  NAND U27430 ( .A(ereg[360]), .B(n19486), .Z(n20926) );
  NANDN U27431 ( .A(n19481), .B(ereg[361]), .Z(n20925) );
  NAND U27432 ( .A(n20927), .B(n20928), .Z(n15015) );
  NANDN U27433 ( .A(init), .B(e[362]), .Z(n20928) );
  AND U27434 ( .A(n20929), .B(n20930), .Z(n20927) );
  NAND U27435 ( .A(ereg[361]), .B(n19486), .Z(n20930) );
  NANDN U27436 ( .A(n19481), .B(ereg[362]), .Z(n20929) );
  NAND U27437 ( .A(n20931), .B(n20932), .Z(n15014) );
  NANDN U27438 ( .A(init), .B(e[363]), .Z(n20932) );
  AND U27439 ( .A(n20933), .B(n20934), .Z(n20931) );
  NAND U27440 ( .A(ereg[362]), .B(n19486), .Z(n20934) );
  NANDN U27441 ( .A(n19481), .B(ereg[363]), .Z(n20933) );
  NAND U27442 ( .A(n20935), .B(n20936), .Z(n15013) );
  NANDN U27443 ( .A(init), .B(e[364]), .Z(n20936) );
  AND U27444 ( .A(n20937), .B(n20938), .Z(n20935) );
  NAND U27445 ( .A(ereg[363]), .B(n19486), .Z(n20938) );
  NANDN U27446 ( .A(n19481), .B(ereg[364]), .Z(n20937) );
  NAND U27447 ( .A(n20939), .B(n20940), .Z(n15012) );
  NANDN U27448 ( .A(init), .B(e[365]), .Z(n20940) );
  AND U27449 ( .A(n20941), .B(n20942), .Z(n20939) );
  NAND U27450 ( .A(ereg[364]), .B(n19486), .Z(n20942) );
  NANDN U27451 ( .A(n19481), .B(ereg[365]), .Z(n20941) );
  NAND U27452 ( .A(n20943), .B(n20944), .Z(n15011) );
  NANDN U27453 ( .A(init), .B(e[366]), .Z(n20944) );
  AND U27454 ( .A(n20945), .B(n20946), .Z(n20943) );
  NAND U27455 ( .A(ereg[365]), .B(n19486), .Z(n20946) );
  NANDN U27456 ( .A(n19481), .B(ereg[366]), .Z(n20945) );
  NAND U27457 ( .A(n20947), .B(n20948), .Z(n15010) );
  NANDN U27458 ( .A(init), .B(e[367]), .Z(n20948) );
  AND U27459 ( .A(n20949), .B(n20950), .Z(n20947) );
  NAND U27460 ( .A(ereg[366]), .B(n19486), .Z(n20950) );
  NANDN U27461 ( .A(n19481), .B(ereg[367]), .Z(n20949) );
  NAND U27462 ( .A(n20951), .B(n20952), .Z(n15009) );
  NANDN U27463 ( .A(init), .B(e[368]), .Z(n20952) );
  AND U27464 ( .A(n20953), .B(n20954), .Z(n20951) );
  NAND U27465 ( .A(ereg[367]), .B(n19486), .Z(n20954) );
  NANDN U27466 ( .A(n19481), .B(ereg[368]), .Z(n20953) );
  NAND U27467 ( .A(n20955), .B(n20956), .Z(n15008) );
  NANDN U27468 ( .A(init), .B(e[369]), .Z(n20956) );
  AND U27469 ( .A(n20957), .B(n20958), .Z(n20955) );
  NAND U27470 ( .A(ereg[368]), .B(n19486), .Z(n20958) );
  NANDN U27471 ( .A(n19481), .B(ereg[369]), .Z(n20957) );
  NAND U27472 ( .A(n20959), .B(n20960), .Z(n15007) );
  NANDN U27473 ( .A(init), .B(e[370]), .Z(n20960) );
  AND U27474 ( .A(n20961), .B(n20962), .Z(n20959) );
  NAND U27475 ( .A(ereg[369]), .B(n19486), .Z(n20962) );
  NANDN U27476 ( .A(n19481), .B(ereg[370]), .Z(n20961) );
  NAND U27477 ( .A(n20963), .B(n20964), .Z(n15006) );
  NANDN U27478 ( .A(init), .B(e[371]), .Z(n20964) );
  AND U27479 ( .A(n20965), .B(n20966), .Z(n20963) );
  NAND U27480 ( .A(ereg[370]), .B(n19486), .Z(n20966) );
  NANDN U27481 ( .A(n19481), .B(ereg[371]), .Z(n20965) );
  NAND U27482 ( .A(n20967), .B(n20968), .Z(n15005) );
  NANDN U27483 ( .A(init), .B(e[372]), .Z(n20968) );
  AND U27484 ( .A(n20969), .B(n20970), .Z(n20967) );
  NAND U27485 ( .A(ereg[371]), .B(n19486), .Z(n20970) );
  NANDN U27486 ( .A(n19481), .B(ereg[372]), .Z(n20969) );
  NAND U27487 ( .A(n20971), .B(n20972), .Z(n15004) );
  NANDN U27488 ( .A(init), .B(e[373]), .Z(n20972) );
  AND U27489 ( .A(n20973), .B(n20974), .Z(n20971) );
  NAND U27490 ( .A(ereg[372]), .B(n19486), .Z(n20974) );
  NANDN U27491 ( .A(n19481), .B(ereg[373]), .Z(n20973) );
  NAND U27492 ( .A(n20975), .B(n20976), .Z(n15003) );
  NANDN U27493 ( .A(init), .B(e[374]), .Z(n20976) );
  AND U27494 ( .A(n20977), .B(n20978), .Z(n20975) );
  NAND U27495 ( .A(ereg[373]), .B(n19486), .Z(n20978) );
  NANDN U27496 ( .A(n19481), .B(ereg[374]), .Z(n20977) );
  NAND U27497 ( .A(n20979), .B(n20980), .Z(n15002) );
  NANDN U27498 ( .A(init), .B(e[375]), .Z(n20980) );
  AND U27499 ( .A(n20981), .B(n20982), .Z(n20979) );
  NAND U27500 ( .A(ereg[374]), .B(n19486), .Z(n20982) );
  NANDN U27501 ( .A(n19481), .B(ereg[375]), .Z(n20981) );
  NAND U27502 ( .A(n20983), .B(n20984), .Z(n15001) );
  NANDN U27503 ( .A(init), .B(e[376]), .Z(n20984) );
  AND U27504 ( .A(n20985), .B(n20986), .Z(n20983) );
  NAND U27505 ( .A(ereg[375]), .B(n19486), .Z(n20986) );
  NANDN U27506 ( .A(n19481), .B(ereg[376]), .Z(n20985) );
  NAND U27507 ( .A(n20987), .B(n20988), .Z(n15000) );
  NANDN U27508 ( .A(init), .B(e[377]), .Z(n20988) );
  AND U27509 ( .A(n20989), .B(n20990), .Z(n20987) );
  NAND U27510 ( .A(ereg[376]), .B(n19486), .Z(n20990) );
  NANDN U27511 ( .A(n19481), .B(ereg[377]), .Z(n20989) );
  NAND U27512 ( .A(n20991), .B(n20992), .Z(n14999) );
  NANDN U27513 ( .A(init), .B(e[378]), .Z(n20992) );
  AND U27514 ( .A(n20993), .B(n20994), .Z(n20991) );
  NAND U27515 ( .A(ereg[377]), .B(n19486), .Z(n20994) );
  NANDN U27516 ( .A(n19481), .B(ereg[378]), .Z(n20993) );
  NAND U27517 ( .A(n20995), .B(n20996), .Z(n14998) );
  NANDN U27518 ( .A(init), .B(e[379]), .Z(n20996) );
  AND U27519 ( .A(n20997), .B(n20998), .Z(n20995) );
  NAND U27520 ( .A(ereg[378]), .B(n19486), .Z(n20998) );
  NANDN U27521 ( .A(n19481), .B(ereg[379]), .Z(n20997) );
  NAND U27522 ( .A(n20999), .B(n21000), .Z(n14997) );
  NANDN U27523 ( .A(init), .B(e[380]), .Z(n21000) );
  AND U27524 ( .A(n21001), .B(n21002), .Z(n20999) );
  NAND U27525 ( .A(ereg[379]), .B(n19486), .Z(n21002) );
  NANDN U27526 ( .A(n19481), .B(ereg[380]), .Z(n21001) );
  NAND U27527 ( .A(n21003), .B(n21004), .Z(n14996) );
  NANDN U27528 ( .A(init), .B(e[381]), .Z(n21004) );
  AND U27529 ( .A(n21005), .B(n21006), .Z(n21003) );
  NAND U27530 ( .A(ereg[380]), .B(n19486), .Z(n21006) );
  NANDN U27531 ( .A(n19481), .B(ereg[381]), .Z(n21005) );
  NAND U27532 ( .A(n21007), .B(n21008), .Z(n14995) );
  NANDN U27533 ( .A(init), .B(e[382]), .Z(n21008) );
  AND U27534 ( .A(n21009), .B(n21010), .Z(n21007) );
  NAND U27535 ( .A(ereg[381]), .B(n19486), .Z(n21010) );
  NANDN U27536 ( .A(n19481), .B(ereg[382]), .Z(n21009) );
  NAND U27537 ( .A(n21011), .B(n21012), .Z(n14994) );
  NANDN U27538 ( .A(init), .B(e[383]), .Z(n21012) );
  AND U27539 ( .A(n21013), .B(n21014), .Z(n21011) );
  NAND U27540 ( .A(ereg[382]), .B(n19486), .Z(n21014) );
  NANDN U27541 ( .A(n19481), .B(ereg[383]), .Z(n21013) );
  NAND U27542 ( .A(n21015), .B(n21016), .Z(n14993) );
  NANDN U27543 ( .A(init), .B(e[384]), .Z(n21016) );
  AND U27544 ( .A(n21017), .B(n21018), .Z(n21015) );
  NAND U27545 ( .A(ereg[383]), .B(n19486), .Z(n21018) );
  NANDN U27546 ( .A(n19481), .B(ereg[384]), .Z(n21017) );
  NAND U27547 ( .A(n21019), .B(n21020), .Z(n14992) );
  NANDN U27548 ( .A(init), .B(e[385]), .Z(n21020) );
  AND U27549 ( .A(n21021), .B(n21022), .Z(n21019) );
  NAND U27550 ( .A(ereg[384]), .B(n19486), .Z(n21022) );
  NANDN U27551 ( .A(n19481), .B(ereg[385]), .Z(n21021) );
  NAND U27552 ( .A(n21023), .B(n21024), .Z(n14991) );
  NANDN U27553 ( .A(init), .B(e[386]), .Z(n21024) );
  AND U27554 ( .A(n21025), .B(n21026), .Z(n21023) );
  NAND U27555 ( .A(ereg[385]), .B(n19486), .Z(n21026) );
  NANDN U27556 ( .A(n19481), .B(ereg[386]), .Z(n21025) );
  NAND U27557 ( .A(n21027), .B(n21028), .Z(n14990) );
  NANDN U27558 ( .A(init), .B(e[387]), .Z(n21028) );
  AND U27559 ( .A(n21029), .B(n21030), .Z(n21027) );
  NAND U27560 ( .A(ereg[386]), .B(n19486), .Z(n21030) );
  NANDN U27561 ( .A(n19481), .B(ereg[387]), .Z(n21029) );
  NAND U27562 ( .A(n21031), .B(n21032), .Z(n14989) );
  NANDN U27563 ( .A(init), .B(e[388]), .Z(n21032) );
  AND U27564 ( .A(n21033), .B(n21034), .Z(n21031) );
  NAND U27565 ( .A(ereg[387]), .B(n19486), .Z(n21034) );
  NANDN U27566 ( .A(n19481), .B(ereg[388]), .Z(n21033) );
  NAND U27567 ( .A(n21035), .B(n21036), .Z(n14988) );
  NANDN U27568 ( .A(init), .B(e[389]), .Z(n21036) );
  AND U27569 ( .A(n21037), .B(n21038), .Z(n21035) );
  NAND U27570 ( .A(ereg[388]), .B(n19486), .Z(n21038) );
  NANDN U27571 ( .A(n19481), .B(ereg[389]), .Z(n21037) );
  NAND U27572 ( .A(n21039), .B(n21040), .Z(n14987) );
  NANDN U27573 ( .A(init), .B(e[390]), .Z(n21040) );
  AND U27574 ( .A(n21041), .B(n21042), .Z(n21039) );
  NAND U27575 ( .A(ereg[389]), .B(n19486), .Z(n21042) );
  NANDN U27576 ( .A(n19481), .B(ereg[390]), .Z(n21041) );
  NAND U27577 ( .A(n21043), .B(n21044), .Z(n14986) );
  NANDN U27578 ( .A(init), .B(e[391]), .Z(n21044) );
  AND U27579 ( .A(n21045), .B(n21046), .Z(n21043) );
  NAND U27580 ( .A(ereg[390]), .B(n19486), .Z(n21046) );
  NANDN U27581 ( .A(n19481), .B(ereg[391]), .Z(n21045) );
  NAND U27582 ( .A(n21047), .B(n21048), .Z(n14985) );
  NANDN U27583 ( .A(init), .B(e[392]), .Z(n21048) );
  AND U27584 ( .A(n21049), .B(n21050), .Z(n21047) );
  NAND U27585 ( .A(ereg[391]), .B(n19486), .Z(n21050) );
  NANDN U27586 ( .A(n19481), .B(ereg[392]), .Z(n21049) );
  NAND U27587 ( .A(n21051), .B(n21052), .Z(n14984) );
  NANDN U27588 ( .A(init), .B(e[393]), .Z(n21052) );
  AND U27589 ( .A(n21053), .B(n21054), .Z(n21051) );
  NAND U27590 ( .A(ereg[392]), .B(n19486), .Z(n21054) );
  NANDN U27591 ( .A(n19481), .B(ereg[393]), .Z(n21053) );
  NAND U27592 ( .A(n21055), .B(n21056), .Z(n14983) );
  NANDN U27593 ( .A(init), .B(e[394]), .Z(n21056) );
  AND U27594 ( .A(n21057), .B(n21058), .Z(n21055) );
  NAND U27595 ( .A(ereg[393]), .B(n19486), .Z(n21058) );
  NANDN U27596 ( .A(n19481), .B(ereg[394]), .Z(n21057) );
  NAND U27597 ( .A(n21059), .B(n21060), .Z(n14982) );
  NANDN U27598 ( .A(init), .B(e[395]), .Z(n21060) );
  AND U27599 ( .A(n21061), .B(n21062), .Z(n21059) );
  NAND U27600 ( .A(ereg[394]), .B(n19486), .Z(n21062) );
  NANDN U27601 ( .A(n19481), .B(ereg[395]), .Z(n21061) );
  NAND U27602 ( .A(n21063), .B(n21064), .Z(n14981) );
  NANDN U27603 ( .A(init), .B(e[396]), .Z(n21064) );
  AND U27604 ( .A(n21065), .B(n21066), .Z(n21063) );
  NAND U27605 ( .A(ereg[395]), .B(n19486), .Z(n21066) );
  NANDN U27606 ( .A(n19481), .B(ereg[396]), .Z(n21065) );
  NAND U27607 ( .A(n21067), .B(n21068), .Z(n14980) );
  NANDN U27608 ( .A(init), .B(e[397]), .Z(n21068) );
  AND U27609 ( .A(n21069), .B(n21070), .Z(n21067) );
  NAND U27610 ( .A(ereg[396]), .B(n19486), .Z(n21070) );
  NANDN U27611 ( .A(n19481), .B(ereg[397]), .Z(n21069) );
  NAND U27612 ( .A(n21071), .B(n21072), .Z(n14979) );
  NANDN U27613 ( .A(init), .B(e[398]), .Z(n21072) );
  AND U27614 ( .A(n21073), .B(n21074), .Z(n21071) );
  NAND U27615 ( .A(ereg[397]), .B(n19486), .Z(n21074) );
  NANDN U27616 ( .A(n19481), .B(ereg[398]), .Z(n21073) );
  NAND U27617 ( .A(n21075), .B(n21076), .Z(n14978) );
  NANDN U27618 ( .A(init), .B(e[399]), .Z(n21076) );
  AND U27619 ( .A(n21077), .B(n21078), .Z(n21075) );
  NAND U27620 ( .A(ereg[398]), .B(n19486), .Z(n21078) );
  NANDN U27621 ( .A(n19481), .B(ereg[399]), .Z(n21077) );
  NAND U27622 ( .A(n21079), .B(n21080), .Z(n14977) );
  NANDN U27623 ( .A(init), .B(e[400]), .Z(n21080) );
  AND U27624 ( .A(n21081), .B(n21082), .Z(n21079) );
  NAND U27625 ( .A(ereg[399]), .B(n19486), .Z(n21082) );
  NANDN U27626 ( .A(n19481), .B(ereg[400]), .Z(n21081) );
  NAND U27627 ( .A(n21083), .B(n21084), .Z(n14976) );
  NANDN U27628 ( .A(init), .B(e[401]), .Z(n21084) );
  AND U27629 ( .A(n21085), .B(n21086), .Z(n21083) );
  NAND U27630 ( .A(ereg[400]), .B(n19486), .Z(n21086) );
  NANDN U27631 ( .A(n19481), .B(ereg[401]), .Z(n21085) );
  NAND U27632 ( .A(n21087), .B(n21088), .Z(n14975) );
  NANDN U27633 ( .A(init), .B(e[402]), .Z(n21088) );
  AND U27634 ( .A(n21089), .B(n21090), .Z(n21087) );
  NAND U27635 ( .A(ereg[401]), .B(n19486), .Z(n21090) );
  NANDN U27636 ( .A(n19481), .B(ereg[402]), .Z(n21089) );
  NAND U27637 ( .A(n21091), .B(n21092), .Z(n14974) );
  NANDN U27638 ( .A(init), .B(e[403]), .Z(n21092) );
  AND U27639 ( .A(n21093), .B(n21094), .Z(n21091) );
  NAND U27640 ( .A(ereg[402]), .B(n19486), .Z(n21094) );
  NANDN U27641 ( .A(n19481), .B(ereg[403]), .Z(n21093) );
  NAND U27642 ( .A(n21095), .B(n21096), .Z(n14973) );
  NANDN U27643 ( .A(init), .B(e[404]), .Z(n21096) );
  AND U27644 ( .A(n21097), .B(n21098), .Z(n21095) );
  NAND U27645 ( .A(ereg[403]), .B(n19486), .Z(n21098) );
  NANDN U27646 ( .A(n19481), .B(ereg[404]), .Z(n21097) );
  NAND U27647 ( .A(n21099), .B(n21100), .Z(n14972) );
  NANDN U27648 ( .A(init), .B(e[405]), .Z(n21100) );
  AND U27649 ( .A(n21101), .B(n21102), .Z(n21099) );
  NAND U27650 ( .A(ereg[404]), .B(n19486), .Z(n21102) );
  NANDN U27651 ( .A(n19481), .B(ereg[405]), .Z(n21101) );
  NAND U27652 ( .A(n21103), .B(n21104), .Z(n14971) );
  NANDN U27653 ( .A(init), .B(e[406]), .Z(n21104) );
  AND U27654 ( .A(n21105), .B(n21106), .Z(n21103) );
  NAND U27655 ( .A(ereg[405]), .B(n19486), .Z(n21106) );
  NANDN U27656 ( .A(n19481), .B(ereg[406]), .Z(n21105) );
  NAND U27657 ( .A(n21107), .B(n21108), .Z(n14970) );
  NANDN U27658 ( .A(init), .B(e[407]), .Z(n21108) );
  AND U27659 ( .A(n21109), .B(n21110), .Z(n21107) );
  NAND U27660 ( .A(ereg[406]), .B(n19486), .Z(n21110) );
  NANDN U27661 ( .A(n19481), .B(ereg[407]), .Z(n21109) );
  NAND U27662 ( .A(n21111), .B(n21112), .Z(n14969) );
  NANDN U27663 ( .A(init), .B(e[408]), .Z(n21112) );
  AND U27664 ( .A(n21113), .B(n21114), .Z(n21111) );
  NAND U27665 ( .A(ereg[407]), .B(n19486), .Z(n21114) );
  NANDN U27666 ( .A(n19481), .B(ereg[408]), .Z(n21113) );
  NAND U27667 ( .A(n21115), .B(n21116), .Z(n14968) );
  NANDN U27668 ( .A(init), .B(e[409]), .Z(n21116) );
  AND U27669 ( .A(n21117), .B(n21118), .Z(n21115) );
  NAND U27670 ( .A(ereg[408]), .B(n19486), .Z(n21118) );
  NANDN U27671 ( .A(n19481), .B(ereg[409]), .Z(n21117) );
  NAND U27672 ( .A(n21119), .B(n21120), .Z(n14967) );
  NANDN U27673 ( .A(init), .B(e[410]), .Z(n21120) );
  AND U27674 ( .A(n21121), .B(n21122), .Z(n21119) );
  NAND U27675 ( .A(ereg[409]), .B(n19486), .Z(n21122) );
  NANDN U27676 ( .A(n19481), .B(ereg[410]), .Z(n21121) );
  NAND U27677 ( .A(n21123), .B(n21124), .Z(n14966) );
  NANDN U27678 ( .A(init), .B(e[411]), .Z(n21124) );
  AND U27679 ( .A(n21125), .B(n21126), .Z(n21123) );
  NAND U27680 ( .A(ereg[410]), .B(n19486), .Z(n21126) );
  NANDN U27681 ( .A(n19481), .B(ereg[411]), .Z(n21125) );
  NAND U27682 ( .A(n21127), .B(n21128), .Z(n14965) );
  NANDN U27683 ( .A(init), .B(e[412]), .Z(n21128) );
  AND U27684 ( .A(n21129), .B(n21130), .Z(n21127) );
  NAND U27685 ( .A(ereg[411]), .B(n19486), .Z(n21130) );
  NANDN U27686 ( .A(n19481), .B(ereg[412]), .Z(n21129) );
  NAND U27687 ( .A(n21131), .B(n21132), .Z(n14964) );
  NANDN U27688 ( .A(init), .B(e[413]), .Z(n21132) );
  AND U27689 ( .A(n21133), .B(n21134), .Z(n21131) );
  NAND U27690 ( .A(ereg[412]), .B(n19486), .Z(n21134) );
  NANDN U27691 ( .A(n19481), .B(ereg[413]), .Z(n21133) );
  NAND U27692 ( .A(n21135), .B(n21136), .Z(n14963) );
  NANDN U27693 ( .A(init), .B(e[414]), .Z(n21136) );
  AND U27694 ( .A(n21137), .B(n21138), .Z(n21135) );
  NAND U27695 ( .A(ereg[413]), .B(n19486), .Z(n21138) );
  NANDN U27696 ( .A(n19481), .B(ereg[414]), .Z(n21137) );
  NAND U27697 ( .A(n21139), .B(n21140), .Z(n14962) );
  NANDN U27698 ( .A(init), .B(e[415]), .Z(n21140) );
  AND U27699 ( .A(n21141), .B(n21142), .Z(n21139) );
  NAND U27700 ( .A(ereg[414]), .B(n19486), .Z(n21142) );
  NANDN U27701 ( .A(n19481), .B(ereg[415]), .Z(n21141) );
  NAND U27702 ( .A(n21143), .B(n21144), .Z(n14961) );
  NANDN U27703 ( .A(init), .B(e[416]), .Z(n21144) );
  AND U27704 ( .A(n21145), .B(n21146), .Z(n21143) );
  NAND U27705 ( .A(ereg[415]), .B(n19486), .Z(n21146) );
  NANDN U27706 ( .A(n19481), .B(ereg[416]), .Z(n21145) );
  NAND U27707 ( .A(n21147), .B(n21148), .Z(n14960) );
  NANDN U27708 ( .A(init), .B(e[417]), .Z(n21148) );
  AND U27709 ( .A(n21149), .B(n21150), .Z(n21147) );
  NAND U27710 ( .A(ereg[416]), .B(n19486), .Z(n21150) );
  NANDN U27711 ( .A(n19481), .B(ereg[417]), .Z(n21149) );
  NAND U27712 ( .A(n21151), .B(n21152), .Z(n14959) );
  NANDN U27713 ( .A(init), .B(e[418]), .Z(n21152) );
  AND U27714 ( .A(n21153), .B(n21154), .Z(n21151) );
  NAND U27715 ( .A(ereg[417]), .B(n19486), .Z(n21154) );
  NANDN U27716 ( .A(n19481), .B(ereg[418]), .Z(n21153) );
  NAND U27717 ( .A(n21155), .B(n21156), .Z(n14958) );
  NANDN U27718 ( .A(init), .B(e[419]), .Z(n21156) );
  AND U27719 ( .A(n21157), .B(n21158), .Z(n21155) );
  NAND U27720 ( .A(ereg[418]), .B(n19486), .Z(n21158) );
  NANDN U27721 ( .A(n19481), .B(ereg[419]), .Z(n21157) );
  NAND U27722 ( .A(n21159), .B(n21160), .Z(n14957) );
  NANDN U27723 ( .A(init), .B(e[420]), .Z(n21160) );
  AND U27724 ( .A(n21161), .B(n21162), .Z(n21159) );
  NAND U27725 ( .A(ereg[419]), .B(n19486), .Z(n21162) );
  NANDN U27726 ( .A(n19481), .B(ereg[420]), .Z(n21161) );
  NAND U27727 ( .A(n21163), .B(n21164), .Z(n14956) );
  NANDN U27728 ( .A(init), .B(e[421]), .Z(n21164) );
  AND U27729 ( .A(n21165), .B(n21166), .Z(n21163) );
  NAND U27730 ( .A(ereg[420]), .B(n19486), .Z(n21166) );
  NANDN U27731 ( .A(n19481), .B(ereg[421]), .Z(n21165) );
  NAND U27732 ( .A(n21167), .B(n21168), .Z(n14955) );
  NANDN U27733 ( .A(init), .B(e[422]), .Z(n21168) );
  AND U27734 ( .A(n21169), .B(n21170), .Z(n21167) );
  NAND U27735 ( .A(ereg[421]), .B(n19486), .Z(n21170) );
  NANDN U27736 ( .A(n19481), .B(ereg[422]), .Z(n21169) );
  NAND U27737 ( .A(n21171), .B(n21172), .Z(n14954) );
  NANDN U27738 ( .A(init), .B(e[423]), .Z(n21172) );
  AND U27739 ( .A(n21173), .B(n21174), .Z(n21171) );
  NAND U27740 ( .A(ereg[422]), .B(n19486), .Z(n21174) );
  NANDN U27741 ( .A(n19481), .B(ereg[423]), .Z(n21173) );
  NAND U27742 ( .A(n21175), .B(n21176), .Z(n14953) );
  NANDN U27743 ( .A(init), .B(e[424]), .Z(n21176) );
  AND U27744 ( .A(n21177), .B(n21178), .Z(n21175) );
  NAND U27745 ( .A(ereg[423]), .B(n19486), .Z(n21178) );
  NANDN U27746 ( .A(n19481), .B(ereg[424]), .Z(n21177) );
  NAND U27747 ( .A(n21179), .B(n21180), .Z(n14952) );
  NANDN U27748 ( .A(init), .B(e[425]), .Z(n21180) );
  AND U27749 ( .A(n21181), .B(n21182), .Z(n21179) );
  NAND U27750 ( .A(ereg[424]), .B(n19486), .Z(n21182) );
  NANDN U27751 ( .A(n19481), .B(ereg[425]), .Z(n21181) );
  NAND U27752 ( .A(n21183), .B(n21184), .Z(n14951) );
  NANDN U27753 ( .A(init), .B(e[426]), .Z(n21184) );
  AND U27754 ( .A(n21185), .B(n21186), .Z(n21183) );
  NAND U27755 ( .A(ereg[425]), .B(n19486), .Z(n21186) );
  NANDN U27756 ( .A(n19481), .B(ereg[426]), .Z(n21185) );
  NAND U27757 ( .A(n21187), .B(n21188), .Z(n14950) );
  NANDN U27758 ( .A(init), .B(e[427]), .Z(n21188) );
  AND U27759 ( .A(n21189), .B(n21190), .Z(n21187) );
  NAND U27760 ( .A(ereg[426]), .B(n19486), .Z(n21190) );
  NANDN U27761 ( .A(n19481), .B(ereg[427]), .Z(n21189) );
  NAND U27762 ( .A(n21191), .B(n21192), .Z(n14949) );
  NANDN U27763 ( .A(init), .B(e[428]), .Z(n21192) );
  AND U27764 ( .A(n21193), .B(n21194), .Z(n21191) );
  NAND U27765 ( .A(ereg[427]), .B(n19486), .Z(n21194) );
  NANDN U27766 ( .A(n19481), .B(ereg[428]), .Z(n21193) );
  NAND U27767 ( .A(n21195), .B(n21196), .Z(n14948) );
  NANDN U27768 ( .A(init), .B(e[429]), .Z(n21196) );
  AND U27769 ( .A(n21197), .B(n21198), .Z(n21195) );
  NAND U27770 ( .A(ereg[428]), .B(n19486), .Z(n21198) );
  NANDN U27771 ( .A(n19481), .B(ereg[429]), .Z(n21197) );
  NAND U27772 ( .A(n21199), .B(n21200), .Z(n14947) );
  NANDN U27773 ( .A(init), .B(e[430]), .Z(n21200) );
  AND U27774 ( .A(n21201), .B(n21202), .Z(n21199) );
  NAND U27775 ( .A(ereg[429]), .B(n19486), .Z(n21202) );
  NANDN U27776 ( .A(n19481), .B(ereg[430]), .Z(n21201) );
  NAND U27777 ( .A(n21203), .B(n21204), .Z(n14946) );
  NANDN U27778 ( .A(init), .B(e[431]), .Z(n21204) );
  AND U27779 ( .A(n21205), .B(n21206), .Z(n21203) );
  NAND U27780 ( .A(ereg[430]), .B(n19486), .Z(n21206) );
  NANDN U27781 ( .A(n19481), .B(ereg[431]), .Z(n21205) );
  NAND U27782 ( .A(n21207), .B(n21208), .Z(n14945) );
  NANDN U27783 ( .A(init), .B(e[432]), .Z(n21208) );
  AND U27784 ( .A(n21209), .B(n21210), .Z(n21207) );
  NAND U27785 ( .A(ereg[431]), .B(n19486), .Z(n21210) );
  NANDN U27786 ( .A(n19481), .B(ereg[432]), .Z(n21209) );
  NAND U27787 ( .A(n21211), .B(n21212), .Z(n14944) );
  NANDN U27788 ( .A(init), .B(e[433]), .Z(n21212) );
  AND U27789 ( .A(n21213), .B(n21214), .Z(n21211) );
  NAND U27790 ( .A(ereg[432]), .B(n19486), .Z(n21214) );
  NANDN U27791 ( .A(n19481), .B(ereg[433]), .Z(n21213) );
  NAND U27792 ( .A(n21215), .B(n21216), .Z(n14943) );
  NANDN U27793 ( .A(init), .B(e[434]), .Z(n21216) );
  AND U27794 ( .A(n21217), .B(n21218), .Z(n21215) );
  NAND U27795 ( .A(ereg[433]), .B(n19486), .Z(n21218) );
  NANDN U27796 ( .A(n19481), .B(ereg[434]), .Z(n21217) );
  NAND U27797 ( .A(n21219), .B(n21220), .Z(n14942) );
  NANDN U27798 ( .A(init), .B(e[435]), .Z(n21220) );
  AND U27799 ( .A(n21221), .B(n21222), .Z(n21219) );
  NAND U27800 ( .A(ereg[434]), .B(n19486), .Z(n21222) );
  NANDN U27801 ( .A(n19481), .B(ereg[435]), .Z(n21221) );
  NAND U27802 ( .A(n21223), .B(n21224), .Z(n14941) );
  NANDN U27803 ( .A(init), .B(e[436]), .Z(n21224) );
  AND U27804 ( .A(n21225), .B(n21226), .Z(n21223) );
  NAND U27805 ( .A(ereg[435]), .B(n19486), .Z(n21226) );
  NANDN U27806 ( .A(n19481), .B(ereg[436]), .Z(n21225) );
  NAND U27807 ( .A(n21227), .B(n21228), .Z(n14940) );
  NANDN U27808 ( .A(init), .B(e[437]), .Z(n21228) );
  AND U27809 ( .A(n21229), .B(n21230), .Z(n21227) );
  NAND U27810 ( .A(ereg[436]), .B(n19486), .Z(n21230) );
  NANDN U27811 ( .A(n19481), .B(ereg[437]), .Z(n21229) );
  NAND U27812 ( .A(n21231), .B(n21232), .Z(n14939) );
  NANDN U27813 ( .A(init), .B(e[438]), .Z(n21232) );
  AND U27814 ( .A(n21233), .B(n21234), .Z(n21231) );
  NAND U27815 ( .A(ereg[437]), .B(n19486), .Z(n21234) );
  NANDN U27816 ( .A(n19481), .B(ereg[438]), .Z(n21233) );
  NAND U27817 ( .A(n21235), .B(n21236), .Z(n14938) );
  NANDN U27818 ( .A(init), .B(e[439]), .Z(n21236) );
  AND U27819 ( .A(n21237), .B(n21238), .Z(n21235) );
  NAND U27820 ( .A(ereg[438]), .B(n19486), .Z(n21238) );
  NANDN U27821 ( .A(n19481), .B(ereg[439]), .Z(n21237) );
  NAND U27822 ( .A(n21239), .B(n21240), .Z(n14937) );
  NANDN U27823 ( .A(init), .B(e[440]), .Z(n21240) );
  AND U27824 ( .A(n21241), .B(n21242), .Z(n21239) );
  NAND U27825 ( .A(ereg[439]), .B(n19486), .Z(n21242) );
  NANDN U27826 ( .A(n19481), .B(ereg[440]), .Z(n21241) );
  NAND U27827 ( .A(n21243), .B(n21244), .Z(n14936) );
  NANDN U27828 ( .A(init), .B(e[441]), .Z(n21244) );
  AND U27829 ( .A(n21245), .B(n21246), .Z(n21243) );
  NAND U27830 ( .A(ereg[440]), .B(n19486), .Z(n21246) );
  NANDN U27831 ( .A(n19481), .B(ereg[441]), .Z(n21245) );
  NAND U27832 ( .A(n21247), .B(n21248), .Z(n14935) );
  NANDN U27833 ( .A(init), .B(e[442]), .Z(n21248) );
  AND U27834 ( .A(n21249), .B(n21250), .Z(n21247) );
  NAND U27835 ( .A(ereg[441]), .B(n19486), .Z(n21250) );
  NANDN U27836 ( .A(n19481), .B(ereg[442]), .Z(n21249) );
  NAND U27837 ( .A(n21251), .B(n21252), .Z(n14934) );
  NANDN U27838 ( .A(init), .B(e[443]), .Z(n21252) );
  AND U27839 ( .A(n21253), .B(n21254), .Z(n21251) );
  NAND U27840 ( .A(ereg[442]), .B(n19486), .Z(n21254) );
  NANDN U27841 ( .A(n19481), .B(ereg[443]), .Z(n21253) );
  NAND U27842 ( .A(n21255), .B(n21256), .Z(n14933) );
  NANDN U27843 ( .A(init), .B(e[444]), .Z(n21256) );
  AND U27844 ( .A(n21257), .B(n21258), .Z(n21255) );
  NAND U27845 ( .A(ereg[443]), .B(n19486), .Z(n21258) );
  NANDN U27846 ( .A(n19481), .B(ereg[444]), .Z(n21257) );
  NAND U27847 ( .A(n21259), .B(n21260), .Z(n14932) );
  NANDN U27848 ( .A(init), .B(e[445]), .Z(n21260) );
  AND U27849 ( .A(n21261), .B(n21262), .Z(n21259) );
  NAND U27850 ( .A(ereg[444]), .B(n19486), .Z(n21262) );
  NANDN U27851 ( .A(n19481), .B(ereg[445]), .Z(n21261) );
  NAND U27852 ( .A(n21263), .B(n21264), .Z(n14931) );
  NANDN U27853 ( .A(init), .B(e[446]), .Z(n21264) );
  AND U27854 ( .A(n21265), .B(n21266), .Z(n21263) );
  NAND U27855 ( .A(ereg[445]), .B(n19486), .Z(n21266) );
  NANDN U27856 ( .A(n19481), .B(ereg[446]), .Z(n21265) );
  NAND U27857 ( .A(n21267), .B(n21268), .Z(n14930) );
  NANDN U27858 ( .A(init), .B(e[447]), .Z(n21268) );
  AND U27859 ( .A(n21269), .B(n21270), .Z(n21267) );
  NAND U27860 ( .A(ereg[446]), .B(n19486), .Z(n21270) );
  NANDN U27861 ( .A(n19481), .B(ereg[447]), .Z(n21269) );
  NAND U27862 ( .A(n21271), .B(n21272), .Z(n14929) );
  NANDN U27863 ( .A(init), .B(e[448]), .Z(n21272) );
  AND U27864 ( .A(n21273), .B(n21274), .Z(n21271) );
  NAND U27865 ( .A(ereg[447]), .B(n19486), .Z(n21274) );
  NANDN U27866 ( .A(n19481), .B(ereg[448]), .Z(n21273) );
  NAND U27867 ( .A(n21275), .B(n21276), .Z(n14928) );
  NANDN U27868 ( .A(init), .B(e[449]), .Z(n21276) );
  AND U27869 ( .A(n21277), .B(n21278), .Z(n21275) );
  NAND U27870 ( .A(ereg[448]), .B(n19486), .Z(n21278) );
  NANDN U27871 ( .A(n19481), .B(ereg[449]), .Z(n21277) );
  NAND U27872 ( .A(n21279), .B(n21280), .Z(n14927) );
  NANDN U27873 ( .A(init), .B(e[450]), .Z(n21280) );
  AND U27874 ( .A(n21281), .B(n21282), .Z(n21279) );
  NAND U27875 ( .A(ereg[449]), .B(n19486), .Z(n21282) );
  NANDN U27876 ( .A(n19481), .B(ereg[450]), .Z(n21281) );
  NAND U27877 ( .A(n21283), .B(n21284), .Z(n14926) );
  NANDN U27878 ( .A(init), .B(e[451]), .Z(n21284) );
  AND U27879 ( .A(n21285), .B(n21286), .Z(n21283) );
  NAND U27880 ( .A(ereg[450]), .B(n19486), .Z(n21286) );
  NANDN U27881 ( .A(n19481), .B(ereg[451]), .Z(n21285) );
  NAND U27882 ( .A(n21287), .B(n21288), .Z(n14925) );
  NANDN U27883 ( .A(init), .B(e[452]), .Z(n21288) );
  AND U27884 ( .A(n21289), .B(n21290), .Z(n21287) );
  NAND U27885 ( .A(ereg[451]), .B(n19486), .Z(n21290) );
  NANDN U27886 ( .A(n19481), .B(ereg[452]), .Z(n21289) );
  NAND U27887 ( .A(n21291), .B(n21292), .Z(n14924) );
  NANDN U27888 ( .A(init), .B(e[453]), .Z(n21292) );
  AND U27889 ( .A(n21293), .B(n21294), .Z(n21291) );
  NAND U27890 ( .A(ereg[452]), .B(n19486), .Z(n21294) );
  NANDN U27891 ( .A(n19481), .B(ereg[453]), .Z(n21293) );
  NAND U27892 ( .A(n21295), .B(n21296), .Z(n14923) );
  NANDN U27893 ( .A(init), .B(e[454]), .Z(n21296) );
  AND U27894 ( .A(n21297), .B(n21298), .Z(n21295) );
  NAND U27895 ( .A(ereg[453]), .B(n19486), .Z(n21298) );
  NANDN U27896 ( .A(n19481), .B(ereg[454]), .Z(n21297) );
  NAND U27897 ( .A(n21299), .B(n21300), .Z(n14922) );
  NANDN U27898 ( .A(init), .B(e[455]), .Z(n21300) );
  AND U27899 ( .A(n21301), .B(n21302), .Z(n21299) );
  NAND U27900 ( .A(ereg[454]), .B(n19486), .Z(n21302) );
  NANDN U27901 ( .A(n19481), .B(ereg[455]), .Z(n21301) );
  NAND U27902 ( .A(n21303), .B(n21304), .Z(n14921) );
  NANDN U27903 ( .A(init), .B(e[456]), .Z(n21304) );
  AND U27904 ( .A(n21305), .B(n21306), .Z(n21303) );
  NAND U27905 ( .A(ereg[455]), .B(n19486), .Z(n21306) );
  NANDN U27906 ( .A(n19481), .B(ereg[456]), .Z(n21305) );
  NAND U27907 ( .A(n21307), .B(n21308), .Z(n14920) );
  NANDN U27908 ( .A(init), .B(e[457]), .Z(n21308) );
  AND U27909 ( .A(n21309), .B(n21310), .Z(n21307) );
  NAND U27910 ( .A(ereg[456]), .B(n19486), .Z(n21310) );
  NANDN U27911 ( .A(n19481), .B(ereg[457]), .Z(n21309) );
  NAND U27912 ( .A(n21311), .B(n21312), .Z(n14919) );
  NANDN U27913 ( .A(init), .B(e[458]), .Z(n21312) );
  AND U27914 ( .A(n21313), .B(n21314), .Z(n21311) );
  NAND U27915 ( .A(ereg[457]), .B(n19486), .Z(n21314) );
  NANDN U27916 ( .A(n19481), .B(ereg[458]), .Z(n21313) );
  NAND U27917 ( .A(n21315), .B(n21316), .Z(n14918) );
  NANDN U27918 ( .A(init), .B(e[459]), .Z(n21316) );
  AND U27919 ( .A(n21317), .B(n21318), .Z(n21315) );
  NAND U27920 ( .A(ereg[458]), .B(n19486), .Z(n21318) );
  NANDN U27921 ( .A(n19481), .B(ereg[459]), .Z(n21317) );
  NAND U27922 ( .A(n21319), .B(n21320), .Z(n14917) );
  NANDN U27923 ( .A(init), .B(e[460]), .Z(n21320) );
  AND U27924 ( .A(n21321), .B(n21322), .Z(n21319) );
  NAND U27925 ( .A(ereg[459]), .B(n19486), .Z(n21322) );
  NANDN U27926 ( .A(n19481), .B(ereg[460]), .Z(n21321) );
  NAND U27927 ( .A(n21323), .B(n21324), .Z(n14916) );
  NANDN U27928 ( .A(init), .B(e[461]), .Z(n21324) );
  AND U27929 ( .A(n21325), .B(n21326), .Z(n21323) );
  NAND U27930 ( .A(ereg[460]), .B(n19486), .Z(n21326) );
  NANDN U27931 ( .A(n19481), .B(ereg[461]), .Z(n21325) );
  NAND U27932 ( .A(n21327), .B(n21328), .Z(n14915) );
  NANDN U27933 ( .A(init), .B(e[462]), .Z(n21328) );
  AND U27934 ( .A(n21329), .B(n21330), .Z(n21327) );
  NAND U27935 ( .A(ereg[461]), .B(n19486), .Z(n21330) );
  NANDN U27936 ( .A(n19481), .B(ereg[462]), .Z(n21329) );
  NAND U27937 ( .A(n21331), .B(n21332), .Z(n14914) );
  NANDN U27938 ( .A(init), .B(e[463]), .Z(n21332) );
  AND U27939 ( .A(n21333), .B(n21334), .Z(n21331) );
  NAND U27940 ( .A(ereg[462]), .B(n19486), .Z(n21334) );
  NANDN U27941 ( .A(n19481), .B(ereg[463]), .Z(n21333) );
  NAND U27942 ( .A(n21335), .B(n21336), .Z(n14913) );
  NANDN U27943 ( .A(init), .B(e[464]), .Z(n21336) );
  AND U27944 ( .A(n21337), .B(n21338), .Z(n21335) );
  NAND U27945 ( .A(ereg[463]), .B(n19486), .Z(n21338) );
  NANDN U27946 ( .A(n19481), .B(ereg[464]), .Z(n21337) );
  NAND U27947 ( .A(n21339), .B(n21340), .Z(n14912) );
  NANDN U27948 ( .A(init), .B(e[465]), .Z(n21340) );
  AND U27949 ( .A(n21341), .B(n21342), .Z(n21339) );
  NAND U27950 ( .A(ereg[464]), .B(n19486), .Z(n21342) );
  NANDN U27951 ( .A(n19481), .B(ereg[465]), .Z(n21341) );
  NAND U27952 ( .A(n21343), .B(n21344), .Z(n14911) );
  NANDN U27953 ( .A(init), .B(e[466]), .Z(n21344) );
  AND U27954 ( .A(n21345), .B(n21346), .Z(n21343) );
  NAND U27955 ( .A(ereg[465]), .B(n19486), .Z(n21346) );
  NANDN U27956 ( .A(n19481), .B(ereg[466]), .Z(n21345) );
  NAND U27957 ( .A(n21347), .B(n21348), .Z(n14910) );
  NANDN U27958 ( .A(init), .B(e[467]), .Z(n21348) );
  AND U27959 ( .A(n21349), .B(n21350), .Z(n21347) );
  NAND U27960 ( .A(ereg[466]), .B(n19486), .Z(n21350) );
  NANDN U27961 ( .A(n19481), .B(ereg[467]), .Z(n21349) );
  NAND U27962 ( .A(n21351), .B(n21352), .Z(n14909) );
  NANDN U27963 ( .A(init), .B(e[468]), .Z(n21352) );
  AND U27964 ( .A(n21353), .B(n21354), .Z(n21351) );
  NAND U27965 ( .A(ereg[467]), .B(n19486), .Z(n21354) );
  NANDN U27966 ( .A(n19481), .B(ereg[468]), .Z(n21353) );
  NAND U27967 ( .A(n21355), .B(n21356), .Z(n14908) );
  NANDN U27968 ( .A(init), .B(e[469]), .Z(n21356) );
  AND U27969 ( .A(n21357), .B(n21358), .Z(n21355) );
  NAND U27970 ( .A(ereg[468]), .B(n19486), .Z(n21358) );
  NANDN U27971 ( .A(n19481), .B(ereg[469]), .Z(n21357) );
  NAND U27972 ( .A(n21359), .B(n21360), .Z(n14907) );
  NANDN U27973 ( .A(init), .B(e[470]), .Z(n21360) );
  AND U27974 ( .A(n21361), .B(n21362), .Z(n21359) );
  NAND U27975 ( .A(ereg[469]), .B(n19486), .Z(n21362) );
  NANDN U27976 ( .A(n19481), .B(ereg[470]), .Z(n21361) );
  NAND U27977 ( .A(n21363), .B(n21364), .Z(n14906) );
  NANDN U27978 ( .A(init), .B(e[471]), .Z(n21364) );
  AND U27979 ( .A(n21365), .B(n21366), .Z(n21363) );
  NAND U27980 ( .A(ereg[470]), .B(n19486), .Z(n21366) );
  NANDN U27981 ( .A(n19481), .B(ereg[471]), .Z(n21365) );
  NAND U27982 ( .A(n21367), .B(n21368), .Z(n14905) );
  NANDN U27983 ( .A(init), .B(e[472]), .Z(n21368) );
  AND U27984 ( .A(n21369), .B(n21370), .Z(n21367) );
  NAND U27985 ( .A(ereg[471]), .B(n19486), .Z(n21370) );
  NANDN U27986 ( .A(n19481), .B(ereg[472]), .Z(n21369) );
  NAND U27987 ( .A(n21371), .B(n21372), .Z(n14904) );
  NANDN U27988 ( .A(init), .B(e[473]), .Z(n21372) );
  AND U27989 ( .A(n21373), .B(n21374), .Z(n21371) );
  NAND U27990 ( .A(ereg[472]), .B(n19486), .Z(n21374) );
  NANDN U27991 ( .A(n19481), .B(ereg[473]), .Z(n21373) );
  NAND U27992 ( .A(n21375), .B(n21376), .Z(n14903) );
  NANDN U27993 ( .A(init), .B(e[474]), .Z(n21376) );
  AND U27994 ( .A(n21377), .B(n21378), .Z(n21375) );
  NAND U27995 ( .A(ereg[473]), .B(n19486), .Z(n21378) );
  NANDN U27996 ( .A(n19481), .B(ereg[474]), .Z(n21377) );
  NAND U27997 ( .A(n21379), .B(n21380), .Z(n14902) );
  NANDN U27998 ( .A(init), .B(e[475]), .Z(n21380) );
  AND U27999 ( .A(n21381), .B(n21382), .Z(n21379) );
  NAND U28000 ( .A(ereg[474]), .B(n19486), .Z(n21382) );
  NANDN U28001 ( .A(n19481), .B(ereg[475]), .Z(n21381) );
  NAND U28002 ( .A(n21383), .B(n21384), .Z(n14901) );
  NANDN U28003 ( .A(init), .B(e[476]), .Z(n21384) );
  AND U28004 ( .A(n21385), .B(n21386), .Z(n21383) );
  NAND U28005 ( .A(ereg[475]), .B(n19486), .Z(n21386) );
  NANDN U28006 ( .A(n19481), .B(ereg[476]), .Z(n21385) );
  NAND U28007 ( .A(n21387), .B(n21388), .Z(n14900) );
  NANDN U28008 ( .A(init), .B(e[477]), .Z(n21388) );
  AND U28009 ( .A(n21389), .B(n21390), .Z(n21387) );
  NAND U28010 ( .A(ereg[476]), .B(n19486), .Z(n21390) );
  NANDN U28011 ( .A(n19481), .B(ereg[477]), .Z(n21389) );
  NAND U28012 ( .A(n21391), .B(n21392), .Z(n14899) );
  NANDN U28013 ( .A(init), .B(e[478]), .Z(n21392) );
  AND U28014 ( .A(n21393), .B(n21394), .Z(n21391) );
  NAND U28015 ( .A(ereg[477]), .B(n19486), .Z(n21394) );
  NANDN U28016 ( .A(n19481), .B(ereg[478]), .Z(n21393) );
  NAND U28017 ( .A(n21395), .B(n21396), .Z(n14898) );
  NANDN U28018 ( .A(init), .B(e[479]), .Z(n21396) );
  AND U28019 ( .A(n21397), .B(n21398), .Z(n21395) );
  NAND U28020 ( .A(ereg[478]), .B(n19486), .Z(n21398) );
  NANDN U28021 ( .A(n19481), .B(ereg[479]), .Z(n21397) );
  NAND U28022 ( .A(n21399), .B(n21400), .Z(n14897) );
  NANDN U28023 ( .A(init), .B(e[480]), .Z(n21400) );
  AND U28024 ( .A(n21401), .B(n21402), .Z(n21399) );
  NAND U28025 ( .A(ereg[479]), .B(n19486), .Z(n21402) );
  NANDN U28026 ( .A(n19481), .B(ereg[480]), .Z(n21401) );
  NAND U28027 ( .A(n21403), .B(n21404), .Z(n14896) );
  NANDN U28028 ( .A(init), .B(e[481]), .Z(n21404) );
  AND U28029 ( .A(n21405), .B(n21406), .Z(n21403) );
  NAND U28030 ( .A(ereg[480]), .B(n19486), .Z(n21406) );
  NANDN U28031 ( .A(n19481), .B(ereg[481]), .Z(n21405) );
  NAND U28032 ( .A(n21407), .B(n21408), .Z(n14895) );
  NANDN U28033 ( .A(init), .B(e[482]), .Z(n21408) );
  AND U28034 ( .A(n21409), .B(n21410), .Z(n21407) );
  NAND U28035 ( .A(ereg[481]), .B(n19486), .Z(n21410) );
  NANDN U28036 ( .A(n19481), .B(ereg[482]), .Z(n21409) );
  NAND U28037 ( .A(n21411), .B(n21412), .Z(n14894) );
  NANDN U28038 ( .A(init), .B(e[483]), .Z(n21412) );
  AND U28039 ( .A(n21413), .B(n21414), .Z(n21411) );
  NAND U28040 ( .A(ereg[482]), .B(n19486), .Z(n21414) );
  NANDN U28041 ( .A(n19481), .B(ereg[483]), .Z(n21413) );
  NAND U28042 ( .A(n21415), .B(n21416), .Z(n14893) );
  NANDN U28043 ( .A(init), .B(e[484]), .Z(n21416) );
  AND U28044 ( .A(n21417), .B(n21418), .Z(n21415) );
  NAND U28045 ( .A(ereg[483]), .B(n19486), .Z(n21418) );
  NANDN U28046 ( .A(n19481), .B(ereg[484]), .Z(n21417) );
  NAND U28047 ( .A(n21419), .B(n21420), .Z(n14892) );
  NANDN U28048 ( .A(init), .B(e[485]), .Z(n21420) );
  AND U28049 ( .A(n21421), .B(n21422), .Z(n21419) );
  NAND U28050 ( .A(ereg[484]), .B(n19486), .Z(n21422) );
  NANDN U28051 ( .A(n19481), .B(ereg[485]), .Z(n21421) );
  NAND U28052 ( .A(n21423), .B(n21424), .Z(n14891) );
  NANDN U28053 ( .A(init), .B(e[486]), .Z(n21424) );
  AND U28054 ( .A(n21425), .B(n21426), .Z(n21423) );
  NAND U28055 ( .A(ereg[485]), .B(n19486), .Z(n21426) );
  NANDN U28056 ( .A(n19481), .B(ereg[486]), .Z(n21425) );
  NAND U28057 ( .A(n21427), .B(n21428), .Z(n14890) );
  NANDN U28058 ( .A(init), .B(e[487]), .Z(n21428) );
  AND U28059 ( .A(n21429), .B(n21430), .Z(n21427) );
  NAND U28060 ( .A(ereg[486]), .B(n19486), .Z(n21430) );
  NANDN U28061 ( .A(n19481), .B(ereg[487]), .Z(n21429) );
  NAND U28062 ( .A(n21431), .B(n21432), .Z(n14889) );
  NANDN U28063 ( .A(init), .B(e[488]), .Z(n21432) );
  AND U28064 ( .A(n21433), .B(n21434), .Z(n21431) );
  NAND U28065 ( .A(ereg[487]), .B(n19486), .Z(n21434) );
  NANDN U28066 ( .A(n19481), .B(ereg[488]), .Z(n21433) );
  NAND U28067 ( .A(n21435), .B(n21436), .Z(n14888) );
  NANDN U28068 ( .A(init), .B(e[489]), .Z(n21436) );
  AND U28069 ( .A(n21437), .B(n21438), .Z(n21435) );
  NAND U28070 ( .A(ereg[488]), .B(n19486), .Z(n21438) );
  NANDN U28071 ( .A(n19481), .B(ereg[489]), .Z(n21437) );
  NAND U28072 ( .A(n21439), .B(n21440), .Z(n14887) );
  NANDN U28073 ( .A(init), .B(e[490]), .Z(n21440) );
  AND U28074 ( .A(n21441), .B(n21442), .Z(n21439) );
  NAND U28075 ( .A(ereg[489]), .B(n19486), .Z(n21442) );
  NANDN U28076 ( .A(n19481), .B(ereg[490]), .Z(n21441) );
  NAND U28077 ( .A(n21443), .B(n21444), .Z(n14886) );
  NANDN U28078 ( .A(init), .B(e[491]), .Z(n21444) );
  AND U28079 ( .A(n21445), .B(n21446), .Z(n21443) );
  NAND U28080 ( .A(ereg[490]), .B(n19486), .Z(n21446) );
  NANDN U28081 ( .A(n19481), .B(ereg[491]), .Z(n21445) );
  NAND U28082 ( .A(n21447), .B(n21448), .Z(n14885) );
  NANDN U28083 ( .A(init), .B(e[492]), .Z(n21448) );
  AND U28084 ( .A(n21449), .B(n21450), .Z(n21447) );
  NAND U28085 ( .A(ereg[491]), .B(n19486), .Z(n21450) );
  NANDN U28086 ( .A(n19481), .B(ereg[492]), .Z(n21449) );
  NAND U28087 ( .A(n21451), .B(n21452), .Z(n14884) );
  NANDN U28088 ( .A(init), .B(e[493]), .Z(n21452) );
  AND U28089 ( .A(n21453), .B(n21454), .Z(n21451) );
  NAND U28090 ( .A(ereg[492]), .B(n19486), .Z(n21454) );
  NANDN U28091 ( .A(n19481), .B(ereg[493]), .Z(n21453) );
  NAND U28092 ( .A(n21455), .B(n21456), .Z(n14883) );
  NANDN U28093 ( .A(init), .B(e[494]), .Z(n21456) );
  AND U28094 ( .A(n21457), .B(n21458), .Z(n21455) );
  NAND U28095 ( .A(ereg[493]), .B(n19486), .Z(n21458) );
  NANDN U28096 ( .A(n19481), .B(ereg[494]), .Z(n21457) );
  NAND U28097 ( .A(n21459), .B(n21460), .Z(n14882) );
  NANDN U28098 ( .A(init), .B(e[495]), .Z(n21460) );
  AND U28099 ( .A(n21461), .B(n21462), .Z(n21459) );
  NAND U28100 ( .A(ereg[494]), .B(n19486), .Z(n21462) );
  NANDN U28101 ( .A(n19481), .B(ereg[495]), .Z(n21461) );
  NAND U28102 ( .A(n21463), .B(n21464), .Z(n14881) );
  NANDN U28103 ( .A(init), .B(e[496]), .Z(n21464) );
  AND U28104 ( .A(n21465), .B(n21466), .Z(n21463) );
  NAND U28105 ( .A(ereg[495]), .B(n19486), .Z(n21466) );
  NANDN U28106 ( .A(n19481), .B(ereg[496]), .Z(n21465) );
  NAND U28107 ( .A(n21467), .B(n21468), .Z(n14880) );
  NANDN U28108 ( .A(init), .B(e[497]), .Z(n21468) );
  AND U28109 ( .A(n21469), .B(n21470), .Z(n21467) );
  NAND U28110 ( .A(ereg[496]), .B(n19486), .Z(n21470) );
  NANDN U28111 ( .A(n19481), .B(ereg[497]), .Z(n21469) );
  NAND U28112 ( .A(n21471), .B(n21472), .Z(n14879) );
  NANDN U28113 ( .A(init), .B(e[498]), .Z(n21472) );
  AND U28114 ( .A(n21473), .B(n21474), .Z(n21471) );
  NAND U28115 ( .A(ereg[497]), .B(n19486), .Z(n21474) );
  NANDN U28116 ( .A(n19481), .B(ereg[498]), .Z(n21473) );
  NAND U28117 ( .A(n21475), .B(n21476), .Z(n14878) );
  NANDN U28118 ( .A(init), .B(e[499]), .Z(n21476) );
  AND U28119 ( .A(n21477), .B(n21478), .Z(n21475) );
  NAND U28120 ( .A(ereg[498]), .B(n19486), .Z(n21478) );
  NANDN U28121 ( .A(n19481), .B(ereg[499]), .Z(n21477) );
  NAND U28122 ( .A(n21479), .B(n21480), .Z(n14877) );
  NANDN U28123 ( .A(init), .B(e[500]), .Z(n21480) );
  AND U28124 ( .A(n21481), .B(n21482), .Z(n21479) );
  NAND U28125 ( .A(ereg[499]), .B(n19486), .Z(n21482) );
  NANDN U28126 ( .A(n19481), .B(ereg[500]), .Z(n21481) );
  NAND U28127 ( .A(n21483), .B(n21484), .Z(n14876) );
  NANDN U28128 ( .A(init), .B(e[501]), .Z(n21484) );
  AND U28129 ( .A(n21485), .B(n21486), .Z(n21483) );
  NAND U28130 ( .A(ereg[500]), .B(n19486), .Z(n21486) );
  NANDN U28131 ( .A(n19481), .B(ereg[501]), .Z(n21485) );
  NAND U28132 ( .A(n21487), .B(n21488), .Z(n14875) );
  NANDN U28133 ( .A(init), .B(e[502]), .Z(n21488) );
  AND U28134 ( .A(n21489), .B(n21490), .Z(n21487) );
  NAND U28135 ( .A(ereg[501]), .B(n19486), .Z(n21490) );
  NANDN U28136 ( .A(n19481), .B(ereg[502]), .Z(n21489) );
  NAND U28137 ( .A(n21491), .B(n21492), .Z(n14874) );
  NANDN U28138 ( .A(init), .B(e[503]), .Z(n21492) );
  AND U28139 ( .A(n21493), .B(n21494), .Z(n21491) );
  NAND U28140 ( .A(ereg[502]), .B(n19486), .Z(n21494) );
  NANDN U28141 ( .A(n19481), .B(ereg[503]), .Z(n21493) );
  NAND U28142 ( .A(n21495), .B(n21496), .Z(n14873) );
  NANDN U28143 ( .A(init), .B(e[504]), .Z(n21496) );
  AND U28144 ( .A(n21497), .B(n21498), .Z(n21495) );
  NAND U28145 ( .A(ereg[503]), .B(n19486), .Z(n21498) );
  NANDN U28146 ( .A(n19481), .B(ereg[504]), .Z(n21497) );
  NAND U28147 ( .A(n21499), .B(n21500), .Z(n14872) );
  NANDN U28148 ( .A(init), .B(e[505]), .Z(n21500) );
  AND U28149 ( .A(n21501), .B(n21502), .Z(n21499) );
  NAND U28150 ( .A(ereg[504]), .B(n19486), .Z(n21502) );
  NANDN U28151 ( .A(n19481), .B(ereg[505]), .Z(n21501) );
  NAND U28152 ( .A(n21503), .B(n21504), .Z(n14871) );
  NANDN U28153 ( .A(init), .B(e[506]), .Z(n21504) );
  AND U28154 ( .A(n21505), .B(n21506), .Z(n21503) );
  NAND U28155 ( .A(ereg[505]), .B(n19486), .Z(n21506) );
  NANDN U28156 ( .A(n19481), .B(ereg[506]), .Z(n21505) );
  NAND U28157 ( .A(n21507), .B(n21508), .Z(n14870) );
  NANDN U28158 ( .A(init), .B(e[507]), .Z(n21508) );
  AND U28159 ( .A(n21509), .B(n21510), .Z(n21507) );
  NAND U28160 ( .A(ereg[506]), .B(n19486), .Z(n21510) );
  NANDN U28161 ( .A(n19481), .B(ereg[507]), .Z(n21509) );
  NAND U28162 ( .A(n21511), .B(n21512), .Z(n14869) );
  NANDN U28163 ( .A(init), .B(e[508]), .Z(n21512) );
  AND U28164 ( .A(n21513), .B(n21514), .Z(n21511) );
  NAND U28165 ( .A(ereg[507]), .B(n19486), .Z(n21514) );
  NANDN U28166 ( .A(n19481), .B(ereg[508]), .Z(n21513) );
  NAND U28167 ( .A(n21515), .B(n21516), .Z(n14868) );
  NANDN U28168 ( .A(init), .B(e[509]), .Z(n21516) );
  AND U28169 ( .A(n21517), .B(n21518), .Z(n21515) );
  NAND U28170 ( .A(ereg[508]), .B(n19486), .Z(n21518) );
  NANDN U28171 ( .A(n19481), .B(ereg[509]), .Z(n21517) );
  NAND U28172 ( .A(n21519), .B(n21520), .Z(n14867) );
  NANDN U28173 ( .A(init), .B(e[510]), .Z(n21520) );
  AND U28174 ( .A(n21521), .B(n21522), .Z(n21519) );
  NAND U28175 ( .A(ereg[509]), .B(n19486), .Z(n21522) );
  NANDN U28176 ( .A(n19481), .B(ereg[510]), .Z(n21521) );
  NAND U28177 ( .A(n21523), .B(n21524), .Z(n14866) );
  NANDN U28178 ( .A(init), .B(e[511]), .Z(n21524) );
  AND U28179 ( .A(n21525), .B(n21526), .Z(n21523) );
  NAND U28180 ( .A(ereg[510]), .B(n19486), .Z(n21526) );
  NANDN U28181 ( .A(n19481), .B(ereg[511]), .Z(n21525) );
  NAND U28182 ( .A(n21527), .B(n21528), .Z(n14865) );
  NANDN U28183 ( .A(init), .B(e[512]), .Z(n21528) );
  AND U28184 ( .A(n21529), .B(n21530), .Z(n21527) );
  NAND U28185 ( .A(ereg[511]), .B(n19486), .Z(n21530) );
  NANDN U28186 ( .A(n19481), .B(ereg[512]), .Z(n21529) );
  NAND U28187 ( .A(n21531), .B(n21532), .Z(n14864) );
  NANDN U28188 ( .A(init), .B(e[513]), .Z(n21532) );
  AND U28189 ( .A(n21533), .B(n21534), .Z(n21531) );
  NAND U28190 ( .A(ereg[512]), .B(n19486), .Z(n21534) );
  NANDN U28191 ( .A(n19481), .B(ereg[513]), .Z(n21533) );
  NAND U28192 ( .A(n21535), .B(n21536), .Z(n14863) );
  NANDN U28193 ( .A(init), .B(e[514]), .Z(n21536) );
  AND U28194 ( .A(n21537), .B(n21538), .Z(n21535) );
  NAND U28195 ( .A(ereg[513]), .B(n19486), .Z(n21538) );
  NANDN U28196 ( .A(n19481), .B(ereg[514]), .Z(n21537) );
  NAND U28197 ( .A(n21539), .B(n21540), .Z(n14862) );
  NANDN U28198 ( .A(init), .B(e[515]), .Z(n21540) );
  AND U28199 ( .A(n21541), .B(n21542), .Z(n21539) );
  NAND U28200 ( .A(ereg[514]), .B(n19486), .Z(n21542) );
  NANDN U28201 ( .A(n19481), .B(ereg[515]), .Z(n21541) );
  NAND U28202 ( .A(n21543), .B(n21544), .Z(n14861) );
  NANDN U28203 ( .A(init), .B(e[516]), .Z(n21544) );
  AND U28204 ( .A(n21545), .B(n21546), .Z(n21543) );
  NAND U28205 ( .A(ereg[515]), .B(n19486), .Z(n21546) );
  NANDN U28206 ( .A(n19481), .B(ereg[516]), .Z(n21545) );
  NAND U28207 ( .A(n21547), .B(n21548), .Z(n14860) );
  NANDN U28208 ( .A(init), .B(e[517]), .Z(n21548) );
  AND U28209 ( .A(n21549), .B(n21550), .Z(n21547) );
  NAND U28210 ( .A(ereg[516]), .B(n19486), .Z(n21550) );
  NANDN U28211 ( .A(n19481), .B(ereg[517]), .Z(n21549) );
  NAND U28212 ( .A(n21551), .B(n21552), .Z(n14859) );
  NANDN U28213 ( .A(init), .B(e[518]), .Z(n21552) );
  AND U28214 ( .A(n21553), .B(n21554), .Z(n21551) );
  NAND U28215 ( .A(ereg[517]), .B(n19486), .Z(n21554) );
  NANDN U28216 ( .A(n19481), .B(ereg[518]), .Z(n21553) );
  NAND U28217 ( .A(n21555), .B(n21556), .Z(n14858) );
  NANDN U28218 ( .A(init), .B(e[519]), .Z(n21556) );
  AND U28219 ( .A(n21557), .B(n21558), .Z(n21555) );
  NAND U28220 ( .A(ereg[518]), .B(n19486), .Z(n21558) );
  NANDN U28221 ( .A(n19481), .B(ereg[519]), .Z(n21557) );
  NAND U28222 ( .A(n21559), .B(n21560), .Z(n14857) );
  NANDN U28223 ( .A(init), .B(e[520]), .Z(n21560) );
  AND U28224 ( .A(n21561), .B(n21562), .Z(n21559) );
  NAND U28225 ( .A(ereg[519]), .B(n19486), .Z(n21562) );
  NANDN U28226 ( .A(n19481), .B(ereg[520]), .Z(n21561) );
  NAND U28227 ( .A(n21563), .B(n21564), .Z(n14856) );
  NANDN U28228 ( .A(init), .B(e[521]), .Z(n21564) );
  AND U28229 ( .A(n21565), .B(n21566), .Z(n21563) );
  NAND U28230 ( .A(ereg[520]), .B(n19486), .Z(n21566) );
  NANDN U28231 ( .A(n19481), .B(ereg[521]), .Z(n21565) );
  NAND U28232 ( .A(n21567), .B(n21568), .Z(n14855) );
  NANDN U28233 ( .A(init), .B(e[522]), .Z(n21568) );
  AND U28234 ( .A(n21569), .B(n21570), .Z(n21567) );
  NAND U28235 ( .A(ereg[521]), .B(n19486), .Z(n21570) );
  NANDN U28236 ( .A(n19481), .B(ereg[522]), .Z(n21569) );
  NAND U28237 ( .A(n21571), .B(n21572), .Z(n14854) );
  NANDN U28238 ( .A(init), .B(e[523]), .Z(n21572) );
  AND U28239 ( .A(n21573), .B(n21574), .Z(n21571) );
  NAND U28240 ( .A(ereg[522]), .B(n19486), .Z(n21574) );
  NANDN U28241 ( .A(n19481), .B(ereg[523]), .Z(n21573) );
  NAND U28242 ( .A(n21575), .B(n21576), .Z(n14853) );
  NANDN U28243 ( .A(init), .B(e[524]), .Z(n21576) );
  AND U28244 ( .A(n21577), .B(n21578), .Z(n21575) );
  NAND U28245 ( .A(ereg[523]), .B(n19486), .Z(n21578) );
  NANDN U28246 ( .A(n19481), .B(ereg[524]), .Z(n21577) );
  NAND U28247 ( .A(n21579), .B(n21580), .Z(n14852) );
  NANDN U28248 ( .A(init), .B(e[525]), .Z(n21580) );
  AND U28249 ( .A(n21581), .B(n21582), .Z(n21579) );
  NAND U28250 ( .A(ereg[524]), .B(n19486), .Z(n21582) );
  NANDN U28251 ( .A(n19481), .B(ereg[525]), .Z(n21581) );
  NAND U28252 ( .A(n21583), .B(n21584), .Z(n14851) );
  NANDN U28253 ( .A(init), .B(e[526]), .Z(n21584) );
  AND U28254 ( .A(n21585), .B(n21586), .Z(n21583) );
  NAND U28255 ( .A(ereg[525]), .B(n19486), .Z(n21586) );
  NANDN U28256 ( .A(n19481), .B(ereg[526]), .Z(n21585) );
  NAND U28257 ( .A(n21587), .B(n21588), .Z(n14850) );
  NANDN U28258 ( .A(init), .B(e[527]), .Z(n21588) );
  AND U28259 ( .A(n21589), .B(n21590), .Z(n21587) );
  NAND U28260 ( .A(ereg[526]), .B(n19486), .Z(n21590) );
  NANDN U28261 ( .A(n19481), .B(ereg[527]), .Z(n21589) );
  NAND U28262 ( .A(n21591), .B(n21592), .Z(n14849) );
  NANDN U28263 ( .A(init), .B(e[528]), .Z(n21592) );
  AND U28264 ( .A(n21593), .B(n21594), .Z(n21591) );
  NAND U28265 ( .A(ereg[527]), .B(n19486), .Z(n21594) );
  NANDN U28266 ( .A(n19481), .B(ereg[528]), .Z(n21593) );
  NAND U28267 ( .A(n21595), .B(n21596), .Z(n14848) );
  NANDN U28268 ( .A(init), .B(e[529]), .Z(n21596) );
  AND U28269 ( .A(n21597), .B(n21598), .Z(n21595) );
  NAND U28270 ( .A(ereg[528]), .B(n19486), .Z(n21598) );
  NANDN U28271 ( .A(n19481), .B(ereg[529]), .Z(n21597) );
  NAND U28272 ( .A(n21599), .B(n21600), .Z(n14847) );
  NANDN U28273 ( .A(init), .B(e[530]), .Z(n21600) );
  AND U28274 ( .A(n21601), .B(n21602), .Z(n21599) );
  NAND U28275 ( .A(ereg[529]), .B(n19486), .Z(n21602) );
  NANDN U28276 ( .A(n19481), .B(ereg[530]), .Z(n21601) );
  NAND U28277 ( .A(n21603), .B(n21604), .Z(n14846) );
  NANDN U28278 ( .A(init), .B(e[531]), .Z(n21604) );
  AND U28279 ( .A(n21605), .B(n21606), .Z(n21603) );
  NAND U28280 ( .A(ereg[530]), .B(n19486), .Z(n21606) );
  NANDN U28281 ( .A(n19481), .B(ereg[531]), .Z(n21605) );
  NAND U28282 ( .A(n21607), .B(n21608), .Z(n14845) );
  NANDN U28283 ( .A(init), .B(e[532]), .Z(n21608) );
  AND U28284 ( .A(n21609), .B(n21610), .Z(n21607) );
  NAND U28285 ( .A(ereg[531]), .B(n19486), .Z(n21610) );
  NANDN U28286 ( .A(n19481), .B(ereg[532]), .Z(n21609) );
  NAND U28287 ( .A(n21611), .B(n21612), .Z(n14844) );
  NANDN U28288 ( .A(init), .B(e[533]), .Z(n21612) );
  AND U28289 ( .A(n21613), .B(n21614), .Z(n21611) );
  NAND U28290 ( .A(ereg[532]), .B(n19486), .Z(n21614) );
  NANDN U28291 ( .A(n19481), .B(ereg[533]), .Z(n21613) );
  NAND U28292 ( .A(n21615), .B(n21616), .Z(n14843) );
  NANDN U28293 ( .A(init), .B(e[534]), .Z(n21616) );
  AND U28294 ( .A(n21617), .B(n21618), .Z(n21615) );
  NAND U28295 ( .A(ereg[533]), .B(n19486), .Z(n21618) );
  NANDN U28296 ( .A(n19481), .B(ereg[534]), .Z(n21617) );
  NAND U28297 ( .A(n21619), .B(n21620), .Z(n14842) );
  NANDN U28298 ( .A(init), .B(e[535]), .Z(n21620) );
  AND U28299 ( .A(n21621), .B(n21622), .Z(n21619) );
  NAND U28300 ( .A(ereg[534]), .B(n19486), .Z(n21622) );
  NANDN U28301 ( .A(n19481), .B(ereg[535]), .Z(n21621) );
  NAND U28302 ( .A(n21623), .B(n21624), .Z(n14841) );
  NANDN U28303 ( .A(init), .B(e[536]), .Z(n21624) );
  AND U28304 ( .A(n21625), .B(n21626), .Z(n21623) );
  NAND U28305 ( .A(ereg[535]), .B(n19486), .Z(n21626) );
  NANDN U28306 ( .A(n19481), .B(ereg[536]), .Z(n21625) );
  NAND U28307 ( .A(n21627), .B(n21628), .Z(n14840) );
  NANDN U28308 ( .A(init), .B(e[537]), .Z(n21628) );
  AND U28309 ( .A(n21629), .B(n21630), .Z(n21627) );
  NAND U28310 ( .A(ereg[536]), .B(n19486), .Z(n21630) );
  NANDN U28311 ( .A(n19481), .B(ereg[537]), .Z(n21629) );
  NAND U28312 ( .A(n21631), .B(n21632), .Z(n14839) );
  NANDN U28313 ( .A(init), .B(e[538]), .Z(n21632) );
  AND U28314 ( .A(n21633), .B(n21634), .Z(n21631) );
  NAND U28315 ( .A(ereg[537]), .B(n19486), .Z(n21634) );
  NANDN U28316 ( .A(n19481), .B(ereg[538]), .Z(n21633) );
  NAND U28317 ( .A(n21635), .B(n21636), .Z(n14838) );
  NANDN U28318 ( .A(init), .B(e[539]), .Z(n21636) );
  AND U28319 ( .A(n21637), .B(n21638), .Z(n21635) );
  NAND U28320 ( .A(ereg[538]), .B(n19486), .Z(n21638) );
  NANDN U28321 ( .A(n19481), .B(ereg[539]), .Z(n21637) );
  NAND U28322 ( .A(n21639), .B(n21640), .Z(n14837) );
  NANDN U28323 ( .A(init), .B(e[540]), .Z(n21640) );
  AND U28324 ( .A(n21641), .B(n21642), .Z(n21639) );
  NAND U28325 ( .A(ereg[539]), .B(n19486), .Z(n21642) );
  NANDN U28326 ( .A(n19481), .B(ereg[540]), .Z(n21641) );
  NAND U28327 ( .A(n21643), .B(n21644), .Z(n14836) );
  NANDN U28328 ( .A(init), .B(e[541]), .Z(n21644) );
  AND U28329 ( .A(n21645), .B(n21646), .Z(n21643) );
  NAND U28330 ( .A(ereg[540]), .B(n19486), .Z(n21646) );
  NANDN U28331 ( .A(n19481), .B(ereg[541]), .Z(n21645) );
  NAND U28332 ( .A(n21647), .B(n21648), .Z(n14835) );
  NANDN U28333 ( .A(init), .B(e[542]), .Z(n21648) );
  AND U28334 ( .A(n21649), .B(n21650), .Z(n21647) );
  NAND U28335 ( .A(ereg[541]), .B(n19486), .Z(n21650) );
  NANDN U28336 ( .A(n19481), .B(ereg[542]), .Z(n21649) );
  NAND U28337 ( .A(n21651), .B(n21652), .Z(n14834) );
  NANDN U28338 ( .A(init), .B(e[543]), .Z(n21652) );
  AND U28339 ( .A(n21653), .B(n21654), .Z(n21651) );
  NAND U28340 ( .A(ereg[542]), .B(n19486), .Z(n21654) );
  NANDN U28341 ( .A(n19481), .B(ereg[543]), .Z(n21653) );
  NAND U28342 ( .A(n21655), .B(n21656), .Z(n14833) );
  NANDN U28343 ( .A(init), .B(e[544]), .Z(n21656) );
  AND U28344 ( .A(n21657), .B(n21658), .Z(n21655) );
  NAND U28345 ( .A(ereg[543]), .B(n19486), .Z(n21658) );
  NANDN U28346 ( .A(n19481), .B(ereg[544]), .Z(n21657) );
  NAND U28347 ( .A(n21659), .B(n21660), .Z(n14832) );
  NANDN U28348 ( .A(init), .B(e[545]), .Z(n21660) );
  AND U28349 ( .A(n21661), .B(n21662), .Z(n21659) );
  NAND U28350 ( .A(ereg[544]), .B(n19486), .Z(n21662) );
  NANDN U28351 ( .A(n19481), .B(ereg[545]), .Z(n21661) );
  NAND U28352 ( .A(n21663), .B(n21664), .Z(n14831) );
  NANDN U28353 ( .A(init), .B(e[546]), .Z(n21664) );
  AND U28354 ( .A(n21665), .B(n21666), .Z(n21663) );
  NAND U28355 ( .A(ereg[545]), .B(n19486), .Z(n21666) );
  NANDN U28356 ( .A(n19481), .B(ereg[546]), .Z(n21665) );
  NAND U28357 ( .A(n21667), .B(n21668), .Z(n14830) );
  NANDN U28358 ( .A(init), .B(e[547]), .Z(n21668) );
  AND U28359 ( .A(n21669), .B(n21670), .Z(n21667) );
  NAND U28360 ( .A(ereg[546]), .B(n19486), .Z(n21670) );
  NANDN U28361 ( .A(n19481), .B(ereg[547]), .Z(n21669) );
  NAND U28362 ( .A(n21671), .B(n21672), .Z(n14829) );
  NANDN U28363 ( .A(init), .B(e[548]), .Z(n21672) );
  AND U28364 ( .A(n21673), .B(n21674), .Z(n21671) );
  NAND U28365 ( .A(ereg[547]), .B(n19486), .Z(n21674) );
  NANDN U28366 ( .A(n19481), .B(ereg[548]), .Z(n21673) );
  NAND U28367 ( .A(n21675), .B(n21676), .Z(n14828) );
  NANDN U28368 ( .A(init), .B(e[549]), .Z(n21676) );
  AND U28369 ( .A(n21677), .B(n21678), .Z(n21675) );
  NAND U28370 ( .A(ereg[548]), .B(n19486), .Z(n21678) );
  NANDN U28371 ( .A(n19481), .B(ereg[549]), .Z(n21677) );
  NAND U28372 ( .A(n21679), .B(n21680), .Z(n14827) );
  NANDN U28373 ( .A(init), .B(e[550]), .Z(n21680) );
  AND U28374 ( .A(n21681), .B(n21682), .Z(n21679) );
  NAND U28375 ( .A(ereg[549]), .B(n19486), .Z(n21682) );
  NANDN U28376 ( .A(n19481), .B(ereg[550]), .Z(n21681) );
  NAND U28377 ( .A(n21683), .B(n21684), .Z(n14826) );
  NANDN U28378 ( .A(init), .B(e[551]), .Z(n21684) );
  AND U28379 ( .A(n21685), .B(n21686), .Z(n21683) );
  NAND U28380 ( .A(ereg[550]), .B(n19486), .Z(n21686) );
  NANDN U28381 ( .A(n19481), .B(ereg[551]), .Z(n21685) );
  NAND U28382 ( .A(n21687), .B(n21688), .Z(n14825) );
  NANDN U28383 ( .A(init), .B(e[552]), .Z(n21688) );
  AND U28384 ( .A(n21689), .B(n21690), .Z(n21687) );
  NAND U28385 ( .A(ereg[551]), .B(n19486), .Z(n21690) );
  NANDN U28386 ( .A(n19481), .B(ereg[552]), .Z(n21689) );
  NAND U28387 ( .A(n21691), .B(n21692), .Z(n14824) );
  NANDN U28388 ( .A(init), .B(e[553]), .Z(n21692) );
  AND U28389 ( .A(n21693), .B(n21694), .Z(n21691) );
  NAND U28390 ( .A(ereg[552]), .B(n19486), .Z(n21694) );
  NANDN U28391 ( .A(n19481), .B(ereg[553]), .Z(n21693) );
  NAND U28392 ( .A(n21695), .B(n21696), .Z(n14823) );
  NANDN U28393 ( .A(init), .B(e[554]), .Z(n21696) );
  AND U28394 ( .A(n21697), .B(n21698), .Z(n21695) );
  NAND U28395 ( .A(ereg[553]), .B(n19486), .Z(n21698) );
  NANDN U28396 ( .A(n19481), .B(ereg[554]), .Z(n21697) );
  NAND U28397 ( .A(n21699), .B(n21700), .Z(n14822) );
  NANDN U28398 ( .A(init), .B(e[555]), .Z(n21700) );
  AND U28399 ( .A(n21701), .B(n21702), .Z(n21699) );
  NAND U28400 ( .A(ereg[554]), .B(n19486), .Z(n21702) );
  NANDN U28401 ( .A(n19481), .B(ereg[555]), .Z(n21701) );
  NAND U28402 ( .A(n21703), .B(n21704), .Z(n14821) );
  NANDN U28403 ( .A(init), .B(e[556]), .Z(n21704) );
  AND U28404 ( .A(n21705), .B(n21706), .Z(n21703) );
  NAND U28405 ( .A(ereg[555]), .B(n19486), .Z(n21706) );
  NANDN U28406 ( .A(n19481), .B(ereg[556]), .Z(n21705) );
  NAND U28407 ( .A(n21707), .B(n21708), .Z(n14820) );
  NANDN U28408 ( .A(init), .B(e[557]), .Z(n21708) );
  AND U28409 ( .A(n21709), .B(n21710), .Z(n21707) );
  NAND U28410 ( .A(ereg[556]), .B(n19486), .Z(n21710) );
  NANDN U28411 ( .A(n19481), .B(ereg[557]), .Z(n21709) );
  NAND U28412 ( .A(n21711), .B(n21712), .Z(n14819) );
  NANDN U28413 ( .A(init), .B(e[558]), .Z(n21712) );
  AND U28414 ( .A(n21713), .B(n21714), .Z(n21711) );
  NAND U28415 ( .A(ereg[557]), .B(n19486), .Z(n21714) );
  NANDN U28416 ( .A(n19481), .B(ereg[558]), .Z(n21713) );
  NAND U28417 ( .A(n21715), .B(n21716), .Z(n14818) );
  NANDN U28418 ( .A(init), .B(e[559]), .Z(n21716) );
  AND U28419 ( .A(n21717), .B(n21718), .Z(n21715) );
  NAND U28420 ( .A(ereg[558]), .B(n19486), .Z(n21718) );
  NANDN U28421 ( .A(n19481), .B(ereg[559]), .Z(n21717) );
  NAND U28422 ( .A(n21719), .B(n21720), .Z(n14817) );
  NANDN U28423 ( .A(init), .B(e[560]), .Z(n21720) );
  AND U28424 ( .A(n21721), .B(n21722), .Z(n21719) );
  NAND U28425 ( .A(ereg[559]), .B(n19486), .Z(n21722) );
  NANDN U28426 ( .A(n19481), .B(ereg[560]), .Z(n21721) );
  NAND U28427 ( .A(n21723), .B(n21724), .Z(n14816) );
  NANDN U28428 ( .A(init), .B(e[561]), .Z(n21724) );
  AND U28429 ( .A(n21725), .B(n21726), .Z(n21723) );
  NAND U28430 ( .A(ereg[560]), .B(n19486), .Z(n21726) );
  NANDN U28431 ( .A(n19481), .B(ereg[561]), .Z(n21725) );
  NAND U28432 ( .A(n21727), .B(n21728), .Z(n14815) );
  NANDN U28433 ( .A(init), .B(e[562]), .Z(n21728) );
  AND U28434 ( .A(n21729), .B(n21730), .Z(n21727) );
  NAND U28435 ( .A(ereg[561]), .B(n19486), .Z(n21730) );
  NANDN U28436 ( .A(n19481), .B(ereg[562]), .Z(n21729) );
  NAND U28437 ( .A(n21731), .B(n21732), .Z(n14814) );
  NANDN U28438 ( .A(init), .B(e[563]), .Z(n21732) );
  AND U28439 ( .A(n21733), .B(n21734), .Z(n21731) );
  NAND U28440 ( .A(ereg[562]), .B(n19486), .Z(n21734) );
  NANDN U28441 ( .A(n19481), .B(ereg[563]), .Z(n21733) );
  NAND U28442 ( .A(n21735), .B(n21736), .Z(n14813) );
  NANDN U28443 ( .A(init), .B(e[564]), .Z(n21736) );
  AND U28444 ( .A(n21737), .B(n21738), .Z(n21735) );
  NAND U28445 ( .A(ereg[563]), .B(n19486), .Z(n21738) );
  NANDN U28446 ( .A(n19481), .B(ereg[564]), .Z(n21737) );
  NAND U28447 ( .A(n21739), .B(n21740), .Z(n14812) );
  NANDN U28448 ( .A(init), .B(e[565]), .Z(n21740) );
  AND U28449 ( .A(n21741), .B(n21742), .Z(n21739) );
  NAND U28450 ( .A(ereg[564]), .B(n19486), .Z(n21742) );
  NANDN U28451 ( .A(n19481), .B(ereg[565]), .Z(n21741) );
  NAND U28452 ( .A(n21743), .B(n21744), .Z(n14811) );
  NANDN U28453 ( .A(init), .B(e[566]), .Z(n21744) );
  AND U28454 ( .A(n21745), .B(n21746), .Z(n21743) );
  NAND U28455 ( .A(ereg[565]), .B(n19486), .Z(n21746) );
  NANDN U28456 ( .A(n19481), .B(ereg[566]), .Z(n21745) );
  NAND U28457 ( .A(n21747), .B(n21748), .Z(n14810) );
  NANDN U28458 ( .A(init), .B(e[567]), .Z(n21748) );
  AND U28459 ( .A(n21749), .B(n21750), .Z(n21747) );
  NAND U28460 ( .A(ereg[566]), .B(n19486), .Z(n21750) );
  NANDN U28461 ( .A(n19481), .B(ereg[567]), .Z(n21749) );
  NAND U28462 ( .A(n21751), .B(n21752), .Z(n14809) );
  NANDN U28463 ( .A(init), .B(e[568]), .Z(n21752) );
  AND U28464 ( .A(n21753), .B(n21754), .Z(n21751) );
  NAND U28465 ( .A(ereg[567]), .B(n19486), .Z(n21754) );
  NANDN U28466 ( .A(n19481), .B(ereg[568]), .Z(n21753) );
  NAND U28467 ( .A(n21755), .B(n21756), .Z(n14808) );
  NANDN U28468 ( .A(init), .B(e[569]), .Z(n21756) );
  AND U28469 ( .A(n21757), .B(n21758), .Z(n21755) );
  NAND U28470 ( .A(ereg[568]), .B(n19486), .Z(n21758) );
  NANDN U28471 ( .A(n19481), .B(ereg[569]), .Z(n21757) );
  NAND U28472 ( .A(n21759), .B(n21760), .Z(n14807) );
  NANDN U28473 ( .A(init), .B(e[570]), .Z(n21760) );
  AND U28474 ( .A(n21761), .B(n21762), .Z(n21759) );
  NAND U28475 ( .A(ereg[569]), .B(n19486), .Z(n21762) );
  NANDN U28476 ( .A(n19481), .B(ereg[570]), .Z(n21761) );
  NAND U28477 ( .A(n21763), .B(n21764), .Z(n14806) );
  NANDN U28478 ( .A(init), .B(e[571]), .Z(n21764) );
  AND U28479 ( .A(n21765), .B(n21766), .Z(n21763) );
  NAND U28480 ( .A(ereg[570]), .B(n19486), .Z(n21766) );
  NANDN U28481 ( .A(n19481), .B(ereg[571]), .Z(n21765) );
  NAND U28482 ( .A(n21767), .B(n21768), .Z(n14805) );
  NANDN U28483 ( .A(init), .B(e[572]), .Z(n21768) );
  AND U28484 ( .A(n21769), .B(n21770), .Z(n21767) );
  NAND U28485 ( .A(ereg[571]), .B(n19486), .Z(n21770) );
  NANDN U28486 ( .A(n19481), .B(ereg[572]), .Z(n21769) );
  NAND U28487 ( .A(n21771), .B(n21772), .Z(n14804) );
  NANDN U28488 ( .A(init), .B(e[573]), .Z(n21772) );
  AND U28489 ( .A(n21773), .B(n21774), .Z(n21771) );
  NAND U28490 ( .A(ereg[572]), .B(n19486), .Z(n21774) );
  NANDN U28491 ( .A(n19481), .B(ereg[573]), .Z(n21773) );
  NAND U28492 ( .A(n21775), .B(n21776), .Z(n14803) );
  NANDN U28493 ( .A(init), .B(e[574]), .Z(n21776) );
  AND U28494 ( .A(n21777), .B(n21778), .Z(n21775) );
  NAND U28495 ( .A(ereg[573]), .B(n19486), .Z(n21778) );
  NANDN U28496 ( .A(n19481), .B(ereg[574]), .Z(n21777) );
  NAND U28497 ( .A(n21779), .B(n21780), .Z(n14802) );
  NANDN U28498 ( .A(init), .B(e[575]), .Z(n21780) );
  AND U28499 ( .A(n21781), .B(n21782), .Z(n21779) );
  NAND U28500 ( .A(ereg[574]), .B(n19486), .Z(n21782) );
  NANDN U28501 ( .A(n19481), .B(ereg[575]), .Z(n21781) );
  NAND U28502 ( .A(n21783), .B(n21784), .Z(n14801) );
  NANDN U28503 ( .A(init), .B(e[576]), .Z(n21784) );
  AND U28504 ( .A(n21785), .B(n21786), .Z(n21783) );
  NAND U28505 ( .A(ereg[575]), .B(n19486), .Z(n21786) );
  NANDN U28506 ( .A(n19481), .B(ereg[576]), .Z(n21785) );
  NAND U28507 ( .A(n21787), .B(n21788), .Z(n14800) );
  NANDN U28508 ( .A(init), .B(e[577]), .Z(n21788) );
  AND U28509 ( .A(n21789), .B(n21790), .Z(n21787) );
  NAND U28510 ( .A(ereg[576]), .B(n19486), .Z(n21790) );
  NANDN U28511 ( .A(n19481), .B(ereg[577]), .Z(n21789) );
  NAND U28512 ( .A(n21791), .B(n21792), .Z(n14799) );
  NANDN U28513 ( .A(init), .B(e[578]), .Z(n21792) );
  AND U28514 ( .A(n21793), .B(n21794), .Z(n21791) );
  NAND U28515 ( .A(ereg[577]), .B(n19486), .Z(n21794) );
  NANDN U28516 ( .A(n19481), .B(ereg[578]), .Z(n21793) );
  NAND U28517 ( .A(n21795), .B(n21796), .Z(n14798) );
  NANDN U28518 ( .A(init), .B(e[579]), .Z(n21796) );
  AND U28519 ( .A(n21797), .B(n21798), .Z(n21795) );
  NAND U28520 ( .A(ereg[578]), .B(n19486), .Z(n21798) );
  NANDN U28521 ( .A(n19481), .B(ereg[579]), .Z(n21797) );
  NAND U28522 ( .A(n21799), .B(n21800), .Z(n14797) );
  NANDN U28523 ( .A(init), .B(e[580]), .Z(n21800) );
  AND U28524 ( .A(n21801), .B(n21802), .Z(n21799) );
  NAND U28525 ( .A(ereg[579]), .B(n19486), .Z(n21802) );
  NANDN U28526 ( .A(n19481), .B(ereg[580]), .Z(n21801) );
  NAND U28527 ( .A(n21803), .B(n21804), .Z(n14796) );
  NANDN U28528 ( .A(init), .B(e[581]), .Z(n21804) );
  AND U28529 ( .A(n21805), .B(n21806), .Z(n21803) );
  NAND U28530 ( .A(ereg[580]), .B(n19486), .Z(n21806) );
  NANDN U28531 ( .A(n19481), .B(ereg[581]), .Z(n21805) );
  NAND U28532 ( .A(n21807), .B(n21808), .Z(n14795) );
  NANDN U28533 ( .A(init), .B(e[582]), .Z(n21808) );
  AND U28534 ( .A(n21809), .B(n21810), .Z(n21807) );
  NAND U28535 ( .A(ereg[581]), .B(n19486), .Z(n21810) );
  NANDN U28536 ( .A(n19481), .B(ereg[582]), .Z(n21809) );
  NAND U28537 ( .A(n21811), .B(n21812), .Z(n14794) );
  NANDN U28538 ( .A(init), .B(e[583]), .Z(n21812) );
  AND U28539 ( .A(n21813), .B(n21814), .Z(n21811) );
  NAND U28540 ( .A(ereg[582]), .B(n19486), .Z(n21814) );
  NANDN U28541 ( .A(n19481), .B(ereg[583]), .Z(n21813) );
  NAND U28542 ( .A(n21815), .B(n21816), .Z(n14793) );
  NANDN U28543 ( .A(init), .B(e[584]), .Z(n21816) );
  AND U28544 ( .A(n21817), .B(n21818), .Z(n21815) );
  NAND U28545 ( .A(ereg[583]), .B(n19486), .Z(n21818) );
  NANDN U28546 ( .A(n19481), .B(ereg[584]), .Z(n21817) );
  NAND U28547 ( .A(n21819), .B(n21820), .Z(n14792) );
  NANDN U28548 ( .A(init), .B(e[585]), .Z(n21820) );
  AND U28549 ( .A(n21821), .B(n21822), .Z(n21819) );
  NAND U28550 ( .A(ereg[584]), .B(n19486), .Z(n21822) );
  NANDN U28551 ( .A(n19481), .B(ereg[585]), .Z(n21821) );
  NAND U28552 ( .A(n21823), .B(n21824), .Z(n14791) );
  NANDN U28553 ( .A(init), .B(e[586]), .Z(n21824) );
  AND U28554 ( .A(n21825), .B(n21826), .Z(n21823) );
  NAND U28555 ( .A(ereg[585]), .B(n19486), .Z(n21826) );
  NANDN U28556 ( .A(n19481), .B(ereg[586]), .Z(n21825) );
  NAND U28557 ( .A(n21827), .B(n21828), .Z(n14790) );
  NANDN U28558 ( .A(init), .B(e[587]), .Z(n21828) );
  AND U28559 ( .A(n21829), .B(n21830), .Z(n21827) );
  NAND U28560 ( .A(ereg[586]), .B(n19486), .Z(n21830) );
  NANDN U28561 ( .A(n19481), .B(ereg[587]), .Z(n21829) );
  NAND U28562 ( .A(n21831), .B(n21832), .Z(n14789) );
  NANDN U28563 ( .A(init), .B(e[588]), .Z(n21832) );
  AND U28564 ( .A(n21833), .B(n21834), .Z(n21831) );
  NAND U28565 ( .A(ereg[587]), .B(n19486), .Z(n21834) );
  NANDN U28566 ( .A(n19481), .B(ereg[588]), .Z(n21833) );
  NAND U28567 ( .A(n21835), .B(n21836), .Z(n14788) );
  NANDN U28568 ( .A(init), .B(e[589]), .Z(n21836) );
  AND U28569 ( .A(n21837), .B(n21838), .Z(n21835) );
  NAND U28570 ( .A(ereg[588]), .B(n19486), .Z(n21838) );
  NANDN U28571 ( .A(n19481), .B(ereg[589]), .Z(n21837) );
  NAND U28572 ( .A(n21839), .B(n21840), .Z(n14787) );
  NANDN U28573 ( .A(init), .B(e[590]), .Z(n21840) );
  AND U28574 ( .A(n21841), .B(n21842), .Z(n21839) );
  NAND U28575 ( .A(ereg[589]), .B(n19486), .Z(n21842) );
  NANDN U28576 ( .A(n19481), .B(ereg[590]), .Z(n21841) );
  NAND U28577 ( .A(n21843), .B(n21844), .Z(n14786) );
  NANDN U28578 ( .A(init), .B(e[591]), .Z(n21844) );
  AND U28579 ( .A(n21845), .B(n21846), .Z(n21843) );
  NAND U28580 ( .A(ereg[590]), .B(n19486), .Z(n21846) );
  NANDN U28581 ( .A(n19481), .B(ereg[591]), .Z(n21845) );
  NAND U28582 ( .A(n21847), .B(n21848), .Z(n14785) );
  NANDN U28583 ( .A(init), .B(e[592]), .Z(n21848) );
  AND U28584 ( .A(n21849), .B(n21850), .Z(n21847) );
  NAND U28585 ( .A(ereg[591]), .B(n19486), .Z(n21850) );
  NANDN U28586 ( .A(n19481), .B(ereg[592]), .Z(n21849) );
  NAND U28587 ( .A(n21851), .B(n21852), .Z(n14784) );
  NANDN U28588 ( .A(init), .B(e[593]), .Z(n21852) );
  AND U28589 ( .A(n21853), .B(n21854), .Z(n21851) );
  NAND U28590 ( .A(ereg[592]), .B(n19486), .Z(n21854) );
  NANDN U28591 ( .A(n19481), .B(ereg[593]), .Z(n21853) );
  NAND U28592 ( .A(n21855), .B(n21856), .Z(n14783) );
  NANDN U28593 ( .A(init), .B(e[594]), .Z(n21856) );
  AND U28594 ( .A(n21857), .B(n21858), .Z(n21855) );
  NAND U28595 ( .A(ereg[593]), .B(n19486), .Z(n21858) );
  NANDN U28596 ( .A(n19481), .B(ereg[594]), .Z(n21857) );
  NAND U28597 ( .A(n21859), .B(n21860), .Z(n14782) );
  NANDN U28598 ( .A(init), .B(e[595]), .Z(n21860) );
  AND U28599 ( .A(n21861), .B(n21862), .Z(n21859) );
  NAND U28600 ( .A(ereg[594]), .B(n19486), .Z(n21862) );
  NANDN U28601 ( .A(n19481), .B(ereg[595]), .Z(n21861) );
  NAND U28602 ( .A(n21863), .B(n21864), .Z(n14781) );
  NANDN U28603 ( .A(init), .B(e[596]), .Z(n21864) );
  AND U28604 ( .A(n21865), .B(n21866), .Z(n21863) );
  NAND U28605 ( .A(ereg[595]), .B(n19486), .Z(n21866) );
  NANDN U28606 ( .A(n19481), .B(ereg[596]), .Z(n21865) );
  NAND U28607 ( .A(n21867), .B(n21868), .Z(n14780) );
  NANDN U28608 ( .A(init), .B(e[597]), .Z(n21868) );
  AND U28609 ( .A(n21869), .B(n21870), .Z(n21867) );
  NAND U28610 ( .A(ereg[596]), .B(n19486), .Z(n21870) );
  NANDN U28611 ( .A(n19481), .B(ereg[597]), .Z(n21869) );
  NAND U28612 ( .A(n21871), .B(n21872), .Z(n14779) );
  NANDN U28613 ( .A(init), .B(e[598]), .Z(n21872) );
  AND U28614 ( .A(n21873), .B(n21874), .Z(n21871) );
  NAND U28615 ( .A(ereg[597]), .B(n19486), .Z(n21874) );
  NANDN U28616 ( .A(n19481), .B(ereg[598]), .Z(n21873) );
  NAND U28617 ( .A(n21875), .B(n21876), .Z(n14778) );
  NANDN U28618 ( .A(init), .B(e[599]), .Z(n21876) );
  AND U28619 ( .A(n21877), .B(n21878), .Z(n21875) );
  NAND U28620 ( .A(ereg[598]), .B(n19486), .Z(n21878) );
  NANDN U28621 ( .A(n19481), .B(ereg[599]), .Z(n21877) );
  NAND U28622 ( .A(n21879), .B(n21880), .Z(n14777) );
  NANDN U28623 ( .A(init), .B(e[600]), .Z(n21880) );
  AND U28624 ( .A(n21881), .B(n21882), .Z(n21879) );
  NAND U28625 ( .A(ereg[599]), .B(n19486), .Z(n21882) );
  NANDN U28626 ( .A(n19481), .B(ereg[600]), .Z(n21881) );
  NAND U28627 ( .A(n21883), .B(n21884), .Z(n14776) );
  NANDN U28628 ( .A(init), .B(e[601]), .Z(n21884) );
  AND U28629 ( .A(n21885), .B(n21886), .Z(n21883) );
  NAND U28630 ( .A(ereg[600]), .B(n19486), .Z(n21886) );
  NANDN U28631 ( .A(n19481), .B(ereg[601]), .Z(n21885) );
  NAND U28632 ( .A(n21887), .B(n21888), .Z(n14775) );
  NANDN U28633 ( .A(init), .B(e[602]), .Z(n21888) );
  AND U28634 ( .A(n21889), .B(n21890), .Z(n21887) );
  NAND U28635 ( .A(ereg[601]), .B(n19486), .Z(n21890) );
  NANDN U28636 ( .A(n19481), .B(ereg[602]), .Z(n21889) );
  NAND U28637 ( .A(n21891), .B(n21892), .Z(n14774) );
  NANDN U28638 ( .A(init), .B(e[603]), .Z(n21892) );
  AND U28639 ( .A(n21893), .B(n21894), .Z(n21891) );
  NAND U28640 ( .A(ereg[602]), .B(n19486), .Z(n21894) );
  NANDN U28641 ( .A(n19481), .B(ereg[603]), .Z(n21893) );
  NAND U28642 ( .A(n21895), .B(n21896), .Z(n14773) );
  NANDN U28643 ( .A(init), .B(e[604]), .Z(n21896) );
  AND U28644 ( .A(n21897), .B(n21898), .Z(n21895) );
  NAND U28645 ( .A(ereg[603]), .B(n19486), .Z(n21898) );
  NANDN U28646 ( .A(n19481), .B(ereg[604]), .Z(n21897) );
  NAND U28647 ( .A(n21899), .B(n21900), .Z(n14772) );
  NANDN U28648 ( .A(init), .B(e[605]), .Z(n21900) );
  AND U28649 ( .A(n21901), .B(n21902), .Z(n21899) );
  NAND U28650 ( .A(ereg[604]), .B(n19486), .Z(n21902) );
  NANDN U28651 ( .A(n19481), .B(ereg[605]), .Z(n21901) );
  NAND U28652 ( .A(n21903), .B(n21904), .Z(n14771) );
  NANDN U28653 ( .A(init), .B(e[606]), .Z(n21904) );
  AND U28654 ( .A(n21905), .B(n21906), .Z(n21903) );
  NAND U28655 ( .A(ereg[605]), .B(n19486), .Z(n21906) );
  NANDN U28656 ( .A(n19481), .B(ereg[606]), .Z(n21905) );
  NAND U28657 ( .A(n21907), .B(n21908), .Z(n14770) );
  NANDN U28658 ( .A(init), .B(e[607]), .Z(n21908) );
  AND U28659 ( .A(n21909), .B(n21910), .Z(n21907) );
  NAND U28660 ( .A(ereg[606]), .B(n19486), .Z(n21910) );
  NANDN U28661 ( .A(n19481), .B(ereg[607]), .Z(n21909) );
  NAND U28662 ( .A(n21911), .B(n21912), .Z(n14769) );
  NANDN U28663 ( .A(init), .B(e[608]), .Z(n21912) );
  AND U28664 ( .A(n21913), .B(n21914), .Z(n21911) );
  NAND U28665 ( .A(ereg[607]), .B(n19486), .Z(n21914) );
  NANDN U28666 ( .A(n19481), .B(ereg[608]), .Z(n21913) );
  NAND U28667 ( .A(n21915), .B(n21916), .Z(n14768) );
  NANDN U28668 ( .A(init), .B(e[609]), .Z(n21916) );
  AND U28669 ( .A(n21917), .B(n21918), .Z(n21915) );
  NAND U28670 ( .A(ereg[608]), .B(n19486), .Z(n21918) );
  NANDN U28671 ( .A(n19481), .B(ereg[609]), .Z(n21917) );
  NAND U28672 ( .A(n21919), .B(n21920), .Z(n14767) );
  NANDN U28673 ( .A(init), .B(e[610]), .Z(n21920) );
  AND U28674 ( .A(n21921), .B(n21922), .Z(n21919) );
  NAND U28675 ( .A(ereg[609]), .B(n19486), .Z(n21922) );
  NANDN U28676 ( .A(n19481), .B(ereg[610]), .Z(n21921) );
  NAND U28677 ( .A(n21923), .B(n21924), .Z(n14766) );
  NANDN U28678 ( .A(init), .B(e[611]), .Z(n21924) );
  AND U28679 ( .A(n21925), .B(n21926), .Z(n21923) );
  NAND U28680 ( .A(ereg[610]), .B(n19486), .Z(n21926) );
  NANDN U28681 ( .A(n19481), .B(ereg[611]), .Z(n21925) );
  NAND U28682 ( .A(n21927), .B(n21928), .Z(n14765) );
  NANDN U28683 ( .A(init), .B(e[612]), .Z(n21928) );
  AND U28684 ( .A(n21929), .B(n21930), .Z(n21927) );
  NAND U28685 ( .A(ereg[611]), .B(n19486), .Z(n21930) );
  NANDN U28686 ( .A(n19481), .B(ereg[612]), .Z(n21929) );
  NAND U28687 ( .A(n21931), .B(n21932), .Z(n14764) );
  NANDN U28688 ( .A(init), .B(e[613]), .Z(n21932) );
  AND U28689 ( .A(n21933), .B(n21934), .Z(n21931) );
  NAND U28690 ( .A(ereg[612]), .B(n19486), .Z(n21934) );
  NANDN U28691 ( .A(n19481), .B(ereg[613]), .Z(n21933) );
  NAND U28692 ( .A(n21935), .B(n21936), .Z(n14763) );
  NANDN U28693 ( .A(init), .B(e[614]), .Z(n21936) );
  AND U28694 ( .A(n21937), .B(n21938), .Z(n21935) );
  NAND U28695 ( .A(ereg[613]), .B(n19486), .Z(n21938) );
  NANDN U28696 ( .A(n19481), .B(ereg[614]), .Z(n21937) );
  NAND U28697 ( .A(n21939), .B(n21940), .Z(n14762) );
  NANDN U28698 ( .A(init), .B(e[615]), .Z(n21940) );
  AND U28699 ( .A(n21941), .B(n21942), .Z(n21939) );
  NAND U28700 ( .A(ereg[614]), .B(n19486), .Z(n21942) );
  NANDN U28701 ( .A(n19481), .B(ereg[615]), .Z(n21941) );
  NAND U28702 ( .A(n21943), .B(n21944), .Z(n14761) );
  NANDN U28703 ( .A(init), .B(e[616]), .Z(n21944) );
  AND U28704 ( .A(n21945), .B(n21946), .Z(n21943) );
  NAND U28705 ( .A(ereg[615]), .B(n19486), .Z(n21946) );
  NANDN U28706 ( .A(n19481), .B(ereg[616]), .Z(n21945) );
  NAND U28707 ( .A(n21947), .B(n21948), .Z(n14760) );
  NANDN U28708 ( .A(init), .B(e[617]), .Z(n21948) );
  AND U28709 ( .A(n21949), .B(n21950), .Z(n21947) );
  NAND U28710 ( .A(ereg[616]), .B(n19486), .Z(n21950) );
  NANDN U28711 ( .A(n19481), .B(ereg[617]), .Z(n21949) );
  NAND U28712 ( .A(n21951), .B(n21952), .Z(n14759) );
  NANDN U28713 ( .A(init), .B(e[618]), .Z(n21952) );
  AND U28714 ( .A(n21953), .B(n21954), .Z(n21951) );
  NAND U28715 ( .A(ereg[617]), .B(n19486), .Z(n21954) );
  NANDN U28716 ( .A(n19481), .B(ereg[618]), .Z(n21953) );
  NAND U28717 ( .A(n21955), .B(n21956), .Z(n14758) );
  NANDN U28718 ( .A(init), .B(e[619]), .Z(n21956) );
  AND U28719 ( .A(n21957), .B(n21958), .Z(n21955) );
  NAND U28720 ( .A(ereg[618]), .B(n19486), .Z(n21958) );
  NANDN U28721 ( .A(n19481), .B(ereg[619]), .Z(n21957) );
  NAND U28722 ( .A(n21959), .B(n21960), .Z(n14757) );
  NANDN U28723 ( .A(init), .B(e[620]), .Z(n21960) );
  AND U28724 ( .A(n21961), .B(n21962), .Z(n21959) );
  NAND U28725 ( .A(ereg[619]), .B(n19486), .Z(n21962) );
  NANDN U28726 ( .A(n19481), .B(ereg[620]), .Z(n21961) );
  NAND U28727 ( .A(n21963), .B(n21964), .Z(n14756) );
  NANDN U28728 ( .A(init), .B(e[621]), .Z(n21964) );
  AND U28729 ( .A(n21965), .B(n21966), .Z(n21963) );
  NAND U28730 ( .A(ereg[620]), .B(n19486), .Z(n21966) );
  NANDN U28731 ( .A(n19481), .B(ereg[621]), .Z(n21965) );
  NAND U28732 ( .A(n21967), .B(n21968), .Z(n14755) );
  NANDN U28733 ( .A(init), .B(e[622]), .Z(n21968) );
  AND U28734 ( .A(n21969), .B(n21970), .Z(n21967) );
  NAND U28735 ( .A(ereg[621]), .B(n19486), .Z(n21970) );
  NANDN U28736 ( .A(n19481), .B(ereg[622]), .Z(n21969) );
  NAND U28737 ( .A(n21971), .B(n21972), .Z(n14754) );
  NANDN U28738 ( .A(init), .B(e[623]), .Z(n21972) );
  AND U28739 ( .A(n21973), .B(n21974), .Z(n21971) );
  NAND U28740 ( .A(ereg[622]), .B(n19486), .Z(n21974) );
  NANDN U28741 ( .A(n19481), .B(ereg[623]), .Z(n21973) );
  NAND U28742 ( .A(n21975), .B(n21976), .Z(n14753) );
  NANDN U28743 ( .A(init), .B(e[624]), .Z(n21976) );
  AND U28744 ( .A(n21977), .B(n21978), .Z(n21975) );
  NAND U28745 ( .A(ereg[623]), .B(n19486), .Z(n21978) );
  NANDN U28746 ( .A(n19481), .B(ereg[624]), .Z(n21977) );
  NAND U28747 ( .A(n21979), .B(n21980), .Z(n14752) );
  NANDN U28748 ( .A(init), .B(e[625]), .Z(n21980) );
  AND U28749 ( .A(n21981), .B(n21982), .Z(n21979) );
  NAND U28750 ( .A(ereg[624]), .B(n19486), .Z(n21982) );
  NANDN U28751 ( .A(n19481), .B(ereg[625]), .Z(n21981) );
  NAND U28752 ( .A(n21983), .B(n21984), .Z(n14751) );
  NANDN U28753 ( .A(init), .B(e[626]), .Z(n21984) );
  AND U28754 ( .A(n21985), .B(n21986), .Z(n21983) );
  NAND U28755 ( .A(ereg[625]), .B(n19486), .Z(n21986) );
  NANDN U28756 ( .A(n19481), .B(ereg[626]), .Z(n21985) );
  NAND U28757 ( .A(n21987), .B(n21988), .Z(n14750) );
  NANDN U28758 ( .A(init), .B(e[627]), .Z(n21988) );
  AND U28759 ( .A(n21989), .B(n21990), .Z(n21987) );
  NAND U28760 ( .A(ereg[626]), .B(n19486), .Z(n21990) );
  NANDN U28761 ( .A(n19481), .B(ereg[627]), .Z(n21989) );
  NAND U28762 ( .A(n21991), .B(n21992), .Z(n14749) );
  NANDN U28763 ( .A(init), .B(e[628]), .Z(n21992) );
  AND U28764 ( .A(n21993), .B(n21994), .Z(n21991) );
  NAND U28765 ( .A(ereg[627]), .B(n19486), .Z(n21994) );
  NANDN U28766 ( .A(n19481), .B(ereg[628]), .Z(n21993) );
  NAND U28767 ( .A(n21995), .B(n21996), .Z(n14748) );
  NANDN U28768 ( .A(init), .B(e[629]), .Z(n21996) );
  AND U28769 ( .A(n21997), .B(n21998), .Z(n21995) );
  NAND U28770 ( .A(ereg[628]), .B(n19486), .Z(n21998) );
  NANDN U28771 ( .A(n19481), .B(ereg[629]), .Z(n21997) );
  NAND U28772 ( .A(n21999), .B(n22000), .Z(n14747) );
  NANDN U28773 ( .A(init), .B(e[630]), .Z(n22000) );
  AND U28774 ( .A(n22001), .B(n22002), .Z(n21999) );
  NAND U28775 ( .A(ereg[629]), .B(n19486), .Z(n22002) );
  NANDN U28776 ( .A(n19481), .B(ereg[630]), .Z(n22001) );
  NAND U28777 ( .A(n22003), .B(n22004), .Z(n14746) );
  NANDN U28778 ( .A(init), .B(e[631]), .Z(n22004) );
  AND U28779 ( .A(n22005), .B(n22006), .Z(n22003) );
  NAND U28780 ( .A(ereg[630]), .B(n19486), .Z(n22006) );
  NANDN U28781 ( .A(n19481), .B(ereg[631]), .Z(n22005) );
  NAND U28782 ( .A(n22007), .B(n22008), .Z(n14745) );
  NANDN U28783 ( .A(init), .B(e[632]), .Z(n22008) );
  AND U28784 ( .A(n22009), .B(n22010), .Z(n22007) );
  NAND U28785 ( .A(ereg[631]), .B(n19486), .Z(n22010) );
  NANDN U28786 ( .A(n19481), .B(ereg[632]), .Z(n22009) );
  NAND U28787 ( .A(n22011), .B(n22012), .Z(n14744) );
  NANDN U28788 ( .A(init), .B(e[633]), .Z(n22012) );
  AND U28789 ( .A(n22013), .B(n22014), .Z(n22011) );
  NAND U28790 ( .A(ereg[632]), .B(n19486), .Z(n22014) );
  NANDN U28791 ( .A(n19481), .B(ereg[633]), .Z(n22013) );
  NAND U28792 ( .A(n22015), .B(n22016), .Z(n14743) );
  NANDN U28793 ( .A(init), .B(e[634]), .Z(n22016) );
  AND U28794 ( .A(n22017), .B(n22018), .Z(n22015) );
  NAND U28795 ( .A(ereg[633]), .B(n19486), .Z(n22018) );
  NANDN U28796 ( .A(n19481), .B(ereg[634]), .Z(n22017) );
  NAND U28797 ( .A(n22019), .B(n22020), .Z(n14742) );
  NANDN U28798 ( .A(init), .B(e[635]), .Z(n22020) );
  AND U28799 ( .A(n22021), .B(n22022), .Z(n22019) );
  NAND U28800 ( .A(ereg[634]), .B(n19486), .Z(n22022) );
  NANDN U28801 ( .A(n19481), .B(ereg[635]), .Z(n22021) );
  NAND U28802 ( .A(n22023), .B(n22024), .Z(n14741) );
  NANDN U28803 ( .A(init), .B(e[636]), .Z(n22024) );
  AND U28804 ( .A(n22025), .B(n22026), .Z(n22023) );
  NAND U28805 ( .A(ereg[635]), .B(n19486), .Z(n22026) );
  NANDN U28806 ( .A(n19481), .B(ereg[636]), .Z(n22025) );
  NAND U28807 ( .A(n22027), .B(n22028), .Z(n14740) );
  NANDN U28808 ( .A(init), .B(e[637]), .Z(n22028) );
  AND U28809 ( .A(n22029), .B(n22030), .Z(n22027) );
  NAND U28810 ( .A(ereg[636]), .B(n19486), .Z(n22030) );
  NANDN U28811 ( .A(n19481), .B(ereg[637]), .Z(n22029) );
  NAND U28812 ( .A(n22031), .B(n22032), .Z(n14739) );
  NANDN U28813 ( .A(init), .B(e[638]), .Z(n22032) );
  AND U28814 ( .A(n22033), .B(n22034), .Z(n22031) );
  NAND U28815 ( .A(ereg[637]), .B(n19486), .Z(n22034) );
  NANDN U28816 ( .A(n19481), .B(ereg[638]), .Z(n22033) );
  NAND U28817 ( .A(n22035), .B(n22036), .Z(n14738) );
  NANDN U28818 ( .A(init), .B(e[639]), .Z(n22036) );
  AND U28819 ( .A(n22037), .B(n22038), .Z(n22035) );
  NAND U28820 ( .A(ereg[638]), .B(n19486), .Z(n22038) );
  NANDN U28821 ( .A(n19481), .B(ereg[639]), .Z(n22037) );
  NAND U28822 ( .A(n22039), .B(n22040), .Z(n14737) );
  NANDN U28823 ( .A(init), .B(e[640]), .Z(n22040) );
  AND U28824 ( .A(n22041), .B(n22042), .Z(n22039) );
  NAND U28825 ( .A(ereg[639]), .B(n19486), .Z(n22042) );
  NANDN U28826 ( .A(n19481), .B(ereg[640]), .Z(n22041) );
  NAND U28827 ( .A(n22043), .B(n22044), .Z(n14736) );
  NANDN U28828 ( .A(init), .B(e[641]), .Z(n22044) );
  AND U28829 ( .A(n22045), .B(n22046), .Z(n22043) );
  NAND U28830 ( .A(ereg[640]), .B(n19486), .Z(n22046) );
  NANDN U28831 ( .A(n19481), .B(ereg[641]), .Z(n22045) );
  NAND U28832 ( .A(n22047), .B(n22048), .Z(n14735) );
  NANDN U28833 ( .A(init), .B(e[642]), .Z(n22048) );
  AND U28834 ( .A(n22049), .B(n22050), .Z(n22047) );
  NAND U28835 ( .A(ereg[641]), .B(n19486), .Z(n22050) );
  NANDN U28836 ( .A(n19481), .B(ereg[642]), .Z(n22049) );
  NAND U28837 ( .A(n22051), .B(n22052), .Z(n14734) );
  NANDN U28838 ( .A(init), .B(e[643]), .Z(n22052) );
  AND U28839 ( .A(n22053), .B(n22054), .Z(n22051) );
  NAND U28840 ( .A(ereg[642]), .B(n19486), .Z(n22054) );
  NANDN U28841 ( .A(n19481), .B(ereg[643]), .Z(n22053) );
  NAND U28842 ( .A(n22055), .B(n22056), .Z(n14733) );
  NANDN U28843 ( .A(init), .B(e[644]), .Z(n22056) );
  AND U28844 ( .A(n22057), .B(n22058), .Z(n22055) );
  NAND U28845 ( .A(ereg[643]), .B(n19486), .Z(n22058) );
  NANDN U28846 ( .A(n19481), .B(ereg[644]), .Z(n22057) );
  NAND U28847 ( .A(n22059), .B(n22060), .Z(n14732) );
  NANDN U28848 ( .A(init), .B(e[645]), .Z(n22060) );
  AND U28849 ( .A(n22061), .B(n22062), .Z(n22059) );
  NAND U28850 ( .A(ereg[644]), .B(n19486), .Z(n22062) );
  NANDN U28851 ( .A(n19481), .B(ereg[645]), .Z(n22061) );
  NAND U28852 ( .A(n22063), .B(n22064), .Z(n14731) );
  NANDN U28853 ( .A(init), .B(e[646]), .Z(n22064) );
  AND U28854 ( .A(n22065), .B(n22066), .Z(n22063) );
  NAND U28855 ( .A(ereg[645]), .B(n19486), .Z(n22066) );
  NANDN U28856 ( .A(n19481), .B(ereg[646]), .Z(n22065) );
  NAND U28857 ( .A(n22067), .B(n22068), .Z(n14730) );
  NANDN U28858 ( .A(init), .B(e[647]), .Z(n22068) );
  AND U28859 ( .A(n22069), .B(n22070), .Z(n22067) );
  NAND U28860 ( .A(ereg[646]), .B(n19486), .Z(n22070) );
  NANDN U28861 ( .A(n19481), .B(ereg[647]), .Z(n22069) );
  NAND U28862 ( .A(n22071), .B(n22072), .Z(n14729) );
  NANDN U28863 ( .A(init), .B(e[648]), .Z(n22072) );
  AND U28864 ( .A(n22073), .B(n22074), .Z(n22071) );
  NAND U28865 ( .A(ereg[647]), .B(n19486), .Z(n22074) );
  NANDN U28866 ( .A(n19481), .B(ereg[648]), .Z(n22073) );
  NAND U28867 ( .A(n22075), .B(n22076), .Z(n14728) );
  NANDN U28868 ( .A(init), .B(e[649]), .Z(n22076) );
  AND U28869 ( .A(n22077), .B(n22078), .Z(n22075) );
  NAND U28870 ( .A(ereg[648]), .B(n19486), .Z(n22078) );
  NANDN U28871 ( .A(n19481), .B(ereg[649]), .Z(n22077) );
  NAND U28872 ( .A(n22079), .B(n22080), .Z(n14727) );
  NANDN U28873 ( .A(init), .B(e[650]), .Z(n22080) );
  AND U28874 ( .A(n22081), .B(n22082), .Z(n22079) );
  NAND U28875 ( .A(ereg[649]), .B(n19486), .Z(n22082) );
  NANDN U28876 ( .A(n19481), .B(ereg[650]), .Z(n22081) );
  NAND U28877 ( .A(n22083), .B(n22084), .Z(n14726) );
  NANDN U28878 ( .A(init), .B(e[651]), .Z(n22084) );
  AND U28879 ( .A(n22085), .B(n22086), .Z(n22083) );
  NAND U28880 ( .A(ereg[650]), .B(n19486), .Z(n22086) );
  NANDN U28881 ( .A(n19481), .B(ereg[651]), .Z(n22085) );
  NAND U28882 ( .A(n22087), .B(n22088), .Z(n14725) );
  NANDN U28883 ( .A(init), .B(e[652]), .Z(n22088) );
  AND U28884 ( .A(n22089), .B(n22090), .Z(n22087) );
  NAND U28885 ( .A(ereg[651]), .B(n19486), .Z(n22090) );
  NANDN U28886 ( .A(n19481), .B(ereg[652]), .Z(n22089) );
  NAND U28887 ( .A(n22091), .B(n22092), .Z(n14724) );
  NANDN U28888 ( .A(init), .B(e[653]), .Z(n22092) );
  AND U28889 ( .A(n22093), .B(n22094), .Z(n22091) );
  NAND U28890 ( .A(ereg[652]), .B(n19486), .Z(n22094) );
  NANDN U28891 ( .A(n19481), .B(ereg[653]), .Z(n22093) );
  NAND U28892 ( .A(n22095), .B(n22096), .Z(n14723) );
  NANDN U28893 ( .A(init), .B(e[654]), .Z(n22096) );
  AND U28894 ( .A(n22097), .B(n22098), .Z(n22095) );
  NAND U28895 ( .A(ereg[653]), .B(n19486), .Z(n22098) );
  NANDN U28896 ( .A(n19481), .B(ereg[654]), .Z(n22097) );
  NAND U28897 ( .A(n22099), .B(n22100), .Z(n14722) );
  NANDN U28898 ( .A(init), .B(e[655]), .Z(n22100) );
  AND U28899 ( .A(n22101), .B(n22102), .Z(n22099) );
  NAND U28900 ( .A(ereg[654]), .B(n19486), .Z(n22102) );
  NANDN U28901 ( .A(n19481), .B(ereg[655]), .Z(n22101) );
  NAND U28902 ( .A(n22103), .B(n22104), .Z(n14721) );
  NANDN U28903 ( .A(init), .B(e[656]), .Z(n22104) );
  AND U28904 ( .A(n22105), .B(n22106), .Z(n22103) );
  NAND U28905 ( .A(ereg[655]), .B(n19486), .Z(n22106) );
  NANDN U28906 ( .A(n19481), .B(ereg[656]), .Z(n22105) );
  NAND U28907 ( .A(n22107), .B(n22108), .Z(n14720) );
  NANDN U28908 ( .A(init), .B(e[657]), .Z(n22108) );
  AND U28909 ( .A(n22109), .B(n22110), .Z(n22107) );
  NAND U28910 ( .A(ereg[656]), .B(n19486), .Z(n22110) );
  NANDN U28911 ( .A(n19481), .B(ereg[657]), .Z(n22109) );
  NAND U28912 ( .A(n22111), .B(n22112), .Z(n14719) );
  NANDN U28913 ( .A(init), .B(e[658]), .Z(n22112) );
  AND U28914 ( .A(n22113), .B(n22114), .Z(n22111) );
  NAND U28915 ( .A(ereg[657]), .B(n19486), .Z(n22114) );
  NANDN U28916 ( .A(n19481), .B(ereg[658]), .Z(n22113) );
  NAND U28917 ( .A(n22115), .B(n22116), .Z(n14718) );
  NANDN U28918 ( .A(init), .B(e[659]), .Z(n22116) );
  AND U28919 ( .A(n22117), .B(n22118), .Z(n22115) );
  NAND U28920 ( .A(ereg[658]), .B(n19486), .Z(n22118) );
  NANDN U28921 ( .A(n19481), .B(ereg[659]), .Z(n22117) );
  NAND U28922 ( .A(n22119), .B(n22120), .Z(n14717) );
  NANDN U28923 ( .A(init), .B(e[660]), .Z(n22120) );
  AND U28924 ( .A(n22121), .B(n22122), .Z(n22119) );
  NAND U28925 ( .A(ereg[659]), .B(n19486), .Z(n22122) );
  NANDN U28926 ( .A(n19481), .B(ereg[660]), .Z(n22121) );
  NAND U28927 ( .A(n22123), .B(n22124), .Z(n14716) );
  NANDN U28928 ( .A(init), .B(e[661]), .Z(n22124) );
  AND U28929 ( .A(n22125), .B(n22126), .Z(n22123) );
  NAND U28930 ( .A(ereg[660]), .B(n19486), .Z(n22126) );
  NANDN U28931 ( .A(n19481), .B(ereg[661]), .Z(n22125) );
  NAND U28932 ( .A(n22127), .B(n22128), .Z(n14715) );
  NANDN U28933 ( .A(init), .B(e[662]), .Z(n22128) );
  AND U28934 ( .A(n22129), .B(n22130), .Z(n22127) );
  NAND U28935 ( .A(ereg[661]), .B(n19486), .Z(n22130) );
  NANDN U28936 ( .A(n19481), .B(ereg[662]), .Z(n22129) );
  NAND U28937 ( .A(n22131), .B(n22132), .Z(n14714) );
  NANDN U28938 ( .A(init), .B(e[663]), .Z(n22132) );
  AND U28939 ( .A(n22133), .B(n22134), .Z(n22131) );
  NAND U28940 ( .A(ereg[662]), .B(n19486), .Z(n22134) );
  NANDN U28941 ( .A(n19481), .B(ereg[663]), .Z(n22133) );
  NAND U28942 ( .A(n22135), .B(n22136), .Z(n14713) );
  NANDN U28943 ( .A(init), .B(e[664]), .Z(n22136) );
  AND U28944 ( .A(n22137), .B(n22138), .Z(n22135) );
  NAND U28945 ( .A(ereg[663]), .B(n19486), .Z(n22138) );
  NANDN U28946 ( .A(n19481), .B(ereg[664]), .Z(n22137) );
  NAND U28947 ( .A(n22139), .B(n22140), .Z(n14712) );
  NANDN U28948 ( .A(init), .B(e[665]), .Z(n22140) );
  AND U28949 ( .A(n22141), .B(n22142), .Z(n22139) );
  NAND U28950 ( .A(ereg[664]), .B(n19486), .Z(n22142) );
  NANDN U28951 ( .A(n19481), .B(ereg[665]), .Z(n22141) );
  NAND U28952 ( .A(n22143), .B(n22144), .Z(n14711) );
  NANDN U28953 ( .A(init), .B(e[666]), .Z(n22144) );
  AND U28954 ( .A(n22145), .B(n22146), .Z(n22143) );
  NAND U28955 ( .A(ereg[665]), .B(n19486), .Z(n22146) );
  NANDN U28956 ( .A(n19481), .B(ereg[666]), .Z(n22145) );
  NAND U28957 ( .A(n22147), .B(n22148), .Z(n14710) );
  NANDN U28958 ( .A(init), .B(e[667]), .Z(n22148) );
  AND U28959 ( .A(n22149), .B(n22150), .Z(n22147) );
  NAND U28960 ( .A(ereg[666]), .B(n19486), .Z(n22150) );
  NANDN U28961 ( .A(n19481), .B(ereg[667]), .Z(n22149) );
  NAND U28962 ( .A(n22151), .B(n22152), .Z(n14709) );
  NANDN U28963 ( .A(init), .B(e[668]), .Z(n22152) );
  AND U28964 ( .A(n22153), .B(n22154), .Z(n22151) );
  NAND U28965 ( .A(ereg[667]), .B(n19486), .Z(n22154) );
  NANDN U28966 ( .A(n19481), .B(ereg[668]), .Z(n22153) );
  NAND U28967 ( .A(n22155), .B(n22156), .Z(n14708) );
  NANDN U28968 ( .A(init), .B(e[669]), .Z(n22156) );
  AND U28969 ( .A(n22157), .B(n22158), .Z(n22155) );
  NAND U28970 ( .A(ereg[668]), .B(n19486), .Z(n22158) );
  NANDN U28971 ( .A(n19481), .B(ereg[669]), .Z(n22157) );
  NAND U28972 ( .A(n22159), .B(n22160), .Z(n14707) );
  NANDN U28973 ( .A(init), .B(e[670]), .Z(n22160) );
  AND U28974 ( .A(n22161), .B(n22162), .Z(n22159) );
  NAND U28975 ( .A(ereg[669]), .B(n19486), .Z(n22162) );
  NANDN U28976 ( .A(n19481), .B(ereg[670]), .Z(n22161) );
  NAND U28977 ( .A(n22163), .B(n22164), .Z(n14706) );
  NANDN U28978 ( .A(init), .B(e[671]), .Z(n22164) );
  AND U28979 ( .A(n22165), .B(n22166), .Z(n22163) );
  NAND U28980 ( .A(ereg[670]), .B(n19486), .Z(n22166) );
  NANDN U28981 ( .A(n19481), .B(ereg[671]), .Z(n22165) );
  NAND U28982 ( .A(n22167), .B(n22168), .Z(n14705) );
  NANDN U28983 ( .A(init), .B(e[672]), .Z(n22168) );
  AND U28984 ( .A(n22169), .B(n22170), .Z(n22167) );
  NAND U28985 ( .A(ereg[671]), .B(n19486), .Z(n22170) );
  NANDN U28986 ( .A(n19481), .B(ereg[672]), .Z(n22169) );
  NAND U28987 ( .A(n22171), .B(n22172), .Z(n14704) );
  NANDN U28988 ( .A(init), .B(e[673]), .Z(n22172) );
  AND U28989 ( .A(n22173), .B(n22174), .Z(n22171) );
  NAND U28990 ( .A(ereg[672]), .B(n19486), .Z(n22174) );
  NANDN U28991 ( .A(n19481), .B(ereg[673]), .Z(n22173) );
  NAND U28992 ( .A(n22175), .B(n22176), .Z(n14703) );
  NANDN U28993 ( .A(init), .B(e[674]), .Z(n22176) );
  AND U28994 ( .A(n22177), .B(n22178), .Z(n22175) );
  NAND U28995 ( .A(ereg[673]), .B(n19486), .Z(n22178) );
  NANDN U28996 ( .A(n19481), .B(ereg[674]), .Z(n22177) );
  NAND U28997 ( .A(n22179), .B(n22180), .Z(n14702) );
  NANDN U28998 ( .A(init), .B(e[675]), .Z(n22180) );
  AND U28999 ( .A(n22181), .B(n22182), .Z(n22179) );
  NAND U29000 ( .A(ereg[674]), .B(n19486), .Z(n22182) );
  NANDN U29001 ( .A(n19481), .B(ereg[675]), .Z(n22181) );
  NAND U29002 ( .A(n22183), .B(n22184), .Z(n14701) );
  NANDN U29003 ( .A(init), .B(e[676]), .Z(n22184) );
  AND U29004 ( .A(n22185), .B(n22186), .Z(n22183) );
  NAND U29005 ( .A(ereg[675]), .B(n19486), .Z(n22186) );
  NANDN U29006 ( .A(n19481), .B(ereg[676]), .Z(n22185) );
  NAND U29007 ( .A(n22187), .B(n22188), .Z(n14700) );
  NANDN U29008 ( .A(init), .B(e[677]), .Z(n22188) );
  AND U29009 ( .A(n22189), .B(n22190), .Z(n22187) );
  NAND U29010 ( .A(ereg[676]), .B(n19486), .Z(n22190) );
  NANDN U29011 ( .A(n19481), .B(ereg[677]), .Z(n22189) );
  NAND U29012 ( .A(n22191), .B(n22192), .Z(n14699) );
  NANDN U29013 ( .A(init), .B(e[678]), .Z(n22192) );
  AND U29014 ( .A(n22193), .B(n22194), .Z(n22191) );
  NAND U29015 ( .A(ereg[677]), .B(n19486), .Z(n22194) );
  NANDN U29016 ( .A(n19481), .B(ereg[678]), .Z(n22193) );
  NAND U29017 ( .A(n22195), .B(n22196), .Z(n14698) );
  NANDN U29018 ( .A(init), .B(e[679]), .Z(n22196) );
  AND U29019 ( .A(n22197), .B(n22198), .Z(n22195) );
  NAND U29020 ( .A(ereg[678]), .B(n19486), .Z(n22198) );
  NANDN U29021 ( .A(n19481), .B(ereg[679]), .Z(n22197) );
  NAND U29022 ( .A(n22199), .B(n22200), .Z(n14697) );
  NANDN U29023 ( .A(init), .B(e[680]), .Z(n22200) );
  AND U29024 ( .A(n22201), .B(n22202), .Z(n22199) );
  NAND U29025 ( .A(ereg[679]), .B(n19486), .Z(n22202) );
  NANDN U29026 ( .A(n19481), .B(ereg[680]), .Z(n22201) );
  NAND U29027 ( .A(n22203), .B(n22204), .Z(n14696) );
  NANDN U29028 ( .A(init), .B(e[681]), .Z(n22204) );
  AND U29029 ( .A(n22205), .B(n22206), .Z(n22203) );
  NAND U29030 ( .A(ereg[680]), .B(n19486), .Z(n22206) );
  NANDN U29031 ( .A(n19481), .B(ereg[681]), .Z(n22205) );
  NAND U29032 ( .A(n22207), .B(n22208), .Z(n14695) );
  NANDN U29033 ( .A(init), .B(e[682]), .Z(n22208) );
  AND U29034 ( .A(n22209), .B(n22210), .Z(n22207) );
  NAND U29035 ( .A(ereg[681]), .B(n19486), .Z(n22210) );
  NANDN U29036 ( .A(n19481), .B(ereg[682]), .Z(n22209) );
  NAND U29037 ( .A(n22211), .B(n22212), .Z(n14694) );
  NANDN U29038 ( .A(init), .B(e[683]), .Z(n22212) );
  AND U29039 ( .A(n22213), .B(n22214), .Z(n22211) );
  NAND U29040 ( .A(ereg[682]), .B(n19486), .Z(n22214) );
  NANDN U29041 ( .A(n19481), .B(ereg[683]), .Z(n22213) );
  NAND U29042 ( .A(n22215), .B(n22216), .Z(n14693) );
  NANDN U29043 ( .A(init), .B(e[684]), .Z(n22216) );
  AND U29044 ( .A(n22217), .B(n22218), .Z(n22215) );
  NAND U29045 ( .A(ereg[683]), .B(n19486), .Z(n22218) );
  NANDN U29046 ( .A(n19481), .B(ereg[684]), .Z(n22217) );
  NAND U29047 ( .A(n22219), .B(n22220), .Z(n14692) );
  NANDN U29048 ( .A(init), .B(e[685]), .Z(n22220) );
  AND U29049 ( .A(n22221), .B(n22222), .Z(n22219) );
  NAND U29050 ( .A(ereg[684]), .B(n19486), .Z(n22222) );
  NANDN U29051 ( .A(n19481), .B(ereg[685]), .Z(n22221) );
  NAND U29052 ( .A(n22223), .B(n22224), .Z(n14691) );
  NANDN U29053 ( .A(init), .B(e[686]), .Z(n22224) );
  AND U29054 ( .A(n22225), .B(n22226), .Z(n22223) );
  NAND U29055 ( .A(ereg[685]), .B(n19486), .Z(n22226) );
  NANDN U29056 ( .A(n19481), .B(ereg[686]), .Z(n22225) );
  NAND U29057 ( .A(n22227), .B(n22228), .Z(n14690) );
  NANDN U29058 ( .A(init), .B(e[687]), .Z(n22228) );
  AND U29059 ( .A(n22229), .B(n22230), .Z(n22227) );
  NAND U29060 ( .A(ereg[686]), .B(n19486), .Z(n22230) );
  NANDN U29061 ( .A(n19481), .B(ereg[687]), .Z(n22229) );
  NAND U29062 ( .A(n22231), .B(n22232), .Z(n14689) );
  NANDN U29063 ( .A(init), .B(e[688]), .Z(n22232) );
  AND U29064 ( .A(n22233), .B(n22234), .Z(n22231) );
  NAND U29065 ( .A(ereg[687]), .B(n19486), .Z(n22234) );
  NANDN U29066 ( .A(n19481), .B(ereg[688]), .Z(n22233) );
  NAND U29067 ( .A(n22235), .B(n22236), .Z(n14688) );
  NANDN U29068 ( .A(init), .B(e[689]), .Z(n22236) );
  AND U29069 ( .A(n22237), .B(n22238), .Z(n22235) );
  NAND U29070 ( .A(ereg[688]), .B(n19486), .Z(n22238) );
  NANDN U29071 ( .A(n19481), .B(ereg[689]), .Z(n22237) );
  NAND U29072 ( .A(n22239), .B(n22240), .Z(n14687) );
  NANDN U29073 ( .A(init), .B(e[690]), .Z(n22240) );
  AND U29074 ( .A(n22241), .B(n22242), .Z(n22239) );
  NAND U29075 ( .A(ereg[689]), .B(n19486), .Z(n22242) );
  NANDN U29076 ( .A(n19481), .B(ereg[690]), .Z(n22241) );
  NAND U29077 ( .A(n22243), .B(n22244), .Z(n14686) );
  NANDN U29078 ( .A(init), .B(e[691]), .Z(n22244) );
  AND U29079 ( .A(n22245), .B(n22246), .Z(n22243) );
  NAND U29080 ( .A(ereg[690]), .B(n19486), .Z(n22246) );
  NANDN U29081 ( .A(n19481), .B(ereg[691]), .Z(n22245) );
  NAND U29082 ( .A(n22247), .B(n22248), .Z(n14685) );
  NANDN U29083 ( .A(init), .B(e[692]), .Z(n22248) );
  AND U29084 ( .A(n22249), .B(n22250), .Z(n22247) );
  NAND U29085 ( .A(ereg[691]), .B(n19486), .Z(n22250) );
  NANDN U29086 ( .A(n19481), .B(ereg[692]), .Z(n22249) );
  NAND U29087 ( .A(n22251), .B(n22252), .Z(n14684) );
  NANDN U29088 ( .A(init), .B(e[693]), .Z(n22252) );
  AND U29089 ( .A(n22253), .B(n22254), .Z(n22251) );
  NAND U29090 ( .A(ereg[692]), .B(n19486), .Z(n22254) );
  NANDN U29091 ( .A(n19481), .B(ereg[693]), .Z(n22253) );
  NAND U29092 ( .A(n22255), .B(n22256), .Z(n14683) );
  NANDN U29093 ( .A(init), .B(e[694]), .Z(n22256) );
  AND U29094 ( .A(n22257), .B(n22258), .Z(n22255) );
  NAND U29095 ( .A(ereg[693]), .B(n19486), .Z(n22258) );
  NANDN U29096 ( .A(n19481), .B(ereg[694]), .Z(n22257) );
  NAND U29097 ( .A(n22259), .B(n22260), .Z(n14682) );
  NANDN U29098 ( .A(init), .B(e[695]), .Z(n22260) );
  AND U29099 ( .A(n22261), .B(n22262), .Z(n22259) );
  NAND U29100 ( .A(ereg[694]), .B(n19486), .Z(n22262) );
  NANDN U29101 ( .A(n19481), .B(ereg[695]), .Z(n22261) );
  NAND U29102 ( .A(n22263), .B(n22264), .Z(n14681) );
  NANDN U29103 ( .A(init), .B(e[696]), .Z(n22264) );
  AND U29104 ( .A(n22265), .B(n22266), .Z(n22263) );
  NAND U29105 ( .A(ereg[695]), .B(n19486), .Z(n22266) );
  NANDN U29106 ( .A(n19481), .B(ereg[696]), .Z(n22265) );
  NAND U29107 ( .A(n22267), .B(n22268), .Z(n14680) );
  NANDN U29108 ( .A(init), .B(e[697]), .Z(n22268) );
  AND U29109 ( .A(n22269), .B(n22270), .Z(n22267) );
  NAND U29110 ( .A(ereg[696]), .B(n19486), .Z(n22270) );
  NANDN U29111 ( .A(n19481), .B(ereg[697]), .Z(n22269) );
  NAND U29112 ( .A(n22271), .B(n22272), .Z(n14679) );
  NANDN U29113 ( .A(init), .B(e[698]), .Z(n22272) );
  AND U29114 ( .A(n22273), .B(n22274), .Z(n22271) );
  NAND U29115 ( .A(ereg[697]), .B(n19486), .Z(n22274) );
  NANDN U29116 ( .A(n19481), .B(ereg[698]), .Z(n22273) );
  NAND U29117 ( .A(n22275), .B(n22276), .Z(n14678) );
  NANDN U29118 ( .A(init), .B(e[699]), .Z(n22276) );
  AND U29119 ( .A(n22277), .B(n22278), .Z(n22275) );
  NAND U29120 ( .A(ereg[698]), .B(n19486), .Z(n22278) );
  NANDN U29121 ( .A(n19481), .B(ereg[699]), .Z(n22277) );
  NAND U29122 ( .A(n22279), .B(n22280), .Z(n14677) );
  NANDN U29123 ( .A(init), .B(e[700]), .Z(n22280) );
  AND U29124 ( .A(n22281), .B(n22282), .Z(n22279) );
  NAND U29125 ( .A(ereg[699]), .B(n19486), .Z(n22282) );
  NANDN U29126 ( .A(n19481), .B(ereg[700]), .Z(n22281) );
  NAND U29127 ( .A(n22283), .B(n22284), .Z(n14676) );
  NANDN U29128 ( .A(init), .B(e[701]), .Z(n22284) );
  AND U29129 ( .A(n22285), .B(n22286), .Z(n22283) );
  NAND U29130 ( .A(ereg[700]), .B(n19486), .Z(n22286) );
  NANDN U29131 ( .A(n19481), .B(ereg[701]), .Z(n22285) );
  NAND U29132 ( .A(n22287), .B(n22288), .Z(n14675) );
  NANDN U29133 ( .A(init), .B(e[702]), .Z(n22288) );
  AND U29134 ( .A(n22289), .B(n22290), .Z(n22287) );
  NAND U29135 ( .A(ereg[701]), .B(n19486), .Z(n22290) );
  NANDN U29136 ( .A(n19481), .B(ereg[702]), .Z(n22289) );
  NAND U29137 ( .A(n22291), .B(n22292), .Z(n14674) );
  NANDN U29138 ( .A(init), .B(e[703]), .Z(n22292) );
  AND U29139 ( .A(n22293), .B(n22294), .Z(n22291) );
  NAND U29140 ( .A(ereg[702]), .B(n19486), .Z(n22294) );
  NANDN U29141 ( .A(n19481), .B(ereg[703]), .Z(n22293) );
  NAND U29142 ( .A(n22295), .B(n22296), .Z(n14673) );
  NANDN U29143 ( .A(init), .B(e[704]), .Z(n22296) );
  AND U29144 ( .A(n22297), .B(n22298), .Z(n22295) );
  NAND U29145 ( .A(ereg[703]), .B(n19486), .Z(n22298) );
  NANDN U29146 ( .A(n19481), .B(ereg[704]), .Z(n22297) );
  NAND U29147 ( .A(n22299), .B(n22300), .Z(n14672) );
  NANDN U29148 ( .A(init), .B(e[705]), .Z(n22300) );
  AND U29149 ( .A(n22301), .B(n22302), .Z(n22299) );
  NAND U29150 ( .A(ereg[704]), .B(n19486), .Z(n22302) );
  NANDN U29151 ( .A(n19481), .B(ereg[705]), .Z(n22301) );
  NAND U29152 ( .A(n22303), .B(n22304), .Z(n14671) );
  NANDN U29153 ( .A(init), .B(e[706]), .Z(n22304) );
  AND U29154 ( .A(n22305), .B(n22306), .Z(n22303) );
  NAND U29155 ( .A(ereg[705]), .B(n19486), .Z(n22306) );
  NANDN U29156 ( .A(n19481), .B(ereg[706]), .Z(n22305) );
  NAND U29157 ( .A(n22307), .B(n22308), .Z(n14670) );
  NANDN U29158 ( .A(init), .B(e[707]), .Z(n22308) );
  AND U29159 ( .A(n22309), .B(n22310), .Z(n22307) );
  NAND U29160 ( .A(ereg[706]), .B(n19486), .Z(n22310) );
  NANDN U29161 ( .A(n19481), .B(ereg[707]), .Z(n22309) );
  NAND U29162 ( .A(n22311), .B(n22312), .Z(n14669) );
  NANDN U29163 ( .A(init), .B(e[708]), .Z(n22312) );
  AND U29164 ( .A(n22313), .B(n22314), .Z(n22311) );
  NAND U29165 ( .A(ereg[707]), .B(n19486), .Z(n22314) );
  NANDN U29166 ( .A(n19481), .B(ereg[708]), .Z(n22313) );
  NAND U29167 ( .A(n22315), .B(n22316), .Z(n14668) );
  NANDN U29168 ( .A(init), .B(e[709]), .Z(n22316) );
  AND U29169 ( .A(n22317), .B(n22318), .Z(n22315) );
  NAND U29170 ( .A(ereg[708]), .B(n19486), .Z(n22318) );
  NANDN U29171 ( .A(n19481), .B(ereg[709]), .Z(n22317) );
  NAND U29172 ( .A(n22319), .B(n22320), .Z(n14667) );
  NANDN U29173 ( .A(init), .B(e[710]), .Z(n22320) );
  AND U29174 ( .A(n22321), .B(n22322), .Z(n22319) );
  NAND U29175 ( .A(ereg[709]), .B(n19486), .Z(n22322) );
  NANDN U29176 ( .A(n19481), .B(ereg[710]), .Z(n22321) );
  NAND U29177 ( .A(n22323), .B(n22324), .Z(n14666) );
  NANDN U29178 ( .A(init), .B(e[711]), .Z(n22324) );
  AND U29179 ( .A(n22325), .B(n22326), .Z(n22323) );
  NAND U29180 ( .A(ereg[710]), .B(n19486), .Z(n22326) );
  NANDN U29181 ( .A(n19481), .B(ereg[711]), .Z(n22325) );
  NAND U29182 ( .A(n22327), .B(n22328), .Z(n14665) );
  NANDN U29183 ( .A(init), .B(e[712]), .Z(n22328) );
  AND U29184 ( .A(n22329), .B(n22330), .Z(n22327) );
  NAND U29185 ( .A(ereg[711]), .B(n19486), .Z(n22330) );
  NANDN U29186 ( .A(n19481), .B(ereg[712]), .Z(n22329) );
  NAND U29187 ( .A(n22331), .B(n22332), .Z(n14664) );
  NANDN U29188 ( .A(init), .B(e[713]), .Z(n22332) );
  AND U29189 ( .A(n22333), .B(n22334), .Z(n22331) );
  NAND U29190 ( .A(ereg[712]), .B(n19486), .Z(n22334) );
  NANDN U29191 ( .A(n19481), .B(ereg[713]), .Z(n22333) );
  NAND U29192 ( .A(n22335), .B(n22336), .Z(n14663) );
  NANDN U29193 ( .A(init), .B(e[714]), .Z(n22336) );
  AND U29194 ( .A(n22337), .B(n22338), .Z(n22335) );
  NAND U29195 ( .A(ereg[713]), .B(n19486), .Z(n22338) );
  NANDN U29196 ( .A(n19481), .B(ereg[714]), .Z(n22337) );
  NAND U29197 ( .A(n22339), .B(n22340), .Z(n14662) );
  NANDN U29198 ( .A(init), .B(e[715]), .Z(n22340) );
  AND U29199 ( .A(n22341), .B(n22342), .Z(n22339) );
  NAND U29200 ( .A(ereg[714]), .B(n19486), .Z(n22342) );
  NANDN U29201 ( .A(n19481), .B(ereg[715]), .Z(n22341) );
  NAND U29202 ( .A(n22343), .B(n22344), .Z(n14661) );
  NANDN U29203 ( .A(init), .B(e[716]), .Z(n22344) );
  AND U29204 ( .A(n22345), .B(n22346), .Z(n22343) );
  NAND U29205 ( .A(ereg[715]), .B(n19486), .Z(n22346) );
  NANDN U29206 ( .A(n19481), .B(ereg[716]), .Z(n22345) );
  NAND U29207 ( .A(n22347), .B(n22348), .Z(n14660) );
  NANDN U29208 ( .A(init), .B(e[717]), .Z(n22348) );
  AND U29209 ( .A(n22349), .B(n22350), .Z(n22347) );
  NAND U29210 ( .A(ereg[716]), .B(n19486), .Z(n22350) );
  NANDN U29211 ( .A(n19481), .B(ereg[717]), .Z(n22349) );
  NAND U29212 ( .A(n22351), .B(n22352), .Z(n14659) );
  NANDN U29213 ( .A(init), .B(e[718]), .Z(n22352) );
  AND U29214 ( .A(n22353), .B(n22354), .Z(n22351) );
  NAND U29215 ( .A(ereg[717]), .B(n19486), .Z(n22354) );
  NANDN U29216 ( .A(n19481), .B(ereg[718]), .Z(n22353) );
  NAND U29217 ( .A(n22355), .B(n22356), .Z(n14658) );
  NANDN U29218 ( .A(init), .B(e[719]), .Z(n22356) );
  AND U29219 ( .A(n22357), .B(n22358), .Z(n22355) );
  NAND U29220 ( .A(ereg[718]), .B(n19486), .Z(n22358) );
  NANDN U29221 ( .A(n19481), .B(ereg[719]), .Z(n22357) );
  NAND U29222 ( .A(n22359), .B(n22360), .Z(n14657) );
  NANDN U29223 ( .A(init), .B(e[720]), .Z(n22360) );
  AND U29224 ( .A(n22361), .B(n22362), .Z(n22359) );
  NAND U29225 ( .A(ereg[719]), .B(n19486), .Z(n22362) );
  NANDN U29226 ( .A(n19481), .B(ereg[720]), .Z(n22361) );
  NAND U29227 ( .A(n22363), .B(n22364), .Z(n14656) );
  NANDN U29228 ( .A(init), .B(e[721]), .Z(n22364) );
  AND U29229 ( .A(n22365), .B(n22366), .Z(n22363) );
  NAND U29230 ( .A(ereg[720]), .B(n19486), .Z(n22366) );
  NANDN U29231 ( .A(n19481), .B(ereg[721]), .Z(n22365) );
  NAND U29232 ( .A(n22367), .B(n22368), .Z(n14655) );
  NANDN U29233 ( .A(init), .B(e[722]), .Z(n22368) );
  AND U29234 ( .A(n22369), .B(n22370), .Z(n22367) );
  NAND U29235 ( .A(ereg[721]), .B(n19486), .Z(n22370) );
  NANDN U29236 ( .A(n19481), .B(ereg[722]), .Z(n22369) );
  NAND U29237 ( .A(n22371), .B(n22372), .Z(n14654) );
  NANDN U29238 ( .A(init), .B(e[723]), .Z(n22372) );
  AND U29239 ( .A(n22373), .B(n22374), .Z(n22371) );
  NAND U29240 ( .A(ereg[722]), .B(n19486), .Z(n22374) );
  NANDN U29241 ( .A(n19481), .B(ereg[723]), .Z(n22373) );
  NAND U29242 ( .A(n22375), .B(n22376), .Z(n14653) );
  NANDN U29243 ( .A(init), .B(e[724]), .Z(n22376) );
  AND U29244 ( .A(n22377), .B(n22378), .Z(n22375) );
  NAND U29245 ( .A(ereg[723]), .B(n19486), .Z(n22378) );
  NANDN U29246 ( .A(n19481), .B(ereg[724]), .Z(n22377) );
  NAND U29247 ( .A(n22379), .B(n22380), .Z(n14652) );
  NANDN U29248 ( .A(init), .B(e[725]), .Z(n22380) );
  AND U29249 ( .A(n22381), .B(n22382), .Z(n22379) );
  NAND U29250 ( .A(ereg[724]), .B(n19486), .Z(n22382) );
  NANDN U29251 ( .A(n19481), .B(ereg[725]), .Z(n22381) );
  NAND U29252 ( .A(n22383), .B(n22384), .Z(n14651) );
  NANDN U29253 ( .A(init), .B(e[726]), .Z(n22384) );
  AND U29254 ( .A(n22385), .B(n22386), .Z(n22383) );
  NAND U29255 ( .A(ereg[725]), .B(n19486), .Z(n22386) );
  NANDN U29256 ( .A(n19481), .B(ereg[726]), .Z(n22385) );
  NAND U29257 ( .A(n22387), .B(n22388), .Z(n14650) );
  NANDN U29258 ( .A(init), .B(e[727]), .Z(n22388) );
  AND U29259 ( .A(n22389), .B(n22390), .Z(n22387) );
  NAND U29260 ( .A(ereg[726]), .B(n19486), .Z(n22390) );
  NANDN U29261 ( .A(n19481), .B(ereg[727]), .Z(n22389) );
  NAND U29262 ( .A(n22391), .B(n22392), .Z(n14649) );
  NANDN U29263 ( .A(init), .B(e[728]), .Z(n22392) );
  AND U29264 ( .A(n22393), .B(n22394), .Z(n22391) );
  NAND U29265 ( .A(ereg[727]), .B(n19486), .Z(n22394) );
  NANDN U29266 ( .A(n19481), .B(ereg[728]), .Z(n22393) );
  NAND U29267 ( .A(n22395), .B(n22396), .Z(n14648) );
  NANDN U29268 ( .A(init), .B(e[729]), .Z(n22396) );
  AND U29269 ( .A(n22397), .B(n22398), .Z(n22395) );
  NAND U29270 ( .A(ereg[728]), .B(n19486), .Z(n22398) );
  NANDN U29271 ( .A(n19481), .B(ereg[729]), .Z(n22397) );
  NAND U29272 ( .A(n22399), .B(n22400), .Z(n14647) );
  NANDN U29273 ( .A(init), .B(e[730]), .Z(n22400) );
  AND U29274 ( .A(n22401), .B(n22402), .Z(n22399) );
  NAND U29275 ( .A(ereg[729]), .B(n19486), .Z(n22402) );
  NANDN U29276 ( .A(n19481), .B(ereg[730]), .Z(n22401) );
  NAND U29277 ( .A(n22403), .B(n22404), .Z(n14646) );
  NANDN U29278 ( .A(init), .B(e[731]), .Z(n22404) );
  AND U29279 ( .A(n22405), .B(n22406), .Z(n22403) );
  NAND U29280 ( .A(ereg[730]), .B(n19486), .Z(n22406) );
  NANDN U29281 ( .A(n19481), .B(ereg[731]), .Z(n22405) );
  NAND U29282 ( .A(n22407), .B(n22408), .Z(n14645) );
  NANDN U29283 ( .A(init), .B(e[732]), .Z(n22408) );
  AND U29284 ( .A(n22409), .B(n22410), .Z(n22407) );
  NAND U29285 ( .A(ereg[731]), .B(n19486), .Z(n22410) );
  NANDN U29286 ( .A(n19481), .B(ereg[732]), .Z(n22409) );
  NAND U29287 ( .A(n22411), .B(n22412), .Z(n14644) );
  NANDN U29288 ( .A(init), .B(e[733]), .Z(n22412) );
  AND U29289 ( .A(n22413), .B(n22414), .Z(n22411) );
  NAND U29290 ( .A(ereg[732]), .B(n19486), .Z(n22414) );
  NANDN U29291 ( .A(n19481), .B(ereg[733]), .Z(n22413) );
  NAND U29292 ( .A(n22415), .B(n22416), .Z(n14643) );
  NANDN U29293 ( .A(init), .B(e[734]), .Z(n22416) );
  AND U29294 ( .A(n22417), .B(n22418), .Z(n22415) );
  NAND U29295 ( .A(ereg[733]), .B(n19486), .Z(n22418) );
  NANDN U29296 ( .A(n19481), .B(ereg[734]), .Z(n22417) );
  NAND U29297 ( .A(n22419), .B(n22420), .Z(n14642) );
  NANDN U29298 ( .A(init), .B(e[735]), .Z(n22420) );
  AND U29299 ( .A(n22421), .B(n22422), .Z(n22419) );
  NAND U29300 ( .A(ereg[734]), .B(n19486), .Z(n22422) );
  NANDN U29301 ( .A(n19481), .B(ereg[735]), .Z(n22421) );
  NAND U29302 ( .A(n22423), .B(n22424), .Z(n14641) );
  NANDN U29303 ( .A(init), .B(e[736]), .Z(n22424) );
  AND U29304 ( .A(n22425), .B(n22426), .Z(n22423) );
  NAND U29305 ( .A(ereg[735]), .B(n19486), .Z(n22426) );
  NANDN U29306 ( .A(n19481), .B(ereg[736]), .Z(n22425) );
  NAND U29307 ( .A(n22427), .B(n22428), .Z(n14640) );
  NANDN U29308 ( .A(init), .B(e[737]), .Z(n22428) );
  AND U29309 ( .A(n22429), .B(n22430), .Z(n22427) );
  NAND U29310 ( .A(ereg[736]), .B(n19486), .Z(n22430) );
  NANDN U29311 ( .A(n19481), .B(ereg[737]), .Z(n22429) );
  NAND U29312 ( .A(n22431), .B(n22432), .Z(n14639) );
  NANDN U29313 ( .A(init), .B(e[738]), .Z(n22432) );
  AND U29314 ( .A(n22433), .B(n22434), .Z(n22431) );
  NAND U29315 ( .A(ereg[737]), .B(n19486), .Z(n22434) );
  NANDN U29316 ( .A(n19481), .B(ereg[738]), .Z(n22433) );
  NAND U29317 ( .A(n22435), .B(n22436), .Z(n14638) );
  NANDN U29318 ( .A(init), .B(e[739]), .Z(n22436) );
  AND U29319 ( .A(n22437), .B(n22438), .Z(n22435) );
  NAND U29320 ( .A(ereg[738]), .B(n19486), .Z(n22438) );
  NANDN U29321 ( .A(n19481), .B(ereg[739]), .Z(n22437) );
  NAND U29322 ( .A(n22439), .B(n22440), .Z(n14637) );
  NANDN U29323 ( .A(init), .B(e[740]), .Z(n22440) );
  AND U29324 ( .A(n22441), .B(n22442), .Z(n22439) );
  NAND U29325 ( .A(ereg[739]), .B(n19486), .Z(n22442) );
  NANDN U29326 ( .A(n19481), .B(ereg[740]), .Z(n22441) );
  NAND U29327 ( .A(n22443), .B(n22444), .Z(n14636) );
  NANDN U29328 ( .A(init), .B(e[741]), .Z(n22444) );
  AND U29329 ( .A(n22445), .B(n22446), .Z(n22443) );
  NAND U29330 ( .A(ereg[740]), .B(n19486), .Z(n22446) );
  NANDN U29331 ( .A(n19481), .B(ereg[741]), .Z(n22445) );
  NAND U29332 ( .A(n22447), .B(n22448), .Z(n14635) );
  NANDN U29333 ( .A(init), .B(e[742]), .Z(n22448) );
  AND U29334 ( .A(n22449), .B(n22450), .Z(n22447) );
  NAND U29335 ( .A(ereg[741]), .B(n19486), .Z(n22450) );
  NANDN U29336 ( .A(n19481), .B(ereg[742]), .Z(n22449) );
  NAND U29337 ( .A(n22451), .B(n22452), .Z(n14634) );
  NANDN U29338 ( .A(init), .B(e[743]), .Z(n22452) );
  AND U29339 ( .A(n22453), .B(n22454), .Z(n22451) );
  NAND U29340 ( .A(ereg[742]), .B(n19486), .Z(n22454) );
  NANDN U29341 ( .A(n19481), .B(ereg[743]), .Z(n22453) );
  NAND U29342 ( .A(n22455), .B(n22456), .Z(n14633) );
  NANDN U29343 ( .A(init), .B(e[744]), .Z(n22456) );
  AND U29344 ( .A(n22457), .B(n22458), .Z(n22455) );
  NAND U29345 ( .A(ereg[743]), .B(n19486), .Z(n22458) );
  NANDN U29346 ( .A(n19481), .B(ereg[744]), .Z(n22457) );
  NAND U29347 ( .A(n22459), .B(n22460), .Z(n14632) );
  NANDN U29348 ( .A(init), .B(e[745]), .Z(n22460) );
  AND U29349 ( .A(n22461), .B(n22462), .Z(n22459) );
  NAND U29350 ( .A(ereg[744]), .B(n19486), .Z(n22462) );
  NANDN U29351 ( .A(n19481), .B(ereg[745]), .Z(n22461) );
  NAND U29352 ( .A(n22463), .B(n22464), .Z(n14631) );
  NANDN U29353 ( .A(init), .B(e[746]), .Z(n22464) );
  AND U29354 ( .A(n22465), .B(n22466), .Z(n22463) );
  NAND U29355 ( .A(ereg[745]), .B(n19486), .Z(n22466) );
  NANDN U29356 ( .A(n19481), .B(ereg[746]), .Z(n22465) );
  NAND U29357 ( .A(n22467), .B(n22468), .Z(n14630) );
  NANDN U29358 ( .A(init), .B(e[747]), .Z(n22468) );
  AND U29359 ( .A(n22469), .B(n22470), .Z(n22467) );
  NAND U29360 ( .A(ereg[746]), .B(n19486), .Z(n22470) );
  NANDN U29361 ( .A(n19481), .B(ereg[747]), .Z(n22469) );
  NAND U29362 ( .A(n22471), .B(n22472), .Z(n14629) );
  NANDN U29363 ( .A(init), .B(e[748]), .Z(n22472) );
  AND U29364 ( .A(n22473), .B(n22474), .Z(n22471) );
  NAND U29365 ( .A(ereg[747]), .B(n19486), .Z(n22474) );
  NANDN U29366 ( .A(n19481), .B(ereg[748]), .Z(n22473) );
  NAND U29367 ( .A(n22475), .B(n22476), .Z(n14628) );
  NANDN U29368 ( .A(init), .B(e[749]), .Z(n22476) );
  AND U29369 ( .A(n22477), .B(n22478), .Z(n22475) );
  NAND U29370 ( .A(ereg[748]), .B(n19486), .Z(n22478) );
  NANDN U29371 ( .A(n19481), .B(ereg[749]), .Z(n22477) );
  NAND U29372 ( .A(n22479), .B(n22480), .Z(n14627) );
  NANDN U29373 ( .A(init), .B(e[750]), .Z(n22480) );
  AND U29374 ( .A(n22481), .B(n22482), .Z(n22479) );
  NAND U29375 ( .A(ereg[749]), .B(n19486), .Z(n22482) );
  NANDN U29376 ( .A(n19481), .B(ereg[750]), .Z(n22481) );
  NAND U29377 ( .A(n22483), .B(n22484), .Z(n14626) );
  NANDN U29378 ( .A(init), .B(e[751]), .Z(n22484) );
  AND U29379 ( .A(n22485), .B(n22486), .Z(n22483) );
  NAND U29380 ( .A(ereg[750]), .B(n19486), .Z(n22486) );
  NANDN U29381 ( .A(n19481), .B(ereg[751]), .Z(n22485) );
  NAND U29382 ( .A(n22487), .B(n22488), .Z(n14625) );
  NANDN U29383 ( .A(init), .B(e[752]), .Z(n22488) );
  AND U29384 ( .A(n22489), .B(n22490), .Z(n22487) );
  NAND U29385 ( .A(ereg[751]), .B(n19486), .Z(n22490) );
  NANDN U29386 ( .A(n19481), .B(ereg[752]), .Z(n22489) );
  NAND U29387 ( .A(n22491), .B(n22492), .Z(n14624) );
  NANDN U29388 ( .A(init), .B(e[753]), .Z(n22492) );
  AND U29389 ( .A(n22493), .B(n22494), .Z(n22491) );
  NAND U29390 ( .A(ereg[752]), .B(n19486), .Z(n22494) );
  NANDN U29391 ( .A(n19481), .B(ereg[753]), .Z(n22493) );
  NAND U29392 ( .A(n22495), .B(n22496), .Z(n14623) );
  NANDN U29393 ( .A(init), .B(e[754]), .Z(n22496) );
  AND U29394 ( .A(n22497), .B(n22498), .Z(n22495) );
  NAND U29395 ( .A(ereg[753]), .B(n19486), .Z(n22498) );
  NANDN U29396 ( .A(n19481), .B(ereg[754]), .Z(n22497) );
  NAND U29397 ( .A(n22499), .B(n22500), .Z(n14622) );
  NANDN U29398 ( .A(init), .B(e[755]), .Z(n22500) );
  AND U29399 ( .A(n22501), .B(n22502), .Z(n22499) );
  NAND U29400 ( .A(ereg[754]), .B(n19486), .Z(n22502) );
  NANDN U29401 ( .A(n19481), .B(ereg[755]), .Z(n22501) );
  NAND U29402 ( .A(n22503), .B(n22504), .Z(n14621) );
  NANDN U29403 ( .A(init), .B(e[756]), .Z(n22504) );
  AND U29404 ( .A(n22505), .B(n22506), .Z(n22503) );
  NAND U29405 ( .A(ereg[755]), .B(n19486), .Z(n22506) );
  NANDN U29406 ( .A(n19481), .B(ereg[756]), .Z(n22505) );
  NAND U29407 ( .A(n22507), .B(n22508), .Z(n14620) );
  NANDN U29408 ( .A(init), .B(e[757]), .Z(n22508) );
  AND U29409 ( .A(n22509), .B(n22510), .Z(n22507) );
  NAND U29410 ( .A(ereg[756]), .B(n19486), .Z(n22510) );
  NANDN U29411 ( .A(n19481), .B(ereg[757]), .Z(n22509) );
  NAND U29412 ( .A(n22511), .B(n22512), .Z(n14619) );
  NANDN U29413 ( .A(init), .B(e[758]), .Z(n22512) );
  AND U29414 ( .A(n22513), .B(n22514), .Z(n22511) );
  NAND U29415 ( .A(ereg[757]), .B(n19486), .Z(n22514) );
  NANDN U29416 ( .A(n19481), .B(ereg[758]), .Z(n22513) );
  NAND U29417 ( .A(n22515), .B(n22516), .Z(n14618) );
  NANDN U29418 ( .A(init), .B(e[759]), .Z(n22516) );
  AND U29419 ( .A(n22517), .B(n22518), .Z(n22515) );
  NAND U29420 ( .A(ereg[758]), .B(n19486), .Z(n22518) );
  NANDN U29421 ( .A(n19481), .B(ereg[759]), .Z(n22517) );
  NAND U29422 ( .A(n22519), .B(n22520), .Z(n14617) );
  NANDN U29423 ( .A(init), .B(e[760]), .Z(n22520) );
  AND U29424 ( .A(n22521), .B(n22522), .Z(n22519) );
  NAND U29425 ( .A(ereg[759]), .B(n19486), .Z(n22522) );
  NANDN U29426 ( .A(n19481), .B(ereg[760]), .Z(n22521) );
  NAND U29427 ( .A(n22523), .B(n22524), .Z(n14616) );
  NANDN U29428 ( .A(init), .B(e[761]), .Z(n22524) );
  AND U29429 ( .A(n22525), .B(n22526), .Z(n22523) );
  NAND U29430 ( .A(ereg[760]), .B(n19486), .Z(n22526) );
  NANDN U29431 ( .A(n19481), .B(ereg[761]), .Z(n22525) );
  NAND U29432 ( .A(n22527), .B(n22528), .Z(n14615) );
  NANDN U29433 ( .A(init), .B(e[762]), .Z(n22528) );
  AND U29434 ( .A(n22529), .B(n22530), .Z(n22527) );
  NAND U29435 ( .A(ereg[761]), .B(n19486), .Z(n22530) );
  NANDN U29436 ( .A(n19481), .B(ereg[762]), .Z(n22529) );
  NAND U29437 ( .A(n22531), .B(n22532), .Z(n14614) );
  NANDN U29438 ( .A(init), .B(e[763]), .Z(n22532) );
  AND U29439 ( .A(n22533), .B(n22534), .Z(n22531) );
  NAND U29440 ( .A(ereg[762]), .B(n19486), .Z(n22534) );
  NANDN U29441 ( .A(n19481), .B(ereg[763]), .Z(n22533) );
  NAND U29442 ( .A(n22535), .B(n22536), .Z(n14613) );
  NANDN U29443 ( .A(init), .B(e[764]), .Z(n22536) );
  AND U29444 ( .A(n22537), .B(n22538), .Z(n22535) );
  NAND U29445 ( .A(ereg[763]), .B(n19486), .Z(n22538) );
  NANDN U29446 ( .A(n19481), .B(ereg[764]), .Z(n22537) );
  NAND U29447 ( .A(n22539), .B(n22540), .Z(n14612) );
  NANDN U29448 ( .A(init), .B(e[765]), .Z(n22540) );
  AND U29449 ( .A(n22541), .B(n22542), .Z(n22539) );
  NAND U29450 ( .A(ereg[764]), .B(n19486), .Z(n22542) );
  NANDN U29451 ( .A(n19481), .B(ereg[765]), .Z(n22541) );
  NAND U29452 ( .A(n22543), .B(n22544), .Z(n14611) );
  NANDN U29453 ( .A(init), .B(e[766]), .Z(n22544) );
  AND U29454 ( .A(n22545), .B(n22546), .Z(n22543) );
  NAND U29455 ( .A(ereg[765]), .B(n19486), .Z(n22546) );
  NANDN U29456 ( .A(n19481), .B(ereg[766]), .Z(n22545) );
  NAND U29457 ( .A(n22547), .B(n22548), .Z(n14610) );
  NANDN U29458 ( .A(init), .B(e[767]), .Z(n22548) );
  AND U29459 ( .A(n22549), .B(n22550), .Z(n22547) );
  NAND U29460 ( .A(ereg[766]), .B(n19486), .Z(n22550) );
  NANDN U29461 ( .A(n19481), .B(ereg[767]), .Z(n22549) );
  NAND U29462 ( .A(n22551), .B(n22552), .Z(n14609) );
  NANDN U29463 ( .A(init), .B(e[768]), .Z(n22552) );
  AND U29464 ( .A(n22553), .B(n22554), .Z(n22551) );
  NAND U29465 ( .A(ereg[767]), .B(n19486), .Z(n22554) );
  NANDN U29466 ( .A(n19481), .B(ereg[768]), .Z(n22553) );
  NAND U29467 ( .A(n22555), .B(n22556), .Z(n14608) );
  NANDN U29468 ( .A(init), .B(e[769]), .Z(n22556) );
  AND U29469 ( .A(n22557), .B(n22558), .Z(n22555) );
  NAND U29470 ( .A(ereg[768]), .B(n19486), .Z(n22558) );
  NANDN U29471 ( .A(n19481), .B(ereg[769]), .Z(n22557) );
  NAND U29472 ( .A(n22559), .B(n22560), .Z(n14607) );
  NANDN U29473 ( .A(init), .B(e[770]), .Z(n22560) );
  AND U29474 ( .A(n22561), .B(n22562), .Z(n22559) );
  NAND U29475 ( .A(ereg[769]), .B(n19486), .Z(n22562) );
  NANDN U29476 ( .A(n19481), .B(ereg[770]), .Z(n22561) );
  NAND U29477 ( .A(n22563), .B(n22564), .Z(n14606) );
  NANDN U29478 ( .A(init), .B(e[771]), .Z(n22564) );
  AND U29479 ( .A(n22565), .B(n22566), .Z(n22563) );
  NAND U29480 ( .A(ereg[770]), .B(n19486), .Z(n22566) );
  NANDN U29481 ( .A(n19481), .B(ereg[771]), .Z(n22565) );
  NAND U29482 ( .A(n22567), .B(n22568), .Z(n14605) );
  NANDN U29483 ( .A(init), .B(e[772]), .Z(n22568) );
  AND U29484 ( .A(n22569), .B(n22570), .Z(n22567) );
  NAND U29485 ( .A(ereg[771]), .B(n19486), .Z(n22570) );
  NANDN U29486 ( .A(n19481), .B(ereg[772]), .Z(n22569) );
  NAND U29487 ( .A(n22571), .B(n22572), .Z(n14604) );
  NANDN U29488 ( .A(init), .B(e[773]), .Z(n22572) );
  AND U29489 ( .A(n22573), .B(n22574), .Z(n22571) );
  NAND U29490 ( .A(ereg[772]), .B(n19486), .Z(n22574) );
  NANDN U29491 ( .A(n19481), .B(ereg[773]), .Z(n22573) );
  NAND U29492 ( .A(n22575), .B(n22576), .Z(n14603) );
  NANDN U29493 ( .A(init), .B(e[774]), .Z(n22576) );
  AND U29494 ( .A(n22577), .B(n22578), .Z(n22575) );
  NAND U29495 ( .A(ereg[773]), .B(n19486), .Z(n22578) );
  NANDN U29496 ( .A(n19481), .B(ereg[774]), .Z(n22577) );
  NAND U29497 ( .A(n22579), .B(n22580), .Z(n14602) );
  NANDN U29498 ( .A(init), .B(e[775]), .Z(n22580) );
  AND U29499 ( .A(n22581), .B(n22582), .Z(n22579) );
  NAND U29500 ( .A(ereg[774]), .B(n19486), .Z(n22582) );
  NANDN U29501 ( .A(n19481), .B(ereg[775]), .Z(n22581) );
  NAND U29502 ( .A(n22583), .B(n22584), .Z(n14601) );
  NANDN U29503 ( .A(init), .B(e[776]), .Z(n22584) );
  AND U29504 ( .A(n22585), .B(n22586), .Z(n22583) );
  NAND U29505 ( .A(ereg[775]), .B(n19486), .Z(n22586) );
  NANDN U29506 ( .A(n19481), .B(ereg[776]), .Z(n22585) );
  NAND U29507 ( .A(n22587), .B(n22588), .Z(n14600) );
  NANDN U29508 ( .A(init), .B(e[777]), .Z(n22588) );
  AND U29509 ( .A(n22589), .B(n22590), .Z(n22587) );
  NAND U29510 ( .A(ereg[776]), .B(n19486), .Z(n22590) );
  NANDN U29511 ( .A(n19481), .B(ereg[777]), .Z(n22589) );
  NAND U29512 ( .A(n22591), .B(n22592), .Z(n14599) );
  NANDN U29513 ( .A(init), .B(e[778]), .Z(n22592) );
  AND U29514 ( .A(n22593), .B(n22594), .Z(n22591) );
  NAND U29515 ( .A(ereg[777]), .B(n19486), .Z(n22594) );
  NANDN U29516 ( .A(n19481), .B(ereg[778]), .Z(n22593) );
  NAND U29517 ( .A(n22595), .B(n22596), .Z(n14598) );
  NANDN U29518 ( .A(init), .B(e[779]), .Z(n22596) );
  AND U29519 ( .A(n22597), .B(n22598), .Z(n22595) );
  NAND U29520 ( .A(ereg[778]), .B(n19486), .Z(n22598) );
  NANDN U29521 ( .A(n19481), .B(ereg[779]), .Z(n22597) );
  NAND U29522 ( .A(n22599), .B(n22600), .Z(n14597) );
  NANDN U29523 ( .A(init), .B(e[780]), .Z(n22600) );
  AND U29524 ( .A(n22601), .B(n22602), .Z(n22599) );
  NAND U29525 ( .A(ereg[779]), .B(n19486), .Z(n22602) );
  NANDN U29526 ( .A(n19481), .B(ereg[780]), .Z(n22601) );
  NAND U29527 ( .A(n22603), .B(n22604), .Z(n14596) );
  NANDN U29528 ( .A(init), .B(e[781]), .Z(n22604) );
  AND U29529 ( .A(n22605), .B(n22606), .Z(n22603) );
  NAND U29530 ( .A(ereg[780]), .B(n19486), .Z(n22606) );
  NANDN U29531 ( .A(n19481), .B(ereg[781]), .Z(n22605) );
  NAND U29532 ( .A(n22607), .B(n22608), .Z(n14595) );
  NANDN U29533 ( .A(init), .B(e[782]), .Z(n22608) );
  AND U29534 ( .A(n22609), .B(n22610), .Z(n22607) );
  NAND U29535 ( .A(ereg[781]), .B(n19486), .Z(n22610) );
  NANDN U29536 ( .A(n19481), .B(ereg[782]), .Z(n22609) );
  NAND U29537 ( .A(n22611), .B(n22612), .Z(n14594) );
  NANDN U29538 ( .A(init), .B(e[783]), .Z(n22612) );
  AND U29539 ( .A(n22613), .B(n22614), .Z(n22611) );
  NAND U29540 ( .A(ereg[782]), .B(n19486), .Z(n22614) );
  NANDN U29541 ( .A(n19481), .B(ereg[783]), .Z(n22613) );
  NAND U29542 ( .A(n22615), .B(n22616), .Z(n14593) );
  NANDN U29543 ( .A(init), .B(e[784]), .Z(n22616) );
  AND U29544 ( .A(n22617), .B(n22618), .Z(n22615) );
  NAND U29545 ( .A(ereg[783]), .B(n19486), .Z(n22618) );
  NANDN U29546 ( .A(n19481), .B(ereg[784]), .Z(n22617) );
  NAND U29547 ( .A(n22619), .B(n22620), .Z(n14592) );
  NANDN U29548 ( .A(init), .B(e[785]), .Z(n22620) );
  AND U29549 ( .A(n22621), .B(n22622), .Z(n22619) );
  NAND U29550 ( .A(ereg[784]), .B(n19486), .Z(n22622) );
  NANDN U29551 ( .A(n19481), .B(ereg[785]), .Z(n22621) );
  NAND U29552 ( .A(n22623), .B(n22624), .Z(n14591) );
  NANDN U29553 ( .A(init), .B(e[786]), .Z(n22624) );
  AND U29554 ( .A(n22625), .B(n22626), .Z(n22623) );
  NAND U29555 ( .A(ereg[785]), .B(n19486), .Z(n22626) );
  NANDN U29556 ( .A(n19481), .B(ereg[786]), .Z(n22625) );
  NAND U29557 ( .A(n22627), .B(n22628), .Z(n14590) );
  NANDN U29558 ( .A(init), .B(e[787]), .Z(n22628) );
  AND U29559 ( .A(n22629), .B(n22630), .Z(n22627) );
  NAND U29560 ( .A(ereg[786]), .B(n19486), .Z(n22630) );
  NANDN U29561 ( .A(n19481), .B(ereg[787]), .Z(n22629) );
  NAND U29562 ( .A(n22631), .B(n22632), .Z(n14589) );
  NANDN U29563 ( .A(init), .B(e[788]), .Z(n22632) );
  AND U29564 ( .A(n22633), .B(n22634), .Z(n22631) );
  NAND U29565 ( .A(ereg[787]), .B(n19486), .Z(n22634) );
  NANDN U29566 ( .A(n19481), .B(ereg[788]), .Z(n22633) );
  NAND U29567 ( .A(n22635), .B(n22636), .Z(n14588) );
  NANDN U29568 ( .A(init), .B(e[789]), .Z(n22636) );
  AND U29569 ( .A(n22637), .B(n22638), .Z(n22635) );
  NAND U29570 ( .A(ereg[788]), .B(n19486), .Z(n22638) );
  NANDN U29571 ( .A(n19481), .B(ereg[789]), .Z(n22637) );
  NAND U29572 ( .A(n22639), .B(n22640), .Z(n14587) );
  NANDN U29573 ( .A(init), .B(e[790]), .Z(n22640) );
  AND U29574 ( .A(n22641), .B(n22642), .Z(n22639) );
  NAND U29575 ( .A(ereg[789]), .B(n19486), .Z(n22642) );
  NANDN U29576 ( .A(n19481), .B(ereg[790]), .Z(n22641) );
  NAND U29577 ( .A(n22643), .B(n22644), .Z(n14586) );
  NANDN U29578 ( .A(init), .B(e[791]), .Z(n22644) );
  AND U29579 ( .A(n22645), .B(n22646), .Z(n22643) );
  NAND U29580 ( .A(ereg[790]), .B(n19486), .Z(n22646) );
  NANDN U29581 ( .A(n19481), .B(ereg[791]), .Z(n22645) );
  NAND U29582 ( .A(n22647), .B(n22648), .Z(n14585) );
  NANDN U29583 ( .A(init), .B(e[792]), .Z(n22648) );
  AND U29584 ( .A(n22649), .B(n22650), .Z(n22647) );
  NAND U29585 ( .A(ereg[791]), .B(n19486), .Z(n22650) );
  NANDN U29586 ( .A(n19481), .B(ereg[792]), .Z(n22649) );
  NAND U29587 ( .A(n22651), .B(n22652), .Z(n14584) );
  NANDN U29588 ( .A(init), .B(e[793]), .Z(n22652) );
  AND U29589 ( .A(n22653), .B(n22654), .Z(n22651) );
  NAND U29590 ( .A(ereg[792]), .B(n19486), .Z(n22654) );
  NANDN U29591 ( .A(n19481), .B(ereg[793]), .Z(n22653) );
  NAND U29592 ( .A(n22655), .B(n22656), .Z(n14583) );
  NANDN U29593 ( .A(init), .B(e[794]), .Z(n22656) );
  AND U29594 ( .A(n22657), .B(n22658), .Z(n22655) );
  NAND U29595 ( .A(ereg[793]), .B(n19486), .Z(n22658) );
  NANDN U29596 ( .A(n19481), .B(ereg[794]), .Z(n22657) );
  NAND U29597 ( .A(n22659), .B(n22660), .Z(n14582) );
  NANDN U29598 ( .A(init), .B(e[795]), .Z(n22660) );
  AND U29599 ( .A(n22661), .B(n22662), .Z(n22659) );
  NAND U29600 ( .A(ereg[794]), .B(n19486), .Z(n22662) );
  NANDN U29601 ( .A(n19481), .B(ereg[795]), .Z(n22661) );
  NAND U29602 ( .A(n22663), .B(n22664), .Z(n14581) );
  NANDN U29603 ( .A(init), .B(e[796]), .Z(n22664) );
  AND U29604 ( .A(n22665), .B(n22666), .Z(n22663) );
  NAND U29605 ( .A(ereg[795]), .B(n19486), .Z(n22666) );
  NANDN U29606 ( .A(n19481), .B(ereg[796]), .Z(n22665) );
  NAND U29607 ( .A(n22667), .B(n22668), .Z(n14580) );
  NANDN U29608 ( .A(init), .B(e[797]), .Z(n22668) );
  AND U29609 ( .A(n22669), .B(n22670), .Z(n22667) );
  NAND U29610 ( .A(ereg[796]), .B(n19486), .Z(n22670) );
  NANDN U29611 ( .A(n19481), .B(ereg[797]), .Z(n22669) );
  NAND U29612 ( .A(n22671), .B(n22672), .Z(n14579) );
  NANDN U29613 ( .A(init), .B(e[798]), .Z(n22672) );
  AND U29614 ( .A(n22673), .B(n22674), .Z(n22671) );
  NAND U29615 ( .A(ereg[797]), .B(n19486), .Z(n22674) );
  NANDN U29616 ( .A(n19481), .B(ereg[798]), .Z(n22673) );
  NAND U29617 ( .A(n22675), .B(n22676), .Z(n14578) );
  NANDN U29618 ( .A(init), .B(e[799]), .Z(n22676) );
  AND U29619 ( .A(n22677), .B(n22678), .Z(n22675) );
  NAND U29620 ( .A(ereg[798]), .B(n19486), .Z(n22678) );
  NANDN U29621 ( .A(n19481), .B(ereg[799]), .Z(n22677) );
  NAND U29622 ( .A(n22679), .B(n22680), .Z(n14577) );
  NANDN U29623 ( .A(init), .B(e[800]), .Z(n22680) );
  AND U29624 ( .A(n22681), .B(n22682), .Z(n22679) );
  NAND U29625 ( .A(ereg[799]), .B(n19486), .Z(n22682) );
  NANDN U29626 ( .A(n19481), .B(ereg[800]), .Z(n22681) );
  NAND U29627 ( .A(n22683), .B(n22684), .Z(n14576) );
  NANDN U29628 ( .A(init), .B(e[801]), .Z(n22684) );
  AND U29629 ( .A(n22685), .B(n22686), .Z(n22683) );
  NAND U29630 ( .A(ereg[800]), .B(n19486), .Z(n22686) );
  NANDN U29631 ( .A(n19481), .B(ereg[801]), .Z(n22685) );
  NAND U29632 ( .A(n22687), .B(n22688), .Z(n14575) );
  NANDN U29633 ( .A(init), .B(e[802]), .Z(n22688) );
  AND U29634 ( .A(n22689), .B(n22690), .Z(n22687) );
  NAND U29635 ( .A(ereg[801]), .B(n19486), .Z(n22690) );
  NANDN U29636 ( .A(n19481), .B(ereg[802]), .Z(n22689) );
  NAND U29637 ( .A(n22691), .B(n22692), .Z(n14574) );
  NANDN U29638 ( .A(init), .B(e[803]), .Z(n22692) );
  AND U29639 ( .A(n22693), .B(n22694), .Z(n22691) );
  NAND U29640 ( .A(ereg[802]), .B(n19486), .Z(n22694) );
  NANDN U29641 ( .A(n19481), .B(ereg[803]), .Z(n22693) );
  NAND U29642 ( .A(n22695), .B(n22696), .Z(n14573) );
  NANDN U29643 ( .A(init), .B(e[804]), .Z(n22696) );
  AND U29644 ( .A(n22697), .B(n22698), .Z(n22695) );
  NAND U29645 ( .A(ereg[803]), .B(n19486), .Z(n22698) );
  NANDN U29646 ( .A(n19481), .B(ereg[804]), .Z(n22697) );
  NAND U29647 ( .A(n22699), .B(n22700), .Z(n14572) );
  NANDN U29648 ( .A(init), .B(e[805]), .Z(n22700) );
  AND U29649 ( .A(n22701), .B(n22702), .Z(n22699) );
  NAND U29650 ( .A(ereg[804]), .B(n19486), .Z(n22702) );
  NANDN U29651 ( .A(n19481), .B(ereg[805]), .Z(n22701) );
  NAND U29652 ( .A(n22703), .B(n22704), .Z(n14571) );
  NANDN U29653 ( .A(init), .B(e[806]), .Z(n22704) );
  AND U29654 ( .A(n22705), .B(n22706), .Z(n22703) );
  NAND U29655 ( .A(ereg[805]), .B(n19486), .Z(n22706) );
  NANDN U29656 ( .A(n19481), .B(ereg[806]), .Z(n22705) );
  NAND U29657 ( .A(n22707), .B(n22708), .Z(n14570) );
  NANDN U29658 ( .A(init), .B(e[807]), .Z(n22708) );
  AND U29659 ( .A(n22709), .B(n22710), .Z(n22707) );
  NAND U29660 ( .A(ereg[806]), .B(n19486), .Z(n22710) );
  NANDN U29661 ( .A(n19481), .B(ereg[807]), .Z(n22709) );
  NAND U29662 ( .A(n22711), .B(n22712), .Z(n14569) );
  NANDN U29663 ( .A(init), .B(e[808]), .Z(n22712) );
  AND U29664 ( .A(n22713), .B(n22714), .Z(n22711) );
  NAND U29665 ( .A(ereg[807]), .B(n19486), .Z(n22714) );
  NANDN U29666 ( .A(n19481), .B(ereg[808]), .Z(n22713) );
  NAND U29667 ( .A(n22715), .B(n22716), .Z(n14568) );
  NANDN U29668 ( .A(init), .B(e[809]), .Z(n22716) );
  AND U29669 ( .A(n22717), .B(n22718), .Z(n22715) );
  NAND U29670 ( .A(ereg[808]), .B(n19486), .Z(n22718) );
  NANDN U29671 ( .A(n19481), .B(ereg[809]), .Z(n22717) );
  NAND U29672 ( .A(n22719), .B(n22720), .Z(n14567) );
  NANDN U29673 ( .A(init), .B(e[810]), .Z(n22720) );
  AND U29674 ( .A(n22721), .B(n22722), .Z(n22719) );
  NAND U29675 ( .A(ereg[809]), .B(n19486), .Z(n22722) );
  NANDN U29676 ( .A(n19481), .B(ereg[810]), .Z(n22721) );
  NAND U29677 ( .A(n22723), .B(n22724), .Z(n14566) );
  NANDN U29678 ( .A(init), .B(e[811]), .Z(n22724) );
  AND U29679 ( .A(n22725), .B(n22726), .Z(n22723) );
  NAND U29680 ( .A(ereg[810]), .B(n19486), .Z(n22726) );
  NANDN U29681 ( .A(n19481), .B(ereg[811]), .Z(n22725) );
  NAND U29682 ( .A(n22727), .B(n22728), .Z(n14565) );
  NANDN U29683 ( .A(init), .B(e[812]), .Z(n22728) );
  AND U29684 ( .A(n22729), .B(n22730), .Z(n22727) );
  NAND U29685 ( .A(ereg[811]), .B(n19486), .Z(n22730) );
  NANDN U29686 ( .A(n19481), .B(ereg[812]), .Z(n22729) );
  NAND U29687 ( .A(n22731), .B(n22732), .Z(n14564) );
  NANDN U29688 ( .A(init), .B(e[813]), .Z(n22732) );
  AND U29689 ( .A(n22733), .B(n22734), .Z(n22731) );
  NAND U29690 ( .A(ereg[812]), .B(n19486), .Z(n22734) );
  NANDN U29691 ( .A(n19481), .B(ereg[813]), .Z(n22733) );
  NAND U29692 ( .A(n22735), .B(n22736), .Z(n14563) );
  NANDN U29693 ( .A(init), .B(e[814]), .Z(n22736) );
  AND U29694 ( .A(n22737), .B(n22738), .Z(n22735) );
  NAND U29695 ( .A(ereg[813]), .B(n19486), .Z(n22738) );
  NANDN U29696 ( .A(n19481), .B(ereg[814]), .Z(n22737) );
  NAND U29697 ( .A(n22739), .B(n22740), .Z(n14562) );
  NANDN U29698 ( .A(init), .B(e[815]), .Z(n22740) );
  AND U29699 ( .A(n22741), .B(n22742), .Z(n22739) );
  NAND U29700 ( .A(ereg[814]), .B(n19486), .Z(n22742) );
  NANDN U29701 ( .A(n19481), .B(ereg[815]), .Z(n22741) );
  NAND U29702 ( .A(n22743), .B(n22744), .Z(n14561) );
  NANDN U29703 ( .A(init), .B(e[816]), .Z(n22744) );
  AND U29704 ( .A(n22745), .B(n22746), .Z(n22743) );
  NAND U29705 ( .A(ereg[815]), .B(n19486), .Z(n22746) );
  NANDN U29706 ( .A(n19481), .B(ereg[816]), .Z(n22745) );
  NAND U29707 ( .A(n22747), .B(n22748), .Z(n14560) );
  NANDN U29708 ( .A(init), .B(e[817]), .Z(n22748) );
  AND U29709 ( .A(n22749), .B(n22750), .Z(n22747) );
  NAND U29710 ( .A(ereg[816]), .B(n19486), .Z(n22750) );
  NANDN U29711 ( .A(n19481), .B(ereg[817]), .Z(n22749) );
  NAND U29712 ( .A(n22751), .B(n22752), .Z(n14559) );
  NANDN U29713 ( .A(init), .B(e[818]), .Z(n22752) );
  AND U29714 ( .A(n22753), .B(n22754), .Z(n22751) );
  NAND U29715 ( .A(ereg[817]), .B(n19486), .Z(n22754) );
  NANDN U29716 ( .A(n19481), .B(ereg[818]), .Z(n22753) );
  NAND U29717 ( .A(n22755), .B(n22756), .Z(n14558) );
  NANDN U29718 ( .A(init), .B(e[819]), .Z(n22756) );
  AND U29719 ( .A(n22757), .B(n22758), .Z(n22755) );
  NAND U29720 ( .A(ereg[818]), .B(n19486), .Z(n22758) );
  NANDN U29721 ( .A(n19481), .B(ereg[819]), .Z(n22757) );
  NAND U29722 ( .A(n22759), .B(n22760), .Z(n14557) );
  NANDN U29723 ( .A(init), .B(e[820]), .Z(n22760) );
  AND U29724 ( .A(n22761), .B(n22762), .Z(n22759) );
  NAND U29725 ( .A(ereg[819]), .B(n19486), .Z(n22762) );
  NANDN U29726 ( .A(n19481), .B(ereg[820]), .Z(n22761) );
  NAND U29727 ( .A(n22763), .B(n22764), .Z(n14556) );
  NANDN U29728 ( .A(init), .B(e[821]), .Z(n22764) );
  AND U29729 ( .A(n22765), .B(n22766), .Z(n22763) );
  NAND U29730 ( .A(ereg[820]), .B(n19486), .Z(n22766) );
  NANDN U29731 ( .A(n19481), .B(ereg[821]), .Z(n22765) );
  NAND U29732 ( .A(n22767), .B(n22768), .Z(n14555) );
  NANDN U29733 ( .A(init), .B(e[822]), .Z(n22768) );
  AND U29734 ( .A(n22769), .B(n22770), .Z(n22767) );
  NAND U29735 ( .A(ereg[821]), .B(n19486), .Z(n22770) );
  NANDN U29736 ( .A(n19481), .B(ereg[822]), .Z(n22769) );
  NAND U29737 ( .A(n22771), .B(n22772), .Z(n14554) );
  NANDN U29738 ( .A(init), .B(e[823]), .Z(n22772) );
  AND U29739 ( .A(n22773), .B(n22774), .Z(n22771) );
  NAND U29740 ( .A(ereg[822]), .B(n19486), .Z(n22774) );
  NANDN U29741 ( .A(n19481), .B(ereg[823]), .Z(n22773) );
  NAND U29742 ( .A(n22775), .B(n22776), .Z(n14553) );
  NANDN U29743 ( .A(init), .B(e[824]), .Z(n22776) );
  AND U29744 ( .A(n22777), .B(n22778), .Z(n22775) );
  NAND U29745 ( .A(ereg[823]), .B(n19486), .Z(n22778) );
  NANDN U29746 ( .A(n19481), .B(ereg[824]), .Z(n22777) );
  NAND U29747 ( .A(n22779), .B(n22780), .Z(n14552) );
  NANDN U29748 ( .A(init), .B(e[825]), .Z(n22780) );
  AND U29749 ( .A(n22781), .B(n22782), .Z(n22779) );
  NAND U29750 ( .A(ereg[824]), .B(n19486), .Z(n22782) );
  NANDN U29751 ( .A(n19481), .B(ereg[825]), .Z(n22781) );
  NAND U29752 ( .A(n22783), .B(n22784), .Z(n14551) );
  NANDN U29753 ( .A(init), .B(e[826]), .Z(n22784) );
  AND U29754 ( .A(n22785), .B(n22786), .Z(n22783) );
  NAND U29755 ( .A(ereg[825]), .B(n19486), .Z(n22786) );
  NANDN U29756 ( .A(n19481), .B(ereg[826]), .Z(n22785) );
  NAND U29757 ( .A(n22787), .B(n22788), .Z(n14550) );
  NANDN U29758 ( .A(init), .B(e[827]), .Z(n22788) );
  AND U29759 ( .A(n22789), .B(n22790), .Z(n22787) );
  NAND U29760 ( .A(ereg[826]), .B(n19486), .Z(n22790) );
  NANDN U29761 ( .A(n19481), .B(ereg[827]), .Z(n22789) );
  NAND U29762 ( .A(n22791), .B(n22792), .Z(n14549) );
  NANDN U29763 ( .A(init), .B(e[828]), .Z(n22792) );
  AND U29764 ( .A(n22793), .B(n22794), .Z(n22791) );
  NAND U29765 ( .A(ereg[827]), .B(n19486), .Z(n22794) );
  NANDN U29766 ( .A(n19481), .B(ereg[828]), .Z(n22793) );
  NAND U29767 ( .A(n22795), .B(n22796), .Z(n14548) );
  NANDN U29768 ( .A(init), .B(e[829]), .Z(n22796) );
  AND U29769 ( .A(n22797), .B(n22798), .Z(n22795) );
  NAND U29770 ( .A(ereg[828]), .B(n19486), .Z(n22798) );
  NANDN U29771 ( .A(n19481), .B(ereg[829]), .Z(n22797) );
  NAND U29772 ( .A(n22799), .B(n22800), .Z(n14547) );
  NANDN U29773 ( .A(init), .B(e[830]), .Z(n22800) );
  AND U29774 ( .A(n22801), .B(n22802), .Z(n22799) );
  NAND U29775 ( .A(ereg[829]), .B(n19486), .Z(n22802) );
  NANDN U29776 ( .A(n19481), .B(ereg[830]), .Z(n22801) );
  NAND U29777 ( .A(n22803), .B(n22804), .Z(n14546) );
  NANDN U29778 ( .A(init), .B(e[831]), .Z(n22804) );
  AND U29779 ( .A(n22805), .B(n22806), .Z(n22803) );
  NAND U29780 ( .A(ereg[830]), .B(n19486), .Z(n22806) );
  NANDN U29781 ( .A(n19481), .B(ereg[831]), .Z(n22805) );
  NAND U29782 ( .A(n22807), .B(n22808), .Z(n14545) );
  NANDN U29783 ( .A(init), .B(e[832]), .Z(n22808) );
  AND U29784 ( .A(n22809), .B(n22810), .Z(n22807) );
  NAND U29785 ( .A(ereg[831]), .B(n19486), .Z(n22810) );
  NANDN U29786 ( .A(n19481), .B(ereg[832]), .Z(n22809) );
  NAND U29787 ( .A(n22811), .B(n22812), .Z(n14544) );
  NANDN U29788 ( .A(init), .B(e[833]), .Z(n22812) );
  AND U29789 ( .A(n22813), .B(n22814), .Z(n22811) );
  NAND U29790 ( .A(ereg[832]), .B(n19486), .Z(n22814) );
  NANDN U29791 ( .A(n19481), .B(ereg[833]), .Z(n22813) );
  NAND U29792 ( .A(n22815), .B(n22816), .Z(n14543) );
  NANDN U29793 ( .A(init), .B(e[834]), .Z(n22816) );
  AND U29794 ( .A(n22817), .B(n22818), .Z(n22815) );
  NAND U29795 ( .A(ereg[833]), .B(n19486), .Z(n22818) );
  NANDN U29796 ( .A(n19481), .B(ereg[834]), .Z(n22817) );
  NAND U29797 ( .A(n22819), .B(n22820), .Z(n14542) );
  NANDN U29798 ( .A(init), .B(e[835]), .Z(n22820) );
  AND U29799 ( .A(n22821), .B(n22822), .Z(n22819) );
  NAND U29800 ( .A(ereg[834]), .B(n19486), .Z(n22822) );
  NANDN U29801 ( .A(n19481), .B(ereg[835]), .Z(n22821) );
  NAND U29802 ( .A(n22823), .B(n22824), .Z(n14541) );
  NANDN U29803 ( .A(init), .B(e[836]), .Z(n22824) );
  AND U29804 ( .A(n22825), .B(n22826), .Z(n22823) );
  NAND U29805 ( .A(ereg[835]), .B(n19486), .Z(n22826) );
  NANDN U29806 ( .A(n19481), .B(ereg[836]), .Z(n22825) );
  NAND U29807 ( .A(n22827), .B(n22828), .Z(n14540) );
  NANDN U29808 ( .A(init), .B(e[837]), .Z(n22828) );
  AND U29809 ( .A(n22829), .B(n22830), .Z(n22827) );
  NAND U29810 ( .A(ereg[836]), .B(n19486), .Z(n22830) );
  NANDN U29811 ( .A(n19481), .B(ereg[837]), .Z(n22829) );
  NAND U29812 ( .A(n22831), .B(n22832), .Z(n14539) );
  NANDN U29813 ( .A(init), .B(e[838]), .Z(n22832) );
  AND U29814 ( .A(n22833), .B(n22834), .Z(n22831) );
  NAND U29815 ( .A(ereg[837]), .B(n19486), .Z(n22834) );
  NANDN U29816 ( .A(n19481), .B(ereg[838]), .Z(n22833) );
  NAND U29817 ( .A(n22835), .B(n22836), .Z(n14538) );
  NANDN U29818 ( .A(init), .B(e[839]), .Z(n22836) );
  AND U29819 ( .A(n22837), .B(n22838), .Z(n22835) );
  NAND U29820 ( .A(ereg[838]), .B(n19486), .Z(n22838) );
  NANDN U29821 ( .A(n19481), .B(ereg[839]), .Z(n22837) );
  NAND U29822 ( .A(n22839), .B(n22840), .Z(n14537) );
  NANDN U29823 ( .A(init), .B(e[840]), .Z(n22840) );
  AND U29824 ( .A(n22841), .B(n22842), .Z(n22839) );
  NAND U29825 ( .A(ereg[839]), .B(n19486), .Z(n22842) );
  NANDN U29826 ( .A(n19481), .B(ereg[840]), .Z(n22841) );
  NAND U29827 ( .A(n22843), .B(n22844), .Z(n14536) );
  NANDN U29828 ( .A(init), .B(e[841]), .Z(n22844) );
  AND U29829 ( .A(n22845), .B(n22846), .Z(n22843) );
  NAND U29830 ( .A(ereg[840]), .B(n19486), .Z(n22846) );
  NANDN U29831 ( .A(n19481), .B(ereg[841]), .Z(n22845) );
  NAND U29832 ( .A(n22847), .B(n22848), .Z(n14535) );
  NANDN U29833 ( .A(init), .B(e[842]), .Z(n22848) );
  AND U29834 ( .A(n22849), .B(n22850), .Z(n22847) );
  NAND U29835 ( .A(ereg[841]), .B(n19486), .Z(n22850) );
  NANDN U29836 ( .A(n19481), .B(ereg[842]), .Z(n22849) );
  NAND U29837 ( .A(n22851), .B(n22852), .Z(n14534) );
  NANDN U29838 ( .A(init), .B(e[843]), .Z(n22852) );
  AND U29839 ( .A(n22853), .B(n22854), .Z(n22851) );
  NAND U29840 ( .A(ereg[842]), .B(n19486), .Z(n22854) );
  NANDN U29841 ( .A(n19481), .B(ereg[843]), .Z(n22853) );
  NAND U29842 ( .A(n22855), .B(n22856), .Z(n14533) );
  NANDN U29843 ( .A(init), .B(e[844]), .Z(n22856) );
  AND U29844 ( .A(n22857), .B(n22858), .Z(n22855) );
  NAND U29845 ( .A(ereg[843]), .B(n19486), .Z(n22858) );
  NANDN U29846 ( .A(n19481), .B(ereg[844]), .Z(n22857) );
  NAND U29847 ( .A(n22859), .B(n22860), .Z(n14532) );
  NANDN U29848 ( .A(init), .B(e[845]), .Z(n22860) );
  AND U29849 ( .A(n22861), .B(n22862), .Z(n22859) );
  NAND U29850 ( .A(ereg[844]), .B(n19486), .Z(n22862) );
  NANDN U29851 ( .A(n19481), .B(ereg[845]), .Z(n22861) );
  NAND U29852 ( .A(n22863), .B(n22864), .Z(n14531) );
  NANDN U29853 ( .A(init), .B(e[846]), .Z(n22864) );
  AND U29854 ( .A(n22865), .B(n22866), .Z(n22863) );
  NAND U29855 ( .A(ereg[845]), .B(n19486), .Z(n22866) );
  NANDN U29856 ( .A(n19481), .B(ereg[846]), .Z(n22865) );
  NAND U29857 ( .A(n22867), .B(n22868), .Z(n14530) );
  NANDN U29858 ( .A(init), .B(e[847]), .Z(n22868) );
  AND U29859 ( .A(n22869), .B(n22870), .Z(n22867) );
  NAND U29860 ( .A(ereg[846]), .B(n19486), .Z(n22870) );
  NANDN U29861 ( .A(n19481), .B(ereg[847]), .Z(n22869) );
  NAND U29862 ( .A(n22871), .B(n22872), .Z(n14529) );
  NANDN U29863 ( .A(init), .B(e[848]), .Z(n22872) );
  AND U29864 ( .A(n22873), .B(n22874), .Z(n22871) );
  NAND U29865 ( .A(ereg[847]), .B(n19486), .Z(n22874) );
  NANDN U29866 ( .A(n19481), .B(ereg[848]), .Z(n22873) );
  NAND U29867 ( .A(n22875), .B(n22876), .Z(n14528) );
  NANDN U29868 ( .A(init), .B(e[849]), .Z(n22876) );
  AND U29869 ( .A(n22877), .B(n22878), .Z(n22875) );
  NAND U29870 ( .A(ereg[848]), .B(n19486), .Z(n22878) );
  NANDN U29871 ( .A(n19481), .B(ereg[849]), .Z(n22877) );
  NAND U29872 ( .A(n22879), .B(n22880), .Z(n14527) );
  NANDN U29873 ( .A(init), .B(e[850]), .Z(n22880) );
  AND U29874 ( .A(n22881), .B(n22882), .Z(n22879) );
  NAND U29875 ( .A(ereg[849]), .B(n19486), .Z(n22882) );
  NANDN U29876 ( .A(n19481), .B(ereg[850]), .Z(n22881) );
  NAND U29877 ( .A(n22883), .B(n22884), .Z(n14526) );
  NANDN U29878 ( .A(init), .B(e[851]), .Z(n22884) );
  AND U29879 ( .A(n22885), .B(n22886), .Z(n22883) );
  NAND U29880 ( .A(ereg[850]), .B(n19486), .Z(n22886) );
  NANDN U29881 ( .A(n19481), .B(ereg[851]), .Z(n22885) );
  NAND U29882 ( .A(n22887), .B(n22888), .Z(n14525) );
  NANDN U29883 ( .A(init), .B(e[852]), .Z(n22888) );
  AND U29884 ( .A(n22889), .B(n22890), .Z(n22887) );
  NAND U29885 ( .A(ereg[851]), .B(n19486), .Z(n22890) );
  NANDN U29886 ( .A(n19481), .B(ereg[852]), .Z(n22889) );
  NAND U29887 ( .A(n22891), .B(n22892), .Z(n14524) );
  NANDN U29888 ( .A(init), .B(e[853]), .Z(n22892) );
  AND U29889 ( .A(n22893), .B(n22894), .Z(n22891) );
  NAND U29890 ( .A(ereg[852]), .B(n19486), .Z(n22894) );
  NANDN U29891 ( .A(n19481), .B(ereg[853]), .Z(n22893) );
  NAND U29892 ( .A(n22895), .B(n22896), .Z(n14523) );
  NANDN U29893 ( .A(init), .B(e[854]), .Z(n22896) );
  AND U29894 ( .A(n22897), .B(n22898), .Z(n22895) );
  NAND U29895 ( .A(ereg[853]), .B(n19486), .Z(n22898) );
  NANDN U29896 ( .A(n19481), .B(ereg[854]), .Z(n22897) );
  NAND U29897 ( .A(n22899), .B(n22900), .Z(n14522) );
  NANDN U29898 ( .A(init), .B(e[855]), .Z(n22900) );
  AND U29899 ( .A(n22901), .B(n22902), .Z(n22899) );
  NAND U29900 ( .A(ereg[854]), .B(n19486), .Z(n22902) );
  NANDN U29901 ( .A(n19481), .B(ereg[855]), .Z(n22901) );
  NAND U29902 ( .A(n22903), .B(n22904), .Z(n14521) );
  NANDN U29903 ( .A(init), .B(e[856]), .Z(n22904) );
  AND U29904 ( .A(n22905), .B(n22906), .Z(n22903) );
  NAND U29905 ( .A(ereg[855]), .B(n19486), .Z(n22906) );
  NANDN U29906 ( .A(n19481), .B(ereg[856]), .Z(n22905) );
  NAND U29907 ( .A(n22907), .B(n22908), .Z(n14520) );
  NANDN U29908 ( .A(init), .B(e[857]), .Z(n22908) );
  AND U29909 ( .A(n22909), .B(n22910), .Z(n22907) );
  NAND U29910 ( .A(ereg[856]), .B(n19486), .Z(n22910) );
  NANDN U29911 ( .A(n19481), .B(ereg[857]), .Z(n22909) );
  NAND U29912 ( .A(n22911), .B(n22912), .Z(n14519) );
  NANDN U29913 ( .A(init), .B(e[858]), .Z(n22912) );
  AND U29914 ( .A(n22913), .B(n22914), .Z(n22911) );
  NAND U29915 ( .A(ereg[857]), .B(n19486), .Z(n22914) );
  NANDN U29916 ( .A(n19481), .B(ereg[858]), .Z(n22913) );
  NAND U29917 ( .A(n22915), .B(n22916), .Z(n14518) );
  NANDN U29918 ( .A(init), .B(e[859]), .Z(n22916) );
  AND U29919 ( .A(n22917), .B(n22918), .Z(n22915) );
  NAND U29920 ( .A(ereg[858]), .B(n19486), .Z(n22918) );
  NANDN U29921 ( .A(n19481), .B(ereg[859]), .Z(n22917) );
  NAND U29922 ( .A(n22919), .B(n22920), .Z(n14517) );
  NANDN U29923 ( .A(init), .B(e[860]), .Z(n22920) );
  AND U29924 ( .A(n22921), .B(n22922), .Z(n22919) );
  NAND U29925 ( .A(ereg[859]), .B(n19486), .Z(n22922) );
  NANDN U29926 ( .A(n19481), .B(ereg[860]), .Z(n22921) );
  NAND U29927 ( .A(n22923), .B(n22924), .Z(n14516) );
  NANDN U29928 ( .A(init), .B(e[861]), .Z(n22924) );
  AND U29929 ( .A(n22925), .B(n22926), .Z(n22923) );
  NAND U29930 ( .A(ereg[860]), .B(n19486), .Z(n22926) );
  NANDN U29931 ( .A(n19481), .B(ereg[861]), .Z(n22925) );
  NAND U29932 ( .A(n22927), .B(n22928), .Z(n14515) );
  NANDN U29933 ( .A(init), .B(e[862]), .Z(n22928) );
  AND U29934 ( .A(n22929), .B(n22930), .Z(n22927) );
  NAND U29935 ( .A(ereg[861]), .B(n19486), .Z(n22930) );
  NANDN U29936 ( .A(n19481), .B(ereg[862]), .Z(n22929) );
  NAND U29937 ( .A(n22931), .B(n22932), .Z(n14514) );
  NANDN U29938 ( .A(init), .B(e[863]), .Z(n22932) );
  AND U29939 ( .A(n22933), .B(n22934), .Z(n22931) );
  NAND U29940 ( .A(ereg[862]), .B(n19486), .Z(n22934) );
  NANDN U29941 ( .A(n19481), .B(ereg[863]), .Z(n22933) );
  NAND U29942 ( .A(n22935), .B(n22936), .Z(n14513) );
  NANDN U29943 ( .A(init), .B(e[864]), .Z(n22936) );
  AND U29944 ( .A(n22937), .B(n22938), .Z(n22935) );
  NAND U29945 ( .A(ereg[863]), .B(n19486), .Z(n22938) );
  NANDN U29946 ( .A(n19481), .B(ereg[864]), .Z(n22937) );
  NAND U29947 ( .A(n22939), .B(n22940), .Z(n14512) );
  NANDN U29948 ( .A(init), .B(e[865]), .Z(n22940) );
  AND U29949 ( .A(n22941), .B(n22942), .Z(n22939) );
  NAND U29950 ( .A(ereg[864]), .B(n19486), .Z(n22942) );
  NANDN U29951 ( .A(n19481), .B(ereg[865]), .Z(n22941) );
  NAND U29952 ( .A(n22943), .B(n22944), .Z(n14511) );
  NANDN U29953 ( .A(init), .B(e[866]), .Z(n22944) );
  AND U29954 ( .A(n22945), .B(n22946), .Z(n22943) );
  NAND U29955 ( .A(ereg[865]), .B(n19486), .Z(n22946) );
  NANDN U29956 ( .A(n19481), .B(ereg[866]), .Z(n22945) );
  NAND U29957 ( .A(n22947), .B(n22948), .Z(n14510) );
  NANDN U29958 ( .A(init), .B(e[867]), .Z(n22948) );
  AND U29959 ( .A(n22949), .B(n22950), .Z(n22947) );
  NAND U29960 ( .A(ereg[866]), .B(n19486), .Z(n22950) );
  NANDN U29961 ( .A(n19481), .B(ereg[867]), .Z(n22949) );
  NAND U29962 ( .A(n22951), .B(n22952), .Z(n14509) );
  NANDN U29963 ( .A(init), .B(e[868]), .Z(n22952) );
  AND U29964 ( .A(n22953), .B(n22954), .Z(n22951) );
  NAND U29965 ( .A(ereg[867]), .B(n19486), .Z(n22954) );
  NANDN U29966 ( .A(n19481), .B(ereg[868]), .Z(n22953) );
  NAND U29967 ( .A(n22955), .B(n22956), .Z(n14508) );
  NANDN U29968 ( .A(init), .B(e[869]), .Z(n22956) );
  AND U29969 ( .A(n22957), .B(n22958), .Z(n22955) );
  NAND U29970 ( .A(ereg[868]), .B(n19486), .Z(n22958) );
  NANDN U29971 ( .A(n19481), .B(ereg[869]), .Z(n22957) );
  NAND U29972 ( .A(n22959), .B(n22960), .Z(n14507) );
  NANDN U29973 ( .A(init), .B(e[870]), .Z(n22960) );
  AND U29974 ( .A(n22961), .B(n22962), .Z(n22959) );
  NAND U29975 ( .A(ereg[869]), .B(n19486), .Z(n22962) );
  NANDN U29976 ( .A(n19481), .B(ereg[870]), .Z(n22961) );
  NAND U29977 ( .A(n22963), .B(n22964), .Z(n14506) );
  NANDN U29978 ( .A(init), .B(e[871]), .Z(n22964) );
  AND U29979 ( .A(n22965), .B(n22966), .Z(n22963) );
  NAND U29980 ( .A(ereg[870]), .B(n19486), .Z(n22966) );
  NANDN U29981 ( .A(n19481), .B(ereg[871]), .Z(n22965) );
  NAND U29982 ( .A(n22967), .B(n22968), .Z(n14505) );
  NANDN U29983 ( .A(init), .B(e[872]), .Z(n22968) );
  AND U29984 ( .A(n22969), .B(n22970), .Z(n22967) );
  NAND U29985 ( .A(ereg[871]), .B(n19486), .Z(n22970) );
  NANDN U29986 ( .A(n19481), .B(ereg[872]), .Z(n22969) );
  NAND U29987 ( .A(n22971), .B(n22972), .Z(n14504) );
  NANDN U29988 ( .A(init), .B(e[873]), .Z(n22972) );
  AND U29989 ( .A(n22973), .B(n22974), .Z(n22971) );
  NAND U29990 ( .A(ereg[872]), .B(n19486), .Z(n22974) );
  NANDN U29991 ( .A(n19481), .B(ereg[873]), .Z(n22973) );
  NAND U29992 ( .A(n22975), .B(n22976), .Z(n14503) );
  NANDN U29993 ( .A(init), .B(e[874]), .Z(n22976) );
  AND U29994 ( .A(n22977), .B(n22978), .Z(n22975) );
  NAND U29995 ( .A(ereg[873]), .B(n19486), .Z(n22978) );
  NANDN U29996 ( .A(n19481), .B(ereg[874]), .Z(n22977) );
  NAND U29997 ( .A(n22979), .B(n22980), .Z(n14502) );
  NANDN U29998 ( .A(init), .B(e[875]), .Z(n22980) );
  AND U29999 ( .A(n22981), .B(n22982), .Z(n22979) );
  NAND U30000 ( .A(ereg[874]), .B(n19486), .Z(n22982) );
  NANDN U30001 ( .A(n19481), .B(ereg[875]), .Z(n22981) );
  NAND U30002 ( .A(n22983), .B(n22984), .Z(n14501) );
  NANDN U30003 ( .A(init), .B(e[876]), .Z(n22984) );
  AND U30004 ( .A(n22985), .B(n22986), .Z(n22983) );
  NAND U30005 ( .A(ereg[875]), .B(n19486), .Z(n22986) );
  NANDN U30006 ( .A(n19481), .B(ereg[876]), .Z(n22985) );
  NAND U30007 ( .A(n22987), .B(n22988), .Z(n14500) );
  NANDN U30008 ( .A(init), .B(e[877]), .Z(n22988) );
  AND U30009 ( .A(n22989), .B(n22990), .Z(n22987) );
  NAND U30010 ( .A(ereg[876]), .B(n19486), .Z(n22990) );
  NANDN U30011 ( .A(n19481), .B(ereg[877]), .Z(n22989) );
  NAND U30012 ( .A(n22991), .B(n22992), .Z(n14499) );
  NANDN U30013 ( .A(init), .B(e[878]), .Z(n22992) );
  AND U30014 ( .A(n22993), .B(n22994), .Z(n22991) );
  NAND U30015 ( .A(ereg[877]), .B(n19486), .Z(n22994) );
  NANDN U30016 ( .A(n19481), .B(ereg[878]), .Z(n22993) );
  NAND U30017 ( .A(n22995), .B(n22996), .Z(n14498) );
  NANDN U30018 ( .A(init), .B(e[879]), .Z(n22996) );
  AND U30019 ( .A(n22997), .B(n22998), .Z(n22995) );
  NAND U30020 ( .A(ereg[878]), .B(n19486), .Z(n22998) );
  NANDN U30021 ( .A(n19481), .B(ereg[879]), .Z(n22997) );
  NAND U30022 ( .A(n22999), .B(n23000), .Z(n14497) );
  NANDN U30023 ( .A(init), .B(e[880]), .Z(n23000) );
  AND U30024 ( .A(n23001), .B(n23002), .Z(n22999) );
  NAND U30025 ( .A(ereg[879]), .B(n19486), .Z(n23002) );
  NANDN U30026 ( .A(n19481), .B(ereg[880]), .Z(n23001) );
  NAND U30027 ( .A(n23003), .B(n23004), .Z(n14496) );
  NANDN U30028 ( .A(init), .B(e[881]), .Z(n23004) );
  AND U30029 ( .A(n23005), .B(n23006), .Z(n23003) );
  NAND U30030 ( .A(ereg[880]), .B(n19486), .Z(n23006) );
  NANDN U30031 ( .A(n19481), .B(ereg[881]), .Z(n23005) );
  NAND U30032 ( .A(n23007), .B(n23008), .Z(n14495) );
  NANDN U30033 ( .A(init), .B(e[882]), .Z(n23008) );
  AND U30034 ( .A(n23009), .B(n23010), .Z(n23007) );
  NAND U30035 ( .A(ereg[881]), .B(n19486), .Z(n23010) );
  NANDN U30036 ( .A(n19481), .B(ereg[882]), .Z(n23009) );
  NAND U30037 ( .A(n23011), .B(n23012), .Z(n14494) );
  NANDN U30038 ( .A(init), .B(e[883]), .Z(n23012) );
  AND U30039 ( .A(n23013), .B(n23014), .Z(n23011) );
  NAND U30040 ( .A(ereg[882]), .B(n19486), .Z(n23014) );
  NANDN U30041 ( .A(n19481), .B(ereg[883]), .Z(n23013) );
  NAND U30042 ( .A(n23015), .B(n23016), .Z(n14493) );
  NANDN U30043 ( .A(init), .B(e[884]), .Z(n23016) );
  AND U30044 ( .A(n23017), .B(n23018), .Z(n23015) );
  NAND U30045 ( .A(ereg[883]), .B(n19486), .Z(n23018) );
  NANDN U30046 ( .A(n19481), .B(ereg[884]), .Z(n23017) );
  NAND U30047 ( .A(n23019), .B(n23020), .Z(n14492) );
  NANDN U30048 ( .A(init), .B(e[885]), .Z(n23020) );
  AND U30049 ( .A(n23021), .B(n23022), .Z(n23019) );
  NAND U30050 ( .A(ereg[884]), .B(n19486), .Z(n23022) );
  NANDN U30051 ( .A(n19481), .B(ereg[885]), .Z(n23021) );
  NAND U30052 ( .A(n23023), .B(n23024), .Z(n14491) );
  NANDN U30053 ( .A(init), .B(e[886]), .Z(n23024) );
  AND U30054 ( .A(n23025), .B(n23026), .Z(n23023) );
  NAND U30055 ( .A(ereg[885]), .B(n19486), .Z(n23026) );
  NANDN U30056 ( .A(n19481), .B(ereg[886]), .Z(n23025) );
  NAND U30057 ( .A(n23027), .B(n23028), .Z(n14490) );
  NANDN U30058 ( .A(init), .B(e[887]), .Z(n23028) );
  AND U30059 ( .A(n23029), .B(n23030), .Z(n23027) );
  NAND U30060 ( .A(ereg[886]), .B(n19486), .Z(n23030) );
  NANDN U30061 ( .A(n19481), .B(ereg[887]), .Z(n23029) );
  NAND U30062 ( .A(n23031), .B(n23032), .Z(n14489) );
  NANDN U30063 ( .A(init), .B(e[888]), .Z(n23032) );
  AND U30064 ( .A(n23033), .B(n23034), .Z(n23031) );
  NAND U30065 ( .A(ereg[887]), .B(n19486), .Z(n23034) );
  NANDN U30066 ( .A(n19481), .B(ereg[888]), .Z(n23033) );
  NAND U30067 ( .A(n23035), .B(n23036), .Z(n14488) );
  NANDN U30068 ( .A(init), .B(e[889]), .Z(n23036) );
  AND U30069 ( .A(n23037), .B(n23038), .Z(n23035) );
  NAND U30070 ( .A(ereg[888]), .B(n19486), .Z(n23038) );
  NANDN U30071 ( .A(n19481), .B(ereg[889]), .Z(n23037) );
  NAND U30072 ( .A(n23039), .B(n23040), .Z(n14487) );
  NANDN U30073 ( .A(init), .B(e[890]), .Z(n23040) );
  AND U30074 ( .A(n23041), .B(n23042), .Z(n23039) );
  NAND U30075 ( .A(ereg[889]), .B(n19486), .Z(n23042) );
  NANDN U30076 ( .A(n19481), .B(ereg[890]), .Z(n23041) );
  NAND U30077 ( .A(n23043), .B(n23044), .Z(n14486) );
  NANDN U30078 ( .A(init), .B(e[891]), .Z(n23044) );
  AND U30079 ( .A(n23045), .B(n23046), .Z(n23043) );
  NAND U30080 ( .A(ereg[890]), .B(n19486), .Z(n23046) );
  NANDN U30081 ( .A(n19481), .B(ereg[891]), .Z(n23045) );
  NAND U30082 ( .A(n23047), .B(n23048), .Z(n14485) );
  NANDN U30083 ( .A(init), .B(e[892]), .Z(n23048) );
  AND U30084 ( .A(n23049), .B(n23050), .Z(n23047) );
  NAND U30085 ( .A(ereg[891]), .B(n19486), .Z(n23050) );
  NANDN U30086 ( .A(n19481), .B(ereg[892]), .Z(n23049) );
  NAND U30087 ( .A(n23051), .B(n23052), .Z(n14484) );
  NANDN U30088 ( .A(init), .B(e[893]), .Z(n23052) );
  AND U30089 ( .A(n23053), .B(n23054), .Z(n23051) );
  NAND U30090 ( .A(ereg[892]), .B(n19486), .Z(n23054) );
  NANDN U30091 ( .A(n19481), .B(ereg[893]), .Z(n23053) );
  NAND U30092 ( .A(n23055), .B(n23056), .Z(n14483) );
  NANDN U30093 ( .A(init), .B(e[894]), .Z(n23056) );
  AND U30094 ( .A(n23057), .B(n23058), .Z(n23055) );
  NAND U30095 ( .A(ereg[893]), .B(n19486), .Z(n23058) );
  NANDN U30096 ( .A(n19481), .B(ereg[894]), .Z(n23057) );
  NAND U30097 ( .A(n23059), .B(n23060), .Z(n14482) );
  NANDN U30098 ( .A(init), .B(e[895]), .Z(n23060) );
  AND U30099 ( .A(n23061), .B(n23062), .Z(n23059) );
  NAND U30100 ( .A(ereg[894]), .B(n19486), .Z(n23062) );
  NANDN U30101 ( .A(n19481), .B(ereg[895]), .Z(n23061) );
  NAND U30102 ( .A(n23063), .B(n23064), .Z(n14481) );
  NANDN U30103 ( .A(init), .B(e[896]), .Z(n23064) );
  AND U30104 ( .A(n23065), .B(n23066), .Z(n23063) );
  NAND U30105 ( .A(ereg[895]), .B(n19486), .Z(n23066) );
  NANDN U30106 ( .A(n19481), .B(ereg[896]), .Z(n23065) );
  NAND U30107 ( .A(n23067), .B(n23068), .Z(n14480) );
  NANDN U30108 ( .A(init), .B(e[897]), .Z(n23068) );
  AND U30109 ( .A(n23069), .B(n23070), .Z(n23067) );
  NAND U30110 ( .A(ereg[896]), .B(n19486), .Z(n23070) );
  NANDN U30111 ( .A(n19481), .B(ereg[897]), .Z(n23069) );
  NAND U30112 ( .A(n23071), .B(n23072), .Z(n14479) );
  NANDN U30113 ( .A(init), .B(e[898]), .Z(n23072) );
  AND U30114 ( .A(n23073), .B(n23074), .Z(n23071) );
  NAND U30115 ( .A(ereg[897]), .B(n19486), .Z(n23074) );
  NANDN U30116 ( .A(n19481), .B(ereg[898]), .Z(n23073) );
  NAND U30117 ( .A(n23075), .B(n23076), .Z(n14478) );
  NANDN U30118 ( .A(init), .B(e[899]), .Z(n23076) );
  AND U30119 ( .A(n23077), .B(n23078), .Z(n23075) );
  NAND U30120 ( .A(ereg[898]), .B(n19486), .Z(n23078) );
  NANDN U30121 ( .A(n19481), .B(ereg[899]), .Z(n23077) );
  NAND U30122 ( .A(n23079), .B(n23080), .Z(n14477) );
  NANDN U30123 ( .A(init), .B(e[900]), .Z(n23080) );
  AND U30124 ( .A(n23081), .B(n23082), .Z(n23079) );
  NAND U30125 ( .A(ereg[899]), .B(n19486), .Z(n23082) );
  NANDN U30126 ( .A(n19481), .B(ereg[900]), .Z(n23081) );
  NAND U30127 ( .A(n23083), .B(n23084), .Z(n14476) );
  NANDN U30128 ( .A(init), .B(e[901]), .Z(n23084) );
  AND U30129 ( .A(n23085), .B(n23086), .Z(n23083) );
  NAND U30130 ( .A(ereg[900]), .B(n19486), .Z(n23086) );
  NANDN U30131 ( .A(n19481), .B(ereg[901]), .Z(n23085) );
  NAND U30132 ( .A(n23087), .B(n23088), .Z(n14475) );
  NANDN U30133 ( .A(init), .B(e[902]), .Z(n23088) );
  AND U30134 ( .A(n23089), .B(n23090), .Z(n23087) );
  NAND U30135 ( .A(ereg[901]), .B(n19486), .Z(n23090) );
  NANDN U30136 ( .A(n19481), .B(ereg[902]), .Z(n23089) );
  NAND U30137 ( .A(n23091), .B(n23092), .Z(n14474) );
  NANDN U30138 ( .A(init), .B(e[903]), .Z(n23092) );
  AND U30139 ( .A(n23093), .B(n23094), .Z(n23091) );
  NAND U30140 ( .A(ereg[902]), .B(n19486), .Z(n23094) );
  NANDN U30141 ( .A(n19481), .B(ereg[903]), .Z(n23093) );
  NAND U30142 ( .A(n23095), .B(n23096), .Z(n14473) );
  NANDN U30143 ( .A(init), .B(e[904]), .Z(n23096) );
  AND U30144 ( .A(n23097), .B(n23098), .Z(n23095) );
  NAND U30145 ( .A(ereg[903]), .B(n19486), .Z(n23098) );
  NANDN U30146 ( .A(n19481), .B(ereg[904]), .Z(n23097) );
  NAND U30147 ( .A(n23099), .B(n23100), .Z(n14472) );
  NANDN U30148 ( .A(init), .B(e[905]), .Z(n23100) );
  AND U30149 ( .A(n23101), .B(n23102), .Z(n23099) );
  NAND U30150 ( .A(ereg[904]), .B(n19486), .Z(n23102) );
  NANDN U30151 ( .A(n19481), .B(ereg[905]), .Z(n23101) );
  NAND U30152 ( .A(n23103), .B(n23104), .Z(n14471) );
  NANDN U30153 ( .A(init), .B(e[906]), .Z(n23104) );
  AND U30154 ( .A(n23105), .B(n23106), .Z(n23103) );
  NAND U30155 ( .A(ereg[905]), .B(n19486), .Z(n23106) );
  NANDN U30156 ( .A(n19481), .B(ereg[906]), .Z(n23105) );
  NAND U30157 ( .A(n23107), .B(n23108), .Z(n14470) );
  NANDN U30158 ( .A(init), .B(e[907]), .Z(n23108) );
  AND U30159 ( .A(n23109), .B(n23110), .Z(n23107) );
  NAND U30160 ( .A(ereg[906]), .B(n19486), .Z(n23110) );
  NANDN U30161 ( .A(n19481), .B(ereg[907]), .Z(n23109) );
  NAND U30162 ( .A(n23111), .B(n23112), .Z(n14469) );
  NANDN U30163 ( .A(init), .B(e[908]), .Z(n23112) );
  AND U30164 ( .A(n23113), .B(n23114), .Z(n23111) );
  NAND U30165 ( .A(ereg[907]), .B(n19486), .Z(n23114) );
  NANDN U30166 ( .A(n19481), .B(ereg[908]), .Z(n23113) );
  NAND U30167 ( .A(n23115), .B(n23116), .Z(n14468) );
  NANDN U30168 ( .A(init), .B(e[909]), .Z(n23116) );
  AND U30169 ( .A(n23117), .B(n23118), .Z(n23115) );
  NAND U30170 ( .A(ereg[908]), .B(n19486), .Z(n23118) );
  NANDN U30171 ( .A(n19481), .B(ereg[909]), .Z(n23117) );
  NAND U30172 ( .A(n23119), .B(n23120), .Z(n14467) );
  NANDN U30173 ( .A(init), .B(e[910]), .Z(n23120) );
  AND U30174 ( .A(n23121), .B(n23122), .Z(n23119) );
  NAND U30175 ( .A(ereg[909]), .B(n19486), .Z(n23122) );
  NANDN U30176 ( .A(n19481), .B(ereg[910]), .Z(n23121) );
  NAND U30177 ( .A(n23123), .B(n23124), .Z(n14466) );
  NANDN U30178 ( .A(init), .B(e[911]), .Z(n23124) );
  AND U30179 ( .A(n23125), .B(n23126), .Z(n23123) );
  NAND U30180 ( .A(ereg[910]), .B(n19486), .Z(n23126) );
  NANDN U30181 ( .A(n19481), .B(ereg[911]), .Z(n23125) );
  NAND U30182 ( .A(n23127), .B(n23128), .Z(n14465) );
  NANDN U30183 ( .A(init), .B(e[912]), .Z(n23128) );
  AND U30184 ( .A(n23129), .B(n23130), .Z(n23127) );
  NAND U30185 ( .A(ereg[911]), .B(n19486), .Z(n23130) );
  NANDN U30186 ( .A(n19481), .B(ereg[912]), .Z(n23129) );
  NAND U30187 ( .A(n23131), .B(n23132), .Z(n14464) );
  NANDN U30188 ( .A(init), .B(e[913]), .Z(n23132) );
  AND U30189 ( .A(n23133), .B(n23134), .Z(n23131) );
  NAND U30190 ( .A(ereg[912]), .B(n19486), .Z(n23134) );
  NANDN U30191 ( .A(n19481), .B(ereg[913]), .Z(n23133) );
  NAND U30192 ( .A(n23135), .B(n23136), .Z(n14463) );
  NANDN U30193 ( .A(init), .B(e[914]), .Z(n23136) );
  AND U30194 ( .A(n23137), .B(n23138), .Z(n23135) );
  NAND U30195 ( .A(ereg[913]), .B(n19486), .Z(n23138) );
  NANDN U30196 ( .A(n19481), .B(ereg[914]), .Z(n23137) );
  NAND U30197 ( .A(n23139), .B(n23140), .Z(n14462) );
  NANDN U30198 ( .A(init), .B(e[915]), .Z(n23140) );
  AND U30199 ( .A(n23141), .B(n23142), .Z(n23139) );
  NAND U30200 ( .A(ereg[914]), .B(n19486), .Z(n23142) );
  NANDN U30201 ( .A(n19481), .B(ereg[915]), .Z(n23141) );
  NAND U30202 ( .A(n23143), .B(n23144), .Z(n14461) );
  NANDN U30203 ( .A(init), .B(e[916]), .Z(n23144) );
  AND U30204 ( .A(n23145), .B(n23146), .Z(n23143) );
  NAND U30205 ( .A(ereg[915]), .B(n19486), .Z(n23146) );
  NANDN U30206 ( .A(n19481), .B(ereg[916]), .Z(n23145) );
  NAND U30207 ( .A(n23147), .B(n23148), .Z(n14460) );
  NANDN U30208 ( .A(init), .B(e[917]), .Z(n23148) );
  AND U30209 ( .A(n23149), .B(n23150), .Z(n23147) );
  NAND U30210 ( .A(ereg[916]), .B(n19486), .Z(n23150) );
  NANDN U30211 ( .A(n19481), .B(ereg[917]), .Z(n23149) );
  NAND U30212 ( .A(n23151), .B(n23152), .Z(n14459) );
  NANDN U30213 ( .A(init), .B(e[918]), .Z(n23152) );
  AND U30214 ( .A(n23153), .B(n23154), .Z(n23151) );
  NAND U30215 ( .A(ereg[917]), .B(n19486), .Z(n23154) );
  NANDN U30216 ( .A(n19481), .B(ereg[918]), .Z(n23153) );
  NAND U30217 ( .A(n23155), .B(n23156), .Z(n14458) );
  NANDN U30218 ( .A(init), .B(e[919]), .Z(n23156) );
  AND U30219 ( .A(n23157), .B(n23158), .Z(n23155) );
  NAND U30220 ( .A(ereg[918]), .B(n19486), .Z(n23158) );
  NANDN U30221 ( .A(n19481), .B(ereg[919]), .Z(n23157) );
  NAND U30222 ( .A(n23159), .B(n23160), .Z(n14457) );
  NANDN U30223 ( .A(init), .B(e[920]), .Z(n23160) );
  AND U30224 ( .A(n23161), .B(n23162), .Z(n23159) );
  NAND U30225 ( .A(ereg[919]), .B(n19486), .Z(n23162) );
  NANDN U30226 ( .A(n19481), .B(ereg[920]), .Z(n23161) );
  NAND U30227 ( .A(n23163), .B(n23164), .Z(n14456) );
  NANDN U30228 ( .A(init), .B(e[921]), .Z(n23164) );
  AND U30229 ( .A(n23165), .B(n23166), .Z(n23163) );
  NAND U30230 ( .A(ereg[920]), .B(n19486), .Z(n23166) );
  NANDN U30231 ( .A(n19481), .B(ereg[921]), .Z(n23165) );
  NAND U30232 ( .A(n23167), .B(n23168), .Z(n14455) );
  NANDN U30233 ( .A(init), .B(e[922]), .Z(n23168) );
  AND U30234 ( .A(n23169), .B(n23170), .Z(n23167) );
  NAND U30235 ( .A(ereg[921]), .B(n19486), .Z(n23170) );
  NANDN U30236 ( .A(n19481), .B(ereg[922]), .Z(n23169) );
  NAND U30237 ( .A(n23171), .B(n23172), .Z(n14454) );
  NANDN U30238 ( .A(init), .B(e[923]), .Z(n23172) );
  AND U30239 ( .A(n23173), .B(n23174), .Z(n23171) );
  NAND U30240 ( .A(ereg[922]), .B(n19486), .Z(n23174) );
  NANDN U30241 ( .A(n19481), .B(ereg[923]), .Z(n23173) );
  NAND U30242 ( .A(n23175), .B(n23176), .Z(n14453) );
  NANDN U30243 ( .A(init), .B(e[924]), .Z(n23176) );
  AND U30244 ( .A(n23177), .B(n23178), .Z(n23175) );
  NAND U30245 ( .A(ereg[923]), .B(n19486), .Z(n23178) );
  NANDN U30246 ( .A(n19481), .B(ereg[924]), .Z(n23177) );
  NAND U30247 ( .A(n23179), .B(n23180), .Z(n14452) );
  NANDN U30248 ( .A(init), .B(e[925]), .Z(n23180) );
  AND U30249 ( .A(n23181), .B(n23182), .Z(n23179) );
  NAND U30250 ( .A(ereg[924]), .B(n19486), .Z(n23182) );
  NANDN U30251 ( .A(n19481), .B(ereg[925]), .Z(n23181) );
  NAND U30252 ( .A(n23183), .B(n23184), .Z(n14451) );
  NANDN U30253 ( .A(init), .B(e[926]), .Z(n23184) );
  AND U30254 ( .A(n23185), .B(n23186), .Z(n23183) );
  NAND U30255 ( .A(ereg[925]), .B(n19486), .Z(n23186) );
  NANDN U30256 ( .A(n19481), .B(ereg[926]), .Z(n23185) );
  NAND U30257 ( .A(n23187), .B(n23188), .Z(n14450) );
  NANDN U30258 ( .A(init), .B(e[927]), .Z(n23188) );
  AND U30259 ( .A(n23189), .B(n23190), .Z(n23187) );
  NAND U30260 ( .A(ereg[926]), .B(n19486), .Z(n23190) );
  NANDN U30261 ( .A(n19481), .B(ereg[927]), .Z(n23189) );
  NAND U30262 ( .A(n23191), .B(n23192), .Z(n14449) );
  NANDN U30263 ( .A(init), .B(e[928]), .Z(n23192) );
  AND U30264 ( .A(n23193), .B(n23194), .Z(n23191) );
  NAND U30265 ( .A(ereg[927]), .B(n19486), .Z(n23194) );
  NANDN U30266 ( .A(n19481), .B(ereg[928]), .Z(n23193) );
  NAND U30267 ( .A(n23195), .B(n23196), .Z(n14448) );
  NANDN U30268 ( .A(init), .B(e[929]), .Z(n23196) );
  AND U30269 ( .A(n23197), .B(n23198), .Z(n23195) );
  NAND U30270 ( .A(ereg[928]), .B(n19486), .Z(n23198) );
  NANDN U30271 ( .A(n19481), .B(ereg[929]), .Z(n23197) );
  NAND U30272 ( .A(n23199), .B(n23200), .Z(n14447) );
  NANDN U30273 ( .A(init), .B(e[930]), .Z(n23200) );
  AND U30274 ( .A(n23201), .B(n23202), .Z(n23199) );
  NAND U30275 ( .A(ereg[929]), .B(n19486), .Z(n23202) );
  NANDN U30276 ( .A(n19481), .B(ereg[930]), .Z(n23201) );
  NAND U30277 ( .A(n23203), .B(n23204), .Z(n14446) );
  NANDN U30278 ( .A(init), .B(e[931]), .Z(n23204) );
  AND U30279 ( .A(n23205), .B(n23206), .Z(n23203) );
  NAND U30280 ( .A(ereg[930]), .B(n19486), .Z(n23206) );
  NANDN U30281 ( .A(n19481), .B(ereg[931]), .Z(n23205) );
  NAND U30282 ( .A(n23207), .B(n23208), .Z(n14445) );
  NANDN U30283 ( .A(init), .B(e[932]), .Z(n23208) );
  AND U30284 ( .A(n23209), .B(n23210), .Z(n23207) );
  NAND U30285 ( .A(ereg[931]), .B(n19486), .Z(n23210) );
  NANDN U30286 ( .A(n19481), .B(ereg[932]), .Z(n23209) );
  NAND U30287 ( .A(n23211), .B(n23212), .Z(n14444) );
  NANDN U30288 ( .A(init), .B(e[933]), .Z(n23212) );
  AND U30289 ( .A(n23213), .B(n23214), .Z(n23211) );
  NAND U30290 ( .A(ereg[932]), .B(n19486), .Z(n23214) );
  NANDN U30291 ( .A(n19481), .B(ereg[933]), .Z(n23213) );
  NAND U30292 ( .A(n23215), .B(n23216), .Z(n14443) );
  NANDN U30293 ( .A(init), .B(e[934]), .Z(n23216) );
  AND U30294 ( .A(n23217), .B(n23218), .Z(n23215) );
  NAND U30295 ( .A(ereg[933]), .B(n19486), .Z(n23218) );
  NANDN U30296 ( .A(n19481), .B(ereg[934]), .Z(n23217) );
  NAND U30297 ( .A(n23219), .B(n23220), .Z(n14442) );
  NANDN U30298 ( .A(init), .B(e[935]), .Z(n23220) );
  AND U30299 ( .A(n23221), .B(n23222), .Z(n23219) );
  NAND U30300 ( .A(ereg[934]), .B(n19486), .Z(n23222) );
  NANDN U30301 ( .A(n19481), .B(ereg[935]), .Z(n23221) );
  NAND U30302 ( .A(n23223), .B(n23224), .Z(n14441) );
  NANDN U30303 ( .A(init), .B(e[936]), .Z(n23224) );
  AND U30304 ( .A(n23225), .B(n23226), .Z(n23223) );
  NAND U30305 ( .A(ereg[935]), .B(n19486), .Z(n23226) );
  NANDN U30306 ( .A(n19481), .B(ereg[936]), .Z(n23225) );
  NAND U30307 ( .A(n23227), .B(n23228), .Z(n14440) );
  NANDN U30308 ( .A(init), .B(e[937]), .Z(n23228) );
  AND U30309 ( .A(n23229), .B(n23230), .Z(n23227) );
  NAND U30310 ( .A(ereg[936]), .B(n19486), .Z(n23230) );
  NANDN U30311 ( .A(n19481), .B(ereg[937]), .Z(n23229) );
  NAND U30312 ( .A(n23231), .B(n23232), .Z(n14439) );
  NANDN U30313 ( .A(init), .B(e[938]), .Z(n23232) );
  AND U30314 ( .A(n23233), .B(n23234), .Z(n23231) );
  NAND U30315 ( .A(ereg[937]), .B(n19486), .Z(n23234) );
  NANDN U30316 ( .A(n19481), .B(ereg[938]), .Z(n23233) );
  NAND U30317 ( .A(n23235), .B(n23236), .Z(n14438) );
  NANDN U30318 ( .A(init), .B(e[939]), .Z(n23236) );
  AND U30319 ( .A(n23237), .B(n23238), .Z(n23235) );
  NAND U30320 ( .A(ereg[938]), .B(n19486), .Z(n23238) );
  NANDN U30321 ( .A(n19481), .B(ereg[939]), .Z(n23237) );
  NAND U30322 ( .A(n23239), .B(n23240), .Z(n14437) );
  NANDN U30323 ( .A(init), .B(e[940]), .Z(n23240) );
  AND U30324 ( .A(n23241), .B(n23242), .Z(n23239) );
  NAND U30325 ( .A(ereg[939]), .B(n19486), .Z(n23242) );
  NANDN U30326 ( .A(n19481), .B(ereg[940]), .Z(n23241) );
  NAND U30327 ( .A(n23243), .B(n23244), .Z(n14436) );
  NANDN U30328 ( .A(init), .B(e[941]), .Z(n23244) );
  AND U30329 ( .A(n23245), .B(n23246), .Z(n23243) );
  NAND U30330 ( .A(ereg[940]), .B(n19486), .Z(n23246) );
  NANDN U30331 ( .A(n19481), .B(ereg[941]), .Z(n23245) );
  NAND U30332 ( .A(n23247), .B(n23248), .Z(n14435) );
  NANDN U30333 ( .A(init), .B(e[942]), .Z(n23248) );
  AND U30334 ( .A(n23249), .B(n23250), .Z(n23247) );
  NAND U30335 ( .A(ereg[941]), .B(n19486), .Z(n23250) );
  NANDN U30336 ( .A(n19481), .B(ereg[942]), .Z(n23249) );
  NAND U30337 ( .A(n23251), .B(n23252), .Z(n14434) );
  NANDN U30338 ( .A(init), .B(e[943]), .Z(n23252) );
  AND U30339 ( .A(n23253), .B(n23254), .Z(n23251) );
  NAND U30340 ( .A(ereg[942]), .B(n19486), .Z(n23254) );
  NANDN U30341 ( .A(n19481), .B(ereg[943]), .Z(n23253) );
  NAND U30342 ( .A(n23255), .B(n23256), .Z(n14433) );
  NANDN U30343 ( .A(init), .B(e[944]), .Z(n23256) );
  AND U30344 ( .A(n23257), .B(n23258), .Z(n23255) );
  NAND U30345 ( .A(ereg[943]), .B(n19486), .Z(n23258) );
  NANDN U30346 ( .A(n19481), .B(ereg[944]), .Z(n23257) );
  NAND U30347 ( .A(n23259), .B(n23260), .Z(n14432) );
  NANDN U30348 ( .A(init), .B(e[945]), .Z(n23260) );
  AND U30349 ( .A(n23261), .B(n23262), .Z(n23259) );
  NAND U30350 ( .A(ereg[944]), .B(n19486), .Z(n23262) );
  NANDN U30351 ( .A(n19481), .B(ereg[945]), .Z(n23261) );
  NAND U30352 ( .A(n23263), .B(n23264), .Z(n14431) );
  NANDN U30353 ( .A(init), .B(e[946]), .Z(n23264) );
  AND U30354 ( .A(n23265), .B(n23266), .Z(n23263) );
  NAND U30355 ( .A(ereg[945]), .B(n19486), .Z(n23266) );
  NANDN U30356 ( .A(n19481), .B(ereg[946]), .Z(n23265) );
  NAND U30357 ( .A(n23267), .B(n23268), .Z(n14430) );
  NANDN U30358 ( .A(init), .B(e[947]), .Z(n23268) );
  AND U30359 ( .A(n23269), .B(n23270), .Z(n23267) );
  NAND U30360 ( .A(ereg[946]), .B(n19486), .Z(n23270) );
  NANDN U30361 ( .A(n19481), .B(ereg[947]), .Z(n23269) );
  NAND U30362 ( .A(n23271), .B(n23272), .Z(n14429) );
  NANDN U30363 ( .A(init), .B(e[948]), .Z(n23272) );
  AND U30364 ( .A(n23273), .B(n23274), .Z(n23271) );
  NAND U30365 ( .A(ereg[947]), .B(n19486), .Z(n23274) );
  NANDN U30366 ( .A(n19481), .B(ereg[948]), .Z(n23273) );
  NAND U30367 ( .A(n23275), .B(n23276), .Z(n14428) );
  NANDN U30368 ( .A(init), .B(e[949]), .Z(n23276) );
  AND U30369 ( .A(n23277), .B(n23278), .Z(n23275) );
  NAND U30370 ( .A(ereg[948]), .B(n19486), .Z(n23278) );
  NANDN U30371 ( .A(n19481), .B(ereg[949]), .Z(n23277) );
  NAND U30372 ( .A(n23279), .B(n23280), .Z(n14427) );
  NANDN U30373 ( .A(init), .B(e[950]), .Z(n23280) );
  AND U30374 ( .A(n23281), .B(n23282), .Z(n23279) );
  NAND U30375 ( .A(ereg[949]), .B(n19486), .Z(n23282) );
  NANDN U30376 ( .A(n19481), .B(ereg[950]), .Z(n23281) );
  NAND U30377 ( .A(n23283), .B(n23284), .Z(n14426) );
  NANDN U30378 ( .A(init), .B(e[951]), .Z(n23284) );
  AND U30379 ( .A(n23285), .B(n23286), .Z(n23283) );
  NAND U30380 ( .A(ereg[950]), .B(n19486), .Z(n23286) );
  NANDN U30381 ( .A(n19481), .B(ereg[951]), .Z(n23285) );
  NAND U30382 ( .A(n23287), .B(n23288), .Z(n14425) );
  NANDN U30383 ( .A(init), .B(e[952]), .Z(n23288) );
  AND U30384 ( .A(n23289), .B(n23290), .Z(n23287) );
  NAND U30385 ( .A(ereg[951]), .B(n19486), .Z(n23290) );
  NANDN U30386 ( .A(n19481), .B(ereg[952]), .Z(n23289) );
  NAND U30387 ( .A(n23291), .B(n23292), .Z(n14424) );
  NANDN U30388 ( .A(init), .B(e[953]), .Z(n23292) );
  AND U30389 ( .A(n23293), .B(n23294), .Z(n23291) );
  NAND U30390 ( .A(ereg[952]), .B(n19486), .Z(n23294) );
  NANDN U30391 ( .A(n19481), .B(ereg[953]), .Z(n23293) );
  NAND U30392 ( .A(n23295), .B(n23296), .Z(n14423) );
  NANDN U30393 ( .A(init), .B(e[954]), .Z(n23296) );
  AND U30394 ( .A(n23297), .B(n23298), .Z(n23295) );
  NAND U30395 ( .A(ereg[953]), .B(n19486), .Z(n23298) );
  NANDN U30396 ( .A(n19481), .B(ereg[954]), .Z(n23297) );
  NAND U30397 ( .A(n23299), .B(n23300), .Z(n14422) );
  NANDN U30398 ( .A(init), .B(e[955]), .Z(n23300) );
  AND U30399 ( .A(n23301), .B(n23302), .Z(n23299) );
  NAND U30400 ( .A(ereg[954]), .B(n19486), .Z(n23302) );
  NANDN U30401 ( .A(n19481), .B(ereg[955]), .Z(n23301) );
  NAND U30402 ( .A(n23303), .B(n23304), .Z(n14421) );
  NANDN U30403 ( .A(init), .B(e[956]), .Z(n23304) );
  AND U30404 ( .A(n23305), .B(n23306), .Z(n23303) );
  NAND U30405 ( .A(ereg[955]), .B(n19486), .Z(n23306) );
  NANDN U30406 ( .A(n19481), .B(ereg[956]), .Z(n23305) );
  NAND U30407 ( .A(n23307), .B(n23308), .Z(n14420) );
  NANDN U30408 ( .A(init), .B(e[957]), .Z(n23308) );
  AND U30409 ( .A(n23309), .B(n23310), .Z(n23307) );
  NAND U30410 ( .A(ereg[956]), .B(n19486), .Z(n23310) );
  NANDN U30411 ( .A(n19481), .B(ereg[957]), .Z(n23309) );
  NAND U30412 ( .A(n23311), .B(n23312), .Z(n14419) );
  NANDN U30413 ( .A(init), .B(e[958]), .Z(n23312) );
  AND U30414 ( .A(n23313), .B(n23314), .Z(n23311) );
  NAND U30415 ( .A(ereg[957]), .B(n19486), .Z(n23314) );
  NANDN U30416 ( .A(n19481), .B(ereg[958]), .Z(n23313) );
  NAND U30417 ( .A(n23315), .B(n23316), .Z(n14418) );
  NANDN U30418 ( .A(init), .B(e[959]), .Z(n23316) );
  AND U30419 ( .A(n23317), .B(n23318), .Z(n23315) );
  NAND U30420 ( .A(ereg[958]), .B(n19486), .Z(n23318) );
  NANDN U30421 ( .A(n19481), .B(ereg[959]), .Z(n23317) );
  NAND U30422 ( .A(n23319), .B(n23320), .Z(n14417) );
  NANDN U30423 ( .A(init), .B(e[960]), .Z(n23320) );
  AND U30424 ( .A(n23321), .B(n23322), .Z(n23319) );
  NAND U30425 ( .A(ereg[959]), .B(n19486), .Z(n23322) );
  NANDN U30426 ( .A(n19481), .B(ereg[960]), .Z(n23321) );
  NAND U30427 ( .A(n23323), .B(n23324), .Z(n14416) );
  NANDN U30428 ( .A(init), .B(e[961]), .Z(n23324) );
  AND U30429 ( .A(n23325), .B(n23326), .Z(n23323) );
  NAND U30430 ( .A(ereg[960]), .B(n19486), .Z(n23326) );
  NANDN U30431 ( .A(n19481), .B(ereg[961]), .Z(n23325) );
  NAND U30432 ( .A(n23327), .B(n23328), .Z(n14415) );
  NANDN U30433 ( .A(init), .B(e[962]), .Z(n23328) );
  AND U30434 ( .A(n23329), .B(n23330), .Z(n23327) );
  NAND U30435 ( .A(ereg[961]), .B(n19486), .Z(n23330) );
  NANDN U30436 ( .A(n19481), .B(ereg[962]), .Z(n23329) );
  NAND U30437 ( .A(n23331), .B(n23332), .Z(n14414) );
  NANDN U30438 ( .A(init), .B(e[963]), .Z(n23332) );
  AND U30439 ( .A(n23333), .B(n23334), .Z(n23331) );
  NAND U30440 ( .A(ereg[962]), .B(n19486), .Z(n23334) );
  NANDN U30441 ( .A(n19481), .B(ereg[963]), .Z(n23333) );
  NAND U30442 ( .A(n23335), .B(n23336), .Z(n14413) );
  NANDN U30443 ( .A(init), .B(e[964]), .Z(n23336) );
  AND U30444 ( .A(n23337), .B(n23338), .Z(n23335) );
  NAND U30445 ( .A(ereg[963]), .B(n19486), .Z(n23338) );
  NANDN U30446 ( .A(n19481), .B(ereg[964]), .Z(n23337) );
  NAND U30447 ( .A(n23339), .B(n23340), .Z(n14412) );
  NANDN U30448 ( .A(init), .B(e[965]), .Z(n23340) );
  AND U30449 ( .A(n23341), .B(n23342), .Z(n23339) );
  NAND U30450 ( .A(ereg[964]), .B(n19486), .Z(n23342) );
  NANDN U30451 ( .A(n19481), .B(ereg[965]), .Z(n23341) );
  NAND U30452 ( .A(n23343), .B(n23344), .Z(n14411) );
  NANDN U30453 ( .A(init), .B(e[966]), .Z(n23344) );
  AND U30454 ( .A(n23345), .B(n23346), .Z(n23343) );
  NAND U30455 ( .A(ereg[965]), .B(n19486), .Z(n23346) );
  NANDN U30456 ( .A(n19481), .B(ereg[966]), .Z(n23345) );
  NAND U30457 ( .A(n23347), .B(n23348), .Z(n14410) );
  NANDN U30458 ( .A(init), .B(e[967]), .Z(n23348) );
  AND U30459 ( .A(n23349), .B(n23350), .Z(n23347) );
  NAND U30460 ( .A(ereg[966]), .B(n19486), .Z(n23350) );
  NANDN U30461 ( .A(n19481), .B(ereg[967]), .Z(n23349) );
  NAND U30462 ( .A(n23351), .B(n23352), .Z(n14409) );
  NANDN U30463 ( .A(init), .B(e[968]), .Z(n23352) );
  AND U30464 ( .A(n23353), .B(n23354), .Z(n23351) );
  NAND U30465 ( .A(ereg[967]), .B(n19486), .Z(n23354) );
  NANDN U30466 ( .A(n19481), .B(ereg[968]), .Z(n23353) );
  NAND U30467 ( .A(n23355), .B(n23356), .Z(n14408) );
  NANDN U30468 ( .A(init), .B(e[969]), .Z(n23356) );
  AND U30469 ( .A(n23357), .B(n23358), .Z(n23355) );
  NAND U30470 ( .A(ereg[968]), .B(n19486), .Z(n23358) );
  NANDN U30471 ( .A(n19481), .B(ereg[969]), .Z(n23357) );
  NAND U30472 ( .A(n23359), .B(n23360), .Z(n14407) );
  NANDN U30473 ( .A(init), .B(e[970]), .Z(n23360) );
  AND U30474 ( .A(n23361), .B(n23362), .Z(n23359) );
  NAND U30475 ( .A(ereg[969]), .B(n19486), .Z(n23362) );
  NANDN U30476 ( .A(n19481), .B(ereg[970]), .Z(n23361) );
  NAND U30477 ( .A(n23363), .B(n23364), .Z(n14406) );
  NANDN U30478 ( .A(init), .B(e[971]), .Z(n23364) );
  AND U30479 ( .A(n23365), .B(n23366), .Z(n23363) );
  NAND U30480 ( .A(ereg[970]), .B(n19486), .Z(n23366) );
  NANDN U30481 ( .A(n19481), .B(ereg[971]), .Z(n23365) );
  NAND U30482 ( .A(n23367), .B(n23368), .Z(n14405) );
  NANDN U30483 ( .A(init), .B(e[972]), .Z(n23368) );
  AND U30484 ( .A(n23369), .B(n23370), .Z(n23367) );
  NAND U30485 ( .A(ereg[971]), .B(n19486), .Z(n23370) );
  NANDN U30486 ( .A(n19481), .B(ereg[972]), .Z(n23369) );
  NAND U30487 ( .A(n23371), .B(n23372), .Z(n14404) );
  NANDN U30488 ( .A(init), .B(e[973]), .Z(n23372) );
  AND U30489 ( .A(n23373), .B(n23374), .Z(n23371) );
  NAND U30490 ( .A(ereg[972]), .B(n19486), .Z(n23374) );
  NANDN U30491 ( .A(n19481), .B(ereg[973]), .Z(n23373) );
  NAND U30492 ( .A(n23375), .B(n23376), .Z(n14403) );
  NANDN U30493 ( .A(init), .B(e[974]), .Z(n23376) );
  AND U30494 ( .A(n23377), .B(n23378), .Z(n23375) );
  NAND U30495 ( .A(ereg[973]), .B(n19486), .Z(n23378) );
  NANDN U30496 ( .A(n19481), .B(ereg[974]), .Z(n23377) );
  NAND U30497 ( .A(n23379), .B(n23380), .Z(n14402) );
  NANDN U30498 ( .A(init), .B(e[975]), .Z(n23380) );
  AND U30499 ( .A(n23381), .B(n23382), .Z(n23379) );
  NAND U30500 ( .A(ereg[974]), .B(n19486), .Z(n23382) );
  NANDN U30501 ( .A(n19481), .B(ereg[975]), .Z(n23381) );
  NAND U30502 ( .A(n23383), .B(n23384), .Z(n14401) );
  NANDN U30503 ( .A(init), .B(e[976]), .Z(n23384) );
  AND U30504 ( .A(n23385), .B(n23386), .Z(n23383) );
  NAND U30505 ( .A(ereg[975]), .B(n19486), .Z(n23386) );
  NANDN U30506 ( .A(n19481), .B(ereg[976]), .Z(n23385) );
  NAND U30507 ( .A(n23387), .B(n23388), .Z(n14400) );
  NANDN U30508 ( .A(init), .B(e[977]), .Z(n23388) );
  AND U30509 ( .A(n23389), .B(n23390), .Z(n23387) );
  NAND U30510 ( .A(ereg[976]), .B(n19486), .Z(n23390) );
  NANDN U30511 ( .A(n19481), .B(ereg[977]), .Z(n23389) );
  NAND U30512 ( .A(n23391), .B(n23392), .Z(n14399) );
  NANDN U30513 ( .A(init), .B(e[978]), .Z(n23392) );
  AND U30514 ( .A(n23393), .B(n23394), .Z(n23391) );
  NAND U30515 ( .A(ereg[977]), .B(n19486), .Z(n23394) );
  NANDN U30516 ( .A(n19481), .B(ereg[978]), .Z(n23393) );
  NAND U30517 ( .A(n23395), .B(n23396), .Z(n14398) );
  NANDN U30518 ( .A(init), .B(e[979]), .Z(n23396) );
  AND U30519 ( .A(n23397), .B(n23398), .Z(n23395) );
  NAND U30520 ( .A(ereg[978]), .B(n19486), .Z(n23398) );
  NANDN U30521 ( .A(n19481), .B(ereg[979]), .Z(n23397) );
  NAND U30522 ( .A(n23399), .B(n23400), .Z(n14397) );
  NANDN U30523 ( .A(init), .B(e[980]), .Z(n23400) );
  AND U30524 ( .A(n23401), .B(n23402), .Z(n23399) );
  NAND U30525 ( .A(ereg[979]), .B(n19486), .Z(n23402) );
  NANDN U30526 ( .A(n19481), .B(ereg[980]), .Z(n23401) );
  NAND U30527 ( .A(n23403), .B(n23404), .Z(n14396) );
  NANDN U30528 ( .A(init), .B(e[981]), .Z(n23404) );
  AND U30529 ( .A(n23405), .B(n23406), .Z(n23403) );
  NAND U30530 ( .A(ereg[980]), .B(n19486), .Z(n23406) );
  NANDN U30531 ( .A(n19481), .B(ereg[981]), .Z(n23405) );
  NAND U30532 ( .A(n23407), .B(n23408), .Z(n14395) );
  NANDN U30533 ( .A(init), .B(e[982]), .Z(n23408) );
  AND U30534 ( .A(n23409), .B(n23410), .Z(n23407) );
  NAND U30535 ( .A(ereg[981]), .B(n19486), .Z(n23410) );
  NANDN U30536 ( .A(n19481), .B(ereg[982]), .Z(n23409) );
  NAND U30537 ( .A(n23411), .B(n23412), .Z(n14394) );
  NANDN U30538 ( .A(init), .B(e[983]), .Z(n23412) );
  AND U30539 ( .A(n23413), .B(n23414), .Z(n23411) );
  NAND U30540 ( .A(ereg[982]), .B(n19486), .Z(n23414) );
  NANDN U30541 ( .A(n19481), .B(ereg[983]), .Z(n23413) );
  NAND U30542 ( .A(n23415), .B(n23416), .Z(n14393) );
  NANDN U30543 ( .A(init), .B(e[984]), .Z(n23416) );
  AND U30544 ( .A(n23417), .B(n23418), .Z(n23415) );
  NAND U30545 ( .A(ereg[983]), .B(n19486), .Z(n23418) );
  NANDN U30546 ( .A(n19481), .B(ereg[984]), .Z(n23417) );
  NAND U30547 ( .A(n23419), .B(n23420), .Z(n14392) );
  NANDN U30548 ( .A(init), .B(e[985]), .Z(n23420) );
  AND U30549 ( .A(n23421), .B(n23422), .Z(n23419) );
  NAND U30550 ( .A(ereg[984]), .B(n19486), .Z(n23422) );
  NANDN U30551 ( .A(n19481), .B(ereg[985]), .Z(n23421) );
  NAND U30552 ( .A(n23423), .B(n23424), .Z(n14391) );
  NANDN U30553 ( .A(init), .B(e[986]), .Z(n23424) );
  AND U30554 ( .A(n23425), .B(n23426), .Z(n23423) );
  NAND U30555 ( .A(ereg[985]), .B(n19486), .Z(n23426) );
  NANDN U30556 ( .A(n19481), .B(ereg[986]), .Z(n23425) );
  NAND U30557 ( .A(n23427), .B(n23428), .Z(n14390) );
  NANDN U30558 ( .A(init), .B(e[987]), .Z(n23428) );
  AND U30559 ( .A(n23429), .B(n23430), .Z(n23427) );
  NAND U30560 ( .A(ereg[986]), .B(n19486), .Z(n23430) );
  NANDN U30561 ( .A(n19481), .B(ereg[987]), .Z(n23429) );
  NAND U30562 ( .A(n23431), .B(n23432), .Z(n14389) );
  NANDN U30563 ( .A(init), .B(e[988]), .Z(n23432) );
  AND U30564 ( .A(n23433), .B(n23434), .Z(n23431) );
  NAND U30565 ( .A(ereg[987]), .B(n19486), .Z(n23434) );
  NANDN U30566 ( .A(n19481), .B(ereg[988]), .Z(n23433) );
  NAND U30567 ( .A(n23435), .B(n23436), .Z(n14388) );
  NANDN U30568 ( .A(init), .B(e[989]), .Z(n23436) );
  AND U30569 ( .A(n23437), .B(n23438), .Z(n23435) );
  NAND U30570 ( .A(ereg[988]), .B(n19486), .Z(n23438) );
  NANDN U30571 ( .A(n19481), .B(ereg[989]), .Z(n23437) );
  NAND U30572 ( .A(n23439), .B(n23440), .Z(n14387) );
  NANDN U30573 ( .A(init), .B(e[990]), .Z(n23440) );
  AND U30574 ( .A(n23441), .B(n23442), .Z(n23439) );
  NAND U30575 ( .A(ereg[989]), .B(n19486), .Z(n23442) );
  NANDN U30576 ( .A(n19481), .B(ereg[990]), .Z(n23441) );
  NAND U30577 ( .A(n23443), .B(n23444), .Z(n14386) );
  NANDN U30578 ( .A(init), .B(e[991]), .Z(n23444) );
  AND U30579 ( .A(n23445), .B(n23446), .Z(n23443) );
  NAND U30580 ( .A(ereg[990]), .B(n19486), .Z(n23446) );
  NANDN U30581 ( .A(n19481), .B(ereg[991]), .Z(n23445) );
  NAND U30582 ( .A(n23447), .B(n23448), .Z(n14385) );
  NANDN U30583 ( .A(init), .B(e[992]), .Z(n23448) );
  AND U30584 ( .A(n23449), .B(n23450), .Z(n23447) );
  NAND U30585 ( .A(ereg[991]), .B(n19486), .Z(n23450) );
  NANDN U30586 ( .A(n19481), .B(ereg[992]), .Z(n23449) );
  NAND U30587 ( .A(n23451), .B(n23452), .Z(n14384) );
  NANDN U30588 ( .A(init), .B(e[993]), .Z(n23452) );
  AND U30589 ( .A(n23453), .B(n23454), .Z(n23451) );
  NAND U30590 ( .A(ereg[992]), .B(n19486), .Z(n23454) );
  NANDN U30591 ( .A(n19481), .B(ereg[993]), .Z(n23453) );
  NAND U30592 ( .A(n23455), .B(n23456), .Z(n14383) );
  NANDN U30593 ( .A(init), .B(e[994]), .Z(n23456) );
  AND U30594 ( .A(n23457), .B(n23458), .Z(n23455) );
  NAND U30595 ( .A(ereg[993]), .B(n19486), .Z(n23458) );
  NANDN U30596 ( .A(n19481), .B(ereg[994]), .Z(n23457) );
  NAND U30597 ( .A(n23459), .B(n23460), .Z(n14382) );
  NANDN U30598 ( .A(init), .B(e[995]), .Z(n23460) );
  AND U30599 ( .A(n23461), .B(n23462), .Z(n23459) );
  NAND U30600 ( .A(ereg[994]), .B(n19486), .Z(n23462) );
  NANDN U30601 ( .A(n19481), .B(ereg[995]), .Z(n23461) );
  NAND U30602 ( .A(n23463), .B(n23464), .Z(n14381) );
  NANDN U30603 ( .A(init), .B(e[996]), .Z(n23464) );
  AND U30604 ( .A(n23465), .B(n23466), .Z(n23463) );
  NAND U30605 ( .A(ereg[995]), .B(n19486), .Z(n23466) );
  NANDN U30606 ( .A(n19481), .B(ereg[996]), .Z(n23465) );
  NAND U30607 ( .A(n23467), .B(n23468), .Z(n14380) );
  NANDN U30608 ( .A(init), .B(e[997]), .Z(n23468) );
  AND U30609 ( .A(n23469), .B(n23470), .Z(n23467) );
  NAND U30610 ( .A(ereg[996]), .B(n19486), .Z(n23470) );
  NANDN U30611 ( .A(n19481), .B(ereg[997]), .Z(n23469) );
  NAND U30612 ( .A(n23471), .B(n23472), .Z(n14379) );
  NANDN U30613 ( .A(init), .B(e[998]), .Z(n23472) );
  AND U30614 ( .A(n23473), .B(n23474), .Z(n23471) );
  NAND U30615 ( .A(ereg[997]), .B(n19486), .Z(n23474) );
  NANDN U30616 ( .A(n19481), .B(ereg[998]), .Z(n23473) );
  NAND U30617 ( .A(n23475), .B(n23476), .Z(n14378) );
  NANDN U30618 ( .A(init), .B(e[999]), .Z(n23476) );
  AND U30619 ( .A(n23477), .B(n23478), .Z(n23475) );
  NAND U30620 ( .A(ereg[998]), .B(n19486), .Z(n23478) );
  NANDN U30621 ( .A(n19481), .B(ereg[999]), .Z(n23477) );
  NAND U30622 ( .A(n23479), .B(n23480), .Z(n14377) );
  NANDN U30623 ( .A(init), .B(e[1000]), .Z(n23480) );
  AND U30624 ( .A(n23481), .B(n23482), .Z(n23479) );
  NAND U30625 ( .A(ereg[999]), .B(n19486), .Z(n23482) );
  NANDN U30626 ( .A(n19481), .B(ereg[1000]), .Z(n23481) );
  NAND U30627 ( .A(n23483), .B(n23484), .Z(n14376) );
  NANDN U30628 ( .A(init), .B(e[1001]), .Z(n23484) );
  AND U30629 ( .A(n23485), .B(n23486), .Z(n23483) );
  NAND U30630 ( .A(ereg[1000]), .B(n19486), .Z(n23486) );
  NANDN U30631 ( .A(n19481), .B(ereg[1001]), .Z(n23485) );
  NAND U30632 ( .A(n23487), .B(n23488), .Z(n14375) );
  NANDN U30633 ( .A(init), .B(e[1002]), .Z(n23488) );
  AND U30634 ( .A(n23489), .B(n23490), .Z(n23487) );
  NAND U30635 ( .A(ereg[1001]), .B(n19486), .Z(n23490) );
  NANDN U30636 ( .A(n19481), .B(ereg[1002]), .Z(n23489) );
  NAND U30637 ( .A(n23491), .B(n23492), .Z(n14374) );
  NANDN U30638 ( .A(init), .B(e[1003]), .Z(n23492) );
  AND U30639 ( .A(n23493), .B(n23494), .Z(n23491) );
  NAND U30640 ( .A(ereg[1002]), .B(n19486), .Z(n23494) );
  NANDN U30641 ( .A(n19481), .B(ereg[1003]), .Z(n23493) );
  NAND U30642 ( .A(n23495), .B(n23496), .Z(n14373) );
  NANDN U30643 ( .A(init), .B(e[1004]), .Z(n23496) );
  AND U30644 ( .A(n23497), .B(n23498), .Z(n23495) );
  NAND U30645 ( .A(ereg[1003]), .B(n19486), .Z(n23498) );
  NANDN U30646 ( .A(n19481), .B(ereg[1004]), .Z(n23497) );
  NAND U30647 ( .A(n23499), .B(n23500), .Z(n14372) );
  NANDN U30648 ( .A(init), .B(e[1005]), .Z(n23500) );
  AND U30649 ( .A(n23501), .B(n23502), .Z(n23499) );
  NAND U30650 ( .A(ereg[1004]), .B(n19486), .Z(n23502) );
  NANDN U30651 ( .A(n19481), .B(ereg[1005]), .Z(n23501) );
  NAND U30652 ( .A(n23503), .B(n23504), .Z(n14371) );
  NANDN U30653 ( .A(init), .B(e[1006]), .Z(n23504) );
  AND U30654 ( .A(n23505), .B(n23506), .Z(n23503) );
  NAND U30655 ( .A(ereg[1005]), .B(n19486), .Z(n23506) );
  NANDN U30656 ( .A(n19481), .B(ereg[1006]), .Z(n23505) );
  NAND U30657 ( .A(n23507), .B(n23508), .Z(n14370) );
  NANDN U30658 ( .A(init), .B(e[1007]), .Z(n23508) );
  AND U30659 ( .A(n23509), .B(n23510), .Z(n23507) );
  NAND U30660 ( .A(ereg[1006]), .B(n19486), .Z(n23510) );
  NANDN U30661 ( .A(n19481), .B(ereg[1007]), .Z(n23509) );
  NAND U30662 ( .A(n23511), .B(n23512), .Z(n14369) );
  NANDN U30663 ( .A(init), .B(e[1008]), .Z(n23512) );
  AND U30664 ( .A(n23513), .B(n23514), .Z(n23511) );
  NAND U30665 ( .A(ereg[1007]), .B(n19486), .Z(n23514) );
  NANDN U30666 ( .A(n19481), .B(ereg[1008]), .Z(n23513) );
  NAND U30667 ( .A(n23515), .B(n23516), .Z(n14368) );
  NANDN U30668 ( .A(init), .B(e[1009]), .Z(n23516) );
  AND U30669 ( .A(n23517), .B(n23518), .Z(n23515) );
  NAND U30670 ( .A(ereg[1008]), .B(n19486), .Z(n23518) );
  NANDN U30671 ( .A(n19481), .B(ereg[1009]), .Z(n23517) );
  NAND U30672 ( .A(n23519), .B(n23520), .Z(n14367) );
  NANDN U30673 ( .A(init), .B(e[1010]), .Z(n23520) );
  AND U30674 ( .A(n23521), .B(n23522), .Z(n23519) );
  NAND U30675 ( .A(ereg[1009]), .B(n19486), .Z(n23522) );
  NANDN U30676 ( .A(n19481), .B(ereg[1010]), .Z(n23521) );
  NAND U30677 ( .A(n23523), .B(n23524), .Z(n14366) );
  NANDN U30678 ( .A(init), .B(e[1011]), .Z(n23524) );
  AND U30679 ( .A(n23525), .B(n23526), .Z(n23523) );
  NAND U30680 ( .A(ereg[1010]), .B(n19486), .Z(n23526) );
  NANDN U30681 ( .A(n19481), .B(ereg[1011]), .Z(n23525) );
  NAND U30682 ( .A(n23527), .B(n23528), .Z(n14365) );
  NANDN U30683 ( .A(init), .B(e[1012]), .Z(n23528) );
  AND U30684 ( .A(n23529), .B(n23530), .Z(n23527) );
  NAND U30685 ( .A(ereg[1011]), .B(n19486), .Z(n23530) );
  NANDN U30686 ( .A(n19481), .B(ereg[1012]), .Z(n23529) );
  NAND U30687 ( .A(n23531), .B(n23532), .Z(n14364) );
  NANDN U30688 ( .A(init), .B(e[1013]), .Z(n23532) );
  AND U30689 ( .A(n23533), .B(n23534), .Z(n23531) );
  NAND U30690 ( .A(ereg[1012]), .B(n19486), .Z(n23534) );
  NANDN U30691 ( .A(n19481), .B(ereg[1013]), .Z(n23533) );
  NAND U30692 ( .A(n23535), .B(n23536), .Z(n14363) );
  NANDN U30693 ( .A(init), .B(e[1014]), .Z(n23536) );
  AND U30694 ( .A(n23537), .B(n23538), .Z(n23535) );
  NAND U30695 ( .A(ereg[1013]), .B(n19486), .Z(n23538) );
  NANDN U30696 ( .A(n19481), .B(ereg[1014]), .Z(n23537) );
  NAND U30697 ( .A(n23539), .B(n23540), .Z(n14362) );
  NANDN U30698 ( .A(init), .B(e[1015]), .Z(n23540) );
  AND U30699 ( .A(n23541), .B(n23542), .Z(n23539) );
  NAND U30700 ( .A(ereg[1014]), .B(n19486), .Z(n23542) );
  NANDN U30701 ( .A(n19481), .B(ereg[1015]), .Z(n23541) );
  NAND U30702 ( .A(n23543), .B(n23544), .Z(n14361) );
  NANDN U30703 ( .A(init), .B(e[1016]), .Z(n23544) );
  AND U30704 ( .A(n23545), .B(n23546), .Z(n23543) );
  NAND U30705 ( .A(ereg[1015]), .B(n19486), .Z(n23546) );
  NANDN U30706 ( .A(n19481), .B(ereg[1016]), .Z(n23545) );
  NAND U30707 ( .A(n23547), .B(n23548), .Z(n14360) );
  NANDN U30708 ( .A(init), .B(e[1017]), .Z(n23548) );
  AND U30709 ( .A(n23549), .B(n23550), .Z(n23547) );
  NAND U30710 ( .A(ereg[1016]), .B(n19486), .Z(n23550) );
  NANDN U30711 ( .A(n19481), .B(ereg[1017]), .Z(n23549) );
  NAND U30712 ( .A(n23551), .B(n23552), .Z(n14359) );
  NANDN U30713 ( .A(init), .B(e[1018]), .Z(n23552) );
  AND U30714 ( .A(n23553), .B(n23554), .Z(n23551) );
  NAND U30715 ( .A(ereg[1017]), .B(n19486), .Z(n23554) );
  NANDN U30716 ( .A(n19481), .B(ereg[1018]), .Z(n23553) );
  NAND U30717 ( .A(n23555), .B(n23556), .Z(n14358) );
  NANDN U30718 ( .A(init), .B(e[1019]), .Z(n23556) );
  AND U30719 ( .A(n23557), .B(n23558), .Z(n23555) );
  NAND U30720 ( .A(ereg[1018]), .B(n19486), .Z(n23558) );
  NANDN U30721 ( .A(n19481), .B(ereg[1019]), .Z(n23557) );
  NAND U30722 ( .A(n23559), .B(n23560), .Z(n14357) );
  NANDN U30723 ( .A(init), .B(e[1020]), .Z(n23560) );
  AND U30724 ( .A(n23561), .B(n23562), .Z(n23559) );
  NAND U30725 ( .A(ereg[1019]), .B(n19486), .Z(n23562) );
  NANDN U30726 ( .A(n19481), .B(ereg[1020]), .Z(n23561) );
  NAND U30727 ( .A(n23563), .B(n23564), .Z(n14356) );
  NANDN U30728 ( .A(init), .B(e[1021]), .Z(n23564) );
  AND U30729 ( .A(n23565), .B(n23566), .Z(n23563) );
  NAND U30730 ( .A(ereg[1020]), .B(n19486), .Z(n23566) );
  NANDN U30731 ( .A(n19481), .B(ereg[1021]), .Z(n23565) );
  NAND U30732 ( .A(n23567), .B(n23568), .Z(n14355) );
  NANDN U30733 ( .A(init), .B(e[1022]), .Z(n23568) );
  AND U30734 ( .A(n23569), .B(n23570), .Z(n23567) );
  NAND U30735 ( .A(ereg[1021]), .B(n19486), .Z(n23570) );
  NANDN U30736 ( .A(n19481), .B(ereg[1022]), .Z(n23569) );
  NAND U30737 ( .A(n23571), .B(n23572), .Z(n14354) );
  NANDN U30738 ( .A(init), .B(e[1023]), .Z(n23572) );
  AND U30739 ( .A(n23573), .B(n23574), .Z(n23571) );
  NAND U30740 ( .A(ereg[1022]), .B(n19486), .Z(n23574) );
  AND U30741 ( .A(start_in[1023]), .B(n19481), .Z(n19486) );
  NANDN U30742 ( .A(n19481), .B(ereg[1023]), .Z(n23573) );
  AND U30743 ( .A(n23575), .B(n15381), .Z(n19481) );
  NANDN U30744 ( .A(mul_pow), .B(init), .Z(n15381) );
  NANDN U30745 ( .A(start_in[1023]), .B(init), .Z(n23575) );
  NAND U30746 ( .A(n23576), .B(n19424), .Z(n14353) );
  NANDN U30747 ( .A(init), .B(m[1023]), .Z(n19424) );
  AND U30748 ( .A(n23577), .B(n23578), .Z(n23576) );
  NAND U30749 ( .A(o[1023]), .B(n23579), .Z(n23578) );
  NANDN U30750 ( .A(n23580), .B(creg[1023]), .Z(n23577) );
  NAND U30751 ( .A(n23581), .B(n19476), .Z(n14352) );
  NANDN U30752 ( .A(init), .B(m[0]), .Z(n19476) );
  AND U30753 ( .A(n23582), .B(n23583), .Z(n23581) );
  NAND U30754 ( .A(o[0]), .B(n23579), .Z(n23583) );
  NANDN U30755 ( .A(n23580), .B(creg[0]), .Z(n23582) );
  NAND U30756 ( .A(n23584), .B(n19206), .Z(n14351) );
  NANDN U30757 ( .A(init), .B(m[1]), .Z(n19206) );
  AND U30758 ( .A(n23585), .B(n23586), .Z(n23584) );
  NAND U30759 ( .A(o[1]), .B(n23579), .Z(n23586) );
  NANDN U30760 ( .A(n23580), .B(creg[1]), .Z(n23585) );
  NAND U30761 ( .A(n23587), .B(n18984), .Z(n14350) );
  NANDN U30762 ( .A(init), .B(m[2]), .Z(n18984) );
  AND U30763 ( .A(n23588), .B(n23589), .Z(n23587) );
  NAND U30764 ( .A(o[2]), .B(n23579), .Z(n23589) );
  NANDN U30765 ( .A(n23580), .B(creg[2]), .Z(n23588) );
  NAND U30766 ( .A(n23590), .B(n18762), .Z(n14349) );
  NANDN U30767 ( .A(init), .B(m[3]), .Z(n18762) );
  AND U30768 ( .A(n23591), .B(n23592), .Z(n23590) );
  NAND U30769 ( .A(o[3]), .B(n23579), .Z(n23592) );
  NANDN U30770 ( .A(n23580), .B(creg[3]), .Z(n23591) );
  NAND U30771 ( .A(n23593), .B(n18540), .Z(n14348) );
  NANDN U30772 ( .A(init), .B(m[4]), .Z(n18540) );
  AND U30773 ( .A(n23594), .B(n23595), .Z(n23593) );
  NAND U30774 ( .A(o[4]), .B(n23579), .Z(n23595) );
  NANDN U30775 ( .A(n23580), .B(creg[4]), .Z(n23594) );
  NAND U30776 ( .A(n23596), .B(n18318), .Z(n14347) );
  NANDN U30777 ( .A(init), .B(m[5]), .Z(n18318) );
  AND U30778 ( .A(n23597), .B(n23598), .Z(n23596) );
  NAND U30779 ( .A(o[5]), .B(n23579), .Z(n23598) );
  NANDN U30780 ( .A(n23580), .B(creg[5]), .Z(n23597) );
  NAND U30781 ( .A(n23599), .B(n18096), .Z(n14346) );
  NANDN U30782 ( .A(init), .B(m[6]), .Z(n18096) );
  AND U30783 ( .A(n23600), .B(n23601), .Z(n23599) );
  NAND U30784 ( .A(o[6]), .B(n23579), .Z(n23601) );
  NANDN U30785 ( .A(n23580), .B(creg[6]), .Z(n23600) );
  NAND U30786 ( .A(n23602), .B(n17874), .Z(n14345) );
  NANDN U30787 ( .A(init), .B(m[7]), .Z(n17874) );
  AND U30788 ( .A(n23603), .B(n23604), .Z(n23602) );
  NAND U30789 ( .A(o[7]), .B(n23579), .Z(n23604) );
  NANDN U30790 ( .A(n23580), .B(creg[7]), .Z(n23603) );
  NAND U30791 ( .A(n23605), .B(n17652), .Z(n14344) );
  NANDN U30792 ( .A(init), .B(m[8]), .Z(n17652) );
  AND U30793 ( .A(n23606), .B(n23607), .Z(n23605) );
  NAND U30794 ( .A(o[8]), .B(n23579), .Z(n23607) );
  NANDN U30795 ( .A(n23580), .B(creg[8]), .Z(n23606) );
  NAND U30796 ( .A(n23608), .B(n17430), .Z(n14343) );
  NANDN U30797 ( .A(init), .B(m[9]), .Z(n17430) );
  AND U30798 ( .A(n23609), .B(n23610), .Z(n23608) );
  NAND U30799 ( .A(o[9]), .B(n23579), .Z(n23610) );
  NANDN U30800 ( .A(n23580), .B(creg[9]), .Z(n23609) );
  NAND U30801 ( .A(n23611), .B(n19406), .Z(n14342) );
  NANDN U30802 ( .A(init), .B(m[10]), .Z(n19406) );
  AND U30803 ( .A(n23612), .B(n23613), .Z(n23611) );
  NAND U30804 ( .A(o[10]), .B(n23579), .Z(n23613) );
  NANDN U30805 ( .A(n23580), .B(creg[10]), .Z(n23612) );
  NAND U30806 ( .A(n23614), .B(n19384), .Z(n14341) );
  NANDN U30807 ( .A(init), .B(m[11]), .Z(n19384) );
  AND U30808 ( .A(n23615), .B(n23616), .Z(n23614) );
  NAND U30809 ( .A(o[11]), .B(n23579), .Z(n23616) );
  NANDN U30810 ( .A(n23580), .B(creg[11]), .Z(n23615) );
  NAND U30811 ( .A(n23617), .B(n19362), .Z(n14340) );
  NANDN U30812 ( .A(init), .B(m[12]), .Z(n19362) );
  AND U30813 ( .A(n23618), .B(n23619), .Z(n23617) );
  NAND U30814 ( .A(o[12]), .B(n23579), .Z(n23619) );
  NANDN U30815 ( .A(n23580), .B(creg[12]), .Z(n23618) );
  NAND U30816 ( .A(n23620), .B(n19340), .Z(n14339) );
  NANDN U30817 ( .A(init), .B(m[13]), .Z(n19340) );
  AND U30818 ( .A(n23621), .B(n23622), .Z(n23620) );
  NAND U30819 ( .A(o[13]), .B(n23579), .Z(n23622) );
  NANDN U30820 ( .A(n23580), .B(creg[13]), .Z(n23621) );
  NAND U30821 ( .A(n23623), .B(n19318), .Z(n14338) );
  NANDN U30822 ( .A(init), .B(m[14]), .Z(n19318) );
  AND U30823 ( .A(n23624), .B(n23625), .Z(n23623) );
  NAND U30824 ( .A(o[14]), .B(n23579), .Z(n23625) );
  NANDN U30825 ( .A(n23580), .B(creg[14]), .Z(n23624) );
  NAND U30826 ( .A(n23626), .B(n19296), .Z(n14337) );
  NANDN U30827 ( .A(init), .B(m[15]), .Z(n19296) );
  AND U30828 ( .A(n23627), .B(n23628), .Z(n23626) );
  NAND U30829 ( .A(o[15]), .B(n23579), .Z(n23628) );
  NANDN U30830 ( .A(n23580), .B(creg[15]), .Z(n23627) );
  NAND U30831 ( .A(n23629), .B(n19274), .Z(n14336) );
  NANDN U30832 ( .A(init), .B(m[16]), .Z(n19274) );
  AND U30833 ( .A(n23630), .B(n23631), .Z(n23629) );
  NAND U30834 ( .A(o[16]), .B(n23579), .Z(n23631) );
  NANDN U30835 ( .A(n23580), .B(creg[16]), .Z(n23630) );
  NAND U30836 ( .A(n23632), .B(n19252), .Z(n14335) );
  NANDN U30837 ( .A(init), .B(m[17]), .Z(n19252) );
  AND U30838 ( .A(n23633), .B(n23634), .Z(n23632) );
  NAND U30839 ( .A(o[17]), .B(n23579), .Z(n23634) );
  NANDN U30840 ( .A(n23580), .B(creg[17]), .Z(n23633) );
  NAND U30841 ( .A(n23635), .B(n19230), .Z(n14334) );
  NANDN U30842 ( .A(init), .B(m[18]), .Z(n19230) );
  AND U30843 ( .A(n23636), .B(n23637), .Z(n23635) );
  NAND U30844 ( .A(o[18]), .B(n23579), .Z(n23637) );
  NANDN U30845 ( .A(n23580), .B(creg[18]), .Z(n23636) );
  NAND U30846 ( .A(n23638), .B(n19208), .Z(n14333) );
  NANDN U30847 ( .A(init), .B(m[19]), .Z(n19208) );
  AND U30848 ( .A(n23639), .B(n23640), .Z(n23638) );
  NAND U30849 ( .A(o[19]), .B(n23579), .Z(n23640) );
  NANDN U30850 ( .A(n23580), .B(creg[19]), .Z(n23639) );
  NAND U30851 ( .A(n23641), .B(n19184), .Z(n14332) );
  NANDN U30852 ( .A(init), .B(m[20]), .Z(n19184) );
  AND U30853 ( .A(n23642), .B(n23643), .Z(n23641) );
  NAND U30854 ( .A(o[20]), .B(n23579), .Z(n23643) );
  NANDN U30855 ( .A(n23580), .B(creg[20]), .Z(n23642) );
  NAND U30856 ( .A(n23644), .B(n19162), .Z(n14331) );
  NANDN U30857 ( .A(init), .B(m[21]), .Z(n19162) );
  AND U30858 ( .A(n23645), .B(n23646), .Z(n23644) );
  NAND U30859 ( .A(o[21]), .B(n23579), .Z(n23646) );
  NANDN U30860 ( .A(n23580), .B(creg[21]), .Z(n23645) );
  NAND U30861 ( .A(n23647), .B(n19140), .Z(n14330) );
  NANDN U30862 ( .A(init), .B(m[22]), .Z(n19140) );
  AND U30863 ( .A(n23648), .B(n23649), .Z(n23647) );
  NAND U30864 ( .A(o[22]), .B(n23579), .Z(n23649) );
  NANDN U30865 ( .A(n23580), .B(creg[22]), .Z(n23648) );
  NAND U30866 ( .A(n23650), .B(n19118), .Z(n14329) );
  NANDN U30867 ( .A(init), .B(m[23]), .Z(n19118) );
  AND U30868 ( .A(n23651), .B(n23652), .Z(n23650) );
  NAND U30869 ( .A(o[23]), .B(n23579), .Z(n23652) );
  NANDN U30870 ( .A(n23580), .B(creg[23]), .Z(n23651) );
  NAND U30871 ( .A(n23653), .B(n19096), .Z(n14328) );
  NANDN U30872 ( .A(init), .B(m[24]), .Z(n19096) );
  AND U30873 ( .A(n23654), .B(n23655), .Z(n23653) );
  NAND U30874 ( .A(o[24]), .B(n23579), .Z(n23655) );
  NANDN U30875 ( .A(n23580), .B(creg[24]), .Z(n23654) );
  NAND U30876 ( .A(n23656), .B(n19074), .Z(n14327) );
  NANDN U30877 ( .A(init), .B(m[25]), .Z(n19074) );
  AND U30878 ( .A(n23657), .B(n23658), .Z(n23656) );
  NAND U30879 ( .A(o[25]), .B(n23579), .Z(n23658) );
  NANDN U30880 ( .A(n23580), .B(creg[25]), .Z(n23657) );
  NAND U30881 ( .A(n23659), .B(n19052), .Z(n14326) );
  NANDN U30882 ( .A(init), .B(m[26]), .Z(n19052) );
  AND U30883 ( .A(n23660), .B(n23661), .Z(n23659) );
  NAND U30884 ( .A(o[26]), .B(n23579), .Z(n23661) );
  NANDN U30885 ( .A(n23580), .B(creg[26]), .Z(n23660) );
  NAND U30886 ( .A(n23662), .B(n19030), .Z(n14325) );
  NANDN U30887 ( .A(init), .B(m[27]), .Z(n19030) );
  AND U30888 ( .A(n23663), .B(n23664), .Z(n23662) );
  NAND U30889 ( .A(o[27]), .B(n23579), .Z(n23664) );
  NANDN U30890 ( .A(n23580), .B(creg[27]), .Z(n23663) );
  NAND U30891 ( .A(n23665), .B(n19008), .Z(n14324) );
  NANDN U30892 ( .A(init), .B(m[28]), .Z(n19008) );
  AND U30893 ( .A(n23666), .B(n23667), .Z(n23665) );
  NAND U30894 ( .A(o[28]), .B(n23579), .Z(n23667) );
  NANDN U30895 ( .A(n23580), .B(creg[28]), .Z(n23666) );
  NAND U30896 ( .A(n23668), .B(n18986), .Z(n14323) );
  NANDN U30897 ( .A(init), .B(m[29]), .Z(n18986) );
  AND U30898 ( .A(n23669), .B(n23670), .Z(n23668) );
  NAND U30899 ( .A(o[29]), .B(n23579), .Z(n23670) );
  NANDN U30900 ( .A(n23580), .B(creg[29]), .Z(n23669) );
  NAND U30901 ( .A(n23671), .B(n18962), .Z(n14322) );
  NANDN U30902 ( .A(init), .B(m[30]), .Z(n18962) );
  AND U30903 ( .A(n23672), .B(n23673), .Z(n23671) );
  NAND U30904 ( .A(o[30]), .B(n23579), .Z(n23673) );
  NANDN U30905 ( .A(n23580), .B(creg[30]), .Z(n23672) );
  NAND U30906 ( .A(n23674), .B(n18940), .Z(n14321) );
  NANDN U30907 ( .A(init), .B(m[31]), .Z(n18940) );
  AND U30908 ( .A(n23675), .B(n23676), .Z(n23674) );
  NAND U30909 ( .A(o[31]), .B(n23579), .Z(n23676) );
  NANDN U30910 ( .A(n23580), .B(creg[31]), .Z(n23675) );
  NAND U30911 ( .A(n23677), .B(n18918), .Z(n14320) );
  NANDN U30912 ( .A(init), .B(m[32]), .Z(n18918) );
  AND U30913 ( .A(n23678), .B(n23679), .Z(n23677) );
  NAND U30914 ( .A(o[32]), .B(n23579), .Z(n23679) );
  NANDN U30915 ( .A(n23580), .B(creg[32]), .Z(n23678) );
  NAND U30916 ( .A(n23680), .B(n18896), .Z(n14319) );
  NANDN U30917 ( .A(init), .B(m[33]), .Z(n18896) );
  AND U30918 ( .A(n23681), .B(n23682), .Z(n23680) );
  NAND U30919 ( .A(o[33]), .B(n23579), .Z(n23682) );
  NANDN U30920 ( .A(n23580), .B(creg[33]), .Z(n23681) );
  NAND U30921 ( .A(n23683), .B(n18874), .Z(n14318) );
  NANDN U30922 ( .A(init), .B(m[34]), .Z(n18874) );
  AND U30923 ( .A(n23684), .B(n23685), .Z(n23683) );
  NAND U30924 ( .A(o[34]), .B(n23579), .Z(n23685) );
  NANDN U30925 ( .A(n23580), .B(creg[34]), .Z(n23684) );
  NAND U30926 ( .A(n23686), .B(n18852), .Z(n14317) );
  NANDN U30927 ( .A(init), .B(m[35]), .Z(n18852) );
  AND U30928 ( .A(n23687), .B(n23688), .Z(n23686) );
  NAND U30929 ( .A(o[35]), .B(n23579), .Z(n23688) );
  NANDN U30930 ( .A(n23580), .B(creg[35]), .Z(n23687) );
  NAND U30931 ( .A(n23689), .B(n18830), .Z(n14316) );
  NANDN U30932 ( .A(init), .B(m[36]), .Z(n18830) );
  AND U30933 ( .A(n23690), .B(n23691), .Z(n23689) );
  NAND U30934 ( .A(o[36]), .B(n23579), .Z(n23691) );
  NANDN U30935 ( .A(n23580), .B(creg[36]), .Z(n23690) );
  NAND U30936 ( .A(n23692), .B(n18808), .Z(n14315) );
  NANDN U30937 ( .A(init), .B(m[37]), .Z(n18808) );
  AND U30938 ( .A(n23693), .B(n23694), .Z(n23692) );
  NAND U30939 ( .A(o[37]), .B(n23579), .Z(n23694) );
  NANDN U30940 ( .A(n23580), .B(creg[37]), .Z(n23693) );
  NAND U30941 ( .A(n23695), .B(n18786), .Z(n14314) );
  NANDN U30942 ( .A(init), .B(m[38]), .Z(n18786) );
  AND U30943 ( .A(n23696), .B(n23697), .Z(n23695) );
  NAND U30944 ( .A(o[38]), .B(n23579), .Z(n23697) );
  NANDN U30945 ( .A(n23580), .B(creg[38]), .Z(n23696) );
  NAND U30946 ( .A(n23698), .B(n18764), .Z(n14313) );
  NANDN U30947 ( .A(init), .B(m[39]), .Z(n18764) );
  AND U30948 ( .A(n23699), .B(n23700), .Z(n23698) );
  NAND U30949 ( .A(o[39]), .B(n23579), .Z(n23700) );
  NANDN U30950 ( .A(n23580), .B(creg[39]), .Z(n23699) );
  NAND U30951 ( .A(n23701), .B(n18740), .Z(n14312) );
  NANDN U30952 ( .A(init), .B(m[40]), .Z(n18740) );
  AND U30953 ( .A(n23702), .B(n23703), .Z(n23701) );
  NAND U30954 ( .A(o[40]), .B(n23579), .Z(n23703) );
  NANDN U30955 ( .A(n23580), .B(creg[40]), .Z(n23702) );
  NAND U30956 ( .A(n23704), .B(n18718), .Z(n14311) );
  NANDN U30957 ( .A(init), .B(m[41]), .Z(n18718) );
  AND U30958 ( .A(n23705), .B(n23706), .Z(n23704) );
  NAND U30959 ( .A(o[41]), .B(n23579), .Z(n23706) );
  NANDN U30960 ( .A(n23580), .B(creg[41]), .Z(n23705) );
  NAND U30961 ( .A(n23707), .B(n18696), .Z(n14310) );
  NANDN U30962 ( .A(init), .B(m[42]), .Z(n18696) );
  AND U30963 ( .A(n23708), .B(n23709), .Z(n23707) );
  NAND U30964 ( .A(o[42]), .B(n23579), .Z(n23709) );
  NANDN U30965 ( .A(n23580), .B(creg[42]), .Z(n23708) );
  NAND U30966 ( .A(n23710), .B(n18674), .Z(n14309) );
  NANDN U30967 ( .A(init), .B(m[43]), .Z(n18674) );
  AND U30968 ( .A(n23711), .B(n23712), .Z(n23710) );
  NAND U30969 ( .A(o[43]), .B(n23579), .Z(n23712) );
  NANDN U30970 ( .A(n23580), .B(creg[43]), .Z(n23711) );
  NAND U30971 ( .A(n23713), .B(n18652), .Z(n14308) );
  NANDN U30972 ( .A(init), .B(m[44]), .Z(n18652) );
  AND U30973 ( .A(n23714), .B(n23715), .Z(n23713) );
  NAND U30974 ( .A(o[44]), .B(n23579), .Z(n23715) );
  NANDN U30975 ( .A(n23580), .B(creg[44]), .Z(n23714) );
  NAND U30976 ( .A(n23716), .B(n18630), .Z(n14307) );
  NANDN U30977 ( .A(init), .B(m[45]), .Z(n18630) );
  AND U30978 ( .A(n23717), .B(n23718), .Z(n23716) );
  NAND U30979 ( .A(o[45]), .B(n23579), .Z(n23718) );
  NANDN U30980 ( .A(n23580), .B(creg[45]), .Z(n23717) );
  NAND U30981 ( .A(n23719), .B(n18608), .Z(n14306) );
  NANDN U30982 ( .A(init), .B(m[46]), .Z(n18608) );
  AND U30983 ( .A(n23720), .B(n23721), .Z(n23719) );
  NAND U30984 ( .A(o[46]), .B(n23579), .Z(n23721) );
  NANDN U30985 ( .A(n23580), .B(creg[46]), .Z(n23720) );
  NAND U30986 ( .A(n23722), .B(n18586), .Z(n14305) );
  NANDN U30987 ( .A(init), .B(m[47]), .Z(n18586) );
  AND U30988 ( .A(n23723), .B(n23724), .Z(n23722) );
  NAND U30989 ( .A(o[47]), .B(n23579), .Z(n23724) );
  NANDN U30990 ( .A(n23580), .B(creg[47]), .Z(n23723) );
  NAND U30991 ( .A(n23725), .B(n18564), .Z(n14304) );
  NANDN U30992 ( .A(init), .B(m[48]), .Z(n18564) );
  AND U30993 ( .A(n23726), .B(n23727), .Z(n23725) );
  NAND U30994 ( .A(o[48]), .B(n23579), .Z(n23727) );
  NANDN U30995 ( .A(n23580), .B(creg[48]), .Z(n23726) );
  NAND U30996 ( .A(n23728), .B(n18542), .Z(n14303) );
  NANDN U30997 ( .A(init), .B(m[49]), .Z(n18542) );
  AND U30998 ( .A(n23729), .B(n23730), .Z(n23728) );
  NAND U30999 ( .A(o[49]), .B(n23579), .Z(n23730) );
  NANDN U31000 ( .A(n23580), .B(creg[49]), .Z(n23729) );
  NAND U31001 ( .A(n23731), .B(n18518), .Z(n14302) );
  NANDN U31002 ( .A(init), .B(m[50]), .Z(n18518) );
  AND U31003 ( .A(n23732), .B(n23733), .Z(n23731) );
  NAND U31004 ( .A(o[50]), .B(n23579), .Z(n23733) );
  NANDN U31005 ( .A(n23580), .B(creg[50]), .Z(n23732) );
  NAND U31006 ( .A(n23734), .B(n18496), .Z(n14301) );
  NANDN U31007 ( .A(init), .B(m[51]), .Z(n18496) );
  AND U31008 ( .A(n23735), .B(n23736), .Z(n23734) );
  NAND U31009 ( .A(o[51]), .B(n23579), .Z(n23736) );
  NANDN U31010 ( .A(n23580), .B(creg[51]), .Z(n23735) );
  NAND U31011 ( .A(n23737), .B(n18474), .Z(n14300) );
  NANDN U31012 ( .A(init), .B(m[52]), .Z(n18474) );
  AND U31013 ( .A(n23738), .B(n23739), .Z(n23737) );
  NAND U31014 ( .A(o[52]), .B(n23579), .Z(n23739) );
  NANDN U31015 ( .A(n23580), .B(creg[52]), .Z(n23738) );
  NAND U31016 ( .A(n23740), .B(n18452), .Z(n14299) );
  NANDN U31017 ( .A(init), .B(m[53]), .Z(n18452) );
  AND U31018 ( .A(n23741), .B(n23742), .Z(n23740) );
  NAND U31019 ( .A(o[53]), .B(n23579), .Z(n23742) );
  NANDN U31020 ( .A(n23580), .B(creg[53]), .Z(n23741) );
  NAND U31021 ( .A(n23743), .B(n18430), .Z(n14298) );
  NANDN U31022 ( .A(init), .B(m[54]), .Z(n18430) );
  AND U31023 ( .A(n23744), .B(n23745), .Z(n23743) );
  NAND U31024 ( .A(o[54]), .B(n23579), .Z(n23745) );
  NANDN U31025 ( .A(n23580), .B(creg[54]), .Z(n23744) );
  NAND U31026 ( .A(n23746), .B(n18408), .Z(n14297) );
  NANDN U31027 ( .A(init), .B(m[55]), .Z(n18408) );
  AND U31028 ( .A(n23747), .B(n23748), .Z(n23746) );
  NAND U31029 ( .A(o[55]), .B(n23579), .Z(n23748) );
  NANDN U31030 ( .A(n23580), .B(creg[55]), .Z(n23747) );
  NAND U31031 ( .A(n23749), .B(n18386), .Z(n14296) );
  NANDN U31032 ( .A(init), .B(m[56]), .Z(n18386) );
  AND U31033 ( .A(n23750), .B(n23751), .Z(n23749) );
  NAND U31034 ( .A(o[56]), .B(n23579), .Z(n23751) );
  NANDN U31035 ( .A(n23580), .B(creg[56]), .Z(n23750) );
  NAND U31036 ( .A(n23752), .B(n18364), .Z(n14295) );
  NANDN U31037 ( .A(init), .B(m[57]), .Z(n18364) );
  AND U31038 ( .A(n23753), .B(n23754), .Z(n23752) );
  NAND U31039 ( .A(o[57]), .B(n23579), .Z(n23754) );
  NANDN U31040 ( .A(n23580), .B(creg[57]), .Z(n23753) );
  NAND U31041 ( .A(n23755), .B(n18342), .Z(n14294) );
  NANDN U31042 ( .A(init), .B(m[58]), .Z(n18342) );
  AND U31043 ( .A(n23756), .B(n23757), .Z(n23755) );
  NAND U31044 ( .A(o[58]), .B(n23579), .Z(n23757) );
  NANDN U31045 ( .A(n23580), .B(creg[58]), .Z(n23756) );
  NAND U31046 ( .A(n23758), .B(n18320), .Z(n14293) );
  NANDN U31047 ( .A(init), .B(m[59]), .Z(n18320) );
  AND U31048 ( .A(n23759), .B(n23760), .Z(n23758) );
  NAND U31049 ( .A(o[59]), .B(n23579), .Z(n23760) );
  NANDN U31050 ( .A(n23580), .B(creg[59]), .Z(n23759) );
  NAND U31051 ( .A(n23761), .B(n18296), .Z(n14292) );
  NANDN U31052 ( .A(init), .B(m[60]), .Z(n18296) );
  AND U31053 ( .A(n23762), .B(n23763), .Z(n23761) );
  NAND U31054 ( .A(o[60]), .B(n23579), .Z(n23763) );
  NANDN U31055 ( .A(n23580), .B(creg[60]), .Z(n23762) );
  NAND U31056 ( .A(n23764), .B(n18274), .Z(n14291) );
  NANDN U31057 ( .A(init), .B(m[61]), .Z(n18274) );
  AND U31058 ( .A(n23765), .B(n23766), .Z(n23764) );
  NAND U31059 ( .A(o[61]), .B(n23579), .Z(n23766) );
  NANDN U31060 ( .A(n23580), .B(creg[61]), .Z(n23765) );
  NAND U31061 ( .A(n23767), .B(n18252), .Z(n14290) );
  NANDN U31062 ( .A(init), .B(m[62]), .Z(n18252) );
  AND U31063 ( .A(n23768), .B(n23769), .Z(n23767) );
  NAND U31064 ( .A(o[62]), .B(n23579), .Z(n23769) );
  NANDN U31065 ( .A(n23580), .B(creg[62]), .Z(n23768) );
  NAND U31066 ( .A(n23770), .B(n18230), .Z(n14289) );
  NANDN U31067 ( .A(init), .B(m[63]), .Z(n18230) );
  AND U31068 ( .A(n23771), .B(n23772), .Z(n23770) );
  NAND U31069 ( .A(o[63]), .B(n23579), .Z(n23772) );
  NANDN U31070 ( .A(n23580), .B(creg[63]), .Z(n23771) );
  NAND U31071 ( .A(n23773), .B(n18208), .Z(n14288) );
  NANDN U31072 ( .A(init), .B(m[64]), .Z(n18208) );
  AND U31073 ( .A(n23774), .B(n23775), .Z(n23773) );
  NAND U31074 ( .A(o[64]), .B(n23579), .Z(n23775) );
  NANDN U31075 ( .A(n23580), .B(creg[64]), .Z(n23774) );
  NAND U31076 ( .A(n23776), .B(n18186), .Z(n14287) );
  NANDN U31077 ( .A(init), .B(m[65]), .Z(n18186) );
  AND U31078 ( .A(n23777), .B(n23778), .Z(n23776) );
  NAND U31079 ( .A(o[65]), .B(n23579), .Z(n23778) );
  NANDN U31080 ( .A(n23580), .B(creg[65]), .Z(n23777) );
  NAND U31081 ( .A(n23779), .B(n18164), .Z(n14286) );
  NANDN U31082 ( .A(init), .B(m[66]), .Z(n18164) );
  AND U31083 ( .A(n23780), .B(n23781), .Z(n23779) );
  NAND U31084 ( .A(o[66]), .B(n23579), .Z(n23781) );
  NANDN U31085 ( .A(n23580), .B(creg[66]), .Z(n23780) );
  NAND U31086 ( .A(n23782), .B(n18142), .Z(n14285) );
  NANDN U31087 ( .A(init), .B(m[67]), .Z(n18142) );
  AND U31088 ( .A(n23783), .B(n23784), .Z(n23782) );
  NAND U31089 ( .A(o[67]), .B(n23579), .Z(n23784) );
  NANDN U31090 ( .A(n23580), .B(creg[67]), .Z(n23783) );
  NAND U31091 ( .A(n23785), .B(n18120), .Z(n14284) );
  NANDN U31092 ( .A(init), .B(m[68]), .Z(n18120) );
  AND U31093 ( .A(n23786), .B(n23787), .Z(n23785) );
  NAND U31094 ( .A(o[68]), .B(n23579), .Z(n23787) );
  NANDN U31095 ( .A(n23580), .B(creg[68]), .Z(n23786) );
  NAND U31096 ( .A(n23788), .B(n18098), .Z(n14283) );
  NANDN U31097 ( .A(init), .B(m[69]), .Z(n18098) );
  AND U31098 ( .A(n23789), .B(n23790), .Z(n23788) );
  NAND U31099 ( .A(o[69]), .B(n23579), .Z(n23790) );
  NANDN U31100 ( .A(n23580), .B(creg[69]), .Z(n23789) );
  NAND U31101 ( .A(n23791), .B(n18074), .Z(n14282) );
  NANDN U31102 ( .A(init), .B(m[70]), .Z(n18074) );
  AND U31103 ( .A(n23792), .B(n23793), .Z(n23791) );
  NAND U31104 ( .A(o[70]), .B(n23579), .Z(n23793) );
  NANDN U31105 ( .A(n23580), .B(creg[70]), .Z(n23792) );
  NAND U31106 ( .A(n23794), .B(n18052), .Z(n14281) );
  NANDN U31107 ( .A(init), .B(m[71]), .Z(n18052) );
  AND U31108 ( .A(n23795), .B(n23796), .Z(n23794) );
  NAND U31109 ( .A(o[71]), .B(n23579), .Z(n23796) );
  NANDN U31110 ( .A(n23580), .B(creg[71]), .Z(n23795) );
  NAND U31111 ( .A(n23797), .B(n18030), .Z(n14280) );
  NANDN U31112 ( .A(init), .B(m[72]), .Z(n18030) );
  AND U31113 ( .A(n23798), .B(n23799), .Z(n23797) );
  NAND U31114 ( .A(o[72]), .B(n23579), .Z(n23799) );
  NANDN U31115 ( .A(n23580), .B(creg[72]), .Z(n23798) );
  NAND U31116 ( .A(n23800), .B(n18008), .Z(n14279) );
  NANDN U31117 ( .A(init), .B(m[73]), .Z(n18008) );
  AND U31118 ( .A(n23801), .B(n23802), .Z(n23800) );
  NAND U31119 ( .A(o[73]), .B(n23579), .Z(n23802) );
  NANDN U31120 ( .A(n23580), .B(creg[73]), .Z(n23801) );
  NAND U31121 ( .A(n23803), .B(n17986), .Z(n14278) );
  NANDN U31122 ( .A(init), .B(m[74]), .Z(n17986) );
  AND U31123 ( .A(n23804), .B(n23805), .Z(n23803) );
  NAND U31124 ( .A(o[74]), .B(n23579), .Z(n23805) );
  NANDN U31125 ( .A(n23580), .B(creg[74]), .Z(n23804) );
  NAND U31126 ( .A(n23806), .B(n17964), .Z(n14277) );
  NANDN U31127 ( .A(init), .B(m[75]), .Z(n17964) );
  AND U31128 ( .A(n23807), .B(n23808), .Z(n23806) );
  NAND U31129 ( .A(o[75]), .B(n23579), .Z(n23808) );
  NANDN U31130 ( .A(n23580), .B(creg[75]), .Z(n23807) );
  NAND U31131 ( .A(n23809), .B(n17942), .Z(n14276) );
  NANDN U31132 ( .A(init), .B(m[76]), .Z(n17942) );
  AND U31133 ( .A(n23810), .B(n23811), .Z(n23809) );
  NAND U31134 ( .A(o[76]), .B(n23579), .Z(n23811) );
  NANDN U31135 ( .A(n23580), .B(creg[76]), .Z(n23810) );
  NAND U31136 ( .A(n23812), .B(n17920), .Z(n14275) );
  NANDN U31137 ( .A(init), .B(m[77]), .Z(n17920) );
  AND U31138 ( .A(n23813), .B(n23814), .Z(n23812) );
  NAND U31139 ( .A(o[77]), .B(n23579), .Z(n23814) );
  NANDN U31140 ( .A(n23580), .B(creg[77]), .Z(n23813) );
  NAND U31141 ( .A(n23815), .B(n17898), .Z(n14274) );
  NANDN U31142 ( .A(init), .B(m[78]), .Z(n17898) );
  AND U31143 ( .A(n23816), .B(n23817), .Z(n23815) );
  NAND U31144 ( .A(o[78]), .B(n23579), .Z(n23817) );
  NANDN U31145 ( .A(n23580), .B(creg[78]), .Z(n23816) );
  NAND U31146 ( .A(n23818), .B(n17876), .Z(n14273) );
  NANDN U31147 ( .A(init), .B(m[79]), .Z(n17876) );
  AND U31148 ( .A(n23819), .B(n23820), .Z(n23818) );
  NAND U31149 ( .A(o[79]), .B(n23579), .Z(n23820) );
  NANDN U31150 ( .A(n23580), .B(creg[79]), .Z(n23819) );
  NAND U31151 ( .A(n23821), .B(n17852), .Z(n14272) );
  NANDN U31152 ( .A(init), .B(m[80]), .Z(n17852) );
  AND U31153 ( .A(n23822), .B(n23823), .Z(n23821) );
  NAND U31154 ( .A(o[80]), .B(n23579), .Z(n23823) );
  NANDN U31155 ( .A(n23580), .B(creg[80]), .Z(n23822) );
  NAND U31156 ( .A(n23824), .B(n17830), .Z(n14271) );
  NANDN U31157 ( .A(init), .B(m[81]), .Z(n17830) );
  AND U31158 ( .A(n23825), .B(n23826), .Z(n23824) );
  NAND U31159 ( .A(o[81]), .B(n23579), .Z(n23826) );
  NANDN U31160 ( .A(n23580), .B(creg[81]), .Z(n23825) );
  NAND U31161 ( .A(n23827), .B(n17808), .Z(n14270) );
  NANDN U31162 ( .A(init), .B(m[82]), .Z(n17808) );
  AND U31163 ( .A(n23828), .B(n23829), .Z(n23827) );
  NAND U31164 ( .A(o[82]), .B(n23579), .Z(n23829) );
  NANDN U31165 ( .A(n23580), .B(creg[82]), .Z(n23828) );
  NAND U31166 ( .A(n23830), .B(n17786), .Z(n14269) );
  NANDN U31167 ( .A(init), .B(m[83]), .Z(n17786) );
  AND U31168 ( .A(n23831), .B(n23832), .Z(n23830) );
  NAND U31169 ( .A(o[83]), .B(n23579), .Z(n23832) );
  NANDN U31170 ( .A(n23580), .B(creg[83]), .Z(n23831) );
  NAND U31171 ( .A(n23833), .B(n17764), .Z(n14268) );
  NANDN U31172 ( .A(init), .B(m[84]), .Z(n17764) );
  AND U31173 ( .A(n23834), .B(n23835), .Z(n23833) );
  NAND U31174 ( .A(o[84]), .B(n23579), .Z(n23835) );
  NANDN U31175 ( .A(n23580), .B(creg[84]), .Z(n23834) );
  NAND U31176 ( .A(n23836), .B(n17742), .Z(n14267) );
  NANDN U31177 ( .A(init), .B(m[85]), .Z(n17742) );
  AND U31178 ( .A(n23837), .B(n23838), .Z(n23836) );
  NAND U31179 ( .A(o[85]), .B(n23579), .Z(n23838) );
  NANDN U31180 ( .A(n23580), .B(creg[85]), .Z(n23837) );
  NAND U31181 ( .A(n23839), .B(n17720), .Z(n14266) );
  NANDN U31182 ( .A(init), .B(m[86]), .Z(n17720) );
  AND U31183 ( .A(n23840), .B(n23841), .Z(n23839) );
  NAND U31184 ( .A(o[86]), .B(n23579), .Z(n23841) );
  NANDN U31185 ( .A(n23580), .B(creg[86]), .Z(n23840) );
  NAND U31186 ( .A(n23842), .B(n17698), .Z(n14265) );
  NANDN U31187 ( .A(init), .B(m[87]), .Z(n17698) );
  AND U31188 ( .A(n23843), .B(n23844), .Z(n23842) );
  NAND U31189 ( .A(o[87]), .B(n23579), .Z(n23844) );
  NANDN U31190 ( .A(n23580), .B(creg[87]), .Z(n23843) );
  NAND U31191 ( .A(n23845), .B(n17676), .Z(n14264) );
  NANDN U31192 ( .A(init), .B(m[88]), .Z(n17676) );
  AND U31193 ( .A(n23846), .B(n23847), .Z(n23845) );
  NAND U31194 ( .A(o[88]), .B(n23579), .Z(n23847) );
  NANDN U31195 ( .A(n23580), .B(creg[88]), .Z(n23846) );
  NAND U31196 ( .A(n23848), .B(n17654), .Z(n14263) );
  NANDN U31197 ( .A(init), .B(m[89]), .Z(n17654) );
  AND U31198 ( .A(n23849), .B(n23850), .Z(n23848) );
  NAND U31199 ( .A(o[89]), .B(n23579), .Z(n23850) );
  NANDN U31200 ( .A(n23580), .B(creg[89]), .Z(n23849) );
  NAND U31201 ( .A(n23851), .B(n17630), .Z(n14262) );
  NANDN U31202 ( .A(init), .B(m[90]), .Z(n17630) );
  AND U31203 ( .A(n23852), .B(n23853), .Z(n23851) );
  NAND U31204 ( .A(o[90]), .B(n23579), .Z(n23853) );
  NANDN U31205 ( .A(n23580), .B(creg[90]), .Z(n23852) );
  NAND U31206 ( .A(n23854), .B(n17608), .Z(n14261) );
  NANDN U31207 ( .A(init), .B(m[91]), .Z(n17608) );
  AND U31208 ( .A(n23855), .B(n23856), .Z(n23854) );
  NAND U31209 ( .A(o[91]), .B(n23579), .Z(n23856) );
  NANDN U31210 ( .A(n23580), .B(creg[91]), .Z(n23855) );
  NAND U31211 ( .A(n23857), .B(n17586), .Z(n14260) );
  NANDN U31212 ( .A(init), .B(m[92]), .Z(n17586) );
  AND U31213 ( .A(n23858), .B(n23859), .Z(n23857) );
  NAND U31214 ( .A(o[92]), .B(n23579), .Z(n23859) );
  NANDN U31215 ( .A(n23580), .B(creg[92]), .Z(n23858) );
  NAND U31216 ( .A(n23860), .B(n17564), .Z(n14259) );
  NANDN U31217 ( .A(init), .B(m[93]), .Z(n17564) );
  AND U31218 ( .A(n23861), .B(n23862), .Z(n23860) );
  NAND U31219 ( .A(o[93]), .B(n23579), .Z(n23862) );
  NANDN U31220 ( .A(n23580), .B(creg[93]), .Z(n23861) );
  NAND U31221 ( .A(n23863), .B(n17542), .Z(n14258) );
  NANDN U31222 ( .A(init), .B(m[94]), .Z(n17542) );
  AND U31223 ( .A(n23864), .B(n23865), .Z(n23863) );
  NAND U31224 ( .A(o[94]), .B(n23579), .Z(n23865) );
  NANDN U31225 ( .A(n23580), .B(creg[94]), .Z(n23864) );
  NAND U31226 ( .A(n23866), .B(n17520), .Z(n14257) );
  NANDN U31227 ( .A(init), .B(m[95]), .Z(n17520) );
  AND U31228 ( .A(n23867), .B(n23868), .Z(n23866) );
  NAND U31229 ( .A(o[95]), .B(n23579), .Z(n23868) );
  NANDN U31230 ( .A(n23580), .B(creg[95]), .Z(n23867) );
  NAND U31231 ( .A(n23869), .B(n17498), .Z(n14256) );
  NANDN U31232 ( .A(init), .B(m[96]), .Z(n17498) );
  AND U31233 ( .A(n23870), .B(n23871), .Z(n23869) );
  NAND U31234 ( .A(o[96]), .B(n23579), .Z(n23871) );
  NANDN U31235 ( .A(n23580), .B(creg[96]), .Z(n23870) );
  NAND U31236 ( .A(n23872), .B(n17476), .Z(n14255) );
  NANDN U31237 ( .A(init), .B(m[97]), .Z(n17476) );
  AND U31238 ( .A(n23873), .B(n23874), .Z(n23872) );
  NAND U31239 ( .A(o[97]), .B(n23579), .Z(n23874) );
  NANDN U31240 ( .A(n23580), .B(creg[97]), .Z(n23873) );
  NAND U31241 ( .A(n23875), .B(n17454), .Z(n14254) );
  NANDN U31242 ( .A(init), .B(m[98]), .Z(n17454) );
  AND U31243 ( .A(n23876), .B(n23877), .Z(n23875) );
  NAND U31244 ( .A(o[98]), .B(n23579), .Z(n23877) );
  NANDN U31245 ( .A(n23580), .B(creg[98]), .Z(n23876) );
  NAND U31246 ( .A(n23878), .B(n17432), .Z(n14253) );
  NANDN U31247 ( .A(init), .B(m[99]), .Z(n17432) );
  AND U31248 ( .A(n23879), .B(n23880), .Z(n23878) );
  NAND U31249 ( .A(o[99]), .B(n23579), .Z(n23880) );
  NANDN U31250 ( .A(n23580), .B(creg[99]), .Z(n23879) );
  NAND U31251 ( .A(n23881), .B(n19454), .Z(n14252) );
  NANDN U31252 ( .A(init), .B(m[100]), .Z(n19454) );
  AND U31253 ( .A(n23882), .B(n23883), .Z(n23881) );
  NAND U31254 ( .A(o[100]), .B(n23579), .Z(n23883) );
  NANDN U31255 ( .A(n23580), .B(creg[100]), .Z(n23882) );
  NAND U31256 ( .A(n23884), .B(n19432), .Z(n14251) );
  NANDN U31257 ( .A(init), .B(m[101]), .Z(n19432) );
  AND U31258 ( .A(n23885), .B(n23886), .Z(n23884) );
  NAND U31259 ( .A(o[101]), .B(n23579), .Z(n23886) );
  NANDN U31260 ( .A(n23580), .B(creg[101]), .Z(n23885) );
  NAND U31261 ( .A(n23887), .B(n19422), .Z(n14250) );
  NANDN U31262 ( .A(init), .B(m[102]), .Z(n19422) );
  AND U31263 ( .A(n23888), .B(n23889), .Z(n23887) );
  NAND U31264 ( .A(o[102]), .B(n23579), .Z(n23889) );
  NANDN U31265 ( .A(n23580), .B(creg[102]), .Z(n23888) );
  NAND U31266 ( .A(n23890), .B(n19420), .Z(n14249) );
  NANDN U31267 ( .A(init), .B(m[103]), .Z(n19420) );
  AND U31268 ( .A(n23891), .B(n23892), .Z(n23890) );
  NAND U31269 ( .A(o[103]), .B(n23579), .Z(n23892) );
  NANDN U31270 ( .A(n23580), .B(creg[103]), .Z(n23891) );
  NAND U31271 ( .A(n23893), .B(n19418), .Z(n14248) );
  NANDN U31272 ( .A(init), .B(m[104]), .Z(n19418) );
  AND U31273 ( .A(n23894), .B(n23895), .Z(n23893) );
  NAND U31274 ( .A(o[104]), .B(n23579), .Z(n23895) );
  NANDN U31275 ( .A(n23580), .B(creg[104]), .Z(n23894) );
  NAND U31276 ( .A(n23896), .B(n19416), .Z(n14247) );
  NANDN U31277 ( .A(init), .B(m[105]), .Z(n19416) );
  AND U31278 ( .A(n23897), .B(n23898), .Z(n23896) );
  NAND U31279 ( .A(o[105]), .B(n23579), .Z(n23898) );
  NANDN U31280 ( .A(n23580), .B(creg[105]), .Z(n23897) );
  NAND U31281 ( .A(n23899), .B(n19414), .Z(n14246) );
  NANDN U31282 ( .A(init), .B(m[106]), .Z(n19414) );
  AND U31283 ( .A(n23900), .B(n23901), .Z(n23899) );
  NAND U31284 ( .A(o[106]), .B(n23579), .Z(n23901) );
  NANDN U31285 ( .A(n23580), .B(creg[106]), .Z(n23900) );
  NAND U31286 ( .A(n23902), .B(n19412), .Z(n14245) );
  NANDN U31287 ( .A(init), .B(m[107]), .Z(n19412) );
  AND U31288 ( .A(n23903), .B(n23904), .Z(n23902) );
  NAND U31289 ( .A(o[107]), .B(n23579), .Z(n23904) );
  NANDN U31290 ( .A(n23580), .B(creg[107]), .Z(n23903) );
  NAND U31291 ( .A(n23905), .B(n19410), .Z(n14244) );
  NANDN U31292 ( .A(init), .B(m[108]), .Z(n19410) );
  AND U31293 ( .A(n23906), .B(n23907), .Z(n23905) );
  NAND U31294 ( .A(o[108]), .B(n23579), .Z(n23907) );
  NANDN U31295 ( .A(n23580), .B(creg[108]), .Z(n23906) );
  NAND U31296 ( .A(n23908), .B(n19408), .Z(n14243) );
  NANDN U31297 ( .A(init), .B(m[109]), .Z(n19408) );
  AND U31298 ( .A(n23909), .B(n23910), .Z(n23908) );
  NAND U31299 ( .A(o[109]), .B(n23579), .Z(n23910) );
  NANDN U31300 ( .A(n23580), .B(creg[109]), .Z(n23909) );
  NAND U31301 ( .A(n23911), .B(n19404), .Z(n14242) );
  NANDN U31302 ( .A(init), .B(m[110]), .Z(n19404) );
  AND U31303 ( .A(n23912), .B(n23913), .Z(n23911) );
  NAND U31304 ( .A(o[110]), .B(n23579), .Z(n23913) );
  NANDN U31305 ( .A(n23580), .B(creg[110]), .Z(n23912) );
  NAND U31306 ( .A(n23914), .B(n19402), .Z(n14241) );
  NANDN U31307 ( .A(init), .B(m[111]), .Z(n19402) );
  AND U31308 ( .A(n23915), .B(n23916), .Z(n23914) );
  NAND U31309 ( .A(o[111]), .B(n23579), .Z(n23916) );
  NANDN U31310 ( .A(n23580), .B(creg[111]), .Z(n23915) );
  NAND U31311 ( .A(n23917), .B(n19400), .Z(n14240) );
  NANDN U31312 ( .A(init), .B(m[112]), .Z(n19400) );
  AND U31313 ( .A(n23918), .B(n23919), .Z(n23917) );
  NAND U31314 ( .A(o[112]), .B(n23579), .Z(n23919) );
  NANDN U31315 ( .A(n23580), .B(creg[112]), .Z(n23918) );
  NAND U31316 ( .A(n23920), .B(n19398), .Z(n14239) );
  NANDN U31317 ( .A(init), .B(m[113]), .Z(n19398) );
  AND U31318 ( .A(n23921), .B(n23922), .Z(n23920) );
  NAND U31319 ( .A(o[113]), .B(n23579), .Z(n23922) );
  NANDN U31320 ( .A(n23580), .B(creg[113]), .Z(n23921) );
  NAND U31321 ( .A(n23923), .B(n19396), .Z(n14238) );
  NANDN U31322 ( .A(init), .B(m[114]), .Z(n19396) );
  AND U31323 ( .A(n23924), .B(n23925), .Z(n23923) );
  NAND U31324 ( .A(o[114]), .B(n23579), .Z(n23925) );
  NANDN U31325 ( .A(n23580), .B(creg[114]), .Z(n23924) );
  NAND U31326 ( .A(n23926), .B(n19394), .Z(n14237) );
  NANDN U31327 ( .A(init), .B(m[115]), .Z(n19394) );
  AND U31328 ( .A(n23927), .B(n23928), .Z(n23926) );
  NAND U31329 ( .A(o[115]), .B(n23579), .Z(n23928) );
  NANDN U31330 ( .A(n23580), .B(creg[115]), .Z(n23927) );
  NAND U31331 ( .A(n23929), .B(n19392), .Z(n14236) );
  NANDN U31332 ( .A(init), .B(m[116]), .Z(n19392) );
  AND U31333 ( .A(n23930), .B(n23931), .Z(n23929) );
  NAND U31334 ( .A(o[116]), .B(n23579), .Z(n23931) );
  NANDN U31335 ( .A(n23580), .B(creg[116]), .Z(n23930) );
  NAND U31336 ( .A(n23932), .B(n19390), .Z(n14235) );
  NANDN U31337 ( .A(init), .B(m[117]), .Z(n19390) );
  AND U31338 ( .A(n23933), .B(n23934), .Z(n23932) );
  NAND U31339 ( .A(o[117]), .B(n23579), .Z(n23934) );
  NANDN U31340 ( .A(n23580), .B(creg[117]), .Z(n23933) );
  NAND U31341 ( .A(n23935), .B(n19388), .Z(n14234) );
  NANDN U31342 ( .A(init), .B(m[118]), .Z(n19388) );
  AND U31343 ( .A(n23936), .B(n23937), .Z(n23935) );
  NAND U31344 ( .A(o[118]), .B(n23579), .Z(n23937) );
  NANDN U31345 ( .A(n23580), .B(creg[118]), .Z(n23936) );
  NAND U31346 ( .A(n23938), .B(n19386), .Z(n14233) );
  NANDN U31347 ( .A(init), .B(m[119]), .Z(n19386) );
  AND U31348 ( .A(n23939), .B(n23940), .Z(n23938) );
  NAND U31349 ( .A(o[119]), .B(n23579), .Z(n23940) );
  NANDN U31350 ( .A(n23580), .B(creg[119]), .Z(n23939) );
  NAND U31351 ( .A(n23941), .B(n19382), .Z(n14232) );
  NANDN U31352 ( .A(init), .B(m[120]), .Z(n19382) );
  AND U31353 ( .A(n23942), .B(n23943), .Z(n23941) );
  NAND U31354 ( .A(o[120]), .B(n23579), .Z(n23943) );
  NANDN U31355 ( .A(n23580), .B(creg[120]), .Z(n23942) );
  NAND U31356 ( .A(n23944), .B(n19380), .Z(n14231) );
  NANDN U31357 ( .A(init), .B(m[121]), .Z(n19380) );
  AND U31358 ( .A(n23945), .B(n23946), .Z(n23944) );
  NAND U31359 ( .A(o[121]), .B(n23579), .Z(n23946) );
  NANDN U31360 ( .A(n23580), .B(creg[121]), .Z(n23945) );
  NAND U31361 ( .A(n23947), .B(n19378), .Z(n14230) );
  NANDN U31362 ( .A(init), .B(m[122]), .Z(n19378) );
  AND U31363 ( .A(n23948), .B(n23949), .Z(n23947) );
  NAND U31364 ( .A(o[122]), .B(n23579), .Z(n23949) );
  NANDN U31365 ( .A(n23580), .B(creg[122]), .Z(n23948) );
  NAND U31366 ( .A(n23950), .B(n19376), .Z(n14229) );
  NANDN U31367 ( .A(init), .B(m[123]), .Z(n19376) );
  AND U31368 ( .A(n23951), .B(n23952), .Z(n23950) );
  NAND U31369 ( .A(o[123]), .B(n23579), .Z(n23952) );
  NANDN U31370 ( .A(n23580), .B(creg[123]), .Z(n23951) );
  NAND U31371 ( .A(n23953), .B(n19374), .Z(n14228) );
  NANDN U31372 ( .A(init), .B(m[124]), .Z(n19374) );
  AND U31373 ( .A(n23954), .B(n23955), .Z(n23953) );
  NAND U31374 ( .A(o[124]), .B(n23579), .Z(n23955) );
  NANDN U31375 ( .A(n23580), .B(creg[124]), .Z(n23954) );
  NAND U31376 ( .A(n23956), .B(n19372), .Z(n14227) );
  NANDN U31377 ( .A(init), .B(m[125]), .Z(n19372) );
  AND U31378 ( .A(n23957), .B(n23958), .Z(n23956) );
  NAND U31379 ( .A(o[125]), .B(n23579), .Z(n23958) );
  NANDN U31380 ( .A(n23580), .B(creg[125]), .Z(n23957) );
  NAND U31381 ( .A(n23959), .B(n19370), .Z(n14226) );
  NANDN U31382 ( .A(init), .B(m[126]), .Z(n19370) );
  AND U31383 ( .A(n23960), .B(n23961), .Z(n23959) );
  NAND U31384 ( .A(o[126]), .B(n23579), .Z(n23961) );
  NANDN U31385 ( .A(n23580), .B(creg[126]), .Z(n23960) );
  NAND U31386 ( .A(n23962), .B(n19368), .Z(n14225) );
  NANDN U31387 ( .A(init), .B(m[127]), .Z(n19368) );
  AND U31388 ( .A(n23963), .B(n23964), .Z(n23962) );
  NAND U31389 ( .A(o[127]), .B(n23579), .Z(n23964) );
  NANDN U31390 ( .A(n23580), .B(creg[127]), .Z(n23963) );
  NAND U31391 ( .A(n23965), .B(n19366), .Z(n14224) );
  NANDN U31392 ( .A(init), .B(m[128]), .Z(n19366) );
  AND U31393 ( .A(n23966), .B(n23967), .Z(n23965) );
  NAND U31394 ( .A(o[128]), .B(n23579), .Z(n23967) );
  NANDN U31395 ( .A(n23580), .B(creg[128]), .Z(n23966) );
  NAND U31396 ( .A(n23968), .B(n19364), .Z(n14223) );
  NANDN U31397 ( .A(init), .B(m[129]), .Z(n19364) );
  AND U31398 ( .A(n23969), .B(n23970), .Z(n23968) );
  NAND U31399 ( .A(o[129]), .B(n23579), .Z(n23970) );
  NANDN U31400 ( .A(n23580), .B(creg[129]), .Z(n23969) );
  NAND U31401 ( .A(n23971), .B(n19360), .Z(n14222) );
  NANDN U31402 ( .A(init), .B(m[130]), .Z(n19360) );
  AND U31403 ( .A(n23972), .B(n23973), .Z(n23971) );
  NAND U31404 ( .A(o[130]), .B(n23579), .Z(n23973) );
  NANDN U31405 ( .A(n23580), .B(creg[130]), .Z(n23972) );
  NAND U31406 ( .A(n23974), .B(n19358), .Z(n14221) );
  NANDN U31407 ( .A(init), .B(m[131]), .Z(n19358) );
  AND U31408 ( .A(n23975), .B(n23976), .Z(n23974) );
  NAND U31409 ( .A(o[131]), .B(n23579), .Z(n23976) );
  NANDN U31410 ( .A(n23580), .B(creg[131]), .Z(n23975) );
  NAND U31411 ( .A(n23977), .B(n19356), .Z(n14220) );
  NANDN U31412 ( .A(init), .B(m[132]), .Z(n19356) );
  AND U31413 ( .A(n23978), .B(n23979), .Z(n23977) );
  NAND U31414 ( .A(o[132]), .B(n23579), .Z(n23979) );
  NANDN U31415 ( .A(n23580), .B(creg[132]), .Z(n23978) );
  NAND U31416 ( .A(n23980), .B(n19354), .Z(n14219) );
  NANDN U31417 ( .A(init), .B(m[133]), .Z(n19354) );
  AND U31418 ( .A(n23981), .B(n23982), .Z(n23980) );
  NAND U31419 ( .A(o[133]), .B(n23579), .Z(n23982) );
  NANDN U31420 ( .A(n23580), .B(creg[133]), .Z(n23981) );
  NAND U31421 ( .A(n23983), .B(n19352), .Z(n14218) );
  NANDN U31422 ( .A(init), .B(m[134]), .Z(n19352) );
  AND U31423 ( .A(n23984), .B(n23985), .Z(n23983) );
  NAND U31424 ( .A(o[134]), .B(n23579), .Z(n23985) );
  NANDN U31425 ( .A(n23580), .B(creg[134]), .Z(n23984) );
  NAND U31426 ( .A(n23986), .B(n19350), .Z(n14217) );
  NANDN U31427 ( .A(init), .B(m[135]), .Z(n19350) );
  AND U31428 ( .A(n23987), .B(n23988), .Z(n23986) );
  NAND U31429 ( .A(o[135]), .B(n23579), .Z(n23988) );
  NANDN U31430 ( .A(n23580), .B(creg[135]), .Z(n23987) );
  NAND U31431 ( .A(n23989), .B(n19348), .Z(n14216) );
  NANDN U31432 ( .A(init), .B(m[136]), .Z(n19348) );
  AND U31433 ( .A(n23990), .B(n23991), .Z(n23989) );
  NAND U31434 ( .A(o[136]), .B(n23579), .Z(n23991) );
  NANDN U31435 ( .A(n23580), .B(creg[136]), .Z(n23990) );
  NAND U31436 ( .A(n23992), .B(n19346), .Z(n14215) );
  NANDN U31437 ( .A(init), .B(m[137]), .Z(n19346) );
  AND U31438 ( .A(n23993), .B(n23994), .Z(n23992) );
  NAND U31439 ( .A(o[137]), .B(n23579), .Z(n23994) );
  NANDN U31440 ( .A(n23580), .B(creg[137]), .Z(n23993) );
  NAND U31441 ( .A(n23995), .B(n19344), .Z(n14214) );
  NANDN U31442 ( .A(init), .B(m[138]), .Z(n19344) );
  AND U31443 ( .A(n23996), .B(n23997), .Z(n23995) );
  NAND U31444 ( .A(o[138]), .B(n23579), .Z(n23997) );
  NANDN U31445 ( .A(n23580), .B(creg[138]), .Z(n23996) );
  NAND U31446 ( .A(n23998), .B(n19342), .Z(n14213) );
  NANDN U31447 ( .A(init), .B(m[139]), .Z(n19342) );
  AND U31448 ( .A(n23999), .B(n24000), .Z(n23998) );
  NAND U31449 ( .A(o[139]), .B(n23579), .Z(n24000) );
  NANDN U31450 ( .A(n23580), .B(creg[139]), .Z(n23999) );
  NAND U31451 ( .A(n24001), .B(n19338), .Z(n14212) );
  NANDN U31452 ( .A(init), .B(m[140]), .Z(n19338) );
  AND U31453 ( .A(n24002), .B(n24003), .Z(n24001) );
  NAND U31454 ( .A(o[140]), .B(n23579), .Z(n24003) );
  NANDN U31455 ( .A(n23580), .B(creg[140]), .Z(n24002) );
  NAND U31456 ( .A(n24004), .B(n19336), .Z(n14211) );
  NANDN U31457 ( .A(init), .B(m[141]), .Z(n19336) );
  AND U31458 ( .A(n24005), .B(n24006), .Z(n24004) );
  NAND U31459 ( .A(o[141]), .B(n23579), .Z(n24006) );
  NANDN U31460 ( .A(n23580), .B(creg[141]), .Z(n24005) );
  NAND U31461 ( .A(n24007), .B(n19334), .Z(n14210) );
  NANDN U31462 ( .A(init), .B(m[142]), .Z(n19334) );
  AND U31463 ( .A(n24008), .B(n24009), .Z(n24007) );
  NAND U31464 ( .A(o[142]), .B(n23579), .Z(n24009) );
  NANDN U31465 ( .A(n23580), .B(creg[142]), .Z(n24008) );
  NAND U31466 ( .A(n24010), .B(n19332), .Z(n14209) );
  NANDN U31467 ( .A(init), .B(m[143]), .Z(n19332) );
  AND U31468 ( .A(n24011), .B(n24012), .Z(n24010) );
  NAND U31469 ( .A(o[143]), .B(n23579), .Z(n24012) );
  NANDN U31470 ( .A(n23580), .B(creg[143]), .Z(n24011) );
  NAND U31471 ( .A(n24013), .B(n19330), .Z(n14208) );
  NANDN U31472 ( .A(init), .B(m[144]), .Z(n19330) );
  AND U31473 ( .A(n24014), .B(n24015), .Z(n24013) );
  NAND U31474 ( .A(o[144]), .B(n23579), .Z(n24015) );
  NANDN U31475 ( .A(n23580), .B(creg[144]), .Z(n24014) );
  NAND U31476 ( .A(n24016), .B(n19328), .Z(n14207) );
  NANDN U31477 ( .A(init), .B(m[145]), .Z(n19328) );
  AND U31478 ( .A(n24017), .B(n24018), .Z(n24016) );
  NAND U31479 ( .A(o[145]), .B(n23579), .Z(n24018) );
  NANDN U31480 ( .A(n23580), .B(creg[145]), .Z(n24017) );
  NAND U31481 ( .A(n24019), .B(n19326), .Z(n14206) );
  NANDN U31482 ( .A(init), .B(m[146]), .Z(n19326) );
  AND U31483 ( .A(n24020), .B(n24021), .Z(n24019) );
  NAND U31484 ( .A(o[146]), .B(n23579), .Z(n24021) );
  NANDN U31485 ( .A(n23580), .B(creg[146]), .Z(n24020) );
  NAND U31486 ( .A(n24022), .B(n19324), .Z(n14205) );
  NANDN U31487 ( .A(init), .B(m[147]), .Z(n19324) );
  AND U31488 ( .A(n24023), .B(n24024), .Z(n24022) );
  NAND U31489 ( .A(o[147]), .B(n23579), .Z(n24024) );
  NANDN U31490 ( .A(n23580), .B(creg[147]), .Z(n24023) );
  NAND U31491 ( .A(n24025), .B(n19322), .Z(n14204) );
  NANDN U31492 ( .A(init), .B(m[148]), .Z(n19322) );
  AND U31493 ( .A(n24026), .B(n24027), .Z(n24025) );
  NAND U31494 ( .A(o[148]), .B(n23579), .Z(n24027) );
  NANDN U31495 ( .A(n23580), .B(creg[148]), .Z(n24026) );
  NAND U31496 ( .A(n24028), .B(n19320), .Z(n14203) );
  NANDN U31497 ( .A(init), .B(m[149]), .Z(n19320) );
  AND U31498 ( .A(n24029), .B(n24030), .Z(n24028) );
  NAND U31499 ( .A(o[149]), .B(n23579), .Z(n24030) );
  NANDN U31500 ( .A(n23580), .B(creg[149]), .Z(n24029) );
  NAND U31501 ( .A(n24031), .B(n19316), .Z(n14202) );
  NANDN U31502 ( .A(init), .B(m[150]), .Z(n19316) );
  AND U31503 ( .A(n24032), .B(n24033), .Z(n24031) );
  NAND U31504 ( .A(o[150]), .B(n23579), .Z(n24033) );
  NANDN U31505 ( .A(n23580), .B(creg[150]), .Z(n24032) );
  NAND U31506 ( .A(n24034), .B(n19314), .Z(n14201) );
  NANDN U31507 ( .A(init), .B(m[151]), .Z(n19314) );
  AND U31508 ( .A(n24035), .B(n24036), .Z(n24034) );
  NAND U31509 ( .A(o[151]), .B(n23579), .Z(n24036) );
  NANDN U31510 ( .A(n23580), .B(creg[151]), .Z(n24035) );
  NAND U31511 ( .A(n24037), .B(n19312), .Z(n14200) );
  NANDN U31512 ( .A(init), .B(m[152]), .Z(n19312) );
  AND U31513 ( .A(n24038), .B(n24039), .Z(n24037) );
  NAND U31514 ( .A(o[152]), .B(n23579), .Z(n24039) );
  NANDN U31515 ( .A(n23580), .B(creg[152]), .Z(n24038) );
  NAND U31516 ( .A(n24040), .B(n19310), .Z(n14199) );
  NANDN U31517 ( .A(init), .B(m[153]), .Z(n19310) );
  AND U31518 ( .A(n24041), .B(n24042), .Z(n24040) );
  NAND U31519 ( .A(o[153]), .B(n23579), .Z(n24042) );
  NANDN U31520 ( .A(n23580), .B(creg[153]), .Z(n24041) );
  NAND U31521 ( .A(n24043), .B(n19308), .Z(n14198) );
  NANDN U31522 ( .A(init), .B(m[154]), .Z(n19308) );
  AND U31523 ( .A(n24044), .B(n24045), .Z(n24043) );
  NAND U31524 ( .A(o[154]), .B(n23579), .Z(n24045) );
  NANDN U31525 ( .A(n23580), .B(creg[154]), .Z(n24044) );
  NAND U31526 ( .A(n24046), .B(n19306), .Z(n14197) );
  NANDN U31527 ( .A(init), .B(m[155]), .Z(n19306) );
  AND U31528 ( .A(n24047), .B(n24048), .Z(n24046) );
  NAND U31529 ( .A(o[155]), .B(n23579), .Z(n24048) );
  NANDN U31530 ( .A(n23580), .B(creg[155]), .Z(n24047) );
  NAND U31531 ( .A(n24049), .B(n19304), .Z(n14196) );
  NANDN U31532 ( .A(init), .B(m[156]), .Z(n19304) );
  AND U31533 ( .A(n24050), .B(n24051), .Z(n24049) );
  NAND U31534 ( .A(o[156]), .B(n23579), .Z(n24051) );
  NANDN U31535 ( .A(n23580), .B(creg[156]), .Z(n24050) );
  NAND U31536 ( .A(n24052), .B(n19302), .Z(n14195) );
  NANDN U31537 ( .A(init), .B(m[157]), .Z(n19302) );
  AND U31538 ( .A(n24053), .B(n24054), .Z(n24052) );
  NAND U31539 ( .A(o[157]), .B(n23579), .Z(n24054) );
  NANDN U31540 ( .A(n23580), .B(creg[157]), .Z(n24053) );
  NAND U31541 ( .A(n24055), .B(n19300), .Z(n14194) );
  NANDN U31542 ( .A(init), .B(m[158]), .Z(n19300) );
  AND U31543 ( .A(n24056), .B(n24057), .Z(n24055) );
  NAND U31544 ( .A(o[158]), .B(n23579), .Z(n24057) );
  NANDN U31545 ( .A(n23580), .B(creg[158]), .Z(n24056) );
  NAND U31546 ( .A(n24058), .B(n19298), .Z(n14193) );
  NANDN U31547 ( .A(init), .B(m[159]), .Z(n19298) );
  AND U31548 ( .A(n24059), .B(n24060), .Z(n24058) );
  NAND U31549 ( .A(o[159]), .B(n23579), .Z(n24060) );
  NANDN U31550 ( .A(n23580), .B(creg[159]), .Z(n24059) );
  NAND U31551 ( .A(n24061), .B(n19294), .Z(n14192) );
  NANDN U31552 ( .A(init), .B(m[160]), .Z(n19294) );
  AND U31553 ( .A(n24062), .B(n24063), .Z(n24061) );
  NAND U31554 ( .A(o[160]), .B(n23579), .Z(n24063) );
  NANDN U31555 ( .A(n23580), .B(creg[160]), .Z(n24062) );
  NAND U31556 ( .A(n24064), .B(n19292), .Z(n14191) );
  NANDN U31557 ( .A(init), .B(m[161]), .Z(n19292) );
  AND U31558 ( .A(n24065), .B(n24066), .Z(n24064) );
  NAND U31559 ( .A(o[161]), .B(n23579), .Z(n24066) );
  NANDN U31560 ( .A(n23580), .B(creg[161]), .Z(n24065) );
  NAND U31561 ( .A(n24067), .B(n19290), .Z(n14190) );
  NANDN U31562 ( .A(init), .B(m[162]), .Z(n19290) );
  AND U31563 ( .A(n24068), .B(n24069), .Z(n24067) );
  NAND U31564 ( .A(o[162]), .B(n23579), .Z(n24069) );
  NANDN U31565 ( .A(n23580), .B(creg[162]), .Z(n24068) );
  NAND U31566 ( .A(n24070), .B(n19288), .Z(n14189) );
  NANDN U31567 ( .A(init), .B(m[163]), .Z(n19288) );
  AND U31568 ( .A(n24071), .B(n24072), .Z(n24070) );
  NAND U31569 ( .A(o[163]), .B(n23579), .Z(n24072) );
  NANDN U31570 ( .A(n23580), .B(creg[163]), .Z(n24071) );
  NAND U31571 ( .A(n24073), .B(n19286), .Z(n14188) );
  NANDN U31572 ( .A(init), .B(m[164]), .Z(n19286) );
  AND U31573 ( .A(n24074), .B(n24075), .Z(n24073) );
  NAND U31574 ( .A(o[164]), .B(n23579), .Z(n24075) );
  NANDN U31575 ( .A(n23580), .B(creg[164]), .Z(n24074) );
  NAND U31576 ( .A(n24076), .B(n19284), .Z(n14187) );
  NANDN U31577 ( .A(init), .B(m[165]), .Z(n19284) );
  AND U31578 ( .A(n24077), .B(n24078), .Z(n24076) );
  NAND U31579 ( .A(o[165]), .B(n23579), .Z(n24078) );
  NANDN U31580 ( .A(n23580), .B(creg[165]), .Z(n24077) );
  NAND U31581 ( .A(n24079), .B(n19282), .Z(n14186) );
  NANDN U31582 ( .A(init), .B(m[166]), .Z(n19282) );
  AND U31583 ( .A(n24080), .B(n24081), .Z(n24079) );
  NAND U31584 ( .A(o[166]), .B(n23579), .Z(n24081) );
  NANDN U31585 ( .A(n23580), .B(creg[166]), .Z(n24080) );
  NAND U31586 ( .A(n24082), .B(n19280), .Z(n14185) );
  NANDN U31587 ( .A(init), .B(m[167]), .Z(n19280) );
  AND U31588 ( .A(n24083), .B(n24084), .Z(n24082) );
  NAND U31589 ( .A(o[167]), .B(n23579), .Z(n24084) );
  NANDN U31590 ( .A(n23580), .B(creg[167]), .Z(n24083) );
  NAND U31591 ( .A(n24085), .B(n19278), .Z(n14184) );
  NANDN U31592 ( .A(init), .B(m[168]), .Z(n19278) );
  AND U31593 ( .A(n24086), .B(n24087), .Z(n24085) );
  NAND U31594 ( .A(o[168]), .B(n23579), .Z(n24087) );
  NANDN U31595 ( .A(n23580), .B(creg[168]), .Z(n24086) );
  NAND U31596 ( .A(n24088), .B(n19276), .Z(n14183) );
  NANDN U31597 ( .A(init), .B(m[169]), .Z(n19276) );
  AND U31598 ( .A(n24089), .B(n24090), .Z(n24088) );
  NAND U31599 ( .A(o[169]), .B(n23579), .Z(n24090) );
  NANDN U31600 ( .A(n23580), .B(creg[169]), .Z(n24089) );
  NAND U31601 ( .A(n24091), .B(n19272), .Z(n14182) );
  NANDN U31602 ( .A(init), .B(m[170]), .Z(n19272) );
  AND U31603 ( .A(n24092), .B(n24093), .Z(n24091) );
  NAND U31604 ( .A(o[170]), .B(n23579), .Z(n24093) );
  NANDN U31605 ( .A(n23580), .B(creg[170]), .Z(n24092) );
  NAND U31606 ( .A(n24094), .B(n19270), .Z(n14181) );
  NANDN U31607 ( .A(init), .B(m[171]), .Z(n19270) );
  AND U31608 ( .A(n24095), .B(n24096), .Z(n24094) );
  NAND U31609 ( .A(o[171]), .B(n23579), .Z(n24096) );
  NANDN U31610 ( .A(n23580), .B(creg[171]), .Z(n24095) );
  NAND U31611 ( .A(n24097), .B(n19268), .Z(n14180) );
  NANDN U31612 ( .A(init), .B(m[172]), .Z(n19268) );
  AND U31613 ( .A(n24098), .B(n24099), .Z(n24097) );
  NAND U31614 ( .A(o[172]), .B(n23579), .Z(n24099) );
  NANDN U31615 ( .A(n23580), .B(creg[172]), .Z(n24098) );
  NAND U31616 ( .A(n24100), .B(n19266), .Z(n14179) );
  NANDN U31617 ( .A(init), .B(m[173]), .Z(n19266) );
  AND U31618 ( .A(n24101), .B(n24102), .Z(n24100) );
  NAND U31619 ( .A(o[173]), .B(n23579), .Z(n24102) );
  NANDN U31620 ( .A(n23580), .B(creg[173]), .Z(n24101) );
  NAND U31621 ( .A(n24103), .B(n19264), .Z(n14178) );
  NANDN U31622 ( .A(init), .B(m[174]), .Z(n19264) );
  AND U31623 ( .A(n24104), .B(n24105), .Z(n24103) );
  NAND U31624 ( .A(o[174]), .B(n23579), .Z(n24105) );
  NANDN U31625 ( .A(n23580), .B(creg[174]), .Z(n24104) );
  NAND U31626 ( .A(n24106), .B(n19262), .Z(n14177) );
  NANDN U31627 ( .A(init), .B(m[175]), .Z(n19262) );
  AND U31628 ( .A(n24107), .B(n24108), .Z(n24106) );
  NAND U31629 ( .A(o[175]), .B(n23579), .Z(n24108) );
  NANDN U31630 ( .A(n23580), .B(creg[175]), .Z(n24107) );
  NAND U31631 ( .A(n24109), .B(n19260), .Z(n14176) );
  NANDN U31632 ( .A(init), .B(m[176]), .Z(n19260) );
  AND U31633 ( .A(n24110), .B(n24111), .Z(n24109) );
  NAND U31634 ( .A(o[176]), .B(n23579), .Z(n24111) );
  NANDN U31635 ( .A(n23580), .B(creg[176]), .Z(n24110) );
  NAND U31636 ( .A(n24112), .B(n19258), .Z(n14175) );
  NANDN U31637 ( .A(init), .B(m[177]), .Z(n19258) );
  AND U31638 ( .A(n24113), .B(n24114), .Z(n24112) );
  NAND U31639 ( .A(o[177]), .B(n23579), .Z(n24114) );
  NANDN U31640 ( .A(n23580), .B(creg[177]), .Z(n24113) );
  NAND U31641 ( .A(n24115), .B(n19256), .Z(n14174) );
  NANDN U31642 ( .A(init), .B(m[178]), .Z(n19256) );
  AND U31643 ( .A(n24116), .B(n24117), .Z(n24115) );
  NAND U31644 ( .A(o[178]), .B(n23579), .Z(n24117) );
  NANDN U31645 ( .A(n23580), .B(creg[178]), .Z(n24116) );
  NAND U31646 ( .A(n24118), .B(n19254), .Z(n14173) );
  NANDN U31647 ( .A(init), .B(m[179]), .Z(n19254) );
  AND U31648 ( .A(n24119), .B(n24120), .Z(n24118) );
  NAND U31649 ( .A(o[179]), .B(n23579), .Z(n24120) );
  NANDN U31650 ( .A(n23580), .B(creg[179]), .Z(n24119) );
  NAND U31651 ( .A(n24121), .B(n19250), .Z(n14172) );
  NANDN U31652 ( .A(init), .B(m[180]), .Z(n19250) );
  AND U31653 ( .A(n24122), .B(n24123), .Z(n24121) );
  NAND U31654 ( .A(o[180]), .B(n23579), .Z(n24123) );
  NANDN U31655 ( .A(n23580), .B(creg[180]), .Z(n24122) );
  NAND U31656 ( .A(n24124), .B(n19248), .Z(n14171) );
  NANDN U31657 ( .A(init), .B(m[181]), .Z(n19248) );
  AND U31658 ( .A(n24125), .B(n24126), .Z(n24124) );
  NAND U31659 ( .A(o[181]), .B(n23579), .Z(n24126) );
  NANDN U31660 ( .A(n23580), .B(creg[181]), .Z(n24125) );
  NAND U31661 ( .A(n24127), .B(n19246), .Z(n14170) );
  NANDN U31662 ( .A(init), .B(m[182]), .Z(n19246) );
  AND U31663 ( .A(n24128), .B(n24129), .Z(n24127) );
  NAND U31664 ( .A(o[182]), .B(n23579), .Z(n24129) );
  NANDN U31665 ( .A(n23580), .B(creg[182]), .Z(n24128) );
  NAND U31666 ( .A(n24130), .B(n19244), .Z(n14169) );
  NANDN U31667 ( .A(init), .B(m[183]), .Z(n19244) );
  AND U31668 ( .A(n24131), .B(n24132), .Z(n24130) );
  NAND U31669 ( .A(o[183]), .B(n23579), .Z(n24132) );
  NANDN U31670 ( .A(n23580), .B(creg[183]), .Z(n24131) );
  NAND U31671 ( .A(n24133), .B(n19242), .Z(n14168) );
  NANDN U31672 ( .A(init), .B(m[184]), .Z(n19242) );
  AND U31673 ( .A(n24134), .B(n24135), .Z(n24133) );
  NAND U31674 ( .A(o[184]), .B(n23579), .Z(n24135) );
  NANDN U31675 ( .A(n23580), .B(creg[184]), .Z(n24134) );
  NAND U31676 ( .A(n24136), .B(n19240), .Z(n14167) );
  NANDN U31677 ( .A(init), .B(m[185]), .Z(n19240) );
  AND U31678 ( .A(n24137), .B(n24138), .Z(n24136) );
  NAND U31679 ( .A(o[185]), .B(n23579), .Z(n24138) );
  NANDN U31680 ( .A(n23580), .B(creg[185]), .Z(n24137) );
  NAND U31681 ( .A(n24139), .B(n19238), .Z(n14166) );
  NANDN U31682 ( .A(init), .B(m[186]), .Z(n19238) );
  AND U31683 ( .A(n24140), .B(n24141), .Z(n24139) );
  NAND U31684 ( .A(o[186]), .B(n23579), .Z(n24141) );
  NANDN U31685 ( .A(n23580), .B(creg[186]), .Z(n24140) );
  NAND U31686 ( .A(n24142), .B(n19236), .Z(n14165) );
  NANDN U31687 ( .A(init), .B(m[187]), .Z(n19236) );
  AND U31688 ( .A(n24143), .B(n24144), .Z(n24142) );
  NAND U31689 ( .A(o[187]), .B(n23579), .Z(n24144) );
  NANDN U31690 ( .A(n23580), .B(creg[187]), .Z(n24143) );
  NAND U31691 ( .A(n24145), .B(n19234), .Z(n14164) );
  NANDN U31692 ( .A(init), .B(m[188]), .Z(n19234) );
  AND U31693 ( .A(n24146), .B(n24147), .Z(n24145) );
  NAND U31694 ( .A(o[188]), .B(n23579), .Z(n24147) );
  NANDN U31695 ( .A(n23580), .B(creg[188]), .Z(n24146) );
  NAND U31696 ( .A(n24148), .B(n19232), .Z(n14163) );
  NANDN U31697 ( .A(init), .B(m[189]), .Z(n19232) );
  AND U31698 ( .A(n24149), .B(n24150), .Z(n24148) );
  NAND U31699 ( .A(o[189]), .B(n23579), .Z(n24150) );
  NANDN U31700 ( .A(n23580), .B(creg[189]), .Z(n24149) );
  NAND U31701 ( .A(n24151), .B(n19228), .Z(n14162) );
  NANDN U31702 ( .A(init), .B(m[190]), .Z(n19228) );
  AND U31703 ( .A(n24152), .B(n24153), .Z(n24151) );
  NAND U31704 ( .A(o[190]), .B(n23579), .Z(n24153) );
  NANDN U31705 ( .A(n23580), .B(creg[190]), .Z(n24152) );
  NAND U31706 ( .A(n24154), .B(n19226), .Z(n14161) );
  NANDN U31707 ( .A(init), .B(m[191]), .Z(n19226) );
  AND U31708 ( .A(n24155), .B(n24156), .Z(n24154) );
  NAND U31709 ( .A(o[191]), .B(n23579), .Z(n24156) );
  NANDN U31710 ( .A(n23580), .B(creg[191]), .Z(n24155) );
  NAND U31711 ( .A(n24157), .B(n19224), .Z(n14160) );
  NANDN U31712 ( .A(init), .B(m[192]), .Z(n19224) );
  AND U31713 ( .A(n24158), .B(n24159), .Z(n24157) );
  NAND U31714 ( .A(o[192]), .B(n23579), .Z(n24159) );
  NANDN U31715 ( .A(n23580), .B(creg[192]), .Z(n24158) );
  NAND U31716 ( .A(n24160), .B(n19222), .Z(n14159) );
  NANDN U31717 ( .A(init), .B(m[193]), .Z(n19222) );
  AND U31718 ( .A(n24161), .B(n24162), .Z(n24160) );
  NAND U31719 ( .A(o[193]), .B(n23579), .Z(n24162) );
  NANDN U31720 ( .A(n23580), .B(creg[193]), .Z(n24161) );
  NAND U31721 ( .A(n24163), .B(n19220), .Z(n14158) );
  NANDN U31722 ( .A(init), .B(m[194]), .Z(n19220) );
  AND U31723 ( .A(n24164), .B(n24165), .Z(n24163) );
  NAND U31724 ( .A(o[194]), .B(n23579), .Z(n24165) );
  NANDN U31725 ( .A(n23580), .B(creg[194]), .Z(n24164) );
  NAND U31726 ( .A(n24166), .B(n19218), .Z(n14157) );
  NANDN U31727 ( .A(init), .B(m[195]), .Z(n19218) );
  AND U31728 ( .A(n24167), .B(n24168), .Z(n24166) );
  NAND U31729 ( .A(o[195]), .B(n23579), .Z(n24168) );
  NANDN U31730 ( .A(n23580), .B(creg[195]), .Z(n24167) );
  NAND U31731 ( .A(n24169), .B(n19216), .Z(n14156) );
  NANDN U31732 ( .A(init), .B(m[196]), .Z(n19216) );
  AND U31733 ( .A(n24170), .B(n24171), .Z(n24169) );
  NAND U31734 ( .A(o[196]), .B(n23579), .Z(n24171) );
  NANDN U31735 ( .A(n23580), .B(creg[196]), .Z(n24170) );
  NAND U31736 ( .A(n24172), .B(n19214), .Z(n14155) );
  NANDN U31737 ( .A(init), .B(m[197]), .Z(n19214) );
  AND U31738 ( .A(n24173), .B(n24174), .Z(n24172) );
  NAND U31739 ( .A(o[197]), .B(n23579), .Z(n24174) );
  NANDN U31740 ( .A(n23580), .B(creg[197]), .Z(n24173) );
  NAND U31741 ( .A(n24175), .B(n19212), .Z(n14154) );
  NANDN U31742 ( .A(init), .B(m[198]), .Z(n19212) );
  AND U31743 ( .A(n24176), .B(n24177), .Z(n24175) );
  NAND U31744 ( .A(o[198]), .B(n23579), .Z(n24177) );
  NANDN U31745 ( .A(n23580), .B(creg[198]), .Z(n24176) );
  NAND U31746 ( .A(n24178), .B(n19210), .Z(n14153) );
  NANDN U31747 ( .A(init), .B(m[199]), .Z(n19210) );
  AND U31748 ( .A(n24179), .B(n24180), .Z(n24178) );
  NAND U31749 ( .A(o[199]), .B(n23579), .Z(n24180) );
  NANDN U31750 ( .A(n23580), .B(creg[199]), .Z(n24179) );
  NAND U31751 ( .A(n24181), .B(n19204), .Z(n14152) );
  NANDN U31752 ( .A(init), .B(m[200]), .Z(n19204) );
  AND U31753 ( .A(n24182), .B(n24183), .Z(n24181) );
  NAND U31754 ( .A(o[200]), .B(n23579), .Z(n24183) );
  NANDN U31755 ( .A(n23580), .B(creg[200]), .Z(n24182) );
  NAND U31756 ( .A(n24184), .B(n19202), .Z(n14151) );
  NANDN U31757 ( .A(init), .B(m[201]), .Z(n19202) );
  AND U31758 ( .A(n24185), .B(n24186), .Z(n24184) );
  NAND U31759 ( .A(o[201]), .B(n23579), .Z(n24186) );
  NANDN U31760 ( .A(n23580), .B(creg[201]), .Z(n24185) );
  NAND U31761 ( .A(n24187), .B(n19200), .Z(n14150) );
  NANDN U31762 ( .A(init), .B(m[202]), .Z(n19200) );
  AND U31763 ( .A(n24188), .B(n24189), .Z(n24187) );
  NAND U31764 ( .A(o[202]), .B(n23579), .Z(n24189) );
  NANDN U31765 ( .A(n23580), .B(creg[202]), .Z(n24188) );
  NAND U31766 ( .A(n24190), .B(n19198), .Z(n14149) );
  NANDN U31767 ( .A(init), .B(m[203]), .Z(n19198) );
  AND U31768 ( .A(n24191), .B(n24192), .Z(n24190) );
  NAND U31769 ( .A(o[203]), .B(n23579), .Z(n24192) );
  NANDN U31770 ( .A(n23580), .B(creg[203]), .Z(n24191) );
  NAND U31771 ( .A(n24193), .B(n19196), .Z(n14148) );
  NANDN U31772 ( .A(init), .B(m[204]), .Z(n19196) );
  AND U31773 ( .A(n24194), .B(n24195), .Z(n24193) );
  NAND U31774 ( .A(o[204]), .B(n23579), .Z(n24195) );
  NANDN U31775 ( .A(n23580), .B(creg[204]), .Z(n24194) );
  NAND U31776 ( .A(n24196), .B(n19194), .Z(n14147) );
  NANDN U31777 ( .A(init), .B(m[205]), .Z(n19194) );
  AND U31778 ( .A(n24197), .B(n24198), .Z(n24196) );
  NAND U31779 ( .A(o[205]), .B(n23579), .Z(n24198) );
  NANDN U31780 ( .A(n23580), .B(creg[205]), .Z(n24197) );
  NAND U31781 ( .A(n24199), .B(n19192), .Z(n14146) );
  NANDN U31782 ( .A(init), .B(m[206]), .Z(n19192) );
  AND U31783 ( .A(n24200), .B(n24201), .Z(n24199) );
  NAND U31784 ( .A(o[206]), .B(n23579), .Z(n24201) );
  NANDN U31785 ( .A(n23580), .B(creg[206]), .Z(n24200) );
  NAND U31786 ( .A(n24202), .B(n19190), .Z(n14145) );
  NANDN U31787 ( .A(init), .B(m[207]), .Z(n19190) );
  AND U31788 ( .A(n24203), .B(n24204), .Z(n24202) );
  NAND U31789 ( .A(o[207]), .B(n23579), .Z(n24204) );
  NANDN U31790 ( .A(n23580), .B(creg[207]), .Z(n24203) );
  NAND U31791 ( .A(n24205), .B(n19188), .Z(n14144) );
  NANDN U31792 ( .A(init), .B(m[208]), .Z(n19188) );
  AND U31793 ( .A(n24206), .B(n24207), .Z(n24205) );
  NAND U31794 ( .A(o[208]), .B(n23579), .Z(n24207) );
  NANDN U31795 ( .A(n23580), .B(creg[208]), .Z(n24206) );
  NAND U31796 ( .A(n24208), .B(n19186), .Z(n14143) );
  NANDN U31797 ( .A(init), .B(m[209]), .Z(n19186) );
  AND U31798 ( .A(n24209), .B(n24210), .Z(n24208) );
  NAND U31799 ( .A(o[209]), .B(n23579), .Z(n24210) );
  NANDN U31800 ( .A(n23580), .B(creg[209]), .Z(n24209) );
  NAND U31801 ( .A(n24211), .B(n19182), .Z(n14142) );
  NANDN U31802 ( .A(init), .B(m[210]), .Z(n19182) );
  AND U31803 ( .A(n24212), .B(n24213), .Z(n24211) );
  NAND U31804 ( .A(o[210]), .B(n23579), .Z(n24213) );
  NANDN U31805 ( .A(n23580), .B(creg[210]), .Z(n24212) );
  NAND U31806 ( .A(n24214), .B(n19180), .Z(n14141) );
  NANDN U31807 ( .A(init), .B(m[211]), .Z(n19180) );
  AND U31808 ( .A(n24215), .B(n24216), .Z(n24214) );
  NAND U31809 ( .A(o[211]), .B(n23579), .Z(n24216) );
  NANDN U31810 ( .A(n23580), .B(creg[211]), .Z(n24215) );
  NAND U31811 ( .A(n24217), .B(n19178), .Z(n14140) );
  NANDN U31812 ( .A(init), .B(m[212]), .Z(n19178) );
  AND U31813 ( .A(n24218), .B(n24219), .Z(n24217) );
  NAND U31814 ( .A(o[212]), .B(n23579), .Z(n24219) );
  NANDN U31815 ( .A(n23580), .B(creg[212]), .Z(n24218) );
  NAND U31816 ( .A(n24220), .B(n19176), .Z(n14139) );
  NANDN U31817 ( .A(init), .B(m[213]), .Z(n19176) );
  AND U31818 ( .A(n24221), .B(n24222), .Z(n24220) );
  NAND U31819 ( .A(o[213]), .B(n23579), .Z(n24222) );
  NANDN U31820 ( .A(n23580), .B(creg[213]), .Z(n24221) );
  NAND U31821 ( .A(n24223), .B(n19174), .Z(n14138) );
  NANDN U31822 ( .A(init), .B(m[214]), .Z(n19174) );
  AND U31823 ( .A(n24224), .B(n24225), .Z(n24223) );
  NAND U31824 ( .A(o[214]), .B(n23579), .Z(n24225) );
  NANDN U31825 ( .A(n23580), .B(creg[214]), .Z(n24224) );
  NAND U31826 ( .A(n24226), .B(n19172), .Z(n14137) );
  NANDN U31827 ( .A(init), .B(m[215]), .Z(n19172) );
  AND U31828 ( .A(n24227), .B(n24228), .Z(n24226) );
  NAND U31829 ( .A(o[215]), .B(n23579), .Z(n24228) );
  NANDN U31830 ( .A(n23580), .B(creg[215]), .Z(n24227) );
  NAND U31831 ( .A(n24229), .B(n19170), .Z(n14136) );
  NANDN U31832 ( .A(init), .B(m[216]), .Z(n19170) );
  AND U31833 ( .A(n24230), .B(n24231), .Z(n24229) );
  NAND U31834 ( .A(o[216]), .B(n23579), .Z(n24231) );
  NANDN U31835 ( .A(n23580), .B(creg[216]), .Z(n24230) );
  NAND U31836 ( .A(n24232), .B(n19168), .Z(n14135) );
  NANDN U31837 ( .A(init), .B(m[217]), .Z(n19168) );
  AND U31838 ( .A(n24233), .B(n24234), .Z(n24232) );
  NAND U31839 ( .A(o[217]), .B(n23579), .Z(n24234) );
  NANDN U31840 ( .A(n23580), .B(creg[217]), .Z(n24233) );
  NAND U31841 ( .A(n24235), .B(n19166), .Z(n14134) );
  NANDN U31842 ( .A(init), .B(m[218]), .Z(n19166) );
  AND U31843 ( .A(n24236), .B(n24237), .Z(n24235) );
  NAND U31844 ( .A(o[218]), .B(n23579), .Z(n24237) );
  NANDN U31845 ( .A(n23580), .B(creg[218]), .Z(n24236) );
  NAND U31846 ( .A(n24238), .B(n19164), .Z(n14133) );
  NANDN U31847 ( .A(init), .B(m[219]), .Z(n19164) );
  AND U31848 ( .A(n24239), .B(n24240), .Z(n24238) );
  NAND U31849 ( .A(o[219]), .B(n23579), .Z(n24240) );
  NANDN U31850 ( .A(n23580), .B(creg[219]), .Z(n24239) );
  NAND U31851 ( .A(n24241), .B(n19160), .Z(n14132) );
  NANDN U31852 ( .A(init), .B(m[220]), .Z(n19160) );
  AND U31853 ( .A(n24242), .B(n24243), .Z(n24241) );
  NAND U31854 ( .A(o[220]), .B(n23579), .Z(n24243) );
  NANDN U31855 ( .A(n23580), .B(creg[220]), .Z(n24242) );
  NAND U31856 ( .A(n24244), .B(n19158), .Z(n14131) );
  NANDN U31857 ( .A(init), .B(m[221]), .Z(n19158) );
  AND U31858 ( .A(n24245), .B(n24246), .Z(n24244) );
  NAND U31859 ( .A(o[221]), .B(n23579), .Z(n24246) );
  NANDN U31860 ( .A(n23580), .B(creg[221]), .Z(n24245) );
  NAND U31861 ( .A(n24247), .B(n19156), .Z(n14130) );
  NANDN U31862 ( .A(init), .B(m[222]), .Z(n19156) );
  AND U31863 ( .A(n24248), .B(n24249), .Z(n24247) );
  NAND U31864 ( .A(o[222]), .B(n23579), .Z(n24249) );
  NANDN U31865 ( .A(n23580), .B(creg[222]), .Z(n24248) );
  NAND U31866 ( .A(n24250), .B(n19154), .Z(n14129) );
  NANDN U31867 ( .A(init), .B(m[223]), .Z(n19154) );
  AND U31868 ( .A(n24251), .B(n24252), .Z(n24250) );
  NAND U31869 ( .A(o[223]), .B(n23579), .Z(n24252) );
  NANDN U31870 ( .A(n23580), .B(creg[223]), .Z(n24251) );
  NAND U31871 ( .A(n24253), .B(n19152), .Z(n14128) );
  NANDN U31872 ( .A(init), .B(m[224]), .Z(n19152) );
  AND U31873 ( .A(n24254), .B(n24255), .Z(n24253) );
  NAND U31874 ( .A(o[224]), .B(n23579), .Z(n24255) );
  NANDN U31875 ( .A(n23580), .B(creg[224]), .Z(n24254) );
  NAND U31876 ( .A(n24256), .B(n19150), .Z(n14127) );
  NANDN U31877 ( .A(init), .B(m[225]), .Z(n19150) );
  AND U31878 ( .A(n24257), .B(n24258), .Z(n24256) );
  NAND U31879 ( .A(o[225]), .B(n23579), .Z(n24258) );
  NANDN U31880 ( .A(n23580), .B(creg[225]), .Z(n24257) );
  NAND U31881 ( .A(n24259), .B(n19148), .Z(n14126) );
  NANDN U31882 ( .A(init), .B(m[226]), .Z(n19148) );
  AND U31883 ( .A(n24260), .B(n24261), .Z(n24259) );
  NAND U31884 ( .A(o[226]), .B(n23579), .Z(n24261) );
  NANDN U31885 ( .A(n23580), .B(creg[226]), .Z(n24260) );
  NAND U31886 ( .A(n24262), .B(n19146), .Z(n14125) );
  NANDN U31887 ( .A(init), .B(m[227]), .Z(n19146) );
  AND U31888 ( .A(n24263), .B(n24264), .Z(n24262) );
  NAND U31889 ( .A(o[227]), .B(n23579), .Z(n24264) );
  NANDN U31890 ( .A(n23580), .B(creg[227]), .Z(n24263) );
  NAND U31891 ( .A(n24265), .B(n19144), .Z(n14124) );
  NANDN U31892 ( .A(init), .B(m[228]), .Z(n19144) );
  AND U31893 ( .A(n24266), .B(n24267), .Z(n24265) );
  NAND U31894 ( .A(o[228]), .B(n23579), .Z(n24267) );
  NANDN U31895 ( .A(n23580), .B(creg[228]), .Z(n24266) );
  NAND U31896 ( .A(n24268), .B(n19142), .Z(n14123) );
  NANDN U31897 ( .A(init), .B(m[229]), .Z(n19142) );
  AND U31898 ( .A(n24269), .B(n24270), .Z(n24268) );
  NAND U31899 ( .A(o[229]), .B(n23579), .Z(n24270) );
  NANDN U31900 ( .A(n23580), .B(creg[229]), .Z(n24269) );
  NAND U31901 ( .A(n24271), .B(n19138), .Z(n14122) );
  NANDN U31902 ( .A(init), .B(m[230]), .Z(n19138) );
  AND U31903 ( .A(n24272), .B(n24273), .Z(n24271) );
  NAND U31904 ( .A(o[230]), .B(n23579), .Z(n24273) );
  NANDN U31905 ( .A(n23580), .B(creg[230]), .Z(n24272) );
  NAND U31906 ( .A(n24274), .B(n19136), .Z(n14121) );
  NANDN U31907 ( .A(init), .B(m[231]), .Z(n19136) );
  AND U31908 ( .A(n24275), .B(n24276), .Z(n24274) );
  NAND U31909 ( .A(o[231]), .B(n23579), .Z(n24276) );
  NANDN U31910 ( .A(n23580), .B(creg[231]), .Z(n24275) );
  NAND U31911 ( .A(n24277), .B(n19134), .Z(n14120) );
  NANDN U31912 ( .A(init), .B(m[232]), .Z(n19134) );
  AND U31913 ( .A(n24278), .B(n24279), .Z(n24277) );
  NAND U31914 ( .A(o[232]), .B(n23579), .Z(n24279) );
  NANDN U31915 ( .A(n23580), .B(creg[232]), .Z(n24278) );
  NAND U31916 ( .A(n24280), .B(n19132), .Z(n14119) );
  NANDN U31917 ( .A(init), .B(m[233]), .Z(n19132) );
  AND U31918 ( .A(n24281), .B(n24282), .Z(n24280) );
  NAND U31919 ( .A(o[233]), .B(n23579), .Z(n24282) );
  NANDN U31920 ( .A(n23580), .B(creg[233]), .Z(n24281) );
  NAND U31921 ( .A(n24283), .B(n19130), .Z(n14118) );
  NANDN U31922 ( .A(init), .B(m[234]), .Z(n19130) );
  AND U31923 ( .A(n24284), .B(n24285), .Z(n24283) );
  NAND U31924 ( .A(o[234]), .B(n23579), .Z(n24285) );
  NANDN U31925 ( .A(n23580), .B(creg[234]), .Z(n24284) );
  NAND U31926 ( .A(n24286), .B(n19128), .Z(n14117) );
  NANDN U31927 ( .A(init), .B(m[235]), .Z(n19128) );
  AND U31928 ( .A(n24287), .B(n24288), .Z(n24286) );
  NAND U31929 ( .A(o[235]), .B(n23579), .Z(n24288) );
  NANDN U31930 ( .A(n23580), .B(creg[235]), .Z(n24287) );
  NAND U31931 ( .A(n24289), .B(n19126), .Z(n14116) );
  NANDN U31932 ( .A(init), .B(m[236]), .Z(n19126) );
  AND U31933 ( .A(n24290), .B(n24291), .Z(n24289) );
  NAND U31934 ( .A(o[236]), .B(n23579), .Z(n24291) );
  NANDN U31935 ( .A(n23580), .B(creg[236]), .Z(n24290) );
  NAND U31936 ( .A(n24292), .B(n19124), .Z(n14115) );
  NANDN U31937 ( .A(init), .B(m[237]), .Z(n19124) );
  AND U31938 ( .A(n24293), .B(n24294), .Z(n24292) );
  NAND U31939 ( .A(o[237]), .B(n23579), .Z(n24294) );
  NANDN U31940 ( .A(n23580), .B(creg[237]), .Z(n24293) );
  NAND U31941 ( .A(n24295), .B(n19122), .Z(n14114) );
  NANDN U31942 ( .A(init), .B(m[238]), .Z(n19122) );
  AND U31943 ( .A(n24296), .B(n24297), .Z(n24295) );
  NAND U31944 ( .A(o[238]), .B(n23579), .Z(n24297) );
  NANDN U31945 ( .A(n23580), .B(creg[238]), .Z(n24296) );
  NAND U31946 ( .A(n24298), .B(n19120), .Z(n14113) );
  NANDN U31947 ( .A(init), .B(m[239]), .Z(n19120) );
  AND U31948 ( .A(n24299), .B(n24300), .Z(n24298) );
  NAND U31949 ( .A(o[239]), .B(n23579), .Z(n24300) );
  NANDN U31950 ( .A(n23580), .B(creg[239]), .Z(n24299) );
  NAND U31951 ( .A(n24301), .B(n19116), .Z(n14112) );
  NANDN U31952 ( .A(init), .B(m[240]), .Z(n19116) );
  AND U31953 ( .A(n24302), .B(n24303), .Z(n24301) );
  NAND U31954 ( .A(o[240]), .B(n23579), .Z(n24303) );
  NANDN U31955 ( .A(n23580), .B(creg[240]), .Z(n24302) );
  NAND U31956 ( .A(n24304), .B(n19114), .Z(n14111) );
  NANDN U31957 ( .A(init), .B(m[241]), .Z(n19114) );
  AND U31958 ( .A(n24305), .B(n24306), .Z(n24304) );
  NAND U31959 ( .A(o[241]), .B(n23579), .Z(n24306) );
  NANDN U31960 ( .A(n23580), .B(creg[241]), .Z(n24305) );
  NAND U31961 ( .A(n24307), .B(n19112), .Z(n14110) );
  NANDN U31962 ( .A(init), .B(m[242]), .Z(n19112) );
  AND U31963 ( .A(n24308), .B(n24309), .Z(n24307) );
  NAND U31964 ( .A(o[242]), .B(n23579), .Z(n24309) );
  NANDN U31965 ( .A(n23580), .B(creg[242]), .Z(n24308) );
  NAND U31966 ( .A(n24310), .B(n19110), .Z(n14109) );
  NANDN U31967 ( .A(init), .B(m[243]), .Z(n19110) );
  AND U31968 ( .A(n24311), .B(n24312), .Z(n24310) );
  NAND U31969 ( .A(o[243]), .B(n23579), .Z(n24312) );
  NANDN U31970 ( .A(n23580), .B(creg[243]), .Z(n24311) );
  NAND U31971 ( .A(n24313), .B(n19108), .Z(n14108) );
  NANDN U31972 ( .A(init), .B(m[244]), .Z(n19108) );
  AND U31973 ( .A(n24314), .B(n24315), .Z(n24313) );
  NAND U31974 ( .A(o[244]), .B(n23579), .Z(n24315) );
  NANDN U31975 ( .A(n23580), .B(creg[244]), .Z(n24314) );
  NAND U31976 ( .A(n24316), .B(n19106), .Z(n14107) );
  NANDN U31977 ( .A(init), .B(m[245]), .Z(n19106) );
  AND U31978 ( .A(n24317), .B(n24318), .Z(n24316) );
  NAND U31979 ( .A(o[245]), .B(n23579), .Z(n24318) );
  NANDN U31980 ( .A(n23580), .B(creg[245]), .Z(n24317) );
  NAND U31981 ( .A(n24319), .B(n19104), .Z(n14106) );
  NANDN U31982 ( .A(init), .B(m[246]), .Z(n19104) );
  AND U31983 ( .A(n24320), .B(n24321), .Z(n24319) );
  NAND U31984 ( .A(o[246]), .B(n23579), .Z(n24321) );
  NANDN U31985 ( .A(n23580), .B(creg[246]), .Z(n24320) );
  NAND U31986 ( .A(n24322), .B(n19102), .Z(n14105) );
  NANDN U31987 ( .A(init), .B(m[247]), .Z(n19102) );
  AND U31988 ( .A(n24323), .B(n24324), .Z(n24322) );
  NAND U31989 ( .A(o[247]), .B(n23579), .Z(n24324) );
  NANDN U31990 ( .A(n23580), .B(creg[247]), .Z(n24323) );
  NAND U31991 ( .A(n24325), .B(n19100), .Z(n14104) );
  NANDN U31992 ( .A(init), .B(m[248]), .Z(n19100) );
  AND U31993 ( .A(n24326), .B(n24327), .Z(n24325) );
  NAND U31994 ( .A(o[248]), .B(n23579), .Z(n24327) );
  NANDN U31995 ( .A(n23580), .B(creg[248]), .Z(n24326) );
  NAND U31996 ( .A(n24328), .B(n19098), .Z(n14103) );
  NANDN U31997 ( .A(init), .B(m[249]), .Z(n19098) );
  AND U31998 ( .A(n24329), .B(n24330), .Z(n24328) );
  NAND U31999 ( .A(o[249]), .B(n23579), .Z(n24330) );
  NANDN U32000 ( .A(n23580), .B(creg[249]), .Z(n24329) );
  NAND U32001 ( .A(n24331), .B(n19094), .Z(n14102) );
  NANDN U32002 ( .A(init), .B(m[250]), .Z(n19094) );
  AND U32003 ( .A(n24332), .B(n24333), .Z(n24331) );
  NAND U32004 ( .A(o[250]), .B(n23579), .Z(n24333) );
  NANDN U32005 ( .A(n23580), .B(creg[250]), .Z(n24332) );
  NAND U32006 ( .A(n24334), .B(n19092), .Z(n14101) );
  NANDN U32007 ( .A(init), .B(m[251]), .Z(n19092) );
  AND U32008 ( .A(n24335), .B(n24336), .Z(n24334) );
  NAND U32009 ( .A(o[251]), .B(n23579), .Z(n24336) );
  NANDN U32010 ( .A(n23580), .B(creg[251]), .Z(n24335) );
  NAND U32011 ( .A(n24337), .B(n19090), .Z(n14100) );
  NANDN U32012 ( .A(init), .B(m[252]), .Z(n19090) );
  AND U32013 ( .A(n24338), .B(n24339), .Z(n24337) );
  NAND U32014 ( .A(o[252]), .B(n23579), .Z(n24339) );
  NANDN U32015 ( .A(n23580), .B(creg[252]), .Z(n24338) );
  NAND U32016 ( .A(n24340), .B(n19088), .Z(n14099) );
  NANDN U32017 ( .A(init), .B(m[253]), .Z(n19088) );
  AND U32018 ( .A(n24341), .B(n24342), .Z(n24340) );
  NAND U32019 ( .A(o[253]), .B(n23579), .Z(n24342) );
  NANDN U32020 ( .A(n23580), .B(creg[253]), .Z(n24341) );
  NAND U32021 ( .A(n24343), .B(n19086), .Z(n14098) );
  NANDN U32022 ( .A(init), .B(m[254]), .Z(n19086) );
  AND U32023 ( .A(n24344), .B(n24345), .Z(n24343) );
  NAND U32024 ( .A(o[254]), .B(n23579), .Z(n24345) );
  NANDN U32025 ( .A(n23580), .B(creg[254]), .Z(n24344) );
  NAND U32026 ( .A(n24346), .B(n19084), .Z(n14097) );
  NANDN U32027 ( .A(init), .B(m[255]), .Z(n19084) );
  AND U32028 ( .A(n24347), .B(n24348), .Z(n24346) );
  NAND U32029 ( .A(o[255]), .B(n23579), .Z(n24348) );
  NANDN U32030 ( .A(n23580), .B(creg[255]), .Z(n24347) );
  NAND U32031 ( .A(n24349), .B(n19082), .Z(n14096) );
  NANDN U32032 ( .A(init), .B(m[256]), .Z(n19082) );
  AND U32033 ( .A(n24350), .B(n24351), .Z(n24349) );
  NAND U32034 ( .A(o[256]), .B(n23579), .Z(n24351) );
  NANDN U32035 ( .A(n23580), .B(creg[256]), .Z(n24350) );
  NAND U32036 ( .A(n24352), .B(n19080), .Z(n14095) );
  NANDN U32037 ( .A(init), .B(m[257]), .Z(n19080) );
  AND U32038 ( .A(n24353), .B(n24354), .Z(n24352) );
  NAND U32039 ( .A(o[257]), .B(n23579), .Z(n24354) );
  NANDN U32040 ( .A(n23580), .B(creg[257]), .Z(n24353) );
  NAND U32041 ( .A(n24355), .B(n19078), .Z(n14094) );
  NANDN U32042 ( .A(init), .B(m[258]), .Z(n19078) );
  AND U32043 ( .A(n24356), .B(n24357), .Z(n24355) );
  NAND U32044 ( .A(o[258]), .B(n23579), .Z(n24357) );
  NANDN U32045 ( .A(n23580), .B(creg[258]), .Z(n24356) );
  NAND U32046 ( .A(n24358), .B(n19076), .Z(n14093) );
  NANDN U32047 ( .A(init), .B(m[259]), .Z(n19076) );
  AND U32048 ( .A(n24359), .B(n24360), .Z(n24358) );
  NAND U32049 ( .A(o[259]), .B(n23579), .Z(n24360) );
  NANDN U32050 ( .A(n23580), .B(creg[259]), .Z(n24359) );
  NAND U32051 ( .A(n24361), .B(n19072), .Z(n14092) );
  NANDN U32052 ( .A(init), .B(m[260]), .Z(n19072) );
  AND U32053 ( .A(n24362), .B(n24363), .Z(n24361) );
  NAND U32054 ( .A(o[260]), .B(n23579), .Z(n24363) );
  NANDN U32055 ( .A(n23580), .B(creg[260]), .Z(n24362) );
  NAND U32056 ( .A(n24364), .B(n19070), .Z(n14091) );
  NANDN U32057 ( .A(init), .B(m[261]), .Z(n19070) );
  AND U32058 ( .A(n24365), .B(n24366), .Z(n24364) );
  NAND U32059 ( .A(o[261]), .B(n23579), .Z(n24366) );
  NANDN U32060 ( .A(n23580), .B(creg[261]), .Z(n24365) );
  NAND U32061 ( .A(n24367), .B(n19068), .Z(n14090) );
  NANDN U32062 ( .A(init), .B(m[262]), .Z(n19068) );
  AND U32063 ( .A(n24368), .B(n24369), .Z(n24367) );
  NAND U32064 ( .A(o[262]), .B(n23579), .Z(n24369) );
  NANDN U32065 ( .A(n23580), .B(creg[262]), .Z(n24368) );
  NAND U32066 ( .A(n24370), .B(n19066), .Z(n14089) );
  NANDN U32067 ( .A(init), .B(m[263]), .Z(n19066) );
  AND U32068 ( .A(n24371), .B(n24372), .Z(n24370) );
  NAND U32069 ( .A(o[263]), .B(n23579), .Z(n24372) );
  NANDN U32070 ( .A(n23580), .B(creg[263]), .Z(n24371) );
  NAND U32071 ( .A(n24373), .B(n19064), .Z(n14088) );
  NANDN U32072 ( .A(init), .B(m[264]), .Z(n19064) );
  AND U32073 ( .A(n24374), .B(n24375), .Z(n24373) );
  NAND U32074 ( .A(o[264]), .B(n23579), .Z(n24375) );
  NANDN U32075 ( .A(n23580), .B(creg[264]), .Z(n24374) );
  NAND U32076 ( .A(n24376), .B(n19062), .Z(n14087) );
  NANDN U32077 ( .A(init), .B(m[265]), .Z(n19062) );
  AND U32078 ( .A(n24377), .B(n24378), .Z(n24376) );
  NAND U32079 ( .A(o[265]), .B(n23579), .Z(n24378) );
  NANDN U32080 ( .A(n23580), .B(creg[265]), .Z(n24377) );
  NAND U32081 ( .A(n24379), .B(n19060), .Z(n14086) );
  NANDN U32082 ( .A(init), .B(m[266]), .Z(n19060) );
  AND U32083 ( .A(n24380), .B(n24381), .Z(n24379) );
  NAND U32084 ( .A(o[266]), .B(n23579), .Z(n24381) );
  NANDN U32085 ( .A(n23580), .B(creg[266]), .Z(n24380) );
  NAND U32086 ( .A(n24382), .B(n19058), .Z(n14085) );
  NANDN U32087 ( .A(init), .B(m[267]), .Z(n19058) );
  AND U32088 ( .A(n24383), .B(n24384), .Z(n24382) );
  NAND U32089 ( .A(o[267]), .B(n23579), .Z(n24384) );
  NANDN U32090 ( .A(n23580), .B(creg[267]), .Z(n24383) );
  NAND U32091 ( .A(n24385), .B(n19056), .Z(n14084) );
  NANDN U32092 ( .A(init), .B(m[268]), .Z(n19056) );
  AND U32093 ( .A(n24386), .B(n24387), .Z(n24385) );
  NAND U32094 ( .A(o[268]), .B(n23579), .Z(n24387) );
  NANDN U32095 ( .A(n23580), .B(creg[268]), .Z(n24386) );
  NAND U32096 ( .A(n24388), .B(n19054), .Z(n14083) );
  NANDN U32097 ( .A(init), .B(m[269]), .Z(n19054) );
  AND U32098 ( .A(n24389), .B(n24390), .Z(n24388) );
  NAND U32099 ( .A(o[269]), .B(n23579), .Z(n24390) );
  NANDN U32100 ( .A(n23580), .B(creg[269]), .Z(n24389) );
  NAND U32101 ( .A(n24391), .B(n19050), .Z(n14082) );
  NANDN U32102 ( .A(init), .B(m[270]), .Z(n19050) );
  AND U32103 ( .A(n24392), .B(n24393), .Z(n24391) );
  NAND U32104 ( .A(o[270]), .B(n23579), .Z(n24393) );
  NANDN U32105 ( .A(n23580), .B(creg[270]), .Z(n24392) );
  NAND U32106 ( .A(n24394), .B(n19048), .Z(n14081) );
  NANDN U32107 ( .A(init), .B(m[271]), .Z(n19048) );
  AND U32108 ( .A(n24395), .B(n24396), .Z(n24394) );
  NAND U32109 ( .A(o[271]), .B(n23579), .Z(n24396) );
  NANDN U32110 ( .A(n23580), .B(creg[271]), .Z(n24395) );
  NAND U32111 ( .A(n24397), .B(n19046), .Z(n14080) );
  NANDN U32112 ( .A(init), .B(m[272]), .Z(n19046) );
  AND U32113 ( .A(n24398), .B(n24399), .Z(n24397) );
  NAND U32114 ( .A(o[272]), .B(n23579), .Z(n24399) );
  NANDN U32115 ( .A(n23580), .B(creg[272]), .Z(n24398) );
  NAND U32116 ( .A(n24400), .B(n19044), .Z(n14079) );
  NANDN U32117 ( .A(init), .B(m[273]), .Z(n19044) );
  AND U32118 ( .A(n24401), .B(n24402), .Z(n24400) );
  NAND U32119 ( .A(o[273]), .B(n23579), .Z(n24402) );
  NANDN U32120 ( .A(n23580), .B(creg[273]), .Z(n24401) );
  NAND U32121 ( .A(n24403), .B(n19042), .Z(n14078) );
  NANDN U32122 ( .A(init), .B(m[274]), .Z(n19042) );
  AND U32123 ( .A(n24404), .B(n24405), .Z(n24403) );
  NAND U32124 ( .A(o[274]), .B(n23579), .Z(n24405) );
  NANDN U32125 ( .A(n23580), .B(creg[274]), .Z(n24404) );
  NAND U32126 ( .A(n24406), .B(n19040), .Z(n14077) );
  NANDN U32127 ( .A(init), .B(m[275]), .Z(n19040) );
  AND U32128 ( .A(n24407), .B(n24408), .Z(n24406) );
  NAND U32129 ( .A(o[275]), .B(n23579), .Z(n24408) );
  NANDN U32130 ( .A(n23580), .B(creg[275]), .Z(n24407) );
  NAND U32131 ( .A(n24409), .B(n19038), .Z(n14076) );
  NANDN U32132 ( .A(init), .B(m[276]), .Z(n19038) );
  AND U32133 ( .A(n24410), .B(n24411), .Z(n24409) );
  NAND U32134 ( .A(o[276]), .B(n23579), .Z(n24411) );
  NANDN U32135 ( .A(n23580), .B(creg[276]), .Z(n24410) );
  NAND U32136 ( .A(n24412), .B(n19036), .Z(n14075) );
  NANDN U32137 ( .A(init), .B(m[277]), .Z(n19036) );
  AND U32138 ( .A(n24413), .B(n24414), .Z(n24412) );
  NAND U32139 ( .A(o[277]), .B(n23579), .Z(n24414) );
  NANDN U32140 ( .A(n23580), .B(creg[277]), .Z(n24413) );
  NAND U32141 ( .A(n24415), .B(n19034), .Z(n14074) );
  NANDN U32142 ( .A(init), .B(m[278]), .Z(n19034) );
  AND U32143 ( .A(n24416), .B(n24417), .Z(n24415) );
  NAND U32144 ( .A(o[278]), .B(n23579), .Z(n24417) );
  NANDN U32145 ( .A(n23580), .B(creg[278]), .Z(n24416) );
  NAND U32146 ( .A(n24418), .B(n19032), .Z(n14073) );
  NANDN U32147 ( .A(init), .B(m[279]), .Z(n19032) );
  AND U32148 ( .A(n24419), .B(n24420), .Z(n24418) );
  NAND U32149 ( .A(o[279]), .B(n23579), .Z(n24420) );
  NANDN U32150 ( .A(n23580), .B(creg[279]), .Z(n24419) );
  NAND U32151 ( .A(n24421), .B(n19028), .Z(n14072) );
  NANDN U32152 ( .A(init), .B(m[280]), .Z(n19028) );
  AND U32153 ( .A(n24422), .B(n24423), .Z(n24421) );
  NAND U32154 ( .A(o[280]), .B(n23579), .Z(n24423) );
  NANDN U32155 ( .A(n23580), .B(creg[280]), .Z(n24422) );
  NAND U32156 ( .A(n24424), .B(n19026), .Z(n14071) );
  NANDN U32157 ( .A(init), .B(m[281]), .Z(n19026) );
  AND U32158 ( .A(n24425), .B(n24426), .Z(n24424) );
  NAND U32159 ( .A(o[281]), .B(n23579), .Z(n24426) );
  NANDN U32160 ( .A(n23580), .B(creg[281]), .Z(n24425) );
  NAND U32161 ( .A(n24427), .B(n19024), .Z(n14070) );
  NANDN U32162 ( .A(init), .B(m[282]), .Z(n19024) );
  AND U32163 ( .A(n24428), .B(n24429), .Z(n24427) );
  NAND U32164 ( .A(o[282]), .B(n23579), .Z(n24429) );
  NANDN U32165 ( .A(n23580), .B(creg[282]), .Z(n24428) );
  NAND U32166 ( .A(n24430), .B(n19022), .Z(n14069) );
  NANDN U32167 ( .A(init), .B(m[283]), .Z(n19022) );
  AND U32168 ( .A(n24431), .B(n24432), .Z(n24430) );
  NAND U32169 ( .A(o[283]), .B(n23579), .Z(n24432) );
  NANDN U32170 ( .A(n23580), .B(creg[283]), .Z(n24431) );
  NAND U32171 ( .A(n24433), .B(n19020), .Z(n14068) );
  NANDN U32172 ( .A(init), .B(m[284]), .Z(n19020) );
  AND U32173 ( .A(n24434), .B(n24435), .Z(n24433) );
  NAND U32174 ( .A(o[284]), .B(n23579), .Z(n24435) );
  NANDN U32175 ( .A(n23580), .B(creg[284]), .Z(n24434) );
  NAND U32176 ( .A(n24436), .B(n19018), .Z(n14067) );
  NANDN U32177 ( .A(init), .B(m[285]), .Z(n19018) );
  AND U32178 ( .A(n24437), .B(n24438), .Z(n24436) );
  NAND U32179 ( .A(o[285]), .B(n23579), .Z(n24438) );
  NANDN U32180 ( .A(n23580), .B(creg[285]), .Z(n24437) );
  NAND U32181 ( .A(n24439), .B(n19016), .Z(n14066) );
  NANDN U32182 ( .A(init), .B(m[286]), .Z(n19016) );
  AND U32183 ( .A(n24440), .B(n24441), .Z(n24439) );
  NAND U32184 ( .A(o[286]), .B(n23579), .Z(n24441) );
  NANDN U32185 ( .A(n23580), .B(creg[286]), .Z(n24440) );
  NAND U32186 ( .A(n24442), .B(n19014), .Z(n14065) );
  NANDN U32187 ( .A(init), .B(m[287]), .Z(n19014) );
  AND U32188 ( .A(n24443), .B(n24444), .Z(n24442) );
  NAND U32189 ( .A(o[287]), .B(n23579), .Z(n24444) );
  NANDN U32190 ( .A(n23580), .B(creg[287]), .Z(n24443) );
  NAND U32191 ( .A(n24445), .B(n19012), .Z(n14064) );
  NANDN U32192 ( .A(init), .B(m[288]), .Z(n19012) );
  AND U32193 ( .A(n24446), .B(n24447), .Z(n24445) );
  NAND U32194 ( .A(o[288]), .B(n23579), .Z(n24447) );
  NANDN U32195 ( .A(n23580), .B(creg[288]), .Z(n24446) );
  NAND U32196 ( .A(n24448), .B(n19010), .Z(n14063) );
  NANDN U32197 ( .A(init), .B(m[289]), .Z(n19010) );
  AND U32198 ( .A(n24449), .B(n24450), .Z(n24448) );
  NAND U32199 ( .A(o[289]), .B(n23579), .Z(n24450) );
  NANDN U32200 ( .A(n23580), .B(creg[289]), .Z(n24449) );
  NAND U32201 ( .A(n24451), .B(n19006), .Z(n14062) );
  NANDN U32202 ( .A(init), .B(m[290]), .Z(n19006) );
  AND U32203 ( .A(n24452), .B(n24453), .Z(n24451) );
  NAND U32204 ( .A(o[290]), .B(n23579), .Z(n24453) );
  NANDN U32205 ( .A(n23580), .B(creg[290]), .Z(n24452) );
  NAND U32206 ( .A(n24454), .B(n19004), .Z(n14061) );
  NANDN U32207 ( .A(init), .B(m[291]), .Z(n19004) );
  AND U32208 ( .A(n24455), .B(n24456), .Z(n24454) );
  NAND U32209 ( .A(o[291]), .B(n23579), .Z(n24456) );
  NANDN U32210 ( .A(n23580), .B(creg[291]), .Z(n24455) );
  NAND U32211 ( .A(n24457), .B(n19002), .Z(n14060) );
  NANDN U32212 ( .A(init), .B(m[292]), .Z(n19002) );
  AND U32213 ( .A(n24458), .B(n24459), .Z(n24457) );
  NAND U32214 ( .A(o[292]), .B(n23579), .Z(n24459) );
  NANDN U32215 ( .A(n23580), .B(creg[292]), .Z(n24458) );
  NAND U32216 ( .A(n24460), .B(n19000), .Z(n14059) );
  NANDN U32217 ( .A(init), .B(m[293]), .Z(n19000) );
  AND U32218 ( .A(n24461), .B(n24462), .Z(n24460) );
  NAND U32219 ( .A(o[293]), .B(n23579), .Z(n24462) );
  NANDN U32220 ( .A(n23580), .B(creg[293]), .Z(n24461) );
  NAND U32221 ( .A(n24463), .B(n18998), .Z(n14058) );
  NANDN U32222 ( .A(init), .B(m[294]), .Z(n18998) );
  AND U32223 ( .A(n24464), .B(n24465), .Z(n24463) );
  NAND U32224 ( .A(o[294]), .B(n23579), .Z(n24465) );
  NANDN U32225 ( .A(n23580), .B(creg[294]), .Z(n24464) );
  NAND U32226 ( .A(n24466), .B(n18996), .Z(n14057) );
  NANDN U32227 ( .A(init), .B(m[295]), .Z(n18996) );
  AND U32228 ( .A(n24467), .B(n24468), .Z(n24466) );
  NAND U32229 ( .A(o[295]), .B(n23579), .Z(n24468) );
  NANDN U32230 ( .A(n23580), .B(creg[295]), .Z(n24467) );
  NAND U32231 ( .A(n24469), .B(n18994), .Z(n14056) );
  NANDN U32232 ( .A(init), .B(m[296]), .Z(n18994) );
  AND U32233 ( .A(n24470), .B(n24471), .Z(n24469) );
  NAND U32234 ( .A(o[296]), .B(n23579), .Z(n24471) );
  NANDN U32235 ( .A(n23580), .B(creg[296]), .Z(n24470) );
  NAND U32236 ( .A(n24472), .B(n18992), .Z(n14055) );
  NANDN U32237 ( .A(init), .B(m[297]), .Z(n18992) );
  AND U32238 ( .A(n24473), .B(n24474), .Z(n24472) );
  NAND U32239 ( .A(o[297]), .B(n23579), .Z(n24474) );
  NANDN U32240 ( .A(n23580), .B(creg[297]), .Z(n24473) );
  NAND U32241 ( .A(n24475), .B(n18990), .Z(n14054) );
  NANDN U32242 ( .A(init), .B(m[298]), .Z(n18990) );
  AND U32243 ( .A(n24476), .B(n24477), .Z(n24475) );
  NAND U32244 ( .A(o[298]), .B(n23579), .Z(n24477) );
  NANDN U32245 ( .A(n23580), .B(creg[298]), .Z(n24476) );
  NAND U32246 ( .A(n24478), .B(n18988), .Z(n14053) );
  NANDN U32247 ( .A(init), .B(m[299]), .Z(n18988) );
  AND U32248 ( .A(n24479), .B(n24480), .Z(n24478) );
  NAND U32249 ( .A(o[299]), .B(n23579), .Z(n24480) );
  NANDN U32250 ( .A(n23580), .B(creg[299]), .Z(n24479) );
  NAND U32251 ( .A(n24481), .B(n18982), .Z(n14052) );
  NANDN U32252 ( .A(init), .B(m[300]), .Z(n18982) );
  AND U32253 ( .A(n24482), .B(n24483), .Z(n24481) );
  NAND U32254 ( .A(o[300]), .B(n23579), .Z(n24483) );
  NANDN U32255 ( .A(n23580), .B(creg[300]), .Z(n24482) );
  NAND U32256 ( .A(n24484), .B(n18980), .Z(n14051) );
  NANDN U32257 ( .A(init), .B(m[301]), .Z(n18980) );
  AND U32258 ( .A(n24485), .B(n24486), .Z(n24484) );
  NAND U32259 ( .A(o[301]), .B(n23579), .Z(n24486) );
  NANDN U32260 ( .A(n23580), .B(creg[301]), .Z(n24485) );
  NAND U32261 ( .A(n24487), .B(n18978), .Z(n14050) );
  NANDN U32262 ( .A(init), .B(m[302]), .Z(n18978) );
  AND U32263 ( .A(n24488), .B(n24489), .Z(n24487) );
  NAND U32264 ( .A(o[302]), .B(n23579), .Z(n24489) );
  NANDN U32265 ( .A(n23580), .B(creg[302]), .Z(n24488) );
  NAND U32266 ( .A(n24490), .B(n18976), .Z(n14049) );
  NANDN U32267 ( .A(init), .B(m[303]), .Z(n18976) );
  AND U32268 ( .A(n24491), .B(n24492), .Z(n24490) );
  NAND U32269 ( .A(o[303]), .B(n23579), .Z(n24492) );
  NANDN U32270 ( .A(n23580), .B(creg[303]), .Z(n24491) );
  NAND U32271 ( .A(n24493), .B(n18974), .Z(n14048) );
  NANDN U32272 ( .A(init), .B(m[304]), .Z(n18974) );
  AND U32273 ( .A(n24494), .B(n24495), .Z(n24493) );
  NAND U32274 ( .A(o[304]), .B(n23579), .Z(n24495) );
  NANDN U32275 ( .A(n23580), .B(creg[304]), .Z(n24494) );
  NAND U32276 ( .A(n24496), .B(n18972), .Z(n14047) );
  NANDN U32277 ( .A(init), .B(m[305]), .Z(n18972) );
  AND U32278 ( .A(n24497), .B(n24498), .Z(n24496) );
  NAND U32279 ( .A(o[305]), .B(n23579), .Z(n24498) );
  NANDN U32280 ( .A(n23580), .B(creg[305]), .Z(n24497) );
  NAND U32281 ( .A(n24499), .B(n18970), .Z(n14046) );
  NANDN U32282 ( .A(init), .B(m[306]), .Z(n18970) );
  AND U32283 ( .A(n24500), .B(n24501), .Z(n24499) );
  NAND U32284 ( .A(o[306]), .B(n23579), .Z(n24501) );
  NANDN U32285 ( .A(n23580), .B(creg[306]), .Z(n24500) );
  NAND U32286 ( .A(n24502), .B(n18968), .Z(n14045) );
  NANDN U32287 ( .A(init), .B(m[307]), .Z(n18968) );
  AND U32288 ( .A(n24503), .B(n24504), .Z(n24502) );
  NAND U32289 ( .A(o[307]), .B(n23579), .Z(n24504) );
  NANDN U32290 ( .A(n23580), .B(creg[307]), .Z(n24503) );
  NAND U32291 ( .A(n24505), .B(n18966), .Z(n14044) );
  NANDN U32292 ( .A(init), .B(m[308]), .Z(n18966) );
  AND U32293 ( .A(n24506), .B(n24507), .Z(n24505) );
  NAND U32294 ( .A(o[308]), .B(n23579), .Z(n24507) );
  NANDN U32295 ( .A(n23580), .B(creg[308]), .Z(n24506) );
  NAND U32296 ( .A(n24508), .B(n18964), .Z(n14043) );
  NANDN U32297 ( .A(init), .B(m[309]), .Z(n18964) );
  AND U32298 ( .A(n24509), .B(n24510), .Z(n24508) );
  NAND U32299 ( .A(o[309]), .B(n23579), .Z(n24510) );
  NANDN U32300 ( .A(n23580), .B(creg[309]), .Z(n24509) );
  NAND U32301 ( .A(n24511), .B(n18960), .Z(n14042) );
  NANDN U32302 ( .A(init), .B(m[310]), .Z(n18960) );
  AND U32303 ( .A(n24512), .B(n24513), .Z(n24511) );
  NAND U32304 ( .A(o[310]), .B(n23579), .Z(n24513) );
  NANDN U32305 ( .A(n23580), .B(creg[310]), .Z(n24512) );
  NAND U32306 ( .A(n24514), .B(n18958), .Z(n14041) );
  NANDN U32307 ( .A(init), .B(m[311]), .Z(n18958) );
  AND U32308 ( .A(n24515), .B(n24516), .Z(n24514) );
  NAND U32309 ( .A(o[311]), .B(n23579), .Z(n24516) );
  NANDN U32310 ( .A(n23580), .B(creg[311]), .Z(n24515) );
  NAND U32311 ( .A(n24517), .B(n18956), .Z(n14040) );
  NANDN U32312 ( .A(init), .B(m[312]), .Z(n18956) );
  AND U32313 ( .A(n24518), .B(n24519), .Z(n24517) );
  NAND U32314 ( .A(o[312]), .B(n23579), .Z(n24519) );
  NANDN U32315 ( .A(n23580), .B(creg[312]), .Z(n24518) );
  NAND U32316 ( .A(n24520), .B(n18954), .Z(n14039) );
  NANDN U32317 ( .A(init), .B(m[313]), .Z(n18954) );
  AND U32318 ( .A(n24521), .B(n24522), .Z(n24520) );
  NAND U32319 ( .A(o[313]), .B(n23579), .Z(n24522) );
  NANDN U32320 ( .A(n23580), .B(creg[313]), .Z(n24521) );
  NAND U32321 ( .A(n24523), .B(n18952), .Z(n14038) );
  NANDN U32322 ( .A(init), .B(m[314]), .Z(n18952) );
  AND U32323 ( .A(n24524), .B(n24525), .Z(n24523) );
  NAND U32324 ( .A(o[314]), .B(n23579), .Z(n24525) );
  NANDN U32325 ( .A(n23580), .B(creg[314]), .Z(n24524) );
  NAND U32326 ( .A(n24526), .B(n18950), .Z(n14037) );
  NANDN U32327 ( .A(init), .B(m[315]), .Z(n18950) );
  AND U32328 ( .A(n24527), .B(n24528), .Z(n24526) );
  NAND U32329 ( .A(o[315]), .B(n23579), .Z(n24528) );
  NANDN U32330 ( .A(n23580), .B(creg[315]), .Z(n24527) );
  NAND U32331 ( .A(n24529), .B(n18948), .Z(n14036) );
  NANDN U32332 ( .A(init), .B(m[316]), .Z(n18948) );
  AND U32333 ( .A(n24530), .B(n24531), .Z(n24529) );
  NAND U32334 ( .A(o[316]), .B(n23579), .Z(n24531) );
  NANDN U32335 ( .A(n23580), .B(creg[316]), .Z(n24530) );
  NAND U32336 ( .A(n24532), .B(n18946), .Z(n14035) );
  NANDN U32337 ( .A(init), .B(m[317]), .Z(n18946) );
  AND U32338 ( .A(n24533), .B(n24534), .Z(n24532) );
  NAND U32339 ( .A(o[317]), .B(n23579), .Z(n24534) );
  NANDN U32340 ( .A(n23580), .B(creg[317]), .Z(n24533) );
  NAND U32341 ( .A(n24535), .B(n18944), .Z(n14034) );
  NANDN U32342 ( .A(init), .B(m[318]), .Z(n18944) );
  AND U32343 ( .A(n24536), .B(n24537), .Z(n24535) );
  NAND U32344 ( .A(o[318]), .B(n23579), .Z(n24537) );
  NANDN U32345 ( .A(n23580), .B(creg[318]), .Z(n24536) );
  NAND U32346 ( .A(n24538), .B(n18942), .Z(n14033) );
  NANDN U32347 ( .A(init), .B(m[319]), .Z(n18942) );
  AND U32348 ( .A(n24539), .B(n24540), .Z(n24538) );
  NAND U32349 ( .A(o[319]), .B(n23579), .Z(n24540) );
  NANDN U32350 ( .A(n23580), .B(creg[319]), .Z(n24539) );
  NAND U32351 ( .A(n24541), .B(n18938), .Z(n14032) );
  NANDN U32352 ( .A(init), .B(m[320]), .Z(n18938) );
  AND U32353 ( .A(n24542), .B(n24543), .Z(n24541) );
  NAND U32354 ( .A(o[320]), .B(n23579), .Z(n24543) );
  NANDN U32355 ( .A(n23580), .B(creg[320]), .Z(n24542) );
  NAND U32356 ( .A(n24544), .B(n18936), .Z(n14031) );
  NANDN U32357 ( .A(init), .B(m[321]), .Z(n18936) );
  AND U32358 ( .A(n24545), .B(n24546), .Z(n24544) );
  NAND U32359 ( .A(o[321]), .B(n23579), .Z(n24546) );
  NANDN U32360 ( .A(n23580), .B(creg[321]), .Z(n24545) );
  NAND U32361 ( .A(n24547), .B(n18934), .Z(n14030) );
  NANDN U32362 ( .A(init), .B(m[322]), .Z(n18934) );
  AND U32363 ( .A(n24548), .B(n24549), .Z(n24547) );
  NAND U32364 ( .A(o[322]), .B(n23579), .Z(n24549) );
  NANDN U32365 ( .A(n23580), .B(creg[322]), .Z(n24548) );
  NAND U32366 ( .A(n24550), .B(n18932), .Z(n14029) );
  NANDN U32367 ( .A(init), .B(m[323]), .Z(n18932) );
  AND U32368 ( .A(n24551), .B(n24552), .Z(n24550) );
  NAND U32369 ( .A(o[323]), .B(n23579), .Z(n24552) );
  NANDN U32370 ( .A(n23580), .B(creg[323]), .Z(n24551) );
  NAND U32371 ( .A(n24553), .B(n18930), .Z(n14028) );
  NANDN U32372 ( .A(init), .B(m[324]), .Z(n18930) );
  AND U32373 ( .A(n24554), .B(n24555), .Z(n24553) );
  NAND U32374 ( .A(o[324]), .B(n23579), .Z(n24555) );
  NANDN U32375 ( .A(n23580), .B(creg[324]), .Z(n24554) );
  NAND U32376 ( .A(n24556), .B(n18928), .Z(n14027) );
  NANDN U32377 ( .A(init), .B(m[325]), .Z(n18928) );
  AND U32378 ( .A(n24557), .B(n24558), .Z(n24556) );
  NAND U32379 ( .A(o[325]), .B(n23579), .Z(n24558) );
  NANDN U32380 ( .A(n23580), .B(creg[325]), .Z(n24557) );
  NAND U32381 ( .A(n24559), .B(n18926), .Z(n14026) );
  NANDN U32382 ( .A(init), .B(m[326]), .Z(n18926) );
  AND U32383 ( .A(n24560), .B(n24561), .Z(n24559) );
  NAND U32384 ( .A(o[326]), .B(n23579), .Z(n24561) );
  NANDN U32385 ( .A(n23580), .B(creg[326]), .Z(n24560) );
  NAND U32386 ( .A(n24562), .B(n18924), .Z(n14025) );
  NANDN U32387 ( .A(init), .B(m[327]), .Z(n18924) );
  AND U32388 ( .A(n24563), .B(n24564), .Z(n24562) );
  NAND U32389 ( .A(o[327]), .B(n23579), .Z(n24564) );
  NANDN U32390 ( .A(n23580), .B(creg[327]), .Z(n24563) );
  NAND U32391 ( .A(n24565), .B(n18922), .Z(n14024) );
  NANDN U32392 ( .A(init), .B(m[328]), .Z(n18922) );
  AND U32393 ( .A(n24566), .B(n24567), .Z(n24565) );
  NAND U32394 ( .A(o[328]), .B(n23579), .Z(n24567) );
  NANDN U32395 ( .A(n23580), .B(creg[328]), .Z(n24566) );
  NAND U32396 ( .A(n24568), .B(n18920), .Z(n14023) );
  NANDN U32397 ( .A(init), .B(m[329]), .Z(n18920) );
  AND U32398 ( .A(n24569), .B(n24570), .Z(n24568) );
  NAND U32399 ( .A(o[329]), .B(n23579), .Z(n24570) );
  NANDN U32400 ( .A(n23580), .B(creg[329]), .Z(n24569) );
  NAND U32401 ( .A(n24571), .B(n18916), .Z(n14022) );
  NANDN U32402 ( .A(init), .B(m[330]), .Z(n18916) );
  AND U32403 ( .A(n24572), .B(n24573), .Z(n24571) );
  NAND U32404 ( .A(o[330]), .B(n23579), .Z(n24573) );
  NANDN U32405 ( .A(n23580), .B(creg[330]), .Z(n24572) );
  NAND U32406 ( .A(n24574), .B(n18914), .Z(n14021) );
  NANDN U32407 ( .A(init), .B(m[331]), .Z(n18914) );
  AND U32408 ( .A(n24575), .B(n24576), .Z(n24574) );
  NAND U32409 ( .A(o[331]), .B(n23579), .Z(n24576) );
  NANDN U32410 ( .A(n23580), .B(creg[331]), .Z(n24575) );
  NAND U32411 ( .A(n24577), .B(n18912), .Z(n14020) );
  NANDN U32412 ( .A(init), .B(m[332]), .Z(n18912) );
  AND U32413 ( .A(n24578), .B(n24579), .Z(n24577) );
  NAND U32414 ( .A(o[332]), .B(n23579), .Z(n24579) );
  NANDN U32415 ( .A(n23580), .B(creg[332]), .Z(n24578) );
  NAND U32416 ( .A(n24580), .B(n18910), .Z(n14019) );
  NANDN U32417 ( .A(init), .B(m[333]), .Z(n18910) );
  AND U32418 ( .A(n24581), .B(n24582), .Z(n24580) );
  NAND U32419 ( .A(o[333]), .B(n23579), .Z(n24582) );
  NANDN U32420 ( .A(n23580), .B(creg[333]), .Z(n24581) );
  NAND U32421 ( .A(n24583), .B(n18908), .Z(n14018) );
  NANDN U32422 ( .A(init), .B(m[334]), .Z(n18908) );
  AND U32423 ( .A(n24584), .B(n24585), .Z(n24583) );
  NAND U32424 ( .A(o[334]), .B(n23579), .Z(n24585) );
  NANDN U32425 ( .A(n23580), .B(creg[334]), .Z(n24584) );
  NAND U32426 ( .A(n24586), .B(n18906), .Z(n14017) );
  NANDN U32427 ( .A(init), .B(m[335]), .Z(n18906) );
  AND U32428 ( .A(n24587), .B(n24588), .Z(n24586) );
  NAND U32429 ( .A(o[335]), .B(n23579), .Z(n24588) );
  NANDN U32430 ( .A(n23580), .B(creg[335]), .Z(n24587) );
  NAND U32431 ( .A(n24589), .B(n18904), .Z(n14016) );
  NANDN U32432 ( .A(init), .B(m[336]), .Z(n18904) );
  AND U32433 ( .A(n24590), .B(n24591), .Z(n24589) );
  NAND U32434 ( .A(o[336]), .B(n23579), .Z(n24591) );
  NANDN U32435 ( .A(n23580), .B(creg[336]), .Z(n24590) );
  NAND U32436 ( .A(n24592), .B(n18902), .Z(n14015) );
  NANDN U32437 ( .A(init), .B(m[337]), .Z(n18902) );
  AND U32438 ( .A(n24593), .B(n24594), .Z(n24592) );
  NAND U32439 ( .A(o[337]), .B(n23579), .Z(n24594) );
  NANDN U32440 ( .A(n23580), .B(creg[337]), .Z(n24593) );
  NAND U32441 ( .A(n24595), .B(n18900), .Z(n14014) );
  NANDN U32442 ( .A(init), .B(m[338]), .Z(n18900) );
  AND U32443 ( .A(n24596), .B(n24597), .Z(n24595) );
  NAND U32444 ( .A(o[338]), .B(n23579), .Z(n24597) );
  NANDN U32445 ( .A(n23580), .B(creg[338]), .Z(n24596) );
  NAND U32446 ( .A(n24598), .B(n18898), .Z(n14013) );
  NANDN U32447 ( .A(init), .B(m[339]), .Z(n18898) );
  AND U32448 ( .A(n24599), .B(n24600), .Z(n24598) );
  NAND U32449 ( .A(o[339]), .B(n23579), .Z(n24600) );
  NANDN U32450 ( .A(n23580), .B(creg[339]), .Z(n24599) );
  NAND U32451 ( .A(n24601), .B(n18894), .Z(n14012) );
  NANDN U32452 ( .A(init), .B(m[340]), .Z(n18894) );
  AND U32453 ( .A(n24602), .B(n24603), .Z(n24601) );
  NAND U32454 ( .A(o[340]), .B(n23579), .Z(n24603) );
  NANDN U32455 ( .A(n23580), .B(creg[340]), .Z(n24602) );
  NAND U32456 ( .A(n24604), .B(n18892), .Z(n14011) );
  NANDN U32457 ( .A(init), .B(m[341]), .Z(n18892) );
  AND U32458 ( .A(n24605), .B(n24606), .Z(n24604) );
  NAND U32459 ( .A(o[341]), .B(n23579), .Z(n24606) );
  NANDN U32460 ( .A(n23580), .B(creg[341]), .Z(n24605) );
  NAND U32461 ( .A(n24607), .B(n18890), .Z(n14010) );
  NANDN U32462 ( .A(init), .B(m[342]), .Z(n18890) );
  AND U32463 ( .A(n24608), .B(n24609), .Z(n24607) );
  NAND U32464 ( .A(o[342]), .B(n23579), .Z(n24609) );
  NANDN U32465 ( .A(n23580), .B(creg[342]), .Z(n24608) );
  NAND U32466 ( .A(n24610), .B(n18888), .Z(n14009) );
  NANDN U32467 ( .A(init), .B(m[343]), .Z(n18888) );
  AND U32468 ( .A(n24611), .B(n24612), .Z(n24610) );
  NAND U32469 ( .A(o[343]), .B(n23579), .Z(n24612) );
  NANDN U32470 ( .A(n23580), .B(creg[343]), .Z(n24611) );
  NAND U32471 ( .A(n24613), .B(n18886), .Z(n14008) );
  NANDN U32472 ( .A(init), .B(m[344]), .Z(n18886) );
  AND U32473 ( .A(n24614), .B(n24615), .Z(n24613) );
  NAND U32474 ( .A(o[344]), .B(n23579), .Z(n24615) );
  NANDN U32475 ( .A(n23580), .B(creg[344]), .Z(n24614) );
  NAND U32476 ( .A(n24616), .B(n18884), .Z(n14007) );
  NANDN U32477 ( .A(init), .B(m[345]), .Z(n18884) );
  AND U32478 ( .A(n24617), .B(n24618), .Z(n24616) );
  NAND U32479 ( .A(o[345]), .B(n23579), .Z(n24618) );
  NANDN U32480 ( .A(n23580), .B(creg[345]), .Z(n24617) );
  NAND U32481 ( .A(n24619), .B(n18882), .Z(n14006) );
  NANDN U32482 ( .A(init), .B(m[346]), .Z(n18882) );
  AND U32483 ( .A(n24620), .B(n24621), .Z(n24619) );
  NAND U32484 ( .A(o[346]), .B(n23579), .Z(n24621) );
  NANDN U32485 ( .A(n23580), .B(creg[346]), .Z(n24620) );
  NAND U32486 ( .A(n24622), .B(n18880), .Z(n14005) );
  NANDN U32487 ( .A(init), .B(m[347]), .Z(n18880) );
  AND U32488 ( .A(n24623), .B(n24624), .Z(n24622) );
  NAND U32489 ( .A(o[347]), .B(n23579), .Z(n24624) );
  NANDN U32490 ( .A(n23580), .B(creg[347]), .Z(n24623) );
  NAND U32491 ( .A(n24625), .B(n18878), .Z(n14004) );
  NANDN U32492 ( .A(init), .B(m[348]), .Z(n18878) );
  AND U32493 ( .A(n24626), .B(n24627), .Z(n24625) );
  NAND U32494 ( .A(o[348]), .B(n23579), .Z(n24627) );
  NANDN U32495 ( .A(n23580), .B(creg[348]), .Z(n24626) );
  NAND U32496 ( .A(n24628), .B(n18876), .Z(n14003) );
  NANDN U32497 ( .A(init), .B(m[349]), .Z(n18876) );
  AND U32498 ( .A(n24629), .B(n24630), .Z(n24628) );
  NAND U32499 ( .A(o[349]), .B(n23579), .Z(n24630) );
  NANDN U32500 ( .A(n23580), .B(creg[349]), .Z(n24629) );
  NAND U32501 ( .A(n24631), .B(n18872), .Z(n14002) );
  NANDN U32502 ( .A(init), .B(m[350]), .Z(n18872) );
  AND U32503 ( .A(n24632), .B(n24633), .Z(n24631) );
  NAND U32504 ( .A(o[350]), .B(n23579), .Z(n24633) );
  NANDN U32505 ( .A(n23580), .B(creg[350]), .Z(n24632) );
  NAND U32506 ( .A(n24634), .B(n18870), .Z(n14001) );
  NANDN U32507 ( .A(init), .B(m[351]), .Z(n18870) );
  AND U32508 ( .A(n24635), .B(n24636), .Z(n24634) );
  NAND U32509 ( .A(o[351]), .B(n23579), .Z(n24636) );
  NANDN U32510 ( .A(n23580), .B(creg[351]), .Z(n24635) );
  NAND U32511 ( .A(n24637), .B(n18868), .Z(n14000) );
  NANDN U32512 ( .A(init), .B(m[352]), .Z(n18868) );
  AND U32513 ( .A(n24638), .B(n24639), .Z(n24637) );
  NAND U32514 ( .A(o[352]), .B(n23579), .Z(n24639) );
  NANDN U32515 ( .A(n23580), .B(creg[352]), .Z(n24638) );
  NAND U32516 ( .A(n24640), .B(n18866), .Z(n13999) );
  NANDN U32517 ( .A(init), .B(m[353]), .Z(n18866) );
  AND U32518 ( .A(n24641), .B(n24642), .Z(n24640) );
  NAND U32519 ( .A(o[353]), .B(n23579), .Z(n24642) );
  NANDN U32520 ( .A(n23580), .B(creg[353]), .Z(n24641) );
  NAND U32521 ( .A(n24643), .B(n18864), .Z(n13998) );
  NANDN U32522 ( .A(init), .B(m[354]), .Z(n18864) );
  AND U32523 ( .A(n24644), .B(n24645), .Z(n24643) );
  NAND U32524 ( .A(o[354]), .B(n23579), .Z(n24645) );
  NANDN U32525 ( .A(n23580), .B(creg[354]), .Z(n24644) );
  NAND U32526 ( .A(n24646), .B(n18862), .Z(n13997) );
  NANDN U32527 ( .A(init), .B(m[355]), .Z(n18862) );
  AND U32528 ( .A(n24647), .B(n24648), .Z(n24646) );
  NAND U32529 ( .A(o[355]), .B(n23579), .Z(n24648) );
  NANDN U32530 ( .A(n23580), .B(creg[355]), .Z(n24647) );
  NAND U32531 ( .A(n24649), .B(n18860), .Z(n13996) );
  NANDN U32532 ( .A(init), .B(m[356]), .Z(n18860) );
  AND U32533 ( .A(n24650), .B(n24651), .Z(n24649) );
  NAND U32534 ( .A(o[356]), .B(n23579), .Z(n24651) );
  NANDN U32535 ( .A(n23580), .B(creg[356]), .Z(n24650) );
  NAND U32536 ( .A(n24652), .B(n18858), .Z(n13995) );
  NANDN U32537 ( .A(init), .B(m[357]), .Z(n18858) );
  AND U32538 ( .A(n24653), .B(n24654), .Z(n24652) );
  NAND U32539 ( .A(o[357]), .B(n23579), .Z(n24654) );
  NANDN U32540 ( .A(n23580), .B(creg[357]), .Z(n24653) );
  NAND U32541 ( .A(n24655), .B(n18856), .Z(n13994) );
  NANDN U32542 ( .A(init), .B(m[358]), .Z(n18856) );
  AND U32543 ( .A(n24656), .B(n24657), .Z(n24655) );
  NAND U32544 ( .A(o[358]), .B(n23579), .Z(n24657) );
  NANDN U32545 ( .A(n23580), .B(creg[358]), .Z(n24656) );
  NAND U32546 ( .A(n24658), .B(n18854), .Z(n13993) );
  NANDN U32547 ( .A(init), .B(m[359]), .Z(n18854) );
  AND U32548 ( .A(n24659), .B(n24660), .Z(n24658) );
  NAND U32549 ( .A(o[359]), .B(n23579), .Z(n24660) );
  NANDN U32550 ( .A(n23580), .B(creg[359]), .Z(n24659) );
  NAND U32551 ( .A(n24661), .B(n18850), .Z(n13992) );
  NANDN U32552 ( .A(init), .B(m[360]), .Z(n18850) );
  AND U32553 ( .A(n24662), .B(n24663), .Z(n24661) );
  NAND U32554 ( .A(o[360]), .B(n23579), .Z(n24663) );
  NANDN U32555 ( .A(n23580), .B(creg[360]), .Z(n24662) );
  NAND U32556 ( .A(n24664), .B(n18848), .Z(n13991) );
  NANDN U32557 ( .A(init), .B(m[361]), .Z(n18848) );
  AND U32558 ( .A(n24665), .B(n24666), .Z(n24664) );
  NAND U32559 ( .A(o[361]), .B(n23579), .Z(n24666) );
  NANDN U32560 ( .A(n23580), .B(creg[361]), .Z(n24665) );
  NAND U32561 ( .A(n24667), .B(n18846), .Z(n13990) );
  NANDN U32562 ( .A(init), .B(m[362]), .Z(n18846) );
  AND U32563 ( .A(n24668), .B(n24669), .Z(n24667) );
  NAND U32564 ( .A(o[362]), .B(n23579), .Z(n24669) );
  NANDN U32565 ( .A(n23580), .B(creg[362]), .Z(n24668) );
  NAND U32566 ( .A(n24670), .B(n18844), .Z(n13989) );
  NANDN U32567 ( .A(init), .B(m[363]), .Z(n18844) );
  AND U32568 ( .A(n24671), .B(n24672), .Z(n24670) );
  NAND U32569 ( .A(o[363]), .B(n23579), .Z(n24672) );
  NANDN U32570 ( .A(n23580), .B(creg[363]), .Z(n24671) );
  NAND U32571 ( .A(n24673), .B(n18842), .Z(n13988) );
  NANDN U32572 ( .A(init), .B(m[364]), .Z(n18842) );
  AND U32573 ( .A(n24674), .B(n24675), .Z(n24673) );
  NAND U32574 ( .A(o[364]), .B(n23579), .Z(n24675) );
  NANDN U32575 ( .A(n23580), .B(creg[364]), .Z(n24674) );
  NAND U32576 ( .A(n24676), .B(n18840), .Z(n13987) );
  NANDN U32577 ( .A(init), .B(m[365]), .Z(n18840) );
  AND U32578 ( .A(n24677), .B(n24678), .Z(n24676) );
  NAND U32579 ( .A(o[365]), .B(n23579), .Z(n24678) );
  NANDN U32580 ( .A(n23580), .B(creg[365]), .Z(n24677) );
  NAND U32581 ( .A(n24679), .B(n18838), .Z(n13986) );
  NANDN U32582 ( .A(init), .B(m[366]), .Z(n18838) );
  AND U32583 ( .A(n24680), .B(n24681), .Z(n24679) );
  NAND U32584 ( .A(o[366]), .B(n23579), .Z(n24681) );
  NANDN U32585 ( .A(n23580), .B(creg[366]), .Z(n24680) );
  NAND U32586 ( .A(n24682), .B(n18836), .Z(n13985) );
  NANDN U32587 ( .A(init), .B(m[367]), .Z(n18836) );
  AND U32588 ( .A(n24683), .B(n24684), .Z(n24682) );
  NAND U32589 ( .A(o[367]), .B(n23579), .Z(n24684) );
  NANDN U32590 ( .A(n23580), .B(creg[367]), .Z(n24683) );
  NAND U32591 ( .A(n24685), .B(n18834), .Z(n13984) );
  NANDN U32592 ( .A(init), .B(m[368]), .Z(n18834) );
  AND U32593 ( .A(n24686), .B(n24687), .Z(n24685) );
  NAND U32594 ( .A(o[368]), .B(n23579), .Z(n24687) );
  NANDN U32595 ( .A(n23580), .B(creg[368]), .Z(n24686) );
  NAND U32596 ( .A(n24688), .B(n18832), .Z(n13983) );
  NANDN U32597 ( .A(init), .B(m[369]), .Z(n18832) );
  AND U32598 ( .A(n24689), .B(n24690), .Z(n24688) );
  NAND U32599 ( .A(o[369]), .B(n23579), .Z(n24690) );
  NANDN U32600 ( .A(n23580), .B(creg[369]), .Z(n24689) );
  NAND U32601 ( .A(n24691), .B(n18828), .Z(n13982) );
  NANDN U32602 ( .A(init), .B(m[370]), .Z(n18828) );
  AND U32603 ( .A(n24692), .B(n24693), .Z(n24691) );
  NAND U32604 ( .A(o[370]), .B(n23579), .Z(n24693) );
  NANDN U32605 ( .A(n23580), .B(creg[370]), .Z(n24692) );
  NAND U32606 ( .A(n24694), .B(n18826), .Z(n13981) );
  NANDN U32607 ( .A(init), .B(m[371]), .Z(n18826) );
  AND U32608 ( .A(n24695), .B(n24696), .Z(n24694) );
  NAND U32609 ( .A(o[371]), .B(n23579), .Z(n24696) );
  NANDN U32610 ( .A(n23580), .B(creg[371]), .Z(n24695) );
  NAND U32611 ( .A(n24697), .B(n18824), .Z(n13980) );
  NANDN U32612 ( .A(init), .B(m[372]), .Z(n18824) );
  AND U32613 ( .A(n24698), .B(n24699), .Z(n24697) );
  NAND U32614 ( .A(o[372]), .B(n23579), .Z(n24699) );
  NANDN U32615 ( .A(n23580), .B(creg[372]), .Z(n24698) );
  NAND U32616 ( .A(n24700), .B(n18822), .Z(n13979) );
  NANDN U32617 ( .A(init), .B(m[373]), .Z(n18822) );
  AND U32618 ( .A(n24701), .B(n24702), .Z(n24700) );
  NAND U32619 ( .A(o[373]), .B(n23579), .Z(n24702) );
  NANDN U32620 ( .A(n23580), .B(creg[373]), .Z(n24701) );
  NAND U32621 ( .A(n24703), .B(n18820), .Z(n13978) );
  NANDN U32622 ( .A(init), .B(m[374]), .Z(n18820) );
  AND U32623 ( .A(n24704), .B(n24705), .Z(n24703) );
  NAND U32624 ( .A(o[374]), .B(n23579), .Z(n24705) );
  NANDN U32625 ( .A(n23580), .B(creg[374]), .Z(n24704) );
  NAND U32626 ( .A(n24706), .B(n18818), .Z(n13977) );
  NANDN U32627 ( .A(init), .B(m[375]), .Z(n18818) );
  AND U32628 ( .A(n24707), .B(n24708), .Z(n24706) );
  NAND U32629 ( .A(o[375]), .B(n23579), .Z(n24708) );
  NANDN U32630 ( .A(n23580), .B(creg[375]), .Z(n24707) );
  NAND U32631 ( .A(n24709), .B(n18816), .Z(n13976) );
  NANDN U32632 ( .A(init), .B(m[376]), .Z(n18816) );
  AND U32633 ( .A(n24710), .B(n24711), .Z(n24709) );
  NAND U32634 ( .A(o[376]), .B(n23579), .Z(n24711) );
  NANDN U32635 ( .A(n23580), .B(creg[376]), .Z(n24710) );
  NAND U32636 ( .A(n24712), .B(n18814), .Z(n13975) );
  NANDN U32637 ( .A(init), .B(m[377]), .Z(n18814) );
  AND U32638 ( .A(n24713), .B(n24714), .Z(n24712) );
  NAND U32639 ( .A(o[377]), .B(n23579), .Z(n24714) );
  NANDN U32640 ( .A(n23580), .B(creg[377]), .Z(n24713) );
  NAND U32641 ( .A(n24715), .B(n18812), .Z(n13974) );
  NANDN U32642 ( .A(init), .B(m[378]), .Z(n18812) );
  AND U32643 ( .A(n24716), .B(n24717), .Z(n24715) );
  NAND U32644 ( .A(o[378]), .B(n23579), .Z(n24717) );
  NANDN U32645 ( .A(n23580), .B(creg[378]), .Z(n24716) );
  NAND U32646 ( .A(n24718), .B(n18810), .Z(n13973) );
  NANDN U32647 ( .A(init), .B(m[379]), .Z(n18810) );
  AND U32648 ( .A(n24719), .B(n24720), .Z(n24718) );
  NAND U32649 ( .A(o[379]), .B(n23579), .Z(n24720) );
  NANDN U32650 ( .A(n23580), .B(creg[379]), .Z(n24719) );
  NAND U32651 ( .A(n24721), .B(n18806), .Z(n13972) );
  NANDN U32652 ( .A(init), .B(m[380]), .Z(n18806) );
  AND U32653 ( .A(n24722), .B(n24723), .Z(n24721) );
  NAND U32654 ( .A(o[380]), .B(n23579), .Z(n24723) );
  NANDN U32655 ( .A(n23580), .B(creg[380]), .Z(n24722) );
  NAND U32656 ( .A(n24724), .B(n18804), .Z(n13971) );
  NANDN U32657 ( .A(init), .B(m[381]), .Z(n18804) );
  AND U32658 ( .A(n24725), .B(n24726), .Z(n24724) );
  NAND U32659 ( .A(o[381]), .B(n23579), .Z(n24726) );
  NANDN U32660 ( .A(n23580), .B(creg[381]), .Z(n24725) );
  NAND U32661 ( .A(n24727), .B(n18802), .Z(n13970) );
  NANDN U32662 ( .A(init), .B(m[382]), .Z(n18802) );
  AND U32663 ( .A(n24728), .B(n24729), .Z(n24727) );
  NAND U32664 ( .A(o[382]), .B(n23579), .Z(n24729) );
  NANDN U32665 ( .A(n23580), .B(creg[382]), .Z(n24728) );
  NAND U32666 ( .A(n24730), .B(n18800), .Z(n13969) );
  NANDN U32667 ( .A(init), .B(m[383]), .Z(n18800) );
  AND U32668 ( .A(n24731), .B(n24732), .Z(n24730) );
  NAND U32669 ( .A(o[383]), .B(n23579), .Z(n24732) );
  NANDN U32670 ( .A(n23580), .B(creg[383]), .Z(n24731) );
  NAND U32671 ( .A(n24733), .B(n18798), .Z(n13968) );
  NANDN U32672 ( .A(init), .B(m[384]), .Z(n18798) );
  AND U32673 ( .A(n24734), .B(n24735), .Z(n24733) );
  NAND U32674 ( .A(o[384]), .B(n23579), .Z(n24735) );
  NANDN U32675 ( .A(n23580), .B(creg[384]), .Z(n24734) );
  NAND U32676 ( .A(n24736), .B(n18796), .Z(n13967) );
  NANDN U32677 ( .A(init), .B(m[385]), .Z(n18796) );
  AND U32678 ( .A(n24737), .B(n24738), .Z(n24736) );
  NAND U32679 ( .A(o[385]), .B(n23579), .Z(n24738) );
  NANDN U32680 ( .A(n23580), .B(creg[385]), .Z(n24737) );
  NAND U32681 ( .A(n24739), .B(n18794), .Z(n13966) );
  NANDN U32682 ( .A(init), .B(m[386]), .Z(n18794) );
  AND U32683 ( .A(n24740), .B(n24741), .Z(n24739) );
  NAND U32684 ( .A(o[386]), .B(n23579), .Z(n24741) );
  NANDN U32685 ( .A(n23580), .B(creg[386]), .Z(n24740) );
  NAND U32686 ( .A(n24742), .B(n18792), .Z(n13965) );
  NANDN U32687 ( .A(init), .B(m[387]), .Z(n18792) );
  AND U32688 ( .A(n24743), .B(n24744), .Z(n24742) );
  NAND U32689 ( .A(o[387]), .B(n23579), .Z(n24744) );
  NANDN U32690 ( .A(n23580), .B(creg[387]), .Z(n24743) );
  NAND U32691 ( .A(n24745), .B(n18790), .Z(n13964) );
  NANDN U32692 ( .A(init), .B(m[388]), .Z(n18790) );
  AND U32693 ( .A(n24746), .B(n24747), .Z(n24745) );
  NAND U32694 ( .A(o[388]), .B(n23579), .Z(n24747) );
  NANDN U32695 ( .A(n23580), .B(creg[388]), .Z(n24746) );
  NAND U32696 ( .A(n24748), .B(n18788), .Z(n13963) );
  NANDN U32697 ( .A(init), .B(m[389]), .Z(n18788) );
  AND U32698 ( .A(n24749), .B(n24750), .Z(n24748) );
  NAND U32699 ( .A(o[389]), .B(n23579), .Z(n24750) );
  NANDN U32700 ( .A(n23580), .B(creg[389]), .Z(n24749) );
  NAND U32701 ( .A(n24751), .B(n18784), .Z(n13962) );
  NANDN U32702 ( .A(init), .B(m[390]), .Z(n18784) );
  AND U32703 ( .A(n24752), .B(n24753), .Z(n24751) );
  NAND U32704 ( .A(o[390]), .B(n23579), .Z(n24753) );
  NANDN U32705 ( .A(n23580), .B(creg[390]), .Z(n24752) );
  NAND U32706 ( .A(n24754), .B(n18782), .Z(n13961) );
  NANDN U32707 ( .A(init), .B(m[391]), .Z(n18782) );
  AND U32708 ( .A(n24755), .B(n24756), .Z(n24754) );
  NAND U32709 ( .A(o[391]), .B(n23579), .Z(n24756) );
  NANDN U32710 ( .A(n23580), .B(creg[391]), .Z(n24755) );
  NAND U32711 ( .A(n24757), .B(n18780), .Z(n13960) );
  NANDN U32712 ( .A(init), .B(m[392]), .Z(n18780) );
  AND U32713 ( .A(n24758), .B(n24759), .Z(n24757) );
  NAND U32714 ( .A(o[392]), .B(n23579), .Z(n24759) );
  NANDN U32715 ( .A(n23580), .B(creg[392]), .Z(n24758) );
  NAND U32716 ( .A(n24760), .B(n18778), .Z(n13959) );
  NANDN U32717 ( .A(init), .B(m[393]), .Z(n18778) );
  AND U32718 ( .A(n24761), .B(n24762), .Z(n24760) );
  NAND U32719 ( .A(o[393]), .B(n23579), .Z(n24762) );
  NANDN U32720 ( .A(n23580), .B(creg[393]), .Z(n24761) );
  NAND U32721 ( .A(n24763), .B(n18776), .Z(n13958) );
  NANDN U32722 ( .A(init), .B(m[394]), .Z(n18776) );
  AND U32723 ( .A(n24764), .B(n24765), .Z(n24763) );
  NAND U32724 ( .A(o[394]), .B(n23579), .Z(n24765) );
  NANDN U32725 ( .A(n23580), .B(creg[394]), .Z(n24764) );
  NAND U32726 ( .A(n24766), .B(n18774), .Z(n13957) );
  NANDN U32727 ( .A(init), .B(m[395]), .Z(n18774) );
  AND U32728 ( .A(n24767), .B(n24768), .Z(n24766) );
  NAND U32729 ( .A(o[395]), .B(n23579), .Z(n24768) );
  NANDN U32730 ( .A(n23580), .B(creg[395]), .Z(n24767) );
  NAND U32731 ( .A(n24769), .B(n18772), .Z(n13956) );
  NANDN U32732 ( .A(init), .B(m[396]), .Z(n18772) );
  AND U32733 ( .A(n24770), .B(n24771), .Z(n24769) );
  NAND U32734 ( .A(o[396]), .B(n23579), .Z(n24771) );
  NANDN U32735 ( .A(n23580), .B(creg[396]), .Z(n24770) );
  NAND U32736 ( .A(n24772), .B(n18770), .Z(n13955) );
  NANDN U32737 ( .A(init), .B(m[397]), .Z(n18770) );
  AND U32738 ( .A(n24773), .B(n24774), .Z(n24772) );
  NAND U32739 ( .A(o[397]), .B(n23579), .Z(n24774) );
  NANDN U32740 ( .A(n23580), .B(creg[397]), .Z(n24773) );
  NAND U32741 ( .A(n24775), .B(n18768), .Z(n13954) );
  NANDN U32742 ( .A(init), .B(m[398]), .Z(n18768) );
  AND U32743 ( .A(n24776), .B(n24777), .Z(n24775) );
  NAND U32744 ( .A(o[398]), .B(n23579), .Z(n24777) );
  NANDN U32745 ( .A(n23580), .B(creg[398]), .Z(n24776) );
  NAND U32746 ( .A(n24778), .B(n18766), .Z(n13953) );
  NANDN U32747 ( .A(init), .B(m[399]), .Z(n18766) );
  AND U32748 ( .A(n24779), .B(n24780), .Z(n24778) );
  NAND U32749 ( .A(o[399]), .B(n23579), .Z(n24780) );
  NANDN U32750 ( .A(n23580), .B(creg[399]), .Z(n24779) );
  NAND U32751 ( .A(n24781), .B(n18760), .Z(n13952) );
  NANDN U32752 ( .A(init), .B(m[400]), .Z(n18760) );
  AND U32753 ( .A(n24782), .B(n24783), .Z(n24781) );
  NAND U32754 ( .A(o[400]), .B(n23579), .Z(n24783) );
  NANDN U32755 ( .A(n23580), .B(creg[400]), .Z(n24782) );
  NAND U32756 ( .A(n24784), .B(n18758), .Z(n13951) );
  NANDN U32757 ( .A(init), .B(m[401]), .Z(n18758) );
  AND U32758 ( .A(n24785), .B(n24786), .Z(n24784) );
  NAND U32759 ( .A(o[401]), .B(n23579), .Z(n24786) );
  NANDN U32760 ( .A(n23580), .B(creg[401]), .Z(n24785) );
  NAND U32761 ( .A(n24787), .B(n18756), .Z(n13950) );
  NANDN U32762 ( .A(init), .B(m[402]), .Z(n18756) );
  AND U32763 ( .A(n24788), .B(n24789), .Z(n24787) );
  NAND U32764 ( .A(o[402]), .B(n23579), .Z(n24789) );
  NANDN U32765 ( .A(n23580), .B(creg[402]), .Z(n24788) );
  NAND U32766 ( .A(n24790), .B(n18754), .Z(n13949) );
  NANDN U32767 ( .A(init), .B(m[403]), .Z(n18754) );
  AND U32768 ( .A(n24791), .B(n24792), .Z(n24790) );
  NAND U32769 ( .A(o[403]), .B(n23579), .Z(n24792) );
  NANDN U32770 ( .A(n23580), .B(creg[403]), .Z(n24791) );
  NAND U32771 ( .A(n24793), .B(n18752), .Z(n13948) );
  NANDN U32772 ( .A(init), .B(m[404]), .Z(n18752) );
  AND U32773 ( .A(n24794), .B(n24795), .Z(n24793) );
  NAND U32774 ( .A(o[404]), .B(n23579), .Z(n24795) );
  NANDN U32775 ( .A(n23580), .B(creg[404]), .Z(n24794) );
  NAND U32776 ( .A(n24796), .B(n18750), .Z(n13947) );
  NANDN U32777 ( .A(init), .B(m[405]), .Z(n18750) );
  AND U32778 ( .A(n24797), .B(n24798), .Z(n24796) );
  NAND U32779 ( .A(o[405]), .B(n23579), .Z(n24798) );
  NANDN U32780 ( .A(n23580), .B(creg[405]), .Z(n24797) );
  NAND U32781 ( .A(n24799), .B(n18748), .Z(n13946) );
  NANDN U32782 ( .A(init), .B(m[406]), .Z(n18748) );
  AND U32783 ( .A(n24800), .B(n24801), .Z(n24799) );
  NAND U32784 ( .A(o[406]), .B(n23579), .Z(n24801) );
  NANDN U32785 ( .A(n23580), .B(creg[406]), .Z(n24800) );
  NAND U32786 ( .A(n24802), .B(n18746), .Z(n13945) );
  NANDN U32787 ( .A(init), .B(m[407]), .Z(n18746) );
  AND U32788 ( .A(n24803), .B(n24804), .Z(n24802) );
  NAND U32789 ( .A(o[407]), .B(n23579), .Z(n24804) );
  NANDN U32790 ( .A(n23580), .B(creg[407]), .Z(n24803) );
  NAND U32791 ( .A(n24805), .B(n18744), .Z(n13944) );
  NANDN U32792 ( .A(init), .B(m[408]), .Z(n18744) );
  AND U32793 ( .A(n24806), .B(n24807), .Z(n24805) );
  NAND U32794 ( .A(o[408]), .B(n23579), .Z(n24807) );
  NANDN U32795 ( .A(n23580), .B(creg[408]), .Z(n24806) );
  NAND U32796 ( .A(n24808), .B(n18742), .Z(n13943) );
  NANDN U32797 ( .A(init), .B(m[409]), .Z(n18742) );
  AND U32798 ( .A(n24809), .B(n24810), .Z(n24808) );
  NAND U32799 ( .A(o[409]), .B(n23579), .Z(n24810) );
  NANDN U32800 ( .A(n23580), .B(creg[409]), .Z(n24809) );
  NAND U32801 ( .A(n24811), .B(n18738), .Z(n13942) );
  NANDN U32802 ( .A(init), .B(m[410]), .Z(n18738) );
  AND U32803 ( .A(n24812), .B(n24813), .Z(n24811) );
  NAND U32804 ( .A(o[410]), .B(n23579), .Z(n24813) );
  NANDN U32805 ( .A(n23580), .B(creg[410]), .Z(n24812) );
  NAND U32806 ( .A(n24814), .B(n18736), .Z(n13941) );
  NANDN U32807 ( .A(init), .B(m[411]), .Z(n18736) );
  AND U32808 ( .A(n24815), .B(n24816), .Z(n24814) );
  NAND U32809 ( .A(o[411]), .B(n23579), .Z(n24816) );
  NANDN U32810 ( .A(n23580), .B(creg[411]), .Z(n24815) );
  NAND U32811 ( .A(n24817), .B(n18734), .Z(n13940) );
  NANDN U32812 ( .A(init), .B(m[412]), .Z(n18734) );
  AND U32813 ( .A(n24818), .B(n24819), .Z(n24817) );
  NAND U32814 ( .A(o[412]), .B(n23579), .Z(n24819) );
  NANDN U32815 ( .A(n23580), .B(creg[412]), .Z(n24818) );
  NAND U32816 ( .A(n24820), .B(n18732), .Z(n13939) );
  NANDN U32817 ( .A(init), .B(m[413]), .Z(n18732) );
  AND U32818 ( .A(n24821), .B(n24822), .Z(n24820) );
  NAND U32819 ( .A(o[413]), .B(n23579), .Z(n24822) );
  NANDN U32820 ( .A(n23580), .B(creg[413]), .Z(n24821) );
  NAND U32821 ( .A(n24823), .B(n18730), .Z(n13938) );
  NANDN U32822 ( .A(init), .B(m[414]), .Z(n18730) );
  AND U32823 ( .A(n24824), .B(n24825), .Z(n24823) );
  NAND U32824 ( .A(o[414]), .B(n23579), .Z(n24825) );
  NANDN U32825 ( .A(n23580), .B(creg[414]), .Z(n24824) );
  NAND U32826 ( .A(n24826), .B(n18728), .Z(n13937) );
  NANDN U32827 ( .A(init), .B(m[415]), .Z(n18728) );
  AND U32828 ( .A(n24827), .B(n24828), .Z(n24826) );
  NAND U32829 ( .A(o[415]), .B(n23579), .Z(n24828) );
  NANDN U32830 ( .A(n23580), .B(creg[415]), .Z(n24827) );
  NAND U32831 ( .A(n24829), .B(n18726), .Z(n13936) );
  NANDN U32832 ( .A(init), .B(m[416]), .Z(n18726) );
  AND U32833 ( .A(n24830), .B(n24831), .Z(n24829) );
  NAND U32834 ( .A(o[416]), .B(n23579), .Z(n24831) );
  NANDN U32835 ( .A(n23580), .B(creg[416]), .Z(n24830) );
  NAND U32836 ( .A(n24832), .B(n18724), .Z(n13935) );
  NANDN U32837 ( .A(init), .B(m[417]), .Z(n18724) );
  AND U32838 ( .A(n24833), .B(n24834), .Z(n24832) );
  NAND U32839 ( .A(o[417]), .B(n23579), .Z(n24834) );
  NANDN U32840 ( .A(n23580), .B(creg[417]), .Z(n24833) );
  NAND U32841 ( .A(n24835), .B(n18722), .Z(n13934) );
  NANDN U32842 ( .A(init), .B(m[418]), .Z(n18722) );
  AND U32843 ( .A(n24836), .B(n24837), .Z(n24835) );
  NAND U32844 ( .A(o[418]), .B(n23579), .Z(n24837) );
  NANDN U32845 ( .A(n23580), .B(creg[418]), .Z(n24836) );
  NAND U32846 ( .A(n24838), .B(n18720), .Z(n13933) );
  NANDN U32847 ( .A(init), .B(m[419]), .Z(n18720) );
  AND U32848 ( .A(n24839), .B(n24840), .Z(n24838) );
  NAND U32849 ( .A(o[419]), .B(n23579), .Z(n24840) );
  NANDN U32850 ( .A(n23580), .B(creg[419]), .Z(n24839) );
  NAND U32851 ( .A(n24841), .B(n18716), .Z(n13932) );
  NANDN U32852 ( .A(init), .B(m[420]), .Z(n18716) );
  AND U32853 ( .A(n24842), .B(n24843), .Z(n24841) );
  NAND U32854 ( .A(o[420]), .B(n23579), .Z(n24843) );
  NANDN U32855 ( .A(n23580), .B(creg[420]), .Z(n24842) );
  NAND U32856 ( .A(n24844), .B(n18714), .Z(n13931) );
  NANDN U32857 ( .A(init), .B(m[421]), .Z(n18714) );
  AND U32858 ( .A(n24845), .B(n24846), .Z(n24844) );
  NAND U32859 ( .A(o[421]), .B(n23579), .Z(n24846) );
  NANDN U32860 ( .A(n23580), .B(creg[421]), .Z(n24845) );
  NAND U32861 ( .A(n24847), .B(n18712), .Z(n13930) );
  NANDN U32862 ( .A(init), .B(m[422]), .Z(n18712) );
  AND U32863 ( .A(n24848), .B(n24849), .Z(n24847) );
  NAND U32864 ( .A(o[422]), .B(n23579), .Z(n24849) );
  NANDN U32865 ( .A(n23580), .B(creg[422]), .Z(n24848) );
  NAND U32866 ( .A(n24850), .B(n18710), .Z(n13929) );
  NANDN U32867 ( .A(init), .B(m[423]), .Z(n18710) );
  AND U32868 ( .A(n24851), .B(n24852), .Z(n24850) );
  NAND U32869 ( .A(o[423]), .B(n23579), .Z(n24852) );
  NANDN U32870 ( .A(n23580), .B(creg[423]), .Z(n24851) );
  NAND U32871 ( .A(n24853), .B(n18708), .Z(n13928) );
  NANDN U32872 ( .A(init), .B(m[424]), .Z(n18708) );
  AND U32873 ( .A(n24854), .B(n24855), .Z(n24853) );
  NAND U32874 ( .A(o[424]), .B(n23579), .Z(n24855) );
  NANDN U32875 ( .A(n23580), .B(creg[424]), .Z(n24854) );
  NAND U32876 ( .A(n24856), .B(n18706), .Z(n13927) );
  NANDN U32877 ( .A(init), .B(m[425]), .Z(n18706) );
  AND U32878 ( .A(n24857), .B(n24858), .Z(n24856) );
  NAND U32879 ( .A(o[425]), .B(n23579), .Z(n24858) );
  NANDN U32880 ( .A(n23580), .B(creg[425]), .Z(n24857) );
  NAND U32881 ( .A(n24859), .B(n18704), .Z(n13926) );
  NANDN U32882 ( .A(init), .B(m[426]), .Z(n18704) );
  AND U32883 ( .A(n24860), .B(n24861), .Z(n24859) );
  NAND U32884 ( .A(o[426]), .B(n23579), .Z(n24861) );
  NANDN U32885 ( .A(n23580), .B(creg[426]), .Z(n24860) );
  NAND U32886 ( .A(n24862), .B(n18702), .Z(n13925) );
  NANDN U32887 ( .A(init), .B(m[427]), .Z(n18702) );
  AND U32888 ( .A(n24863), .B(n24864), .Z(n24862) );
  NAND U32889 ( .A(o[427]), .B(n23579), .Z(n24864) );
  NANDN U32890 ( .A(n23580), .B(creg[427]), .Z(n24863) );
  NAND U32891 ( .A(n24865), .B(n18700), .Z(n13924) );
  NANDN U32892 ( .A(init), .B(m[428]), .Z(n18700) );
  AND U32893 ( .A(n24866), .B(n24867), .Z(n24865) );
  NAND U32894 ( .A(o[428]), .B(n23579), .Z(n24867) );
  NANDN U32895 ( .A(n23580), .B(creg[428]), .Z(n24866) );
  NAND U32896 ( .A(n24868), .B(n18698), .Z(n13923) );
  NANDN U32897 ( .A(init), .B(m[429]), .Z(n18698) );
  AND U32898 ( .A(n24869), .B(n24870), .Z(n24868) );
  NAND U32899 ( .A(o[429]), .B(n23579), .Z(n24870) );
  NANDN U32900 ( .A(n23580), .B(creg[429]), .Z(n24869) );
  NAND U32901 ( .A(n24871), .B(n18694), .Z(n13922) );
  NANDN U32902 ( .A(init), .B(m[430]), .Z(n18694) );
  AND U32903 ( .A(n24872), .B(n24873), .Z(n24871) );
  NAND U32904 ( .A(o[430]), .B(n23579), .Z(n24873) );
  NANDN U32905 ( .A(n23580), .B(creg[430]), .Z(n24872) );
  NAND U32906 ( .A(n24874), .B(n18692), .Z(n13921) );
  NANDN U32907 ( .A(init), .B(m[431]), .Z(n18692) );
  AND U32908 ( .A(n24875), .B(n24876), .Z(n24874) );
  NAND U32909 ( .A(o[431]), .B(n23579), .Z(n24876) );
  NANDN U32910 ( .A(n23580), .B(creg[431]), .Z(n24875) );
  NAND U32911 ( .A(n24877), .B(n18690), .Z(n13920) );
  NANDN U32912 ( .A(init), .B(m[432]), .Z(n18690) );
  AND U32913 ( .A(n24878), .B(n24879), .Z(n24877) );
  NAND U32914 ( .A(o[432]), .B(n23579), .Z(n24879) );
  NANDN U32915 ( .A(n23580), .B(creg[432]), .Z(n24878) );
  NAND U32916 ( .A(n24880), .B(n18688), .Z(n13919) );
  NANDN U32917 ( .A(init), .B(m[433]), .Z(n18688) );
  AND U32918 ( .A(n24881), .B(n24882), .Z(n24880) );
  NAND U32919 ( .A(o[433]), .B(n23579), .Z(n24882) );
  NANDN U32920 ( .A(n23580), .B(creg[433]), .Z(n24881) );
  NAND U32921 ( .A(n24883), .B(n18686), .Z(n13918) );
  NANDN U32922 ( .A(init), .B(m[434]), .Z(n18686) );
  AND U32923 ( .A(n24884), .B(n24885), .Z(n24883) );
  NAND U32924 ( .A(o[434]), .B(n23579), .Z(n24885) );
  NANDN U32925 ( .A(n23580), .B(creg[434]), .Z(n24884) );
  NAND U32926 ( .A(n24886), .B(n18684), .Z(n13917) );
  NANDN U32927 ( .A(init), .B(m[435]), .Z(n18684) );
  AND U32928 ( .A(n24887), .B(n24888), .Z(n24886) );
  NAND U32929 ( .A(o[435]), .B(n23579), .Z(n24888) );
  NANDN U32930 ( .A(n23580), .B(creg[435]), .Z(n24887) );
  NAND U32931 ( .A(n24889), .B(n18682), .Z(n13916) );
  NANDN U32932 ( .A(init), .B(m[436]), .Z(n18682) );
  AND U32933 ( .A(n24890), .B(n24891), .Z(n24889) );
  NAND U32934 ( .A(o[436]), .B(n23579), .Z(n24891) );
  NANDN U32935 ( .A(n23580), .B(creg[436]), .Z(n24890) );
  NAND U32936 ( .A(n24892), .B(n18680), .Z(n13915) );
  NANDN U32937 ( .A(init), .B(m[437]), .Z(n18680) );
  AND U32938 ( .A(n24893), .B(n24894), .Z(n24892) );
  NAND U32939 ( .A(o[437]), .B(n23579), .Z(n24894) );
  NANDN U32940 ( .A(n23580), .B(creg[437]), .Z(n24893) );
  NAND U32941 ( .A(n24895), .B(n18678), .Z(n13914) );
  NANDN U32942 ( .A(init), .B(m[438]), .Z(n18678) );
  AND U32943 ( .A(n24896), .B(n24897), .Z(n24895) );
  NAND U32944 ( .A(o[438]), .B(n23579), .Z(n24897) );
  NANDN U32945 ( .A(n23580), .B(creg[438]), .Z(n24896) );
  NAND U32946 ( .A(n24898), .B(n18676), .Z(n13913) );
  NANDN U32947 ( .A(init), .B(m[439]), .Z(n18676) );
  AND U32948 ( .A(n24899), .B(n24900), .Z(n24898) );
  NAND U32949 ( .A(o[439]), .B(n23579), .Z(n24900) );
  NANDN U32950 ( .A(n23580), .B(creg[439]), .Z(n24899) );
  NAND U32951 ( .A(n24901), .B(n18672), .Z(n13912) );
  NANDN U32952 ( .A(init), .B(m[440]), .Z(n18672) );
  AND U32953 ( .A(n24902), .B(n24903), .Z(n24901) );
  NAND U32954 ( .A(o[440]), .B(n23579), .Z(n24903) );
  NANDN U32955 ( .A(n23580), .B(creg[440]), .Z(n24902) );
  NAND U32956 ( .A(n24904), .B(n18670), .Z(n13911) );
  NANDN U32957 ( .A(init), .B(m[441]), .Z(n18670) );
  AND U32958 ( .A(n24905), .B(n24906), .Z(n24904) );
  NAND U32959 ( .A(o[441]), .B(n23579), .Z(n24906) );
  NANDN U32960 ( .A(n23580), .B(creg[441]), .Z(n24905) );
  NAND U32961 ( .A(n24907), .B(n18668), .Z(n13910) );
  NANDN U32962 ( .A(init), .B(m[442]), .Z(n18668) );
  AND U32963 ( .A(n24908), .B(n24909), .Z(n24907) );
  NAND U32964 ( .A(o[442]), .B(n23579), .Z(n24909) );
  NANDN U32965 ( .A(n23580), .B(creg[442]), .Z(n24908) );
  NAND U32966 ( .A(n24910), .B(n18666), .Z(n13909) );
  NANDN U32967 ( .A(init), .B(m[443]), .Z(n18666) );
  AND U32968 ( .A(n24911), .B(n24912), .Z(n24910) );
  NAND U32969 ( .A(o[443]), .B(n23579), .Z(n24912) );
  NANDN U32970 ( .A(n23580), .B(creg[443]), .Z(n24911) );
  NAND U32971 ( .A(n24913), .B(n18664), .Z(n13908) );
  NANDN U32972 ( .A(init), .B(m[444]), .Z(n18664) );
  AND U32973 ( .A(n24914), .B(n24915), .Z(n24913) );
  NAND U32974 ( .A(o[444]), .B(n23579), .Z(n24915) );
  NANDN U32975 ( .A(n23580), .B(creg[444]), .Z(n24914) );
  NAND U32976 ( .A(n24916), .B(n18662), .Z(n13907) );
  NANDN U32977 ( .A(init), .B(m[445]), .Z(n18662) );
  AND U32978 ( .A(n24917), .B(n24918), .Z(n24916) );
  NAND U32979 ( .A(o[445]), .B(n23579), .Z(n24918) );
  NANDN U32980 ( .A(n23580), .B(creg[445]), .Z(n24917) );
  NAND U32981 ( .A(n24919), .B(n18660), .Z(n13906) );
  NANDN U32982 ( .A(init), .B(m[446]), .Z(n18660) );
  AND U32983 ( .A(n24920), .B(n24921), .Z(n24919) );
  NAND U32984 ( .A(o[446]), .B(n23579), .Z(n24921) );
  NANDN U32985 ( .A(n23580), .B(creg[446]), .Z(n24920) );
  NAND U32986 ( .A(n24922), .B(n18658), .Z(n13905) );
  NANDN U32987 ( .A(init), .B(m[447]), .Z(n18658) );
  AND U32988 ( .A(n24923), .B(n24924), .Z(n24922) );
  NAND U32989 ( .A(o[447]), .B(n23579), .Z(n24924) );
  NANDN U32990 ( .A(n23580), .B(creg[447]), .Z(n24923) );
  NAND U32991 ( .A(n24925), .B(n18656), .Z(n13904) );
  NANDN U32992 ( .A(init), .B(m[448]), .Z(n18656) );
  AND U32993 ( .A(n24926), .B(n24927), .Z(n24925) );
  NAND U32994 ( .A(o[448]), .B(n23579), .Z(n24927) );
  NANDN U32995 ( .A(n23580), .B(creg[448]), .Z(n24926) );
  NAND U32996 ( .A(n24928), .B(n18654), .Z(n13903) );
  NANDN U32997 ( .A(init), .B(m[449]), .Z(n18654) );
  AND U32998 ( .A(n24929), .B(n24930), .Z(n24928) );
  NAND U32999 ( .A(o[449]), .B(n23579), .Z(n24930) );
  NANDN U33000 ( .A(n23580), .B(creg[449]), .Z(n24929) );
  NAND U33001 ( .A(n24931), .B(n18650), .Z(n13902) );
  NANDN U33002 ( .A(init), .B(m[450]), .Z(n18650) );
  AND U33003 ( .A(n24932), .B(n24933), .Z(n24931) );
  NAND U33004 ( .A(o[450]), .B(n23579), .Z(n24933) );
  NANDN U33005 ( .A(n23580), .B(creg[450]), .Z(n24932) );
  NAND U33006 ( .A(n24934), .B(n18648), .Z(n13901) );
  NANDN U33007 ( .A(init), .B(m[451]), .Z(n18648) );
  AND U33008 ( .A(n24935), .B(n24936), .Z(n24934) );
  NAND U33009 ( .A(o[451]), .B(n23579), .Z(n24936) );
  NANDN U33010 ( .A(n23580), .B(creg[451]), .Z(n24935) );
  NAND U33011 ( .A(n24937), .B(n18646), .Z(n13900) );
  NANDN U33012 ( .A(init), .B(m[452]), .Z(n18646) );
  AND U33013 ( .A(n24938), .B(n24939), .Z(n24937) );
  NAND U33014 ( .A(o[452]), .B(n23579), .Z(n24939) );
  NANDN U33015 ( .A(n23580), .B(creg[452]), .Z(n24938) );
  NAND U33016 ( .A(n24940), .B(n18644), .Z(n13899) );
  NANDN U33017 ( .A(init), .B(m[453]), .Z(n18644) );
  AND U33018 ( .A(n24941), .B(n24942), .Z(n24940) );
  NAND U33019 ( .A(o[453]), .B(n23579), .Z(n24942) );
  NANDN U33020 ( .A(n23580), .B(creg[453]), .Z(n24941) );
  NAND U33021 ( .A(n24943), .B(n18642), .Z(n13898) );
  NANDN U33022 ( .A(init), .B(m[454]), .Z(n18642) );
  AND U33023 ( .A(n24944), .B(n24945), .Z(n24943) );
  NAND U33024 ( .A(o[454]), .B(n23579), .Z(n24945) );
  NANDN U33025 ( .A(n23580), .B(creg[454]), .Z(n24944) );
  NAND U33026 ( .A(n24946), .B(n18640), .Z(n13897) );
  NANDN U33027 ( .A(init), .B(m[455]), .Z(n18640) );
  AND U33028 ( .A(n24947), .B(n24948), .Z(n24946) );
  NAND U33029 ( .A(o[455]), .B(n23579), .Z(n24948) );
  NANDN U33030 ( .A(n23580), .B(creg[455]), .Z(n24947) );
  NAND U33031 ( .A(n24949), .B(n18638), .Z(n13896) );
  NANDN U33032 ( .A(init), .B(m[456]), .Z(n18638) );
  AND U33033 ( .A(n24950), .B(n24951), .Z(n24949) );
  NAND U33034 ( .A(o[456]), .B(n23579), .Z(n24951) );
  NANDN U33035 ( .A(n23580), .B(creg[456]), .Z(n24950) );
  NAND U33036 ( .A(n24952), .B(n18636), .Z(n13895) );
  NANDN U33037 ( .A(init), .B(m[457]), .Z(n18636) );
  AND U33038 ( .A(n24953), .B(n24954), .Z(n24952) );
  NAND U33039 ( .A(o[457]), .B(n23579), .Z(n24954) );
  NANDN U33040 ( .A(n23580), .B(creg[457]), .Z(n24953) );
  NAND U33041 ( .A(n24955), .B(n18634), .Z(n13894) );
  NANDN U33042 ( .A(init), .B(m[458]), .Z(n18634) );
  AND U33043 ( .A(n24956), .B(n24957), .Z(n24955) );
  NAND U33044 ( .A(o[458]), .B(n23579), .Z(n24957) );
  NANDN U33045 ( .A(n23580), .B(creg[458]), .Z(n24956) );
  NAND U33046 ( .A(n24958), .B(n18632), .Z(n13893) );
  NANDN U33047 ( .A(init), .B(m[459]), .Z(n18632) );
  AND U33048 ( .A(n24959), .B(n24960), .Z(n24958) );
  NAND U33049 ( .A(o[459]), .B(n23579), .Z(n24960) );
  NANDN U33050 ( .A(n23580), .B(creg[459]), .Z(n24959) );
  NAND U33051 ( .A(n24961), .B(n18628), .Z(n13892) );
  NANDN U33052 ( .A(init), .B(m[460]), .Z(n18628) );
  AND U33053 ( .A(n24962), .B(n24963), .Z(n24961) );
  NAND U33054 ( .A(o[460]), .B(n23579), .Z(n24963) );
  NANDN U33055 ( .A(n23580), .B(creg[460]), .Z(n24962) );
  NAND U33056 ( .A(n24964), .B(n18626), .Z(n13891) );
  NANDN U33057 ( .A(init), .B(m[461]), .Z(n18626) );
  AND U33058 ( .A(n24965), .B(n24966), .Z(n24964) );
  NAND U33059 ( .A(o[461]), .B(n23579), .Z(n24966) );
  NANDN U33060 ( .A(n23580), .B(creg[461]), .Z(n24965) );
  NAND U33061 ( .A(n24967), .B(n18624), .Z(n13890) );
  NANDN U33062 ( .A(init), .B(m[462]), .Z(n18624) );
  AND U33063 ( .A(n24968), .B(n24969), .Z(n24967) );
  NAND U33064 ( .A(o[462]), .B(n23579), .Z(n24969) );
  NANDN U33065 ( .A(n23580), .B(creg[462]), .Z(n24968) );
  NAND U33066 ( .A(n24970), .B(n18622), .Z(n13889) );
  NANDN U33067 ( .A(init), .B(m[463]), .Z(n18622) );
  AND U33068 ( .A(n24971), .B(n24972), .Z(n24970) );
  NAND U33069 ( .A(o[463]), .B(n23579), .Z(n24972) );
  NANDN U33070 ( .A(n23580), .B(creg[463]), .Z(n24971) );
  NAND U33071 ( .A(n24973), .B(n18620), .Z(n13888) );
  NANDN U33072 ( .A(init), .B(m[464]), .Z(n18620) );
  AND U33073 ( .A(n24974), .B(n24975), .Z(n24973) );
  NAND U33074 ( .A(o[464]), .B(n23579), .Z(n24975) );
  NANDN U33075 ( .A(n23580), .B(creg[464]), .Z(n24974) );
  NAND U33076 ( .A(n24976), .B(n18618), .Z(n13887) );
  NANDN U33077 ( .A(init), .B(m[465]), .Z(n18618) );
  AND U33078 ( .A(n24977), .B(n24978), .Z(n24976) );
  NAND U33079 ( .A(o[465]), .B(n23579), .Z(n24978) );
  NANDN U33080 ( .A(n23580), .B(creg[465]), .Z(n24977) );
  NAND U33081 ( .A(n24979), .B(n18616), .Z(n13886) );
  NANDN U33082 ( .A(init), .B(m[466]), .Z(n18616) );
  AND U33083 ( .A(n24980), .B(n24981), .Z(n24979) );
  NAND U33084 ( .A(o[466]), .B(n23579), .Z(n24981) );
  NANDN U33085 ( .A(n23580), .B(creg[466]), .Z(n24980) );
  NAND U33086 ( .A(n24982), .B(n18614), .Z(n13885) );
  NANDN U33087 ( .A(init), .B(m[467]), .Z(n18614) );
  AND U33088 ( .A(n24983), .B(n24984), .Z(n24982) );
  NAND U33089 ( .A(o[467]), .B(n23579), .Z(n24984) );
  NANDN U33090 ( .A(n23580), .B(creg[467]), .Z(n24983) );
  NAND U33091 ( .A(n24985), .B(n18612), .Z(n13884) );
  NANDN U33092 ( .A(init), .B(m[468]), .Z(n18612) );
  AND U33093 ( .A(n24986), .B(n24987), .Z(n24985) );
  NAND U33094 ( .A(o[468]), .B(n23579), .Z(n24987) );
  NANDN U33095 ( .A(n23580), .B(creg[468]), .Z(n24986) );
  NAND U33096 ( .A(n24988), .B(n18610), .Z(n13883) );
  NANDN U33097 ( .A(init), .B(m[469]), .Z(n18610) );
  AND U33098 ( .A(n24989), .B(n24990), .Z(n24988) );
  NAND U33099 ( .A(o[469]), .B(n23579), .Z(n24990) );
  NANDN U33100 ( .A(n23580), .B(creg[469]), .Z(n24989) );
  NAND U33101 ( .A(n24991), .B(n18606), .Z(n13882) );
  NANDN U33102 ( .A(init), .B(m[470]), .Z(n18606) );
  AND U33103 ( .A(n24992), .B(n24993), .Z(n24991) );
  NAND U33104 ( .A(o[470]), .B(n23579), .Z(n24993) );
  NANDN U33105 ( .A(n23580), .B(creg[470]), .Z(n24992) );
  NAND U33106 ( .A(n24994), .B(n18604), .Z(n13881) );
  NANDN U33107 ( .A(init), .B(m[471]), .Z(n18604) );
  AND U33108 ( .A(n24995), .B(n24996), .Z(n24994) );
  NAND U33109 ( .A(o[471]), .B(n23579), .Z(n24996) );
  NANDN U33110 ( .A(n23580), .B(creg[471]), .Z(n24995) );
  NAND U33111 ( .A(n24997), .B(n18602), .Z(n13880) );
  NANDN U33112 ( .A(init), .B(m[472]), .Z(n18602) );
  AND U33113 ( .A(n24998), .B(n24999), .Z(n24997) );
  NAND U33114 ( .A(o[472]), .B(n23579), .Z(n24999) );
  NANDN U33115 ( .A(n23580), .B(creg[472]), .Z(n24998) );
  NAND U33116 ( .A(n25000), .B(n18600), .Z(n13879) );
  NANDN U33117 ( .A(init), .B(m[473]), .Z(n18600) );
  AND U33118 ( .A(n25001), .B(n25002), .Z(n25000) );
  NAND U33119 ( .A(o[473]), .B(n23579), .Z(n25002) );
  NANDN U33120 ( .A(n23580), .B(creg[473]), .Z(n25001) );
  NAND U33121 ( .A(n25003), .B(n18598), .Z(n13878) );
  NANDN U33122 ( .A(init), .B(m[474]), .Z(n18598) );
  AND U33123 ( .A(n25004), .B(n25005), .Z(n25003) );
  NAND U33124 ( .A(o[474]), .B(n23579), .Z(n25005) );
  NANDN U33125 ( .A(n23580), .B(creg[474]), .Z(n25004) );
  NAND U33126 ( .A(n25006), .B(n18596), .Z(n13877) );
  NANDN U33127 ( .A(init), .B(m[475]), .Z(n18596) );
  AND U33128 ( .A(n25007), .B(n25008), .Z(n25006) );
  NAND U33129 ( .A(o[475]), .B(n23579), .Z(n25008) );
  NANDN U33130 ( .A(n23580), .B(creg[475]), .Z(n25007) );
  NAND U33131 ( .A(n25009), .B(n18594), .Z(n13876) );
  NANDN U33132 ( .A(init), .B(m[476]), .Z(n18594) );
  AND U33133 ( .A(n25010), .B(n25011), .Z(n25009) );
  NAND U33134 ( .A(o[476]), .B(n23579), .Z(n25011) );
  NANDN U33135 ( .A(n23580), .B(creg[476]), .Z(n25010) );
  NAND U33136 ( .A(n25012), .B(n18592), .Z(n13875) );
  NANDN U33137 ( .A(init), .B(m[477]), .Z(n18592) );
  AND U33138 ( .A(n25013), .B(n25014), .Z(n25012) );
  NAND U33139 ( .A(o[477]), .B(n23579), .Z(n25014) );
  NANDN U33140 ( .A(n23580), .B(creg[477]), .Z(n25013) );
  NAND U33141 ( .A(n25015), .B(n18590), .Z(n13874) );
  NANDN U33142 ( .A(init), .B(m[478]), .Z(n18590) );
  AND U33143 ( .A(n25016), .B(n25017), .Z(n25015) );
  NAND U33144 ( .A(o[478]), .B(n23579), .Z(n25017) );
  NANDN U33145 ( .A(n23580), .B(creg[478]), .Z(n25016) );
  NAND U33146 ( .A(n25018), .B(n18588), .Z(n13873) );
  NANDN U33147 ( .A(init), .B(m[479]), .Z(n18588) );
  AND U33148 ( .A(n25019), .B(n25020), .Z(n25018) );
  NAND U33149 ( .A(o[479]), .B(n23579), .Z(n25020) );
  NANDN U33150 ( .A(n23580), .B(creg[479]), .Z(n25019) );
  NAND U33151 ( .A(n25021), .B(n18584), .Z(n13872) );
  NANDN U33152 ( .A(init), .B(m[480]), .Z(n18584) );
  AND U33153 ( .A(n25022), .B(n25023), .Z(n25021) );
  NAND U33154 ( .A(o[480]), .B(n23579), .Z(n25023) );
  NANDN U33155 ( .A(n23580), .B(creg[480]), .Z(n25022) );
  NAND U33156 ( .A(n25024), .B(n18582), .Z(n13871) );
  NANDN U33157 ( .A(init), .B(m[481]), .Z(n18582) );
  AND U33158 ( .A(n25025), .B(n25026), .Z(n25024) );
  NAND U33159 ( .A(o[481]), .B(n23579), .Z(n25026) );
  NANDN U33160 ( .A(n23580), .B(creg[481]), .Z(n25025) );
  NAND U33161 ( .A(n25027), .B(n18580), .Z(n13870) );
  NANDN U33162 ( .A(init), .B(m[482]), .Z(n18580) );
  AND U33163 ( .A(n25028), .B(n25029), .Z(n25027) );
  NAND U33164 ( .A(o[482]), .B(n23579), .Z(n25029) );
  NANDN U33165 ( .A(n23580), .B(creg[482]), .Z(n25028) );
  NAND U33166 ( .A(n25030), .B(n18578), .Z(n13869) );
  NANDN U33167 ( .A(init), .B(m[483]), .Z(n18578) );
  AND U33168 ( .A(n25031), .B(n25032), .Z(n25030) );
  NAND U33169 ( .A(o[483]), .B(n23579), .Z(n25032) );
  NANDN U33170 ( .A(n23580), .B(creg[483]), .Z(n25031) );
  NAND U33171 ( .A(n25033), .B(n18576), .Z(n13868) );
  NANDN U33172 ( .A(init), .B(m[484]), .Z(n18576) );
  AND U33173 ( .A(n25034), .B(n25035), .Z(n25033) );
  NAND U33174 ( .A(o[484]), .B(n23579), .Z(n25035) );
  NANDN U33175 ( .A(n23580), .B(creg[484]), .Z(n25034) );
  NAND U33176 ( .A(n25036), .B(n18574), .Z(n13867) );
  NANDN U33177 ( .A(init), .B(m[485]), .Z(n18574) );
  AND U33178 ( .A(n25037), .B(n25038), .Z(n25036) );
  NAND U33179 ( .A(o[485]), .B(n23579), .Z(n25038) );
  NANDN U33180 ( .A(n23580), .B(creg[485]), .Z(n25037) );
  NAND U33181 ( .A(n25039), .B(n18572), .Z(n13866) );
  NANDN U33182 ( .A(init), .B(m[486]), .Z(n18572) );
  AND U33183 ( .A(n25040), .B(n25041), .Z(n25039) );
  NAND U33184 ( .A(o[486]), .B(n23579), .Z(n25041) );
  NANDN U33185 ( .A(n23580), .B(creg[486]), .Z(n25040) );
  NAND U33186 ( .A(n25042), .B(n18570), .Z(n13865) );
  NANDN U33187 ( .A(init), .B(m[487]), .Z(n18570) );
  AND U33188 ( .A(n25043), .B(n25044), .Z(n25042) );
  NAND U33189 ( .A(o[487]), .B(n23579), .Z(n25044) );
  NANDN U33190 ( .A(n23580), .B(creg[487]), .Z(n25043) );
  NAND U33191 ( .A(n25045), .B(n18568), .Z(n13864) );
  NANDN U33192 ( .A(init), .B(m[488]), .Z(n18568) );
  AND U33193 ( .A(n25046), .B(n25047), .Z(n25045) );
  NAND U33194 ( .A(o[488]), .B(n23579), .Z(n25047) );
  NANDN U33195 ( .A(n23580), .B(creg[488]), .Z(n25046) );
  NAND U33196 ( .A(n25048), .B(n18566), .Z(n13863) );
  NANDN U33197 ( .A(init), .B(m[489]), .Z(n18566) );
  AND U33198 ( .A(n25049), .B(n25050), .Z(n25048) );
  NAND U33199 ( .A(o[489]), .B(n23579), .Z(n25050) );
  NANDN U33200 ( .A(n23580), .B(creg[489]), .Z(n25049) );
  NAND U33201 ( .A(n25051), .B(n18562), .Z(n13862) );
  NANDN U33202 ( .A(init), .B(m[490]), .Z(n18562) );
  AND U33203 ( .A(n25052), .B(n25053), .Z(n25051) );
  NAND U33204 ( .A(o[490]), .B(n23579), .Z(n25053) );
  NANDN U33205 ( .A(n23580), .B(creg[490]), .Z(n25052) );
  NAND U33206 ( .A(n25054), .B(n18560), .Z(n13861) );
  NANDN U33207 ( .A(init), .B(m[491]), .Z(n18560) );
  AND U33208 ( .A(n25055), .B(n25056), .Z(n25054) );
  NAND U33209 ( .A(o[491]), .B(n23579), .Z(n25056) );
  NANDN U33210 ( .A(n23580), .B(creg[491]), .Z(n25055) );
  NAND U33211 ( .A(n25057), .B(n18558), .Z(n13860) );
  NANDN U33212 ( .A(init), .B(m[492]), .Z(n18558) );
  AND U33213 ( .A(n25058), .B(n25059), .Z(n25057) );
  NAND U33214 ( .A(o[492]), .B(n23579), .Z(n25059) );
  NANDN U33215 ( .A(n23580), .B(creg[492]), .Z(n25058) );
  NAND U33216 ( .A(n25060), .B(n18556), .Z(n13859) );
  NANDN U33217 ( .A(init), .B(m[493]), .Z(n18556) );
  AND U33218 ( .A(n25061), .B(n25062), .Z(n25060) );
  NAND U33219 ( .A(o[493]), .B(n23579), .Z(n25062) );
  NANDN U33220 ( .A(n23580), .B(creg[493]), .Z(n25061) );
  NAND U33221 ( .A(n25063), .B(n18554), .Z(n13858) );
  NANDN U33222 ( .A(init), .B(m[494]), .Z(n18554) );
  AND U33223 ( .A(n25064), .B(n25065), .Z(n25063) );
  NAND U33224 ( .A(o[494]), .B(n23579), .Z(n25065) );
  NANDN U33225 ( .A(n23580), .B(creg[494]), .Z(n25064) );
  NAND U33226 ( .A(n25066), .B(n18552), .Z(n13857) );
  NANDN U33227 ( .A(init), .B(m[495]), .Z(n18552) );
  AND U33228 ( .A(n25067), .B(n25068), .Z(n25066) );
  NAND U33229 ( .A(o[495]), .B(n23579), .Z(n25068) );
  NANDN U33230 ( .A(n23580), .B(creg[495]), .Z(n25067) );
  NAND U33231 ( .A(n25069), .B(n18550), .Z(n13856) );
  NANDN U33232 ( .A(init), .B(m[496]), .Z(n18550) );
  AND U33233 ( .A(n25070), .B(n25071), .Z(n25069) );
  NAND U33234 ( .A(o[496]), .B(n23579), .Z(n25071) );
  NANDN U33235 ( .A(n23580), .B(creg[496]), .Z(n25070) );
  NAND U33236 ( .A(n25072), .B(n18548), .Z(n13855) );
  NANDN U33237 ( .A(init), .B(m[497]), .Z(n18548) );
  AND U33238 ( .A(n25073), .B(n25074), .Z(n25072) );
  NAND U33239 ( .A(o[497]), .B(n23579), .Z(n25074) );
  NANDN U33240 ( .A(n23580), .B(creg[497]), .Z(n25073) );
  NAND U33241 ( .A(n25075), .B(n18546), .Z(n13854) );
  NANDN U33242 ( .A(init), .B(m[498]), .Z(n18546) );
  AND U33243 ( .A(n25076), .B(n25077), .Z(n25075) );
  NAND U33244 ( .A(o[498]), .B(n23579), .Z(n25077) );
  NANDN U33245 ( .A(n23580), .B(creg[498]), .Z(n25076) );
  NAND U33246 ( .A(n25078), .B(n18544), .Z(n13853) );
  NANDN U33247 ( .A(init), .B(m[499]), .Z(n18544) );
  AND U33248 ( .A(n25079), .B(n25080), .Z(n25078) );
  NAND U33249 ( .A(o[499]), .B(n23579), .Z(n25080) );
  NANDN U33250 ( .A(n23580), .B(creg[499]), .Z(n25079) );
  NAND U33251 ( .A(n25081), .B(n18538), .Z(n13852) );
  NANDN U33252 ( .A(init), .B(m[500]), .Z(n18538) );
  AND U33253 ( .A(n25082), .B(n25083), .Z(n25081) );
  NAND U33254 ( .A(o[500]), .B(n23579), .Z(n25083) );
  NANDN U33255 ( .A(n23580), .B(creg[500]), .Z(n25082) );
  NAND U33256 ( .A(n25084), .B(n18536), .Z(n13851) );
  NANDN U33257 ( .A(init), .B(m[501]), .Z(n18536) );
  AND U33258 ( .A(n25085), .B(n25086), .Z(n25084) );
  NAND U33259 ( .A(o[501]), .B(n23579), .Z(n25086) );
  NANDN U33260 ( .A(n23580), .B(creg[501]), .Z(n25085) );
  NAND U33261 ( .A(n25087), .B(n18534), .Z(n13850) );
  NANDN U33262 ( .A(init), .B(m[502]), .Z(n18534) );
  AND U33263 ( .A(n25088), .B(n25089), .Z(n25087) );
  NAND U33264 ( .A(o[502]), .B(n23579), .Z(n25089) );
  NANDN U33265 ( .A(n23580), .B(creg[502]), .Z(n25088) );
  NAND U33266 ( .A(n25090), .B(n18532), .Z(n13849) );
  NANDN U33267 ( .A(init), .B(m[503]), .Z(n18532) );
  AND U33268 ( .A(n25091), .B(n25092), .Z(n25090) );
  NAND U33269 ( .A(o[503]), .B(n23579), .Z(n25092) );
  NANDN U33270 ( .A(n23580), .B(creg[503]), .Z(n25091) );
  NAND U33271 ( .A(n25093), .B(n18530), .Z(n13848) );
  NANDN U33272 ( .A(init), .B(m[504]), .Z(n18530) );
  AND U33273 ( .A(n25094), .B(n25095), .Z(n25093) );
  NAND U33274 ( .A(o[504]), .B(n23579), .Z(n25095) );
  NANDN U33275 ( .A(n23580), .B(creg[504]), .Z(n25094) );
  NAND U33276 ( .A(n25096), .B(n18528), .Z(n13847) );
  NANDN U33277 ( .A(init), .B(m[505]), .Z(n18528) );
  AND U33278 ( .A(n25097), .B(n25098), .Z(n25096) );
  NAND U33279 ( .A(o[505]), .B(n23579), .Z(n25098) );
  NANDN U33280 ( .A(n23580), .B(creg[505]), .Z(n25097) );
  NAND U33281 ( .A(n25099), .B(n18526), .Z(n13846) );
  NANDN U33282 ( .A(init), .B(m[506]), .Z(n18526) );
  AND U33283 ( .A(n25100), .B(n25101), .Z(n25099) );
  NAND U33284 ( .A(o[506]), .B(n23579), .Z(n25101) );
  NANDN U33285 ( .A(n23580), .B(creg[506]), .Z(n25100) );
  NAND U33286 ( .A(n25102), .B(n18524), .Z(n13845) );
  NANDN U33287 ( .A(init), .B(m[507]), .Z(n18524) );
  AND U33288 ( .A(n25103), .B(n25104), .Z(n25102) );
  NAND U33289 ( .A(o[507]), .B(n23579), .Z(n25104) );
  NANDN U33290 ( .A(n23580), .B(creg[507]), .Z(n25103) );
  NAND U33291 ( .A(n25105), .B(n18522), .Z(n13844) );
  NANDN U33292 ( .A(init), .B(m[508]), .Z(n18522) );
  AND U33293 ( .A(n25106), .B(n25107), .Z(n25105) );
  NAND U33294 ( .A(o[508]), .B(n23579), .Z(n25107) );
  NANDN U33295 ( .A(n23580), .B(creg[508]), .Z(n25106) );
  NAND U33296 ( .A(n25108), .B(n18520), .Z(n13843) );
  NANDN U33297 ( .A(init), .B(m[509]), .Z(n18520) );
  AND U33298 ( .A(n25109), .B(n25110), .Z(n25108) );
  NAND U33299 ( .A(o[509]), .B(n23579), .Z(n25110) );
  NANDN U33300 ( .A(n23580), .B(creg[509]), .Z(n25109) );
  NAND U33301 ( .A(n25111), .B(n18516), .Z(n13842) );
  NANDN U33302 ( .A(init), .B(m[510]), .Z(n18516) );
  AND U33303 ( .A(n25112), .B(n25113), .Z(n25111) );
  NAND U33304 ( .A(o[510]), .B(n23579), .Z(n25113) );
  NANDN U33305 ( .A(n23580), .B(creg[510]), .Z(n25112) );
  NAND U33306 ( .A(n25114), .B(n18514), .Z(n13841) );
  NANDN U33307 ( .A(init), .B(m[511]), .Z(n18514) );
  AND U33308 ( .A(n25115), .B(n25116), .Z(n25114) );
  NAND U33309 ( .A(o[511]), .B(n23579), .Z(n25116) );
  NANDN U33310 ( .A(n23580), .B(creg[511]), .Z(n25115) );
  NAND U33311 ( .A(n25117), .B(n18512), .Z(n13840) );
  NANDN U33312 ( .A(init), .B(m[512]), .Z(n18512) );
  AND U33313 ( .A(n25118), .B(n25119), .Z(n25117) );
  NAND U33314 ( .A(o[512]), .B(n23579), .Z(n25119) );
  NANDN U33315 ( .A(n23580), .B(creg[512]), .Z(n25118) );
  NAND U33316 ( .A(n25120), .B(n18510), .Z(n13839) );
  NANDN U33317 ( .A(init), .B(m[513]), .Z(n18510) );
  AND U33318 ( .A(n25121), .B(n25122), .Z(n25120) );
  NAND U33319 ( .A(o[513]), .B(n23579), .Z(n25122) );
  NANDN U33320 ( .A(n23580), .B(creg[513]), .Z(n25121) );
  NAND U33321 ( .A(n25123), .B(n18508), .Z(n13838) );
  NANDN U33322 ( .A(init), .B(m[514]), .Z(n18508) );
  AND U33323 ( .A(n25124), .B(n25125), .Z(n25123) );
  NAND U33324 ( .A(o[514]), .B(n23579), .Z(n25125) );
  NANDN U33325 ( .A(n23580), .B(creg[514]), .Z(n25124) );
  NAND U33326 ( .A(n25126), .B(n18506), .Z(n13837) );
  NANDN U33327 ( .A(init), .B(m[515]), .Z(n18506) );
  AND U33328 ( .A(n25127), .B(n25128), .Z(n25126) );
  NAND U33329 ( .A(o[515]), .B(n23579), .Z(n25128) );
  NANDN U33330 ( .A(n23580), .B(creg[515]), .Z(n25127) );
  NAND U33331 ( .A(n25129), .B(n18504), .Z(n13836) );
  NANDN U33332 ( .A(init), .B(m[516]), .Z(n18504) );
  AND U33333 ( .A(n25130), .B(n25131), .Z(n25129) );
  NAND U33334 ( .A(o[516]), .B(n23579), .Z(n25131) );
  NANDN U33335 ( .A(n23580), .B(creg[516]), .Z(n25130) );
  NAND U33336 ( .A(n25132), .B(n18502), .Z(n13835) );
  NANDN U33337 ( .A(init), .B(m[517]), .Z(n18502) );
  AND U33338 ( .A(n25133), .B(n25134), .Z(n25132) );
  NAND U33339 ( .A(o[517]), .B(n23579), .Z(n25134) );
  NANDN U33340 ( .A(n23580), .B(creg[517]), .Z(n25133) );
  NAND U33341 ( .A(n25135), .B(n18500), .Z(n13834) );
  NANDN U33342 ( .A(init), .B(m[518]), .Z(n18500) );
  AND U33343 ( .A(n25136), .B(n25137), .Z(n25135) );
  NAND U33344 ( .A(o[518]), .B(n23579), .Z(n25137) );
  NANDN U33345 ( .A(n23580), .B(creg[518]), .Z(n25136) );
  NAND U33346 ( .A(n25138), .B(n18498), .Z(n13833) );
  NANDN U33347 ( .A(init), .B(m[519]), .Z(n18498) );
  AND U33348 ( .A(n25139), .B(n25140), .Z(n25138) );
  NAND U33349 ( .A(o[519]), .B(n23579), .Z(n25140) );
  NANDN U33350 ( .A(n23580), .B(creg[519]), .Z(n25139) );
  NAND U33351 ( .A(n25141), .B(n18494), .Z(n13832) );
  NANDN U33352 ( .A(init), .B(m[520]), .Z(n18494) );
  AND U33353 ( .A(n25142), .B(n25143), .Z(n25141) );
  NAND U33354 ( .A(o[520]), .B(n23579), .Z(n25143) );
  NANDN U33355 ( .A(n23580), .B(creg[520]), .Z(n25142) );
  NAND U33356 ( .A(n25144), .B(n18492), .Z(n13831) );
  NANDN U33357 ( .A(init), .B(m[521]), .Z(n18492) );
  AND U33358 ( .A(n25145), .B(n25146), .Z(n25144) );
  NAND U33359 ( .A(o[521]), .B(n23579), .Z(n25146) );
  NANDN U33360 ( .A(n23580), .B(creg[521]), .Z(n25145) );
  NAND U33361 ( .A(n25147), .B(n18490), .Z(n13830) );
  NANDN U33362 ( .A(init), .B(m[522]), .Z(n18490) );
  AND U33363 ( .A(n25148), .B(n25149), .Z(n25147) );
  NAND U33364 ( .A(o[522]), .B(n23579), .Z(n25149) );
  NANDN U33365 ( .A(n23580), .B(creg[522]), .Z(n25148) );
  NAND U33366 ( .A(n25150), .B(n18488), .Z(n13829) );
  NANDN U33367 ( .A(init), .B(m[523]), .Z(n18488) );
  AND U33368 ( .A(n25151), .B(n25152), .Z(n25150) );
  NAND U33369 ( .A(o[523]), .B(n23579), .Z(n25152) );
  NANDN U33370 ( .A(n23580), .B(creg[523]), .Z(n25151) );
  NAND U33371 ( .A(n25153), .B(n18486), .Z(n13828) );
  NANDN U33372 ( .A(init), .B(m[524]), .Z(n18486) );
  AND U33373 ( .A(n25154), .B(n25155), .Z(n25153) );
  NAND U33374 ( .A(o[524]), .B(n23579), .Z(n25155) );
  NANDN U33375 ( .A(n23580), .B(creg[524]), .Z(n25154) );
  NAND U33376 ( .A(n25156), .B(n18484), .Z(n13827) );
  NANDN U33377 ( .A(init), .B(m[525]), .Z(n18484) );
  AND U33378 ( .A(n25157), .B(n25158), .Z(n25156) );
  NAND U33379 ( .A(o[525]), .B(n23579), .Z(n25158) );
  NANDN U33380 ( .A(n23580), .B(creg[525]), .Z(n25157) );
  NAND U33381 ( .A(n25159), .B(n18482), .Z(n13826) );
  NANDN U33382 ( .A(init), .B(m[526]), .Z(n18482) );
  AND U33383 ( .A(n25160), .B(n25161), .Z(n25159) );
  NAND U33384 ( .A(o[526]), .B(n23579), .Z(n25161) );
  NANDN U33385 ( .A(n23580), .B(creg[526]), .Z(n25160) );
  NAND U33386 ( .A(n25162), .B(n18480), .Z(n13825) );
  NANDN U33387 ( .A(init), .B(m[527]), .Z(n18480) );
  AND U33388 ( .A(n25163), .B(n25164), .Z(n25162) );
  NAND U33389 ( .A(o[527]), .B(n23579), .Z(n25164) );
  NANDN U33390 ( .A(n23580), .B(creg[527]), .Z(n25163) );
  NAND U33391 ( .A(n25165), .B(n18478), .Z(n13824) );
  NANDN U33392 ( .A(init), .B(m[528]), .Z(n18478) );
  AND U33393 ( .A(n25166), .B(n25167), .Z(n25165) );
  NAND U33394 ( .A(o[528]), .B(n23579), .Z(n25167) );
  NANDN U33395 ( .A(n23580), .B(creg[528]), .Z(n25166) );
  NAND U33396 ( .A(n25168), .B(n18476), .Z(n13823) );
  NANDN U33397 ( .A(init), .B(m[529]), .Z(n18476) );
  AND U33398 ( .A(n25169), .B(n25170), .Z(n25168) );
  NAND U33399 ( .A(o[529]), .B(n23579), .Z(n25170) );
  NANDN U33400 ( .A(n23580), .B(creg[529]), .Z(n25169) );
  NAND U33401 ( .A(n25171), .B(n18472), .Z(n13822) );
  NANDN U33402 ( .A(init), .B(m[530]), .Z(n18472) );
  AND U33403 ( .A(n25172), .B(n25173), .Z(n25171) );
  NAND U33404 ( .A(o[530]), .B(n23579), .Z(n25173) );
  NANDN U33405 ( .A(n23580), .B(creg[530]), .Z(n25172) );
  NAND U33406 ( .A(n25174), .B(n18470), .Z(n13821) );
  NANDN U33407 ( .A(init), .B(m[531]), .Z(n18470) );
  AND U33408 ( .A(n25175), .B(n25176), .Z(n25174) );
  NAND U33409 ( .A(o[531]), .B(n23579), .Z(n25176) );
  NANDN U33410 ( .A(n23580), .B(creg[531]), .Z(n25175) );
  NAND U33411 ( .A(n25177), .B(n18468), .Z(n13820) );
  NANDN U33412 ( .A(init), .B(m[532]), .Z(n18468) );
  AND U33413 ( .A(n25178), .B(n25179), .Z(n25177) );
  NAND U33414 ( .A(o[532]), .B(n23579), .Z(n25179) );
  NANDN U33415 ( .A(n23580), .B(creg[532]), .Z(n25178) );
  NAND U33416 ( .A(n25180), .B(n18466), .Z(n13819) );
  NANDN U33417 ( .A(init), .B(m[533]), .Z(n18466) );
  AND U33418 ( .A(n25181), .B(n25182), .Z(n25180) );
  NAND U33419 ( .A(o[533]), .B(n23579), .Z(n25182) );
  NANDN U33420 ( .A(n23580), .B(creg[533]), .Z(n25181) );
  NAND U33421 ( .A(n25183), .B(n18464), .Z(n13818) );
  NANDN U33422 ( .A(init), .B(m[534]), .Z(n18464) );
  AND U33423 ( .A(n25184), .B(n25185), .Z(n25183) );
  NAND U33424 ( .A(o[534]), .B(n23579), .Z(n25185) );
  NANDN U33425 ( .A(n23580), .B(creg[534]), .Z(n25184) );
  NAND U33426 ( .A(n25186), .B(n18462), .Z(n13817) );
  NANDN U33427 ( .A(init), .B(m[535]), .Z(n18462) );
  AND U33428 ( .A(n25187), .B(n25188), .Z(n25186) );
  NAND U33429 ( .A(o[535]), .B(n23579), .Z(n25188) );
  NANDN U33430 ( .A(n23580), .B(creg[535]), .Z(n25187) );
  NAND U33431 ( .A(n25189), .B(n18460), .Z(n13816) );
  NANDN U33432 ( .A(init), .B(m[536]), .Z(n18460) );
  AND U33433 ( .A(n25190), .B(n25191), .Z(n25189) );
  NAND U33434 ( .A(o[536]), .B(n23579), .Z(n25191) );
  NANDN U33435 ( .A(n23580), .B(creg[536]), .Z(n25190) );
  NAND U33436 ( .A(n25192), .B(n18458), .Z(n13815) );
  NANDN U33437 ( .A(init), .B(m[537]), .Z(n18458) );
  AND U33438 ( .A(n25193), .B(n25194), .Z(n25192) );
  NAND U33439 ( .A(o[537]), .B(n23579), .Z(n25194) );
  NANDN U33440 ( .A(n23580), .B(creg[537]), .Z(n25193) );
  NAND U33441 ( .A(n25195), .B(n18456), .Z(n13814) );
  NANDN U33442 ( .A(init), .B(m[538]), .Z(n18456) );
  AND U33443 ( .A(n25196), .B(n25197), .Z(n25195) );
  NAND U33444 ( .A(o[538]), .B(n23579), .Z(n25197) );
  NANDN U33445 ( .A(n23580), .B(creg[538]), .Z(n25196) );
  NAND U33446 ( .A(n25198), .B(n18454), .Z(n13813) );
  NANDN U33447 ( .A(init), .B(m[539]), .Z(n18454) );
  AND U33448 ( .A(n25199), .B(n25200), .Z(n25198) );
  NAND U33449 ( .A(o[539]), .B(n23579), .Z(n25200) );
  NANDN U33450 ( .A(n23580), .B(creg[539]), .Z(n25199) );
  NAND U33451 ( .A(n25201), .B(n18450), .Z(n13812) );
  NANDN U33452 ( .A(init), .B(m[540]), .Z(n18450) );
  AND U33453 ( .A(n25202), .B(n25203), .Z(n25201) );
  NAND U33454 ( .A(o[540]), .B(n23579), .Z(n25203) );
  NANDN U33455 ( .A(n23580), .B(creg[540]), .Z(n25202) );
  NAND U33456 ( .A(n25204), .B(n18448), .Z(n13811) );
  NANDN U33457 ( .A(init), .B(m[541]), .Z(n18448) );
  AND U33458 ( .A(n25205), .B(n25206), .Z(n25204) );
  NAND U33459 ( .A(o[541]), .B(n23579), .Z(n25206) );
  NANDN U33460 ( .A(n23580), .B(creg[541]), .Z(n25205) );
  NAND U33461 ( .A(n25207), .B(n18446), .Z(n13810) );
  NANDN U33462 ( .A(init), .B(m[542]), .Z(n18446) );
  AND U33463 ( .A(n25208), .B(n25209), .Z(n25207) );
  NAND U33464 ( .A(o[542]), .B(n23579), .Z(n25209) );
  NANDN U33465 ( .A(n23580), .B(creg[542]), .Z(n25208) );
  NAND U33466 ( .A(n25210), .B(n18444), .Z(n13809) );
  NANDN U33467 ( .A(init), .B(m[543]), .Z(n18444) );
  AND U33468 ( .A(n25211), .B(n25212), .Z(n25210) );
  NAND U33469 ( .A(o[543]), .B(n23579), .Z(n25212) );
  NANDN U33470 ( .A(n23580), .B(creg[543]), .Z(n25211) );
  NAND U33471 ( .A(n25213), .B(n18442), .Z(n13808) );
  NANDN U33472 ( .A(init), .B(m[544]), .Z(n18442) );
  AND U33473 ( .A(n25214), .B(n25215), .Z(n25213) );
  NAND U33474 ( .A(o[544]), .B(n23579), .Z(n25215) );
  NANDN U33475 ( .A(n23580), .B(creg[544]), .Z(n25214) );
  NAND U33476 ( .A(n25216), .B(n18440), .Z(n13807) );
  NANDN U33477 ( .A(init), .B(m[545]), .Z(n18440) );
  AND U33478 ( .A(n25217), .B(n25218), .Z(n25216) );
  NAND U33479 ( .A(o[545]), .B(n23579), .Z(n25218) );
  NANDN U33480 ( .A(n23580), .B(creg[545]), .Z(n25217) );
  NAND U33481 ( .A(n25219), .B(n18438), .Z(n13806) );
  NANDN U33482 ( .A(init), .B(m[546]), .Z(n18438) );
  AND U33483 ( .A(n25220), .B(n25221), .Z(n25219) );
  NAND U33484 ( .A(o[546]), .B(n23579), .Z(n25221) );
  NANDN U33485 ( .A(n23580), .B(creg[546]), .Z(n25220) );
  NAND U33486 ( .A(n25222), .B(n18436), .Z(n13805) );
  NANDN U33487 ( .A(init), .B(m[547]), .Z(n18436) );
  AND U33488 ( .A(n25223), .B(n25224), .Z(n25222) );
  NAND U33489 ( .A(o[547]), .B(n23579), .Z(n25224) );
  NANDN U33490 ( .A(n23580), .B(creg[547]), .Z(n25223) );
  NAND U33491 ( .A(n25225), .B(n18434), .Z(n13804) );
  NANDN U33492 ( .A(init), .B(m[548]), .Z(n18434) );
  AND U33493 ( .A(n25226), .B(n25227), .Z(n25225) );
  NAND U33494 ( .A(o[548]), .B(n23579), .Z(n25227) );
  NANDN U33495 ( .A(n23580), .B(creg[548]), .Z(n25226) );
  NAND U33496 ( .A(n25228), .B(n18432), .Z(n13803) );
  NANDN U33497 ( .A(init), .B(m[549]), .Z(n18432) );
  AND U33498 ( .A(n25229), .B(n25230), .Z(n25228) );
  NAND U33499 ( .A(o[549]), .B(n23579), .Z(n25230) );
  NANDN U33500 ( .A(n23580), .B(creg[549]), .Z(n25229) );
  NAND U33501 ( .A(n25231), .B(n18428), .Z(n13802) );
  NANDN U33502 ( .A(init), .B(m[550]), .Z(n18428) );
  AND U33503 ( .A(n25232), .B(n25233), .Z(n25231) );
  NAND U33504 ( .A(o[550]), .B(n23579), .Z(n25233) );
  NANDN U33505 ( .A(n23580), .B(creg[550]), .Z(n25232) );
  NAND U33506 ( .A(n25234), .B(n18426), .Z(n13801) );
  NANDN U33507 ( .A(init), .B(m[551]), .Z(n18426) );
  AND U33508 ( .A(n25235), .B(n25236), .Z(n25234) );
  NAND U33509 ( .A(o[551]), .B(n23579), .Z(n25236) );
  NANDN U33510 ( .A(n23580), .B(creg[551]), .Z(n25235) );
  NAND U33511 ( .A(n25237), .B(n18424), .Z(n13800) );
  NANDN U33512 ( .A(init), .B(m[552]), .Z(n18424) );
  AND U33513 ( .A(n25238), .B(n25239), .Z(n25237) );
  NAND U33514 ( .A(o[552]), .B(n23579), .Z(n25239) );
  NANDN U33515 ( .A(n23580), .B(creg[552]), .Z(n25238) );
  NAND U33516 ( .A(n25240), .B(n18422), .Z(n13799) );
  NANDN U33517 ( .A(init), .B(m[553]), .Z(n18422) );
  AND U33518 ( .A(n25241), .B(n25242), .Z(n25240) );
  NAND U33519 ( .A(o[553]), .B(n23579), .Z(n25242) );
  NANDN U33520 ( .A(n23580), .B(creg[553]), .Z(n25241) );
  NAND U33521 ( .A(n25243), .B(n18420), .Z(n13798) );
  NANDN U33522 ( .A(init), .B(m[554]), .Z(n18420) );
  AND U33523 ( .A(n25244), .B(n25245), .Z(n25243) );
  NAND U33524 ( .A(o[554]), .B(n23579), .Z(n25245) );
  NANDN U33525 ( .A(n23580), .B(creg[554]), .Z(n25244) );
  NAND U33526 ( .A(n25246), .B(n18418), .Z(n13797) );
  NANDN U33527 ( .A(init), .B(m[555]), .Z(n18418) );
  AND U33528 ( .A(n25247), .B(n25248), .Z(n25246) );
  NAND U33529 ( .A(o[555]), .B(n23579), .Z(n25248) );
  NANDN U33530 ( .A(n23580), .B(creg[555]), .Z(n25247) );
  NAND U33531 ( .A(n25249), .B(n18416), .Z(n13796) );
  NANDN U33532 ( .A(init), .B(m[556]), .Z(n18416) );
  AND U33533 ( .A(n25250), .B(n25251), .Z(n25249) );
  NAND U33534 ( .A(o[556]), .B(n23579), .Z(n25251) );
  NANDN U33535 ( .A(n23580), .B(creg[556]), .Z(n25250) );
  NAND U33536 ( .A(n25252), .B(n18414), .Z(n13795) );
  NANDN U33537 ( .A(init), .B(m[557]), .Z(n18414) );
  AND U33538 ( .A(n25253), .B(n25254), .Z(n25252) );
  NAND U33539 ( .A(o[557]), .B(n23579), .Z(n25254) );
  NANDN U33540 ( .A(n23580), .B(creg[557]), .Z(n25253) );
  NAND U33541 ( .A(n25255), .B(n18412), .Z(n13794) );
  NANDN U33542 ( .A(init), .B(m[558]), .Z(n18412) );
  AND U33543 ( .A(n25256), .B(n25257), .Z(n25255) );
  NAND U33544 ( .A(o[558]), .B(n23579), .Z(n25257) );
  NANDN U33545 ( .A(n23580), .B(creg[558]), .Z(n25256) );
  NAND U33546 ( .A(n25258), .B(n18410), .Z(n13793) );
  NANDN U33547 ( .A(init), .B(m[559]), .Z(n18410) );
  AND U33548 ( .A(n25259), .B(n25260), .Z(n25258) );
  NAND U33549 ( .A(o[559]), .B(n23579), .Z(n25260) );
  NANDN U33550 ( .A(n23580), .B(creg[559]), .Z(n25259) );
  NAND U33551 ( .A(n25261), .B(n18406), .Z(n13792) );
  NANDN U33552 ( .A(init), .B(m[560]), .Z(n18406) );
  AND U33553 ( .A(n25262), .B(n25263), .Z(n25261) );
  NAND U33554 ( .A(o[560]), .B(n23579), .Z(n25263) );
  NANDN U33555 ( .A(n23580), .B(creg[560]), .Z(n25262) );
  NAND U33556 ( .A(n25264), .B(n18404), .Z(n13791) );
  NANDN U33557 ( .A(init), .B(m[561]), .Z(n18404) );
  AND U33558 ( .A(n25265), .B(n25266), .Z(n25264) );
  NAND U33559 ( .A(o[561]), .B(n23579), .Z(n25266) );
  NANDN U33560 ( .A(n23580), .B(creg[561]), .Z(n25265) );
  NAND U33561 ( .A(n25267), .B(n18402), .Z(n13790) );
  NANDN U33562 ( .A(init), .B(m[562]), .Z(n18402) );
  AND U33563 ( .A(n25268), .B(n25269), .Z(n25267) );
  NAND U33564 ( .A(o[562]), .B(n23579), .Z(n25269) );
  NANDN U33565 ( .A(n23580), .B(creg[562]), .Z(n25268) );
  NAND U33566 ( .A(n25270), .B(n18400), .Z(n13789) );
  NANDN U33567 ( .A(init), .B(m[563]), .Z(n18400) );
  AND U33568 ( .A(n25271), .B(n25272), .Z(n25270) );
  NAND U33569 ( .A(o[563]), .B(n23579), .Z(n25272) );
  NANDN U33570 ( .A(n23580), .B(creg[563]), .Z(n25271) );
  NAND U33571 ( .A(n25273), .B(n18398), .Z(n13788) );
  NANDN U33572 ( .A(init), .B(m[564]), .Z(n18398) );
  AND U33573 ( .A(n25274), .B(n25275), .Z(n25273) );
  NAND U33574 ( .A(o[564]), .B(n23579), .Z(n25275) );
  NANDN U33575 ( .A(n23580), .B(creg[564]), .Z(n25274) );
  NAND U33576 ( .A(n25276), .B(n18396), .Z(n13787) );
  NANDN U33577 ( .A(init), .B(m[565]), .Z(n18396) );
  AND U33578 ( .A(n25277), .B(n25278), .Z(n25276) );
  NAND U33579 ( .A(o[565]), .B(n23579), .Z(n25278) );
  NANDN U33580 ( .A(n23580), .B(creg[565]), .Z(n25277) );
  NAND U33581 ( .A(n25279), .B(n18394), .Z(n13786) );
  NANDN U33582 ( .A(init), .B(m[566]), .Z(n18394) );
  AND U33583 ( .A(n25280), .B(n25281), .Z(n25279) );
  NAND U33584 ( .A(o[566]), .B(n23579), .Z(n25281) );
  NANDN U33585 ( .A(n23580), .B(creg[566]), .Z(n25280) );
  NAND U33586 ( .A(n25282), .B(n18392), .Z(n13785) );
  NANDN U33587 ( .A(init), .B(m[567]), .Z(n18392) );
  AND U33588 ( .A(n25283), .B(n25284), .Z(n25282) );
  NAND U33589 ( .A(o[567]), .B(n23579), .Z(n25284) );
  NANDN U33590 ( .A(n23580), .B(creg[567]), .Z(n25283) );
  NAND U33591 ( .A(n25285), .B(n18390), .Z(n13784) );
  NANDN U33592 ( .A(init), .B(m[568]), .Z(n18390) );
  AND U33593 ( .A(n25286), .B(n25287), .Z(n25285) );
  NAND U33594 ( .A(o[568]), .B(n23579), .Z(n25287) );
  NANDN U33595 ( .A(n23580), .B(creg[568]), .Z(n25286) );
  NAND U33596 ( .A(n25288), .B(n18388), .Z(n13783) );
  NANDN U33597 ( .A(init), .B(m[569]), .Z(n18388) );
  AND U33598 ( .A(n25289), .B(n25290), .Z(n25288) );
  NAND U33599 ( .A(o[569]), .B(n23579), .Z(n25290) );
  NANDN U33600 ( .A(n23580), .B(creg[569]), .Z(n25289) );
  NAND U33601 ( .A(n25291), .B(n18384), .Z(n13782) );
  NANDN U33602 ( .A(init), .B(m[570]), .Z(n18384) );
  AND U33603 ( .A(n25292), .B(n25293), .Z(n25291) );
  NAND U33604 ( .A(o[570]), .B(n23579), .Z(n25293) );
  NANDN U33605 ( .A(n23580), .B(creg[570]), .Z(n25292) );
  NAND U33606 ( .A(n25294), .B(n18382), .Z(n13781) );
  NANDN U33607 ( .A(init), .B(m[571]), .Z(n18382) );
  AND U33608 ( .A(n25295), .B(n25296), .Z(n25294) );
  NAND U33609 ( .A(o[571]), .B(n23579), .Z(n25296) );
  NANDN U33610 ( .A(n23580), .B(creg[571]), .Z(n25295) );
  NAND U33611 ( .A(n25297), .B(n18380), .Z(n13780) );
  NANDN U33612 ( .A(init), .B(m[572]), .Z(n18380) );
  AND U33613 ( .A(n25298), .B(n25299), .Z(n25297) );
  NAND U33614 ( .A(o[572]), .B(n23579), .Z(n25299) );
  NANDN U33615 ( .A(n23580), .B(creg[572]), .Z(n25298) );
  NAND U33616 ( .A(n25300), .B(n18378), .Z(n13779) );
  NANDN U33617 ( .A(init), .B(m[573]), .Z(n18378) );
  AND U33618 ( .A(n25301), .B(n25302), .Z(n25300) );
  NAND U33619 ( .A(o[573]), .B(n23579), .Z(n25302) );
  NANDN U33620 ( .A(n23580), .B(creg[573]), .Z(n25301) );
  NAND U33621 ( .A(n25303), .B(n18376), .Z(n13778) );
  NANDN U33622 ( .A(init), .B(m[574]), .Z(n18376) );
  AND U33623 ( .A(n25304), .B(n25305), .Z(n25303) );
  NAND U33624 ( .A(o[574]), .B(n23579), .Z(n25305) );
  NANDN U33625 ( .A(n23580), .B(creg[574]), .Z(n25304) );
  NAND U33626 ( .A(n25306), .B(n18374), .Z(n13777) );
  NANDN U33627 ( .A(init), .B(m[575]), .Z(n18374) );
  AND U33628 ( .A(n25307), .B(n25308), .Z(n25306) );
  NAND U33629 ( .A(o[575]), .B(n23579), .Z(n25308) );
  NANDN U33630 ( .A(n23580), .B(creg[575]), .Z(n25307) );
  NAND U33631 ( .A(n25309), .B(n18372), .Z(n13776) );
  NANDN U33632 ( .A(init), .B(m[576]), .Z(n18372) );
  AND U33633 ( .A(n25310), .B(n25311), .Z(n25309) );
  NAND U33634 ( .A(o[576]), .B(n23579), .Z(n25311) );
  NANDN U33635 ( .A(n23580), .B(creg[576]), .Z(n25310) );
  NAND U33636 ( .A(n25312), .B(n18370), .Z(n13775) );
  NANDN U33637 ( .A(init), .B(m[577]), .Z(n18370) );
  AND U33638 ( .A(n25313), .B(n25314), .Z(n25312) );
  NAND U33639 ( .A(o[577]), .B(n23579), .Z(n25314) );
  NANDN U33640 ( .A(n23580), .B(creg[577]), .Z(n25313) );
  NAND U33641 ( .A(n25315), .B(n18368), .Z(n13774) );
  NANDN U33642 ( .A(init), .B(m[578]), .Z(n18368) );
  AND U33643 ( .A(n25316), .B(n25317), .Z(n25315) );
  NAND U33644 ( .A(o[578]), .B(n23579), .Z(n25317) );
  NANDN U33645 ( .A(n23580), .B(creg[578]), .Z(n25316) );
  NAND U33646 ( .A(n25318), .B(n18366), .Z(n13773) );
  NANDN U33647 ( .A(init), .B(m[579]), .Z(n18366) );
  AND U33648 ( .A(n25319), .B(n25320), .Z(n25318) );
  NAND U33649 ( .A(o[579]), .B(n23579), .Z(n25320) );
  NANDN U33650 ( .A(n23580), .B(creg[579]), .Z(n25319) );
  NAND U33651 ( .A(n25321), .B(n18362), .Z(n13772) );
  NANDN U33652 ( .A(init), .B(m[580]), .Z(n18362) );
  AND U33653 ( .A(n25322), .B(n25323), .Z(n25321) );
  NAND U33654 ( .A(o[580]), .B(n23579), .Z(n25323) );
  NANDN U33655 ( .A(n23580), .B(creg[580]), .Z(n25322) );
  NAND U33656 ( .A(n25324), .B(n18360), .Z(n13771) );
  NANDN U33657 ( .A(init), .B(m[581]), .Z(n18360) );
  AND U33658 ( .A(n25325), .B(n25326), .Z(n25324) );
  NAND U33659 ( .A(o[581]), .B(n23579), .Z(n25326) );
  NANDN U33660 ( .A(n23580), .B(creg[581]), .Z(n25325) );
  NAND U33661 ( .A(n25327), .B(n18358), .Z(n13770) );
  NANDN U33662 ( .A(init), .B(m[582]), .Z(n18358) );
  AND U33663 ( .A(n25328), .B(n25329), .Z(n25327) );
  NAND U33664 ( .A(o[582]), .B(n23579), .Z(n25329) );
  NANDN U33665 ( .A(n23580), .B(creg[582]), .Z(n25328) );
  NAND U33666 ( .A(n25330), .B(n18356), .Z(n13769) );
  NANDN U33667 ( .A(init), .B(m[583]), .Z(n18356) );
  AND U33668 ( .A(n25331), .B(n25332), .Z(n25330) );
  NAND U33669 ( .A(o[583]), .B(n23579), .Z(n25332) );
  NANDN U33670 ( .A(n23580), .B(creg[583]), .Z(n25331) );
  NAND U33671 ( .A(n25333), .B(n18354), .Z(n13768) );
  NANDN U33672 ( .A(init), .B(m[584]), .Z(n18354) );
  AND U33673 ( .A(n25334), .B(n25335), .Z(n25333) );
  NAND U33674 ( .A(o[584]), .B(n23579), .Z(n25335) );
  NANDN U33675 ( .A(n23580), .B(creg[584]), .Z(n25334) );
  NAND U33676 ( .A(n25336), .B(n18352), .Z(n13767) );
  NANDN U33677 ( .A(init), .B(m[585]), .Z(n18352) );
  AND U33678 ( .A(n25337), .B(n25338), .Z(n25336) );
  NAND U33679 ( .A(o[585]), .B(n23579), .Z(n25338) );
  NANDN U33680 ( .A(n23580), .B(creg[585]), .Z(n25337) );
  NAND U33681 ( .A(n25339), .B(n18350), .Z(n13766) );
  NANDN U33682 ( .A(init), .B(m[586]), .Z(n18350) );
  AND U33683 ( .A(n25340), .B(n25341), .Z(n25339) );
  NAND U33684 ( .A(o[586]), .B(n23579), .Z(n25341) );
  NANDN U33685 ( .A(n23580), .B(creg[586]), .Z(n25340) );
  NAND U33686 ( .A(n25342), .B(n18348), .Z(n13765) );
  NANDN U33687 ( .A(init), .B(m[587]), .Z(n18348) );
  AND U33688 ( .A(n25343), .B(n25344), .Z(n25342) );
  NAND U33689 ( .A(o[587]), .B(n23579), .Z(n25344) );
  NANDN U33690 ( .A(n23580), .B(creg[587]), .Z(n25343) );
  NAND U33691 ( .A(n25345), .B(n18346), .Z(n13764) );
  NANDN U33692 ( .A(init), .B(m[588]), .Z(n18346) );
  AND U33693 ( .A(n25346), .B(n25347), .Z(n25345) );
  NAND U33694 ( .A(o[588]), .B(n23579), .Z(n25347) );
  NANDN U33695 ( .A(n23580), .B(creg[588]), .Z(n25346) );
  NAND U33696 ( .A(n25348), .B(n18344), .Z(n13763) );
  NANDN U33697 ( .A(init), .B(m[589]), .Z(n18344) );
  AND U33698 ( .A(n25349), .B(n25350), .Z(n25348) );
  NAND U33699 ( .A(o[589]), .B(n23579), .Z(n25350) );
  NANDN U33700 ( .A(n23580), .B(creg[589]), .Z(n25349) );
  NAND U33701 ( .A(n25351), .B(n18340), .Z(n13762) );
  NANDN U33702 ( .A(init), .B(m[590]), .Z(n18340) );
  AND U33703 ( .A(n25352), .B(n25353), .Z(n25351) );
  NAND U33704 ( .A(o[590]), .B(n23579), .Z(n25353) );
  NANDN U33705 ( .A(n23580), .B(creg[590]), .Z(n25352) );
  NAND U33706 ( .A(n25354), .B(n18338), .Z(n13761) );
  NANDN U33707 ( .A(init), .B(m[591]), .Z(n18338) );
  AND U33708 ( .A(n25355), .B(n25356), .Z(n25354) );
  NAND U33709 ( .A(o[591]), .B(n23579), .Z(n25356) );
  NANDN U33710 ( .A(n23580), .B(creg[591]), .Z(n25355) );
  NAND U33711 ( .A(n25357), .B(n18336), .Z(n13760) );
  NANDN U33712 ( .A(init), .B(m[592]), .Z(n18336) );
  AND U33713 ( .A(n25358), .B(n25359), .Z(n25357) );
  NAND U33714 ( .A(o[592]), .B(n23579), .Z(n25359) );
  NANDN U33715 ( .A(n23580), .B(creg[592]), .Z(n25358) );
  NAND U33716 ( .A(n25360), .B(n18334), .Z(n13759) );
  NANDN U33717 ( .A(init), .B(m[593]), .Z(n18334) );
  AND U33718 ( .A(n25361), .B(n25362), .Z(n25360) );
  NAND U33719 ( .A(o[593]), .B(n23579), .Z(n25362) );
  NANDN U33720 ( .A(n23580), .B(creg[593]), .Z(n25361) );
  NAND U33721 ( .A(n25363), .B(n18332), .Z(n13758) );
  NANDN U33722 ( .A(init), .B(m[594]), .Z(n18332) );
  AND U33723 ( .A(n25364), .B(n25365), .Z(n25363) );
  NAND U33724 ( .A(o[594]), .B(n23579), .Z(n25365) );
  NANDN U33725 ( .A(n23580), .B(creg[594]), .Z(n25364) );
  NAND U33726 ( .A(n25366), .B(n18330), .Z(n13757) );
  NANDN U33727 ( .A(init), .B(m[595]), .Z(n18330) );
  AND U33728 ( .A(n25367), .B(n25368), .Z(n25366) );
  NAND U33729 ( .A(o[595]), .B(n23579), .Z(n25368) );
  NANDN U33730 ( .A(n23580), .B(creg[595]), .Z(n25367) );
  NAND U33731 ( .A(n25369), .B(n18328), .Z(n13756) );
  NANDN U33732 ( .A(init), .B(m[596]), .Z(n18328) );
  AND U33733 ( .A(n25370), .B(n25371), .Z(n25369) );
  NAND U33734 ( .A(o[596]), .B(n23579), .Z(n25371) );
  NANDN U33735 ( .A(n23580), .B(creg[596]), .Z(n25370) );
  NAND U33736 ( .A(n25372), .B(n18326), .Z(n13755) );
  NANDN U33737 ( .A(init), .B(m[597]), .Z(n18326) );
  AND U33738 ( .A(n25373), .B(n25374), .Z(n25372) );
  NAND U33739 ( .A(o[597]), .B(n23579), .Z(n25374) );
  NANDN U33740 ( .A(n23580), .B(creg[597]), .Z(n25373) );
  NAND U33741 ( .A(n25375), .B(n18324), .Z(n13754) );
  NANDN U33742 ( .A(init), .B(m[598]), .Z(n18324) );
  AND U33743 ( .A(n25376), .B(n25377), .Z(n25375) );
  NAND U33744 ( .A(o[598]), .B(n23579), .Z(n25377) );
  NANDN U33745 ( .A(n23580), .B(creg[598]), .Z(n25376) );
  NAND U33746 ( .A(n25378), .B(n18322), .Z(n13753) );
  NANDN U33747 ( .A(init), .B(m[599]), .Z(n18322) );
  AND U33748 ( .A(n25379), .B(n25380), .Z(n25378) );
  NAND U33749 ( .A(o[599]), .B(n23579), .Z(n25380) );
  NANDN U33750 ( .A(n23580), .B(creg[599]), .Z(n25379) );
  NAND U33751 ( .A(n25381), .B(n18316), .Z(n13752) );
  NANDN U33752 ( .A(init), .B(m[600]), .Z(n18316) );
  AND U33753 ( .A(n25382), .B(n25383), .Z(n25381) );
  NAND U33754 ( .A(o[600]), .B(n23579), .Z(n25383) );
  NANDN U33755 ( .A(n23580), .B(creg[600]), .Z(n25382) );
  NAND U33756 ( .A(n25384), .B(n18314), .Z(n13751) );
  NANDN U33757 ( .A(init), .B(m[601]), .Z(n18314) );
  AND U33758 ( .A(n25385), .B(n25386), .Z(n25384) );
  NAND U33759 ( .A(o[601]), .B(n23579), .Z(n25386) );
  NANDN U33760 ( .A(n23580), .B(creg[601]), .Z(n25385) );
  NAND U33761 ( .A(n25387), .B(n18312), .Z(n13750) );
  NANDN U33762 ( .A(init), .B(m[602]), .Z(n18312) );
  AND U33763 ( .A(n25388), .B(n25389), .Z(n25387) );
  NAND U33764 ( .A(o[602]), .B(n23579), .Z(n25389) );
  NANDN U33765 ( .A(n23580), .B(creg[602]), .Z(n25388) );
  NAND U33766 ( .A(n25390), .B(n18310), .Z(n13749) );
  NANDN U33767 ( .A(init), .B(m[603]), .Z(n18310) );
  AND U33768 ( .A(n25391), .B(n25392), .Z(n25390) );
  NAND U33769 ( .A(o[603]), .B(n23579), .Z(n25392) );
  NANDN U33770 ( .A(n23580), .B(creg[603]), .Z(n25391) );
  NAND U33771 ( .A(n25393), .B(n18308), .Z(n13748) );
  NANDN U33772 ( .A(init), .B(m[604]), .Z(n18308) );
  AND U33773 ( .A(n25394), .B(n25395), .Z(n25393) );
  NAND U33774 ( .A(o[604]), .B(n23579), .Z(n25395) );
  NANDN U33775 ( .A(n23580), .B(creg[604]), .Z(n25394) );
  NAND U33776 ( .A(n25396), .B(n18306), .Z(n13747) );
  NANDN U33777 ( .A(init), .B(m[605]), .Z(n18306) );
  AND U33778 ( .A(n25397), .B(n25398), .Z(n25396) );
  NAND U33779 ( .A(o[605]), .B(n23579), .Z(n25398) );
  NANDN U33780 ( .A(n23580), .B(creg[605]), .Z(n25397) );
  NAND U33781 ( .A(n25399), .B(n18304), .Z(n13746) );
  NANDN U33782 ( .A(init), .B(m[606]), .Z(n18304) );
  AND U33783 ( .A(n25400), .B(n25401), .Z(n25399) );
  NAND U33784 ( .A(o[606]), .B(n23579), .Z(n25401) );
  NANDN U33785 ( .A(n23580), .B(creg[606]), .Z(n25400) );
  NAND U33786 ( .A(n25402), .B(n18302), .Z(n13745) );
  NANDN U33787 ( .A(init), .B(m[607]), .Z(n18302) );
  AND U33788 ( .A(n25403), .B(n25404), .Z(n25402) );
  NAND U33789 ( .A(o[607]), .B(n23579), .Z(n25404) );
  NANDN U33790 ( .A(n23580), .B(creg[607]), .Z(n25403) );
  NAND U33791 ( .A(n25405), .B(n18300), .Z(n13744) );
  NANDN U33792 ( .A(init), .B(m[608]), .Z(n18300) );
  AND U33793 ( .A(n25406), .B(n25407), .Z(n25405) );
  NAND U33794 ( .A(o[608]), .B(n23579), .Z(n25407) );
  NANDN U33795 ( .A(n23580), .B(creg[608]), .Z(n25406) );
  NAND U33796 ( .A(n25408), .B(n18298), .Z(n13743) );
  NANDN U33797 ( .A(init), .B(m[609]), .Z(n18298) );
  AND U33798 ( .A(n25409), .B(n25410), .Z(n25408) );
  NAND U33799 ( .A(o[609]), .B(n23579), .Z(n25410) );
  NANDN U33800 ( .A(n23580), .B(creg[609]), .Z(n25409) );
  NAND U33801 ( .A(n25411), .B(n18294), .Z(n13742) );
  NANDN U33802 ( .A(init), .B(m[610]), .Z(n18294) );
  AND U33803 ( .A(n25412), .B(n25413), .Z(n25411) );
  NAND U33804 ( .A(o[610]), .B(n23579), .Z(n25413) );
  NANDN U33805 ( .A(n23580), .B(creg[610]), .Z(n25412) );
  NAND U33806 ( .A(n25414), .B(n18292), .Z(n13741) );
  NANDN U33807 ( .A(init), .B(m[611]), .Z(n18292) );
  AND U33808 ( .A(n25415), .B(n25416), .Z(n25414) );
  NAND U33809 ( .A(o[611]), .B(n23579), .Z(n25416) );
  NANDN U33810 ( .A(n23580), .B(creg[611]), .Z(n25415) );
  NAND U33811 ( .A(n25417), .B(n18290), .Z(n13740) );
  NANDN U33812 ( .A(init), .B(m[612]), .Z(n18290) );
  AND U33813 ( .A(n25418), .B(n25419), .Z(n25417) );
  NAND U33814 ( .A(o[612]), .B(n23579), .Z(n25419) );
  NANDN U33815 ( .A(n23580), .B(creg[612]), .Z(n25418) );
  NAND U33816 ( .A(n25420), .B(n18288), .Z(n13739) );
  NANDN U33817 ( .A(init), .B(m[613]), .Z(n18288) );
  AND U33818 ( .A(n25421), .B(n25422), .Z(n25420) );
  NAND U33819 ( .A(o[613]), .B(n23579), .Z(n25422) );
  NANDN U33820 ( .A(n23580), .B(creg[613]), .Z(n25421) );
  NAND U33821 ( .A(n25423), .B(n18286), .Z(n13738) );
  NANDN U33822 ( .A(init), .B(m[614]), .Z(n18286) );
  AND U33823 ( .A(n25424), .B(n25425), .Z(n25423) );
  NAND U33824 ( .A(o[614]), .B(n23579), .Z(n25425) );
  NANDN U33825 ( .A(n23580), .B(creg[614]), .Z(n25424) );
  NAND U33826 ( .A(n25426), .B(n18284), .Z(n13737) );
  NANDN U33827 ( .A(init), .B(m[615]), .Z(n18284) );
  AND U33828 ( .A(n25427), .B(n25428), .Z(n25426) );
  NAND U33829 ( .A(o[615]), .B(n23579), .Z(n25428) );
  NANDN U33830 ( .A(n23580), .B(creg[615]), .Z(n25427) );
  NAND U33831 ( .A(n25429), .B(n18282), .Z(n13736) );
  NANDN U33832 ( .A(init), .B(m[616]), .Z(n18282) );
  AND U33833 ( .A(n25430), .B(n25431), .Z(n25429) );
  NAND U33834 ( .A(o[616]), .B(n23579), .Z(n25431) );
  NANDN U33835 ( .A(n23580), .B(creg[616]), .Z(n25430) );
  NAND U33836 ( .A(n25432), .B(n18280), .Z(n13735) );
  NANDN U33837 ( .A(init), .B(m[617]), .Z(n18280) );
  AND U33838 ( .A(n25433), .B(n25434), .Z(n25432) );
  NAND U33839 ( .A(o[617]), .B(n23579), .Z(n25434) );
  NANDN U33840 ( .A(n23580), .B(creg[617]), .Z(n25433) );
  NAND U33841 ( .A(n25435), .B(n18278), .Z(n13734) );
  NANDN U33842 ( .A(init), .B(m[618]), .Z(n18278) );
  AND U33843 ( .A(n25436), .B(n25437), .Z(n25435) );
  NAND U33844 ( .A(o[618]), .B(n23579), .Z(n25437) );
  NANDN U33845 ( .A(n23580), .B(creg[618]), .Z(n25436) );
  NAND U33846 ( .A(n25438), .B(n18276), .Z(n13733) );
  NANDN U33847 ( .A(init), .B(m[619]), .Z(n18276) );
  AND U33848 ( .A(n25439), .B(n25440), .Z(n25438) );
  NAND U33849 ( .A(o[619]), .B(n23579), .Z(n25440) );
  NANDN U33850 ( .A(n23580), .B(creg[619]), .Z(n25439) );
  NAND U33851 ( .A(n25441), .B(n18272), .Z(n13732) );
  NANDN U33852 ( .A(init), .B(m[620]), .Z(n18272) );
  AND U33853 ( .A(n25442), .B(n25443), .Z(n25441) );
  NAND U33854 ( .A(o[620]), .B(n23579), .Z(n25443) );
  NANDN U33855 ( .A(n23580), .B(creg[620]), .Z(n25442) );
  NAND U33856 ( .A(n25444), .B(n18270), .Z(n13731) );
  NANDN U33857 ( .A(init), .B(m[621]), .Z(n18270) );
  AND U33858 ( .A(n25445), .B(n25446), .Z(n25444) );
  NAND U33859 ( .A(o[621]), .B(n23579), .Z(n25446) );
  NANDN U33860 ( .A(n23580), .B(creg[621]), .Z(n25445) );
  NAND U33861 ( .A(n25447), .B(n18268), .Z(n13730) );
  NANDN U33862 ( .A(init), .B(m[622]), .Z(n18268) );
  AND U33863 ( .A(n25448), .B(n25449), .Z(n25447) );
  NAND U33864 ( .A(o[622]), .B(n23579), .Z(n25449) );
  NANDN U33865 ( .A(n23580), .B(creg[622]), .Z(n25448) );
  NAND U33866 ( .A(n25450), .B(n18266), .Z(n13729) );
  NANDN U33867 ( .A(init), .B(m[623]), .Z(n18266) );
  AND U33868 ( .A(n25451), .B(n25452), .Z(n25450) );
  NAND U33869 ( .A(o[623]), .B(n23579), .Z(n25452) );
  NANDN U33870 ( .A(n23580), .B(creg[623]), .Z(n25451) );
  NAND U33871 ( .A(n25453), .B(n18264), .Z(n13728) );
  NANDN U33872 ( .A(init), .B(m[624]), .Z(n18264) );
  AND U33873 ( .A(n25454), .B(n25455), .Z(n25453) );
  NAND U33874 ( .A(o[624]), .B(n23579), .Z(n25455) );
  NANDN U33875 ( .A(n23580), .B(creg[624]), .Z(n25454) );
  NAND U33876 ( .A(n25456), .B(n18262), .Z(n13727) );
  NANDN U33877 ( .A(init), .B(m[625]), .Z(n18262) );
  AND U33878 ( .A(n25457), .B(n25458), .Z(n25456) );
  NAND U33879 ( .A(o[625]), .B(n23579), .Z(n25458) );
  NANDN U33880 ( .A(n23580), .B(creg[625]), .Z(n25457) );
  NAND U33881 ( .A(n25459), .B(n18260), .Z(n13726) );
  NANDN U33882 ( .A(init), .B(m[626]), .Z(n18260) );
  AND U33883 ( .A(n25460), .B(n25461), .Z(n25459) );
  NAND U33884 ( .A(o[626]), .B(n23579), .Z(n25461) );
  NANDN U33885 ( .A(n23580), .B(creg[626]), .Z(n25460) );
  NAND U33886 ( .A(n25462), .B(n18258), .Z(n13725) );
  NANDN U33887 ( .A(init), .B(m[627]), .Z(n18258) );
  AND U33888 ( .A(n25463), .B(n25464), .Z(n25462) );
  NAND U33889 ( .A(o[627]), .B(n23579), .Z(n25464) );
  NANDN U33890 ( .A(n23580), .B(creg[627]), .Z(n25463) );
  NAND U33891 ( .A(n25465), .B(n18256), .Z(n13724) );
  NANDN U33892 ( .A(init), .B(m[628]), .Z(n18256) );
  AND U33893 ( .A(n25466), .B(n25467), .Z(n25465) );
  NAND U33894 ( .A(o[628]), .B(n23579), .Z(n25467) );
  NANDN U33895 ( .A(n23580), .B(creg[628]), .Z(n25466) );
  NAND U33896 ( .A(n25468), .B(n18254), .Z(n13723) );
  NANDN U33897 ( .A(init), .B(m[629]), .Z(n18254) );
  AND U33898 ( .A(n25469), .B(n25470), .Z(n25468) );
  NAND U33899 ( .A(o[629]), .B(n23579), .Z(n25470) );
  NANDN U33900 ( .A(n23580), .B(creg[629]), .Z(n25469) );
  NAND U33901 ( .A(n25471), .B(n18250), .Z(n13722) );
  NANDN U33902 ( .A(init), .B(m[630]), .Z(n18250) );
  AND U33903 ( .A(n25472), .B(n25473), .Z(n25471) );
  NAND U33904 ( .A(o[630]), .B(n23579), .Z(n25473) );
  NANDN U33905 ( .A(n23580), .B(creg[630]), .Z(n25472) );
  NAND U33906 ( .A(n25474), .B(n18248), .Z(n13721) );
  NANDN U33907 ( .A(init), .B(m[631]), .Z(n18248) );
  AND U33908 ( .A(n25475), .B(n25476), .Z(n25474) );
  NAND U33909 ( .A(o[631]), .B(n23579), .Z(n25476) );
  NANDN U33910 ( .A(n23580), .B(creg[631]), .Z(n25475) );
  NAND U33911 ( .A(n25477), .B(n18246), .Z(n13720) );
  NANDN U33912 ( .A(init), .B(m[632]), .Z(n18246) );
  AND U33913 ( .A(n25478), .B(n25479), .Z(n25477) );
  NAND U33914 ( .A(o[632]), .B(n23579), .Z(n25479) );
  NANDN U33915 ( .A(n23580), .B(creg[632]), .Z(n25478) );
  NAND U33916 ( .A(n25480), .B(n18244), .Z(n13719) );
  NANDN U33917 ( .A(init), .B(m[633]), .Z(n18244) );
  AND U33918 ( .A(n25481), .B(n25482), .Z(n25480) );
  NAND U33919 ( .A(o[633]), .B(n23579), .Z(n25482) );
  NANDN U33920 ( .A(n23580), .B(creg[633]), .Z(n25481) );
  NAND U33921 ( .A(n25483), .B(n18242), .Z(n13718) );
  NANDN U33922 ( .A(init), .B(m[634]), .Z(n18242) );
  AND U33923 ( .A(n25484), .B(n25485), .Z(n25483) );
  NAND U33924 ( .A(o[634]), .B(n23579), .Z(n25485) );
  NANDN U33925 ( .A(n23580), .B(creg[634]), .Z(n25484) );
  NAND U33926 ( .A(n25486), .B(n18240), .Z(n13717) );
  NANDN U33927 ( .A(init), .B(m[635]), .Z(n18240) );
  AND U33928 ( .A(n25487), .B(n25488), .Z(n25486) );
  NAND U33929 ( .A(o[635]), .B(n23579), .Z(n25488) );
  NANDN U33930 ( .A(n23580), .B(creg[635]), .Z(n25487) );
  NAND U33931 ( .A(n25489), .B(n18238), .Z(n13716) );
  NANDN U33932 ( .A(init), .B(m[636]), .Z(n18238) );
  AND U33933 ( .A(n25490), .B(n25491), .Z(n25489) );
  NAND U33934 ( .A(o[636]), .B(n23579), .Z(n25491) );
  NANDN U33935 ( .A(n23580), .B(creg[636]), .Z(n25490) );
  NAND U33936 ( .A(n25492), .B(n18236), .Z(n13715) );
  NANDN U33937 ( .A(init), .B(m[637]), .Z(n18236) );
  AND U33938 ( .A(n25493), .B(n25494), .Z(n25492) );
  NAND U33939 ( .A(o[637]), .B(n23579), .Z(n25494) );
  NANDN U33940 ( .A(n23580), .B(creg[637]), .Z(n25493) );
  NAND U33941 ( .A(n25495), .B(n18234), .Z(n13714) );
  NANDN U33942 ( .A(init), .B(m[638]), .Z(n18234) );
  AND U33943 ( .A(n25496), .B(n25497), .Z(n25495) );
  NAND U33944 ( .A(o[638]), .B(n23579), .Z(n25497) );
  NANDN U33945 ( .A(n23580), .B(creg[638]), .Z(n25496) );
  NAND U33946 ( .A(n25498), .B(n18232), .Z(n13713) );
  NANDN U33947 ( .A(init), .B(m[639]), .Z(n18232) );
  AND U33948 ( .A(n25499), .B(n25500), .Z(n25498) );
  NAND U33949 ( .A(o[639]), .B(n23579), .Z(n25500) );
  NANDN U33950 ( .A(n23580), .B(creg[639]), .Z(n25499) );
  NAND U33951 ( .A(n25501), .B(n18228), .Z(n13712) );
  NANDN U33952 ( .A(init), .B(m[640]), .Z(n18228) );
  AND U33953 ( .A(n25502), .B(n25503), .Z(n25501) );
  NAND U33954 ( .A(o[640]), .B(n23579), .Z(n25503) );
  NANDN U33955 ( .A(n23580), .B(creg[640]), .Z(n25502) );
  NAND U33956 ( .A(n25504), .B(n18226), .Z(n13711) );
  NANDN U33957 ( .A(init), .B(m[641]), .Z(n18226) );
  AND U33958 ( .A(n25505), .B(n25506), .Z(n25504) );
  NAND U33959 ( .A(o[641]), .B(n23579), .Z(n25506) );
  NANDN U33960 ( .A(n23580), .B(creg[641]), .Z(n25505) );
  NAND U33961 ( .A(n25507), .B(n18224), .Z(n13710) );
  NANDN U33962 ( .A(init), .B(m[642]), .Z(n18224) );
  AND U33963 ( .A(n25508), .B(n25509), .Z(n25507) );
  NAND U33964 ( .A(o[642]), .B(n23579), .Z(n25509) );
  NANDN U33965 ( .A(n23580), .B(creg[642]), .Z(n25508) );
  NAND U33966 ( .A(n25510), .B(n18222), .Z(n13709) );
  NANDN U33967 ( .A(init), .B(m[643]), .Z(n18222) );
  AND U33968 ( .A(n25511), .B(n25512), .Z(n25510) );
  NAND U33969 ( .A(o[643]), .B(n23579), .Z(n25512) );
  NANDN U33970 ( .A(n23580), .B(creg[643]), .Z(n25511) );
  NAND U33971 ( .A(n25513), .B(n18220), .Z(n13708) );
  NANDN U33972 ( .A(init), .B(m[644]), .Z(n18220) );
  AND U33973 ( .A(n25514), .B(n25515), .Z(n25513) );
  NAND U33974 ( .A(o[644]), .B(n23579), .Z(n25515) );
  NANDN U33975 ( .A(n23580), .B(creg[644]), .Z(n25514) );
  NAND U33976 ( .A(n25516), .B(n18218), .Z(n13707) );
  NANDN U33977 ( .A(init), .B(m[645]), .Z(n18218) );
  AND U33978 ( .A(n25517), .B(n25518), .Z(n25516) );
  NAND U33979 ( .A(o[645]), .B(n23579), .Z(n25518) );
  NANDN U33980 ( .A(n23580), .B(creg[645]), .Z(n25517) );
  NAND U33981 ( .A(n25519), .B(n18216), .Z(n13706) );
  NANDN U33982 ( .A(init), .B(m[646]), .Z(n18216) );
  AND U33983 ( .A(n25520), .B(n25521), .Z(n25519) );
  NAND U33984 ( .A(o[646]), .B(n23579), .Z(n25521) );
  NANDN U33985 ( .A(n23580), .B(creg[646]), .Z(n25520) );
  NAND U33986 ( .A(n25522), .B(n18214), .Z(n13705) );
  NANDN U33987 ( .A(init), .B(m[647]), .Z(n18214) );
  AND U33988 ( .A(n25523), .B(n25524), .Z(n25522) );
  NAND U33989 ( .A(o[647]), .B(n23579), .Z(n25524) );
  NANDN U33990 ( .A(n23580), .B(creg[647]), .Z(n25523) );
  NAND U33991 ( .A(n25525), .B(n18212), .Z(n13704) );
  NANDN U33992 ( .A(init), .B(m[648]), .Z(n18212) );
  AND U33993 ( .A(n25526), .B(n25527), .Z(n25525) );
  NAND U33994 ( .A(o[648]), .B(n23579), .Z(n25527) );
  NANDN U33995 ( .A(n23580), .B(creg[648]), .Z(n25526) );
  NAND U33996 ( .A(n25528), .B(n18210), .Z(n13703) );
  NANDN U33997 ( .A(init), .B(m[649]), .Z(n18210) );
  AND U33998 ( .A(n25529), .B(n25530), .Z(n25528) );
  NAND U33999 ( .A(o[649]), .B(n23579), .Z(n25530) );
  NANDN U34000 ( .A(n23580), .B(creg[649]), .Z(n25529) );
  NAND U34001 ( .A(n25531), .B(n18206), .Z(n13702) );
  NANDN U34002 ( .A(init), .B(m[650]), .Z(n18206) );
  AND U34003 ( .A(n25532), .B(n25533), .Z(n25531) );
  NAND U34004 ( .A(o[650]), .B(n23579), .Z(n25533) );
  NANDN U34005 ( .A(n23580), .B(creg[650]), .Z(n25532) );
  NAND U34006 ( .A(n25534), .B(n18204), .Z(n13701) );
  NANDN U34007 ( .A(init), .B(m[651]), .Z(n18204) );
  AND U34008 ( .A(n25535), .B(n25536), .Z(n25534) );
  NAND U34009 ( .A(o[651]), .B(n23579), .Z(n25536) );
  NANDN U34010 ( .A(n23580), .B(creg[651]), .Z(n25535) );
  NAND U34011 ( .A(n25537), .B(n18202), .Z(n13700) );
  NANDN U34012 ( .A(init), .B(m[652]), .Z(n18202) );
  AND U34013 ( .A(n25538), .B(n25539), .Z(n25537) );
  NAND U34014 ( .A(o[652]), .B(n23579), .Z(n25539) );
  NANDN U34015 ( .A(n23580), .B(creg[652]), .Z(n25538) );
  NAND U34016 ( .A(n25540), .B(n18200), .Z(n13699) );
  NANDN U34017 ( .A(init), .B(m[653]), .Z(n18200) );
  AND U34018 ( .A(n25541), .B(n25542), .Z(n25540) );
  NAND U34019 ( .A(o[653]), .B(n23579), .Z(n25542) );
  NANDN U34020 ( .A(n23580), .B(creg[653]), .Z(n25541) );
  NAND U34021 ( .A(n25543), .B(n18198), .Z(n13698) );
  NANDN U34022 ( .A(init), .B(m[654]), .Z(n18198) );
  AND U34023 ( .A(n25544), .B(n25545), .Z(n25543) );
  NAND U34024 ( .A(o[654]), .B(n23579), .Z(n25545) );
  NANDN U34025 ( .A(n23580), .B(creg[654]), .Z(n25544) );
  NAND U34026 ( .A(n25546), .B(n18196), .Z(n13697) );
  NANDN U34027 ( .A(init), .B(m[655]), .Z(n18196) );
  AND U34028 ( .A(n25547), .B(n25548), .Z(n25546) );
  NAND U34029 ( .A(o[655]), .B(n23579), .Z(n25548) );
  NANDN U34030 ( .A(n23580), .B(creg[655]), .Z(n25547) );
  NAND U34031 ( .A(n25549), .B(n18194), .Z(n13696) );
  NANDN U34032 ( .A(init), .B(m[656]), .Z(n18194) );
  AND U34033 ( .A(n25550), .B(n25551), .Z(n25549) );
  NAND U34034 ( .A(o[656]), .B(n23579), .Z(n25551) );
  NANDN U34035 ( .A(n23580), .B(creg[656]), .Z(n25550) );
  NAND U34036 ( .A(n25552), .B(n18192), .Z(n13695) );
  NANDN U34037 ( .A(init), .B(m[657]), .Z(n18192) );
  AND U34038 ( .A(n25553), .B(n25554), .Z(n25552) );
  NAND U34039 ( .A(o[657]), .B(n23579), .Z(n25554) );
  NANDN U34040 ( .A(n23580), .B(creg[657]), .Z(n25553) );
  NAND U34041 ( .A(n25555), .B(n18190), .Z(n13694) );
  NANDN U34042 ( .A(init), .B(m[658]), .Z(n18190) );
  AND U34043 ( .A(n25556), .B(n25557), .Z(n25555) );
  NAND U34044 ( .A(o[658]), .B(n23579), .Z(n25557) );
  NANDN U34045 ( .A(n23580), .B(creg[658]), .Z(n25556) );
  NAND U34046 ( .A(n25558), .B(n18188), .Z(n13693) );
  NANDN U34047 ( .A(init), .B(m[659]), .Z(n18188) );
  AND U34048 ( .A(n25559), .B(n25560), .Z(n25558) );
  NAND U34049 ( .A(o[659]), .B(n23579), .Z(n25560) );
  NANDN U34050 ( .A(n23580), .B(creg[659]), .Z(n25559) );
  NAND U34051 ( .A(n25561), .B(n18184), .Z(n13692) );
  NANDN U34052 ( .A(init), .B(m[660]), .Z(n18184) );
  AND U34053 ( .A(n25562), .B(n25563), .Z(n25561) );
  NAND U34054 ( .A(o[660]), .B(n23579), .Z(n25563) );
  NANDN U34055 ( .A(n23580), .B(creg[660]), .Z(n25562) );
  NAND U34056 ( .A(n25564), .B(n18182), .Z(n13691) );
  NANDN U34057 ( .A(init), .B(m[661]), .Z(n18182) );
  AND U34058 ( .A(n25565), .B(n25566), .Z(n25564) );
  NAND U34059 ( .A(o[661]), .B(n23579), .Z(n25566) );
  NANDN U34060 ( .A(n23580), .B(creg[661]), .Z(n25565) );
  NAND U34061 ( .A(n25567), .B(n18180), .Z(n13690) );
  NANDN U34062 ( .A(init), .B(m[662]), .Z(n18180) );
  AND U34063 ( .A(n25568), .B(n25569), .Z(n25567) );
  NAND U34064 ( .A(o[662]), .B(n23579), .Z(n25569) );
  NANDN U34065 ( .A(n23580), .B(creg[662]), .Z(n25568) );
  NAND U34066 ( .A(n25570), .B(n18178), .Z(n13689) );
  NANDN U34067 ( .A(init), .B(m[663]), .Z(n18178) );
  AND U34068 ( .A(n25571), .B(n25572), .Z(n25570) );
  NAND U34069 ( .A(o[663]), .B(n23579), .Z(n25572) );
  NANDN U34070 ( .A(n23580), .B(creg[663]), .Z(n25571) );
  NAND U34071 ( .A(n25573), .B(n18176), .Z(n13688) );
  NANDN U34072 ( .A(init), .B(m[664]), .Z(n18176) );
  AND U34073 ( .A(n25574), .B(n25575), .Z(n25573) );
  NAND U34074 ( .A(o[664]), .B(n23579), .Z(n25575) );
  NANDN U34075 ( .A(n23580), .B(creg[664]), .Z(n25574) );
  NAND U34076 ( .A(n25576), .B(n18174), .Z(n13687) );
  NANDN U34077 ( .A(init), .B(m[665]), .Z(n18174) );
  AND U34078 ( .A(n25577), .B(n25578), .Z(n25576) );
  NAND U34079 ( .A(o[665]), .B(n23579), .Z(n25578) );
  NANDN U34080 ( .A(n23580), .B(creg[665]), .Z(n25577) );
  NAND U34081 ( .A(n25579), .B(n18172), .Z(n13686) );
  NANDN U34082 ( .A(init), .B(m[666]), .Z(n18172) );
  AND U34083 ( .A(n25580), .B(n25581), .Z(n25579) );
  NAND U34084 ( .A(o[666]), .B(n23579), .Z(n25581) );
  NANDN U34085 ( .A(n23580), .B(creg[666]), .Z(n25580) );
  NAND U34086 ( .A(n25582), .B(n18170), .Z(n13685) );
  NANDN U34087 ( .A(init), .B(m[667]), .Z(n18170) );
  AND U34088 ( .A(n25583), .B(n25584), .Z(n25582) );
  NAND U34089 ( .A(o[667]), .B(n23579), .Z(n25584) );
  NANDN U34090 ( .A(n23580), .B(creg[667]), .Z(n25583) );
  NAND U34091 ( .A(n25585), .B(n18168), .Z(n13684) );
  NANDN U34092 ( .A(init), .B(m[668]), .Z(n18168) );
  AND U34093 ( .A(n25586), .B(n25587), .Z(n25585) );
  NAND U34094 ( .A(o[668]), .B(n23579), .Z(n25587) );
  NANDN U34095 ( .A(n23580), .B(creg[668]), .Z(n25586) );
  NAND U34096 ( .A(n25588), .B(n18166), .Z(n13683) );
  NANDN U34097 ( .A(init), .B(m[669]), .Z(n18166) );
  AND U34098 ( .A(n25589), .B(n25590), .Z(n25588) );
  NAND U34099 ( .A(o[669]), .B(n23579), .Z(n25590) );
  NANDN U34100 ( .A(n23580), .B(creg[669]), .Z(n25589) );
  NAND U34101 ( .A(n25591), .B(n18162), .Z(n13682) );
  NANDN U34102 ( .A(init), .B(m[670]), .Z(n18162) );
  AND U34103 ( .A(n25592), .B(n25593), .Z(n25591) );
  NAND U34104 ( .A(o[670]), .B(n23579), .Z(n25593) );
  NANDN U34105 ( .A(n23580), .B(creg[670]), .Z(n25592) );
  NAND U34106 ( .A(n25594), .B(n18160), .Z(n13681) );
  NANDN U34107 ( .A(init), .B(m[671]), .Z(n18160) );
  AND U34108 ( .A(n25595), .B(n25596), .Z(n25594) );
  NAND U34109 ( .A(o[671]), .B(n23579), .Z(n25596) );
  NANDN U34110 ( .A(n23580), .B(creg[671]), .Z(n25595) );
  NAND U34111 ( .A(n25597), .B(n18158), .Z(n13680) );
  NANDN U34112 ( .A(init), .B(m[672]), .Z(n18158) );
  AND U34113 ( .A(n25598), .B(n25599), .Z(n25597) );
  NAND U34114 ( .A(o[672]), .B(n23579), .Z(n25599) );
  NANDN U34115 ( .A(n23580), .B(creg[672]), .Z(n25598) );
  NAND U34116 ( .A(n25600), .B(n18156), .Z(n13679) );
  NANDN U34117 ( .A(init), .B(m[673]), .Z(n18156) );
  AND U34118 ( .A(n25601), .B(n25602), .Z(n25600) );
  NAND U34119 ( .A(o[673]), .B(n23579), .Z(n25602) );
  NANDN U34120 ( .A(n23580), .B(creg[673]), .Z(n25601) );
  NAND U34121 ( .A(n25603), .B(n18154), .Z(n13678) );
  NANDN U34122 ( .A(init), .B(m[674]), .Z(n18154) );
  AND U34123 ( .A(n25604), .B(n25605), .Z(n25603) );
  NAND U34124 ( .A(o[674]), .B(n23579), .Z(n25605) );
  NANDN U34125 ( .A(n23580), .B(creg[674]), .Z(n25604) );
  NAND U34126 ( .A(n25606), .B(n18152), .Z(n13677) );
  NANDN U34127 ( .A(init), .B(m[675]), .Z(n18152) );
  AND U34128 ( .A(n25607), .B(n25608), .Z(n25606) );
  NAND U34129 ( .A(o[675]), .B(n23579), .Z(n25608) );
  NANDN U34130 ( .A(n23580), .B(creg[675]), .Z(n25607) );
  NAND U34131 ( .A(n25609), .B(n18150), .Z(n13676) );
  NANDN U34132 ( .A(init), .B(m[676]), .Z(n18150) );
  AND U34133 ( .A(n25610), .B(n25611), .Z(n25609) );
  NAND U34134 ( .A(o[676]), .B(n23579), .Z(n25611) );
  NANDN U34135 ( .A(n23580), .B(creg[676]), .Z(n25610) );
  NAND U34136 ( .A(n25612), .B(n18148), .Z(n13675) );
  NANDN U34137 ( .A(init), .B(m[677]), .Z(n18148) );
  AND U34138 ( .A(n25613), .B(n25614), .Z(n25612) );
  NAND U34139 ( .A(o[677]), .B(n23579), .Z(n25614) );
  NANDN U34140 ( .A(n23580), .B(creg[677]), .Z(n25613) );
  NAND U34141 ( .A(n25615), .B(n18146), .Z(n13674) );
  NANDN U34142 ( .A(init), .B(m[678]), .Z(n18146) );
  AND U34143 ( .A(n25616), .B(n25617), .Z(n25615) );
  NAND U34144 ( .A(o[678]), .B(n23579), .Z(n25617) );
  NANDN U34145 ( .A(n23580), .B(creg[678]), .Z(n25616) );
  NAND U34146 ( .A(n25618), .B(n18144), .Z(n13673) );
  NANDN U34147 ( .A(init), .B(m[679]), .Z(n18144) );
  AND U34148 ( .A(n25619), .B(n25620), .Z(n25618) );
  NAND U34149 ( .A(o[679]), .B(n23579), .Z(n25620) );
  NANDN U34150 ( .A(n23580), .B(creg[679]), .Z(n25619) );
  NAND U34151 ( .A(n25621), .B(n18140), .Z(n13672) );
  NANDN U34152 ( .A(init), .B(m[680]), .Z(n18140) );
  AND U34153 ( .A(n25622), .B(n25623), .Z(n25621) );
  NAND U34154 ( .A(o[680]), .B(n23579), .Z(n25623) );
  NANDN U34155 ( .A(n23580), .B(creg[680]), .Z(n25622) );
  NAND U34156 ( .A(n25624), .B(n18138), .Z(n13671) );
  NANDN U34157 ( .A(init), .B(m[681]), .Z(n18138) );
  AND U34158 ( .A(n25625), .B(n25626), .Z(n25624) );
  NAND U34159 ( .A(o[681]), .B(n23579), .Z(n25626) );
  NANDN U34160 ( .A(n23580), .B(creg[681]), .Z(n25625) );
  NAND U34161 ( .A(n25627), .B(n18136), .Z(n13670) );
  NANDN U34162 ( .A(init), .B(m[682]), .Z(n18136) );
  AND U34163 ( .A(n25628), .B(n25629), .Z(n25627) );
  NAND U34164 ( .A(o[682]), .B(n23579), .Z(n25629) );
  NANDN U34165 ( .A(n23580), .B(creg[682]), .Z(n25628) );
  NAND U34166 ( .A(n25630), .B(n18134), .Z(n13669) );
  NANDN U34167 ( .A(init), .B(m[683]), .Z(n18134) );
  AND U34168 ( .A(n25631), .B(n25632), .Z(n25630) );
  NAND U34169 ( .A(o[683]), .B(n23579), .Z(n25632) );
  NANDN U34170 ( .A(n23580), .B(creg[683]), .Z(n25631) );
  NAND U34171 ( .A(n25633), .B(n18132), .Z(n13668) );
  NANDN U34172 ( .A(init), .B(m[684]), .Z(n18132) );
  AND U34173 ( .A(n25634), .B(n25635), .Z(n25633) );
  NAND U34174 ( .A(o[684]), .B(n23579), .Z(n25635) );
  NANDN U34175 ( .A(n23580), .B(creg[684]), .Z(n25634) );
  NAND U34176 ( .A(n25636), .B(n18130), .Z(n13667) );
  NANDN U34177 ( .A(init), .B(m[685]), .Z(n18130) );
  AND U34178 ( .A(n25637), .B(n25638), .Z(n25636) );
  NAND U34179 ( .A(o[685]), .B(n23579), .Z(n25638) );
  NANDN U34180 ( .A(n23580), .B(creg[685]), .Z(n25637) );
  NAND U34181 ( .A(n25639), .B(n18128), .Z(n13666) );
  NANDN U34182 ( .A(init), .B(m[686]), .Z(n18128) );
  AND U34183 ( .A(n25640), .B(n25641), .Z(n25639) );
  NAND U34184 ( .A(o[686]), .B(n23579), .Z(n25641) );
  NANDN U34185 ( .A(n23580), .B(creg[686]), .Z(n25640) );
  NAND U34186 ( .A(n25642), .B(n18126), .Z(n13665) );
  NANDN U34187 ( .A(init), .B(m[687]), .Z(n18126) );
  AND U34188 ( .A(n25643), .B(n25644), .Z(n25642) );
  NAND U34189 ( .A(o[687]), .B(n23579), .Z(n25644) );
  NANDN U34190 ( .A(n23580), .B(creg[687]), .Z(n25643) );
  NAND U34191 ( .A(n25645), .B(n18124), .Z(n13664) );
  NANDN U34192 ( .A(init), .B(m[688]), .Z(n18124) );
  AND U34193 ( .A(n25646), .B(n25647), .Z(n25645) );
  NAND U34194 ( .A(o[688]), .B(n23579), .Z(n25647) );
  NANDN U34195 ( .A(n23580), .B(creg[688]), .Z(n25646) );
  NAND U34196 ( .A(n25648), .B(n18122), .Z(n13663) );
  NANDN U34197 ( .A(init), .B(m[689]), .Z(n18122) );
  AND U34198 ( .A(n25649), .B(n25650), .Z(n25648) );
  NAND U34199 ( .A(o[689]), .B(n23579), .Z(n25650) );
  NANDN U34200 ( .A(n23580), .B(creg[689]), .Z(n25649) );
  NAND U34201 ( .A(n25651), .B(n18118), .Z(n13662) );
  NANDN U34202 ( .A(init), .B(m[690]), .Z(n18118) );
  AND U34203 ( .A(n25652), .B(n25653), .Z(n25651) );
  NAND U34204 ( .A(o[690]), .B(n23579), .Z(n25653) );
  NANDN U34205 ( .A(n23580), .B(creg[690]), .Z(n25652) );
  NAND U34206 ( .A(n25654), .B(n18116), .Z(n13661) );
  NANDN U34207 ( .A(init), .B(m[691]), .Z(n18116) );
  AND U34208 ( .A(n25655), .B(n25656), .Z(n25654) );
  NAND U34209 ( .A(o[691]), .B(n23579), .Z(n25656) );
  NANDN U34210 ( .A(n23580), .B(creg[691]), .Z(n25655) );
  NAND U34211 ( .A(n25657), .B(n18114), .Z(n13660) );
  NANDN U34212 ( .A(init), .B(m[692]), .Z(n18114) );
  AND U34213 ( .A(n25658), .B(n25659), .Z(n25657) );
  NAND U34214 ( .A(o[692]), .B(n23579), .Z(n25659) );
  NANDN U34215 ( .A(n23580), .B(creg[692]), .Z(n25658) );
  NAND U34216 ( .A(n25660), .B(n18112), .Z(n13659) );
  NANDN U34217 ( .A(init), .B(m[693]), .Z(n18112) );
  AND U34218 ( .A(n25661), .B(n25662), .Z(n25660) );
  NAND U34219 ( .A(o[693]), .B(n23579), .Z(n25662) );
  NANDN U34220 ( .A(n23580), .B(creg[693]), .Z(n25661) );
  NAND U34221 ( .A(n25663), .B(n18110), .Z(n13658) );
  NANDN U34222 ( .A(init), .B(m[694]), .Z(n18110) );
  AND U34223 ( .A(n25664), .B(n25665), .Z(n25663) );
  NAND U34224 ( .A(o[694]), .B(n23579), .Z(n25665) );
  NANDN U34225 ( .A(n23580), .B(creg[694]), .Z(n25664) );
  NAND U34226 ( .A(n25666), .B(n18108), .Z(n13657) );
  NANDN U34227 ( .A(init), .B(m[695]), .Z(n18108) );
  AND U34228 ( .A(n25667), .B(n25668), .Z(n25666) );
  NAND U34229 ( .A(o[695]), .B(n23579), .Z(n25668) );
  NANDN U34230 ( .A(n23580), .B(creg[695]), .Z(n25667) );
  NAND U34231 ( .A(n25669), .B(n18106), .Z(n13656) );
  NANDN U34232 ( .A(init), .B(m[696]), .Z(n18106) );
  AND U34233 ( .A(n25670), .B(n25671), .Z(n25669) );
  NAND U34234 ( .A(o[696]), .B(n23579), .Z(n25671) );
  NANDN U34235 ( .A(n23580), .B(creg[696]), .Z(n25670) );
  NAND U34236 ( .A(n25672), .B(n18104), .Z(n13655) );
  NANDN U34237 ( .A(init), .B(m[697]), .Z(n18104) );
  AND U34238 ( .A(n25673), .B(n25674), .Z(n25672) );
  NAND U34239 ( .A(o[697]), .B(n23579), .Z(n25674) );
  NANDN U34240 ( .A(n23580), .B(creg[697]), .Z(n25673) );
  NAND U34241 ( .A(n25675), .B(n18102), .Z(n13654) );
  NANDN U34242 ( .A(init), .B(m[698]), .Z(n18102) );
  AND U34243 ( .A(n25676), .B(n25677), .Z(n25675) );
  NAND U34244 ( .A(o[698]), .B(n23579), .Z(n25677) );
  NANDN U34245 ( .A(n23580), .B(creg[698]), .Z(n25676) );
  NAND U34246 ( .A(n25678), .B(n18100), .Z(n13653) );
  NANDN U34247 ( .A(init), .B(m[699]), .Z(n18100) );
  AND U34248 ( .A(n25679), .B(n25680), .Z(n25678) );
  NAND U34249 ( .A(o[699]), .B(n23579), .Z(n25680) );
  NANDN U34250 ( .A(n23580), .B(creg[699]), .Z(n25679) );
  NAND U34251 ( .A(n25681), .B(n18094), .Z(n13652) );
  NANDN U34252 ( .A(init), .B(m[700]), .Z(n18094) );
  AND U34253 ( .A(n25682), .B(n25683), .Z(n25681) );
  NAND U34254 ( .A(o[700]), .B(n23579), .Z(n25683) );
  NANDN U34255 ( .A(n23580), .B(creg[700]), .Z(n25682) );
  NAND U34256 ( .A(n25684), .B(n18092), .Z(n13651) );
  NANDN U34257 ( .A(init), .B(m[701]), .Z(n18092) );
  AND U34258 ( .A(n25685), .B(n25686), .Z(n25684) );
  NAND U34259 ( .A(o[701]), .B(n23579), .Z(n25686) );
  NANDN U34260 ( .A(n23580), .B(creg[701]), .Z(n25685) );
  NAND U34261 ( .A(n25687), .B(n18090), .Z(n13650) );
  NANDN U34262 ( .A(init), .B(m[702]), .Z(n18090) );
  AND U34263 ( .A(n25688), .B(n25689), .Z(n25687) );
  NAND U34264 ( .A(o[702]), .B(n23579), .Z(n25689) );
  NANDN U34265 ( .A(n23580), .B(creg[702]), .Z(n25688) );
  NAND U34266 ( .A(n25690), .B(n18088), .Z(n13649) );
  NANDN U34267 ( .A(init), .B(m[703]), .Z(n18088) );
  AND U34268 ( .A(n25691), .B(n25692), .Z(n25690) );
  NAND U34269 ( .A(o[703]), .B(n23579), .Z(n25692) );
  NANDN U34270 ( .A(n23580), .B(creg[703]), .Z(n25691) );
  NAND U34271 ( .A(n25693), .B(n18086), .Z(n13648) );
  NANDN U34272 ( .A(init), .B(m[704]), .Z(n18086) );
  AND U34273 ( .A(n25694), .B(n25695), .Z(n25693) );
  NAND U34274 ( .A(o[704]), .B(n23579), .Z(n25695) );
  NANDN U34275 ( .A(n23580), .B(creg[704]), .Z(n25694) );
  NAND U34276 ( .A(n25696), .B(n18084), .Z(n13647) );
  NANDN U34277 ( .A(init), .B(m[705]), .Z(n18084) );
  AND U34278 ( .A(n25697), .B(n25698), .Z(n25696) );
  NAND U34279 ( .A(o[705]), .B(n23579), .Z(n25698) );
  NANDN U34280 ( .A(n23580), .B(creg[705]), .Z(n25697) );
  NAND U34281 ( .A(n25699), .B(n18082), .Z(n13646) );
  NANDN U34282 ( .A(init), .B(m[706]), .Z(n18082) );
  AND U34283 ( .A(n25700), .B(n25701), .Z(n25699) );
  NAND U34284 ( .A(o[706]), .B(n23579), .Z(n25701) );
  NANDN U34285 ( .A(n23580), .B(creg[706]), .Z(n25700) );
  NAND U34286 ( .A(n25702), .B(n18080), .Z(n13645) );
  NANDN U34287 ( .A(init), .B(m[707]), .Z(n18080) );
  AND U34288 ( .A(n25703), .B(n25704), .Z(n25702) );
  NAND U34289 ( .A(o[707]), .B(n23579), .Z(n25704) );
  NANDN U34290 ( .A(n23580), .B(creg[707]), .Z(n25703) );
  NAND U34291 ( .A(n25705), .B(n18078), .Z(n13644) );
  NANDN U34292 ( .A(init), .B(m[708]), .Z(n18078) );
  AND U34293 ( .A(n25706), .B(n25707), .Z(n25705) );
  NAND U34294 ( .A(o[708]), .B(n23579), .Z(n25707) );
  NANDN U34295 ( .A(n23580), .B(creg[708]), .Z(n25706) );
  NAND U34296 ( .A(n25708), .B(n18076), .Z(n13643) );
  NANDN U34297 ( .A(init), .B(m[709]), .Z(n18076) );
  AND U34298 ( .A(n25709), .B(n25710), .Z(n25708) );
  NAND U34299 ( .A(o[709]), .B(n23579), .Z(n25710) );
  NANDN U34300 ( .A(n23580), .B(creg[709]), .Z(n25709) );
  NAND U34301 ( .A(n25711), .B(n18072), .Z(n13642) );
  NANDN U34302 ( .A(init), .B(m[710]), .Z(n18072) );
  AND U34303 ( .A(n25712), .B(n25713), .Z(n25711) );
  NAND U34304 ( .A(o[710]), .B(n23579), .Z(n25713) );
  NANDN U34305 ( .A(n23580), .B(creg[710]), .Z(n25712) );
  NAND U34306 ( .A(n25714), .B(n18070), .Z(n13641) );
  NANDN U34307 ( .A(init), .B(m[711]), .Z(n18070) );
  AND U34308 ( .A(n25715), .B(n25716), .Z(n25714) );
  NAND U34309 ( .A(o[711]), .B(n23579), .Z(n25716) );
  NANDN U34310 ( .A(n23580), .B(creg[711]), .Z(n25715) );
  NAND U34311 ( .A(n25717), .B(n18068), .Z(n13640) );
  NANDN U34312 ( .A(init), .B(m[712]), .Z(n18068) );
  AND U34313 ( .A(n25718), .B(n25719), .Z(n25717) );
  NAND U34314 ( .A(o[712]), .B(n23579), .Z(n25719) );
  NANDN U34315 ( .A(n23580), .B(creg[712]), .Z(n25718) );
  NAND U34316 ( .A(n25720), .B(n18066), .Z(n13639) );
  NANDN U34317 ( .A(init), .B(m[713]), .Z(n18066) );
  AND U34318 ( .A(n25721), .B(n25722), .Z(n25720) );
  NAND U34319 ( .A(o[713]), .B(n23579), .Z(n25722) );
  NANDN U34320 ( .A(n23580), .B(creg[713]), .Z(n25721) );
  NAND U34321 ( .A(n25723), .B(n18064), .Z(n13638) );
  NANDN U34322 ( .A(init), .B(m[714]), .Z(n18064) );
  AND U34323 ( .A(n25724), .B(n25725), .Z(n25723) );
  NAND U34324 ( .A(o[714]), .B(n23579), .Z(n25725) );
  NANDN U34325 ( .A(n23580), .B(creg[714]), .Z(n25724) );
  NAND U34326 ( .A(n25726), .B(n18062), .Z(n13637) );
  NANDN U34327 ( .A(init), .B(m[715]), .Z(n18062) );
  AND U34328 ( .A(n25727), .B(n25728), .Z(n25726) );
  NAND U34329 ( .A(o[715]), .B(n23579), .Z(n25728) );
  NANDN U34330 ( .A(n23580), .B(creg[715]), .Z(n25727) );
  NAND U34331 ( .A(n25729), .B(n18060), .Z(n13636) );
  NANDN U34332 ( .A(init), .B(m[716]), .Z(n18060) );
  AND U34333 ( .A(n25730), .B(n25731), .Z(n25729) );
  NAND U34334 ( .A(o[716]), .B(n23579), .Z(n25731) );
  NANDN U34335 ( .A(n23580), .B(creg[716]), .Z(n25730) );
  NAND U34336 ( .A(n25732), .B(n18058), .Z(n13635) );
  NANDN U34337 ( .A(init), .B(m[717]), .Z(n18058) );
  AND U34338 ( .A(n25733), .B(n25734), .Z(n25732) );
  NAND U34339 ( .A(o[717]), .B(n23579), .Z(n25734) );
  NANDN U34340 ( .A(n23580), .B(creg[717]), .Z(n25733) );
  NAND U34341 ( .A(n25735), .B(n18056), .Z(n13634) );
  NANDN U34342 ( .A(init), .B(m[718]), .Z(n18056) );
  AND U34343 ( .A(n25736), .B(n25737), .Z(n25735) );
  NAND U34344 ( .A(o[718]), .B(n23579), .Z(n25737) );
  NANDN U34345 ( .A(n23580), .B(creg[718]), .Z(n25736) );
  NAND U34346 ( .A(n25738), .B(n18054), .Z(n13633) );
  NANDN U34347 ( .A(init), .B(m[719]), .Z(n18054) );
  AND U34348 ( .A(n25739), .B(n25740), .Z(n25738) );
  NAND U34349 ( .A(o[719]), .B(n23579), .Z(n25740) );
  NANDN U34350 ( .A(n23580), .B(creg[719]), .Z(n25739) );
  NAND U34351 ( .A(n25741), .B(n18050), .Z(n13632) );
  NANDN U34352 ( .A(init), .B(m[720]), .Z(n18050) );
  AND U34353 ( .A(n25742), .B(n25743), .Z(n25741) );
  NAND U34354 ( .A(o[720]), .B(n23579), .Z(n25743) );
  NANDN U34355 ( .A(n23580), .B(creg[720]), .Z(n25742) );
  NAND U34356 ( .A(n25744), .B(n18048), .Z(n13631) );
  NANDN U34357 ( .A(init), .B(m[721]), .Z(n18048) );
  AND U34358 ( .A(n25745), .B(n25746), .Z(n25744) );
  NAND U34359 ( .A(o[721]), .B(n23579), .Z(n25746) );
  NANDN U34360 ( .A(n23580), .B(creg[721]), .Z(n25745) );
  NAND U34361 ( .A(n25747), .B(n18046), .Z(n13630) );
  NANDN U34362 ( .A(init), .B(m[722]), .Z(n18046) );
  AND U34363 ( .A(n25748), .B(n25749), .Z(n25747) );
  NAND U34364 ( .A(o[722]), .B(n23579), .Z(n25749) );
  NANDN U34365 ( .A(n23580), .B(creg[722]), .Z(n25748) );
  NAND U34366 ( .A(n25750), .B(n18044), .Z(n13629) );
  NANDN U34367 ( .A(init), .B(m[723]), .Z(n18044) );
  AND U34368 ( .A(n25751), .B(n25752), .Z(n25750) );
  NAND U34369 ( .A(o[723]), .B(n23579), .Z(n25752) );
  NANDN U34370 ( .A(n23580), .B(creg[723]), .Z(n25751) );
  NAND U34371 ( .A(n25753), .B(n18042), .Z(n13628) );
  NANDN U34372 ( .A(init), .B(m[724]), .Z(n18042) );
  AND U34373 ( .A(n25754), .B(n25755), .Z(n25753) );
  NAND U34374 ( .A(o[724]), .B(n23579), .Z(n25755) );
  NANDN U34375 ( .A(n23580), .B(creg[724]), .Z(n25754) );
  NAND U34376 ( .A(n25756), .B(n18040), .Z(n13627) );
  NANDN U34377 ( .A(init), .B(m[725]), .Z(n18040) );
  AND U34378 ( .A(n25757), .B(n25758), .Z(n25756) );
  NAND U34379 ( .A(o[725]), .B(n23579), .Z(n25758) );
  NANDN U34380 ( .A(n23580), .B(creg[725]), .Z(n25757) );
  NAND U34381 ( .A(n25759), .B(n18038), .Z(n13626) );
  NANDN U34382 ( .A(init), .B(m[726]), .Z(n18038) );
  AND U34383 ( .A(n25760), .B(n25761), .Z(n25759) );
  NAND U34384 ( .A(o[726]), .B(n23579), .Z(n25761) );
  NANDN U34385 ( .A(n23580), .B(creg[726]), .Z(n25760) );
  NAND U34386 ( .A(n25762), .B(n18036), .Z(n13625) );
  NANDN U34387 ( .A(init), .B(m[727]), .Z(n18036) );
  AND U34388 ( .A(n25763), .B(n25764), .Z(n25762) );
  NAND U34389 ( .A(o[727]), .B(n23579), .Z(n25764) );
  NANDN U34390 ( .A(n23580), .B(creg[727]), .Z(n25763) );
  NAND U34391 ( .A(n25765), .B(n18034), .Z(n13624) );
  NANDN U34392 ( .A(init), .B(m[728]), .Z(n18034) );
  AND U34393 ( .A(n25766), .B(n25767), .Z(n25765) );
  NAND U34394 ( .A(o[728]), .B(n23579), .Z(n25767) );
  NANDN U34395 ( .A(n23580), .B(creg[728]), .Z(n25766) );
  NAND U34396 ( .A(n25768), .B(n18032), .Z(n13623) );
  NANDN U34397 ( .A(init), .B(m[729]), .Z(n18032) );
  AND U34398 ( .A(n25769), .B(n25770), .Z(n25768) );
  NAND U34399 ( .A(o[729]), .B(n23579), .Z(n25770) );
  NANDN U34400 ( .A(n23580), .B(creg[729]), .Z(n25769) );
  NAND U34401 ( .A(n25771), .B(n18028), .Z(n13622) );
  NANDN U34402 ( .A(init), .B(m[730]), .Z(n18028) );
  AND U34403 ( .A(n25772), .B(n25773), .Z(n25771) );
  NAND U34404 ( .A(o[730]), .B(n23579), .Z(n25773) );
  NANDN U34405 ( .A(n23580), .B(creg[730]), .Z(n25772) );
  NAND U34406 ( .A(n25774), .B(n18026), .Z(n13621) );
  NANDN U34407 ( .A(init), .B(m[731]), .Z(n18026) );
  AND U34408 ( .A(n25775), .B(n25776), .Z(n25774) );
  NAND U34409 ( .A(o[731]), .B(n23579), .Z(n25776) );
  NANDN U34410 ( .A(n23580), .B(creg[731]), .Z(n25775) );
  NAND U34411 ( .A(n25777), .B(n18024), .Z(n13620) );
  NANDN U34412 ( .A(init), .B(m[732]), .Z(n18024) );
  AND U34413 ( .A(n25778), .B(n25779), .Z(n25777) );
  NAND U34414 ( .A(o[732]), .B(n23579), .Z(n25779) );
  NANDN U34415 ( .A(n23580), .B(creg[732]), .Z(n25778) );
  NAND U34416 ( .A(n25780), .B(n18022), .Z(n13619) );
  NANDN U34417 ( .A(init), .B(m[733]), .Z(n18022) );
  AND U34418 ( .A(n25781), .B(n25782), .Z(n25780) );
  NAND U34419 ( .A(o[733]), .B(n23579), .Z(n25782) );
  NANDN U34420 ( .A(n23580), .B(creg[733]), .Z(n25781) );
  NAND U34421 ( .A(n25783), .B(n18020), .Z(n13618) );
  NANDN U34422 ( .A(init), .B(m[734]), .Z(n18020) );
  AND U34423 ( .A(n25784), .B(n25785), .Z(n25783) );
  NAND U34424 ( .A(o[734]), .B(n23579), .Z(n25785) );
  NANDN U34425 ( .A(n23580), .B(creg[734]), .Z(n25784) );
  NAND U34426 ( .A(n25786), .B(n18018), .Z(n13617) );
  NANDN U34427 ( .A(init), .B(m[735]), .Z(n18018) );
  AND U34428 ( .A(n25787), .B(n25788), .Z(n25786) );
  NAND U34429 ( .A(o[735]), .B(n23579), .Z(n25788) );
  NANDN U34430 ( .A(n23580), .B(creg[735]), .Z(n25787) );
  NAND U34431 ( .A(n25789), .B(n18016), .Z(n13616) );
  NANDN U34432 ( .A(init), .B(m[736]), .Z(n18016) );
  AND U34433 ( .A(n25790), .B(n25791), .Z(n25789) );
  NAND U34434 ( .A(o[736]), .B(n23579), .Z(n25791) );
  NANDN U34435 ( .A(n23580), .B(creg[736]), .Z(n25790) );
  NAND U34436 ( .A(n25792), .B(n18014), .Z(n13615) );
  NANDN U34437 ( .A(init), .B(m[737]), .Z(n18014) );
  AND U34438 ( .A(n25793), .B(n25794), .Z(n25792) );
  NAND U34439 ( .A(o[737]), .B(n23579), .Z(n25794) );
  NANDN U34440 ( .A(n23580), .B(creg[737]), .Z(n25793) );
  NAND U34441 ( .A(n25795), .B(n18012), .Z(n13614) );
  NANDN U34442 ( .A(init), .B(m[738]), .Z(n18012) );
  AND U34443 ( .A(n25796), .B(n25797), .Z(n25795) );
  NAND U34444 ( .A(o[738]), .B(n23579), .Z(n25797) );
  NANDN U34445 ( .A(n23580), .B(creg[738]), .Z(n25796) );
  NAND U34446 ( .A(n25798), .B(n18010), .Z(n13613) );
  NANDN U34447 ( .A(init), .B(m[739]), .Z(n18010) );
  AND U34448 ( .A(n25799), .B(n25800), .Z(n25798) );
  NAND U34449 ( .A(o[739]), .B(n23579), .Z(n25800) );
  NANDN U34450 ( .A(n23580), .B(creg[739]), .Z(n25799) );
  NAND U34451 ( .A(n25801), .B(n18006), .Z(n13612) );
  NANDN U34452 ( .A(init), .B(m[740]), .Z(n18006) );
  AND U34453 ( .A(n25802), .B(n25803), .Z(n25801) );
  NAND U34454 ( .A(o[740]), .B(n23579), .Z(n25803) );
  NANDN U34455 ( .A(n23580), .B(creg[740]), .Z(n25802) );
  NAND U34456 ( .A(n25804), .B(n18004), .Z(n13611) );
  NANDN U34457 ( .A(init), .B(m[741]), .Z(n18004) );
  AND U34458 ( .A(n25805), .B(n25806), .Z(n25804) );
  NAND U34459 ( .A(o[741]), .B(n23579), .Z(n25806) );
  NANDN U34460 ( .A(n23580), .B(creg[741]), .Z(n25805) );
  NAND U34461 ( .A(n25807), .B(n18002), .Z(n13610) );
  NANDN U34462 ( .A(init), .B(m[742]), .Z(n18002) );
  AND U34463 ( .A(n25808), .B(n25809), .Z(n25807) );
  NAND U34464 ( .A(o[742]), .B(n23579), .Z(n25809) );
  NANDN U34465 ( .A(n23580), .B(creg[742]), .Z(n25808) );
  NAND U34466 ( .A(n25810), .B(n18000), .Z(n13609) );
  NANDN U34467 ( .A(init), .B(m[743]), .Z(n18000) );
  AND U34468 ( .A(n25811), .B(n25812), .Z(n25810) );
  NAND U34469 ( .A(o[743]), .B(n23579), .Z(n25812) );
  NANDN U34470 ( .A(n23580), .B(creg[743]), .Z(n25811) );
  NAND U34471 ( .A(n25813), .B(n17998), .Z(n13608) );
  NANDN U34472 ( .A(init), .B(m[744]), .Z(n17998) );
  AND U34473 ( .A(n25814), .B(n25815), .Z(n25813) );
  NAND U34474 ( .A(o[744]), .B(n23579), .Z(n25815) );
  NANDN U34475 ( .A(n23580), .B(creg[744]), .Z(n25814) );
  NAND U34476 ( .A(n25816), .B(n17996), .Z(n13607) );
  NANDN U34477 ( .A(init), .B(m[745]), .Z(n17996) );
  AND U34478 ( .A(n25817), .B(n25818), .Z(n25816) );
  NAND U34479 ( .A(o[745]), .B(n23579), .Z(n25818) );
  NANDN U34480 ( .A(n23580), .B(creg[745]), .Z(n25817) );
  NAND U34481 ( .A(n25819), .B(n17994), .Z(n13606) );
  NANDN U34482 ( .A(init), .B(m[746]), .Z(n17994) );
  AND U34483 ( .A(n25820), .B(n25821), .Z(n25819) );
  NAND U34484 ( .A(o[746]), .B(n23579), .Z(n25821) );
  NANDN U34485 ( .A(n23580), .B(creg[746]), .Z(n25820) );
  NAND U34486 ( .A(n25822), .B(n17992), .Z(n13605) );
  NANDN U34487 ( .A(init), .B(m[747]), .Z(n17992) );
  AND U34488 ( .A(n25823), .B(n25824), .Z(n25822) );
  NAND U34489 ( .A(o[747]), .B(n23579), .Z(n25824) );
  NANDN U34490 ( .A(n23580), .B(creg[747]), .Z(n25823) );
  NAND U34491 ( .A(n25825), .B(n17990), .Z(n13604) );
  NANDN U34492 ( .A(init), .B(m[748]), .Z(n17990) );
  AND U34493 ( .A(n25826), .B(n25827), .Z(n25825) );
  NAND U34494 ( .A(o[748]), .B(n23579), .Z(n25827) );
  NANDN U34495 ( .A(n23580), .B(creg[748]), .Z(n25826) );
  NAND U34496 ( .A(n25828), .B(n17988), .Z(n13603) );
  NANDN U34497 ( .A(init), .B(m[749]), .Z(n17988) );
  AND U34498 ( .A(n25829), .B(n25830), .Z(n25828) );
  NAND U34499 ( .A(o[749]), .B(n23579), .Z(n25830) );
  NANDN U34500 ( .A(n23580), .B(creg[749]), .Z(n25829) );
  NAND U34501 ( .A(n25831), .B(n17984), .Z(n13602) );
  NANDN U34502 ( .A(init), .B(m[750]), .Z(n17984) );
  AND U34503 ( .A(n25832), .B(n25833), .Z(n25831) );
  NAND U34504 ( .A(o[750]), .B(n23579), .Z(n25833) );
  NANDN U34505 ( .A(n23580), .B(creg[750]), .Z(n25832) );
  NAND U34506 ( .A(n25834), .B(n17982), .Z(n13601) );
  NANDN U34507 ( .A(init), .B(m[751]), .Z(n17982) );
  AND U34508 ( .A(n25835), .B(n25836), .Z(n25834) );
  NAND U34509 ( .A(o[751]), .B(n23579), .Z(n25836) );
  NANDN U34510 ( .A(n23580), .B(creg[751]), .Z(n25835) );
  NAND U34511 ( .A(n25837), .B(n17980), .Z(n13600) );
  NANDN U34512 ( .A(init), .B(m[752]), .Z(n17980) );
  AND U34513 ( .A(n25838), .B(n25839), .Z(n25837) );
  NAND U34514 ( .A(o[752]), .B(n23579), .Z(n25839) );
  NANDN U34515 ( .A(n23580), .B(creg[752]), .Z(n25838) );
  NAND U34516 ( .A(n25840), .B(n17978), .Z(n13599) );
  NANDN U34517 ( .A(init), .B(m[753]), .Z(n17978) );
  AND U34518 ( .A(n25841), .B(n25842), .Z(n25840) );
  NAND U34519 ( .A(o[753]), .B(n23579), .Z(n25842) );
  NANDN U34520 ( .A(n23580), .B(creg[753]), .Z(n25841) );
  NAND U34521 ( .A(n25843), .B(n17976), .Z(n13598) );
  NANDN U34522 ( .A(init), .B(m[754]), .Z(n17976) );
  AND U34523 ( .A(n25844), .B(n25845), .Z(n25843) );
  NAND U34524 ( .A(o[754]), .B(n23579), .Z(n25845) );
  NANDN U34525 ( .A(n23580), .B(creg[754]), .Z(n25844) );
  NAND U34526 ( .A(n25846), .B(n17974), .Z(n13597) );
  NANDN U34527 ( .A(init), .B(m[755]), .Z(n17974) );
  AND U34528 ( .A(n25847), .B(n25848), .Z(n25846) );
  NAND U34529 ( .A(o[755]), .B(n23579), .Z(n25848) );
  NANDN U34530 ( .A(n23580), .B(creg[755]), .Z(n25847) );
  NAND U34531 ( .A(n25849), .B(n17972), .Z(n13596) );
  NANDN U34532 ( .A(init), .B(m[756]), .Z(n17972) );
  AND U34533 ( .A(n25850), .B(n25851), .Z(n25849) );
  NAND U34534 ( .A(o[756]), .B(n23579), .Z(n25851) );
  NANDN U34535 ( .A(n23580), .B(creg[756]), .Z(n25850) );
  NAND U34536 ( .A(n25852), .B(n17970), .Z(n13595) );
  NANDN U34537 ( .A(init), .B(m[757]), .Z(n17970) );
  AND U34538 ( .A(n25853), .B(n25854), .Z(n25852) );
  NAND U34539 ( .A(o[757]), .B(n23579), .Z(n25854) );
  NANDN U34540 ( .A(n23580), .B(creg[757]), .Z(n25853) );
  NAND U34541 ( .A(n25855), .B(n17968), .Z(n13594) );
  NANDN U34542 ( .A(init), .B(m[758]), .Z(n17968) );
  AND U34543 ( .A(n25856), .B(n25857), .Z(n25855) );
  NAND U34544 ( .A(o[758]), .B(n23579), .Z(n25857) );
  NANDN U34545 ( .A(n23580), .B(creg[758]), .Z(n25856) );
  NAND U34546 ( .A(n25858), .B(n17966), .Z(n13593) );
  NANDN U34547 ( .A(init), .B(m[759]), .Z(n17966) );
  AND U34548 ( .A(n25859), .B(n25860), .Z(n25858) );
  NAND U34549 ( .A(o[759]), .B(n23579), .Z(n25860) );
  NANDN U34550 ( .A(n23580), .B(creg[759]), .Z(n25859) );
  NAND U34551 ( .A(n25861), .B(n17962), .Z(n13592) );
  NANDN U34552 ( .A(init), .B(m[760]), .Z(n17962) );
  AND U34553 ( .A(n25862), .B(n25863), .Z(n25861) );
  NAND U34554 ( .A(o[760]), .B(n23579), .Z(n25863) );
  NANDN U34555 ( .A(n23580), .B(creg[760]), .Z(n25862) );
  NAND U34556 ( .A(n25864), .B(n17960), .Z(n13591) );
  NANDN U34557 ( .A(init), .B(m[761]), .Z(n17960) );
  AND U34558 ( .A(n25865), .B(n25866), .Z(n25864) );
  NAND U34559 ( .A(o[761]), .B(n23579), .Z(n25866) );
  NANDN U34560 ( .A(n23580), .B(creg[761]), .Z(n25865) );
  NAND U34561 ( .A(n25867), .B(n17958), .Z(n13590) );
  NANDN U34562 ( .A(init), .B(m[762]), .Z(n17958) );
  AND U34563 ( .A(n25868), .B(n25869), .Z(n25867) );
  NAND U34564 ( .A(o[762]), .B(n23579), .Z(n25869) );
  NANDN U34565 ( .A(n23580), .B(creg[762]), .Z(n25868) );
  NAND U34566 ( .A(n25870), .B(n17956), .Z(n13589) );
  NANDN U34567 ( .A(init), .B(m[763]), .Z(n17956) );
  AND U34568 ( .A(n25871), .B(n25872), .Z(n25870) );
  NAND U34569 ( .A(o[763]), .B(n23579), .Z(n25872) );
  NANDN U34570 ( .A(n23580), .B(creg[763]), .Z(n25871) );
  NAND U34571 ( .A(n25873), .B(n17954), .Z(n13588) );
  NANDN U34572 ( .A(init), .B(m[764]), .Z(n17954) );
  AND U34573 ( .A(n25874), .B(n25875), .Z(n25873) );
  NAND U34574 ( .A(o[764]), .B(n23579), .Z(n25875) );
  NANDN U34575 ( .A(n23580), .B(creg[764]), .Z(n25874) );
  NAND U34576 ( .A(n25876), .B(n17952), .Z(n13587) );
  NANDN U34577 ( .A(init), .B(m[765]), .Z(n17952) );
  AND U34578 ( .A(n25877), .B(n25878), .Z(n25876) );
  NAND U34579 ( .A(o[765]), .B(n23579), .Z(n25878) );
  NANDN U34580 ( .A(n23580), .B(creg[765]), .Z(n25877) );
  NAND U34581 ( .A(n25879), .B(n17950), .Z(n13586) );
  NANDN U34582 ( .A(init), .B(m[766]), .Z(n17950) );
  AND U34583 ( .A(n25880), .B(n25881), .Z(n25879) );
  NAND U34584 ( .A(o[766]), .B(n23579), .Z(n25881) );
  NANDN U34585 ( .A(n23580), .B(creg[766]), .Z(n25880) );
  NAND U34586 ( .A(n25882), .B(n17948), .Z(n13585) );
  NANDN U34587 ( .A(init), .B(m[767]), .Z(n17948) );
  AND U34588 ( .A(n25883), .B(n25884), .Z(n25882) );
  NAND U34589 ( .A(o[767]), .B(n23579), .Z(n25884) );
  NANDN U34590 ( .A(n23580), .B(creg[767]), .Z(n25883) );
  NAND U34591 ( .A(n25885), .B(n17946), .Z(n13584) );
  NANDN U34592 ( .A(init), .B(m[768]), .Z(n17946) );
  AND U34593 ( .A(n25886), .B(n25887), .Z(n25885) );
  NAND U34594 ( .A(o[768]), .B(n23579), .Z(n25887) );
  NANDN U34595 ( .A(n23580), .B(creg[768]), .Z(n25886) );
  NAND U34596 ( .A(n25888), .B(n17944), .Z(n13583) );
  NANDN U34597 ( .A(init), .B(m[769]), .Z(n17944) );
  AND U34598 ( .A(n25889), .B(n25890), .Z(n25888) );
  NAND U34599 ( .A(o[769]), .B(n23579), .Z(n25890) );
  NANDN U34600 ( .A(n23580), .B(creg[769]), .Z(n25889) );
  NAND U34601 ( .A(n25891), .B(n17940), .Z(n13582) );
  NANDN U34602 ( .A(init), .B(m[770]), .Z(n17940) );
  AND U34603 ( .A(n25892), .B(n25893), .Z(n25891) );
  NAND U34604 ( .A(o[770]), .B(n23579), .Z(n25893) );
  NANDN U34605 ( .A(n23580), .B(creg[770]), .Z(n25892) );
  NAND U34606 ( .A(n25894), .B(n17938), .Z(n13581) );
  NANDN U34607 ( .A(init), .B(m[771]), .Z(n17938) );
  AND U34608 ( .A(n25895), .B(n25896), .Z(n25894) );
  NAND U34609 ( .A(o[771]), .B(n23579), .Z(n25896) );
  NANDN U34610 ( .A(n23580), .B(creg[771]), .Z(n25895) );
  NAND U34611 ( .A(n25897), .B(n17936), .Z(n13580) );
  NANDN U34612 ( .A(init), .B(m[772]), .Z(n17936) );
  AND U34613 ( .A(n25898), .B(n25899), .Z(n25897) );
  NAND U34614 ( .A(o[772]), .B(n23579), .Z(n25899) );
  NANDN U34615 ( .A(n23580), .B(creg[772]), .Z(n25898) );
  NAND U34616 ( .A(n25900), .B(n17934), .Z(n13579) );
  NANDN U34617 ( .A(init), .B(m[773]), .Z(n17934) );
  AND U34618 ( .A(n25901), .B(n25902), .Z(n25900) );
  NAND U34619 ( .A(o[773]), .B(n23579), .Z(n25902) );
  NANDN U34620 ( .A(n23580), .B(creg[773]), .Z(n25901) );
  NAND U34621 ( .A(n25903), .B(n17932), .Z(n13578) );
  NANDN U34622 ( .A(init), .B(m[774]), .Z(n17932) );
  AND U34623 ( .A(n25904), .B(n25905), .Z(n25903) );
  NAND U34624 ( .A(o[774]), .B(n23579), .Z(n25905) );
  NANDN U34625 ( .A(n23580), .B(creg[774]), .Z(n25904) );
  NAND U34626 ( .A(n25906), .B(n17930), .Z(n13577) );
  NANDN U34627 ( .A(init), .B(m[775]), .Z(n17930) );
  AND U34628 ( .A(n25907), .B(n25908), .Z(n25906) );
  NAND U34629 ( .A(o[775]), .B(n23579), .Z(n25908) );
  NANDN U34630 ( .A(n23580), .B(creg[775]), .Z(n25907) );
  NAND U34631 ( .A(n25909), .B(n17928), .Z(n13576) );
  NANDN U34632 ( .A(init), .B(m[776]), .Z(n17928) );
  AND U34633 ( .A(n25910), .B(n25911), .Z(n25909) );
  NAND U34634 ( .A(o[776]), .B(n23579), .Z(n25911) );
  NANDN U34635 ( .A(n23580), .B(creg[776]), .Z(n25910) );
  NAND U34636 ( .A(n25912), .B(n17926), .Z(n13575) );
  NANDN U34637 ( .A(init), .B(m[777]), .Z(n17926) );
  AND U34638 ( .A(n25913), .B(n25914), .Z(n25912) );
  NAND U34639 ( .A(o[777]), .B(n23579), .Z(n25914) );
  NANDN U34640 ( .A(n23580), .B(creg[777]), .Z(n25913) );
  NAND U34641 ( .A(n25915), .B(n17924), .Z(n13574) );
  NANDN U34642 ( .A(init), .B(m[778]), .Z(n17924) );
  AND U34643 ( .A(n25916), .B(n25917), .Z(n25915) );
  NAND U34644 ( .A(o[778]), .B(n23579), .Z(n25917) );
  NANDN U34645 ( .A(n23580), .B(creg[778]), .Z(n25916) );
  NAND U34646 ( .A(n25918), .B(n17922), .Z(n13573) );
  NANDN U34647 ( .A(init), .B(m[779]), .Z(n17922) );
  AND U34648 ( .A(n25919), .B(n25920), .Z(n25918) );
  NAND U34649 ( .A(o[779]), .B(n23579), .Z(n25920) );
  NANDN U34650 ( .A(n23580), .B(creg[779]), .Z(n25919) );
  NAND U34651 ( .A(n25921), .B(n17918), .Z(n13572) );
  NANDN U34652 ( .A(init), .B(m[780]), .Z(n17918) );
  AND U34653 ( .A(n25922), .B(n25923), .Z(n25921) );
  NAND U34654 ( .A(o[780]), .B(n23579), .Z(n25923) );
  NANDN U34655 ( .A(n23580), .B(creg[780]), .Z(n25922) );
  NAND U34656 ( .A(n25924), .B(n17916), .Z(n13571) );
  NANDN U34657 ( .A(init), .B(m[781]), .Z(n17916) );
  AND U34658 ( .A(n25925), .B(n25926), .Z(n25924) );
  NAND U34659 ( .A(o[781]), .B(n23579), .Z(n25926) );
  NANDN U34660 ( .A(n23580), .B(creg[781]), .Z(n25925) );
  NAND U34661 ( .A(n25927), .B(n17914), .Z(n13570) );
  NANDN U34662 ( .A(init), .B(m[782]), .Z(n17914) );
  AND U34663 ( .A(n25928), .B(n25929), .Z(n25927) );
  NAND U34664 ( .A(o[782]), .B(n23579), .Z(n25929) );
  NANDN U34665 ( .A(n23580), .B(creg[782]), .Z(n25928) );
  NAND U34666 ( .A(n25930), .B(n17912), .Z(n13569) );
  NANDN U34667 ( .A(init), .B(m[783]), .Z(n17912) );
  AND U34668 ( .A(n25931), .B(n25932), .Z(n25930) );
  NAND U34669 ( .A(o[783]), .B(n23579), .Z(n25932) );
  NANDN U34670 ( .A(n23580), .B(creg[783]), .Z(n25931) );
  NAND U34671 ( .A(n25933), .B(n17910), .Z(n13568) );
  NANDN U34672 ( .A(init), .B(m[784]), .Z(n17910) );
  AND U34673 ( .A(n25934), .B(n25935), .Z(n25933) );
  NAND U34674 ( .A(o[784]), .B(n23579), .Z(n25935) );
  NANDN U34675 ( .A(n23580), .B(creg[784]), .Z(n25934) );
  NAND U34676 ( .A(n25936), .B(n17908), .Z(n13567) );
  NANDN U34677 ( .A(init), .B(m[785]), .Z(n17908) );
  AND U34678 ( .A(n25937), .B(n25938), .Z(n25936) );
  NAND U34679 ( .A(o[785]), .B(n23579), .Z(n25938) );
  NANDN U34680 ( .A(n23580), .B(creg[785]), .Z(n25937) );
  NAND U34681 ( .A(n25939), .B(n17906), .Z(n13566) );
  NANDN U34682 ( .A(init), .B(m[786]), .Z(n17906) );
  AND U34683 ( .A(n25940), .B(n25941), .Z(n25939) );
  NAND U34684 ( .A(o[786]), .B(n23579), .Z(n25941) );
  NANDN U34685 ( .A(n23580), .B(creg[786]), .Z(n25940) );
  NAND U34686 ( .A(n25942), .B(n17904), .Z(n13565) );
  NANDN U34687 ( .A(init), .B(m[787]), .Z(n17904) );
  AND U34688 ( .A(n25943), .B(n25944), .Z(n25942) );
  NAND U34689 ( .A(o[787]), .B(n23579), .Z(n25944) );
  NANDN U34690 ( .A(n23580), .B(creg[787]), .Z(n25943) );
  NAND U34691 ( .A(n25945), .B(n17902), .Z(n13564) );
  NANDN U34692 ( .A(init), .B(m[788]), .Z(n17902) );
  AND U34693 ( .A(n25946), .B(n25947), .Z(n25945) );
  NAND U34694 ( .A(o[788]), .B(n23579), .Z(n25947) );
  NANDN U34695 ( .A(n23580), .B(creg[788]), .Z(n25946) );
  NAND U34696 ( .A(n25948), .B(n17900), .Z(n13563) );
  NANDN U34697 ( .A(init), .B(m[789]), .Z(n17900) );
  AND U34698 ( .A(n25949), .B(n25950), .Z(n25948) );
  NAND U34699 ( .A(o[789]), .B(n23579), .Z(n25950) );
  NANDN U34700 ( .A(n23580), .B(creg[789]), .Z(n25949) );
  NAND U34701 ( .A(n25951), .B(n17896), .Z(n13562) );
  NANDN U34702 ( .A(init), .B(m[790]), .Z(n17896) );
  AND U34703 ( .A(n25952), .B(n25953), .Z(n25951) );
  NAND U34704 ( .A(o[790]), .B(n23579), .Z(n25953) );
  NANDN U34705 ( .A(n23580), .B(creg[790]), .Z(n25952) );
  NAND U34706 ( .A(n25954), .B(n17894), .Z(n13561) );
  NANDN U34707 ( .A(init), .B(m[791]), .Z(n17894) );
  AND U34708 ( .A(n25955), .B(n25956), .Z(n25954) );
  NAND U34709 ( .A(o[791]), .B(n23579), .Z(n25956) );
  NANDN U34710 ( .A(n23580), .B(creg[791]), .Z(n25955) );
  NAND U34711 ( .A(n25957), .B(n17892), .Z(n13560) );
  NANDN U34712 ( .A(init), .B(m[792]), .Z(n17892) );
  AND U34713 ( .A(n25958), .B(n25959), .Z(n25957) );
  NAND U34714 ( .A(o[792]), .B(n23579), .Z(n25959) );
  NANDN U34715 ( .A(n23580), .B(creg[792]), .Z(n25958) );
  NAND U34716 ( .A(n25960), .B(n17890), .Z(n13559) );
  NANDN U34717 ( .A(init), .B(m[793]), .Z(n17890) );
  AND U34718 ( .A(n25961), .B(n25962), .Z(n25960) );
  NAND U34719 ( .A(o[793]), .B(n23579), .Z(n25962) );
  NANDN U34720 ( .A(n23580), .B(creg[793]), .Z(n25961) );
  NAND U34721 ( .A(n25963), .B(n17888), .Z(n13558) );
  NANDN U34722 ( .A(init), .B(m[794]), .Z(n17888) );
  AND U34723 ( .A(n25964), .B(n25965), .Z(n25963) );
  NAND U34724 ( .A(o[794]), .B(n23579), .Z(n25965) );
  NANDN U34725 ( .A(n23580), .B(creg[794]), .Z(n25964) );
  NAND U34726 ( .A(n25966), .B(n17886), .Z(n13557) );
  NANDN U34727 ( .A(init), .B(m[795]), .Z(n17886) );
  AND U34728 ( .A(n25967), .B(n25968), .Z(n25966) );
  NAND U34729 ( .A(o[795]), .B(n23579), .Z(n25968) );
  NANDN U34730 ( .A(n23580), .B(creg[795]), .Z(n25967) );
  NAND U34731 ( .A(n25969), .B(n17884), .Z(n13556) );
  NANDN U34732 ( .A(init), .B(m[796]), .Z(n17884) );
  AND U34733 ( .A(n25970), .B(n25971), .Z(n25969) );
  NAND U34734 ( .A(o[796]), .B(n23579), .Z(n25971) );
  NANDN U34735 ( .A(n23580), .B(creg[796]), .Z(n25970) );
  NAND U34736 ( .A(n25972), .B(n17882), .Z(n13555) );
  NANDN U34737 ( .A(init), .B(m[797]), .Z(n17882) );
  AND U34738 ( .A(n25973), .B(n25974), .Z(n25972) );
  NAND U34739 ( .A(o[797]), .B(n23579), .Z(n25974) );
  NANDN U34740 ( .A(n23580), .B(creg[797]), .Z(n25973) );
  NAND U34741 ( .A(n25975), .B(n17880), .Z(n13554) );
  NANDN U34742 ( .A(init), .B(m[798]), .Z(n17880) );
  AND U34743 ( .A(n25976), .B(n25977), .Z(n25975) );
  NAND U34744 ( .A(o[798]), .B(n23579), .Z(n25977) );
  NANDN U34745 ( .A(n23580), .B(creg[798]), .Z(n25976) );
  NAND U34746 ( .A(n25978), .B(n17878), .Z(n13553) );
  NANDN U34747 ( .A(init), .B(m[799]), .Z(n17878) );
  AND U34748 ( .A(n25979), .B(n25980), .Z(n25978) );
  NAND U34749 ( .A(o[799]), .B(n23579), .Z(n25980) );
  NANDN U34750 ( .A(n23580), .B(creg[799]), .Z(n25979) );
  NAND U34751 ( .A(n25981), .B(n17872), .Z(n13552) );
  NANDN U34752 ( .A(init), .B(m[800]), .Z(n17872) );
  AND U34753 ( .A(n25982), .B(n25983), .Z(n25981) );
  NAND U34754 ( .A(o[800]), .B(n23579), .Z(n25983) );
  NANDN U34755 ( .A(n23580), .B(creg[800]), .Z(n25982) );
  NAND U34756 ( .A(n25984), .B(n17870), .Z(n13551) );
  NANDN U34757 ( .A(init), .B(m[801]), .Z(n17870) );
  AND U34758 ( .A(n25985), .B(n25986), .Z(n25984) );
  NAND U34759 ( .A(o[801]), .B(n23579), .Z(n25986) );
  NANDN U34760 ( .A(n23580), .B(creg[801]), .Z(n25985) );
  NAND U34761 ( .A(n25987), .B(n17868), .Z(n13550) );
  NANDN U34762 ( .A(init), .B(m[802]), .Z(n17868) );
  AND U34763 ( .A(n25988), .B(n25989), .Z(n25987) );
  NAND U34764 ( .A(o[802]), .B(n23579), .Z(n25989) );
  NANDN U34765 ( .A(n23580), .B(creg[802]), .Z(n25988) );
  NAND U34766 ( .A(n25990), .B(n17866), .Z(n13549) );
  NANDN U34767 ( .A(init), .B(m[803]), .Z(n17866) );
  AND U34768 ( .A(n25991), .B(n25992), .Z(n25990) );
  NAND U34769 ( .A(o[803]), .B(n23579), .Z(n25992) );
  NANDN U34770 ( .A(n23580), .B(creg[803]), .Z(n25991) );
  NAND U34771 ( .A(n25993), .B(n17864), .Z(n13548) );
  NANDN U34772 ( .A(init), .B(m[804]), .Z(n17864) );
  AND U34773 ( .A(n25994), .B(n25995), .Z(n25993) );
  NAND U34774 ( .A(o[804]), .B(n23579), .Z(n25995) );
  NANDN U34775 ( .A(n23580), .B(creg[804]), .Z(n25994) );
  NAND U34776 ( .A(n25996), .B(n17862), .Z(n13547) );
  NANDN U34777 ( .A(init), .B(m[805]), .Z(n17862) );
  AND U34778 ( .A(n25997), .B(n25998), .Z(n25996) );
  NAND U34779 ( .A(o[805]), .B(n23579), .Z(n25998) );
  NANDN U34780 ( .A(n23580), .B(creg[805]), .Z(n25997) );
  NAND U34781 ( .A(n25999), .B(n17860), .Z(n13546) );
  NANDN U34782 ( .A(init), .B(m[806]), .Z(n17860) );
  AND U34783 ( .A(n26000), .B(n26001), .Z(n25999) );
  NAND U34784 ( .A(o[806]), .B(n23579), .Z(n26001) );
  NANDN U34785 ( .A(n23580), .B(creg[806]), .Z(n26000) );
  NAND U34786 ( .A(n26002), .B(n17858), .Z(n13545) );
  NANDN U34787 ( .A(init), .B(m[807]), .Z(n17858) );
  AND U34788 ( .A(n26003), .B(n26004), .Z(n26002) );
  NAND U34789 ( .A(o[807]), .B(n23579), .Z(n26004) );
  NANDN U34790 ( .A(n23580), .B(creg[807]), .Z(n26003) );
  NAND U34791 ( .A(n26005), .B(n17856), .Z(n13544) );
  NANDN U34792 ( .A(init), .B(m[808]), .Z(n17856) );
  AND U34793 ( .A(n26006), .B(n26007), .Z(n26005) );
  NAND U34794 ( .A(o[808]), .B(n23579), .Z(n26007) );
  NANDN U34795 ( .A(n23580), .B(creg[808]), .Z(n26006) );
  NAND U34796 ( .A(n26008), .B(n17854), .Z(n13543) );
  NANDN U34797 ( .A(init), .B(m[809]), .Z(n17854) );
  AND U34798 ( .A(n26009), .B(n26010), .Z(n26008) );
  NAND U34799 ( .A(o[809]), .B(n23579), .Z(n26010) );
  NANDN U34800 ( .A(n23580), .B(creg[809]), .Z(n26009) );
  NAND U34801 ( .A(n26011), .B(n17850), .Z(n13542) );
  NANDN U34802 ( .A(init), .B(m[810]), .Z(n17850) );
  AND U34803 ( .A(n26012), .B(n26013), .Z(n26011) );
  NAND U34804 ( .A(o[810]), .B(n23579), .Z(n26013) );
  NANDN U34805 ( .A(n23580), .B(creg[810]), .Z(n26012) );
  NAND U34806 ( .A(n26014), .B(n17848), .Z(n13541) );
  NANDN U34807 ( .A(init), .B(m[811]), .Z(n17848) );
  AND U34808 ( .A(n26015), .B(n26016), .Z(n26014) );
  NAND U34809 ( .A(o[811]), .B(n23579), .Z(n26016) );
  NANDN U34810 ( .A(n23580), .B(creg[811]), .Z(n26015) );
  NAND U34811 ( .A(n26017), .B(n17846), .Z(n13540) );
  NANDN U34812 ( .A(init), .B(m[812]), .Z(n17846) );
  AND U34813 ( .A(n26018), .B(n26019), .Z(n26017) );
  NAND U34814 ( .A(o[812]), .B(n23579), .Z(n26019) );
  NANDN U34815 ( .A(n23580), .B(creg[812]), .Z(n26018) );
  NAND U34816 ( .A(n26020), .B(n17844), .Z(n13539) );
  NANDN U34817 ( .A(init), .B(m[813]), .Z(n17844) );
  AND U34818 ( .A(n26021), .B(n26022), .Z(n26020) );
  NAND U34819 ( .A(o[813]), .B(n23579), .Z(n26022) );
  NANDN U34820 ( .A(n23580), .B(creg[813]), .Z(n26021) );
  NAND U34821 ( .A(n26023), .B(n17842), .Z(n13538) );
  NANDN U34822 ( .A(init), .B(m[814]), .Z(n17842) );
  AND U34823 ( .A(n26024), .B(n26025), .Z(n26023) );
  NAND U34824 ( .A(o[814]), .B(n23579), .Z(n26025) );
  NANDN U34825 ( .A(n23580), .B(creg[814]), .Z(n26024) );
  NAND U34826 ( .A(n26026), .B(n17840), .Z(n13537) );
  NANDN U34827 ( .A(init), .B(m[815]), .Z(n17840) );
  AND U34828 ( .A(n26027), .B(n26028), .Z(n26026) );
  NAND U34829 ( .A(o[815]), .B(n23579), .Z(n26028) );
  NANDN U34830 ( .A(n23580), .B(creg[815]), .Z(n26027) );
  NAND U34831 ( .A(n26029), .B(n17838), .Z(n13536) );
  NANDN U34832 ( .A(init), .B(m[816]), .Z(n17838) );
  AND U34833 ( .A(n26030), .B(n26031), .Z(n26029) );
  NAND U34834 ( .A(o[816]), .B(n23579), .Z(n26031) );
  NANDN U34835 ( .A(n23580), .B(creg[816]), .Z(n26030) );
  NAND U34836 ( .A(n26032), .B(n17836), .Z(n13535) );
  NANDN U34837 ( .A(init), .B(m[817]), .Z(n17836) );
  AND U34838 ( .A(n26033), .B(n26034), .Z(n26032) );
  NAND U34839 ( .A(o[817]), .B(n23579), .Z(n26034) );
  NANDN U34840 ( .A(n23580), .B(creg[817]), .Z(n26033) );
  NAND U34841 ( .A(n26035), .B(n17834), .Z(n13534) );
  NANDN U34842 ( .A(init), .B(m[818]), .Z(n17834) );
  AND U34843 ( .A(n26036), .B(n26037), .Z(n26035) );
  NAND U34844 ( .A(o[818]), .B(n23579), .Z(n26037) );
  NANDN U34845 ( .A(n23580), .B(creg[818]), .Z(n26036) );
  NAND U34846 ( .A(n26038), .B(n17832), .Z(n13533) );
  NANDN U34847 ( .A(init), .B(m[819]), .Z(n17832) );
  AND U34848 ( .A(n26039), .B(n26040), .Z(n26038) );
  NAND U34849 ( .A(o[819]), .B(n23579), .Z(n26040) );
  NANDN U34850 ( .A(n23580), .B(creg[819]), .Z(n26039) );
  NAND U34851 ( .A(n26041), .B(n17828), .Z(n13532) );
  NANDN U34852 ( .A(init), .B(m[820]), .Z(n17828) );
  AND U34853 ( .A(n26042), .B(n26043), .Z(n26041) );
  NAND U34854 ( .A(o[820]), .B(n23579), .Z(n26043) );
  NANDN U34855 ( .A(n23580), .B(creg[820]), .Z(n26042) );
  NAND U34856 ( .A(n26044), .B(n17826), .Z(n13531) );
  NANDN U34857 ( .A(init), .B(m[821]), .Z(n17826) );
  AND U34858 ( .A(n26045), .B(n26046), .Z(n26044) );
  NAND U34859 ( .A(o[821]), .B(n23579), .Z(n26046) );
  NANDN U34860 ( .A(n23580), .B(creg[821]), .Z(n26045) );
  NAND U34861 ( .A(n26047), .B(n17824), .Z(n13530) );
  NANDN U34862 ( .A(init), .B(m[822]), .Z(n17824) );
  AND U34863 ( .A(n26048), .B(n26049), .Z(n26047) );
  NAND U34864 ( .A(o[822]), .B(n23579), .Z(n26049) );
  NANDN U34865 ( .A(n23580), .B(creg[822]), .Z(n26048) );
  NAND U34866 ( .A(n26050), .B(n17822), .Z(n13529) );
  NANDN U34867 ( .A(init), .B(m[823]), .Z(n17822) );
  AND U34868 ( .A(n26051), .B(n26052), .Z(n26050) );
  NAND U34869 ( .A(o[823]), .B(n23579), .Z(n26052) );
  NANDN U34870 ( .A(n23580), .B(creg[823]), .Z(n26051) );
  NAND U34871 ( .A(n26053), .B(n17820), .Z(n13528) );
  NANDN U34872 ( .A(init), .B(m[824]), .Z(n17820) );
  AND U34873 ( .A(n26054), .B(n26055), .Z(n26053) );
  NAND U34874 ( .A(o[824]), .B(n23579), .Z(n26055) );
  NANDN U34875 ( .A(n23580), .B(creg[824]), .Z(n26054) );
  NAND U34876 ( .A(n26056), .B(n17818), .Z(n13527) );
  NANDN U34877 ( .A(init), .B(m[825]), .Z(n17818) );
  AND U34878 ( .A(n26057), .B(n26058), .Z(n26056) );
  NAND U34879 ( .A(o[825]), .B(n23579), .Z(n26058) );
  NANDN U34880 ( .A(n23580), .B(creg[825]), .Z(n26057) );
  NAND U34881 ( .A(n26059), .B(n17816), .Z(n13526) );
  NANDN U34882 ( .A(init), .B(m[826]), .Z(n17816) );
  AND U34883 ( .A(n26060), .B(n26061), .Z(n26059) );
  NAND U34884 ( .A(o[826]), .B(n23579), .Z(n26061) );
  NANDN U34885 ( .A(n23580), .B(creg[826]), .Z(n26060) );
  NAND U34886 ( .A(n26062), .B(n17814), .Z(n13525) );
  NANDN U34887 ( .A(init), .B(m[827]), .Z(n17814) );
  AND U34888 ( .A(n26063), .B(n26064), .Z(n26062) );
  NAND U34889 ( .A(o[827]), .B(n23579), .Z(n26064) );
  NANDN U34890 ( .A(n23580), .B(creg[827]), .Z(n26063) );
  NAND U34891 ( .A(n26065), .B(n17812), .Z(n13524) );
  NANDN U34892 ( .A(init), .B(m[828]), .Z(n17812) );
  AND U34893 ( .A(n26066), .B(n26067), .Z(n26065) );
  NAND U34894 ( .A(o[828]), .B(n23579), .Z(n26067) );
  NANDN U34895 ( .A(n23580), .B(creg[828]), .Z(n26066) );
  NAND U34896 ( .A(n26068), .B(n17810), .Z(n13523) );
  NANDN U34897 ( .A(init), .B(m[829]), .Z(n17810) );
  AND U34898 ( .A(n26069), .B(n26070), .Z(n26068) );
  NAND U34899 ( .A(o[829]), .B(n23579), .Z(n26070) );
  NANDN U34900 ( .A(n23580), .B(creg[829]), .Z(n26069) );
  NAND U34901 ( .A(n26071), .B(n17806), .Z(n13522) );
  NANDN U34902 ( .A(init), .B(m[830]), .Z(n17806) );
  AND U34903 ( .A(n26072), .B(n26073), .Z(n26071) );
  NAND U34904 ( .A(o[830]), .B(n23579), .Z(n26073) );
  NANDN U34905 ( .A(n23580), .B(creg[830]), .Z(n26072) );
  NAND U34906 ( .A(n26074), .B(n17804), .Z(n13521) );
  NANDN U34907 ( .A(init), .B(m[831]), .Z(n17804) );
  AND U34908 ( .A(n26075), .B(n26076), .Z(n26074) );
  NAND U34909 ( .A(o[831]), .B(n23579), .Z(n26076) );
  NANDN U34910 ( .A(n23580), .B(creg[831]), .Z(n26075) );
  NAND U34911 ( .A(n26077), .B(n17802), .Z(n13520) );
  NANDN U34912 ( .A(init), .B(m[832]), .Z(n17802) );
  AND U34913 ( .A(n26078), .B(n26079), .Z(n26077) );
  NAND U34914 ( .A(o[832]), .B(n23579), .Z(n26079) );
  NANDN U34915 ( .A(n23580), .B(creg[832]), .Z(n26078) );
  NAND U34916 ( .A(n26080), .B(n17800), .Z(n13519) );
  NANDN U34917 ( .A(init), .B(m[833]), .Z(n17800) );
  AND U34918 ( .A(n26081), .B(n26082), .Z(n26080) );
  NAND U34919 ( .A(o[833]), .B(n23579), .Z(n26082) );
  NANDN U34920 ( .A(n23580), .B(creg[833]), .Z(n26081) );
  NAND U34921 ( .A(n26083), .B(n17798), .Z(n13518) );
  NANDN U34922 ( .A(init), .B(m[834]), .Z(n17798) );
  AND U34923 ( .A(n26084), .B(n26085), .Z(n26083) );
  NAND U34924 ( .A(o[834]), .B(n23579), .Z(n26085) );
  NANDN U34925 ( .A(n23580), .B(creg[834]), .Z(n26084) );
  NAND U34926 ( .A(n26086), .B(n17796), .Z(n13517) );
  NANDN U34927 ( .A(init), .B(m[835]), .Z(n17796) );
  AND U34928 ( .A(n26087), .B(n26088), .Z(n26086) );
  NAND U34929 ( .A(o[835]), .B(n23579), .Z(n26088) );
  NANDN U34930 ( .A(n23580), .B(creg[835]), .Z(n26087) );
  NAND U34931 ( .A(n26089), .B(n17794), .Z(n13516) );
  NANDN U34932 ( .A(init), .B(m[836]), .Z(n17794) );
  AND U34933 ( .A(n26090), .B(n26091), .Z(n26089) );
  NAND U34934 ( .A(o[836]), .B(n23579), .Z(n26091) );
  NANDN U34935 ( .A(n23580), .B(creg[836]), .Z(n26090) );
  NAND U34936 ( .A(n26092), .B(n17792), .Z(n13515) );
  NANDN U34937 ( .A(init), .B(m[837]), .Z(n17792) );
  AND U34938 ( .A(n26093), .B(n26094), .Z(n26092) );
  NAND U34939 ( .A(o[837]), .B(n23579), .Z(n26094) );
  NANDN U34940 ( .A(n23580), .B(creg[837]), .Z(n26093) );
  NAND U34941 ( .A(n26095), .B(n17790), .Z(n13514) );
  NANDN U34942 ( .A(init), .B(m[838]), .Z(n17790) );
  AND U34943 ( .A(n26096), .B(n26097), .Z(n26095) );
  NAND U34944 ( .A(o[838]), .B(n23579), .Z(n26097) );
  NANDN U34945 ( .A(n23580), .B(creg[838]), .Z(n26096) );
  NAND U34946 ( .A(n26098), .B(n17788), .Z(n13513) );
  NANDN U34947 ( .A(init), .B(m[839]), .Z(n17788) );
  AND U34948 ( .A(n26099), .B(n26100), .Z(n26098) );
  NAND U34949 ( .A(o[839]), .B(n23579), .Z(n26100) );
  NANDN U34950 ( .A(n23580), .B(creg[839]), .Z(n26099) );
  NAND U34951 ( .A(n26101), .B(n17784), .Z(n13512) );
  NANDN U34952 ( .A(init), .B(m[840]), .Z(n17784) );
  AND U34953 ( .A(n26102), .B(n26103), .Z(n26101) );
  NAND U34954 ( .A(o[840]), .B(n23579), .Z(n26103) );
  NANDN U34955 ( .A(n23580), .B(creg[840]), .Z(n26102) );
  NAND U34956 ( .A(n26104), .B(n17782), .Z(n13511) );
  NANDN U34957 ( .A(init), .B(m[841]), .Z(n17782) );
  AND U34958 ( .A(n26105), .B(n26106), .Z(n26104) );
  NAND U34959 ( .A(o[841]), .B(n23579), .Z(n26106) );
  NANDN U34960 ( .A(n23580), .B(creg[841]), .Z(n26105) );
  NAND U34961 ( .A(n26107), .B(n17780), .Z(n13510) );
  NANDN U34962 ( .A(init), .B(m[842]), .Z(n17780) );
  AND U34963 ( .A(n26108), .B(n26109), .Z(n26107) );
  NAND U34964 ( .A(o[842]), .B(n23579), .Z(n26109) );
  NANDN U34965 ( .A(n23580), .B(creg[842]), .Z(n26108) );
  NAND U34966 ( .A(n26110), .B(n17778), .Z(n13509) );
  NANDN U34967 ( .A(init), .B(m[843]), .Z(n17778) );
  AND U34968 ( .A(n26111), .B(n26112), .Z(n26110) );
  NAND U34969 ( .A(o[843]), .B(n23579), .Z(n26112) );
  NANDN U34970 ( .A(n23580), .B(creg[843]), .Z(n26111) );
  NAND U34971 ( .A(n26113), .B(n17776), .Z(n13508) );
  NANDN U34972 ( .A(init), .B(m[844]), .Z(n17776) );
  AND U34973 ( .A(n26114), .B(n26115), .Z(n26113) );
  NAND U34974 ( .A(o[844]), .B(n23579), .Z(n26115) );
  NANDN U34975 ( .A(n23580), .B(creg[844]), .Z(n26114) );
  NAND U34976 ( .A(n26116), .B(n17774), .Z(n13507) );
  NANDN U34977 ( .A(init), .B(m[845]), .Z(n17774) );
  AND U34978 ( .A(n26117), .B(n26118), .Z(n26116) );
  NAND U34979 ( .A(o[845]), .B(n23579), .Z(n26118) );
  NANDN U34980 ( .A(n23580), .B(creg[845]), .Z(n26117) );
  NAND U34981 ( .A(n26119), .B(n17772), .Z(n13506) );
  NANDN U34982 ( .A(init), .B(m[846]), .Z(n17772) );
  AND U34983 ( .A(n26120), .B(n26121), .Z(n26119) );
  NAND U34984 ( .A(o[846]), .B(n23579), .Z(n26121) );
  NANDN U34985 ( .A(n23580), .B(creg[846]), .Z(n26120) );
  NAND U34986 ( .A(n26122), .B(n17770), .Z(n13505) );
  NANDN U34987 ( .A(init), .B(m[847]), .Z(n17770) );
  AND U34988 ( .A(n26123), .B(n26124), .Z(n26122) );
  NAND U34989 ( .A(o[847]), .B(n23579), .Z(n26124) );
  NANDN U34990 ( .A(n23580), .B(creg[847]), .Z(n26123) );
  NAND U34991 ( .A(n26125), .B(n17768), .Z(n13504) );
  NANDN U34992 ( .A(init), .B(m[848]), .Z(n17768) );
  AND U34993 ( .A(n26126), .B(n26127), .Z(n26125) );
  NAND U34994 ( .A(o[848]), .B(n23579), .Z(n26127) );
  NANDN U34995 ( .A(n23580), .B(creg[848]), .Z(n26126) );
  NAND U34996 ( .A(n26128), .B(n17766), .Z(n13503) );
  NANDN U34997 ( .A(init), .B(m[849]), .Z(n17766) );
  AND U34998 ( .A(n26129), .B(n26130), .Z(n26128) );
  NAND U34999 ( .A(o[849]), .B(n23579), .Z(n26130) );
  NANDN U35000 ( .A(n23580), .B(creg[849]), .Z(n26129) );
  NAND U35001 ( .A(n26131), .B(n17762), .Z(n13502) );
  NANDN U35002 ( .A(init), .B(m[850]), .Z(n17762) );
  AND U35003 ( .A(n26132), .B(n26133), .Z(n26131) );
  NAND U35004 ( .A(o[850]), .B(n23579), .Z(n26133) );
  NANDN U35005 ( .A(n23580), .B(creg[850]), .Z(n26132) );
  NAND U35006 ( .A(n26134), .B(n17760), .Z(n13501) );
  NANDN U35007 ( .A(init), .B(m[851]), .Z(n17760) );
  AND U35008 ( .A(n26135), .B(n26136), .Z(n26134) );
  NAND U35009 ( .A(o[851]), .B(n23579), .Z(n26136) );
  NANDN U35010 ( .A(n23580), .B(creg[851]), .Z(n26135) );
  NAND U35011 ( .A(n26137), .B(n17758), .Z(n13500) );
  NANDN U35012 ( .A(init), .B(m[852]), .Z(n17758) );
  AND U35013 ( .A(n26138), .B(n26139), .Z(n26137) );
  NAND U35014 ( .A(o[852]), .B(n23579), .Z(n26139) );
  NANDN U35015 ( .A(n23580), .B(creg[852]), .Z(n26138) );
  NAND U35016 ( .A(n26140), .B(n17756), .Z(n13499) );
  NANDN U35017 ( .A(init), .B(m[853]), .Z(n17756) );
  AND U35018 ( .A(n26141), .B(n26142), .Z(n26140) );
  NAND U35019 ( .A(o[853]), .B(n23579), .Z(n26142) );
  NANDN U35020 ( .A(n23580), .B(creg[853]), .Z(n26141) );
  NAND U35021 ( .A(n26143), .B(n17754), .Z(n13498) );
  NANDN U35022 ( .A(init), .B(m[854]), .Z(n17754) );
  AND U35023 ( .A(n26144), .B(n26145), .Z(n26143) );
  NAND U35024 ( .A(o[854]), .B(n23579), .Z(n26145) );
  NANDN U35025 ( .A(n23580), .B(creg[854]), .Z(n26144) );
  NAND U35026 ( .A(n26146), .B(n17752), .Z(n13497) );
  NANDN U35027 ( .A(init), .B(m[855]), .Z(n17752) );
  AND U35028 ( .A(n26147), .B(n26148), .Z(n26146) );
  NAND U35029 ( .A(o[855]), .B(n23579), .Z(n26148) );
  NANDN U35030 ( .A(n23580), .B(creg[855]), .Z(n26147) );
  NAND U35031 ( .A(n26149), .B(n17750), .Z(n13496) );
  NANDN U35032 ( .A(init), .B(m[856]), .Z(n17750) );
  AND U35033 ( .A(n26150), .B(n26151), .Z(n26149) );
  NAND U35034 ( .A(o[856]), .B(n23579), .Z(n26151) );
  NANDN U35035 ( .A(n23580), .B(creg[856]), .Z(n26150) );
  NAND U35036 ( .A(n26152), .B(n17748), .Z(n13495) );
  NANDN U35037 ( .A(init), .B(m[857]), .Z(n17748) );
  AND U35038 ( .A(n26153), .B(n26154), .Z(n26152) );
  NAND U35039 ( .A(o[857]), .B(n23579), .Z(n26154) );
  NANDN U35040 ( .A(n23580), .B(creg[857]), .Z(n26153) );
  NAND U35041 ( .A(n26155), .B(n17746), .Z(n13494) );
  NANDN U35042 ( .A(init), .B(m[858]), .Z(n17746) );
  AND U35043 ( .A(n26156), .B(n26157), .Z(n26155) );
  NAND U35044 ( .A(o[858]), .B(n23579), .Z(n26157) );
  NANDN U35045 ( .A(n23580), .B(creg[858]), .Z(n26156) );
  NAND U35046 ( .A(n26158), .B(n17744), .Z(n13493) );
  NANDN U35047 ( .A(init), .B(m[859]), .Z(n17744) );
  AND U35048 ( .A(n26159), .B(n26160), .Z(n26158) );
  NAND U35049 ( .A(o[859]), .B(n23579), .Z(n26160) );
  NANDN U35050 ( .A(n23580), .B(creg[859]), .Z(n26159) );
  NAND U35051 ( .A(n26161), .B(n17740), .Z(n13492) );
  NANDN U35052 ( .A(init), .B(m[860]), .Z(n17740) );
  AND U35053 ( .A(n26162), .B(n26163), .Z(n26161) );
  NAND U35054 ( .A(o[860]), .B(n23579), .Z(n26163) );
  NANDN U35055 ( .A(n23580), .B(creg[860]), .Z(n26162) );
  NAND U35056 ( .A(n26164), .B(n17738), .Z(n13491) );
  NANDN U35057 ( .A(init), .B(m[861]), .Z(n17738) );
  AND U35058 ( .A(n26165), .B(n26166), .Z(n26164) );
  NAND U35059 ( .A(o[861]), .B(n23579), .Z(n26166) );
  NANDN U35060 ( .A(n23580), .B(creg[861]), .Z(n26165) );
  NAND U35061 ( .A(n26167), .B(n17736), .Z(n13490) );
  NANDN U35062 ( .A(init), .B(m[862]), .Z(n17736) );
  AND U35063 ( .A(n26168), .B(n26169), .Z(n26167) );
  NAND U35064 ( .A(o[862]), .B(n23579), .Z(n26169) );
  NANDN U35065 ( .A(n23580), .B(creg[862]), .Z(n26168) );
  NAND U35066 ( .A(n26170), .B(n17734), .Z(n13489) );
  NANDN U35067 ( .A(init), .B(m[863]), .Z(n17734) );
  AND U35068 ( .A(n26171), .B(n26172), .Z(n26170) );
  NAND U35069 ( .A(o[863]), .B(n23579), .Z(n26172) );
  NANDN U35070 ( .A(n23580), .B(creg[863]), .Z(n26171) );
  NAND U35071 ( .A(n26173), .B(n17732), .Z(n13488) );
  NANDN U35072 ( .A(init), .B(m[864]), .Z(n17732) );
  AND U35073 ( .A(n26174), .B(n26175), .Z(n26173) );
  NAND U35074 ( .A(o[864]), .B(n23579), .Z(n26175) );
  NANDN U35075 ( .A(n23580), .B(creg[864]), .Z(n26174) );
  NAND U35076 ( .A(n26176), .B(n17730), .Z(n13487) );
  NANDN U35077 ( .A(init), .B(m[865]), .Z(n17730) );
  AND U35078 ( .A(n26177), .B(n26178), .Z(n26176) );
  NAND U35079 ( .A(o[865]), .B(n23579), .Z(n26178) );
  NANDN U35080 ( .A(n23580), .B(creg[865]), .Z(n26177) );
  NAND U35081 ( .A(n26179), .B(n17728), .Z(n13486) );
  NANDN U35082 ( .A(init), .B(m[866]), .Z(n17728) );
  AND U35083 ( .A(n26180), .B(n26181), .Z(n26179) );
  NAND U35084 ( .A(o[866]), .B(n23579), .Z(n26181) );
  NANDN U35085 ( .A(n23580), .B(creg[866]), .Z(n26180) );
  NAND U35086 ( .A(n26182), .B(n17726), .Z(n13485) );
  NANDN U35087 ( .A(init), .B(m[867]), .Z(n17726) );
  AND U35088 ( .A(n26183), .B(n26184), .Z(n26182) );
  NAND U35089 ( .A(o[867]), .B(n23579), .Z(n26184) );
  NANDN U35090 ( .A(n23580), .B(creg[867]), .Z(n26183) );
  NAND U35091 ( .A(n26185), .B(n17724), .Z(n13484) );
  NANDN U35092 ( .A(init), .B(m[868]), .Z(n17724) );
  AND U35093 ( .A(n26186), .B(n26187), .Z(n26185) );
  NAND U35094 ( .A(o[868]), .B(n23579), .Z(n26187) );
  NANDN U35095 ( .A(n23580), .B(creg[868]), .Z(n26186) );
  NAND U35096 ( .A(n26188), .B(n17722), .Z(n13483) );
  NANDN U35097 ( .A(init), .B(m[869]), .Z(n17722) );
  AND U35098 ( .A(n26189), .B(n26190), .Z(n26188) );
  NAND U35099 ( .A(o[869]), .B(n23579), .Z(n26190) );
  NANDN U35100 ( .A(n23580), .B(creg[869]), .Z(n26189) );
  NAND U35101 ( .A(n26191), .B(n17718), .Z(n13482) );
  NANDN U35102 ( .A(init), .B(m[870]), .Z(n17718) );
  AND U35103 ( .A(n26192), .B(n26193), .Z(n26191) );
  NAND U35104 ( .A(o[870]), .B(n23579), .Z(n26193) );
  NANDN U35105 ( .A(n23580), .B(creg[870]), .Z(n26192) );
  NAND U35106 ( .A(n26194), .B(n17716), .Z(n13481) );
  NANDN U35107 ( .A(init), .B(m[871]), .Z(n17716) );
  AND U35108 ( .A(n26195), .B(n26196), .Z(n26194) );
  NAND U35109 ( .A(o[871]), .B(n23579), .Z(n26196) );
  NANDN U35110 ( .A(n23580), .B(creg[871]), .Z(n26195) );
  NAND U35111 ( .A(n26197), .B(n17714), .Z(n13480) );
  NANDN U35112 ( .A(init), .B(m[872]), .Z(n17714) );
  AND U35113 ( .A(n26198), .B(n26199), .Z(n26197) );
  NAND U35114 ( .A(o[872]), .B(n23579), .Z(n26199) );
  NANDN U35115 ( .A(n23580), .B(creg[872]), .Z(n26198) );
  NAND U35116 ( .A(n26200), .B(n17712), .Z(n13479) );
  NANDN U35117 ( .A(init), .B(m[873]), .Z(n17712) );
  AND U35118 ( .A(n26201), .B(n26202), .Z(n26200) );
  NAND U35119 ( .A(o[873]), .B(n23579), .Z(n26202) );
  NANDN U35120 ( .A(n23580), .B(creg[873]), .Z(n26201) );
  NAND U35121 ( .A(n26203), .B(n17710), .Z(n13478) );
  NANDN U35122 ( .A(init), .B(m[874]), .Z(n17710) );
  AND U35123 ( .A(n26204), .B(n26205), .Z(n26203) );
  NAND U35124 ( .A(o[874]), .B(n23579), .Z(n26205) );
  NANDN U35125 ( .A(n23580), .B(creg[874]), .Z(n26204) );
  NAND U35126 ( .A(n26206), .B(n17708), .Z(n13477) );
  NANDN U35127 ( .A(init), .B(m[875]), .Z(n17708) );
  AND U35128 ( .A(n26207), .B(n26208), .Z(n26206) );
  NAND U35129 ( .A(o[875]), .B(n23579), .Z(n26208) );
  NANDN U35130 ( .A(n23580), .B(creg[875]), .Z(n26207) );
  NAND U35131 ( .A(n26209), .B(n17706), .Z(n13476) );
  NANDN U35132 ( .A(init), .B(m[876]), .Z(n17706) );
  AND U35133 ( .A(n26210), .B(n26211), .Z(n26209) );
  NAND U35134 ( .A(o[876]), .B(n23579), .Z(n26211) );
  NANDN U35135 ( .A(n23580), .B(creg[876]), .Z(n26210) );
  NAND U35136 ( .A(n26212), .B(n17704), .Z(n13475) );
  NANDN U35137 ( .A(init), .B(m[877]), .Z(n17704) );
  AND U35138 ( .A(n26213), .B(n26214), .Z(n26212) );
  NAND U35139 ( .A(o[877]), .B(n23579), .Z(n26214) );
  NANDN U35140 ( .A(n23580), .B(creg[877]), .Z(n26213) );
  NAND U35141 ( .A(n26215), .B(n17702), .Z(n13474) );
  NANDN U35142 ( .A(init), .B(m[878]), .Z(n17702) );
  AND U35143 ( .A(n26216), .B(n26217), .Z(n26215) );
  NAND U35144 ( .A(o[878]), .B(n23579), .Z(n26217) );
  NANDN U35145 ( .A(n23580), .B(creg[878]), .Z(n26216) );
  NAND U35146 ( .A(n26218), .B(n17700), .Z(n13473) );
  NANDN U35147 ( .A(init), .B(m[879]), .Z(n17700) );
  AND U35148 ( .A(n26219), .B(n26220), .Z(n26218) );
  NAND U35149 ( .A(o[879]), .B(n23579), .Z(n26220) );
  NANDN U35150 ( .A(n23580), .B(creg[879]), .Z(n26219) );
  NAND U35151 ( .A(n26221), .B(n17696), .Z(n13472) );
  NANDN U35152 ( .A(init), .B(m[880]), .Z(n17696) );
  AND U35153 ( .A(n26222), .B(n26223), .Z(n26221) );
  NAND U35154 ( .A(o[880]), .B(n23579), .Z(n26223) );
  NANDN U35155 ( .A(n23580), .B(creg[880]), .Z(n26222) );
  NAND U35156 ( .A(n26224), .B(n17694), .Z(n13471) );
  NANDN U35157 ( .A(init), .B(m[881]), .Z(n17694) );
  AND U35158 ( .A(n26225), .B(n26226), .Z(n26224) );
  NAND U35159 ( .A(o[881]), .B(n23579), .Z(n26226) );
  NANDN U35160 ( .A(n23580), .B(creg[881]), .Z(n26225) );
  NAND U35161 ( .A(n26227), .B(n17692), .Z(n13470) );
  NANDN U35162 ( .A(init), .B(m[882]), .Z(n17692) );
  AND U35163 ( .A(n26228), .B(n26229), .Z(n26227) );
  NAND U35164 ( .A(o[882]), .B(n23579), .Z(n26229) );
  NANDN U35165 ( .A(n23580), .B(creg[882]), .Z(n26228) );
  NAND U35166 ( .A(n26230), .B(n17690), .Z(n13469) );
  NANDN U35167 ( .A(init), .B(m[883]), .Z(n17690) );
  AND U35168 ( .A(n26231), .B(n26232), .Z(n26230) );
  NAND U35169 ( .A(o[883]), .B(n23579), .Z(n26232) );
  NANDN U35170 ( .A(n23580), .B(creg[883]), .Z(n26231) );
  NAND U35171 ( .A(n26233), .B(n17688), .Z(n13468) );
  NANDN U35172 ( .A(init), .B(m[884]), .Z(n17688) );
  AND U35173 ( .A(n26234), .B(n26235), .Z(n26233) );
  NAND U35174 ( .A(o[884]), .B(n23579), .Z(n26235) );
  NANDN U35175 ( .A(n23580), .B(creg[884]), .Z(n26234) );
  NAND U35176 ( .A(n26236), .B(n17686), .Z(n13467) );
  NANDN U35177 ( .A(init), .B(m[885]), .Z(n17686) );
  AND U35178 ( .A(n26237), .B(n26238), .Z(n26236) );
  NAND U35179 ( .A(o[885]), .B(n23579), .Z(n26238) );
  NANDN U35180 ( .A(n23580), .B(creg[885]), .Z(n26237) );
  NAND U35181 ( .A(n26239), .B(n17684), .Z(n13466) );
  NANDN U35182 ( .A(init), .B(m[886]), .Z(n17684) );
  AND U35183 ( .A(n26240), .B(n26241), .Z(n26239) );
  NAND U35184 ( .A(o[886]), .B(n23579), .Z(n26241) );
  NANDN U35185 ( .A(n23580), .B(creg[886]), .Z(n26240) );
  NAND U35186 ( .A(n26242), .B(n17682), .Z(n13465) );
  NANDN U35187 ( .A(init), .B(m[887]), .Z(n17682) );
  AND U35188 ( .A(n26243), .B(n26244), .Z(n26242) );
  NAND U35189 ( .A(o[887]), .B(n23579), .Z(n26244) );
  NANDN U35190 ( .A(n23580), .B(creg[887]), .Z(n26243) );
  NAND U35191 ( .A(n26245), .B(n17680), .Z(n13464) );
  NANDN U35192 ( .A(init), .B(m[888]), .Z(n17680) );
  AND U35193 ( .A(n26246), .B(n26247), .Z(n26245) );
  NAND U35194 ( .A(o[888]), .B(n23579), .Z(n26247) );
  NANDN U35195 ( .A(n23580), .B(creg[888]), .Z(n26246) );
  NAND U35196 ( .A(n26248), .B(n17678), .Z(n13463) );
  NANDN U35197 ( .A(init), .B(m[889]), .Z(n17678) );
  AND U35198 ( .A(n26249), .B(n26250), .Z(n26248) );
  NAND U35199 ( .A(o[889]), .B(n23579), .Z(n26250) );
  NANDN U35200 ( .A(n23580), .B(creg[889]), .Z(n26249) );
  NAND U35201 ( .A(n26251), .B(n17674), .Z(n13462) );
  NANDN U35202 ( .A(init), .B(m[890]), .Z(n17674) );
  AND U35203 ( .A(n26252), .B(n26253), .Z(n26251) );
  NAND U35204 ( .A(o[890]), .B(n23579), .Z(n26253) );
  NANDN U35205 ( .A(n23580), .B(creg[890]), .Z(n26252) );
  NAND U35206 ( .A(n26254), .B(n17672), .Z(n13461) );
  NANDN U35207 ( .A(init), .B(m[891]), .Z(n17672) );
  AND U35208 ( .A(n26255), .B(n26256), .Z(n26254) );
  NAND U35209 ( .A(o[891]), .B(n23579), .Z(n26256) );
  NANDN U35210 ( .A(n23580), .B(creg[891]), .Z(n26255) );
  NAND U35211 ( .A(n26257), .B(n17670), .Z(n13460) );
  NANDN U35212 ( .A(init), .B(m[892]), .Z(n17670) );
  AND U35213 ( .A(n26258), .B(n26259), .Z(n26257) );
  NAND U35214 ( .A(o[892]), .B(n23579), .Z(n26259) );
  NANDN U35215 ( .A(n23580), .B(creg[892]), .Z(n26258) );
  NAND U35216 ( .A(n26260), .B(n17668), .Z(n13459) );
  NANDN U35217 ( .A(init), .B(m[893]), .Z(n17668) );
  AND U35218 ( .A(n26261), .B(n26262), .Z(n26260) );
  NAND U35219 ( .A(o[893]), .B(n23579), .Z(n26262) );
  NANDN U35220 ( .A(n23580), .B(creg[893]), .Z(n26261) );
  NAND U35221 ( .A(n26263), .B(n17666), .Z(n13458) );
  NANDN U35222 ( .A(init), .B(m[894]), .Z(n17666) );
  AND U35223 ( .A(n26264), .B(n26265), .Z(n26263) );
  NAND U35224 ( .A(o[894]), .B(n23579), .Z(n26265) );
  NANDN U35225 ( .A(n23580), .B(creg[894]), .Z(n26264) );
  NAND U35226 ( .A(n26266), .B(n17664), .Z(n13457) );
  NANDN U35227 ( .A(init), .B(m[895]), .Z(n17664) );
  AND U35228 ( .A(n26267), .B(n26268), .Z(n26266) );
  NAND U35229 ( .A(o[895]), .B(n23579), .Z(n26268) );
  NANDN U35230 ( .A(n23580), .B(creg[895]), .Z(n26267) );
  NAND U35231 ( .A(n26269), .B(n17662), .Z(n13456) );
  NANDN U35232 ( .A(init), .B(m[896]), .Z(n17662) );
  AND U35233 ( .A(n26270), .B(n26271), .Z(n26269) );
  NAND U35234 ( .A(o[896]), .B(n23579), .Z(n26271) );
  NANDN U35235 ( .A(n23580), .B(creg[896]), .Z(n26270) );
  NAND U35236 ( .A(n26272), .B(n17660), .Z(n13455) );
  NANDN U35237 ( .A(init), .B(m[897]), .Z(n17660) );
  AND U35238 ( .A(n26273), .B(n26274), .Z(n26272) );
  NAND U35239 ( .A(o[897]), .B(n23579), .Z(n26274) );
  NANDN U35240 ( .A(n23580), .B(creg[897]), .Z(n26273) );
  NAND U35241 ( .A(n26275), .B(n17658), .Z(n13454) );
  NANDN U35242 ( .A(init), .B(m[898]), .Z(n17658) );
  AND U35243 ( .A(n26276), .B(n26277), .Z(n26275) );
  NAND U35244 ( .A(o[898]), .B(n23579), .Z(n26277) );
  NANDN U35245 ( .A(n23580), .B(creg[898]), .Z(n26276) );
  NAND U35246 ( .A(n26278), .B(n17656), .Z(n13453) );
  NANDN U35247 ( .A(init), .B(m[899]), .Z(n17656) );
  AND U35248 ( .A(n26279), .B(n26280), .Z(n26278) );
  NAND U35249 ( .A(o[899]), .B(n23579), .Z(n26280) );
  NANDN U35250 ( .A(n23580), .B(creg[899]), .Z(n26279) );
  NAND U35251 ( .A(n26281), .B(n17650), .Z(n13452) );
  NANDN U35252 ( .A(init), .B(m[900]), .Z(n17650) );
  AND U35253 ( .A(n26282), .B(n26283), .Z(n26281) );
  NAND U35254 ( .A(o[900]), .B(n23579), .Z(n26283) );
  NANDN U35255 ( .A(n23580), .B(creg[900]), .Z(n26282) );
  NAND U35256 ( .A(n26284), .B(n17648), .Z(n13451) );
  NANDN U35257 ( .A(init), .B(m[901]), .Z(n17648) );
  AND U35258 ( .A(n26285), .B(n26286), .Z(n26284) );
  NAND U35259 ( .A(o[901]), .B(n23579), .Z(n26286) );
  NANDN U35260 ( .A(n23580), .B(creg[901]), .Z(n26285) );
  NAND U35261 ( .A(n26287), .B(n17646), .Z(n13450) );
  NANDN U35262 ( .A(init), .B(m[902]), .Z(n17646) );
  AND U35263 ( .A(n26288), .B(n26289), .Z(n26287) );
  NAND U35264 ( .A(o[902]), .B(n23579), .Z(n26289) );
  NANDN U35265 ( .A(n23580), .B(creg[902]), .Z(n26288) );
  NAND U35266 ( .A(n26290), .B(n17644), .Z(n13449) );
  NANDN U35267 ( .A(init), .B(m[903]), .Z(n17644) );
  AND U35268 ( .A(n26291), .B(n26292), .Z(n26290) );
  NAND U35269 ( .A(o[903]), .B(n23579), .Z(n26292) );
  NANDN U35270 ( .A(n23580), .B(creg[903]), .Z(n26291) );
  NAND U35271 ( .A(n26293), .B(n17642), .Z(n13448) );
  NANDN U35272 ( .A(init), .B(m[904]), .Z(n17642) );
  AND U35273 ( .A(n26294), .B(n26295), .Z(n26293) );
  NAND U35274 ( .A(o[904]), .B(n23579), .Z(n26295) );
  NANDN U35275 ( .A(n23580), .B(creg[904]), .Z(n26294) );
  NAND U35276 ( .A(n26296), .B(n17640), .Z(n13447) );
  NANDN U35277 ( .A(init), .B(m[905]), .Z(n17640) );
  AND U35278 ( .A(n26297), .B(n26298), .Z(n26296) );
  NAND U35279 ( .A(o[905]), .B(n23579), .Z(n26298) );
  NANDN U35280 ( .A(n23580), .B(creg[905]), .Z(n26297) );
  NAND U35281 ( .A(n26299), .B(n17638), .Z(n13446) );
  NANDN U35282 ( .A(init), .B(m[906]), .Z(n17638) );
  AND U35283 ( .A(n26300), .B(n26301), .Z(n26299) );
  NAND U35284 ( .A(o[906]), .B(n23579), .Z(n26301) );
  NANDN U35285 ( .A(n23580), .B(creg[906]), .Z(n26300) );
  NAND U35286 ( .A(n26302), .B(n17636), .Z(n13445) );
  NANDN U35287 ( .A(init), .B(m[907]), .Z(n17636) );
  AND U35288 ( .A(n26303), .B(n26304), .Z(n26302) );
  NAND U35289 ( .A(o[907]), .B(n23579), .Z(n26304) );
  NANDN U35290 ( .A(n23580), .B(creg[907]), .Z(n26303) );
  NAND U35291 ( .A(n26305), .B(n17634), .Z(n13444) );
  NANDN U35292 ( .A(init), .B(m[908]), .Z(n17634) );
  AND U35293 ( .A(n26306), .B(n26307), .Z(n26305) );
  NAND U35294 ( .A(o[908]), .B(n23579), .Z(n26307) );
  NANDN U35295 ( .A(n23580), .B(creg[908]), .Z(n26306) );
  NAND U35296 ( .A(n26308), .B(n17632), .Z(n13443) );
  NANDN U35297 ( .A(init), .B(m[909]), .Z(n17632) );
  AND U35298 ( .A(n26309), .B(n26310), .Z(n26308) );
  NAND U35299 ( .A(o[909]), .B(n23579), .Z(n26310) );
  NANDN U35300 ( .A(n23580), .B(creg[909]), .Z(n26309) );
  NAND U35301 ( .A(n26311), .B(n17628), .Z(n13442) );
  NANDN U35302 ( .A(init), .B(m[910]), .Z(n17628) );
  AND U35303 ( .A(n26312), .B(n26313), .Z(n26311) );
  NAND U35304 ( .A(o[910]), .B(n23579), .Z(n26313) );
  NANDN U35305 ( .A(n23580), .B(creg[910]), .Z(n26312) );
  NAND U35306 ( .A(n26314), .B(n17626), .Z(n13441) );
  NANDN U35307 ( .A(init), .B(m[911]), .Z(n17626) );
  AND U35308 ( .A(n26315), .B(n26316), .Z(n26314) );
  NAND U35309 ( .A(o[911]), .B(n23579), .Z(n26316) );
  NANDN U35310 ( .A(n23580), .B(creg[911]), .Z(n26315) );
  NAND U35311 ( .A(n26317), .B(n17624), .Z(n13440) );
  NANDN U35312 ( .A(init), .B(m[912]), .Z(n17624) );
  AND U35313 ( .A(n26318), .B(n26319), .Z(n26317) );
  NAND U35314 ( .A(o[912]), .B(n23579), .Z(n26319) );
  NANDN U35315 ( .A(n23580), .B(creg[912]), .Z(n26318) );
  NAND U35316 ( .A(n26320), .B(n17622), .Z(n13439) );
  NANDN U35317 ( .A(init), .B(m[913]), .Z(n17622) );
  AND U35318 ( .A(n26321), .B(n26322), .Z(n26320) );
  NAND U35319 ( .A(o[913]), .B(n23579), .Z(n26322) );
  NANDN U35320 ( .A(n23580), .B(creg[913]), .Z(n26321) );
  NAND U35321 ( .A(n26323), .B(n17620), .Z(n13438) );
  NANDN U35322 ( .A(init), .B(m[914]), .Z(n17620) );
  AND U35323 ( .A(n26324), .B(n26325), .Z(n26323) );
  NAND U35324 ( .A(o[914]), .B(n23579), .Z(n26325) );
  NANDN U35325 ( .A(n23580), .B(creg[914]), .Z(n26324) );
  NAND U35326 ( .A(n26326), .B(n17618), .Z(n13437) );
  NANDN U35327 ( .A(init), .B(m[915]), .Z(n17618) );
  AND U35328 ( .A(n26327), .B(n26328), .Z(n26326) );
  NAND U35329 ( .A(o[915]), .B(n23579), .Z(n26328) );
  NANDN U35330 ( .A(n23580), .B(creg[915]), .Z(n26327) );
  NAND U35331 ( .A(n26329), .B(n17616), .Z(n13436) );
  NANDN U35332 ( .A(init), .B(m[916]), .Z(n17616) );
  AND U35333 ( .A(n26330), .B(n26331), .Z(n26329) );
  NAND U35334 ( .A(o[916]), .B(n23579), .Z(n26331) );
  NANDN U35335 ( .A(n23580), .B(creg[916]), .Z(n26330) );
  NAND U35336 ( .A(n26332), .B(n17614), .Z(n13435) );
  NANDN U35337 ( .A(init), .B(m[917]), .Z(n17614) );
  AND U35338 ( .A(n26333), .B(n26334), .Z(n26332) );
  NAND U35339 ( .A(o[917]), .B(n23579), .Z(n26334) );
  NANDN U35340 ( .A(n23580), .B(creg[917]), .Z(n26333) );
  NAND U35341 ( .A(n26335), .B(n17612), .Z(n13434) );
  NANDN U35342 ( .A(init), .B(m[918]), .Z(n17612) );
  AND U35343 ( .A(n26336), .B(n26337), .Z(n26335) );
  NAND U35344 ( .A(o[918]), .B(n23579), .Z(n26337) );
  NANDN U35345 ( .A(n23580), .B(creg[918]), .Z(n26336) );
  NAND U35346 ( .A(n26338), .B(n17610), .Z(n13433) );
  NANDN U35347 ( .A(init), .B(m[919]), .Z(n17610) );
  AND U35348 ( .A(n26339), .B(n26340), .Z(n26338) );
  NAND U35349 ( .A(o[919]), .B(n23579), .Z(n26340) );
  NANDN U35350 ( .A(n23580), .B(creg[919]), .Z(n26339) );
  NAND U35351 ( .A(n26341), .B(n17606), .Z(n13432) );
  NANDN U35352 ( .A(init), .B(m[920]), .Z(n17606) );
  AND U35353 ( .A(n26342), .B(n26343), .Z(n26341) );
  NAND U35354 ( .A(o[920]), .B(n23579), .Z(n26343) );
  NANDN U35355 ( .A(n23580), .B(creg[920]), .Z(n26342) );
  NAND U35356 ( .A(n26344), .B(n17604), .Z(n13431) );
  NANDN U35357 ( .A(init), .B(m[921]), .Z(n17604) );
  AND U35358 ( .A(n26345), .B(n26346), .Z(n26344) );
  NAND U35359 ( .A(o[921]), .B(n23579), .Z(n26346) );
  NANDN U35360 ( .A(n23580), .B(creg[921]), .Z(n26345) );
  NAND U35361 ( .A(n26347), .B(n17602), .Z(n13430) );
  NANDN U35362 ( .A(init), .B(m[922]), .Z(n17602) );
  AND U35363 ( .A(n26348), .B(n26349), .Z(n26347) );
  NAND U35364 ( .A(o[922]), .B(n23579), .Z(n26349) );
  NANDN U35365 ( .A(n23580), .B(creg[922]), .Z(n26348) );
  NAND U35366 ( .A(n26350), .B(n17600), .Z(n13429) );
  NANDN U35367 ( .A(init), .B(m[923]), .Z(n17600) );
  AND U35368 ( .A(n26351), .B(n26352), .Z(n26350) );
  NAND U35369 ( .A(o[923]), .B(n23579), .Z(n26352) );
  NANDN U35370 ( .A(n23580), .B(creg[923]), .Z(n26351) );
  NAND U35371 ( .A(n26353), .B(n17598), .Z(n13428) );
  NANDN U35372 ( .A(init), .B(m[924]), .Z(n17598) );
  AND U35373 ( .A(n26354), .B(n26355), .Z(n26353) );
  NAND U35374 ( .A(o[924]), .B(n23579), .Z(n26355) );
  NANDN U35375 ( .A(n23580), .B(creg[924]), .Z(n26354) );
  NAND U35376 ( .A(n26356), .B(n17596), .Z(n13427) );
  NANDN U35377 ( .A(init), .B(m[925]), .Z(n17596) );
  AND U35378 ( .A(n26357), .B(n26358), .Z(n26356) );
  NAND U35379 ( .A(o[925]), .B(n23579), .Z(n26358) );
  NANDN U35380 ( .A(n23580), .B(creg[925]), .Z(n26357) );
  NAND U35381 ( .A(n26359), .B(n17594), .Z(n13426) );
  NANDN U35382 ( .A(init), .B(m[926]), .Z(n17594) );
  AND U35383 ( .A(n26360), .B(n26361), .Z(n26359) );
  NAND U35384 ( .A(o[926]), .B(n23579), .Z(n26361) );
  NANDN U35385 ( .A(n23580), .B(creg[926]), .Z(n26360) );
  NAND U35386 ( .A(n26362), .B(n17592), .Z(n13425) );
  NANDN U35387 ( .A(init), .B(m[927]), .Z(n17592) );
  AND U35388 ( .A(n26363), .B(n26364), .Z(n26362) );
  NAND U35389 ( .A(o[927]), .B(n23579), .Z(n26364) );
  NANDN U35390 ( .A(n23580), .B(creg[927]), .Z(n26363) );
  NAND U35391 ( .A(n26365), .B(n17590), .Z(n13424) );
  NANDN U35392 ( .A(init), .B(m[928]), .Z(n17590) );
  AND U35393 ( .A(n26366), .B(n26367), .Z(n26365) );
  NAND U35394 ( .A(o[928]), .B(n23579), .Z(n26367) );
  NANDN U35395 ( .A(n23580), .B(creg[928]), .Z(n26366) );
  NAND U35396 ( .A(n26368), .B(n17588), .Z(n13423) );
  NANDN U35397 ( .A(init), .B(m[929]), .Z(n17588) );
  AND U35398 ( .A(n26369), .B(n26370), .Z(n26368) );
  NAND U35399 ( .A(o[929]), .B(n23579), .Z(n26370) );
  NANDN U35400 ( .A(n23580), .B(creg[929]), .Z(n26369) );
  NAND U35401 ( .A(n26371), .B(n17584), .Z(n13422) );
  NANDN U35402 ( .A(init), .B(m[930]), .Z(n17584) );
  AND U35403 ( .A(n26372), .B(n26373), .Z(n26371) );
  NAND U35404 ( .A(o[930]), .B(n23579), .Z(n26373) );
  NANDN U35405 ( .A(n23580), .B(creg[930]), .Z(n26372) );
  NAND U35406 ( .A(n26374), .B(n17582), .Z(n13421) );
  NANDN U35407 ( .A(init), .B(m[931]), .Z(n17582) );
  AND U35408 ( .A(n26375), .B(n26376), .Z(n26374) );
  NAND U35409 ( .A(o[931]), .B(n23579), .Z(n26376) );
  NANDN U35410 ( .A(n23580), .B(creg[931]), .Z(n26375) );
  NAND U35411 ( .A(n26377), .B(n17580), .Z(n13420) );
  NANDN U35412 ( .A(init), .B(m[932]), .Z(n17580) );
  AND U35413 ( .A(n26378), .B(n26379), .Z(n26377) );
  NAND U35414 ( .A(o[932]), .B(n23579), .Z(n26379) );
  NANDN U35415 ( .A(n23580), .B(creg[932]), .Z(n26378) );
  NAND U35416 ( .A(n26380), .B(n17578), .Z(n13419) );
  NANDN U35417 ( .A(init), .B(m[933]), .Z(n17578) );
  AND U35418 ( .A(n26381), .B(n26382), .Z(n26380) );
  NAND U35419 ( .A(o[933]), .B(n23579), .Z(n26382) );
  NANDN U35420 ( .A(n23580), .B(creg[933]), .Z(n26381) );
  NAND U35421 ( .A(n26383), .B(n17576), .Z(n13418) );
  NANDN U35422 ( .A(init), .B(m[934]), .Z(n17576) );
  AND U35423 ( .A(n26384), .B(n26385), .Z(n26383) );
  NAND U35424 ( .A(o[934]), .B(n23579), .Z(n26385) );
  NANDN U35425 ( .A(n23580), .B(creg[934]), .Z(n26384) );
  NAND U35426 ( .A(n26386), .B(n17574), .Z(n13417) );
  NANDN U35427 ( .A(init), .B(m[935]), .Z(n17574) );
  AND U35428 ( .A(n26387), .B(n26388), .Z(n26386) );
  NAND U35429 ( .A(o[935]), .B(n23579), .Z(n26388) );
  NANDN U35430 ( .A(n23580), .B(creg[935]), .Z(n26387) );
  NAND U35431 ( .A(n26389), .B(n17572), .Z(n13416) );
  NANDN U35432 ( .A(init), .B(m[936]), .Z(n17572) );
  AND U35433 ( .A(n26390), .B(n26391), .Z(n26389) );
  NAND U35434 ( .A(o[936]), .B(n23579), .Z(n26391) );
  NANDN U35435 ( .A(n23580), .B(creg[936]), .Z(n26390) );
  NAND U35436 ( .A(n26392), .B(n17570), .Z(n13415) );
  NANDN U35437 ( .A(init), .B(m[937]), .Z(n17570) );
  AND U35438 ( .A(n26393), .B(n26394), .Z(n26392) );
  NAND U35439 ( .A(o[937]), .B(n23579), .Z(n26394) );
  NANDN U35440 ( .A(n23580), .B(creg[937]), .Z(n26393) );
  NAND U35441 ( .A(n26395), .B(n17568), .Z(n13414) );
  NANDN U35442 ( .A(init), .B(m[938]), .Z(n17568) );
  AND U35443 ( .A(n26396), .B(n26397), .Z(n26395) );
  NAND U35444 ( .A(o[938]), .B(n23579), .Z(n26397) );
  NANDN U35445 ( .A(n23580), .B(creg[938]), .Z(n26396) );
  NAND U35446 ( .A(n26398), .B(n17566), .Z(n13413) );
  NANDN U35447 ( .A(init), .B(m[939]), .Z(n17566) );
  AND U35448 ( .A(n26399), .B(n26400), .Z(n26398) );
  NAND U35449 ( .A(o[939]), .B(n23579), .Z(n26400) );
  NANDN U35450 ( .A(n23580), .B(creg[939]), .Z(n26399) );
  NAND U35451 ( .A(n26401), .B(n17562), .Z(n13412) );
  NANDN U35452 ( .A(init), .B(m[940]), .Z(n17562) );
  AND U35453 ( .A(n26402), .B(n26403), .Z(n26401) );
  NAND U35454 ( .A(o[940]), .B(n23579), .Z(n26403) );
  NANDN U35455 ( .A(n23580), .B(creg[940]), .Z(n26402) );
  NAND U35456 ( .A(n26404), .B(n17560), .Z(n13411) );
  NANDN U35457 ( .A(init), .B(m[941]), .Z(n17560) );
  AND U35458 ( .A(n26405), .B(n26406), .Z(n26404) );
  NAND U35459 ( .A(o[941]), .B(n23579), .Z(n26406) );
  NANDN U35460 ( .A(n23580), .B(creg[941]), .Z(n26405) );
  NAND U35461 ( .A(n26407), .B(n17558), .Z(n13410) );
  NANDN U35462 ( .A(init), .B(m[942]), .Z(n17558) );
  AND U35463 ( .A(n26408), .B(n26409), .Z(n26407) );
  NAND U35464 ( .A(o[942]), .B(n23579), .Z(n26409) );
  NANDN U35465 ( .A(n23580), .B(creg[942]), .Z(n26408) );
  NAND U35466 ( .A(n26410), .B(n17556), .Z(n13409) );
  NANDN U35467 ( .A(init), .B(m[943]), .Z(n17556) );
  AND U35468 ( .A(n26411), .B(n26412), .Z(n26410) );
  NAND U35469 ( .A(o[943]), .B(n23579), .Z(n26412) );
  NANDN U35470 ( .A(n23580), .B(creg[943]), .Z(n26411) );
  NAND U35471 ( .A(n26413), .B(n17554), .Z(n13408) );
  NANDN U35472 ( .A(init), .B(m[944]), .Z(n17554) );
  AND U35473 ( .A(n26414), .B(n26415), .Z(n26413) );
  NAND U35474 ( .A(o[944]), .B(n23579), .Z(n26415) );
  NANDN U35475 ( .A(n23580), .B(creg[944]), .Z(n26414) );
  NAND U35476 ( .A(n26416), .B(n17552), .Z(n13407) );
  NANDN U35477 ( .A(init), .B(m[945]), .Z(n17552) );
  AND U35478 ( .A(n26417), .B(n26418), .Z(n26416) );
  NAND U35479 ( .A(o[945]), .B(n23579), .Z(n26418) );
  NANDN U35480 ( .A(n23580), .B(creg[945]), .Z(n26417) );
  NAND U35481 ( .A(n26419), .B(n17550), .Z(n13406) );
  NANDN U35482 ( .A(init), .B(m[946]), .Z(n17550) );
  AND U35483 ( .A(n26420), .B(n26421), .Z(n26419) );
  NAND U35484 ( .A(o[946]), .B(n23579), .Z(n26421) );
  NANDN U35485 ( .A(n23580), .B(creg[946]), .Z(n26420) );
  NAND U35486 ( .A(n26422), .B(n17548), .Z(n13405) );
  NANDN U35487 ( .A(init), .B(m[947]), .Z(n17548) );
  AND U35488 ( .A(n26423), .B(n26424), .Z(n26422) );
  NAND U35489 ( .A(o[947]), .B(n23579), .Z(n26424) );
  NANDN U35490 ( .A(n23580), .B(creg[947]), .Z(n26423) );
  NAND U35491 ( .A(n26425), .B(n17546), .Z(n13404) );
  NANDN U35492 ( .A(init), .B(m[948]), .Z(n17546) );
  AND U35493 ( .A(n26426), .B(n26427), .Z(n26425) );
  NAND U35494 ( .A(o[948]), .B(n23579), .Z(n26427) );
  NANDN U35495 ( .A(n23580), .B(creg[948]), .Z(n26426) );
  NAND U35496 ( .A(n26428), .B(n17544), .Z(n13403) );
  NANDN U35497 ( .A(init), .B(m[949]), .Z(n17544) );
  AND U35498 ( .A(n26429), .B(n26430), .Z(n26428) );
  NAND U35499 ( .A(o[949]), .B(n23579), .Z(n26430) );
  NANDN U35500 ( .A(n23580), .B(creg[949]), .Z(n26429) );
  NAND U35501 ( .A(n26431), .B(n17540), .Z(n13402) );
  NANDN U35502 ( .A(init), .B(m[950]), .Z(n17540) );
  AND U35503 ( .A(n26432), .B(n26433), .Z(n26431) );
  NAND U35504 ( .A(o[950]), .B(n23579), .Z(n26433) );
  NANDN U35505 ( .A(n23580), .B(creg[950]), .Z(n26432) );
  NAND U35506 ( .A(n26434), .B(n17538), .Z(n13401) );
  NANDN U35507 ( .A(init), .B(m[951]), .Z(n17538) );
  AND U35508 ( .A(n26435), .B(n26436), .Z(n26434) );
  NAND U35509 ( .A(o[951]), .B(n23579), .Z(n26436) );
  NANDN U35510 ( .A(n23580), .B(creg[951]), .Z(n26435) );
  NAND U35511 ( .A(n26437), .B(n17536), .Z(n13400) );
  NANDN U35512 ( .A(init), .B(m[952]), .Z(n17536) );
  AND U35513 ( .A(n26438), .B(n26439), .Z(n26437) );
  NAND U35514 ( .A(o[952]), .B(n23579), .Z(n26439) );
  NANDN U35515 ( .A(n23580), .B(creg[952]), .Z(n26438) );
  NAND U35516 ( .A(n26440), .B(n17534), .Z(n13399) );
  NANDN U35517 ( .A(init), .B(m[953]), .Z(n17534) );
  AND U35518 ( .A(n26441), .B(n26442), .Z(n26440) );
  NAND U35519 ( .A(o[953]), .B(n23579), .Z(n26442) );
  NANDN U35520 ( .A(n23580), .B(creg[953]), .Z(n26441) );
  NAND U35521 ( .A(n26443), .B(n17532), .Z(n13398) );
  NANDN U35522 ( .A(init), .B(m[954]), .Z(n17532) );
  AND U35523 ( .A(n26444), .B(n26445), .Z(n26443) );
  NAND U35524 ( .A(o[954]), .B(n23579), .Z(n26445) );
  NANDN U35525 ( .A(n23580), .B(creg[954]), .Z(n26444) );
  NAND U35526 ( .A(n26446), .B(n17530), .Z(n13397) );
  NANDN U35527 ( .A(init), .B(m[955]), .Z(n17530) );
  AND U35528 ( .A(n26447), .B(n26448), .Z(n26446) );
  NAND U35529 ( .A(o[955]), .B(n23579), .Z(n26448) );
  NANDN U35530 ( .A(n23580), .B(creg[955]), .Z(n26447) );
  NAND U35531 ( .A(n26449), .B(n17528), .Z(n13396) );
  NANDN U35532 ( .A(init), .B(m[956]), .Z(n17528) );
  AND U35533 ( .A(n26450), .B(n26451), .Z(n26449) );
  NAND U35534 ( .A(o[956]), .B(n23579), .Z(n26451) );
  NANDN U35535 ( .A(n23580), .B(creg[956]), .Z(n26450) );
  NAND U35536 ( .A(n26452), .B(n17526), .Z(n13395) );
  NANDN U35537 ( .A(init), .B(m[957]), .Z(n17526) );
  AND U35538 ( .A(n26453), .B(n26454), .Z(n26452) );
  NAND U35539 ( .A(o[957]), .B(n23579), .Z(n26454) );
  NANDN U35540 ( .A(n23580), .B(creg[957]), .Z(n26453) );
  NAND U35541 ( .A(n26455), .B(n17524), .Z(n13394) );
  NANDN U35542 ( .A(init), .B(m[958]), .Z(n17524) );
  AND U35543 ( .A(n26456), .B(n26457), .Z(n26455) );
  NAND U35544 ( .A(o[958]), .B(n23579), .Z(n26457) );
  NANDN U35545 ( .A(n23580), .B(creg[958]), .Z(n26456) );
  NAND U35546 ( .A(n26458), .B(n17522), .Z(n13393) );
  NANDN U35547 ( .A(init), .B(m[959]), .Z(n17522) );
  AND U35548 ( .A(n26459), .B(n26460), .Z(n26458) );
  NAND U35549 ( .A(o[959]), .B(n23579), .Z(n26460) );
  NANDN U35550 ( .A(n23580), .B(creg[959]), .Z(n26459) );
  NAND U35551 ( .A(n26461), .B(n17518), .Z(n13392) );
  NANDN U35552 ( .A(init), .B(m[960]), .Z(n17518) );
  AND U35553 ( .A(n26462), .B(n26463), .Z(n26461) );
  NAND U35554 ( .A(o[960]), .B(n23579), .Z(n26463) );
  NANDN U35555 ( .A(n23580), .B(creg[960]), .Z(n26462) );
  NAND U35556 ( .A(n26464), .B(n17516), .Z(n13391) );
  NANDN U35557 ( .A(init), .B(m[961]), .Z(n17516) );
  AND U35558 ( .A(n26465), .B(n26466), .Z(n26464) );
  NAND U35559 ( .A(o[961]), .B(n23579), .Z(n26466) );
  NANDN U35560 ( .A(n23580), .B(creg[961]), .Z(n26465) );
  NAND U35561 ( .A(n26467), .B(n17514), .Z(n13390) );
  NANDN U35562 ( .A(init), .B(m[962]), .Z(n17514) );
  AND U35563 ( .A(n26468), .B(n26469), .Z(n26467) );
  NAND U35564 ( .A(o[962]), .B(n23579), .Z(n26469) );
  NANDN U35565 ( .A(n23580), .B(creg[962]), .Z(n26468) );
  NAND U35566 ( .A(n26470), .B(n17512), .Z(n13389) );
  NANDN U35567 ( .A(init), .B(m[963]), .Z(n17512) );
  AND U35568 ( .A(n26471), .B(n26472), .Z(n26470) );
  NAND U35569 ( .A(o[963]), .B(n23579), .Z(n26472) );
  NANDN U35570 ( .A(n23580), .B(creg[963]), .Z(n26471) );
  NAND U35571 ( .A(n26473), .B(n17510), .Z(n13388) );
  NANDN U35572 ( .A(init), .B(m[964]), .Z(n17510) );
  AND U35573 ( .A(n26474), .B(n26475), .Z(n26473) );
  NAND U35574 ( .A(o[964]), .B(n23579), .Z(n26475) );
  NANDN U35575 ( .A(n23580), .B(creg[964]), .Z(n26474) );
  NAND U35576 ( .A(n26476), .B(n17508), .Z(n13387) );
  NANDN U35577 ( .A(init), .B(m[965]), .Z(n17508) );
  AND U35578 ( .A(n26477), .B(n26478), .Z(n26476) );
  NAND U35579 ( .A(o[965]), .B(n23579), .Z(n26478) );
  NANDN U35580 ( .A(n23580), .B(creg[965]), .Z(n26477) );
  NAND U35581 ( .A(n26479), .B(n17506), .Z(n13386) );
  NANDN U35582 ( .A(init), .B(m[966]), .Z(n17506) );
  AND U35583 ( .A(n26480), .B(n26481), .Z(n26479) );
  NAND U35584 ( .A(o[966]), .B(n23579), .Z(n26481) );
  NANDN U35585 ( .A(n23580), .B(creg[966]), .Z(n26480) );
  NAND U35586 ( .A(n26482), .B(n17504), .Z(n13385) );
  NANDN U35587 ( .A(init), .B(m[967]), .Z(n17504) );
  AND U35588 ( .A(n26483), .B(n26484), .Z(n26482) );
  NAND U35589 ( .A(o[967]), .B(n23579), .Z(n26484) );
  NANDN U35590 ( .A(n23580), .B(creg[967]), .Z(n26483) );
  NAND U35591 ( .A(n26485), .B(n17502), .Z(n13384) );
  NANDN U35592 ( .A(init), .B(m[968]), .Z(n17502) );
  AND U35593 ( .A(n26486), .B(n26487), .Z(n26485) );
  NAND U35594 ( .A(o[968]), .B(n23579), .Z(n26487) );
  NANDN U35595 ( .A(n23580), .B(creg[968]), .Z(n26486) );
  NAND U35596 ( .A(n26488), .B(n17500), .Z(n13383) );
  NANDN U35597 ( .A(init), .B(m[969]), .Z(n17500) );
  AND U35598 ( .A(n26489), .B(n26490), .Z(n26488) );
  NAND U35599 ( .A(o[969]), .B(n23579), .Z(n26490) );
  NANDN U35600 ( .A(n23580), .B(creg[969]), .Z(n26489) );
  NAND U35601 ( .A(n26491), .B(n17496), .Z(n13382) );
  NANDN U35602 ( .A(init), .B(m[970]), .Z(n17496) );
  AND U35603 ( .A(n26492), .B(n26493), .Z(n26491) );
  NAND U35604 ( .A(o[970]), .B(n23579), .Z(n26493) );
  NANDN U35605 ( .A(n23580), .B(creg[970]), .Z(n26492) );
  NAND U35606 ( .A(n26494), .B(n17494), .Z(n13381) );
  NANDN U35607 ( .A(init), .B(m[971]), .Z(n17494) );
  AND U35608 ( .A(n26495), .B(n26496), .Z(n26494) );
  NAND U35609 ( .A(o[971]), .B(n23579), .Z(n26496) );
  NANDN U35610 ( .A(n23580), .B(creg[971]), .Z(n26495) );
  NAND U35611 ( .A(n26497), .B(n17492), .Z(n13380) );
  NANDN U35612 ( .A(init), .B(m[972]), .Z(n17492) );
  AND U35613 ( .A(n26498), .B(n26499), .Z(n26497) );
  NAND U35614 ( .A(o[972]), .B(n23579), .Z(n26499) );
  NANDN U35615 ( .A(n23580), .B(creg[972]), .Z(n26498) );
  NAND U35616 ( .A(n26500), .B(n17490), .Z(n13379) );
  NANDN U35617 ( .A(init), .B(m[973]), .Z(n17490) );
  AND U35618 ( .A(n26501), .B(n26502), .Z(n26500) );
  NAND U35619 ( .A(o[973]), .B(n23579), .Z(n26502) );
  NANDN U35620 ( .A(n23580), .B(creg[973]), .Z(n26501) );
  NAND U35621 ( .A(n26503), .B(n17488), .Z(n13378) );
  NANDN U35622 ( .A(init), .B(m[974]), .Z(n17488) );
  AND U35623 ( .A(n26504), .B(n26505), .Z(n26503) );
  NAND U35624 ( .A(o[974]), .B(n23579), .Z(n26505) );
  NANDN U35625 ( .A(n23580), .B(creg[974]), .Z(n26504) );
  NAND U35626 ( .A(n26506), .B(n17486), .Z(n13377) );
  NANDN U35627 ( .A(init), .B(m[975]), .Z(n17486) );
  AND U35628 ( .A(n26507), .B(n26508), .Z(n26506) );
  NAND U35629 ( .A(o[975]), .B(n23579), .Z(n26508) );
  NANDN U35630 ( .A(n23580), .B(creg[975]), .Z(n26507) );
  NAND U35631 ( .A(n26509), .B(n17484), .Z(n13376) );
  NANDN U35632 ( .A(init), .B(m[976]), .Z(n17484) );
  AND U35633 ( .A(n26510), .B(n26511), .Z(n26509) );
  NAND U35634 ( .A(o[976]), .B(n23579), .Z(n26511) );
  NANDN U35635 ( .A(n23580), .B(creg[976]), .Z(n26510) );
  NAND U35636 ( .A(n26512), .B(n17482), .Z(n13375) );
  NANDN U35637 ( .A(init), .B(m[977]), .Z(n17482) );
  AND U35638 ( .A(n26513), .B(n26514), .Z(n26512) );
  NAND U35639 ( .A(o[977]), .B(n23579), .Z(n26514) );
  NANDN U35640 ( .A(n23580), .B(creg[977]), .Z(n26513) );
  NAND U35641 ( .A(n26515), .B(n17480), .Z(n13374) );
  NANDN U35642 ( .A(init), .B(m[978]), .Z(n17480) );
  AND U35643 ( .A(n26516), .B(n26517), .Z(n26515) );
  NAND U35644 ( .A(o[978]), .B(n23579), .Z(n26517) );
  NANDN U35645 ( .A(n23580), .B(creg[978]), .Z(n26516) );
  NAND U35646 ( .A(n26518), .B(n17478), .Z(n13373) );
  NANDN U35647 ( .A(init), .B(m[979]), .Z(n17478) );
  AND U35648 ( .A(n26519), .B(n26520), .Z(n26518) );
  NAND U35649 ( .A(o[979]), .B(n23579), .Z(n26520) );
  NANDN U35650 ( .A(n23580), .B(creg[979]), .Z(n26519) );
  NAND U35651 ( .A(n26521), .B(n17474), .Z(n13372) );
  NANDN U35652 ( .A(init), .B(m[980]), .Z(n17474) );
  AND U35653 ( .A(n26522), .B(n26523), .Z(n26521) );
  NAND U35654 ( .A(o[980]), .B(n23579), .Z(n26523) );
  NANDN U35655 ( .A(n23580), .B(creg[980]), .Z(n26522) );
  NAND U35656 ( .A(n26524), .B(n17472), .Z(n13371) );
  NANDN U35657 ( .A(init), .B(m[981]), .Z(n17472) );
  AND U35658 ( .A(n26525), .B(n26526), .Z(n26524) );
  NAND U35659 ( .A(o[981]), .B(n23579), .Z(n26526) );
  NANDN U35660 ( .A(n23580), .B(creg[981]), .Z(n26525) );
  NAND U35661 ( .A(n26527), .B(n17470), .Z(n13370) );
  NANDN U35662 ( .A(init), .B(m[982]), .Z(n17470) );
  AND U35663 ( .A(n26528), .B(n26529), .Z(n26527) );
  NAND U35664 ( .A(o[982]), .B(n23579), .Z(n26529) );
  NANDN U35665 ( .A(n23580), .B(creg[982]), .Z(n26528) );
  NAND U35666 ( .A(n26530), .B(n17468), .Z(n13369) );
  NANDN U35667 ( .A(init), .B(m[983]), .Z(n17468) );
  AND U35668 ( .A(n26531), .B(n26532), .Z(n26530) );
  NAND U35669 ( .A(o[983]), .B(n23579), .Z(n26532) );
  NANDN U35670 ( .A(n23580), .B(creg[983]), .Z(n26531) );
  NAND U35671 ( .A(n26533), .B(n17466), .Z(n13368) );
  NANDN U35672 ( .A(init), .B(m[984]), .Z(n17466) );
  AND U35673 ( .A(n26534), .B(n26535), .Z(n26533) );
  NAND U35674 ( .A(o[984]), .B(n23579), .Z(n26535) );
  NANDN U35675 ( .A(n23580), .B(creg[984]), .Z(n26534) );
  NAND U35676 ( .A(n26536), .B(n17464), .Z(n13367) );
  NANDN U35677 ( .A(init), .B(m[985]), .Z(n17464) );
  AND U35678 ( .A(n26537), .B(n26538), .Z(n26536) );
  NAND U35679 ( .A(o[985]), .B(n23579), .Z(n26538) );
  NANDN U35680 ( .A(n23580), .B(creg[985]), .Z(n26537) );
  NAND U35681 ( .A(n26539), .B(n17462), .Z(n13366) );
  NANDN U35682 ( .A(init), .B(m[986]), .Z(n17462) );
  AND U35683 ( .A(n26540), .B(n26541), .Z(n26539) );
  NAND U35684 ( .A(o[986]), .B(n23579), .Z(n26541) );
  NANDN U35685 ( .A(n23580), .B(creg[986]), .Z(n26540) );
  NAND U35686 ( .A(n26542), .B(n17460), .Z(n13365) );
  NANDN U35687 ( .A(init), .B(m[987]), .Z(n17460) );
  AND U35688 ( .A(n26543), .B(n26544), .Z(n26542) );
  NAND U35689 ( .A(o[987]), .B(n23579), .Z(n26544) );
  NANDN U35690 ( .A(n23580), .B(creg[987]), .Z(n26543) );
  NAND U35691 ( .A(n26545), .B(n17458), .Z(n13364) );
  NANDN U35692 ( .A(init), .B(m[988]), .Z(n17458) );
  AND U35693 ( .A(n26546), .B(n26547), .Z(n26545) );
  NAND U35694 ( .A(o[988]), .B(n23579), .Z(n26547) );
  NANDN U35695 ( .A(n23580), .B(creg[988]), .Z(n26546) );
  NAND U35696 ( .A(n26548), .B(n17456), .Z(n13363) );
  NANDN U35697 ( .A(init), .B(m[989]), .Z(n17456) );
  AND U35698 ( .A(n26549), .B(n26550), .Z(n26548) );
  NAND U35699 ( .A(o[989]), .B(n23579), .Z(n26550) );
  NANDN U35700 ( .A(n23580), .B(creg[989]), .Z(n26549) );
  NAND U35701 ( .A(n26551), .B(n17452), .Z(n13362) );
  NANDN U35702 ( .A(init), .B(m[990]), .Z(n17452) );
  AND U35703 ( .A(n26552), .B(n26553), .Z(n26551) );
  NAND U35704 ( .A(o[990]), .B(n23579), .Z(n26553) );
  NANDN U35705 ( .A(n23580), .B(creg[990]), .Z(n26552) );
  NAND U35706 ( .A(n26554), .B(n17450), .Z(n13361) );
  NANDN U35707 ( .A(init), .B(m[991]), .Z(n17450) );
  AND U35708 ( .A(n26555), .B(n26556), .Z(n26554) );
  NAND U35709 ( .A(o[991]), .B(n23579), .Z(n26556) );
  NANDN U35710 ( .A(n23580), .B(creg[991]), .Z(n26555) );
  NAND U35711 ( .A(n26557), .B(n17448), .Z(n13360) );
  NANDN U35712 ( .A(init), .B(m[992]), .Z(n17448) );
  AND U35713 ( .A(n26558), .B(n26559), .Z(n26557) );
  NAND U35714 ( .A(o[992]), .B(n23579), .Z(n26559) );
  NANDN U35715 ( .A(n23580), .B(creg[992]), .Z(n26558) );
  NAND U35716 ( .A(n26560), .B(n17446), .Z(n13359) );
  NANDN U35717 ( .A(init), .B(m[993]), .Z(n17446) );
  AND U35718 ( .A(n26561), .B(n26562), .Z(n26560) );
  NAND U35719 ( .A(o[993]), .B(n23579), .Z(n26562) );
  NANDN U35720 ( .A(n23580), .B(creg[993]), .Z(n26561) );
  NAND U35721 ( .A(n26563), .B(n17444), .Z(n13358) );
  NANDN U35722 ( .A(init), .B(m[994]), .Z(n17444) );
  AND U35723 ( .A(n26564), .B(n26565), .Z(n26563) );
  NAND U35724 ( .A(o[994]), .B(n23579), .Z(n26565) );
  NANDN U35725 ( .A(n23580), .B(creg[994]), .Z(n26564) );
  NAND U35726 ( .A(n26566), .B(n17442), .Z(n13357) );
  NANDN U35727 ( .A(init), .B(m[995]), .Z(n17442) );
  AND U35728 ( .A(n26567), .B(n26568), .Z(n26566) );
  NAND U35729 ( .A(o[995]), .B(n23579), .Z(n26568) );
  NANDN U35730 ( .A(n23580), .B(creg[995]), .Z(n26567) );
  NAND U35731 ( .A(n26569), .B(n17440), .Z(n13356) );
  NANDN U35732 ( .A(init), .B(m[996]), .Z(n17440) );
  AND U35733 ( .A(n26570), .B(n26571), .Z(n26569) );
  NAND U35734 ( .A(o[996]), .B(n23579), .Z(n26571) );
  NANDN U35735 ( .A(n23580), .B(creg[996]), .Z(n26570) );
  NAND U35736 ( .A(n26572), .B(n17438), .Z(n13355) );
  NANDN U35737 ( .A(init), .B(m[997]), .Z(n17438) );
  AND U35738 ( .A(n26573), .B(n26574), .Z(n26572) );
  NAND U35739 ( .A(o[997]), .B(n23579), .Z(n26574) );
  NANDN U35740 ( .A(n23580), .B(creg[997]), .Z(n26573) );
  NAND U35741 ( .A(n26575), .B(n17436), .Z(n13354) );
  NANDN U35742 ( .A(init), .B(m[998]), .Z(n17436) );
  AND U35743 ( .A(n26576), .B(n26577), .Z(n26575) );
  NAND U35744 ( .A(o[998]), .B(n23579), .Z(n26577) );
  NANDN U35745 ( .A(n23580), .B(creg[998]), .Z(n26576) );
  NAND U35746 ( .A(n26578), .B(n17434), .Z(n13353) );
  NANDN U35747 ( .A(init), .B(m[999]), .Z(n17434) );
  AND U35748 ( .A(n26579), .B(n26580), .Z(n26578) );
  NAND U35749 ( .A(o[999]), .B(n23579), .Z(n26580) );
  NANDN U35750 ( .A(n23580), .B(creg[999]), .Z(n26579) );
  NAND U35751 ( .A(n26581), .B(n19474), .Z(n13352) );
  NANDN U35752 ( .A(init), .B(m[1000]), .Z(n19474) );
  AND U35753 ( .A(n26582), .B(n26583), .Z(n26581) );
  NAND U35754 ( .A(o[1000]), .B(n23579), .Z(n26583) );
  NANDN U35755 ( .A(n23580), .B(creg[1000]), .Z(n26582) );
  NAND U35756 ( .A(n26584), .B(n19472), .Z(n13351) );
  NANDN U35757 ( .A(init), .B(m[1001]), .Z(n19472) );
  AND U35758 ( .A(n26585), .B(n26586), .Z(n26584) );
  NAND U35759 ( .A(o[1001]), .B(n23579), .Z(n26586) );
  NANDN U35760 ( .A(n23580), .B(creg[1001]), .Z(n26585) );
  NAND U35761 ( .A(n26587), .B(n19470), .Z(n13350) );
  NANDN U35762 ( .A(init), .B(m[1002]), .Z(n19470) );
  AND U35763 ( .A(n26588), .B(n26589), .Z(n26587) );
  NAND U35764 ( .A(o[1002]), .B(n23579), .Z(n26589) );
  NANDN U35765 ( .A(n23580), .B(creg[1002]), .Z(n26588) );
  NAND U35766 ( .A(n26590), .B(n19468), .Z(n13349) );
  NANDN U35767 ( .A(init), .B(m[1003]), .Z(n19468) );
  AND U35768 ( .A(n26591), .B(n26592), .Z(n26590) );
  NAND U35769 ( .A(o[1003]), .B(n23579), .Z(n26592) );
  NANDN U35770 ( .A(n23580), .B(creg[1003]), .Z(n26591) );
  NAND U35771 ( .A(n26593), .B(n19466), .Z(n13348) );
  NANDN U35772 ( .A(init), .B(m[1004]), .Z(n19466) );
  AND U35773 ( .A(n26594), .B(n26595), .Z(n26593) );
  NAND U35774 ( .A(o[1004]), .B(n23579), .Z(n26595) );
  NANDN U35775 ( .A(n23580), .B(creg[1004]), .Z(n26594) );
  NAND U35776 ( .A(n26596), .B(n19464), .Z(n13347) );
  NANDN U35777 ( .A(init), .B(m[1005]), .Z(n19464) );
  AND U35778 ( .A(n26597), .B(n26598), .Z(n26596) );
  NAND U35779 ( .A(o[1005]), .B(n23579), .Z(n26598) );
  NANDN U35780 ( .A(n23580), .B(creg[1005]), .Z(n26597) );
  NAND U35781 ( .A(n26599), .B(n19462), .Z(n13346) );
  NANDN U35782 ( .A(init), .B(m[1006]), .Z(n19462) );
  AND U35783 ( .A(n26600), .B(n26601), .Z(n26599) );
  NAND U35784 ( .A(o[1006]), .B(n23579), .Z(n26601) );
  NANDN U35785 ( .A(n23580), .B(creg[1006]), .Z(n26600) );
  NAND U35786 ( .A(n26602), .B(n19460), .Z(n13345) );
  NANDN U35787 ( .A(init), .B(m[1007]), .Z(n19460) );
  AND U35788 ( .A(n26603), .B(n26604), .Z(n26602) );
  NAND U35789 ( .A(o[1007]), .B(n23579), .Z(n26604) );
  NANDN U35790 ( .A(n23580), .B(creg[1007]), .Z(n26603) );
  NAND U35791 ( .A(n26605), .B(n19458), .Z(n13344) );
  NANDN U35792 ( .A(init), .B(m[1008]), .Z(n19458) );
  AND U35793 ( .A(n26606), .B(n26607), .Z(n26605) );
  NAND U35794 ( .A(o[1008]), .B(n23579), .Z(n26607) );
  NANDN U35795 ( .A(n23580), .B(creg[1008]), .Z(n26606) );
  NAND U35796 ( .A(n26608), .B(n19456), .Z(n13343) );
  NANDN U35797 ( .A(init), .B(m[1009]), .Z(n19456) );
  AND U35798 ( .A(n26609), .B(n26610), .Z(n26608) );
  NAND U35799 ( .A(o[1009]), .B(n23579), .Z(n26610) );
  NANDN U35800 ( .A(n23580), .B(creg[1009]), .Z(n26609) );
  NAND U35801 ( .A(n26611), .B(n19452), .Z(n13342) );
  NANDN U35802 ( .A(init), .B(m[1010]), .Z(n19452) );
  AND U35803 ( .A(n26612), .B(n26613), .Z(n26611) );
  NAND U35804 ( .A(o[1010]), .B(n23579), .Z(n26613) );
  NANDN U35805 ( .A(n23580), .B(creg[1010]), .Z(n26612) );
  NAND U35806 ( .A(n26614), .B(n19450), .Z(n13341) );
  NANDN U35807 ( .A(init), .B(m[1011]), .Z(n19450) );
  AND U35808 ( .A(n26615), .B(n26616), .Z(n26614) );
  NAND U35809 ( .A(o[1011]), .B(n23579), .Z(n26616) );
  NANDN U35810 ( .A(n23580), .B(creg[1011]), .Z(n26615) );
  NAND U35811 ( .A(n26617), .B(n19448), .Z(n13340) );
  NANDN U35812 ( .A(init), .B(m[1012]), .Z(n19448) );
  AND U35813 ( .A(n26618), .B(n26619), .Z(n26617) );
  NAND U35814 ( .A(o[1012]), .B(n23579), .Z(n26619) );
  NANDN U35815 ( .A(n23580), .B(creg[1012]), .Z(n26618) );
  NAND U35816 ( .A(n26620), .B(n19446), .Z(n13339) );
  NANDN U35817 ( .A(init), .B(m[1013]), .Z(n19446) );
  AND U35818 ( .A(n26621), .B(n26622), .Z(n26620) );
  NAND U35819 ( .A(o[1013]), .B(n23579), .Z(n26622) );
  NANDN U35820 ( .A(n23580), .B(creg[1013]), .Z(n26621) );
  NAND U35821 ( .A(n26623), .B(n19444), .Z(n13338) );
  NANDN U35822 ( .A(init), .B(m[1014]), .Z(n19444) );
  AND U35823 ( .A(n26624), .B(n26625), .Z(n26623) );
  NAND U35824 ( .A(o[1014]), .B(n23579), .Z(n26625) );
  NANDN U35825 ( .A(n23580), .B(creg[1014]), .Z(n26624) );
  NAND U35826 ( .A(n26626), .B(n19442), .Z(n13337) );
  NANDN U35827 ( .A(init), .B(m[1015]), .Z(n19442) );
  AND U35828 ( .A(n26627), .B(n26628), .Z(n26626) );
  NAND U35829 ( .A(o[1015]), .B(n23579), .Z(n26628) );
  NANDN U35830 ( .A(n23580), .B(creg[1015]), .Z(n26627) );
  NAND U35831 ( .A(n26629), .B(n19440), .Z(n13336) );
  NANDN U35832 ( .A(init), .B(m[1016]), .Z(n19440) );
  AND U35833 ( .A(n26630), .B(n26631), .Z(n26629) );
  NAND U35834 ( .A(o[1016]), .B(n23579), .Z(n26631) );
  NANDN U35835 ( .A(n23580), .B(creg[1016]), .Z(n26630) );
  NAND U35836 ( .A(n26632), .B(n19438), .Z(n13335) );
  NANDN U35837 ( .A(init), .B(m[1017]), .Z(n19438) );
  AND U35838 ( .A(n26633), .B(n26634), .Z(n26632) );
  NAND U35839 ( .A(o[1017]), .B(n23579), .Z(n26634) );
  NANDN U35840 ( .A(n23580), .B(creg[1017]), .Z(n26633) );
  NAND U35841 ( .A(n26635), .B(n19436), .Z(n13334) );
  NANDN U35842 ( .A(init), .B(m[1018]), .Z(n19436) );
  AND U35843 ( .A(n26636), .B(n26637), .Z(n26635) );
  NAND U35844 ( .A(o[1018]), .B(n23579), .Z(n26637) );
  NANDN U35845 ( .A(n23580), .B(creg[1018]), .Z(n26636) );
  NAND U35846 ( .A(n26638), .B(n19434), .Z(n13333) );
  NANDN U35847 ( .A(init), .B(m[1019]), .Z(n19434) );
  AND U35848 ( .A(n26639), .B(n26640), .Z(n26638) );
  NAND U35849 ( .A(o[1019]), .B(n23579), .Z(n26640) );
  NANDN U35850 ( .A(n23580), .B(creg[1019]), .Z(n26639) );
  NAND U35851 ( .A(n26641), .B(n19430), .Z(n13332) );
  NANDN U35852 ( .A(init), .B(m[1020]), .Z(n19430) );
  AND U35853 ( .A(n26642), .B(n26643), .Z(n26641) );
  NAND U35854 ( .A(o[1020]), .B(n23579), .Z(n26643) );
  NANDN U35855 ( .A(n23580), .B(creg[1020]), .Z(n26642) );
  NAND U35856 ( .A(n26644), .B(n19428), .Z(n13331) );
  NANDN U35857 ( .A(init), .B(m[1021]), .Z(n19428) );
  AND U35858 ( .A(n26645), .B(n26646), .Z(n26644) );
  NAND U35859 ( .A(o[1021]), .B(n23579), .Z(n26646) );
  NANDN U35860 ( .A(n23580), .B(creg[1021]), .Z(n26645) );
  NAND U35861 ( .A(n26647), .B(n19426), .Z(n13330) );
  NANDN U35862 ( .A(init), .B(m[1022]), .Z(n19426) );
  AND U35863 ( .A(n26648), .B(n26649), .Z(n26647) );
  NAND U35864 ( .A(o[1022]), .B(n23579), .Z(n26649) );
  AND U35865 ( .A(start_in[1023]), .B(n23580), .Z(n23579) );
  NANDN U35866 ( .A(n23580), .B(creg[1022]), .Z(n26648) );
  NAND U35867 ( .A(init), .B(n26650), .Z(n23580) );
  NAND U35868 ( .A(first_one), .B(n26651), .Z(n26650) );
  AND U35869 ( .A(start_in[1023]), .B(n26652), .Z(n26651) );
  NAND U35870 ( .A(n26653), .B(mul_pow), .Z(n26652) );
  NANDN U35871 ( .A(first_one), .B(n26654), .Z(n13329) );
  NAND U35872 ( .A(n26655), .B(ereg[1023]), .Z(n26654) );
  AND U35873 ( .A(start_in[1023]), .B(mul_pow), .Z(n26655) );
  AND U35874 ( .A(start_reg[1023]), .B(init), .Z(start_in[1023]) );
  NAND U35875 ( .A(n26656), .B(n26657), .Z(c[9]) );
  NAND U35876 ( .A(n26658), .B(o[9]), .Z(n26657) );
  NAND U35877 ( .A(n26653), .B(creg[9]), .Z(n26656) );
  NAND U35878 ( .A(n26659), .B(n26660), .Z(c[99]) );
  NAND U35879 ( .A(n26658), .B(o[99]), .Z(n26660) );
  NAND U35880 ( .A(n26653), .B(creg[99]), .Z(n26659) );
  NAND U35881 ( .A(n26661), .B(n26662), .Z(c[999]) );
  NAND U35882 ( .A(n26658), .B(o[999]), .Z(n26662) );
  NAND U35883 ( .A(n26653), .B(creg[999]), .Z(n26661) );
  NAND U35884 ( .A(n26663), .B(n26664), .Z(c[998]) );
  NAND U35885 ( .A(n26658), .B(o[998]), .Z(n26664) );
  NAND U35886 ( .A(n26653), .B(creg[998]), .Z(n26663) );
  NAND U35887 ( .A(n26665), .B(n26666), .Z(c[997]) );
  NAND U35888 ( .A(n26658), .B(o[997]), .Z(n26666) );
  NAND U35889 ( .A(n26653), .B(creg[997]), .Z(n26665) );
  NAND U35890 ( .A(n26667), .B(n26668), .Z(c[996]) );
  NAND U35891 ( .A(n26658), .B(o[996]), .Z(n26668) );
  NAND U35892 ( .A(n26653), .B(creg[996]), .Z(n26667) );
  NAND U35893 ( .A(n26669), .B(n26670), .Z(c[995]) );
  NAND U35894 ( .A(n26658), .B(o[995]), .Z(n26670) );
  NAND U35895 ( .A(n26653), .B(creg[995]), .Z(n26669) );
  NAND U35896 ( .A(n26671), .B(n26672), .Z(c[994]) );
  NAND U35897 ( .A(n26658), .B(o[994]), .Z(n26672) );
  NAND U35898 ( .A(n26653), .B(creg[994]), .Z(n26671) );
  NAND U35899 ( .A(n26673), .B(n26674), .Z(c[993]) );
  NAND U35900 ( .A(n26658), .B(o[993]), .Z(n26674) );
  NAND U35901 ( .A(n26653), .B(creg[993]), .Z(n26673) );
  NAND U35902 ( .A(n26675), .B(n26676), .Z(c[992]) );
  NAND U35903 ( .A(n26658), .B(o[992]), .Z(n26676) );
  NAND U35904 ( .A(n26653), .B(creg[992]), .Z(n26675) );
  NAND U35905 ( .A(n26677), .B(n26678), .Z(c[991]) );
  NAND U35906 ( .A(n26658), .B(o[991]), .Z(n26678) );
  NAND U35907 ( .A(n26653), .B(creg[991]), .Z(n26677) );
  NAND U35908 ( .A(n26679), .B(n26680), .Z(c[990]) );
  NAND U35909 ( .A(n26658), .B(o[990]), .Z(n26680) );
  NAND U35910 ( .A(n26653), .B(creg[990]), .Z(n26679) );
  NAND U35911 ( .A(n26681), .B(n26682), .Z(c[98]) );
  NAND U35912 ( .A(n26658), .B(o[98]), .Z(n26682) );
  NAND U35913 ( .A(n26653), .B(creg[98]), .Z(n26681) );
  NAND U35914 ( .A(n26683), .B(n26684), .Z(c[989]) );
  NAND U35915 ( .A(n26658), .B(o[989]), .Z(n26684) );
  NAND U35916 ( .A(n26653), .B(creg[989]), .Z(n26683) );
  NAND U35917 ( .A(n26685), .B(n26686), .Z(c[988]) );
  NAND U35918 ( .A(n26658), .B(o[988]), .Z(n26686) );
  NAND U35919 ( .A(n26653), .B(creg[988]), .Z(n26685) );
  NAND U35920 ( .A(n26687), .B(n26688), .Z(c[987]) );
  NAND U35921 ( .A(n26658), .B(o[987]), .Z(n26688) );
  NAND U35922 ( .A(n26653), .B(creg[987]), .Z(n26687) );
  NAND U35923 ( .A(n26689), .B(n26690), .Z(c[986]) );
  NAND U35924 ( .A(n26658), .B(o[986]), .Z(n26690) );
  NAND U35925 ( .A(n26653), .B(creg[986]), .Z(n26689) );
  NAND U35926 ( .A(n26691), .B(n26692), .Z(c[985]) );
  NAND U35927 ( .A(n26658), .B(o[985]), .Z(n26692) );
  NAND U35928 ( .A(n26653), .B(creg[985]), .Z(n26691) );
  NAND U35929 ( .A(n26693), .B(n26694), .Z(c[984]) );
  NAND U35930 ( .A(n26658), .B(o[984]), .Z(n26694) );
  NAND U35931 ( .A(n26653), .B(creg[984]), .Z(n26693) );
  NAND U35932 ( .A(n26695), .B(n26696), .Z(c[983]) );
  NAND U35933 ( .A(n26658), .B(o[983]), .Z(n26696) );
  NAND U35934 ( .A(n26653), .B(creg[983]), .Z(n26695) );
  NAND U35935 ( .A(n26697), .B(n26698), .Z(c[982]) );
  NAND U35936 ( .A(n26658), .B(o[982]), .Z(n26698) );
  NAND U35937 ( .A(n26653), .B(creg[982]), .Z(n26697) );
  NAND U35938 ( .A(n26699), .B(n26700), .Z(c[981]) );
  NAND U35939 ( .A(n26658), .B(o[981]), .Z(n26700) );
  NAND U35940 ( .A(n26653), .B(creg[981]), .Z(n26699) );
  NAND U35941 ( .A(n26701), .B(n26702), .Z(c[980]) );
  NAND U35942 ( .A(n26658), .B(o[980]), .Z(n26702) );
  NAND U35943 ( .A(n26653), .B(creg[980]), .Z(n26701) );
  NAND U35944 ( .A(n26703), .B(n26704), .Z(c[97]) );
  NAND U35945 ( .A(n26658), .B(o[97]), .Z(n26704) );
  NAND U35946 ( .A(n26653), .B(creg[97]), .Z(n26703) );
  NAND U35947 ( .A(n26705), .B(n26706), .Z(c[979]) );
  NAND U35948 ( .A(n26658), .B(o[979]), .Z(n26706) );
  NAND U35949 ( .A(n26653), .B(creg[979]), .Z(n26705) );
  NAND U35950 ( .A(n26707), .B(n26708), .Z(c[978]) );
  NAND U35951 ( .A(n26658), .B(o[978]), .Z(n26708) );
  NAND U35952 ( .A(n26653), .B(creg[978]), .Z(n26707) );
  NAND U35953 ( .A(n26709), .B(n26710), .Z(c[977]) );
  NAND U35954 ( .A(n26658), .B(o[977]), .Z(n26710) );
  NAND U35955 ( .A(n26653), .B(creg[977]), .Z(n26709) );
  NAND U35956 ( .A(n26711), .B(n26712), .Z(c[976]) );
  NAND U35957 ( .A(n26658), .B(o[976]), .Z(n26712) );
  NAND U35958 ( .A(n26653), .B(creg[976]), .Z(n26711) );
  NAND U35959 ( .A(n26713), .B(n26714), .Z(c[975]) );
  NAND U35960 ( .A(n26658), .B(o[975]), .Z(n26714) );
  NAND U35961 ( .A(n26653), .B(creg[975]), .Z(n26713) );
  NAND U35962 ( .A(n26715), .B(n26716), .Z(c[974]) );
  NAND U35963 ( .A(n26658), .B(o[974]), .Z(n26716) );
  NAND U35964 ( .A(n26653), .B(creg[974]), .Z(n26715) );
  NAND U35965 ( .A(n26717), .B(n26718), .Z(c[973]) );
  NAND U35966 ( .A(n26658), .B(o[973]), .Z(n26718) );
  NAND U35967 ( .A(n26653), .B(creg[973]), .Z(n26717) );
  NAND U35968 ( .A(n26719), .B(n26720), .Z(c[972]) );
  NAND U35969 ( .A(n26658), .B(o[972]), .Z(n26720) );
  NAND U35970 ( .A(n26653), .B(creg[972]), .Z(n26719) );
  NAND U35971 ( .A(n26721), .B(n26722), .Z(c[971]) );
  NAND U35972 ( .A(n26658), .B(o[971]), .Z(n26722) );
  NAND U35973 ( .A(n26653), .B(creg[971]), .Z(n26721) );
  NAND U35974 ( .A(n26723), .B(n26724), .Z(c[970]) );
  NAND U35975 ( .A(n26658), .B(o[970]), .Z(n26724) );
  NAND U35976 ( .A(n26653), .B(creg[970]), .Z(n26723) );
  NAND U35977 ( .A(n26725), .B(n26726), .Z(c[96]) );
  NAND U35978 ( .A(n26658), .B(o[96]), .Z(n26726) );
  NAND U35979 ( .A(n26653), .B(creg[96]), .Z(n26725) );
  NAND U35980 ( .A(n26727), .B(n26728), .Z(c[969]) );
  NAND U35981 ( .A(n26658), .B(o[969]), .Z(n26728) );
  NAND U35982 ( .A(n26653), .B(creg[969]), .Z(n26727) );
  NAND U35983 ( .A(n26729), .B(n26730), .Z(c[968]) );
  NAND U35984 ( .A(n26658), .B(o[968]), .Z(n26730) );
  NAND U35985 ( .A(n26653), .B(creg[968]), .Z(n26729) );
  NAND U35986 ( .A(n26731), .B(n26732), .Z(c[967]) );
  NAND U35987 ( .A(n26658), .B(o[967]), .Z(n26732) );
  NAND U35988 ( .A(n26653), .B(creg[967]), .Z(n26731) );
  NAND U35989 ( .A(n26733), .B(n26734), .Z(c[966]) );
  NAND U35990 ( .A(n26658), .B(o[966]), .Z(n26734) );
  NAND U35991 ( .A(n26653), .B(creg[966]), .Z(n26733) );
  NAND U35992 ( .A(n26735), .B(n26736), .Z(c[965]) );
  NAND U35993 ( .A(n26658), .B(o[965]), .Z(n26736) );
  NAND U35994 ( .A(n26653), .B(creg[965]), .Z(n26735) );
  NAND U35995 ( .A(n26737), .B(n26738), .Z(c[964]) );
  NAND U35996 ( .A(n26658), .B(o[964]), .Z(n26738) );
  NAND U35997 ( .A(n26653), .B(creg[964]), .Z(n26737) );
  NAND U35998 ( .A(n26739), .B(n26740), .Z(c[963]) );
  NAND U35999 ( .A(n26658), .B(o[963]), .Z(n26740) );
  NAND U36000 ( .A(n26653), .B(creg[963]), .Z(n26739) );
  NAND U36001 ( .A(n26741), .B(n26742), .Z(c[962]) );
  NAND U36002 ( .A(n26658), .B(o[962]), .Z(n26742) );
  NAND U36003 ( .A(n26653), .B(creg[962]), .Z(n26741) );
  NAND U36004 ( .A(n26743), .B(n26744), .Z(c[961]) );
  NAND U36005 ( .A(n26658), .B(o[961]), .Z(n26744) );
  NAND U36006 ( .A(n26653), .B(creg[961]), .Z(n26743) );
  NAND U36007 ( .A(n26745), .B(n26746), .Z(c[960]) );
  NAND U36008 ( .A(n26658), .B(o[960]), .Z(n26746) );
  NAND U36009 ( .A(n26653), .B(creg[960]), .Z(n26745) );
  NAND U36010 ( .A(n26747), .B(n26748), .Z(c[95]) );
  NAND U36011 ( .A(n26658), .B(o[95]), .Z(n26748) );
  NAND U36012 ( .A(n26653), .B(creg[95]), .Z(n26747) );
  NAND U36013 ( .A(n26749), .B(n26750), .Z(c[959]) );
  NAND U36014 ( .A(n26658), .B(o[959]), .Z(n26750) );
  NAND U36015 ( .A(n26653), .B(creg[959]), .Z(n26749) );
  NAND U36016 ( .A(n26751), .B(n26752), .Z(c[958]) );
  NAND U36017 ( .A(n26658), .B(o[958]), .Z(n26752) );
  NAND U36018 ( .A(n26653), .B(creg[958]), .Z(n26751) );
  NAND U36019 ( .A(n26753), .B(n26754), .Z(c[957]) );
  NAND U36020 ( .A(n26658), .B(o[957]), .Z(n26754) );
  NAND U36021 ( .A(n26653), .B(creg[957]), .Z(n26753) );
  NAND U36022 ( .A(n26755), .B(n26756), .Z(c[956]) );
  NAND U36023 ( .A(n26658), .B(o[956]), .Z(n26756) );
  NAND U36024 ( .A(n26653), .B(creg[956]), .Z(n26755) );
  NAND U36025 ( .A(n26757), .B(n26758), .Z(c[955]) );
  NAND U36026 ( .A(n26658), .B(o[955]), .Z(n26758) );
  NAND U36027 ( .A(n26653), .B(creg[955]), .Z(n26757) );
  NAND U36028 ( .A(n26759), .B(n26760), .Z(c[954]) );
  NAND U36029 ( .A(n26658), .B(o[954]), .Z(n26760) );
  NAND U36030 ( .A(n26653), .B(creg[954]), .Z(n26759) );
  NAND U36031 ( .A(n26761), .B(n26762), .Z(c[953]) );
  NAND U36032 ( .A(n26658), .B(o[953]), .Z(n26762) );
  NAND U36033 ( .A(n26653), .B(creg[953]), .Z(n26761) );
  NAND U36034 ( .A(n26763), .B(n26764), .Z(c[952]) );
  NAND U36035 ( .A(n26658), .B(o[952]), .Z(n26764) );
  NAND U36036 ( .A(n26653), .B(creg[952]), .Z(n26763) );
  NAND U36037 ( .A(n26765), .B(n26766), .Z(c[951]) );
  NAND U36038 ( .A(n26658), .B(o[951]), .Z(n26766) );
  NAND U36039 ( .A(n26653), .B(creg[951]), .Z(n26765) );
  NAND U36040 ( .A(n26767), .B(n26768), .Z(c[950]) );
  NAND U36041 ( .A(n26658), .B(o[950]), .Z(n26768) );
  NAND U36042 ( .A(n26653), .B(creg[950]), .Z(n26767) );
  NAND U36043 ( .A(n26769), .B(n26770), .Z(c[94]) );
  NAND U36044 ( .A(n26658), .B(o[94]), .Z(n26770) );
  NAND U36045 ( .A(n26653), .B(creg[94]), .Z(n26769) );
  NAND U36046 ( .A(n26771), .B(n26772), .Z(c[949]) );
  NAND U36047 ( .A(n26658), .B(o[949]), .Z(n26772) );
  NAND U36048 ( .A(n26653), .B(creg[949]), .Z(n26771) );
  NAND U36049 ( .A(n26773), .B(n26774), .Z(c[948]) );
  NAND U36050 ( .A(n26658), .B(o[948]), .Z(n26774) );
  NAND U36051 ( .A(n26653), .B(creg[948]), .Z(n26773) );
  NAND U36052 ( .A(n26775), .B(n26776), .Z(c[947]) );
  NAND U36053 ( .A(n26658), .B(o[947]), .Z(n26776) );
  NAND U36054 ( .A(n26653), .B(creg[947]), .Z(n26775) );
  NAND U36055 ( .A(n26777), .B(n26778), .Z(c[946]) );
  NAND U36056 ( .A(n26658), .B(o[946]), .Z(n26778) );
  NAND U36057 ( .A(n26653), .B(creg[946]), .Z(n26777) );
  NAND U36058 ( .A(n26779), .B(n26780), .Z(c[945]) );
  NAND U36059 ( .A(n26658), .B(o[945]), .Z(n26780) );
  NAND U36060 ( .A(n26653), .B(creg[945]), .Z(n26779) );
  NAND U36061 ( .A(n26781), .B(n26782), .Z(c[944]) );
  NAND U36062 ( .A(n26658), .B(o[944]), .Z(n26782) );
  NAND U36063 ( .A(n26653), .B(creg[944]), .Z(n26781) );
  NAND U36064 ( .A(n26783), .B(n26784), .Z(c[943]) );
  NAND U36065 ( .A(n26658), .B(o[943]), .Z(n26784) );
  NAND U36066 ( .A(n26653), .B(creg[943]), .Z(n26783) );
  NAND U36067 ( .A(n26785), .B(n26786), .Z(c[942]) );
  NAND U36068 ( .A(n26658), .B(o[942]), .Z(n26786) );
  NAND U36069 ( .A(n26653), .B(creg[942]), .Z(n26785) );
  NAND U36070 ( .A(n26787), .B(n26788), .Z(c[941]) );
  NAND U36071 ( .A(n26658), .B(o[941]), .Z(n26788) );
  NAND U36072 ( .A(n26653), .B(creg[941]), .Z(n26787) );
  NAND U36073 ( .A(n26789), .B(n26790), .Z(c[940]) );
  NAND U36074 ( .A(n26658), .B(o[940]), .Z(n26790) );
  NAND U36075 ( .A(n26653), .B(creg[940]), .Z(n26789) );
  NAND U36076 ( .A(n26791), .B(n26792), .Z(c[93]) );
  NAND U36077 ( .A(n26658), .B(o[93]), .Z(n26792) );
  NAND U36078 ( .A(n26653), .B(creg[93]), .Z(n26791) );
  NAND U36079 ( .A(n26793), .B(n26794), .Z(c[939]) );
  NAND U36080 ( .A(n26658), .B(o[939]), .Z(n26794) );
  NAND U36081 ( .A(n26653), .B(creg[939]), .Z(n26793) );
  NAND U36082 ( .A(n26795), .B(n26796), .Z(c[938]) );
  NAND U36083 ( .A(n26658), .B(o[938]), .Z(n26796) );
  NAND U36084 ( .A(n26653), .B(creg[938]), .Z(n26795) );
  NAND U36085 ( .A(n26797), .B(n26798), .Z(c[937]) );
  NAND U36086 ( .A(n26658), .B(o[937]), .Z(n26798) );
  NAND U36087 ( .A(n26653), .B(creg[937]), .Z(n26797) );
  NAND U36088 ( .A(n26799), .B(n26800), .Z(c[936]) );
  NAND U36089 ( .A(n26658), .B(o[936]), .Z(n26800) );
  NAND U36090 ( .A(n26653), .B(creg[936]), .Z(n26799) );
  NAND U36091 ( .A(n26801), .B(n26802), .Z(c[935]) );
  NAND U36092 ( .A(n26658), .B(o[935]), .Z(n26802) );
  NAND U36093 ( .A(n26653), .B(creg[935]), .Z(n26801) );
  NAND U36094 ( .A(n26803), .B(n26804), .Z(c[934]) );
  NAND U36095 ( .A(n26658), .B(o[934]), .Z(n26804) );
  NAND U36096 ( .A(n26653), .B(creg[934]), .Z(n26803) );
  NAND U36097 ( .A(n26805), .B(n26806), .Z(c[933]) );
  NAND U36098 ( .A(n26658), .B(o[933]), .Z(n26806) );
  NAND U36099 ( .A(n26653), .B(creg[933]), .Z(n26805) );
  NAND U36100 ( .A(n26807), .B(n26808), .Z(c[932]) );
  NAND U36101 ( .A(n26658), .B(o[932]), .Z(n26808) );
  NAND U36102 ( .A(n26653), .B(creg[932]), .Z(n26807) );
  NAND U36103 ( .A(n26809), .B(n26810), .Z(c[931]) );
  NAND U36104 ( .A(n26658), .B(o[931]), .Z(n26810) );
  NAND U36105 ( .A(n26653), .B(creg[931]), .Z(n26809) );
  NAND U36106 ( .A(n26811), .B(n26812), .Z(c[930]) );
  NAND U36107 ( .A(n26658), .B(o[930]), .Z(n26812) );
  NAND U36108 ( .A(n26653), .B(creg[930]), .Z(n26811) );
  NAND U36109 ( .A(n26813), .B(n26814), .Z(c[92]) );
  NAND U36110 ( .A(n26658), .B(o[92]), .Z(n26814) );
  NAND U36111 ( .A(n26653), .B(creg[92]), .Z(n26813) );
  NAND U36112 ( .A(n26815), .B(n26816), .Z(c[929]) );
  NAND U36113 ( .A(n26658), .B(o[929]), .Z(n26816) );
  NAND U36114 ( .A(n26653), .B(creg[929]), .Z(n26815) );
  NAND U36115 ( .A(n26817), .B(n26818), .Z(c[928]) );
  NAND U36116 ( .A(n26658), .B(o[928]), .Z(n26818) );
  NAND U36117 ( .A(n26653), .B(creg[928]), .Z(n26817) );
  NAND U36118 ( .A(n26819), .B(n26820), .Z(c[927]) );
  NAND U36119 ( .A(n26658), .B(o[927]), .Z(n26820) );
  NAND U36120 ( .A(n26653), .B(creg[927]), .Z(n26819) );
  NAND U36121 ( .A(n26821), .B(n26822), .Z(c[926]) );
  NAND U36122 ( .A(n26658), .B(o[926]), .Z(n26822) );
  NAND U36123 ( .A(n26653), .B(creg[926]), .Z(n26821) );
  NAND U36124 ( .A(n26823), .B(n26824), .Z(c[925]) );
  NAND U36125 ( .A(n26658), .B(o[925]), .Z(n26824) );
  NAND U36126 ( .A(n26653), .B(creg[925]), .Z(n26823) );
  NAND U36127 ( .A(n26825), .B(n26826), .Z(c[924]) );
  NAND U36128 ( .A(n26658), .B(o[924]), .Z(n26826) );
  NAND U36129 ( .A(n26653), .B(creg[924]), .Z(n26825) );
  NAND U36130 ( .A(n26827), .B(n26828), .Z(c[923]) );
  NAND U36131 ( .A(n26658), .B(o[923]), .Z(n26828) );
  NAND U36132 ( .A(n26653), .B(creg[923]), .Z(n26827) );
  NAND U36133 ( .A(n26829), .B(n26830), .Z(c[922]) );
  NAND U36134 ( .A(n26658), .B(o[922]), .Z(n26830) );
  NAND U36135 ( .A(n26653), .B(creg[922]), .Z(n26829) );
  NAND U36136 ( .A(n26831), .B(n26832), .Z(c[921]) );
  NAND U36137 ( .A(n26658), .B(o[921]), .Z(n26832) );
  NAND U36138 ( .A(n26653), .B(creg[921]), .Z(n26831) );
  NAND U36139 ( .A(n26833), .B(n26834), .Z(c[920]) );
  NAND U36140 ( .A(n26658), .B(o[920]), .Z(n26834) );
  NAND U36141 ( .A(n26653), .B(creg[920]), .Z(n26833) );
  NAND U36142 ( .A(n26835), .B(n26836), .Z(c[91]) );
  NAND U36143 ( .A(n26658), .B(o[91]), .Z(n26836) );
  NAND U36144 ( .A(n26653), .B(creg[91]), .Z(n26835) );
  NAND U36145 ( .A(n26837), .B(n26838), .Z(c[919]) );
  NAND U36146 ( .A(n26658), .B(o[919]), .Z(n26838) );
  NAND U36147 ( .A(n26653), .B(creg[919]), .Z(n26837) );
  NAND U36148 ( .A(n26839), .B(n26840), .Z(c[918]) );
  NAND U36149 ( .A(n26658), .B(o[918]), .Z(n26840) );
  NAND U36150 ( .A(n26653), .B(creg[918]), .Z(n26839) );
  NAND U36151 ( .A(n26841), .B(n26842), .Z(c[917]) );
  NAND U36152 ( .A(n26658), .B(o[917]), .Z(n26842) );
  NAND U36153 ( .A(n26653), .B(creg[917]), .Z(n26841) );
  NAND U36154 ( .A(n26843), .B(n26844), .Z(c[916]) );
  NAND U36155 ( .A(n26658), .B(o[916]), .Z(n26844) );
  NAND U36156 ( .A(n26653), .B(creg[916]), .Z(n26843) );
  NAND U36157 ( .A(n26845), .B(n26846), .Z(c[915]) );
  NAND U36158 ( .A(n26658), .B(o[915]), .Z(n26846) );
  NAND U36159 ( .A(n26653), .B(creg[915]), .Z(n26845) );
  NAND U36160 ( .A(n26847), .B(n26848), .Z(c[914]) );
  NAND U36161 ( .A(n26658), .B(o[914]), .Z(n26848) );
  NAND U36162 ( .A(n26653), .B(creg[914]), .Z(n26847) );
  NAND U36163 ( .A(n26849), .B(n26850), .Z(c[913]) );
  NAND U36164 ( .A(n26658), .B(o[913]), .Z(n26850) );
  NAND U36165 ( .A(n26653), .B(creg[913]), .Z(n26849) );
  NAND U36166 ( .A(n26851), .B(n26852), .Z(c[912]) );
  NAND U36167 ( .A(n26658), .B(o[912]), .Z(n26852) );
  NAND U36168 ( .A(n26653), .B(creg[912]), .Z(n26851) );
  NAND U36169 ( .A(n26853), .B(n26854), .Z(c[911]) );
  NAND U36170 ( .A(n26658), .B(o[911]), .Z(n26854) );
  NAND U36171 ( .A(n26653), .B(creg[911]), .Z(n26853) );
  NAND U36172 ( .A(n26855), .B(n26856), .Z(c[910]) );
  NAND U36173 ( .A(n26658), .B(o[910]), .Z(n26856) );
  NAND U36174 ( .A(n26653), .B(creg[910]), .Z(n26855) );
  NAND U36175 ( .A(n26857), .B(n26858), .Z(c[90]) );
  NAND U36176 ( .A(n26658), .B(o[90]), .Z(n26858) );
  NAND U36177 ( .A(n26653), .B(creg[90]), .Z(n26857) );
  NAND U36178 ( .A(n26859), .B(n26860), .Z(c[909]) );
  NAND U36179 ( .A(n26658), .B(o[909]), .Z(n26860) );
  NAND U36180 ( .A(n26653), .B(creg[909]), .Z(n26859) );
  NAND U36181 ( .A(n26861), .B(n26862), .Z(c[908]) );
  NAND U36182 ( .A(n26658), .B(o[908]), .Z(n26862) );
  NAND U36183 ( .A(n26653), .B(creg[908]), .Z(n26861) );
  NAND U36184 ( .A(n26863), .B(n26864), .Z(c[907]) );
  NAND U36185 ( .A(n26658), .B(o[907]), .Z(n26864) );
  NAND U36186 ( .A(n26653), .B(creg[907]), .Z(n26863) );
  NAND U36187 ( .A(n26865), .B(n26866), .Z(c[906]) );
  NAND U36188 ( .A(n26658), .B(o[906]), .Z(n26866) );
  NAND U36189 ( .A(n26653), .B(creg[906]), .Z(n26865) );
  NAND U36190 ( .A(n26867), .B(n26868), .Z(c[905]) );
  NAND U36191 ( .A(n26658), .B(o[905]), .Z(n26868) );
  NAND U36192 ( .A(n26653), .B(creg[905]), .Z(n26867) );
  NAND U36193 ( .A(n26869), .B(n26870), .Z(c[904]) );
  NAND U36194 ( .A(n26658), .B(o[904]), .Z(n26870) );
  NAND U36195 ( .A(n26653), .B(creg[904]), .Z(n26869) );
  NAND U36196 ( .A(n26871), .B(n26872), .Z(c[903]) );
  NAND U36197 ( .A(n26658), .B(o[903]), .Z(n26872) );
  NAND U36198 ( .A(n26653), .B(creg[903]), .Z(n26871) );
  NAND U36199 ( .A(n26873), .B(n26874), .Z(c[902]) );
  NAND U36200 ( .A(n26658), .B(o[902]), .Z(n26874) );
  NAND U36201 ( .A(n26653), .B(creg[902]), .Z(n26873) );
  NAND U36202 ( .A(n26875), .B(n26876), .Z(c[901]) );
  NAND U36203 ( .A(n26658), .B(o[901]), .Z(n26876) );
  NAND U36204 ( .A(n26653), .B(creg[901]), .Z(n26875) );
  NAND U36205 ( .A(n26877), .B(n26878), .Z(c[900]) );
  NAND U36206 ( .A(n26658), .B(o[900]), .Z(n26878) );
  NAND U36207 ( .A(n26653), .B(creg[900]), .Z(n26877) );
  NAND U36208 ( .A(n26879), .B(n26880), .Z(c[8]) );
  NAND U36209 ( .A(n26658), .B(o[8]), .Z(n26880) );
  NAND U36210 ( .A(n26653), .B(creg[8]), .Z(n26879) );
  NAND U36211 ( .A(n26881), .B(n26882), .Z(c[89]) );
  NAND U36212 ( .A(n26658), .B(o[89]), .Z(n26882) );
  NAND U36213 ( .A(n26653), .B(creg[89]), .Z(n26881) );
  NAND U36214 ( .A(n26883), .B(n26884), .Z(c[899]) );
  NAND U36215 ( .A(n26658), .B(o[899]), .Z(n26884) );
  NAND U36216 ( .A(n26653), .B(creg[899]), .Z(n26883) );
  NAND U36217 ( .A(n26885), .B(n26886), .Z(c[898]) );
  NAND U36218 ( .A(n26658), .B(o[898]), .Z(n26886) );
  NAND U36219 ( .A(n26653), .B(creg[898]), .Z(n26885) );
  NAND U36220 ( .A(n26887), .B(n26888), .Z(c[897]) );
  NAND U36221 ( .A(n26658), .B(o[897]), .Z(n26888) );
  NAND U36222 ( .A(n26653), .B(creg[897]), .Z(n26887) );
  NAND U36223 ( .A(n26889), .B(n26890), .Z(c[896]) );
  NAND U36224 ( .A(n26658), .B(o[896]), .Z(n26890) );
  NAND U36225 ( .A(n26653), .B(creg[896]), .Z(n26889) );
  NAND U36226 ( .A(n26891), .B(n26892), .Z(c[895]) );
  NAND U36227 ( .A(n26658), .B(o[895]), .Z(n26892) );
  NAND U36228 ( .A(n26653), .B(creg[895]), .Z(n26891) );
  NAND U36229 ( .A(n26893), .B(n26894), .Z(c[894]) );
  NAND U36230 ( .A(n26658), .B(o[894]), .Z(n26894) );
  NAND U36231 ( .A(n26653), .B(creg[894]), .Z(n26893) );
  NAND U36232 ( .A(n26895), .B(n26896), .Z(c[893]) );
  NAND U36233 ( .A(n26658), .B(o[893]), .Z(n26896) );
  NAND U36234 ( .A(n26653), .B(creg[893]), .Z(n26895) );
  NAND U36235 ( .A(n26897), .B(n26898), .Z(c[892]) );
  NAND U36236 ( .A(n26658), .B(o[892]), .Z(n26898) );
  NAND U36237 ( .A(n26653), .B(creg[892]), .Z(n26897) );
  NAND U36238 ( .A(n26899), .B(n26900), .Z(c[891]) );
  NAND U36239 ( .A(n26658), .B(o[891]), .Z(n26900) );
  NAND U36240 ( .A(n26653), .B(creg[891]), .Z(n26899) );
  NAND U36241 ( .A(n26901), .B(n26902), .Z(c[890]) );
  NAND U36242 ( .A(n26658), .B(o[890]), .Z(n26902) );
  NAND U36243 ( .A(n26653), .B(creg[890]), .Z(n26901) );
  NAND U36244 ( .A(n26903), .B(n26904), .Z(c[88]) );
  NAND U36245 ( .A(n26658), .B(o[88]), .Z(n26904) );
  NAND U36246 ( .A(n26653), .B(creg[88]), .Z(n26903) );
  NAND U36247 ( .A(n26905), .B(n26906), .Z(c[889]) );
  NAND U36248 ( .A(n26658), .B(o[889]), .Z(n26906) );
  NAND U36249 ( .A(n26653), .B(creg[889]), .Z(n26905) );
  NAND U36250 ( .A(n26907), .B(n26908), .Z(c[888]) );
  NAND U36251 ( .A(n26658), .B(o[888]), .Z(n26908) );
  NAND U36252 ( .A(n26653), .B(creg[888]), .Z(n26907) );
  NAND U36253 ( .A(n26909), .B(n26910), .Z(c[887]) );
  NAND U36254 ( .A(n26658), .B(o[887]), .Z(n26910) );
  NAND U36255 ( .A(n26653), .B(creg[887]), .Z(n26909) );
  NAND U36256 ( .A(n26911), .B(n26912), .Z(c[886]) );
  NAND U36257 ( .A(n26658), .B(o[886]), .Z(n26912) );
  NAND U36258 ( .A(n26653), .B(creg[886]), .Z(n26911) );
  NAND U36259 ( .A(n26913), .B(n26914), .Z(c[885]) );
  NAND U36260 ( .A(n26658), .B(o[885]), .Z(n26914) );
  NAND U36261 ( .A(n26653), .B(creg[885]), .Z(n26913) );
  NAND U36262 ( .A(n26915), .B(n26916), .Z(c[884]) );
  NAND U36263 ( .A(n26658), .B(o[884]), .Z(n26916) );
  NAND U36264 ( .A(n26653), .B(creg[884]), .Z(n26915) );
  NAND U36265 ( .A(n26917), .B(n26918), .Z(c[883]) );
  NAND U36266 ( .A(n26658), .B(o[883]), .Z(n26918) );
  NAND U36267 ( .A(n26653), .B(creg[883]), .Z(n26917) );
  NAND U36268 ( .A(n26919), .B(n26920), .Z(c[882]) );
  NAND U36269 ( .A(n26658), .B(o[882]), .Z(n26920) );
  NAND U36270 ( .A(n26653), .B(creg[882]), .Z(n26919) );
  NAND U36271 ( .A(n26921), .B(n26922), .Z(c[881]) );
  NAND U36272 ( .A(n26658), .B(o[881]), .Z(n26922) );
  NAND U36273 ( .A(n26653), .B(creg[881]), .Z(n26921) );
  NAND U36274 ( .A(n26923), .B(n26924), .Z(c[880]) );
  NAND U36275 ( .A(n26658), .B(o[880]), .Z(n26924) );
  NAND U36276 ( .A(n26653), .B(creg[880]), .Z(n26923) );
  NAND U36277 ( .A(n26925), .B(n26926), .Z(c[87]) );
  NAND U36278 ( .A(n26658), .B(o[87]), .Z(n26926) );
  NAND U36279 ( .A(n26653), .B(creg[87]), .Z(n26925) );
  NAND U36280 ( .A(n26927), .B(n26928), .Z(c[879]) );
  NAND U36281 ( .A(n26658), .B(o[879]), .Z(n26928) );
  NAND U36282 ( .A(n26653), .B(creg[879]), .Z(n26927) );
  NAND U36283 ( .A(n26929), .B(n26930), .Z(c[878]) );
  NAND U36284 ( .A(n26658), .B(o[878]), .Z(n26930) );
  NAND U36285 ( .A(n26653), .B(creg[878]), .Z(n26929) );
  NAND U36286 ( .A(n26931), .B(n26932), .Z(c[877]) );
  NAND U36287 ( .A(n26658), .B(o[877]), .Z(n26932) );
  NAND U36288 ( .A(n26653), .B(creg[877]), .Z(n26931) );
  NAND U36289 ( .A(n26933), .B(n26934), .Z(c[876]) );
  NAND U36290 ( .A(n26658), .B(o[876]), .Z(n26934) );
  NAND U36291 ( .A(n26653), .B(creg[876]), .Z(n26933) );
  NAND U36292 ( .A(n26935), .B(n26936), .Z(c[875]) );
  NAND U36293 ( .A(n26658), .B(o[875]), .Z(n26936) );
  NAND U36294 ( .A(n26653), .B(creg[875]), .Z(n26935) );
  NAND U36295 ( .A(n26937), .B(n26938), .Z(c[874]) );
  NAND U36296 ( .A(n26658), .B(o[874]), .Z(n26938) );
  NAND U36297 ( .A(n26653), .B(creg[874]), .Z(n26937) );
  NAND U36298 ( .A(n26939), .B(n26940), .Z(c[873]) );
  NAND U36299 ( .A(n26658), .B(o[873]), .Z(n26940) );
  NAND U36300 ( .A(n26653), .B(creg[873]), .Z(n26939) );
  NAND U36301 ( .A(n26941), .B(n26942), .Z(c[872]) );
  NAND U36302 ( .A(n26658), .B(o[872]), .Z(n26942) );
  NAND U36303 ( .A(n26653), .B(creg[872]), .Z(n26941) );
  NAND U36304 ( .A(n26943), .B(n26944), .Z(c[871]) );
  NAND U36305 ( .A(n26658), .B(o[871]), .Z(n26944) );
  NAND U36306 ( .A(n26653), .B(creg[871]), .Z(n26943) );
  NAND U36307 ( .A(n26945), .B(n26946), .Z(c[870]) );
  NAND U36308 ( .A(n26658), .B(o[870]), .Z(n26946) );
  NAND U36309 ( .A(n26653), .B(creg[870]), .Z(n26945) );
  NAND U36310 ( .A(n26947), .B(n26948), .Z(c[86]) );
  NAND U36311 ( .A(n26658), .B(o[86]), .Z(n26948) );
  NAND U36312 ( .A(n26653), .B(creg[86]), .Z(n26947) );
  NAND U36313 ( .A(n26949), .B(n26950), .Z(c[869]) );
  NAND U36314 ( .A(n26658), .B(o[869]), .Z(n26950) );
  NAND U36315 ( .A(n26653), .B(creg[869]), .Z(n26949) );
  NAND U36316 ( .A(n26951), .B(n26952), .Z(c[868]) );
  NAND U36317 ( .A(n26658), .B(o[868]), .Z(n26952) );
  NAND U36318 ( .A(n26653), .B(creg[868]), .Z(n26951) );
  NAND U36319 ( .A(n26953), .B(n26954), .Z(c[867]) );
  NAND U36320 ( .A(n26658), .B(o[867]), .Z(n26954) );
  NAND U36321 ( .A(n26653), .B(creg[867]), .Z(n26953) );
  NAND U36322 ( .A(n26955), .B(n26956), .Z(c[866]) );
  NAND U36323 ( .A(n26658), .B(o[866]), .Z(n26956) );
  NAND U36324 ( .A(n26653), .B(creg[866]), .Z(n26955) );
  NAND U36325 ( .A(n26957), .B(n26958), .Z(c[865]) );
  NAND U36326 ( .A(n26658), .B(o[865]), .Z(n26958) );
  NAND U36327 ( .A(n26653), .B(creg[865]), .Z(n26957) );
  NAND U36328 ( .A(n26959), .B(n26960), .Z(c[864]) );
  NAND U36329 ( .A(n26658), .B(o[864]), .Z(n26960) );
  NAND U36330 ( .A(n26653), .B(creg[864]), .Z(n26959) );
  NAND U36331 ( .A(n26961), .B(n26962), .Z(c[863]) );
  NAND U36332 ( .A(n26658), .B(o[863]), .Z(n26962) );
  NAND U36333 ( .A(n26653), .B(creg[863]), .Z(n26961) );
  NAND U36334 ( .A(n26963), .B(n26964), .Z(c[862]) );
  NAND U36335 ( .A(n26658), .B(o[862]), .Z(n26964) );
  NAND U36336 ( .A(n26653), .B(creg[862]), .Z(n26963) );
  NAND U36337 ( .A(n26965), .B(n26966), .Z(c[861]) );
  NAND U36338 ( .A(n26658), .B(o[861]), .Z(n26966) );
  NAND U36339 ( .A(n26653), .B(creg[861]), .Z(n26965) );
  NAND U36340 ( .A(n26967), .B(n26968), .Z(c[860]) );
  NAND U36341 ( .A(n26658), .B(o[860]), .Z(n26968) );
  NAND U36342 ( .A(n26653), .B(creg[860]), .Z(n26967) );
  NAND U36343 ( .A(n26969), .B(n26970), .Z(c[85]) );
  NAND U36344 ( .A(n26658), .B(o[85]), .Z(n26970) );
  NAND U36345 ( .A(n26653), .B(creg[85]), .Z(n26969) );
  NAND U36346 ( .A(n26971), .B(n26972), .Z(c[859]) );
  NAND U36347 ( .A(n26658), .B(o[859]), .Z(n26972) );
  NAND U36348 ( .A(n26653), .B(creg[859]), .Z(n26971) );
  NAND U36349 ( .A(n26973), .B(n26974), .Z(c[858]) );
  NAND U36350 ( .A(n26658), .B(o[858]), .Z(n26974) );
  NAND U36351 ( .A(n26653), .B(creg[858]), .Z(n26973) );
  NAND U36352 ( .A(n26975), .B(n26976), .Z(c[857]) );
  NAND U36353 ( .A(n26658), .B(o[857]), .Z(n26976) );
  NAND U36354 ( .A(n26653), .B(creg[857]), .Z(n26975) );
  NAND U36355 ( .A(n26977), .B(n26978), .Z(c[856]) );
  NAND U36356 ( .A(n26658), .B(o[856]), .Z(n26978) );
  NAND U36357 ( .A(n26653), .B(creg[856]), .Z(n26977) );
  NAND U36358 ( .A(n26979), .B(n26980), .Z(c[855]) );
  NAND U36359 ( .A(n26658), .B(o[855]), .Z(n26980) );
  NAND U36360 ( .A(n26653), .B(creg[855]), .Z(n26979) );
  NAND U36361 ( .A(n26981), .B(n26982), .Z(c[854]) );
  NAND U36362 ( .A(n26658), .B(o[854]), .Z(n26982) );
  NAND U36363 ( .A(n26653), .B(creg[854]), .Z(n26981) );
  NAND U36364 ( .A(n26983), .B(n26984), .Z(c[853]) );
  NAND U36365 ( .A(n26658), .B(o[853]), .Z(n26984) );
  NAND U36366 ( .A(n26653), .B(creg[853]), .Z(n26983) );
  NAND U36367 ( .A(n26985), .B(n26986), .Z(c[852]) );
  NAND U36368 ( .A(n26658), .B(o[852]), .Z(n26986) );
  NAND U36369 ( .A(n26653), .B(creg[852]), .Z(n26985) );
  NAND U36370 ( .A(n26987), .B(n26988), .Z(c[851]) );
  NAND U36371 ( .A(n26658), .B(o[851]), .Z(n26988) );
  NAND U36372 ( .A(n26653), .B(creg[851]), .Z(n26987) );
  NAND U36373 ( .A(n26989), .B(n26990), .Z(c[850]) );
  NAND U36374 ( .A(n26658), .B(o[850]), .Z(n26990) );
  NAND U36375 ( .A(n26653), .B(creg[850]), .Z(n26989) );
  NAND U36376 ( .A(n26991), .B(n26992), .Z(c[84]) );
  NAND U36377 ( .A(n26658), .B(o[84]), .Z(n26992) );
  NAND U36378 ( .A(n26653), .B(creg[84]), .Z(n26991) );
  NAND U36379 ( .A(n26993), .B(n26994), .Z(c[849]) );
  NAND U36380 ( .A(n26658), .B(o[849]), .Z(n26994) );
  NAND U36381 ( .A(n26653), .B(creg[849]), .Z(n26993) );
  NAND U36382 ( .A(n26995), .B(n26996), .Z(c[848]) );
  NAND U36383 ( .A(n26658), .B(o[848]), .Z(n26996) );
  NAND U36384 ( .A(n26653), .B(creg[848]), .Z(n26995) );
  NAND U36385 ( .A(n26997), .B(n26998), .Z(c[847]) );
  NAND U36386 ( .A(n26658), .B(o[847]), .Z(n26998) );
  NAND U36387 ( .A(n26653), .B(creg[847]), .Z(n26997) );
  NAND U36388 ( .A(n26999), .B(n27000), .Z(c[846]) );
  NAND U36389 ( .A(n26658), .B(o[846]), .Z(n27000) );
  NAND U36390 ( .A(n26653), .B(creg[846]), .Z(n26999) );
  NAND U36391 ( .A(n27001), .B(n27002), .Z(c[845]) );
  NAND U36392 ( .A(n26658), .B(o[845]), .Z(n27002) );
  NAND U36393 ( .A(n26653), .B(creg[845]), .Z(n27001) );
  NAND U36394 ( .A(n27003), .B(n27004), .Z(c[844]) );
  NAND U36395 ( .A(n26658), .B(o[844]), .Z(n27004) );
  NAND U36396 ( .A(n26653), .B(creg[844]), .Z(n27003) );
  NAND U36397 ( .A(n27005), .B(n27006), .Z(c[843]) );
  NAND U36398 ( .A(n26658), .B(o[843]), .Z(n27006) );
  NAND U36399 ( .A(n26653), .B(creg[843]), .Z(n27005) );
  NAND U36400 ( .A(n27007), .B(n27008), .Z(c[842]) );
  NAND U36401 ( .A(n26658), .B(o[842]), .Z(n27008) );
  NAND U36402 ( .A(n26653), .B(creg[842]), .Z(n27007) );
  NAND U36403 ( .A(n27009), .B(n27010), .Z(c[841]) );
  NAND U36404 ( .A(n26658), .B(o[841]), .Z(n27010) );
  NAND U36405 ( .A(n26653), .B(creg[841]), .Z(n27009) );
  NAND U36406 ( .A(n27011), .B(n27012), .Z(c[840]) );
  NAND U36407 ( .A(n26658), .B(o[840]), .Z(n27012) );
  NAND U36408 ( .A(n26653), .B(creg[840]), .Z(n27011) );
  NAND U36409 ( .A(n27013), .B(n27014), .Z(c[83]) );
  NAND U36410 ( .A(n26658), .B(o[83]), .Z(n27014) );
  NAND U36411 ( .A(n26653), .B(creg[83]), .Z(n27013) );
  NAND U36412 ( .A(n27015), .B(n27016), .Z(c[839]) );
  NAND U36413 ( .A(n26658), .B(o[839]), .Z(n27016) );
  NAND U36414 ( .A(n26653), .B(creg[839]), .Z(n27015) );
  NAND U36415 ( .A(n27017), .B(n27018), .Z(c[838]) );
  NAND U36416 ( .A(n26658), .B(o[838]), .Z(n27018) );
  NAND U36417 ( .A(n26653), .B(creg[838]), .Z(n27017) );
  NAND U36418 ( .A(n27019), .B(n27020), .Z(c[837]) );
  NAND U36419 ( .A(n26658), .B(o[837]), .Z(n27020) );
  NAND U36420 ( .A(n26653), .B(creg[837]), .Z(n27019) );
  NAND U36421 ( .A(n27021), .B(n27022), .Z(c[836]) );
  NAND U36422 ( .A(n26658), .B(o[836]), .Z(n27022) );
  NAND U36423 ( .A(n26653), .B(creg[836]), .Z(n27021) );
  NAND U36424 ( .A(n27023), .B(n27024), .Z(c[835]) );
  NAND U36425 ( .A(n26658), .B(o[835]), .Z(n27024) );
  NAND U36426 ( .A(n26653), .B(creg[835]), .Z(n27023) );
  NAND U36427 ( .A(n27025), .B(n27026), .Z(c[834]) );
  NAND U36428 ( .A(n26658), .B(o[834]), .Z(n27026) );
  NAND U36429 ( .A(n26653), .B(creg[834]), .Z(n27025) );
  NAND U36430 ( .A(n27027), .B(n27028), .Z(c[833]) );
  NAND U36431 ( .A(n26658), .B(o[833]), .Z(n27028) );
  NAND U36432 ( .A(n26653), .B(creg[833]), .Z(n27027) );
  NAND U36433 ( .A(n27029), .B(n27030), .Z(c[832]) );
  NAND U36434 ( .A(n26658), .B(o[832]), .Z(n27030) );
  NAND U36435 ( .A(n26653), .B(creg[832]), .Z(n27029) );
  NAND U36436 ( .A(n27031), .B(n27032), .Z(c[831]) );
  NAND U36437 ( .A(n26658), .B(o[831]), .Z(n27032) );
  NAND U36438 ( .A(n26653), .B(creg[831]), .Z(n27031) );
  NAND U36439 ( .A(n27033), .B(n27034), .Z(c[830]) );
  NAND U36440 ( .A(n26658), .B(o[830]), .Z(n27034) );
  NAND U36441 ( .A(n26653), .B(creg[830]), .Z(n27033) );
  NAND U36442 ( .A(n27035), .B(n27036), .Z(c[82]) );
  NAND U36443 ( .A(n26658), .B(o[82]), .Z(n27036) );
  NAND U36444 ( .A(n26653), .B(creg[82]), .Z(n27035) );
  NAND U36445 ( .A(n27037), .B(n27038), .Z(c[829]) );
  NAND U36446 ( .A(n26658), .B(o[829]), .Z(n27038) );
  NAND U36447 ( .A(n26653), .B(creg[829]), .Z(n27037) );
  NAND U36448 ( .A(n27039), .B(n27040), .Z(c[828]) );
  NAND U36449 ( .A(n26658), .B(o[828]), .Z(n27040) );
  NAND U36450 ( .A(n26653), .B(creg[828]), .Z(n27039) );
  NAND U36451 ( .A(n27041), .B(n27042), .Z(c[827]) );
  NAND U36452 ( .A(n26658), .B(o[827]), .Z(n27042) );
  NAND U36453 ( .A(n26653), .B(creg[827]), .Z(n27041) );
  NAND U36454 ( .A(n27043), .B(n27044), .Z(c[826]) );
  NAND U36455 ( .A(n26658), .B(o[826]), .Z(n27044) );
  NAND U36456 ( .A(n26653), .B(creg[826]), .Z(n27043) );
  NAND U36457 ( .A(n27045), .B(n27046), .Z(c[825]) );
  NAND U36458 ( .A(n26658), .B(o[825]), .Z(n27046) );
  NAND U36459 ( .A(n26653), .B(creg[825]), .Z(n27045) );
  NAND U36460 ( .A(n27047), .B(n27048), .Z(c[824]) );
  NAND U36461 ( .A(n26658), .B(o[824]), .Z(n27048) );
  NAND U36462 ( .A(n26653), .B(creg[824]), .Z(n27047) );
  NAND U36463 ( .A(n27049), .B(n27050), .Z(c[823]) );
  NAND U36464 ( .A(n26658), .B(o[823]), .Z(n27050) );
  NAND U36465 ( .A(n26653), .B(creg[823]), .Z(n27049) );
  NAND U36466 ( .A(n27051), .B(n27052), .Z(c[822]) );
  NAND U36467 ( .A(n26658), .B(o[822]), .Z(n27052) );
  NAND U36468 ( .A(n26653), .B(creg[822]), .Z(n27051) );
  NAND U36469 ( .A(n27053), .B(n27054), .Z(c[821]) );
  NAND U36470 ( .A(n26658), .B(o[821]), .Z(n27054) );
  NAND U36471 ( .A(n26653), .B(creg[821]), .Z(n27053) );
  NAND U36472 ( .A(n27055), .B(n27056), .Z(c[820]) );
  NAND U36473 ( .A(n26658), .B(o[820]), .Z(n27056) );
  NAND U36474 ( .A(n26653), .B(creg[820]), .Z(n27055) );
  NAND U36475 ( .A(n27057), .B(n27058), .Z(c[81]) );
  NAND U36476 ( .A(n26658), .B(o[81]), .Z(n27058) );
  NAND U36477 ( .A(n26653), .B(creg[81]), .Z(n27057) );
  NAND U36478 ( .A(n27059), .B(n27060), .Z(c[819]) );
  NAND U36479 ( .A(n26658), .B(o[819]), .Z(n27060) );
  NAND U36480 ( .A(n26653), .B(creg[819]), .Z(n27059) );
  NAND U36481 ( .A(n27061), .B(n27062), .Z(c[818]) );
  NAND U36482 ( .A(n26658), .B(o[818]), .Z(n27062) );
  NAND U36483 ( .A(n26653), .B(creg[818]), .Z(n27061) );
  NAND U36484 ( .A(n27063), .B(n27064), .Z(c[817]) );
  NAND U36485 ( .A(n26658), .B(o[817]), .Z(n27064) );
  NAND U36486 ( .A(n26653), .B(creg[817]), .Z(n27063) );
  NAND U36487 ( .A(n27065), .B(n27066), .Z(c[816]) );
  NAND U36488 ( .A(n26658), .B(o[816]), .Z(n27066) );
  NAND U36489 ( .A(n26653), .B(creg[816]), .Z(n27065) );
  NAND U36490 ( .A(n27067), .B(n27068), .Z(c[815]) );
  NAND U36491 ( .A(n26658), .B(o[815]), .Z(n27068) );
  NAND U36492 ( .A(n26653), .B(creg[815]), .Z(n27067) );
  NAND U36493 ( .A(n27069), .B(n27070), .Z(c[814]) );
  NAND U36494 ( .A(n26658), .B(o[814]), .Z(n27070) );
  NAND U36495 ( .A(n26653), .B(creg[814]), .Z(n27069) );
  NAND U36496 ( .A(n27071), .B(n27072), .Z(c[813]) );
  NAND U36497 ( .A(n26658), .B(o[813]), .Z(n27072) );
  NAND U36498 ( .A(n26653), .B(creg[813]), .Z(n27071) );
  NAND U36499 ( .A(n27073), .B(n27074), .Z(c[812]) );
  NAND U36500 ( .A(n26658), .B(o[812]), .Z(n27074) );
  NAND U36501 ( .A(n26653), .B(creg[812]), .Z(n27073) );
  NAND U36502 ( .A(n27075), .B(n27076), .Z(c[811]) );
  NAND U36503 ( .A(n26658), .B(o[811]), .Z(n27076) );
  NAND U36504 ( .A(n26653), .B(creg[811]), .Z(n27075) );
  NAND U36505 ( .A(n27077), .B(n27078), .Z(c[810]) );
  NAND U36506 ( .A(n26658), .B(o[810]), .Z(n27078) );
  NAND U36507 ( .A(n26653), .B(creg[810]), .Z(n27077) );
  NAND U36508 ( .A(n27079), .B(n27080), .Z(c[80]) );
  NAND U36509 ( .A(n26658), .B(o[80]), .Z(n27080) );
  NAND U36510 ( .A(n26653), .B(creg[80]), .Z(n27079) );
  NAND U36511 ( .A(n27081), .B(n27082), .Z(c[809]) );
  NAND U36512 ( .A(n26658), .B(o[809]), .Z(n27082) );
  NAND U36513 ( .A(n26653), .B(creg[809]), .Z(n27081) );
  NAND U36514 ( .A(n27083), .B(n27084), .Z(c[808]) );
  NAND U36515 ( .A(n26658), .B(o[808]), .Z(n27084) );
  NAND U36516 ( .A(n26653), .B(creg[808]), .Z(n27083) );
  NAND U36517 ( .A(n27085), .B(n27086), .Z(c[807]) );
  NAND U36518 ( .A(n26658), .B(o[807]), .Z(n27086) );
  NAND U36519 ( .A(n26653), .B(creg[807]), .Z(n27085) );
  NAND U36520 ( .A(n27087), .B(n27088), .Z(c[806]) );
  NAND U36521 ( .A(n26658), .B(o[806]), .Z(n27088) );
  NAND U36522 ( .A(n26653), .B(creg[806]), .Z(n27087) );
  NAND U36523 ( .A(n27089), .B(n27090), .Z(c[805]) );
  NAND U36524 ( .A(n26658), .B(o[805]), .Z(n27090) );
  NAND U36525 ( .A(n26653), .B(creg[805]), .Z(n27089) );
  NAND U36526 ( .A(n27091), .B(n27092), .Z(c[804]) );
  NAND U36527 ( .A(n26658), .B(o[804]), .Z(n27092) );
  NAND U36528 ( .A(n26653), .B(creg[804]), .Z(n27091) );
  NAND U36529 ( .A(n27093), .B(n27094), .Z(c[803]) );
  NAND U36530 ( .A(n26658), .B(o[803]), .Z(n27094) );
  NAND U36531 ( .A(n26653), .B(creg[803]), .Z(n27093) );
  NAND U36532 ( .A(n27095), .B(n27096), .Z(c[802]) );
  NAND U36533 ( .A(n26658), .B(o[802]), .Z(n27096) );
  NAND U36534 ( .A(n26653), .B(creg[802]), .Z(n27095) );
  NAND U36535 ( .A(n27097), .B(n27098), .Z(c[801]) );
  NAND U36536 ( .A(n26658), .B(o[801]), .Z(n27098) );
  NAND U36537 ( .A(n26653), .B(creg[801]), .Z(n27097) );
  NAND U36538 ( .A(n27099), .B(n27100), .Z(c[800]) );
  NAND U36539 ( .A(n26658), .B(o[800]), .Z(n27100) );
  NAND U36540 ( .A(n26653), .B(creg[800]), .Z(n27099) );
  NAND U36541 ( .A(n27101), .B(n27102), .Z(c[7]) );
  NAND U36542 ( .A(n26658), .B(o[7]), .Z(n27102) );
  NAND U36543 ( .A(n26653), .B(creg[7]), .Z(n27101) );
  NAND U36544 ( .A(n27103), .B(n27104), .Z(c[79]) );
  NAND U36545 ( .A(n26658), .B(o[79]), .Z(n27104) );
  NAND U36546 ( .A(n26653), .B(creg[79]), .Z(n27103) );
  NAND U36547 ( .A(n27105), .B(n27106), .Z(c[799]) );
  NAND U36548 ( .A(n26658), .B(o[799]), .Z(n27106) );
  NAND U36549 ( .A(n26653), .B(creg[799]), .Z(n27105) );
  NAND U36550 ( .A(n27107), .B(n27108), .Z(c[798]) );
  NAND U36551 ( .A(n26658), .B(o[798]), .Z(n27108) );
  NAND U36552 ( .A(n26653), .B(creg[798]), .Z(n27107) );
  NAND U36553 ( .A(n27109), .B(n27110), .Z(c[797]) );
  NAND U36554 ( .A(n26658), .B(o[797]), .Z(n27110) );
  NAND U36555 ( .A(n26653), .B(creg[797]), .Z(n27109) );
  NAND U36556 ( .A(n27111), .B(n27112), .Z(c[796]) );
  NAND U36557 ( .A(n26658), .B(o[796]), .Z(n27112) );
  NAND U36558 ( .A(n26653), .B(creg[796]), .Z(n27111) );
  NAND U36559 ( .A(n27113), .B(n27114), .Z(c[795]) );
  NAND U36560 ( .A(n26658), .B(o[795]), .Z(n27114) );
  NAND U36561 ( .A(n26653), .B(creg[795]), .Z(n27113) );
  NAND U36562 ( .A(n27115), .B(n27116), .Z(c[794]) );
  NAND U36563 ( .A(n26658), .B(o[794]), .Z(n27116) );
  NAND U36564 ( .A(n26653), .B(creg[794]), .Z(n27115) );
  NAND U36565 ( .A(n27117), .B(n27118), .Z(c[793]) );
  NAND U36566 ( .A(n26658), .B(o[793]), .Z(n27118) );
  NAND U36567 ( .A(n26653), .B(creg[793]), .Z(n27117) );
  NAND U36568 ( .A(n27119), .B(n27120), .Z(c[792]) );
  NAND U36569 ( .A(n26658), .B(o[792]), .Z(n27120) );
  NAND U36570 ( .A(n26653), .B(creg[792]), .Z(n27119) );
  NAND U36571 ( .A(n27121), .B(n27122), .Z(c[791]) );
  NAND U36572 ( .A(n26658), .B(o[791]), .Z(n27122) );
  NAND U36573 ( .A(n26653), .B(creg[791]), .Z(n27121) );
  NAND U36574 ( .A(n27123), .B(n27124), .Z(c[790]) );
  NAND U36575 ( .A(n26658), .B(o[790]), .Z(n27124) );
  NAND U36576 ( .A(n26653), .B(creg[790]), .Z(n27123) );
  NAND U36577 ( .A(n27125), .B(n27126), .Z(c[78]) );
  NAND U36578 ( .A(n26658), .B(o[78]), .Z(n27126) );
  NAND U36579 ( .A(n26653), .B(creg[78]), .Z(n27125) );
  NAND U36580 ( .A(n27127), .B(n27128), .Z(c[789]) );
  NAND U36581 ( .A(n26658), .B(o[789]), .Z(n27128) );
  NAND U36582 ( .A(n26653), .B(creg[789]), .Z(n27127) );
  NAND U36583 ( .A(n27129), .B(n27130), .Z(c[788]) );
  NAND U36584 ( .A(n26658), .B(o[788]), .Z(n27130) );
  NAND U36585 ( .A(n26653), .B(creg[788]), .Z(n27129) );
  NAND U36586 ( .A(n27131), .B(n27132), .Z(c[787]) );
  NAND U36587 ( .A(n26658), .B(o[787]), .Z(n27132) );
  NAND U36588 ( .A(n26653), .B(creg[787]), .Z(n27131) );
  NAND U36589 ( .A(n27133), .B(n27134), .Z(c[786]) );
  NAND U36590 ( .A(n26658), .B(o[786]), .Z(n27134) );
  NAND U36591 ( .A(n26653), .B(creg[786]), .Z(n27133) );
  NAND U36592 ( .A(n27135), .B(n27136), .Z(c[785]) );
  NAND U36593 ( .A(n26658), .B(o[785]), .Z(n27136) );
  NAND U36594 ( .A(n26653), .B(creg[785]), .Z(n27135) );
  NAND U36595 ( .A(n27137), .B(n27138), .Z(c[784]) );
  NAND U36596 ( .A(n26658), .B(o[784]), .Z(n27138) );
  NAND U36597 ( .A(n26653), .B(creg[784]), .Z(n27137) );
  NAND U36598 ( .A(n27139), .B(n27140), .Z(c[783]) );
  NAND U36599 ( .A(n26658), .B(o[783]), .Z(n27140) );
  NAND U36600 ( .A(n26653), .B(creg[783]), .Z(n27139) );
  NAND U36601 ( .A(n27141), .B(n27142), .Z(c[782]) );
  NAND U36602 ( .A(n26658), .B(o[782]), .Z(n27142) );
  NAND U36603 ( .A(n26653), .B(creg[782]), .Z(n27141) );
  NAND U36604 ( .A(n27143), .B(n27144), .Z(c[781]) );
  NAND U36605 ( .A(n26658), .B(o[781]), .Z(n27144) );
  NAND U36606 ( .A(n26653), .B(creg[781]), .Z(n27143) );
  NAND U36607 ( .A(n27145), .B(n27146), .Z(c[780]) );
  NAND U36608 ( .A(n26658), .B(o[780]), .Z(n27146) );
  NAND U36609 ( .A(n26653), .B(creg[780]), .Z(n27145) );
  NAND U36610 ( .A(n27147), .B(n27148), .Z(c[77]) );
  NAND U36611 ( .A(n26658), .B(o[77]), .Z(n27148) );
  NAND U36612 ( .A(n26653), .B(creg[77]), .Z(n27147) );
  NAND U36613 ( .A(n27149), .B(n27150), .Z(c[779]) );
  NAND U36614 ( .A(n26658), .B(o[779]), .Z(n27150) );
  NAND U36615 ( .A(n26653), .B(creg[779]), .Z(n27149) );
  NAND U36616 ( .A(n27151), .B(n27152), .Z(c[778]) );
  NAND U36617 ( .A(n26658), .B(o[778]), .Z(n27152) );
  NAND U36618 ( .A(n26653), .B(creg[778]), .Z(n27151) );
  NAND U36619 ( .A(n27153), .B(n27154), .Z(c[777]) );
  NAND U36620 ( .A(n26658), .B(o[777]), .Z(n27154) );
  NAND U36621 ( .A(n26653), .B(creg[777]), .Z(n27153) );
  NAND U36622 ( .A(n27155), .B(n27156), .Z(c[776]) );
  NAND U36623 ( .A(n26658), .B(o[776]), .Z(n27156) );
  NAND U36624 ( .A(n26653), .B(creg[776]), .Z(n27155) );
  NAND U36625 ( .A(n27157), .B(n27158), .Z(c[775]) );
  NAND U36626 ( .A(n26658), .B(o[775]), .Z(n27158) );
  NAND U36627 ( .A(n26653), .B(creg[775]), .Z(n27157) );
  NAND U36628 ( .A(n27159), .B(n27160), .Z(c[774]) );
  NAND U36629 ( .A(n26658), .B(o[774]), .Z(n27160) );
  NAND U36630 ( .A(n26653), .B(creg[774]), .Z(n27159) );
  NAND U36631 ( .A(n27161), .B(n27162), .Z(c[773]) );
  NAND U36632 ( .A(n26658), .B(o[773]), .Z(n27162) );
  NAND U36633 ( .A(n26653), .B(creg[773]), .Z(n27161) );
  NAND U36634 ( .A(n27163), .B(n27164), .Z(c[772]) );
  NAND U36635 ( .A(n26658), .B(o[772]), .Z(n27164) );
  NAND U36636 ( .A(n26653), .B(creg[772]), .Z(n27163) );
  NAND U36637 ( .A(n27165), .B(n27166), .Z(c[771]) );
  NAND U36638 ( .A(n26658), .B(o[771]), .Z(n27166) );
  NAND U36639 ( .A(n26653), .B(creg[771]), .Z(n27165) );
  NAND U36640 ( .A(n27167), .B(n27168), .Z(c[770]) );
  NAND U36641 ( .A(n26658), .B(o[770]), .Z(n27168) );
  NAND U36642 ( .A(n26653), .B(creg[770]), .Z(n27167) );
  NAND U36643 ( .A(n27169), .B(n27170), .Z(c[76]) );
  NAND U36644 ( .A(n26658), .B(o[76]), .Z(n27170) );
  NAND U36645 ( .A(n26653), .B(creg[76]), .Z(n27169) );
  NAND U36646 ( .A(n27171), .B(n27172), .Z(c[769]) );
  NAND U36647 ( .A(n26658), .B(o[769]), .Z(n27172) );
  NAND U36648 ( .A(n26653), .B(creg[769]), .Z(n27171) );
  NAND U36649 ( .A(n27173), .B(n27174), .Z(c[768]) );
  NAND U36650 ( .A(n26658), .B(o[768]), .Z(n27174) );
  NAND U36651 ( .A(n26653), .B(creg[768]), .Z(n27173) );
  NAND U36652 ( .A(n27175), .B(n27176), .Z(c[767]) );
  NAND U36653 ( .A(n26658), .B(o[767]), .Z(n27176) );
  NAND U36654 ( .A(n26653), .B(creg[767]), .Z(n27175) );
  NAND U36655 ( .A(n27177), .B(n27178), .Z(c[766]) );
  NAND U36656 ( .A(n26658), .B(o[766]), .Z(n27178) );
  NAND U36657 ( .A(n26653), .B(creg[766]), .Z(n27177) );
  NAND U36658 ( .A(n27179), .B(n27180), .Z(c[765]) );
  NAND U36659 ( .A(n26658), .B(o[765]), .Z(n27180) );
  NAND U36660 ( .A(n26653), .B(creg[765]), .Z(n27179) );
  NAND U36661 ( .A(n27181), .B(n27182), .Z(c[764]) );
  NAND U36662 ( .A(n26658), .B(o[764]), .Z(n27182) );
  NAND U36663 ( .A(n26653), .B(creg[764]), .Z(n27181) );
  NAND U36664 ( .A(n27183), .B(n27184), .Z(c[763]) );
  NAND U36665 ( .A(n26658), .B(o[763]), .Z(n27184) );
  NAND U36666 ( .A(n26653), .B(creg[763]), .Z(n27183) );
  NAND U36667 ( .A(n27185), .B(n27186), .Z(c[762]) );
  NAND U36668 ( .A(n26658), .B(o[762]), .Z(n27186) );
  NAND U36669 ( .A(n26653), .B(creg[762]), .Z(n27185) );
  NAND U36670 ( .A(n27187), .B(n27188), .Z(c[761]) );
  NAND U36671 ( .A(n26658), .B(o[761]), .Z(n27188) );
  NAND U36672 ( .A(n26653), .B(creg[761]), .Z(n27187) );
  NAND U36673 ( .A(n27189), .B(n27190), .Z(c[760]) );
  NAND U36674 ( .A(n26658), .B(o[760]), .Z(n27190) );
  NAND U36675 ( .A(n26653), .B(creg[760]), .Z(n27189) );
  NAND U36676 ( .A(n27191), .B(n27192), .Z(c[75]) );
  NAND U36677 ( .A(n26658), .B(o[75]), .Z(n27192) );
  NAND U36678 ( .A(n26653), .B(creg[75]), .Z(n27191) );
  NAND U36679 ( .A(n27193), .B(n27194), .Z(c[759]) );
  NAND U36680 ( .A(n26658), .B(o[759]), .Z(n27194) );
  NAND U36681 ( .A(n26653), .B(creg[759]), .Z(n27193) );
  NAND U36682 ( .A(n27195), .B(n27196), .Z(c[758]) );
  NAND U36683 ( .A(n26658), .B(o[758]), .Z(n27196) );
  NAND U36684 ( .A(n26653), .B(creg[758]), .Z(n27195) );
  NAND U36685 ( .A(n27197), .B(n27198), .Z(c[757]) );
  NAND U36686 ( .A(n26658), .B(o[757]), .Z(n27198) );
  NAND U36687 ( .A(n26653), .B(creg[757]), .Z(n27197) );
  NAND U36688 ( .A(n27199), .B(n27200), .Z(c[756]) );
  NAND U36689 ( .A(n26658), .B(o[756]), .Z(n27200) );
  NAND U36690 ( .A(n26653), .B(creg[756]), .Z(n27199) );
  NAND U36691 ( .A(n27201), .B(n27202), .Z(c[755]) );
  NAND U36692 ( .A(n26658), .B(o[755]), .Z(n27202) );
  NAND U36693 ( .A(n26653), .B(creg[755]), .Z(n27201) );
  NAND U36694 ( .A(n27203), .B(n27204), .Z(c[754]) );
  NAND U36695 ( .A(n26658), .B(o[754]), .Z(n27204) );
  NAND U36696 ( .A(n26653), .B(creg[754]), .Z(n27203) );
  NAND U36697 ( .A(n27205), .B(n27206), .Z(c[753]) );
  NAND U36698 ( .A(n26658), .B(o[753]), .Z(n27206) );
  NAND U36699 ( .A(n26653), .B(creg[753]), .Z(n27205) );
  NAND U36700 ( .A(n27207), .B(n27208), .Z(c[752]) );
  NAND U36701 ( .A(n26658), .B(o[752]), .Z(n27208) );
  NAND U36702 ( .A(n26653), .B(creg[752]), .Z(n27207) );
  NAND U36703 ( .A(n27209), .B(n27210), .Z(c[751]) );
  NAND U36704 ( .A(n26658), .B(o[751]), .Z(n27210) );
  NAND U36705 ( .A(n26653), .B(creg[751]), .Z(n27209) );
  NAND U36706 ( .A(n27211), .B(n27212), .Z(c[750]) );
  NAND U36707 ( .A(n26658), .B(o[750]), .Z(n27212) );
  NAND U36708 ( .A(n26653), .B(creg[750]), .Z(n27211) );
  NAND U36709 ( .A(n27213), .B(n27214), .Z(c[74]) );
  NAND U36710 ( .A(n26658), .B(o[74]), .Z(n27214) );
  NAND U36711 ( .A(n26653), .B(creg[74]), .Z(n27213) );
  NAND U36712 ( .A(n27215), .B(n27216), .Z(c[749]) );
  NAND U36713 ( .A(n26658), .B(o[749]), .Z(n27216) );
  NAND U36714 ( .A(n26653), .B(creg[749]), .Z(n27215) );
  NAND U36715 ( .A(n27217), .B(n27218), .Z(c[748]) );
  NAND U36716 ( .A(n26658), .B(o[748]), .Z(n27218) );
  NAND U36717 ( .A(n26653), .B(creg[748]), .Z(n27217) );
  NAND U36718 ( .A(n27219), .B(n27220), .Z(c[747]) );
  NAND U36719 ( .A(n26658), .B(o[747]), .Z(n27220) );
  NAND U36720 ( .A(n26653), .B(creg[747]), .Z(n27219) );
  NAND U36721 ( .A(n27221), .B(n27222), .Z(c[746]) );
  NAND U36722 ( .A(n26658), .B(o[746]), .Z(n27222) );
  NAND U36723 ( .A(n26653), .B(creg[746]), .Z(n27221) );
  NAND U36724 ( .A(n27223), .B(n27224), .Z(c[745]) );
  NAND U36725 ( .A(n26658), .B(o[745]), .Z(n27224) );
  NAND U36726 ( .A(n26653), .B(creg[745]), .Z(n27223) );
  NAND U36727 ( .A(n27225), .B(n27226), .Z(c[744]) );
  NAND U36728 ( .A(n26658), .B(o[744]), .Z(n27226) );
  NAND U36729 ( .A(n26653), .B(creg[744]), .Z(n27225) );
  NAND U36730 ( .A(n27227), .B(n27228), .Z(c[743]) );
  NAND U36731 ( .A(n26658), .B(o[743]), .Z(n27228) );
  NAND U36732 ( .A(n26653), .B(creg[743]), .Z(n27227) );
  NAND U36733 ( .A(n27229), .B(n27230), .Z(c[742]) );
  NAND U36734 ( .A(n26658), .B(o[742]), .Z(n27230) );
  NAND U36735 ( .A(n26653), .B(creg[742]), .Z(n27229) );
  NAND U36736 ( .A(n27231), .B(n27232), .Z(c[741]) );
  NAND U36737 ( .A(n26658), .B(o[741]), .Z(n27232) );
  NAND U36738 ( .A(n26653), .B(creg[741]), .Z(n27231) );
  NAND U36739 ( .A(n27233), .B(n27234), .Z(c[740]) );
  NAND U36740 ( .A(n26658), .B(o[740]), .Z(n27234) );
  NAND U36741 ( .A(n26653), .B(creg[740]), .Z(n27233) );
  NAND U36742 ( .A(n27235), .B(n27236), .Z(c[73]) );
  NAND U36743 ( .A(n26658), .B(o[73]), .Z(n27236) );
  NAND U36744 ( .A(n26653), .B(creg[73]), .Z(n27235) );
  NAND U36745 ( .A(n27237), .B(n27238), .Z(c[739]) );
  NAND U36746 ( .A(n26658), .B(o[739]), .Z(n27238) );
  NAND U36747 ( .A(n26653), .B(creg[739]), .Z(n27237) );
  NAND U36748 ( .A(n27239), .B(n27240), .Z(c[738]) );
  NAND U36749 ( .A(n26658), .B(o[738]), .Z(n27240) );
  NAND U36750 ( .A(n26653), .B(creg[738]), .Z(n27239) );
  NAND U36751 ( .A(n27241), .B(n27242), .Z(c[737]) );
  NAND U36752 ( .A(n26658), .B(o[737]), .Z(n27242) );
  NAND U36753 ( .A(n26653), .B(creg[737]), .Z(n27241) );
  NAND U36754 ( .A(n27243), .B(n27244), .Z(c[736]) );
  NAND U36755 ( .A(n26658), .B(o[736]), .Z(n27244) );
  NAND U36756 ( .A(n26653), .B(creg[736]), .Z(n27243) );
  NAND U36757 ( .A(n27245), .B(n27246), .Z(c[735]) );
  NAND U36758 ( .A(n26658), .B(o[735]), .Z(n27246) );
  NAND U36759 ( .A(n26653), .B(creg[735]), .Z(n27245) );
  NAND U36760 ( .A(n27247), .B(n27248), .Z(c[734]) );
  NAND U36761 ( .A(n26658), .B(o[734]), .Z(n27248) );
  NAND U36762 ( .A(n26653), .B(creg[734]), .Z(n27247) );
  NAND U36763 ( .A(n27249), .B(n27250), .Z(c[733]) );
  NAND U36764 ( .A(n26658), .B(o[733]), .Z(n27250) );
  NAND U36765 ( .A(n26653), .B(creg[733]), .Z(n27249) );
  NAND U36766 ( .A(n27251), .B(n27252), .Z(c[732]) );
  NAND U36767 ( .A(n26658), .B(o[732]), .Z(n27252) );
  NAND U36768 ( .A(n26653), .B(creg[732]), .Z(n27251) );
  NAND U36769 ( .A(n27253), .B(n27254), .Z(c[731]) );
  NAND U36770 ( .A(n26658), .B(o[731]), .Z(n27254) );
  NAND U36771 ( .A(n26653), .B(creg[731]), .Z(n27253) );
  NAND U36772 ( .A(n27255), .B(n27256), .Z(c[730]) );
  NAND U36773 ( .A(n26658), .B(o[730]), .Z(n27256) );
  NAND U36774 ( .A(n26653), .B(creg[730]), .Z(n27255) );
  NAND U36775 ( .A(n27257), .B(n27258), .Z(c[72]) );
  NAND U36776 ( .A(n26658), .B(o[72]), .Z(n27258) );
  NAND U36777 ( .A(n26653), .B(creg[72]), .Z(n27257) );
  NAND U36778 ( .A(n27259), .B(n27260), .Z(c[729]) );
  NAND U36779 ( .A(n26658), .B(o[729]), .Z(n27260) );
  NAND U36780 ( .A(n26653), .B(creg[729]), .Z(n27259) );
  NAND U36781 ( .A(n27261), .B(n27262), .Z(c[728]) );
  NAND U36782 ( .A(n26658), .B(o[728]), .Z(n27262) );
  NAND U36783 ( .A(n26653), .B(creg[728]), .Z(n27261) );
  NAND U36784 ( .A(n27263), .B(n27264), .Z(c[727]) );
  NAND U36785 ( .A(n26658), .B(o[727]), .Z(n27264) );
  NAND U36786 ( .A(n26653), .B(creg[727]), .Z(n27263) );
  NAND U36787 ( .A(n27265), .B(n27266), .Z(c[726]) );
  NAND U36788 ( .A(n26658), .B(o[726]), .Z(n27266) );
  NAND U36789 ( .A(n26653), .B(creg[726]), .Z(n27265) );
  NAND U36790 ( .A(n27267), .B(n27268), .Z(c[725]) );
  NAND U36791 ( .A(n26658), .B(o[725]), .Z(n27268) );
  NAND U36792 ( .A(n26653), .B(creg[725]), .Z(n27267) );
  NAND U36793 ( .A(n27269), .B(n27270), .Z(c[724]) );
  NAND U36794 ( .A(n26658), .B(o[724]), .Z(n27270) );
  NAND U36795 ( .A(n26653), .B(creg[724]), .Z(n27269) );
  NAND U36796 ( .A(n27271), .B(n27272), .Z(c[723]) );
  NAND U36797 ( .A(n26658), .B(o[723]), .Z(n27272) );
  NAND U36798 ( .A(n26653), .B(creg[723]), .Z(n27271) );
  NAND U36799 ( .A(n27273), .B(n27274), .Z(c[722]) );
  NAND U36800 ( .A(n26658), .B(o[722]), .Z(n27274) );
  NAND U36801 ( .A(n26653), .B(creg[722]), .Z(n27273) );
  NAND U36802 ( .A(n27275), .B(n27276), .Z(c[721]) );
  NAND U36803 ( .A(n26658), .B(o[721]), .Z(n27276) );
  NAND U36804 ( .A(n26653), .B(creg[721]), .Z(n27275) );
  NAND U36805 ( .A(n27277), .B(n27278), .Z(c[720]) );
  NAND U36806 ( .A(n26658), .B(o[720]), .Z(n27278) );
  NAND U36807 ( .A(n26653), .B(creg[720]), .Z(n27277) );
  NAND U36808 ( .A(n27279), .B(n27280), .Z(c[71]) );
  NAND U36809 ( .A(n26658), .B(o[71]), .Z(n27280) );
  NAND U36810 ( .A(n26653), .B(creg[71]), .Z(n27279) );
  NAND U36811 ( .A(n27281), .B(n27282), .Z(c[719]) );
  NAND U36812 ( .A(n26658), .B(o[719]), .Z(n27282) );
  NAND U36813 ( .A(n26653), .B(creg[719]), .Z(n27281) );
  NAND U36814 ( .A(n27283), .B(n27284), .Z(c[718]) );
  NAND U36815 ( .A(n26658), .B(o[718]), .Z(n27284) );
  NAND U36816 ( .A(n26653), .B(creg[718]), .Z(n27283) );
  NAND U36817 ( .A(n27285), .B(n27286), .Z(c[717]) );
  NAND U36818 ( .A(n26658), .B(o[717]), .Z(n27286) );
  NAND U36819 ( .A(n26653), .B(creg[717]), .Z(n27285) );
  NAND U36820 ( .A(n27287), .B(n27288), .Z(c[716]) );
  NAND U36821 ( .A(n26658), .B(o[716]), .Z(n27288) );
  NAND U36822 ( .A(n26653), .B(creg[716]), .Z(n27287) );
  NAND U36823 ( .A(n27289), .B(n27290), .Z(c[715]) );
  NAND U36824 ( .A(n26658), .B(o[715]), .Z(n27290) );
  NAND U36825 ( .A(n26653), .B(creg[715]), .Z(n27289) );
  NAND U36826 ( .A(n27291), .B(n27292), .Z(c[714]) );
  NAND U36827 ( .A(n26658), .B(o[714]), .Z(n27292) );
  NAND U36828 ( .A(n26653), .B(creg[714]), .Z(n27291) );
  NAND U36829 ( .A(n27293), .B(n27294), .Z(c[713]) );
  NAND U36830 ( .A(n26658), .B(o[713]), .Z(n27294) );
  NAND U36831 ( .A(n26653), .B(creg[713]), .Z(n27293) );
  NAND U36832 ( .A(n27295), .B(n27296), .Z(c[712]) );
  NAND U36833 ( .A(n26658), .B(o[712]), .Z(n27296) );
  NAND U36834 ( .A(n26653), .B(creg[712]), .Z(n27295) );
  NAND U36835 ( .A(n27297), .B(n27298), .Z(c[711]) );
  NAND U36836 ( .A(n26658), .B(o[711]), .Z(n27298) );
  NAND U36837 ( .A(n26653), .B(creg[711]), .Z(n27297) );
  NAND U36838 ( .A(n27299), .B(n27300), .Z(c[710]) );
  NAND U36839 ( .A(n26658), .B(o[710]), .Z(n27300) );
  NAND U36840 ( .A(n26653), .B(creg[710]), .Z(n27299) );
  NAND U36841 ( .A(n27301), .B(n27302), .Z(c[70]) );
  NAND U36842 ( .A(n26658), .B(o[70]), .Z(n27302) );
  NAND U36843 ( .A(n26653), .B(creg[70]), .Z(n27301) );
  NAND U36844 ( .A(n27303), .B(n27304), .Z(c[709]) );
  NAND U36845 ( .A(n26658), .B(o[709]), .Z(n27304) );
  NAND U36846 ( .A(n26653), .B(creg[709]), .Z(n27303) );
  NAND U36847 ( .A(n27305), .B(n27306), .Z(c[708]) );
  NAND U36848 ( .A(n26658), .B(o[708]), .Z(n27306) );
  NAND U36849 ( .A(n26653), .B(creg[708]), .Z(n27305) );
  NAND U36850 ( .A(n27307), .B(n27308), .Z(c[707]) );
  NAND U36851 ( .A(n26658), .B(o[707]), .Z(n27308) );
  NAND U36852 ( .A(n26653), .B(creg[707]), .Z(n27307) );
  NAND U36853 ( .A(n27309), .B(n27310), .Z(c[706]) );
  NAND U36854 ( .A(n26658), .B(o[706]), .Z(n27310) );
  NAND U36855 ( .A(n26653), .B(creg[706]), .Z(n27309) );
  NAND U36856 ( .A(n27311), .B(n27312), .Z(c[705]) );
  NAND U36857 ( .A(n26658), .B(o[705]), .Z(n27312) );
  NAND U36858 ( .A(n26653), .B(creg[705]), .Z(n27311) );
  NAND U36859 ( .A(n27313), .B(n27314), .Z(c[704]) );
  NAND U36860 ( .A(n26658), .B(o[704]), .Z(n27314) );
  NAND U36861 ( .A(n26653), .B(creg[704]), .Z(n27313) );
  NAND U36862 ( .A(n27315), .B(n27316), .Z(c[703]) );
  NAND U36863 ( .A(n26658), .B(o[703]), .Z(n27316) );
  NAND U36864 ( .A(n26653), .B(creg[703]), .Z(n27315) );
  NAND U36865 ( .A(n27317), .B(n27318), .Z(c[702]) );
  NAND U36866 ( .A(n26658), .B(o[702]), .Z(n27318) );
  NAND U36867 ( .A(n26653), .B(creg[702]), .Z(n27317) );
  NAND U36868 ( .A(n27319), .B(n27320), .Z(c[701]) );
  NAND U36869 ( .A(n26658), .B(o[701]), .Z(n27320) );
  NAND U36870 ( .A(n26653), .B(creg[701]), .Z(n27319) );
  NAND U36871 ( .A(n27321), .B(n27322), .Z(c[700]) );
  NAND U36872 ( .A(n26658), .B(o[700]), .Z(n27322) );
  NAND U36873 ( .A(n26653), .B(creg[700]), .Z(n27321) );
  NAND U36874 ( .A(n27323), .B(n27324), .Z(c[6]) );
  NAND U36875 ( .A(n26658), .B(o[6]), .Z(n27324) );
  NAND U36876 ( .A(n26653), .B(creg[6]), .Z(n27323) );
  NAND U36877 ( .A(n27325), .B(n27326), .Z(c[69]) );
  NAND U36878 ( .A(n26658), .B(o[69]), .Z(n27326) );
  NAND U36879 ( .A(n26653), .B(creg[69]), .Z(n27325) );
  NAND U36880 ( .A(n27327), .B(n27328), .Z(c[699]) );
  NAND U36881 ( .A(n26658), .B(o[699]), .Z(n27328) );
  NAND U36882 ( .A(n26653), .B(creg[699]), .Z(n27327) );
  NAND U36883 ( .A(n27329), .B(n27330), .Z(c[698]) );
  NAND U36884 ( .A(n26658), .B(o[698]), .Z(n27330) );
  NAND U36885 ( .A(n26653), .B(creg[698]), .Z(n27329) );
  NAND U36886 ( .A(n27331), .B(n27332), .Z(c[697]) );
  NAND U36887 ( .A(n26658), .B(o[697]), .Z(n27332) );
  NAND U36888 ( .A(n26653), .B(creg[697]), .Z(n27331) );
  NAND U36889 ( .A(n27333), .B(n27334), .Z(c[696]) );
  NAND U36890 ( .A(n26658), .B(o[696]), .Z(n27334) );
  NAND U36891 ( .A(n26653), .B(creg[696]), .Z(n27333) );
  NAND U36892 ( .A(n27335), .B(n27336), .Z(c[695]) );
  NAND U36893 ( .A(n26658), .B(o[695]), .Z(n27336) );
  NAND U36894 ( .A(n26653), .B(creg[695]), .Z(n27335) );
  NAND U36895 ( .A(n27337), .B(n27338), .Z(c[694]) );
  NAND U36896 ( .A(n26658), .B(o[694]), .Z(n27338) );
  NAND U36897 ( .A(n26653), .B(creg[694]), .Z(n27337) );
  NAND U36898 ( .A(n27339), .B(n27340), .Z(c[693]) );
  NAND U36899 ( .A(n26658), .B(o[693]), .Z(n27340) );
  NAND U36900 ( .A(n26653), .B(creg[693]), .Z(n27339) );
  NAND U36901 ( .A(n27341), .B(n27342), .Z(c[692]) );
  NAND U36902 ( .A(n26658), .B(o[692]), .Z(n27342) );
  NAND U36903 ( .A(n26653), .B(creg[692]), .Z(n27341) );
  NAND U36904 ( .A(n27343), .B(n27344), .Z(c[691]) );
  NAND U36905 ( .A(n26658), .B(o[691]), .Z(n27344) );
  NAND U36906 ( .A(n26653), .B(creg[691]), .Z(n27343) );
  NAND U36907 ( .A(n27345), .B(n27346), .Z(c[690]) );
  NAND U36908 ( .A(n26658), .B(o[690]), .Z(n27346) );
  NAND U36909 ( .A(n26653), .B(creg[690]), .Z(n27345) );
  NAND U36910 ( .A(n27347), .B(n27348), .Z(c[68]) );
  NAND U36911 ( .A(n26658), .B(o[68]), .Z(n27348) );
  NAND U36912 ( .A(n26653), .B(creg[68]), .Z(n27347) );
  NAND U36913 ( .A(n27349), .B(n27350), .Z(c[689]) );
  NAND U36914 ( .A(n26658), .B(o[689]), .Z(n27350) );
  NAND U36915 ( .A(n26653), .B(creg[689]), .Z(n27349) );
  NAND U36916 ( .A(n27351), .B(n27352), .Z(c[688]) );
  NAND U36917 ( .A(n26658), .B(o[688]), .Z(n27352) );
  NAND U36918 ( .A(n26653), .B(creg[688]), .Z(n27351) );
  NAND U36919 ( .A(n27353), .B(n27354), .Z(c[687]) );
  NAND U36920 ( .A(n26658), .B(o[687]), .Z(n27354) );
  NAND U36921 ( .A(n26653), .B(creg[687]), .Z(n27353) );
  NAND U36922 ( .A(n27355), .B(n27356), .Z(c[686]) );
  NAND U36923 ( .A(n26658), .B(o[686]), .Z(n27356) );
  NAND U36924 ( .A(n26653), .B(creg[686]), .Z(n27355) );
  NAND U36925 ( .A(n27357), .B(n27358), .Z(c[685]) );
  NAND U36926 ( .A(n26658), .B(o[685]), .Z(n27358) );
  NAND U36927 ( .A(n26653), .B(creg[685]), .Z(n27357) );
  NAND U36928 ( .A(n27359), .B(n27360), .Z(c[684]) );
  NAND U36929 ( .A(n26658), .B(o[684]), .Z(n27360) );
  NAND U36930 ( .A(n26653), .B(creg[684]), .Z(n27359) );
  NAND U36931 ( .A(n27361), .B(n27362), .Z(c[683]) );
  NAND U36932 ( .A(n26658), .B(o[683]), .Z(n27362) );
  NAND U36933 ( .A(n26653), .B(creg[683]), .Z(n27361) );
  NAND U36934 ( .A(n27363), .B(n27364), .Z(c[682]) );
  NAND U36935 ( .A(n26658), .B(o[682]), .Z(n27364) );
  NAND U36936 ( .A(n26653), .B(creg[682]), .Z(n27363) );
  NAND U36937 ( .A(n27365), .B(n27366), .Z(c[681]) );
  NAND U36938 ( .A(n26658), .B(o[681]), .Z(n27366) );
  NAND U36939 ( .A(n26653), .B(creg[681]), .Z(n27365) );
  NAND U36940 ( .A(n27367), .B(n27368), .Z(c[680]) );
  NAND U36941 ( .A(n26658), .B(o[680]), .Z(n27368) );
  NAND U36942 ( .A(n26653), .B(creg[680]), .Z(n27367) );
  NAND U36943 ( .A(n27369), .B(n27370), .Z(c[67]) );
  NAND U36944 ( .A(n26658), .B(o[67]), .Z(n27370) );
  NAND U36945 ( .A(n26653), .B(creg[67]), .Z(n27369) );
  NAND U36946 ( .A(n27371), .B(n27372), .Z(c[679]) );
  NAND U36947 ( .A(n26658), .B(o[679]), .Z(n27372) );
  NAND U36948 ( .A(n26653), .B(creg[679]), .Z(n27371) );
  NAND U36949 ( .A(n27373), .B(n27374), .Z(c[678]) );
  NAND U36950 ( .A(n26658), .B(o[678]), .Z(n27374) );
  NAND U36951 ( .A(n26653), .B(creg[678]), .Z(n27373) );
  NAND U36952 ( .A(n27375), .B(n27376), .Z(c[677]) );
  NAND U36953 ( .A(n26658), .B(o[677]), .Z(n27376) );
  NAND U36954 ( .A(n26653), .B(creg[677]), .Z(n27375) );
  NAND U36955 ( .A(n27377), .B(n27378), .Z(c[676]) );
  NAND U36956 ( .A(n26658), .B(o[676]), .Z(n27378) );
  NAND U36957 ( .A(n26653), .B(creg[676]), .Z(n27377) );
  NAND U36958 ( .A(n27379), .B(n27380), .Z(c[675]) );
  NAND U36959 ( .A(n26658), .B(o[675]), .Z(n27380) );
  NAND U36960 ( .A(n26653), .B(creg[675]), .Z(n27379) );
  NAND U36961 ( .A(n27381), .B(n27382), .Z(c[674]) );
  NAND U36962 ( .A(n26658), .B(o[674]), .Z(n27382) );
  NAND U36963 ( .A(n26653), .B(creg[674]), .Z(n27381) );
  NAND U36964 ( .A(n27383), .B(n27384), .Z(c[673]) );
  NAND U36965 ( .A(n26658), .B(o[673]), .Z(n27384) );
  NAND U36966 ( .A(n26653), .B(creg[673]), .Z(n27383) );
  NAND U36967 ( .A(n27385), .B(n27386), .Z(c[672]) );
  NAND U36968 ( .A(n26658), .B(o[672]), .Z(n27386) );
  NAND U36969 ( .A(n26653), .B(creg[672]), .Z(n27385) );
  NAND U36970 ( .A(n27387), .B(n27388), .Z(c[671]) );
  NAND U36971 ( .A(n26658), .B(o[671]), .Z(n27388) );
  NAND U36972 ( .A(n26653), .B(creg[671]), .Z(n27387) );
  NAND U36973 ( .A(n27389), .B(n27390), .Z(c[670]) );
  NAND U36974 ( .A(n26658), .B(o[670]), .Z(n27390) );
  NAND U36975 ( .A(n26653), .B(creg[670]), .Z(n27389) );
  NAND U36976 ( .A(n27391), .B(n27392), .Z(c[66]) );
  NAND U36977 ( .A(n26658), .B(o[66]), .Z(n27392) );
  NAND U36978 ( .A(n26653), .B(creg[66]), .Z(n27391) );
  NAND U36979 ( .A(n27393), .B(n27394), .Z(c[669]) );
  NAND U36980 ( .A(n26658), .B(o[669]), .Z(n27394) );
  NAND U36981 ( .A(n26653), .B(creg[669]), .Z(n27393) );
  NAND U36982 ( .A(n27395), .B(n27396), .Z(c[668]) );
  NAND U36983 ( .A(n26658), .B(o[668]), .Z(n27396) );
  NAND U36984 ( .A(n26653), .B(creg[668]), .Z(n27395) );
  NAND U36985 ( .A(n27397), .B(n27398), .Z(c[667]) );
  NAND U36986 ( .A(n26658), .B(o[667]), .Z(n27398) );
  NAND U36987 ( .A(n26653), .B(creg[667]), .Z(n27397) );
  NAND U36988 ( .A(n27399), .B(n27400), .Z(c[666]) );
  NAND U36989 ( .A(n26658), .B(o[666]), .Z(n27400) );
  NAND U36990 ( .A(n26653), .B(creg[666]), .Z(n27399) );
  NAND U36991 ( .A(n27401), .B(n27402), .Z(c[665]) );
  NAND U36992 ( .A(n26658), .B(o[665]), .Z(n27402) );
  NAND U36993 ( .A(n26653), .B(creg[665]), .Z(n27401) );
  NAND U36994 ( .A(n27403), .B(n27404), .Z(c[664]) );
  NAND U36995 ( .A(n26658), .B(o[664]), .Z(n27404) );
  NAND U36996 ( .A(n26653), .B(creg[664]), .Z(n27403) );
  NAND U36997 ( .A(n27405), .B(n27406), .Z(c[663]) );
  NAND U36998 ( .A(n26658), .B(o[663]), .Z(n27406) );
  NAND U36999 ( .A(n26653), .B(creg[663]), .Z(n27405) );
  NAND U37000 ( .A(n27407), .B(n27408), .Z(c[662]) );
  NAND U37001 ( .A(n26658), .B(o[662]), .Z(n27408) );
  NAND U37002 ( .A(n26653), .B(creg[662]), .Z(n27407) );
  NAND U37003 ( .A(n27409), .B(n27410), .Z(c[661]) );
  NAND U37004 ( .A(n26658), .B(o[661]), .Z(n27410) );
  NAND U37005 ( .A(n26653), .B(creg[661]), .Z(n27409) );
  NAND U37006 ( .A(n27411), .B(n27412), .Z(c[660]) );
  NAND U37007 ( .A(n26658), .B(o[660]), .Z(n27412) );
  NAND U37008 ( .A(n26653), .B(creg[660]), .Z(n27411) );
  NAND U37009 ( .A(n27413), .B(n27414), .Z(c[65]) );
  NAND U37010 ( .A(n26658), .B(o[65]), .Z(n27414) );
  NAND U37011 ( .A(n26653), .B(creg[65]), .Z(n27413) );
  NAND U37012 ( .A(n27415), .B(n27416), .Z(c[659]) );
  NAND U37013 ( .A(n26658), .B(o[659]), .Z(n27416) );
  NAND U37014 ( .A(n26653), .B(creg[659]), .Z(n27415) );
  NAND U37015 ( .A(n27417), .B(n27418), .Z(c[658]) );
  NAND U37016 ( .A(n26658), .B(o[658]), .Z(n27418) );
  NAND U37017 ( .A(n26653), .B(creg[658]), .Z(n27417) );
  NAND U37018 ( .A(n27419), .B(n27420), .Z(c[657]) );
  NAND U37019 ( .A(n26658), .B(o[657]), .Z(n27420) );
  NAND U37020 ( .A(n26653), .B(creg[657]), .Z(n27419) );
  NAND U37021 ( .A(n27421), .B(n27422), .Z(c[656]) );
  NAND U37022 ( .A(n26658), .B(o[656]), .Z(n27422) );
  NAND U37023 ( .A(n26653), .B(creg[656]), .Z(n27421) );
  NAND U37024 ( .A(n27423), .B(n27424), .Z(c[655]) );
  NAND U37025 ( .A(n26658), .B(o[655]), .Z(n27424) );
  NAND U37026 ( .A(n26653), .B(creg[655]), .Z(n27423) );
  NAND U37027 ( .A(n27425), .B(n27426), .Z(c[654]) );
  NAND U37028 ( .A(n26658), .B(o[654]), .Z(n27426) );
  NAND U37029 ( .A(n26653), .B(creg[654]), .Z(n27425) );
  NAND U37030 ( .A(n27427), .B(n27428), .Z(c[653]) );
  NAND U37031 ( .A(n26658), .B(o[653]), .Z(n27428) );
  NAND U37032 ( .A(n26653), .B(creg[653]), .Z(n27427) );
  NAND U37033 ( .A(n27429), .B(n27430), .Z(c[652]) );
  NAND U37034 ( .A(n26658), .B(o[652]), .Z(n27430) );
  NAND U37035 ( .A(n26653), .B(creg[652]), .Z(n27429) );
  NAND U37036 ( .A(n27431), .B(n27432), .Z(c[651]) );
  NAND U37037 ( .A(n26658), .B(o[651]), .Z(n27432) );
  NAND U37038 ( .A(n26653), .B(creg[651]), .Z(n27431) );
  NAND U37039 ( .A(n27433), .B(n27434), .Z(c[650]) );
  NAND U37040 ( .A(n26658), .B(o[650]), .Z(n27434) );
  NAND U37041 ( .A(n26653), .B(creg[650]), .Z(n27433) );
  NAND U37042 ( .A(n27435), .B(n27436), .Z(c[64]) );
  NAND U37043 ( .A(n26658), .B(o[64]), .Z(n27436) );
  NAND U37044 ( .A(n26653), .B(creg[64]), .Z(n27435) );
  NAND U37045 ( .A(n27437), .B(n27438), .Z(c[649]) );
  NAND U37046 ( .A(n26658), .B(o[649]), .Z(n27438) );
  NAND U37047 ( .A(n26653), .B(creg[649]), .Z(n27437) );
  NAND U37048 ( .A(n27439), .B(n27440), .Z(c[648]) );
  NAND U37049 ( .A(n26658), .B(o[648]), .Z(n27440) );
  NAND U37050 ( .A(n26653), .B(creg[648]), .Z(n27439) );
  NAND U37051 ( .A(n27441), .B(n27442), .Z(c[647]) );
  NAND U37052 ( .A(n26658), .B(o[647]), .Z(n27442) );
  NAND U37053 ( .A(n26653), .B(creg[647]), .Z(n27441) );
  NAND U37054 ( .A(n27443), .B(n27444), .Z(c[646]) );
  NAND U37055 ( .A(n26658), .B(o[646]), .Z(n27444) );
  NAND U37056 ( .A(n26653), .B(creg[646]), .Z(n27443) );
  NAND U37057 ( .A(n27445), .B(n27446), .Z(c[645]) );
  NAND U37058 ( .A(n26658), .B(o[645]), .Z(n27446) );
  NAND U37059 ( .A(n26653), .B(creg[645]), .Z(n27445) );
  NAND U37060 ( .A(n27447), .B(n27448), .Z(c[644]) );
  NAND U37061 ( .A(n26658), .B(o[644]), .Z(n27448) );
  NAND U37062 ( .A(n26653), .B(creg[644]), .Z(n27447) );
  NAND U37063 ( .A(n27449), .B(n27450), .Z(c[643]) );
  NAND U37064 ( .A(n26658), .B(o[643]), .Z(n27450) );
  NAND U37065 ( .A(n26653), .B(creg[643]), .Z(n27449) );
  NAND U37066 ( .A(n27451), .B(n27452), .Z(c[642]) );
  NAND U37067 ( .A(n26658), .B(o[642]), .Z(n27452) );
  NAND U37068 ( .A(n26653), .B(creg[642]), .Z(n27451) );
  NAND U37069 ( .A(n27453), .B(n27454), .Z(c[641]) );
  NAND U37070 ( .A(n26658), .B(o[641]), .Z(n27454) );
  NAND U37071 ( .A(n26653), .B(creg[641]), .Z(n27453) );
  NAND U37072 ( .A(n27455), .B(n27456), .Z(c[640]) );
  NAND U37073 ( .A(n26658), .B(o[640]), .Z(n27456) );
  NAND U37074 ( .A(n26653), .B(creg[640]), .Z(n27455) );
  NAND U37075 ( .A(n27457), .B(n27458), .Z(c[63]) );
  NAND U37076 ( .A(n26658), .B(o[63]), .Z(n27458) );
  NAND U37077 ( .A(n26653), .B(creg[63]), .Z(n27457) );
  NAND U37078 ( .A(n27459), .B(n27460), .Z(c[639]) );
  NAND U37079 ( .A(n26658), .B(o[639]), .Z(n27460) );
  NAND U37080 ( .A(n26653), .B(creg[639]), .Z(n27459) );
  NAND U37081 ( .A(n27461), .B(n27462), .Z(c[638]) );
  NAND U37082 ( .A(n26658), .B(o[638]), .Z(n27462) );
  NAND U37083 ( .A(n26653), .B(creg[638]), .Z(n27461) );
  NAND U37084 ( .A(n27463), .B(n27464), .Z(c[637]) );
  NAND U37085 ( .A(n26658), .B(o[637]), .Z(n27464) );
  NAND U37086 ( .A(n26653), .B(creg[637]), .Z(n27463) );
  NAND U37087 ( .A(n27465), .B(n27466), .Z(c[636]) );
  NAND U37088 ( .A(n26658), .B(o[636]), .Z(n27466) );
  NAND U37089 ( .A(n26653), .B(creg[636]), .Z(n27465) );
  NAND U37090 ( .A(n27467), .B(n27468), .Z(c[635]) );
  NAND U37091 ( .A(n26658), .B(o[635]), .Z(n27468) );
  NAND U37092 ( .A(n26653), .B(creg[635]), .Z(n27467) );
  NAND U37093 ( .A(n27469), .B(n27470), .Z(c[634]) );
  NAND U37094 ( .A(n26658), .B(o[634]), .Z(n27470) );
  NAND U37095 ( .A(n26653), .B(creg[634]), .Z(n27469) );
  NAND U37096 ( .A(n27471), .B(n27472), .Z(c[633]) );
  NAND U37097 ( .A(n26658), .B(o[633]), .Z(n27472) );
  NAND U37098 ( .A(n26653), .B(creg[633]), .Z(n27471) );
  NAND U37099 ( .A(n27473), .B(n27474), .Z(c[632]) );
  NAND U37100 ( .A(n26658), .B(o[632]), .Z(n27474) );
  NAND U37101 ( .A(n26653), .B(creg[632]), .Z(n27473) );
  NAND U37102 ( .A(n27475), .B(n27476), .Z(c[631]) );
  NAND U37103 ( .A(n26658), .B(o[631]), .Z(n27476) );
  NAND U37104 ( .A(n26653), .B(creg[631]), .Z(n27475) );
  NAND U37105 ( .A(n27477), .B(n27478), .Z(c[630]) );
  NAND U37106 ( .A(n26658), .B(o[630]), .Z(n27478) );
  NAND U37107 ( .A(n26653), .B(creg[630]), .Z(n27477) );
  NAND U37108 ( .A(n27479), .B(n27480), .Z(c[62]) );
  NAND U37109 ( .A(n26658), .B(o[62]), .Z(n27480) );
  NAND U37110 ( .A(n26653), .B(creg[62]), .Z(n27479) );
  NAND U37111 ( .A(n27481), .B(n27482), .Z(c[629]) );
  NAND U37112 ( .A(n26658), .B(o[629]), .Z(n27482) );
  NAND U37113 ( .A(n26653), .B(creg[629]), .Z(n27481) );
  NAND U37114 ( .A(n27483), .B(n27484), .Z(c[628]) );
  NAND U37115 ( .A(n26658), .B(o[628]), .Z(n27484) );
  NAND U37116 ( .A(n26653), .B(creg[628]), .Z(n27483) );
  NAND U37117 ( .A(n27485), .B(n27486), .Z(c[627]) );
  NAND U37118 ( .A(n26658), .B(o[627]), .Z(n27486) );
  NAND U37119 ( .A(n26653), .B(creg[627]), .Z(n27485) );
  NAND U37120 ( .A(n27487), .B(n27488), .Z(c[626]) );
  NAND U37121 ( .A(n26658), .B(o[626]), .Z(n27488) );
  NAND U37122 ( .A(n26653), .B(creg[626]), .Z(n27487) );
  NAND U37123 ( .A(n27489), .B(n27490), .Z(c[625]) );
  NAND U37124 ( .A(n26658), .B(o[625]), .Z(n27490) );
  NAND U37125 ( .A(n26653), .B(creg[625]), .Z(n27489) );
  NAND U37126 ( .A(n27491), .B(n27492), .Z(c[624]) );
  NAND U37127 ( .A(n26658), .B(o[624]), .Z(n27492) );
  NAND U37128 ( .A(n26653), .B(creg[624]), .Z(n27491) );
  NAND U37129 ( .A(n27493), .B(n27494), .Z(c[623]) );
  NAND U37130 ( .A(n26658), .B(o[623]), .Z(n27494) );
  NAND U37131 ( .A(n26653), .B(creg[623]), .Z(n27493) );
  NAND U37132 ( .A(n27495), .B(n27496), .Z(c[622]) );
  NAND U37133 ( .A(n26658), .B(o[622]), .Z(n27496) );
  NAND U37134 ( .A(n26653), .B(creg[622]), .Z(n27495) );
  NAND U37135 ( .A(n27497), .B(n27498), .Z(c[621]) );
  NAND U37136 ( .A(n26658), .B(o[621]), .Z(n27498) );
  NAND U37137 ( .A(n26653), .B(creg[621]), .Z(n27497) );
  NAND U37138 ( .A(n27499), .B(n27500), .Z(c[620]) );
  NAND U37139 ( .A(n26658), .B(o[620]), .Z(n27500) );
  NAND U37140 ( .A(n26653), .B(creg[620]), .Z(n27499) );
  NAND U37141 ( .A(n27501), .B(n27502), .Z(c[61]) );
  NAND U37142 ( .A(n26658), .B(o[61]), .Z(n27502) );
  NAND U37143 ( .A(n26653), .B(creg[61]), .Z(n27501) );
  NAND U37144 ( .A(n27503), .B(n27504), .Z(c[619]) );
  NAND U37145 ( .A(n26658), .B(o[619]), .Z(n27504) );
  NAND U37146 ( .A(n26653), .B(creg[619]), .Z(n27503) );
  NAND U37147 ( .A(n27505), .B(n27506), .Z(c[618]) );
  NAND U37148 ( .A(n26658), .B(o[618]), .Z(n27506) );
  NAND U37149 ( .A(n26653), .B(creg[618]), .Z(n27505) );
  NAND U37150 ( .A(n27507), .B(n27508), .Z(c[617]) );
  NAND U37151 ( .A(n26658), .B(o[617]), .Z(n27508) );
  NAND U37152 ( .A(n26653), .B(creg[617]), .Z(n27507) );
  NAND U37153 ( .A(n27509), .B(n27510), .Z(c[616]) );
  NAND U37154 ( .A(n26658), .B(o[616]), .Z(n27510) );
  NAND U37155 ( .A(n26653), .B(creg[616]), .Z(n27509) );
  NAND U37156 ( .A(n27511), .B(n27512), .Z(c[615]) );
  NAND U37157 ( .A(n26658), .B(o[615]), .Z(n27512) );
  NAND U37158 ( .A(n26653), .B(creg[615]), .Z(n27511) );
  NAND U37159 ( .A(n27513), .B(n27514), .Z(c[614]) );
  NAND U37160 ( .A(n26658), .B(o[614]), .Z(n27514) );
  NAND U37161 ( .A(n26653), .B(creg[614]), .Z(n27513) );
  NAND U37162 ( .A(n27515), .B(n27516), .Z(c[613]) );
  NAND U37163 ( .A(n26658), .B(o[613]), .Z(n27516) );
  NAND U37164 ( .A(n26653), .B(creg[613]), .Z(n27515) );
  NAND U37165 ( .A(n27517), .B(n27518), .Z(c[612]) );
  NAND U37166 ( .A(n26658), .B(o[612]), .Z(n27518) );
  NAND U37167 ( .A(n26653), .B(creg[612]), .Z(n27517) );
  NAND U37168 ( .A(n27519), .B(n27520), .Z(c[611]) );
  NAND U37169 ( .A(n26658), .B(o[611]), .Z(n27520) );
  NAND U37170 ( .A(n26653), .B(creg[611]), .Z(n27519) );
  NAND U37171 ( .A(n27521), .B(n27522), .Z(c[610]) );
  NAND U37172 ( .A(n26658), .B(o[610]), .Z(n27522) );
  NAND U37173 ( .A(n26653), .B(creg[610]), .Z(n27521) );
  NAND U37174 ( .A(n27523), .B(n27524), .Z(c[60]) );
  NAND U37175 ( .A(n26658), .B(o[60]), .Z(n27524) );
  NAND U37176 ( .A(n26653), .B(creg[60]), .Z(n27523) );
  NAND U37177 ( .A(n27525), .B(n27526), .Z(c[609]) );
  NAND U37178 ( .A(n26658), .B(o[609]), .Z(n27526) );
  NAND U37179 ( .A(n26653), .B(creg[609]), .Z(n27525) );
  NAND U37180 ( .A(n27527), .B(n27528), .Z(c[608]) );
  NAND U37181 ( .A(n26658), .B(o[608]), .Z(n27528) );
  NAND U37182 ( .A(n26653), .B(creg[608]), .Z(n27527) );
  NAND U37183 ( .A(n27529), .B(n27530), .Z(c[607]) );
  NAND U37184 ( .A(n26658), .B(o[607]), .Z(n27530) );
  NAND U37185 ( .A(n26653), .B(creg[607]), .Z(n27529) );
  NAND U37186 ( .A(n27531), .B(n27532), .Z(c[606]) );
  NAND U37187 ( .A(n26658), .B(o[606]), .Z(n27532) );
  NAND U37188 ( .A(n26653), .B(creg[606]), .Z(n27531) );
  NAND U37189 ( .A(n27533), .B(n27534), .Z(c[605]) );
  NAND U37190 ( .A(n26658), .B(o[605]), .Z(n27534) );
  NAND U37191 ( .A(n26653), .B(creg[605]), .Z(n27533) );
  NAND U37192 ( .A(n27535), .B(n27536), .Z(c[604]) );
  NAND U37193 ( .A(n26658), .B(o[604]), .Z(n27536) );
  NAND U37194 ( .A(n26653), .B(creg[604]), .Z(n27535) );
  NAND U37195 ( .A(n27537), .B(n27538), .Z(c[603]) );
  NAND U37196 ( .A(n26658), .B(o[603]), .Z(n27538) );
  NAND U37197 ( .A(n26653), .B(creg[603]), .Z(n27537) );
  NAND U37198 ( .A(n27539), .B(n27540), .Z(c[602]) );
  NAND U37199 ( .A(n26658), .B(o[602]), .Z(n27540) );
  NAND U37200 ( .A(n26653), .B(creg[602]), .Z(n27539) );
  NAND U37201 ( .A(n27541), .B(n27542), .Z(c[601]) );
  NAND U37202 ( .A(n26658), .B(o[601]), .Z(n27542) );
  NAND U37203 ( .A(n26653), .B(creg[601]), .Z(n27541) );
  NAND U37204 ( .A(n27543), .B(n27544), .Z(c[600]) );
  NAND U37205 ( .A(n26658), .B(o[600]), .Z(n27544) );
  NAND U37206 ( .A(n26653), .B(creg[600]), .Z(n27543) );
  NAND U37207 ( .A(n27545), .B(n27546), .Z(c[5]) );
  NAND U37208 ( .A(n26658), .B(o[5]), .Z(n27546) );
  NAND U37209 ( .A(n26653), .B(creg[5]), .Z(n27545) );
  NAND U37210 ( .A(n27547), .B(n27548), .Z(c[59]) );
  NAND U37211 ( .A(n26658), .B(o[59]), .Z(n27548) );
  NAND U37212 ( .A(n26653), .B(creg[59]), .Z(n27547) );
  NAND U37213 ( .A(n27549), .B(n27550), .Z(c[599]) );
  NAND U37214 ( .A(n26658), .B(o[599]), .Z(n27550) );
  NAND U37215 ( .A(n26653), .B(creg[599]), .Z(n27549) );
  NAND U37216 ( .A(n27551), .B(n27552), .Z(c[598]) );
  NAND U37217 ( .A(n26658), .B(o[598]), .Z(n27552) );
  NAND U37218 ( .A(n26653), .B(creg[598]), .Z(n27551) );
  NAND U37219 ( .A(n27553), .B(n27554), .Z(c[597]) );
  NAND U37220 ( .A(n26658), .B(o[597]), .Z(n27554) );
  NAND U37221 ( .A(n26653), .B(creg[597]), .Z(n27553) );
  NAND U37222 ( .A(n27555), .B(n27556), .Z(c[596]) );
  NAND U37223 ( .A(n26658), .B(o[596]), .Z(n27556) );
  NAND U37224 ( .A(n26653), .B(creg[596]), .Z(n27555) );
  NAND U37225 ( .A(n27557), .B(n27558), .Z(c[595]) );
  NAND U37226 ( .A(n26658), .B(o[595]), .Z(n27558) );
  NAND U37227 ( .A(n26653), .B(creg[595]), .Z(n27557) );
  NAND U37228 ( .A(n27559), .B(n27560), .Z(c[594]) );
  NAND U37229 ( .A(n26658), .B(o[594]), .Z(n27560) );
  NAND U37230 ( .A(n26653), .B(creg[594]), .Z(n27559) );
  NAND U37231 ( .A(n27561), .B(n27562), .Z(c[593]) );
  NAND U37232 ( .A(n26658), .B(o[593]), .Z(n27562) );
  NAND U37233 ( .A(n26653), .B(creg[593]), .Z(n27561) );
  NAND U37234 ( .A(n27563), .B(n27564), .Z(c[592]) );
  NAND U37235 ( .A(n26658), .B(o[592]), .Z(n27564) );
  NAND U37236 ( .A(n26653), .B(creg[592]), .Z(n27563) );
  NAND U37237 ( .A(n27565), .B(n27566), .Z(c[591]) );
  NAND U37238 ( .A(n26658), .B(o[591]), .Z(n27566) );
  NAND U37239 ( .A(n26653), .B(creg[591]), .Z(n27565) );
  NAND U37240 ( .A(n27567), .B(n27568), .Z(c[590]) );
  NAND U37241 ( .A(n26658), .B(o[590]), .Z(n27568) );
  NAND U37242 ( .A(n26653), .B(creg[590]), .Z(n27567) );
  NAND U37243 ( .A(n27569), .B(n27570), .Z(c[58]) );
  NAND U37244 ( .A(n26658), .B(o[58]), .Z(n27570) );
  NAND U37245 ( .A(n26653), .B(creg[58]), .Z(n27569) );
  NAND U37246 ( .A(n27571), .B(n27572), .Z(c[589]) );
  NAND U37247 ( .A(n26658), .B(o[589]), .Z(n27572) );
  NAND U37248 ( .A(n26653), .B(creg[589]), .Z(n27571) );
  NAND U37249 ( .A(n27573), .B(n27574), .Z(c[588]) );
  NAND U37250 ( .A(n26658), .B(o[588]), .Z(n27574) );
  NAND U37251 ( .A(n26653), .B(creg[588]), .Z(n27573) );
  NAND U37252 ( .A(n27575), .B(n27576), .Z(c[587]) );
  NAND U37253 ( .A(n26658), .B(o[587]), .Z(n27576) );
  NAND U37254 ( .A(n26653), .B(creg[587]), .Z(n27575) );
  NAND U37255 ( .A(n27577), .B(n27578), .Z(c[586]) );
  NAND U37256 ( .A(n26658), .B(o[586]), .Z(n27578) );
  NAND U37257 ( .A(n26653), .B(creg[586]), .Z(n27577) );
  NAND U37258 ( .A(n27579), .B(n27580), .Z(c[585]) );
  NAND U37259 ( .A(n26658), .B(o[585]), .Z(n27580) );
  NAND U37260 ( .A(n26653), .B(creg[585]), .Z(n27579) );
  NAND U37261 ( .A(n27581), .B(n27582), .Z(c[584]) );
  NAND U37262 ( .A(n26658), .B(o[584]), .Z(n27582) );
  NAND U37263 ( .A(n26653), .B(creg[584]), .Z(n27581) );
  NAND U37264 ( .A(n27583), .B(n27584), .Z(c[583]) );
  NAND U37265 ( .A(n26658), .B(o[583]), .Z(n27584) );
  NAND U37266 ( .A(n26653), .B(creg[583]), .Z(n27583) );
  NAND U37267 ( .A(n27585), .B(n27586), .Z(c[582]) );
  NAND U37268 ( .A(n26658), .B(o[582]), .Z(n27586) );
  NAND U37269 ( .A(n26653), .B(creg[582]), .Z(n27585) );
  NAND U37270 ( .A(n27587), .B(n27588), .Z(c[581]) );
  NAND U37271 ( .A(n26658), .B(o[581]), .Z(n27588) );
  NAND U37272 ( .A(n26653), .B(creg[581]), .Z(n27587) );
  NAND U37273 ( .A(n27589), .B(n27590), .Z(c[580]) );
  NAND U37274 ( .A(n26658), .B(o[580]), .Z(n27590) );
  NAND U37275 ( .A(n26653), .B(creg[580]), .Z(n27589) );
  NAND U37276 ( .A(n27591), .B(n27592), .Z(c[57]) );
  NAND U37277 ( .A(n26658), .B(o[57]), .Z(n27592) );
  NAND U37278 ( .A(n26653), .B(creg[57]), .Z(n27591) );
  NAND U37279 ( .A(n27593), .B(n27594), .Z(c[579]) );
  NAND U37280 ( .A(n26658), .B(o[579]), .Z(n27594) );
  NAND U37281 ( .A(n26653), .B(creg[579]), .Z(n27593) );
  NAND U37282 ( .A(n27595), .B(n27596), .Z(c[578]) );
  NAND U37283 ( .A(n26658), .B(o[578]), .Z(n27596) );
  NAND U37284 ( .A(n26653), .B(creg[578]), .Z(n27595) );
  NAND U37285 ( .A(n27597), .B(n27598), .Z(c[577]) );
  NAND U37286 ( .A(n26658), .B(o[577]), .Z(n27598) );
  NAND U37287 ( .A(n26653), .B(creg[577]), .Z(n27597) );
  NAND U37288 ( .A(n27599), .B(n27600), .Z(c[576]) );
  NAND U37289 ( .A(n26658), .B(o[576]), .Z(n27600) );
  NAND U37290 ( .A(n26653), .B(creg[576]), .Z(n27599) );
  NAND U37291 ( .A(n27601), .B(n27602), .Z(c[575]) );
  NAND U37292 ( .A(n26658), .B(o[575]), .Z(n27602) );
  NAND U37293 ( .A(n26653), .B(creg[575]), .Z(n27601) );
  NAND U37294 ( .A(n27603), .B(n27604), .Z(c[574]) );
  NAND U37295 ( .A(n26658), .B(o[574]), .Z(n27604) );
  NAND U37296 ( .A(n26653), .B(creg[574]), .Z(n27603) );
  NAND U37297 ( .A(n27605), .B(n27606), .Z(c[573]) );
  NAND U37298 ( .A(n26658), .B(o[573]), .Z(n27606) );
  NAND U37299 ( .A(n26653), .B(creg[573]), .Z(n27605) );
  NAND U37300 ( .A(n27607), .B(n27608), .Z(c[572]) );
  NAND U37301 ( .A(n26658), .B(o[572]), .Z(n27608) );
  NAND U37302 ( .A(n26653), .B(creg[572]), .Z(n27607) );
  NAND U37303 ( .A(n27609), .B(n27610), .Z(c[571]) );
  NAND U37304 ( .A(n26658), .B(o[571]), .Z(n27610) );
  NAND U37305 ( .A(n26653), .B(creg[571]), .Z(n27609) );
  NAND U37306 ( .A(n27611), .B(n27612), .Z(c[570]) );
  NAND U37307 ( .A(n26658), .B(o[570]), .Z(n27612) );
  NAND U37308 ( .A(n26653), .B(creg[570]), .Z(n27611) );
  NAND U37309 ( .A(n27613), .B(n27614), .Z(c[56]) );
  NAND U37310 ( .A(n26658), .B(o[56]), .Z(n27614) );
  NAND U37311 ( .A(n26653), .B(creg[56]), .Z(n27613) );
  NAND U37312 ( .A(n27615), .B(n27616), .Z(c[569]) );
  NAND U37313 ( .A(n26658), .B(o[569]), .Z(n27616) );
  NAND U37314 ( .A(n26653), .B(creg[569]), .Z(n27615) );
  NAND U37315 ( .A(n27617), .B(n27618), .Z(c[568]) );
  NAND U37316 ( .A(n26658), .B(o[568]), .Z(n27618) );
  NAND U37317 ( .A(n26653), .B(creg[568]), .Z(n27617) );
  NAND U37318 ( .A(n27619), .B(n27620), .Z(c[567]) );
  NAND U37319 ( .A(n26658), .B(o[567]), .Z(n27620) );
  NAND U37320 ( .A(n26653), .B(creg[567]), .Z(n27619) );
  NAND U37321 ( .A(n27621), .B(n27622), .Z(c[566]) );
  NAND U37322 ( .A(n26658), .B(o[566]), .Z(n27622) );
  NAND U37323 ( .A(n26653), .B(creg[566]), .Z(n27621) );
  NAND U37324 ( .A(n27623), .B(n27624), .Z(c[565]) );
  NAND U37325 ( .A(n26658), .B(o[565]), .Z(n27624) );
  NAND U37326 ( .A(n26653), .B(creg[565]), .Z(n27623) );
  NAND U37327 ( .A(n27625), .B(n27626), .Z(c[564]) );
  NAND U37328 ( .A(n26658), .B(o[564]), .Z(n27626) );
  NAND U37329 ( .A(n26653), .B(creg[564]), .Z(n27625) );
  NAND U37330 ( .A(n27627), .B(n27628), .Z(c[563]) );
  NAND U37331 ( .A(n26658), .B(o[563]), .Z(n27628) );
  NAND U37332 ( .A(n26653), .B(creg[563]), .Z(n27627) );
  NAND U37333 ( .A(n27629), .B(n27630), .Z(c[562]) );
  NAND U37334 ( .A(n26658), .B(o[562]), .Z(n27630) );
  NAND U37335 ( .A(n26653), .B(creg[562]), .Z(n27629) );
  NAND U37336 ( .A(n27631), .B(n27632), .Z(c[561]) );
  NAND U37337 ( .A(n26658), .B(o[561]), .Z(n27632) );
  NAND U37338 ( .A(n26653), .B(creg[561]), .Z(n27631) );
  NAND U37339 ( .A(n27633), .B(n27634), .Z(c[560]) );
  NAND U37340 ( .A(n26658), .B(o[560]), .Z(n27634) );
  NAND U37341 ( .A(n26653), .B(creg[560]), .Z(n27633) );
  NAND U37342 ( .A(n27635), .B(n27636), .Z(c[55]) );
  NAND U37343 ( .A(n26658), .B(o[55]), .Z(n27636) );
  NAND U37344 ( .A(n26653), .B(creg[55]), .Z(n27635) );
  NAND U37345 ( .A(n27637), .B(n27638), .Z(c[559]) );
  NAND U37346 ( .A(n26658), .B(o[559]), .Z(n27638) );
  NAND U37347 ( .A(n26653), .B(creg[559]), .Z(n27637) );
  NAND U37348 ( .A(n27639), .B(n27640), .Z(c[558]) );
  NAND U37349 ( .A(n26658), .B(o[558]), .Z(n27640) );
  NAND U37350 ( .A(n26653), .B(creg[558]), .Z(n27639) );
  NAND U37351 ( .A(n27641), .B(n27642), .Z(c[557]) );
  NAND U37352 ( .A(n26658), .B(o[557]), .Z(n27642) );
  NAND U37353 ( .A(n26653), .B(creg[557]), .Z(n27641) );
  NAND U37354 ( .A(n27643), .B(n27644), .Z(c[556]) );
  NAND U37355 ( .A(n26658), .B(o[556]), .Z(n27644) );
  NAND U37356 ( .A(n26653), .B(creg[556]), .Z(n27643) );
  NAND U37357 ( .A(n27645), .B(n27646), .Z(c[555]) );
  NAND U37358 ( .A(n26658), .B(o[555]), .Z(n27646) );
  NAND U37359 ( .A(n26653), .B(creg[555]), .Z(n27645) );
  NAND U37360 ( .A(n27647), .B(n27648), .Z(c[554]) );
  NAND U37361 ( .A(n26658), .B(o[554]), .Z(n27648) );
  NAND U37362 ( .A(n26653), .B(creg[554]), .Z(n27647) );
  NAND U37363 ( .A(n27649), .B(n27650), .Z(c[553]) );
  NAND U37364 ( .A(n26658), .B(o[553]), .Z(n27650) );
  NAND U37365 ( .A(n26653), .B(creg[553]), .Z(n27649) );
  NAND U37366 ( .A(n27651), .B(n27652), .Z(c[552]) );
  NAND U37367 ( .A(n26658), .B(o[552]), .Z(n27652) );
  NAND U37368 ( .A(n26653), .B(creg[552]), .Z(n27651) );
  NAND U37369 ( .A(n27653), .B(n27654), .Z(c[551]) );
  NAND U37370 ( .A(n26658), .B(o[551]), .Z(n27654) );
  NAND U37371 ( .A(n26653), .B(creg[551]), .Z(n27653) );
  NAND U37372 ( .A(n27655), .B(n27656), .Z(c[550]) );
  NAND U37373 ( .A(n26658), .B(o[550]), .Z(n27656) );
  NAND U37374 ( .A(n26653), .B(creg[550]), .Z(n27655) );
  NAND U37375 ( .A(n27657), .B(n27658), .Z(c[54]) );
  NAND U37376 ( .A(n26658), .B(o[54]), .Z(n27658) );
  NAND U37377 ( .A(n26653), .B(creg[54]), .Z(n27657) );
  NAND U37378 ( .A(n27659), .B(n27660), .Z(c[549]) );
  NAND U37379 ( .A(n26658), .B(o[549]), .Z(n27660) );
  NAND U37380 ( .A(n26653), .B(creg[549]), .Z(n27659) );
  NAND U37381 ( .A(n27661), .B(n27662), .Z(c[548]) );
  NAND U37382 ( .A(n26658), .B(o[548]), .Z(n27662) );
  NAND U37383 ( .A(n26653), .B(creg[548]), .Z(n27661) );
  NAND U37384 ( .A(n27663), .B(n27664), .Z(c[547]) );
  NAND U37385 ( .A(n26658), .B(o[547]), .Z(n27664) );
  NAND U37386 ( .A(n26653), .B(creg[547]), .Z(n27663) );
  NAND U37387 ( .A(n27665), .B(n27666), .Z(c[546]) );
  NAND U37388 ( .A(n26658), .B(o[546]), .Z(n27666) );
  NAND U37389 ( .A(n26653), .B(creg[546]), .Z(n27665) );
  NAND U37390 ( .A(n27667), .B(n27668), .Z(c[545]) );
  NAND U37391 ( .A(n26658), .B(o[545]), .Z(n27668) );
  NAND U37392 ( .A(n26653), .B(creg[545]), .Z(n27667) );
  NAND U37393 ( .A(n27669), .B(n27670), .Z(c[544]) );
  NAND U37394 ( .A(n26658), .B(o[544]), .Z(n27670) );
  NAND U37395 ( .A(n26653), .B(creg[544]), .Z(n27669) );
  NAND U37396 ( .A(n27671), .B(n27672), .Z(c[543]) );
  NAND U37397 ( .A(n26658), .B(o[543]), .Z(n27672) );
  NAND U37398 ( .A(n26653), .B(creg[543]), .Z(n27671) );
  NAND U37399 ( .A(n27673), .B(n27674), .Z(c[542]) );
  NAND U37400 ( .A(n26658), .B(o[542]), .Z(n27674) );
  NAND U37401 ( .A(n26653), .B(creg[542]), .Z(n27673) );
  NAND U37402 ( .A(n27675), .B(n27676), .Z(c[541]) );
  NAND U37403 ( .A(n26658), .B(o[541]), .Z(n27676) );
  NAND U37404 ( .A(n26653), .B(creg[541]), .Z(n27675) );
  NAND U37405 ( .A(n27677), .B(n27678), .Z(c[540]) );
  NAND U37406 ( .A(n26658), .B(o[540]), .Z(n27678) );
  NAND U37407 ( .A(n26653), .B(creg[540]), .Z(n27677) );
  NAND U37408 ( .A(n27679), .B(n27680), .Z(c[53]) );
  NAND U37409 ( .A(n26658), .B(o[53]), .Z(n27680) );
  NAND U37410 ( .A(n26653), .B(creg[53]), .Z(n27679) );
  NAND U37411 ( .A(n27681), .B(n27682), .Z(c[539]) );
  NAND U37412 ( .A(n26658), .B(o[539]), .Z(n27682) );
  NAND U37413 ( .A(n26653), .B(creg[539]), .Z(n27681) );
  NAND U37414 ( .A(n27683), .B(n27684), .Z(c[538]) );
  NAND U37415 ( .A(n26658), .B(o[538]), .Z(n27684) );
  NAND U37416 ( .A(n26653), .B(creg[538]), .Z(n27683) );
  NAND U37417 ( .A(n27685), .B(n27686), .Z(c[537]) );
  NAND U37418 ( .A(n26658), .B(o[537]), .Z(n27686) );
  NAND U37419 ( .A(n26653), .B(creg[537]), .Z(n27685) );
  NAND U37420 ( .A(n27687), .B(n27688), .Z(c[536]) );
  NAND U37421 ( .A(n26658), .B(o[536]), .Z(n27688) );
  NAND U37422 ( .A(n26653), .B(creg[536]), .Z(n27687) );
  NAND U37423 ( .A(n27689), .B(n27690), .Z(c[535]) );
  NAND U37424 ( .A(n26658), .B(o[535]), .Z(n27690) );
  NAND U37425 ( .A(n26653), .B(creg[535]), .Z(n27689) );
  NAND U37426 ( .A(n27691), .B(n27692), .Z(c[534]) );
  NAND U37427 ( .A(n26658), .B(o[534]), .Z(n27692) );
  NAND U37428 ( .A(n26653), .B(creg[534]), .Z(n27691) );
  NAND U37429 ( .A(n27693), .B(n27694), .Z(c[533]) );
  NAND U37430 ( .A(n26658), .B(o[533]), .Z(n27694) );
  NAND U37431 ( .A(n26653), .B(creg[533]), .Z(n27693) );
  NAND U37432 ( .A(n27695), .B(n27696), .Z(c[532]) );
  NAND U37433 ( .A(n26658), .B(o[532]), .Z(n27696) );
  NAND U37434 ( .A(n26653), .B(creg[532]), .Z(n27695) );
  NAND U37435 ( .A(n27697), .B(n27698), .Z(c[531]) );
  NAND U37436 ( .A(n26658), .B(o[531]), .Z(n27698) );
  NAND U37437 ( .A(n26653), .B(creg[531]), .Z(n27697) );
  NAND U37438 ( .A(n27699), .B(n27700), .Z(c[530]) );
  NAND U37439 ( .A(n26658), .B(o[530]), .Z(n27700) );
  NAND U37440 ( .A(n26653), .B(creg[530]), .Z(n27699) );
  NAND U37441 ( .A(n27701), .B(n27702), .Z(c[52]) );
  NAND U37442 ( .A(n26658), .B(o[52]), .Z(n27702) );
  NAND U37443 ( .A(n26653), .B(creg[52]), .Z(n27701) );
  NAND U37444 ( .A(n27703), .B(n27704), .Z(c[529]) );
  NAND U37445 ( .A(n26658), .B(o[529]), .Z(n27704) );
  NAND U37446 ( .A(n26653), .B(creg[529]), .Z(n27703) );
  NAND U37447 ( .A(n27705), .B(n27706), .Z(c[528]) );
  NAND U37448 ( .A(n26658), .B(o[528]), .Z(n27706) );
  NAND U37449 ( .A(n26653), .B(creg[528]), .Z(n27705) );
  NAND U37450 ( .A(n27707), .B(n27708), .Z(c[527]) );
  NAND U37451 ( .A(n26658), .B(o[527]), .Z(n27708) );
  NAND U37452 ( .A(n26653), .B(creg[527]), .Z(n27707) );
  NAND U37453 ( .A(n27709), .B(n27710), .Z(c[526]) );
  NAND U37454 ( .A(n26658), .B(o[526]), .Z(n27710) );
  NAND U37455 ( .A(n26653), .B(creg[526]), .Z(n27709) );
  NAND U37456 ( .A(n27711), .B(n27712), .Z(c[525]) );
  NAND U37457 ( .A(n26658), .B(o[525]), .Z(n27712) );
  NAND U37458 ( .A(n26653), .B(creg[525]), .Z(n27711) );
  NAND U37459 ( .A(n27713), .B(n27714), .Z(c[524]) );
  NAND U37460 ( .A(n26658), .B(o[524]), .Z(n27714) );
  NAND U37461 ( .A(n26653), .B(creg[524]), .Z(n27713) );
  NAND U37462 ( .A(n27715), .B(n27716), .Z(c[523]) );
  NAND U37463 ( .A(n26658), .B(o[523]), .Z(n27716) );
  NAND U37464 ( .A(n26653), .B(creg[523]), .Z(n27715) );
  NAND U37465 ( .A(n27717), .B(n27718), .Z(c[522]) );
  NAND U37466 ( .A(n26658), .B(o[522]), .Z(n27718) );
  NAND U37467 ( .A(n26653), .B(creg[522]), .Z(n27717) );
  NAND U37468 ( .A(n27719), .B(n27720), .Z(c[521]) );
  NAND U37469 ( .A(n26658), .B(o[521]), .Z(n27720) );
  NAND U37470 ( .A(n26653), .B(creg[521]), .Z(n27719) );
  NAND U37471 ( .A(n27721), .B(n27722), .Z(c[520]) );
  NAND U37472 ( .A(n26658), .B(o[520]), .Z(n27722) );
  NAND U37473 ( .A(n26653), .B(creg[520]), .Z(n27721) );
  NAND U37474 ( .A(n27723), .B(n27724), .Z(c[51]) );
  NAND U37475 ( .A(n26658), .B(o[51]), .Z(n27724) );
  NAND U37476 ( .A(n26653), .B(creg[51]), .Z(n27723) );
  NAND U37477 ( .A(n27725), .B(n27726), .Z(c[519]) );
  NAND U37478 ( .A(n26658), .B(o[519]), .Z(n27726) );
  NAND U37479 ( .A(n26653), .B(creg[519]), .Z(n27725) );
  NAND U37480 ( .A(n27727), .B(n27728), .Z(c[518]) );
  NAND U37481 ( .A(n26658), .B(o[518]), .Z(n27728) );
  NAND U37482 ( .A(n26653), .B(creg[518]), .Z(n27727) );
  NAND U37483 ( .A(n27729), .B(n27730), .Z(c[517]) );
  NAND U37484 ( .A(n26658), .B(o[517]), .Z(n27730) );
  NAND U37485 ( .A(n26653), .B(creg[517]), .Z(n27729) );
  NAND U37486 ( .A(n27731), .B(n27732), .Z(c[516]) );
  NAND U37487 ( .A(n26658), .B(o[516]), .Z(n27732) );
  NAND U37488 ( .A(n26653), .B(creg[516]), .Z(n27731) );
  NAND U37489 ( .A(n27733), .B(n27734), .Z(c[515]) );
  NAND U37490 ( .A(n26658), .B(o[515]), .Z(n27734) );
  NAND U37491 ( .A(n26653), .B(creg[515]), .Z(n27733) );
  NAND U37492 ( .A(n27735), .B(n27736), .Z(c[514]) );
  NAND U37493 ( .A(n26658), .B(o[514]), .Z(n27736) );
  NAND U37494 ( .A(n26653), .B(creg[514]), .Z(n27735) );
  NAND U37495 ( .A(n27737), .B(n27738), .Z(c[513]) );
  NAND U37496 ( .A(n26658), .B(o[513]), .Z(n27738) );
  NAND U37497 ( .A(n26653), .B(creg[513]), .Z(n27737) );
  NAND U37498 ( .A(n27739), .B(n27740), .Z(c[512]) );
  NAND U37499 ( .A(n26658), .B(o[512]), .Z(n27740) );
  NAND U37500 ( .A(n26653), .B(creg[512]), .Z(n27739) );
  NAND U37501 ( .A(n27741), .B(n27742), .Z(c[511]) );
  NAND U37502 ( .A(n26658), .B(o[511]), .Z(n27742) );
  NAND U37503 ( .A(n26653), .B(creg[511]), .Z(n27741) );
  NAND U37504 ( .A(n27743), .B(n27744), .Z(c[510]) );
  NAND U37505 ( .A(n26658), .B(o[510]), .Z(n27744) );
  NAND U37506 ( .A(n26653), .B(creg[510]), .Z(n27743) );
  NAND U37507 ( .A(n27745), .B(n27746), .Z(c[50]) );
  NAND U37508 ( .A(n26658), .B(o[50]), .Z(n27746) );
  NAND U37509 ( .A(n26653), .B(creg[50]), .Z(n27745) );
  NAND U37510 ( .A(n27747), .B(n27748), .Z(c[509]) );
  NAND U37511 ( .A(n26658), .B(o[509]), .Z(n27748) );
  NAND U37512 ( .A(n26653), .B(creg[509]), .Z(n27747) );
  NAND U37513 ( .A(n27749), .B(n27750), .Z(c[508]) );
  NAND U37514 ( .A(n26658), .B(o[508]), .Z(n27750) );
  NAND U37515 ( .A(n26653), .B(creg[508]), .Z(n27749) );
  NAND U37516 ( .A(n27751), .B(n27752), .Z(c[507]) );
  NAND U37517 ( .A(n26658), .B(o[507]), .Z(n27752) );
  NAND U37518 ( .A(n26653), .B(creg[507]), .Z(n27751) );
  NAND U37519 ( .A(n27753), .B(n27754), .Z(c[506]) );
  NAND U37520 ( .A(n26658), .B(o[506]), .Z(n27754) );
  NAND U37521 ( .A(n26653), .B(creg[506]), .Z(n27753) );
  NAND U37522 ( .A(n27755), .B(n27756), .Z(c[505]) );
  NAND U37523 ( .A(n26658), .B(o[505]), .Z(n27756) );
  NAND U37524 ( .A(n26653), .B(creg[505]), .Z(n27755) );
  NAND U37525 ( .A(n27757), .B(n27758), .Z(c[504]) );
  NAND U37526 ( .A(n26658), .B(o[504]), .Z(n27758) );
  NAND U37527 ( .A(n26653), .B(creg[504]), .Z(n27757) );
  NAND U37528 ( .A(n27759), .B(n27760), .Z(c[503]) );
  NAND U37529 ( .A(n26658), .B(o[503]), .Z(n27760) );
  NAND U37530 ( .A(n26653), .B(creg[503]), .Z(n27759) );
  NAND U37531 ( .A(n27761), .B(n27762), .Z(c[502]) );
  NAND U37532 ( .A(n26658), .B(o[502]), .Z(n27762) );
  NAND U37533 ( .A(n26653), .B(creg[502]), .Z(n27761) );
  NAND U37534 ( .A(n27763), .B(n27764), .Z(c[501]) );
  NAND U37535 ( .A(n26658), .B(o[501]), .Z(n27764) );
  NAND U37536 ( .A(n26653), .B(creg[501]), .Z(n27763) );
  NAND U37537 ( .A(n27765), .B(n27766), .Z(c[500]) );
  NAND U37538 ( .A(n26658), .B(o[500]), .Z(n27766) );
  NAND U37539 ( .A(n26653), .B(creg[500]), .Z(n27765) );
  NAND U37540 ( .A(n27767), .B(n27768), .Z(c[4]) );
  NAND U37541 ( .A(n26658), .B(o[4]), .Z(n27768) );
  NAND U37542 ( .A(n26653), .B(creg[4]), .Z(n27767) );
  NAND U37543 ( .A(n27769), .B(n27770), .Z(c[49]) );
  NAND U37544 ( .A(n26658), .B(o[49]), .Z(n27770) );
  NAND U37545 ( .A(n26653), .B(creg[49]), .Z(n27769) );
  NAND U37546 ( .A(n27771), .B(n27772), .Z(c[499]) );
  NAND U37547 ( .A(n26658), .B(o[499]), .Z(n27772) );
  NAND U37548 ( .A(n26653), .B(creg[499]), .Z(n27771) );
  NAND U37549 ( .A(n27773), .B(n27774), .Z(c[498]) );
  NAND U37550 ( .A(n26658), .B(o[498]), .Z(n27774) );
  NAND U37551 ( .A(n26653), .B(creg[498]), .Z(n27773) );
  NAND U37552 ( .A(n27775), .B(n27776), .Z(c[497]) );
  NAND U37553 ( .A(n26658), .B(o[497]), .Z(n27776) );
  NAND U37554 ( .A(n26653), .B(creg[497]), .Z(n27775) );
  NAND U37555 ( .A(n27777), .B(n27778), .Z(c[496]) );
  NAND U37556 ( .A(n26658), .B(o[496]), .Z(n27778) );
  NAND U37557 ( .A(n26653), .B(creg[496]), .Z(n27777) );
  NAND U37558 ( .A(n27779), .B(n27780), .Z(c[495]) );
  NAND U37559 ( .A(n26658), .B(o[495]), .Z(n27780) );
  NAND U37560 ( .A(n26653), .B(creg[495]), .Z(n27779) );
  NAND U37561 ( .A(n27781), .B(n27782), .Z(c[494]) );
  NAND U37562 ( .A(n26658), .B(o[494]), .Z(n27782) );
  NAND U37563 ( .A(n26653), .B(creg[494]), .Z(n27781) );
  NAND U37564 ( .A(n27783), .B(n27784), .Z(c[493]) );
  NAND U37565 ( .A(n26658), .B(o[493]), .Z(n27784) );
  NAND U37566 ( .A(n26653), .B(creg[493]), .Z(n27783) );
  NAND U37567 ( .A(n27785), .B(n27786), .Z(c[492]) );
  NAND U37568 ( .A(n26658), .B(o[492]), .Z(n27786) );
  NAND U37569 ( .A(n26653), .B(creg[492]), .Z(n27785) );
  NAND U37570 ( .A(n27787), .B(n27788), .Z(c[491]) );
  NAND U37571 ( .A(n26658), .B(o[491]), .Z(n27788) );
  NAND U37572 ( .A(n26653), .B(creg[491]), .Z(n27787) );
  NAND U37573 ( .A(n27789), .B(n27790), .Z(c[490]) );
  NAND U37574 ( .A(n26658), .B(o[490]), .Z(n27790) );
  NAND U37575 ( .A(n26653), .B(creg[490]), .Z(n27789) );
  NAND U37576 ( .A(n27791), .B(n27792), .Z(c[48]) );
  NAND U37577 ( .A(n26658), .B(o[48]), .Z(n27792) );
  NAND U37578 ( .A(n26653), .B(creg[48]), .Z(n27791) );
  NAND U37579 ( .A(n27793), .B(n27794), .Z(c[489]) );
  NAND U37580 ( .A(n26658), .B(o[489]), .Z(n27794) );
  NAND U37581 ( .A(n26653), .B(creg[489]), .Z(n27793) );
  NAND U37582 ( .A(n27795), .B(n27796), .Z(c[488]) );
  NAND U37583 ( .A(n26658), .B(o[488]), .Z(n27796) );
  NAND U37584 ( .A(n26653), .B(creg[488]), .Z(n27795) );
  NAND U37585 ( .A(n27797), .B(n27798), .Z(c[487]) );
  NAND U37586 ( .A(n26658), .B(o[487]), .Z(n27798) );
  NAND U37587 ( .A(n26653), .B(creg[487]), .Z(n27797) );
  NAND U37588 ( .A(n27799), .B(n27800), .Z(c[486]) );
  NAND U37589 ( .A(n26658), .B(o[486]), .Z(n27800) );
  NAND U37590 ( .A(n26653), .B(creg[486]), .Z(n27799) );
  NAND U37591 ( .A(n27801), .B(n27802), .Z(c[485]) );
  NAND U37592 ( .A(n26658), .B(o[485]), .Z(n27802) );
  NAND U37593 ( .A(n26653), .B(creg[485]), .Z(n27801) );
  NAND U37594 ( .A(n27803), .B(n27804), .Z(c[484]) );
  NAND U37595 ( .A(n26658), .B(o[484]), .Z(n27804) );
  NAND U37596 ( .A(n26653), .B(creg[484]), .Z(n27803) );
  NAND U37597 ( .A(n27805), .B(n27806), .Z(c[483]) );
  NAND U37598 ( .A(n26658), .B(o[483]), .Z(n27806) );
  NAND U37599 ( .A(n26653), .B(creg[483]), .Z(n27805) );
  NAND U37600 ( .A(n27807), .B(n27808), .Z(c[482]) );
  NAND U37601 ( .A(n26658), .B(o[482]), .Z(n27808) );
  NAND U37602 ( .A(n26653), .B(creg[482]), .Z(n27807) );
  NAND U37603 ( .A(n27809), .B(n27810), .Z(c[481]) );
  NAND U37604 ( .A(n26658), .B(o[481]), .Z(n27810) );
  NAND U37605 ( .A(n26653), .B(creg[481]), .Z(n27809) );
  NAND U37606 ( .A(n27811), .B(n27812), .Z(c[480]) );
  NAND U37607 ( .A(n26658), .B(o[480]), .Z(n27812) );
  NAND U37608 ( .A(n26653), .B(creg[480]), .Z(n27811) );
  NAND U37609 ( .A(n27813), .B(n27814), .Z(c[47]) );
  NAND U37610 ( .A(n26658), .B(o[47]), .Z(n27814) );
  NAND U37611 ( .A(n26653), .B(creg[47]), .Z(n27813) );
  NAND U37612 ( .A(n27815), .B(n27816), .Z(c[479]) );
  NAND U37613 ( .A(n26658), .B(o[479]), .Z(n27816) );
  NAND U37614 ( .A(n26653), .B(creg[479]), .Z(n27815) );
  NAND U37615 ( .A(n27817), .B(n27818), .Z(c[478]) );
  NAND U37616 ( .A(n26658), .B(o[478]), .Z(n27818) );
  NAND U37617 ( .A(n26653), .B(creg[478]), .Z(n27817) );
  NAND U37618 ( .A(n27819), .B(n27820), .Z(c[477]) );
  NAND U37619 ( .A(n26658), .B(o[477]), .Z(n27820) );
  NAND U37620 ( .A(n26653), .B(creg[477]), .Z(n27819) );
  NAND U37621 ( .A(n27821), .B(n27822), .Z(c[476]) );
  NAND U37622 ( .A(n26658), .B(o[476]), .Z(n27822) );
  NAND U37623 ( .A(n26653), .B(creg[476]), .Z(n27821) );
  NAND U37624 ( .A(n27823), .B(n27824), .Z(c[475]) );
  NAND U37625 ( .A(n26658), .B(o[475]), .Z(n27824) );
  NAND U37626 ( .A(n26653), .B(creg[475]), .Z(n27823) );
  NAND U37627 ( .A(n27825), .B(n27826), .Z(c[474]) );
  NAND U37628 ( .A(n26658), .B(o[474]), .Z(n27826) );
  NAND U37629 ( .A(n26653), .B(creg[474]), .Z(n27825) );
  NAND U37630 ( .A(n27827), .B(n27828), .Z(c[473]) );
  NAND U37631 ( .A(n26658), .B(o[473]), .Z(n27828) );
  NAND U37632 ( .A(n26653), .B(creg[473]), .Z(n27827) );
  NAND U37633 ( .A(n27829), .B(n27830), .Z(c[472]) );
  NAND U37634 ( .A(n26658), .B(o[472]), .Z(n27830) );
  NAND U37635 ( .A(n26653), .B(creg[472]), .Z(n27829) );
  NAND U37636 ( .A(n27831), .B(n27832), .Z(c[471]) );
  NAND U37637 ( .A(n26658), .B(o[471]), .Z(n27832) );
  NAND U37638 ( .A(n26653), .B(creg[471]), .Z(n27831) );
  NAND U37639 ( .A(n27833), .B(n27834), .Z(c[470]) );
  NAND U37640 ( .A(n26658), .B(o[470]), .Z(n27834) );
  NAND U37641 ( .A(n26653), .B(creg[470]), .Z(n27833) );
  NAND U37642 ( .A(n27835), .B(n27836), .Z(c[46]) );
  NAND U37643 ( .A(n26658), .B(o[46]), .Z(n27836) );
  NAND U37644 ( .A(n26653), .B(creg[46]), .Z(n27835) );
  NAND U37645 ( .A(n27837), .B(n27838), .Z(c[469]) );
  NAND U37646 ( .A(n26658), .B(o[469]), .Z(n27838) );
  NAND U37647 ( .A(n26653), .B(creg[469]), .Z(n27837) );
  NAND U37648 ( .A(n27839), .B(n27840), .Z(c[468]) );
  NAND U37649 ( .A(n26658), .B(o[468]), .Z(n27840) );
  NAND U37650 ( .A(n26653), .B(creg[468]), .Z(n27839) );
  NAND U37651 ( .A(n27841), .B(n27842), .Z(c[467]) );
  NAND U37652 ( .A(n26658), .B(o[467]), .Z(n27842) );
  NAND U37653 ( .A(n26653), .B(creg[467]), .Z(n27841) );
  NAND U37654 ( .A(n27843), .B(n27844), .Z(c[466]) );
  NAND U37655 ( .A(n26658), .B(o[466]), .Z(n27844) );
  NAND U37656 ( .A(n26653), .B(creg[466]), .Z(n27843) );
  NAND U37657 ( .A(n27845), .B(n27846), .Z(c[465]) );
  NAND U37658 ( .A(n26658), .B(o[465]), .Z(n27846) );
  NAND U37659 ( .A(n26653), .B(creg[465]), .Z(n27845) );
  NAND U37660 ( .A(n27847), .B(n27848), .Z(c[464]) );
  NAND U37661 ( .A(n26658), .B(o[464]), .Z(n27848) );
  NAND U37662 ( .A(n26653), .B(creg[464]), .Z(n27847) );
  NAND U37663 ( .A(n27849), .B(n27850), .Z(c[463]) );
  NAND U37664 ( .A(n26658), .B(o[463]), .Z(n27850) );
  NAND U37665 ( .A(n26653), .B(creg[463]), .Z(n27849) );
  NAND U37666 ( .A(n27851), .B(n27852), .Z(c[462]) );
  NAND U37667 ( .A(n26658), .B(o[462]), .Z(n27852) );
  NAND U37668 ( .A(n26653), .B(creg[462]), .Z(n27851) );
  NAND U37669 ( .A(n27853), .B(n27854), .Z(c[461]) );
  NAND U37670 ( .A(n26658), .B(o[461]), .Z(n27854) );
  NAND U37671 ( .A(n26653), .B(creg[461]), .Z(n27853) );
  NAND U37672 ( .A(n27855), .B(n27856), .Z(c[460]) );
  NAND U37673 ( .A(n26658), .B(o[460]), .Z(n27856) );
  NAND U37674 ( .A(n26653), .B(creg[460]), .Z(n27855) );
  NAND U37675 ( .A(n27857), .B(n27858), .Z(c[45]) );
  NAND U37676 ( .A(n26658), .B(o[45]), .Z(n27858) );
  NAND U37677 ( .A(n26653), .B(creg[45]), .Z(n27857) );
  NAND U37678 ( .A(n27859), .B(n27860), .Z(c[459]) );
  NAND U37679 ( .A(n26658), .B(o[459]), .Z(n27860) );
  NAND U37680 ( .A(n26653), .B(creg[459]), .Z(n27859) );
  NAND U37681 ( .A(n27861), .B(n27862), .Z(c[458]) );
  NAND U37682 ( .A(n26658), .B(o[458]), .Z(n27862) );
  NAND U37683 ( .A(n26653), .B(creg[458]), .Z(n27861) );
  NAND U37684 ( .A(n27863), .B(n27864), .Z(c[457]) );
  NAND U37685 ( .A(n26658), .B(o[457]), .Z(n27864) );
  NAND U37686 ( .A(n26653), .B(creg[457]), .Z(n27863) );
  NAND U37687 ( .A(n27865), .B(n27866), .Z(c[456]) );
  NAND U37688 ( .A(n26658), .B(o[456]), .Z(n27866) );
  NAND U37689 ( .A(n26653), .B(creg[456]), .Z(n27865) );
  NAND U37690 ( .A(n27867), .B(n27868), .Z(c[455]) );
  NAND U37691 ( .A(n26658), .B(o[455]), .Z(n27868) );
  NAND U37692 ( .A(n26653), .B(creg[455]), .Z(n27867) );
  NAND U37693 ( .A(n27869), .B(n27870), .Z(c[454]) );
  NAND U37694 ( .A(n26658), .B(o[454]), .Z(n27870) );
  NAND U37695 ( .A(n26653), .B(creg[454]), .Z(n27869) );
  NAND U37696 ( .A(n27871), .B(n27872), .Z(c[453]) );
  NAND U37697 ( .A(n26658), .B(o[453]), .Z(n27872) );
  NAND U37698 ( .A(n26653), .B(creg[453]), .Z(n27871) );
  NAND U37699 ( .A(n27873), .B(n27874), .Z(c[452]) );
  NAND U37700 ( .A(n26658), .B(o[452]), .Z(n27874) );
  NAND U37701 ( .A(n26653), .B(creg[452]), .Z(n27873) );
  NAND U37702 ( .A(n27875), .B(n27876), .Z(c[451]) );
  NAND U37703 ( .A(n26658), .B(o[451]), .Z(n27876) );
  NAND U37704 ( .A(n26653), .B(creg[451]), .Z(n27875) );
  NAND U37705 ( .A(n27877), .B(n27878), .Z(c[450]) );
  NAND U37706 ( .A(n26658), .B(o[450]), .Z(n27878) );
  NAND U37707 ( .A(n26653), .B(creg[450]), .Z(n27877) );
  NAND U37708 ( .A(n27879), .B(n27880), .Z(c[44]) );
  NAND U37709 ( .A(n26658), .B(o[44]), .Z(n27880) );
  NAND U37710 ( .A(n26653), .B(creg[44]), .Z(n27879) );
  NAND U37711 ( .A(n27881), .B(n27882), .Z(c[449]) );
  NAND U37712 ( .A(n26658), .B(o[449]), .Z(n27882) );
  NAND U37713 ( .A(n26653), .B(creg[449]), .Z(n27881) );
  NAND U37714 ( .A(n27883), .B(n27884), .Z(c[448]) );
  NAND U37715 ( .A(n26658), .B(o[448]), .Z(n27884) );
  NAND U37716 ( .A(n26653), .B(creg[448]), .Z(n27883) );
  NAND U37717 ( .A(n27885), .B(n27886), .Z(c[447]) );
  NAND U37718 ( .A(n26658), .B(o[447]), .Z(n27886) );
  NAND U37719 ( .A(n26653), .B(creg[447]), .Z(n27885) );
  NAND U37720 ( .A(n27887), .B(n27888), .Z(c[446]) );
  NAND U37721 ( .A(n26658), .B(o[446]), .Z(n27888) );
  NAND U37722 ( .A(n26653), .B(creg[446]), .Z(n27887) );
  NAND U37723 ( .A(n27889), .B(n27890), .Z(c[445]) );
  NAND U37724 ( .A(n26658), .B(o[445]), .Z(n27890) );
  NAND U37725 ( .A(n26653), .B(creg[445]), .Z(n27889) );
  NAND U37726 ( .A(n27891), .B(n27892), .Z(c[444]) );
  NAND U37727 ( .A(n26658), .B(o[444]), .Z(n27892) );
  NAND U37728 ( .A(n26653), .B(creg[444]), .Z(n27891) );
  NAND U37729 ( .A(n27893), .B(n27894), .Z(c[443]) );
  NAND U37730 ( .A(n26658), .B(o[443]), .Z(n27894) );
  NAND U37731 ( .A(n26653), .B(creg[443]), .Z(n27893) );
  NAND U37732 ( .A(n27895), .B(n27896), .Z(c[442]) );
  NAND U37733 ( .A(n26658), .B(o[442]), .Z(n27896) );
  NAND U37734 ( .A(n26653), .B(creg[442]), .Z(n27895) );
  NAND U37735 ( .A(n27897), .B(n27898), .Z(c[441]) );
  NAND U37736 ( .A(n26658), .B(o[441]), .Z(n27898) );
  NAND U37737 ( .A(n26653), .B(creg[441]), .Z(n27897) );
  NAND U37738 ( .A(n27899), .B(n27900), .Z(c[440]) );
  NAND U37739 ( .A(n26658), .B(o[440]), .Z(n27900) );
  NAND U37740 ( .A(n26653), .B(creg[440]), .Z(n27899) );
  NAND U37741 ( .A(n27901), .B(n27902), .Z(c[43]) );
  NAND U37742 ( .A(n26658), .B(o[43]), .Z(n27902) );
  NAND U37743 ( .A(n26653), .B(creg[43]), .Z(n27901) );
  NAND U37744 ( .A(n27903), .B(n27904), .Z(c[439]) );
  NAND U37745 ( .A(n26658), .B(o[439]), .Z(n27904) );
  NAND U37746 ( .A(n26653), .B(creg[439]), .Z(n27903) );
  NAND U37747 ( .A(n27905), .B(n27906), .Z(c[438]) );
  NAND U37748 ( .A(n26658), .B(o[438]), .Z(n27906) );
  NAND U37749 ( .A(n26653), .B(creg[438]), .Z(n27905) );
  NAND U37750 ( .A(n27907), .B(n27908), .Z(c[437]) );
  NAND U37751 ( .A(n26658), .B(o[437]), .Z(n27908) );
  NAND U37752 ( .A(n26653), .B(creg[437]), .Z(n27907) );
  NAND U37753 ( .A(n27909), .B(n27910), .Z(c[436]) );
  NAND U37754 ( .A(n26658), .B(o[436]), .Z(n27910) );
  NAND U37755 ( .A(n26653), .B(creg[436]), .Z(n27909) );
  NAND U37756 ( .A(n27911), .B(n27912), .Z(c[435]) );
  NAND U37757 ( .A(n26658), .B(o[435]), .Z(n27912) );
  NAND U37758 ( .A(n26653), .B(creg[435]), .Z(n27911) );
  NAND U37759 ( .A(n27913), .B(n27914), .Z(c[434]) );
  NAND U37760 ( .A(n26658), .B(o[434]), .Z(n27914) );
  NAND U37761 ( .A(n26653), .B(creg[434]), .Z(n27913) );
  NAND U37762 ( .A(n27915), .B(n27916), .Z(c[433]) );
  NAND U37763 ( .A(n26658), .B(o[433]), .Z(n27916) );
  NAND U37764 ( .A(n26653), .B(creg[433]), .Z(n27915) );
  NAND U37765 ( .A(n27917), .B(n27918), .Z(c[432]) );
  NAND U37766 ( .A(n26658), .B(o[432]), .Z(n27918) );
  NAND U37767 ( .A(n26653), .B(creg[432]), .Z(n27917) );
  NAND U37768 ( .A(n27919), .B(n27920), .Z(c[431]) );
  NAND U37769 ( .A(n26658), .B(o[431]), .Z(n27920) );
  NAND U37770 ( .A(n26653), .B(creg[431]), .Z(n27919) );
  NAND U37771 ( .A(n27921), .B(n27922), .Z(c[430]) );
  NAND U37772 ( .A(n26658), .B(o[430]), .Z(n27922) );
  NAND U37773 ( .A(n26653), .B(creg[430]), .Z(n27921) );
  NAND U37774 ( .A(n27923), .B(n27924), .Z(c[42]) );
  NAND U37775 ( .A(n26658), .B(o[42]), .Z(n27924) );
  NAND U37776 ( .A(n26653), .B(creg[42]), .Z(n27923) );
  NAND U37777 ( .A(n27925), .B(n27926), .Z(c[429]) );
  NAND U37778 ( .A(n26658), .B(o[429]), .Z(n27926) );
  NAND U37779 ( .A(n26653), .B(creg[429]), .Z(n27925) );
  NAND U37780 ( .A(n27927), .B(n27928), .Z(c[428]) );
  NAND U37781 ( .A(n26658), .B(o[428]), .Z(n27928) );
  NAND U37782 ( .A(n26653), .B(creg[428]), .Z(n27927) );
  NAND U37783 ( .A(n27929), .B(n27930), .Z(c[427]) );
  NAND U37784 ( .A(n26658), .B(o[427]), .Z(n27930) );
  NAND U37785 ( .A(n26653), .B(creg[427]), .Z(n27929) );
  NAND U37786 ( .A(n27931), .B(n27932), .Z(c[426]) );
  NAND U37787 ( .A(n26658), .B(o[426]), .Z(n27932) );
  NAND U37788 ( .A(n26653), .B(creg[426]), .Z(n27931) );
  NAND U37789 ( .A(n27933), .B(n27934), .Z(c[425]) );
  NAND U37790 ( .A(n26658), .B(o[425]), .Z(n27934) );
  NAND U37791 ( .A(n26653), .B(creg[425]), .Z(n27933) );
  NAND U37792 ( .A(n27935), .B(n27936), .Z(c[424]) );
  NAND U37793 ( .A(n26658), .B(o[424]), .Z(n27936) );
  NAND U37794 ( .A(n26653), .B(creg[424]), .Z(n27935) );
  NAND U37795 ( .A(n27937), .B(n27938), .Z(c[423]) );
  NAND U37796 ( .A(n26658), .B(o[423]), .Z(n27938) );
  NAND U37797 ( .A(n26653), .B(creg[423]), .Z(n27937) );
  NAND U37798 ( .A(n27939), .B(n27940), .Z(c[422]) );
  NAND U37799 ( .A(n26658), .B(o[422]), .Z(n27940) );
  NAND U37800 ( .A(n26653), .B(creg[422]), .Z(n27939) );
  NAND U37801 ( .A(n27941), .B(n27942), .Z(c[421]) );
  NAND U37802 ( .A(n26658), .B(o[421]), .Z(n27942) );
  NAND U37803 ( .A(n26653), .B(creg[421]), .Z(n27941) );
  NAND U37804 ( .A(n27943), .B(n27944), .Z(c[420]) );
  NAND U37805 ( .A(n26658), .B(o[420]), .Z(n27944) );
  NAND U37806 ( .A(n26653), .B(creg[420]), .Z(n27943) );
  NAND U37807 ( .A(n27945), .B(n27946), .Z(c[41]) );
  NAND U37808 ( .A(n26658), .B(o[41]), .Z(n27946) );
  NAND U37809 ( .A(n26653), .B(creg[41]), .Z(n27945) );
  NAND U37810 ( .A(n27947), .B(n27948), .Z(c[419]) );
  NAND U37811 ( .A(n26658), .B(o[419]), .Z(n27948) );
  NAND U37812 ( .A(n26653), .B(creg[419]), .Z(n27947) );
  NAND U37813 ( .A(n27949), .B(n27950), .Z(c[418]) );
  NAND U37814 ( .A(n26658), .B(o[418]), .Z(n27950) );
  NAND U37815 ( .A(n26653), .B(creg[418]), .Z(n27949) );
  NAND U37816 ( .A(n27951), .B(n27952), .Z(c[417]) );
  NAND U37817 ( .A(n26658), .B(o[417]), .Z(n27952) );
  NAND U37818 ( .A(n26653), .B(creg[417]), .Z(n27951) );
  NAND U37819 ( .A(n27953), .B(n27954), .Z(c[416]) );
  NAND U37820 ( .A(n26658), .B(o[416]), .Z(n27954) );
  NAND U37821 ( .A(n26653), .B(creg[416]), .Z(n27953) );
  NAND U37822 ( .A(n27955), .B(n27956), .Z(c[415]) );
  NAND U37823 ( .A(n26658), .B(o[415]), .Z(n27956) );
  NAND U37824 ( .A(n26653), .B(creg[415]), .Z(n27955) );
  NAND U37825 ( .A(n27957), .B(n27958), .Z(c[414]) );
  NAND U37826 ( .A(n26658), .B(o[414]), .Z(n27958) );
  NAND U37827 ( .A(n26653), .B(creg[414]), .Z(n27957) );
  NAND U37828 ( .A(n27959), .B(n27960), .Z(c[413]) );
  NAND U37829 ( .A(n26658), .B(o[413]), .Z(n27960) );
  NAND U37830 ( .A(n26653), .B(creg[413]), .Z(n27959) );
  NAND U37831 ( .A(n27961), .B(n27962), .Z(c[412]) );
  NAND U37832 ( .A(n26658), .B(o[412]), .Z(n27962) );
  NAND U37833 ( .A(n26653), .B(creg[412]), .Z(n27961) );
  NAND U37834 ( .A(n27963), .B(n27964), .Z(c[411]) );
  NAND U37835 ( .A(n26658), .B(o[411]), .Z(n27964) );
  NAND U37836 ( .A(n26653), .B(creg[411]), .Z(n27963) );
  NAND U37837 ( .A(n27965), .B(n27966), .Z(c[410]) );
  NAND U37838 ( .A(n26658), .B(o[410]), .Z(n27966) );
  NAND U37839 ( .A(n26653), .B(creg[410]), .Z(n27965) );
  NAND U37840 ( .A(n27967), .B(n27968), .Z(c[40]) );
  NAND U37841 ( .A(n26658), .B(o[40]), .Z(n27968) );
  NAND U37842 ( .A(n26653), .B(creg[40]), .Z(n27967) );
  NAND U37843 ( .A(n27969), .B(n27970), .Z(c[409]) );
  NAND U37844 ( .A(n26658), .B(o[409]), .Z(n27970) );
  NAND U37845 ( .A(n26653), .B(creg[409]), .Z(n27969) );
  NAND U37846 ( .A(n27971), .B(n27972), .Z(c[408]) );
  NAND U37847 ( .A(n26658), .B(o[408]), .Z(n27972) );
  NAND U37848 ( .A(n26653), .B(creg[408]), .Z(n27971) );
  NAND U37849 ( .A(n27973), .B(n27974), .Z(c[407]) );
  NAND U37850 ( .A(n26658), .B(o[407]), .Z(n27974) );
  NAND U37851 ( .A(n26653), .B(creg[407]), .Z(n27973) );
  NAND U37852 ( .A(n27975), .B(n27976), .Z(c[406]) );
  NAND U37853 ( .A(n26658), .B(o[406]), .Z(n27976) );
  NAND U37854 ( .A(n26653), .B(creg[406]), .Z(n27975) );
  NAND U37855 ( .A(n27977), .B(n27978), .Z(c[405]) );
  NAND U37856 ( .A(n26658), .B(o[405]), .Z(n27978) );
  NAND U37857 ( .A(n26653), .B(creg[405]), .Z(n27977) );
  NAND U37858 ( .A(n27979), .B(n27980), .Z(c[404]) );
  NAND U37859 ( .A(n26658), .B(o[404]), .Z(n27980) );
  NAND U37860 ( .A(n26653), .B(creg[404]), .Z(n27979) );
  NAND U37861 ( .A(n27981), .B(n27982), .Z(c[403]) );
  NAND U37862 ( .A(n26658), .B(o[403]), .Z(n27982) );
  NAND U37863 ( .A(n26653), .B(creg[403]), .Z(n27981) );
  NAND U37864 ( .A(n27983), .B(n27984), .Z(c[402]) );
  NAND U37865 ( .A(n26658), .B(o[402]), .Z(n27984) );
  NAND U37866 ( .A(n26653), .B(creg[402]), .Z(n27983) );
  NAND U37867 ( .A(n27985), .B(n27986), .Z(c[401]) );
  NAND U37868 ( .A(n26658), .B(o[401]), .Z(n27986) );
  NAND U37869 ( .A(n26653), .B(creg[401]), .Z(n27985) );
  NAND U37870 ( .A(n27987), .B(n27988), .Z(c[400]) );
  NAND U37871 ( .A(n26658), .B(o[400]), .Z(n27988) );
  NAND U37872 ( .A(n26653), .B(creg[400]), .Z(n27987) );
  NAND U37873 ( .A(n27989), .B(n27990), .Z(c[3]) );
  NAND U37874 ( .A(n26658), .B(o[3]), .Z(n27990) );
  NAND U37875 ( .A(n26653), .B(creg[3]), .Z(n27989) );
  NAND U37876 ( .A(n27991), .B(n27992), .Z(c[39]) );
  NAND U37877 ( .A(n26658), .B(o[39]), .Z(n27992) );
  NAND U37878 ( .A(n26653), .B(creg[39]), .Z(n27991) );
  NAND U37879 ( .A(n27993), .B(n27994), .Z(c[399]) );
  NAND U37880 ( .A(n26658), .B(o[399]), .Z(n27994) );
  NAND U37881 ( .A(n26653), .B(creg[399]), .Z(n27993) );
  NAND U37882 ( .A(n27995), .B(n27996), .Z(c[398]) );
  NAND U37883 ( .A(n26658), .B(o[398]), .Z(n27996) );
  NAND U37884 ( .A(n26653), .B(creg[398]), .Z(n27995) );
  NAND U37885 ( .A(n27997), .B(n27998), .Z(c[397]) );
  NAND U37886 ( .A(n26658), .B(o[397]), .Z(n27998) );
  NAND U37887 ( .A(n26653), .B(creg[397]), .Z(n27997) );
  NAND U37888 ( .A(n27999), .B(n28000), .Z(c[396]) );
  NAND U37889 ( .A(n26658), .B(o[396]), .Z(n28000) );
  NAND U37890 ( .A(n26653), .B(creg[396]), .Z(n27999) );
  NAND U37891 ( .A(n28001), .B(n28002), .Z(c[395]) );
  NAND U37892 ( .A(n26658), .B(o[395]), .Z(n28002) );
  NAND U37893 ( .A(n26653), .B(creg[395]), .Z(n28001) );
  NAND U37894 ( .A(n28003), .B(n28004), .Z(c[394]) );
  NAND U37895 ( .A(n26658), .B(o[394]), .Z(n28004) );
  NAND U37896 ( .A(n26653), .B(creg[394]), .Z(n28003) );
  NAND U37897 ( .A(n28005), .B(n28006), .Z(c[393]) );
  NAND U37898 ( .A(n26658), .B(o[393]), .Z(n28006) );
  NAND U37899 ( .A(n26653), .B(creg[393]), .Z(n28005) );
  NAND U37900 ( .A(n28007), .B(n28008), .Z(c[392]) );
  NAND U37901 ( .A(n26658), .B(o[392]), .Z(n28008) );
  NAND U37902 ( .A(n26653), .B(creg[392]), .Z(n28007) );
  NAND U37903 ( .A(n28009), .B(n28010), .Z(c[391]) );
  NAND U37904 ( .A(n26658), .B(o[391]), .Z(n28010) );
  NAND U37905 ( .A(n26653), .B(creg[391]), .Z(n28009) );
  NAND U37906 ( .A(n28011), .B(n28012), .Z(c[390]) );
  NAND U37907 ( .A(n26658), .B(o[390]), .Z(n28012) );
  NAND U37908 ( .A(n26653), .B(creg[390]), .Z(n28011) );
  NAND U37909 ( .A(n28013), .B(n28014), .Z(c[38]) );
  NAND U37910 ( .A(n26658), .B(o[38]), .Z(n28014) );
  NAND U37911 ( .A(n26653), .B(creg[38]), .Z(n28013) );
  NAND U37912 ( .A(n28015), .B(n28016), .Z(c[389]) );
  NAND U37913 ( .A(n26658), .B(o[389]), .Z(n28016) );
  NAND U37914 ( .A(n26653), .B(creg[389]), .Z(n28015) );
  NAND U37915 ( .A(n28017), .B(n28018), .Z(c[388]) );
  NAND U37916 ( .A(n26658), .B(o[388]), .Z(n28018) );
  NAND U37917 ( .A(n26653), .B(creg[388]), .Z(n28017) );
  NAND U37918 ( .A(n28019), .B(n28020), .Z(c[387]) );
  NAND U37919 ( .A(n26658), .B(o[387]), .Z(n28020) );
  NAND U37920 ( .A(n26653), .B(creg[387]), .Z(n28019) );
  NAND U37921 ( .A(n28021), .B(n28022), .Z(c[386]) );
  NAND U37922 ( .A(n26658), .B(o[386]), .Z(n28022) );
  NAND U37923 ( .A(n26653), .B(creg[386]), .Z(n28021) );
  NAND U37924 ( .A(n28023), .B(n28024), .Z(c[385]) );
  NAND U37925 ( .A(n26658), .B(o[385]), .Z(n28024) );
  NAND U37926 ( .A(n26653), .B(creg[385]), .Z(n28023) );
  NAND U37927 ( .A(n28025), .B(n28026), .Z(c[384]) );
  NAND U37928 ( .A(n26658), .B(o[384]), .Z(n28026) );
  NAND U37929 ( .A(n26653), .B(creg[384]), .Z(n28025) );
  NAND U37930 ( .A(n28027), .B(n28028), .Z(c[383]) );
  NAND U37931 ( .A(n26658), .B(o[383]), .Z(n28028) );
  NAND U37932 ( .A(n26653), .B(creg[383]), .Z(n28027) );
  NAND U37933 ( .A(n28029), .B(n28030), .Z(c[382]) );
  NAND U37934 ( .A(n26658), .B(o[382]), .Z(n28030) );
  NAND U37935 ( .A(n26653), .B(creg[382]), .Z(n28029) );
  NAND U37936 ( .A(n28031), .B(n28032), .Z(c[381]) );
  NAND U37937 ( .A(n26658), .B(o[381]), .Z(n28032) );
  NAND U37938 ( .A(n26653), .B(creg[381]), .Z(n28031) );
  NAND U37939 ( .A(n28033), .B(n28034), .Z(c[380]) );
  NAND U37940 ( .A(n26658), .B(o[380]), .Z(n28034) );
  NAND U37941 ( .A(n26653), .B(creg[380]), .Z(n28033) );
  NAND U37942 ( .A(n28035), .B(n28036), .Z(c[37]) );
  NAND U37943 ( .A(n26658), .B(o[37]), .Z(n28036) );
  NAND U37944 ( .A(n26653), .B(creg[37]), .Z(n28035) );
  NAND U37945 ( .A(n28037), .B(n28038), .Z(c[379]) );
  NAND U37946 ( .A(n26658), .B(o[379]), .Z(n28038) );
  NAND U37947 ( .A(n26653), .B(creg[379]), .Z(n28037) );
  NAND U37948 ( .A(n28039), .B(n28040), .Z(c[378]) );
  NAND U37949 ( .A(n26658), .B(o[378]), .Z(n28040) );
  NAND U37950 ( .A(n26653), .B(creg[378]), .Z(n28039) );
  NAND U37951 ( .A(n28041), .B(n28042), .Z(c[377]) );
  NAND U37952 ( .A(n26658), .B(o[377]), .Z(n28042) );
  NAND U37953 ( .A(n26653), .B(creg[377]), .Z(n28041) );
  NAND U37954 ( .A(n28043), .B(n28044), .Z(c[376]) );
  NAND U37955 ( .A(n26658), .B(o[376]), .Z(n28044) );
  NAND U37956 ( .A(n26653), .B(creg[376]), .Z(n28043) );
  NAND U37957 ( .A(n28045), .B(n28046), .Z(c[375]) );
  NAND U37958 ( .A(n26658), .B(o[375]), .Z(n28046) );
  NAND U37959 ( .A(n26653), .B(creg[375]), .Z(n28045) );
  NAND U37960 ( .A(n28047), .B(n28048), .Z(c[374]) );
  NAND U37961 ( .A(n26658), .B(o[374]), .Z(n28048) );
  NAND U37962 ( .A(n26653), .B(creg[374]), .Z(n28047) );
  NAND U37963 ( .A(n28049), .B(n28050), .Z(c[373]) );
  NAND U37964 ( .A(n26658), .B(o[373]), .Z(n28050) );
  NAND U37965 ( .A(n26653), .B(creg[373]), .Z(n28049) );
  NAND U37966 ( .A(n28051), .B(n28052), .Z(c[372]) );
  NAND U37967 ( .A(n26658), .B(o[372]), .Z(n28052) );
  NAND U37968 ( .A(n26653), .B(creg[372]), .Z(n28051) );
  NAND U37969 ( .A(n28053), .B(n28054), .Z(c[371]) );
  NAND U37970 ( .A(n26658), .B(o[371]), .Z(n28054) );
  NAND U37971 ( .A(n26653), .B(creg[371]), .Z(n28053) );
  NAND U37972 ( .A(n28055), .B(n28056), .Z(c[370]) );
  NAND U37973 ( .A(n26658), .B(o[370]), .Z(n28056) );
  NAND U37974 ( .A(n26653), .B(creg[370]), .Z(n28055) );
  NAND U37975 ( .A(n28057), .B(n28058), .Z(c[36]) );
  NAND U37976 ( .A(n26658), .B(o[36]), .Z(n28058) );
  NAND U37977 ( .A(n26653), .B(creg[36]), .Z(n28057) );
  NAND U37978 ( .A(n28059), .B(n28060), .Z(c[369]) );
  NAND U37979 ( .A(n26658), .B(o[369]), .Z(n28060) );
  NAND U37980 ( .A(n26653), .B(creg[369]), .Z(n28059) );
  NAND U37981 ( .A(n28061), .B(n28062), .Z(c[368]) );
  NAND U37982 ( .A(n26658), .B(o[368]), .Z(n28062) );
  NAND U37983 ( .A(n26653), .B(creg[368]), .Z(n28061) );
  NAND U37984 ( .A(n28063), .B(n28064), .Z(c[367]) );
  NAND U37985 ( .A(n26658), .B(o[367]), .Z(n28064) );
  NAND U37986 ( .A(n26653), .B(creg[367]), .Z(n28063) );
  NAND U37987 ( .A(n28065), .B(n28066), .Z(c[366]) );
  NAND U37988 ( .A(n26658), .B(o[366]), .Z(n28066) );
  NAND U37989 ( .A(n26653), .B(creg[366]), .Z(n28065) );
  NAND U37990 ( .A(n28067), .B(n28068), .Z(c[365]) );
  NAND U37991 ( .A(n26658), .B(o[365]), .Z(n28068) );
  NAND U37992 ( .A(n26653), .B(creg[365]), .Z(n28067) );
  NAND U37993 ( .A(n28069), .B(n28070), .Z(c[364]) );
  NAND U37994 ( .A(n26658), .B(o[364]), .Z(n28070) );
  NAND U37995 ( .A(n26653), .B(creg[364]), .Z(n28069) );
  NAND U37996 ( .A(n28071), .B(n28072), .Z(c[363]) );
  NAND U37997 ( .A(n26658), .B(o[363]), .Z(n28072) );
  NAND U37998 ( .A(n26653), .B(creg[363]), .Z(n28071) );
  NAND U37999 ( .A(n28073), .B(n28074), .Z(c[362]) );
  NAND U38000 ( .A(n26658), .B(o[362]), .Z(n28074) );
  NAND U38001 ( .A(n26653), .B(creg[362]), .Z(n28073) );
  NAND U38002 ( .A(n28075), .B(n28076), .Z(c[361]) );
  NAND U38003 ( .A(n26658), .B(o[361]), .Z(n28076) );
  NAND U38004 ( .A(n26653), .B(creg[361]), .Z(n28075) );
  NAND U38005 ( .A(n28077), .B(n28078), .Z(c[360]) );
  NAND U38006 ( .A(n26658), .B(o[360]), .Z(n28078) );
  NAND U38007 ( .A(n26653), .B(creg[360]), .Z(n28077) );
  NAND U38008 ( .A(n28079), .B(n28080), .Z(c[35]) );
  NAND U38009 ( .A(n26658), .B(o[35]), .Z(n28080) );
  NAND U38010 ( .A(n26653), .B(creg[35]), .Z(n28079) );
  NAND U38011 ( .A(n28081), .B(n28082), .Z(c[359]) );
  NAND U38012 ( .A(n26658), .B(o[359]), .Z(n28082) );
  NAND U38013 ( .A(n26653), .B(creg[359]), .Z(n28081) );
  NAND U38014 ( .A(n28083), .B(n28084), .Z(c[358]) );
  NAND U38015 ( .A(n26658), .B(o[358]), .Z(n28084) );
  NAND U38016 ( .A(n26653), .B(creg[358]), .Z(n28083) );
  NAND U38017 ( .A(n28085), .B(n28086), .Z(c[357]) );
  NAND U38018 ( .A(n26658), .B(o[357]), .Z(n28086) );
  NAND U38019 ( .A(n26653), .B(creg[357]), .Z(n28085) );
  NAND U38020 ( .A(n28087), .B(n28088), .Z(c[356]) );
  NAND U38021 ( .A(n26658), .B(o[356]), .Z(n28088) );
  NAND U38022 ( .A(n26653), .B(creg[356]), .Z(n28087) );
  NAND U38023 ( .A(n28089), .B(n28090), .Z(c[355]) );
  NAND U38024 ( .A(n26658), .B(o[355]), .Z(n28090) );
  NAND U38025 ( .A(n26653), .B(creg[355]), .Z(n28089) );
  NAND U38026 ( .A(n28091), .B(n28092), .Z(c[354]) );
  NAND U38027 ( .A(n26658), .B(o[354]), .Z(n28092) );
  NAND U38028 ( .A(n26653), .B(creg[354]), .Z(n28091) );
  NAND U38029 ( .A(n28093), .B(n28094), .Z(c[353]) );
  NAND U38030 ( .A(n26658), .B(o[353]), .Z(n28094) );
  NAND U38031 ( .A(n26653), .B(creg[353]), .Z(n28093) );
  NAND U38032 ( .A(n28095), .B(n28096), .Z(c[352]) );
  NAND U38033 ( .A(n26658), .B(o[352]), .Z(n28096) );
  NAND U38034 ( .A(n26653), .B(creg[352]), .Z(n28095) );
  NAND U38035 ( .A(n28097), .B(n28098), .Z(c[351]) );
  NAND U38036 ( .A(n26658), .B(o[351]), .Z(n28098) );
  NAND U38037 ( .A(n26653), .B(creg[351]), .Z(n28097) );
  NAND U38038 ( .A(n28099), .B(n28100), .Z(c[350]) );
  NAND U38039 ( .A(n26658), .B(o[350]), .Z(n28100) );
  NAND U38040 ( .A(n26653), .B(creg[350]), .Z(n28099) );
  NAND U38041 ( .A(n28101), .B(n28102), .Z(c[34]) );
  NAND U38042 ( .A(n26658), .B(o[34]), .Z(n28102) );
  NAND U38043 ( .A(n26653), .B(creg[34]), .Z(n28101) );
  NAND U38044 ( .A(n28103), .B(n28104), .Z(c[349]) );
  NAND U38045 ( .A(n26658), .B(o[349]), .Z(n28104) );
  NAND U38046 ( .A(n26653), .B(creg[349]), .Z(n28103) );
  NAND U38047 ( .A(n28105), .B(n28106), .Z(c[348]) );
  NAND U38048 ( .A(n26658), .B(o[348]), .Z(n28106) );
  NAND U38049 ( .A(n26653), .B(creg[348]), .Z(n28105) );
  NAND U38050 ( .A(n28107), .B(n28108), .Z(c[347]) );
  NAND U38051 ( .A(n26658), .B(o[347]), .Z(n28108) );
  NAND U38052 ( .A(n26653), .B(creg[347]), .Z(n28107) );
  NAND U38053 ( .A(n28109), .B(n28110), .Z(c[346]) );
  NAND U38054 ( .A(n26658), .B(o[346]), .Z(n28110) );
  NAND U38055 ( .A(n26653), .B(creg[346]), .Z(n28109) );
  NAND U38056 ( .A(n28111), .B(n28112), .Z(c[345]) );
  NAND U38057 ( .A(n26658), .B(o[345]), .Z(n28112) );
  NAND U38058 ( .A(n26653), .B(creg[345]), .Z(n28111) );
  NAND U38059 ( .A(n28113), .B(n28114), .Z(c[344]) );
  NAND U38060 ( .A(n26658), .B(o[344]), .Z(n28114) );
  NAND U38061 ( .A(n26653), .B(creg[344]), .Z(n28113) );
  NAND U38062 ( .A(n28115), .B(n28116), .Z(c[343]) );
  NAND U38063 ( .A(n26658), .B(o[343]), .Z(n28116) );
  NAND U38064 ( .A(n26653), .B(creg[343]), .Z(n28115) );
  NAND U38065 ( .A(n28117), .B(n28118), .Z(c[342]) );
  NAND U38066 ( .A(n26658), .B(o[342]), .Z(n28118) );
  NAND U38067 ( .A(n26653), .B(creg[342]), .Z(n28117) );
  NAND U38068 ( .A(n28119), .B(n28120), .Z(c[341]) );
  NAND U38069 ( .A(n26658), .B(o[341]), .Z(n28120) );
  NAND U38070 ( .A(n26653), .B(creg[341]), .Z(n28119) );
  NAND U38071 ( .A(n28121), .B(n28122), .Z(c[340]) );
  NAND U38072 ( .A(n26658), .B(o[340]), .Z(n28122) );
  NAND U38073 ( .A(n26653), .B(creg[340]), .Z(n28121) );
  NAND U38074 ( .A(n28123), .B(n28124), .Z(c[33]) );
  NAND U38075 ( .A(n26658), .B(o[33]), .Z(n28124) );
  NAND U38076 ( .A(n26653), .B(creg[33]), .Z(n28123) );
  NAND U38077 ( .A(n28125), .B(n28126), .Z(c[339]) );
  NAND U38078 ( .A(n26658), .B(o[339]), .Z(n28126) );
  NAND U38079 ( .A(n26653), .B(creg[339]), .Z(n28125) );
  NAND U38080 ( .A(n28127), .B(n28128), .Z(c[338]) );
  NAND U38081 ( .A(n26658), .B(o[338]), .Z(n28128) );
  NAND U38082 ( .A(n26653), .B(creg[338]), .Z(n28127) );
  NAND U38083 ( .A(n28129), .B(n28130), .Z(c[337]) );
  NAND U38084 ( .A(n26658), .B(o[337]), .Z(n28130) );
  NAND U38085 ( .A(n26653), .B(creg[337]), .Z(n28129) );
  NAND U38086 ( .A(n28131), .B(n28132), .Z(c[336]) );
  NAND U38087 ( .A(n26658), .B(o[336]), .Z(n28132) );
  NAND U38088 ( .A(n26653), .B(creg[336]), .Z(n28131) );
  NAND U38089 ( .A(n28133), .B(n28134), .Z(c[335]) );
  NAND U38090 ( .A(n26658), .B(o[335]), .Z(n28134) );
  NAND U38091 ( .A(n26653), .B(creg[335]), .Z(n28133) );
  NAND U38092 ( .A(n28135), .B(n28136), .Z(c[334]) );
  NAND U38093 ( .A(n26658), .B(o[334]), .Z(n28136) );
  NAND U38094 ( .A(n26653), .B(creg[334]), .Z(n28135) );
  NAND U38095 ( .A(n28137), .B(n28138), .Z(c[333]) );
  NAND U38096 ( .A(n26658), .B(o[333]), .Z(n28138) );
  NAND U38097 ( .A(n26653), .B(creg[333]), .Z(n28137) );
  NAND U38098 ( .A(n28139), .B(n28140), .Z(c[332]) );
  NAND U38099 ( .A(n26658), .B(o[332]), .Z(n28140) );
  NAND U38100 ( .A(n26653), .B(creg[332]), .Z(n28139) );
  NAND U38101 ( .A(n28141), .B(n28142), .Z(c[331]) );
  NAND U38102 ( .A(n26658), .B(o[331]), .Z(n28142) );
  NAND U38103 ( .A(n26653), .B(creg[331]), .Z(n28141) );
  NAND U38104 ( .A(n28143), .B(n28144), .Z(c[330]) );
  NAND U38105 ( .A(n26658), .B(o[330]), .Z(n28144) );
  NAND U38106 ( .A(n26653), .B(creg[330]), .Z(n28143) );
  NAND U38107 ( .A(n28145), .B(n28146), .Z(c[32]) );
  NAND U38108 ( .A(n26658), .B(o[32]), .Z(n28146) );
  NAND U38109 ( .A(n26653), .B(creg[32]), .Z(n28145) );
  NAND U38110 ( .A(n28147), .B(n28148), .Z(c[329]) );
  NAND U38111 ( .A(n26658), .B(o[329]), .Z(n28148) );
  NAND U38112 ( .A(n26653), .B(creg[329]), .Z(n28147) );
  NAND U38113 ( .A(n28149), .B(n28150), .Z(c[328]) );
  NAND U38114 ( .A(n26658), .B(o[328]), .Z(n28150) );
  NAND U38115 ( .A(n26653), .B(creg[328]), .Z(n28149) );
  NAND U38116 ( .A(n28151), .B(n28152), .Z(c[327]) );
  NAND U38117 ( .A(n26658), .B(o[327]), .Z(n28152) );
  NAND U38118 ( .A(n26653), .B(creg[327]), .Z(n28151) );
  NAND U38119 ( .A(n28153), .B(n28154), .Z(c[326]) );
  NAND U38120 ( .A(n26658), .B(o[326]), .Z(n28154) );
  NAND U38121 ( .A(n26653), .B(creg[326]), .Z(n28153) );
  NAND U38122 ( .A(n28155), .B(n28156), .Z(c[325]) );
  NAND U38123 ( .A(n26658), .B(o[325]), .Z(n28156) );
  NAND U38124 ( .A(n26653), .B(creg[325]), .Z(n28155) );
  NAND U38125 ( .A(n28157), .B(n28158), .Z(c[324]) );
  NAND U38126 ( .A(n26658), .B(o[324]), .Z(n28158) );
  NAND U38127 ( .A(n26653), .B(creg[324]), .Z(n28157) );
  NAND U38128 ( .A(n28159), .B(n28160), .Z(c[323]) );
  NAND U38129 ( .A(n26658), .B(o[323]), .Z(n28160) );
  NAND U38130 ( .A(n26653), .B(creg[323]), .Z(n28159) );
  NAND U38131 ( .A(n28161), .B(n28162), .Z(c[322]) );
  NAND U38132 ( .A(n26658), .B(o[322]), .Z(n28162) );
  NAND U38133 ( .A(n26653), .B(creg[322]), .Z(n28161) );
  NAND U38134 ( .A(n28163), .B(n28164), .Z(c[321]) );
  NAND U38135 ( .A(n26658), .B(o[321]), .Z(n28164) );
  NAND U38136 ( .A(n26653), .B(creg[321]), .Z(n28163) );
  NAND U38137 ( .A(n28165), .B(n28166), .Z(c[320]) );
  NAND U38138 ( .A(n26658), .B(o[320]), .Z(n28166) );
  NAND U38139 ( .A(n26653), .B(creg[320]), .Z(n28165) );
  NAND U38140 ( .A(n28167), .B(n28168), .Z(c[31]) );
  NAND U38141 ( .A(n26658), .B(o[31]), .Z(n28168) );
  NAND U38142 ( .A(n26653), .B(creg[31]), .Z(n28167) );
  NAND U38143 ( .A(n28169), .B(n28170), .Z(c[319]) );
  NAND U38144 ( .A(n26658), .B(o[319]), .Z(n28170) );
  NAND U38145 ( .A(n26653), .B(creg[319]), .Z(n28169) );
  NAND U38146 ( .A(n28171), .B(n28172), .Z(c[318]) );
  NAND U38147 ( .A(n26658), .B(o[318]), .Z(n28172) );
  NAND U38148 ( .A(n26653), .B(creg[318]), .Z(n28171) );
  NAND U38149 ( .A(n28173), .B(n28174), .Z(c[317]) );
  NAND U38150 ( .A(n26658), .B(o[317]), .Z(n28174) );
  NAND U38151 ( .A(n26653), .B(creg[317]), .Z(n28173) );
  NAND U38152 ( .A(n28175), .B(n28176), .Z(c[316]) );
  NAND U38153 ( .A(n26658), .B(o[316]), .Z(n28176) );
  NAND U38154 ( .A(n26653), .B(creg[316]), .Z(n28175) );
  NAND U38155 ( .A(n28177), .B(n28178), .Z(c[315]) );
  NAND U38156 ( .A(n26658), .B(o[315]), .Z(n28178) );
  NAND U38157 ( .A(n26653), .B(creg[315]), .Z(n28177) );
  NAND U38158 ( .A(n28179), .B(n28180), .Z(c[314]) );
  NAND U38159 ( .A(n26658), .B(o[314]), .Z(n28180) );
  NAND U38160 ( .A(n26653), .B(creg[314]), .Z(n28179) );
  NAND U38161 ( .A(n28181), .B(n28182), .Z(c[313]) );
  NAND U38162 ( .A(n26658), .B(o[313]), .Z(n28182) );
  NAND U38163 ( .A(n26653), .B(creg[313]), .Z(n28181) );
  NAND U38164 ( .A(n28183), .B(n28184), .Z(c[312]) );
  NAND U38165 ( .A(n26658), .B(o[312]), .Z(n28184) );
  NAND U38166 ( .A(n26653), .B(creg[312]), .Z(n28183) );
  NAND U38167 ( .A(n28185), .B(n28186), .Z(c[311]) );
  NAND U38168 ( .A(n26658), .B(o[311]), .Z(n28186) );
  NAND U38169 ( .A(n26653), .B(creg[311]), .Z(n28185) );
  NAND U38170 ( .A(n28187), .B(n28188), .Z(c[310]) );
  NAND U38171 ( .A(n26658), .B(o[310]), .Z(n28188) );
  NAND U38172 ( .A(n26653), .B(creg[310]), .Z(n28187) );
  NAND U38173 ( .A(n28189), .B(n28190), .Z(c[30]) );
  NAND U38174 ( .A(n26658), .B(o[30]), .Z(n28190) );
  NAND U38175 ( .A(n26653), .B(creg[30]), .Z(n28189) );
  NAND U38176 ( .A(n28191), .B(n28192), .Z(c[309]) );
  NAND U38177 ( .A(n26658), .B(o[309]), .Z(n28192) );
  NAND U38178 ( .A(n26653), .B(creg[309]), .Z(n28191) );
  NAND U38179 ( .A(n28193), .B(n28194), .Z(c[308]) );
  NAND U38180 ( .A(n26658), .B(o[308]), .Z(n28194) );
  NAND U38181 ( .A(n26653), .B(creg[308]), .Z(n28193) );
  NAND U38182 ( .A(n28195), .B(n28196), .Z(c[307]) );
  NAND U38183 ( .A(n26658), .B(o[307]), .Z(n28196) );
  NAND U38184 ( .A(n26653), .B(creg[307]), .Z(n28195) );
  NAND U38185 ( .A(n28197), .B(n28198), .Z(c[306]) );
  NAND U38186 ( .A(n26658), .B(o[306]), .Z(n28198) );
  NAND U38187 ( .A(n26653), .B(creg[306]), .Z(n28197) );
  NAND U38188 ( .A(n28199), .B(n28200), .Z(c[305]) );
  NAND U38189 ( .A(n26658), .B(o[305]), .Z(n28200) );
  NAND U38190 ( .A(n26653), .B(creg[305]), .Z(n28199) );
  NAND U38191 ( .A(n28201), .B(n28202), .Z(c[304]) );
  NAND U38192 ( .A(n26658), .B(o[304]), .Z(n28202) );
  NAND U38193 ( .A(n26653), .B(creg[304]), .Z(n28201) );
  NAND U38194 ( .A(n28203), .B(n28204), .Z(c[303]) );
  NAND U38195 ( .A(n26658), .B(o[303]), .Z(n28204) );
  NAND U38196 ( .A(n26653), .B(creg[303]), .Z(n28203) );
  NAND U38197 ( .A(n28205), .B(n28206), .Z(c[302]) );
  NAND U38198 ( .A(n26658), .B(o[302]), .Z(n28206) );
  NAND U38199 ( .A(n26653), .B(creg[302]), .Z(n28205) );
  NAND U38200 ( .A(n28207), .B(n28208), .Z(c[301]) );
  NAND U38201 ( .A(n26658), .B(o[301]), .Z(n28208) );
  NAND U38202 ( .A(n26653), .B(creg[301]), .Z(n28207) );
  NAND U38203 ( .A(n28209), .B(n28210), .Z(c[300]) );
  NAND U38204 ( .A(n26658), .B(o[300]), .Z(n28210) );
  NAND U38205 ( .A(n26653), .B(creg[300]), .Z(n28209) );
  NAND U38206 ( .A(n28211), .B(n28212), .Z(c[2]) );
  NAND U38207 ( .A(n26658), .B(o[2]), .Z(n28212) );
  NAND U38208 ( .A(n26653), .B(creg[2]), .Z(n28211) );
  NAND U38209 ( .A(n28213), .B(n28214), .Z(c[29]) );
  NAND U38210 ( .A(n26658), .B(o[29]), .Z(n28214) );
  NAND U38211 ( .A(n26653), .B(creg[29]), .Z(n28213) );
  NAND U38212 ( .A(n28215), .B(n28216), .Z(c[299]) );
  NAND U38213 ( .A(n26658), .B(o[299]), .Z(n28216) );
  NAND U38214 ( .A(n26653), .B(creg[299]), .Z(n28215) );
  NAND U38215 ( .A(n28217), .B(n28218), .Z(c[298]) );
  NAND U38216 ( .A(n26658), .B(o[298]), .Z(n28218) );
  NAND U38217 ( .A(n26653), .B(creg[298]), .Z(n28217) );
  NAND U38218 ( .A(n28219), .B(n28220), .Z(c[297]) );
  NAND U38219 ( .A(n26658), .B(o[297]), .Z(n28220) );
  NAND U38220 ( .A(n26653), .B(creg[297]), .Z(n28219) );
  NAND U38221 ( .A(n28221), .B(n28222), .Z(c[296]) );
  NAND U38222 ( .A(n26658), .B(o[296]), .Z(n28222) );
  NAND U38223 ( .A(n26653), .B(creg[296]), .Z(n28221) );
  NAND U38224 ( .A(n28223), .B(n28224), .Z(c[295]) );
  NAND U38225 ( .A(n26658), .B(o[295]), .Z(n28224) );
  NAND U38226 ( .A(n26653), .B(creg[295]), .Z(n28223) );
  NAND U38227 ( .A(n28225), .B(n28226), .Z(c[294]) );
  NAND U38228 ( .A(n26658), .B(o[294]), .Z(n28226) );
  NAND U38229 ( .A(n26653), .B(creg[294]), .Z(n28225) );
  NAND U38230 ( .A(n28227), .B(n28228), .Z(c[293]) );
  NAND U38231 ( .A(n26658), .B(o[293]), .Z(n28228) );
  NAND U38232 ( .A(n26653), .B(creg[293]), .Z(n28227) );
  NAND U38233 ( .A(n28229), .B(n28230), .Z(c[292]) );
  NAND U38234 ( .A(n26658), .B(o[292]), .Z(n28230) );
  NAND U38235 ( .A(n26653), .B(creg[292]), .Z(n28229) );
  NAND U38236 ( .A(n28231), .B(n28232), .Z(c[291]) );
  NAND U38237 ( .A(n26658), .B(o[291]), .Z(n28232) );
  NAND U38238 ( .A(n26653), .B(creg[291]), .Z(n28231) );
  NAND U38239 ( .A(n28233), .B(n28234), .Z(c[290]) );
  NAND U38240 ( .A(n26658), .B(o[290]), .Z(n28234) );
  NAND U38241 ( .A(n26653), .B(creg[290]), .Z(n28233) );
  NAND U38242 ( .A(n28235), .B(n28236), .Z(c[28]) );
  NAND U38243 ( .A(n26658), .B(o[28]), .Z(n28236) );
  NAND U38244 ( .A(n26653), .B(creg[28]), .Z(n28235) );
  NAND U38245 ( .A(n28237), .B(n28238), .Z(c[289]) );
  NAND U38246 ( .A(n26658), .B(o[289]), .Z(n28238) );
  NAND U38247 ( .A(n26653), .B(creg[289]), .Z(n28237) );
  NAND U38248 ( .A(n28239), .B(n28240), .Z(c[288]) );
  NAND U38249 ( .A(n26658), .B(o[288]), .Z(n28240) );
  NAND U38250 ( .A(n26653), .B(creg[288]), .Z(n28239) );
  NAND U38251 ( .A(n28241), .B(n28242), .Z(c[287]) );
  NAND U38252 ( .A(n26658), .B(o[287]), .Z(n28242) );
  NAND U38253 ( .A(n26653), .B(creg[287]), .Z(n28241) );
  NAND U38254 ( .A(n28243), .B(n28244), .Z(c[286]) );
  NAND U38255 ( .A(n26658), .B(o[286]), .Z(n28244) );
  NAND U38256 ( .A(n26653), .B(creg[286]), .Z(n28243) );
  NAND U38257 ( .A(n28245), .B(n28246), .Z(c[285]) );
  NAND U38258 ( .A(n26658), .B(o[285]), .Z(n28246) );
  NAND U38259 ( .A(n26653), .B(creg[285]), .Z(n28245) );
  NAND U38260 ( .A(n28247), .B(n28248), .Z(c[284]) );
  NAND U38261 ( .A(n26658), .B(o[284]), .Z(n28248) );
  NAND U38262 ( .A(n26653), .B(creg[284]), .Z(n28247) );
  NAND U38263 ( .A(n28249), .B(n28250), .Z(c[283]) );
  NAND U38264 ( .A(n26658), .B(o[283]), .Z(n28250) );
  NAND U38265 ( .A(n26653), .B(creg[283]), .Z(n28249) );
  NAND U38266 ( .A(n28251), .B(n28252), .Z(c[282]) );
  NAND U38267 ( .A(n26658), .B(o[282]), .Z(n28252) );
  NAND U38268 ( .A(n26653), .B(creg[282]), .Z(n28251) );
  NAND U38269 ( .A(n28253), .B(n28254), .Z(c[281]) );
  NAND U38270 ( .A(n26658), .B(o[281]), .Z(n28254) );
  NAND U38271 ( .A(n26653), .B(creg[281]), .Z(n28253) );
  NAND U38272 ( .A(n28255), .B(n28256), .Z(c[280]) );
  NAND U38273 ( .A(n26658), .B(o[280]), .Z(n28256) );
  NAND U38274 ( .A(n26653), .B(creg[280]), .Z(n28255) );
  NAND U38275 ( .A(n28257), .B(n28258), .Z(c[27]) );
  NAND U38276 ( .A(n26658), .B(o[27]), .Z(n28258) );
  NAND U38277 ( .A(n26653), .B(creg[27]), .Z(n28257) );
  NAND U38278 ( .A(n28259), .B(n28260), .Z(c[279]) );
  NAND U38279 ( .A(n26658), .B(o[279]), .Z(n28260) );
  NAND U38280 ( .A(n26653), .B(creg[279]), .Z(n28259) );
  NAND U38281 ( .A(n28261), .B(n28262), .Z(c[278]) );
  NAND U38282 ( .A(n26658), .B(o[278]), .Z(n28262) );
  NAND U38283 ( .A(n26653), .B(creg[278]), .Z(n28261) );
  NAND U38284 ( .A(n28263), .B(n28264), .Z(c[277]) );
  NAND U38285 ( .A(n26658), .B(o[277]), .Z(n28264) );
  NAND U38286 ( .A(n26653), .B(creg[277]), .Z(n28263) );
  NAND U38287 ( .A(n28265), .B(n28266), .Z(c[276]) );
  NAND U38288 ( .A(n26658), .B(o[276]), .Z(n28266) );
  NAND U38289 ( .A(n26653), .B(creg[276]), .Z(n28265) );
  NAND U38290 ( .A(n28267), .B(n28268), .Z(c[275]) );
  NAND U38291 ( .A(n26658), .B(o[275]), .Z(n28268) );
  NAND U38292 ( .A(n26653), .B(creg[275]), .Z(n28267) );
  NAND U38293 ( .A(n28269), .B(n28270), .Z(c[274]) );
  NAND U38294 ( .A(n26658), .B(o[274]), .Z(n28270) );
  NAND U38295 ( .A(n26653), .B(creg[274]), .Z(n28269) );
  NAND U38296 ( .A(n28271), .B(n28272), .Z(c[273]) );
  NAND U38297 ( .A(n26658), .B(o[273]), .Z(n28272) );
  NAND U38298 ( .A(n26653), .B(creg[273]), .Z(n28271) );
  NAND U38299 ( .A(n28273), .B(n28274), .Z(c[272]) );
  NAND U38300 ( .A(n26658), .B(o[272]), .Z(n28274) );
  NAND U38301 ( .A(n26653), .B(creg[272]), .Z(n28273) );
  NAND U38302 ( .A(n28275), .B(n28276), .Z(c[271]) );
  NAND U38303 ( .A(n26658), .B(o[271]), .Z(n28276) );
  NAND U38304 ( .A(n26653), .B(creg[271]), .Z(n28275) );
  NAND U38305 ( .A(n28277), .B(n28278), .Z(c[270]) );
  NAND U38306 ( .A(n26658), .B(o[270]), .Z(n28278) );
  NAND U38307 ( .A(n26653), .B(creg[270]), .Z(n28277) );
  NAND U38308 ( .A(n28279), .B(n28280), .Z(c[26]) );
  NAND U38309 ( .A(n26658), .B(o[26]), .Z(n28280) );
  NAND U38310 ( .A(n26653), .B(creg[26]), .Z(n28279) );
  NAND U38311 ( .A(n28281), .B(n28282), .Z(c[269]) );
  NAND U38312 ( .A(n26658), .B(o[269]), .Z(n28282) );
  NAND U38313 ( .A(n26653), .B(creg[269]), .Z(n28281) );
  NAND U38314 ( .A(n28283), .B(n28284), .Z(c[268]) );
  NAND U38315 ( .A(n26658), .B(o[268]), .Z(n28284) );
  NAND U38316 ( .A(n26653), .B(creg[268]), .Z(n28283) );
  NAND U38317 ( .A(n28285), .B(n28286), .Z(c[267]) );
  NAND U38318 ( .A(n26658), .B(o[267]), .Z(n28286) );
  NAND U38319 ( .A(n26653), .B(creg[267]), .Z(n28285) );
  NAND U38320 ( .A(n28287), .B(n28288), .Z(c[266]) );
  NAND U38321 ( .A(n26658), .B(o[266]), .Z(n28288) );
  NAND U38322 ( .A(n26653), .B(creg[266]), .Z(n28287) );
  NAND U38323 ( .A(n28289), .B(n28290), .Z(c[265]) );
  NAND U38324 ( .A(n26658), .B(o[265]), .Z(n28290) );
  NAND U38325 ( .A(n26653), .B(creg[265]), .Z(n28289) );
  NAND U38326 ( .A(n28291), .B(n28292), .Z(c[264]) );
  NAND U38327 ( .A(n26658), .B(o[264]), .Z(n28292) );
  NAND U38328 ( .A(n26653), .B(creg[264]), .Z(n28291) );
  NAND U38329 ( .A(n28293), .B(n28294), .Z(c[263]) );
  NAND U38330 ( .A(n26658), .B(o[263]), .Z(n28294) );
  NAND U38331 ( .A(n26653), .B(creg[263]), .Z(n28293) );
  NAND U38332 ( .A(n28295), .B(n28296), .Z(c[262]) );
  NAND U38333 ( .A(n26658), .B(o[262]), .Z(n28296) );
  NAND U38334 ( .A(n26653), .B(creg[262]), .Z(n28295) );
  NAND U38335 ( .A(n28297), .B(n28298), .Z(c[261]) );
  NAND U38336 ( .A(n26658), .B(o[261]), .Z(n28298) );
  NAND U38337 ( .A(n26653), .B(creg[261]), .Z(n28297) );
  NAND U38338 ( .A(n28299), .B(n28300), .Z(c[260]) );
  NAND U38339 ( .A(n26658), .B(o[260]), .Z(n28300) );
  NAND U38340 ( .A(n26653), .B(creg[260]), .Z(n28299) );
  NAND U38341 ( .A(n28301), .B(n28302), .Z(c[25]) );
  NAND U38342 ( .A(n26658), .B(o[25]), .Z(n28302) );
  NAND U38343 ( .A(n26653), .B(creg[25]), .Z(n28301) );
  NAND U38344 ( .A(n28303), .B(n28304), .Z(c[259]) );
  NAND U38345 ( .A(n26658), .B(o[259]), .Z(n28304) );
  NAND U38346 ( .A(n26653), .B(creg[259]), .Z(n28303) );
  NAND U38347 ( .A(n28305), .B(n28306), .Z(c[258]) );
  NAND U38348 ( .A(n26658), .B(o[258]), .Z(n28306) );
  NAND U38349 ( .A(n26653), .B(creg[258]), .Z(n28305) );
  NAND U38350 ( .A(n28307), .B(n28308), .Z(c[257]) );
  NAND U38351 ( .A(n26658), .B(o[257]), .Z(n28308) );
  NAND U38352 ( .A(n26653), .B(creg[257]), .Z(n28307) );
  NAND U38353 ( .A(n28309), .B(n28310), .Z(c[256]) );
  NAND U38354 ( .A(n26658), .B(o[256]), .Z(n28310) );
  NAND U38355 ( .A(n26653), .B(creg[256]), .Z(n28309) );
  NAND U38356 ( .A(n28311), .B(n28312), .Z(c[255]) );
  NAND U38357 ( .A(n26658), .B(o[255]), .Z(n28312) );
  NAND U38358 ( .A(n26653), .B(creg[255]), .Z(n28311) );
  NAND U38359 ( .A(n28313), .B(n28314), .Z(c[254]) );
  NAND U38360 ( .A(n26658), .B(o[254]), .Z(n28314) );
  NAND U38361 ( .A(n26653), .B(creg[254]), .Z(n28313) );
  NAND U38362 ( .A(n28315), .B(n28316), .Z(c[253]) );
  NAND U38363 ( .A(n26658), .B(o[253]), .Z(n28316) );
  NAND U38364 ( .A(n26653), .B(creg[253]), .Z(n28315) );
  NAND U38365 ( .A(n28317), .B(n28318), .Z(c[252]) );
  NAND U38366 ( .A(n26658), .B(o[252]), .Z(n28318) );
  NAND U38367 ( .A(n26653), .B(creg[252]), .Z(n28317) );
  NAND U38368 ( .A(n28319), .B(n28320), .Z(c[251]) );
  NAND U38369 ( .A(n26658), .B(o[251]), .Z(n28320) );
  NAND U38370 ( .A(n26653), .B(creg[251]), .Z(n28319) );
  NAND U38371 ( .A(n28321), .B(n28322), .Z(c[250]) );
  NAND U38372 ( .A(n26658), .B(o[250]), .Z(n28322) );
  NAND U38373 ( .A(n26653), .B(creg[250]), .Z(n28321) );
  NAND U38374 ( .A(n28323), .B(n28324), .Z(c[24]) );
  NAND U38375 ( .A(n26658), .B(o[24]), .Z(n28324) );
  NAND U38376 ( .A(n26653), .B(creg[24]), .Z(n28323) );
  NAND U38377 ( .A(n28325), .B(n28326), .Z(c[249]) );
  NAND U38378 ( .A(n26658), .B(o[249]), .Z(n28326) );
  NAND U38379 ( .A(n26653), .B(creg[249]), .Z(n28325) );
  NAND U38380 ( .A(n28327), .B(n28328), .Z(c[248]) );
  NAND U38381 ( .A(n26658), .B(o[248]), .Z(n28328) );
  NAND U38382 ( .A(n26653), .B(creg[248]), .Z(n28327) );
  NAND U38383 ( .A(n28329), .B(n28330), .Z(c[247]) );
  NAND U38384 ( .A(n26658), .B(o[247]), .Z(n28330) );
  NAND U38385 ( .A(n26653), .B(creg[247]), .Z(n28329) );
  NAND U38386 ( .A(n28331), .B(n28332), .Z(c[246]) );
  NAND U38387 ( .A(n26658), .B(o[246]), .Z(n28332) );
  NAND U38388 ( .A(n26653), .B(creg[246]), .Z(n28331) );
  NAND U38389 ( .A(n28333), .B(n28334), .Z(c[245]) );
  NAND U38390 ( .A(n26658), .B(o[245]), .Z(n28334) );
  NAND U38391 ( .A(n26653), .B(creg[245]), .Z(n28333) );
  NAND U38392 ( .A(n28335), .B(n28336), .Z(c[244]) );
  NAND U38393 ( .A(n26658), .B(o[244]), .Z(n28336) );
  NAND U38394 ( .A(n26653), .B(creg[244]), .Z(n28335) );
  NAND U38395 ( .A(n28337), .B(n28338), .Z(c[243]) );
  NAND U38396 ( .A(n26658), .B(o[243]), .Z(n28338) );
  NAND U38397 ( .A(n26653), .B(creg[243]), .Z(n28337) );
  NAND U38398 ( .A(n28339), .B(n28340), .Z(c[242]) );
  NAND U38399 ( .A(n26658), .B(o[242]), .Z(n28340) );
  NAND U38400 ( .A(n26653), .B(creg[242]), .Z(n28339) );
  NAND U38401 ( .A(n28341), .B(n28342), .Z(c[241]) );
  NAND U38402 ( .A(n26658), .B(o[241]), .Z(n28342) );
  NAND U38403 ( .A(n26653), .B(creg[241]), .Z(n28341) );
  NAND U38404 ( .A(n28343), .B(n28344), .Z(c[240]) );
  NAND U38405 ( .A(n26658), .B(o[240]), .Z(n28344) );
  NAND U38406 ( .A(n26653), .B(creg[240]), .Z(n28343) );
  NAND U38407 ( .A(n28345), .B(n28346), .Z(c[23]) );
  NAND U38408 ( .A(n26658), .B(o[23]), .Z(n28346) );
  NAND U38409 ( .A(n26653), .B(creg[23]), .Z(n28345) );
  NAND U38410 ( .A(n28347), .B(n28348), .Z(c[239]) );
  NAND U38411 ( .A(n26658), .B(o[239]), .Z(n28348) );
  NAND U38412 ( .A(n26653), .B(creg[239]), .Z(n28347) );
  NAND U38413 ( .A(n28349), .B(n28350), .Z(c[238]) );
  NAND U38414 ( .A(n26658), .B(o[238]), .Z(n28350) );
  NAND U38415 ( .A(n26653), .B(creg[238]), .Z(n28349) );
  NAND U38416 ( .A(n28351), .B(n28352), .Z(c[237]) );
  NAND U38417 ( .A(n26658), .B(o[237]), .Z(n28352) );
  NAND U38418 ( .A(n26653), .B(creg[237]), .Z(n28351) );
  NAND U38419 ( .A(n28353), .B(n28354), .Z(c[236]) );
  NAND U38420 ( .A(n26658), .B(o[236]), .Z(n28354) );
  NAND U38421 ( .A(n26653), .B(creg[236]), .Z(n28353) );
  NAND U38422 ( .A(n28355), .B(n28356), .Z(c[235]) );
  NAND U38423 ( .A(n26658), .B(o[235]), .Z(n28356) );
  NAND U38424 ( .A(n26653), .B(creg[235]), .Z(n28355) );
  NAND U38425 ( .A(n28357), .B(n28358), .Z(c[234]) );
  NAND U38426 ( .A(n26658), .B(o[234]), .Z(n28358) );
  NAND U38427 ( .A(n26653), .B(creg[234]), .Z(n28357) );
  NAND U38428 ( .A(n28359), .B(n28360), .Z(c[233]) );
  NAND U38429 ( .A(n26658), .B(o[233]), .Z(n28360) );
  NAND U38430 ( .A(n26653), .B(creg[233]), .Z(n28359) );
  NAND U38431 ( .A(n28361), .B(n28362), .Z(c[232]) );
  NAND U38432 ( .A(n26658), .B(o[232]), .Z(n28362) );
  NAND U38433 ( .A(n26653), .B(creg[232]), .Z(n28361) );
  NAND U38434 ( .A(n28363), .B(n28364), .Z(c[231]) );
  NAND U38435 ( .A(n26658), .B(o[231]), .Z(n28364) );
  NAND U38436 ( .A(n26653), .B(creg[231]), .Z(n28363) );
  NAND U38437 ( .A(n28365), .B(n28366), .Z(c[230]) );
  NAND U38438 ( .A(n26658), .B(o[230]), .Z(n28366) );
  NAND U38439 ( .A(n26653), .B(creg[230]), .Z(n28365) );
  NAND U38440 ( .A(n28367), .B(n28368), .Z(c[22]) );
  NAND U38441 ( .A(n26658), .B(o[22]), .Z(n28368) );
  NAND U38442 ( .A(n26653), .B(creg[22]), .Z(n28367) );
  NAND U38443 ( .A(n28369), .B(n28370), .Z(c[229]) );
  NAND U38444 ( .A(n26658), .B(o[229]), .Z(n28370) );
  NAND U38445 ( .A(n26653), .B(creg[229]), .Z(n28369) );
  NAND U38446 ( .A(n28371), .B(n28372), .Z(c[228]) );
  NAND U38447 ( .A(n26658), .B(o[228]), .Z(n28372) );
  NAND U38448 ( .A(n26653), .B(creg[228]), .Z(n28371) );
  NAND U38449 ( .A(n28373), .B(n28374), .Z(c[227]) );
  NAND U38450 ( .A(n26658), .B(o[227]), .Z(n28374) );
  NAND U38451 ( .A(n26653), .B(creg[227]), .Z(n28373) );
  NAND U38452 ( .A(n28375), .B(n28376), .Z(c[226]) );
  NAND U38453 ( .A(n26658), .B(o[226]), .Z(n28376) );
  NAND U38454 ( .A(n26653), .B(creg[226]), .Z(n28375) );
  NAND U38455 ( .A(n28377), .B(n28378), .Z(c[225]) );
  NAND U38456 ( .A(n26658), .B(o[225]), .Z(n28378) );
  NAND U38457 ( .A(n26653), .B(creg[225]), .Z(n28377) );
  NAND U38458 ( .A(n28379), .B(n28380), .Z(c[224]) );
  NAND U38459 ( .A(n26658), .B(o[224]), .Z(n28380) );
  NAND U38460 ( .A(n26653), .B(creg[224]), .Z(n28379) );
  NAND U38461 ( .A(n28381), .B(n28382), .Z(c[223]) );
  NAND U38462 ( .A(n26658), .B(o[223]), .Z(n28382) );
  NAND U38463 ( .A(n26653), .B(creg[223]), .Z(n28381) );
  NAND U38464 ( .A(n28383), .B(n28384), .Z(c[222]) );
  NAND U38465 ( .A(n26658), .B(o[222]), .Z(n28384) );
  NAND U38466 ( .A(n26653), .B(creg[222]), .Z(n28383) );
  NAND U38467 ( .A(n28385), .B(n28386), .Z(c[221]) );
  NAND U38468 ( .A(n26658), .B(o[221]), .Z(n28386) );
  NAND U38469 ( .A(n26653), .B(creg[221]), .Z(n28385) );
  NAND U38470 ( .A(n28387), .B(n28388), .Z(c[220]) );
  NAND U38471 ( .A(n26658), .B(o[220]), .Z(n28388) );
  NAND U38472 ( .A(n26653), .B(creg[220]), .Z(n28387) );
  NAND U38473 ( .A(n28389), .B(n28390), .Z(c[21]) );
  NAND U38474 ( .A(n26658), .B(o[21]), .Z(n28390) );
  NAND U38475 ( .A(n26653), .B(creg[21]), .Z(n28389) );
  NAND U38476 ( .A(n28391), .B(n28392), .Z(c[219]) );
  NAND U38477 ( .A(n26658), .B(o[219]), .Z(n28392) );
  NAND U38478 ( .A(n26653), .B(creg[219]), .Z(n28391) );
  NAND U38479 ( .A(n28393), .B(n28394), .Z(c[218]) );
  NAND U38480 ( .A(n26658), .B(o[218]), .Z(n28394) );
  NAND U38481 ( .A(n26653), .B(creg[218]), .Z(n28393) );
  NAND U38482 ( .A(n28395), .B(n28396), .Z(c[217]) );
  NAND U38483 ( .A(n26658), .B(o[217]), .Z(n28396) );
  NAND U38484 ( .A(n26653), .B(creg[217]), .Z(n28395) );
  NAND U38485 ( .A(n28397), .B(n28398), .Z(c[216]) );
  NAND U38486 ( .A(n26658), .B(o[216]), .Z(n28398) );
  NAND U38487 ( .A(n26653), .B(creg[216]), .Z(n28397) );
  NAND U38488 ( .A(n28399), .B(n28400), .Z(c[215]) );
  NAND U38489 ( .A(n26658), .B(o[215]), .Z(n28400) );
  NAND U38490 ( .A(n26653), .B(creg[215]), .Z(n28399) );
  NAND U38491 ( .A(n28401), .B(n28402), .Z(c[214]) );
  NAND U38492 ( .A(n26658), .B(o[214]), .Z(n28402) );
  NAND U38493 ( .A(n26653), .B(creg[214]), .Z(n28401) );
  NAND U38494 ( .A(n28403), .B(n28404), .Z(c[213]) );
  NAND U38495 ( .A(n26658), .B(o[213]), .Z(n28404) );
  NAND U38496 ( .A(n26653), .B(creg[213]), .Z(n28403) );
  NAND U38497 ( .A(n28405), .B(n28406), .Z(c[212]) );
  NAND U38498 ( .A(n26658), .B(o[212]), .Z(n28406) );
  NAND U38499 ( .A(n26653), .B(creg[212]), .Z(n28405) );
  NAND U38500 ( .A(n28407), .B(n28408), .Z(c[211]) );
  NAND U38501 ( .A(n26658), .B(o[211]), .Z(n28408) );
  NAND U38502 ( .A(n26653), .B(creg[211]), .Z(n28407) );
  NAND U38503 ( .A(n28409), .B(n28410), .Z(c[210]) );
  NAND U38504 ( .A(n26658), .B(o[210]), .Z(n28410) );
  NAND U38505 ( .A(n26653), .B(creg[210]), .Z(n28409) );
  NAND U38506 ( .A(n28411), .B(n28412), .Z(c[20]) );
  NAND U38507 ( .A(n26658), .B(o[20]), .Z(n28412) );
  NAND U38508 ( .A(n26653), .B(creg[20]), .Z(n28411) );
  NAND U38509 ( .A(n28413), .B(n28414), .Z(c[209]) );
  NAND U38510 ( .A(n26658), .B(o[209]), .Z(n28414) );
  NAND U38511 ( .A(n26653), .B(creg[209]), .Z(n28413) );
  NAND U38512 ( .A(n28415), .B(n28416), .Z(c[208]) );
  NAND U38513 ( .A(n26658), .B(o[208]), .Z(n28416) );
  NAND U38514 ( .A(n26653), .B(creg[208]), .Z(n28415) );
  NAND U38515 ( .A(n28417), .B(n28418), .Z(c[207]) );
  NAND U38516 ( .A(n26658), .B(o[207]), .Z(n28418) );
  NAND U38517 ( .A(n26653), .B(creg[207]), .Z(n28417) );
  NAND U38518 ( .A(n28419), .B(n28420), .Z(c[206]) );
  NAND U38519 ( .A(n26658), .B(o[206]), .Z(n28420) );
  NAND U38520 ( .A(n26653), .B(creg[206]), .Z(n28419) );
  NAND U38521 ( .A(n28421), .B(n28422), .Z(c[205]) );
  NAND U38522 ( .A(n26658), .B(o[205]), .Z(n28422) );
  NAND U38523 ( .A(n26653), .B(creg[205]), .Z(n28421) );
  NAND U38524 ( .A(n28423), .B(n28424), .Z(c[204]) );
  NAND U38525 ( .A(n26658), .B(o[204]), .Z(n28424) );
  NAND U38526 ( .A(n26653), .B(creg[204]), .Z(n28423) );
  NAND U38527 ( .A(n28425), .B(n28426), .Z(c[203]) );
  NAND U38528 ( .A(n26658), .B(o[203]), .Z(n28426) );
  NAND U38529 ( .A(n26653), .B(creg[203]), .Z(n28425) );
  NAND U38530 ( .A(n28427), .B(n28428), .Z(c[202]) );
  NAND U38531 ( .A(n26658), .B(o[202]), .Z(n28428) );
  NAND U38532 ( .A(n26653), .B(creg[202]), .Z(n28427) );
  NAND U38533 ( .A(n28429), .B(n28430), .Z(c[201]) );
  NAND U38534 ( .A(n26658), .B(o[201]), .Z(n28430) );
  NAND U38535 ( .A(n26653), .B(creg[201]), .Z(n28429) );
  NAND U38536 ( .A(n28431), .B(n28432), .Z(c[200]) );
  NAND U38537 ( .A(n26658), .B(o[200]), .Z(n28432) );
  NAND U38538 ( .A(n26653), .B(creg[200]), .Z(n28431) );
  NAND U38539 ( .A(n28433), .B(n28434), .Z(c[1]) );
  NAND U38540 ( .A(n26658), .B(o[1]), .Z(n28434) );
  NAND U38541 ( .A(n26653), .B(creg[1]), .Z(n28433) );
  NAND U38542 ( .A(n28435), .B(n28436), .Z(c[19]) );
  NAND U38543 ( .A(n26658), .B(o[19]), .Z(n28436) );
  NAND U38544 ( .A(n26653), .B(creg[19]), .Z(n28435) );
  NAND U38545 ( .A(n28437), .B(n28438), .Z(c[199]) );
  NAND U38546 ( .A(n26658), .B(o[199]), .Z(n28438) );
  NAND U38547 ( .A(n26653), .B(creg[199]), .Z(n28437) );
  NAND U38548 ( .A(n28439), .B(n28440), .Z(c[198]) );
  NAND U38549 ( .A(n26658), .B(o[198]), .Z(n28440) );
  NAND U38550 ( .A(n26653), .B(creg[198]), .Z(n28439) );
  NAND U38551 ( .A(n28441), .B(n28442), .Z(c[197]) );
  NAND U38552 ( .A(n26658), .B(o[197]), .Z(n28442) );
  NAND U38553 ( .A(n26653), .B(creg[197]), .Z(n28441) );
  NAND U38554 ( .A(n28443), .B(n28444), .Z(c[196]) );
  NAND U38555 ( .A(n26658), .B(o[196]), .Z(n28444) );
  NAND U38556 ( .A(n26653), .B(creg[196]), .Z(n28443) );
  NAND U38557 ( .A(n28445), .B(n28446), .Z(c[195]) );
  NAND U38558 ( .A(n26658), .B(o[195]), .Z(n28446) );
  NAND U38559 ( .A(n26653), .B(creg[195]), .Z(n28445) );
  NAND U38560 ( .A(n28447), .B(n28448), .Z(c[194]) );
  NAND U38561 ( .A(n26658), .B(o[194]), .Z(n28448) );
  NAND U38562 ( .A(n26653), .B(creg[194]), .Z(n28447) );
  NAND U38563 ( .A(n28449), .B(n28450), .Z(c[193]) );
  NAND U38564 ( .A(n26658), .B(o[193]), .Z(n28450) );
  NAND U38565 ( .A(n26653), .B(creg[193]), .Z(n28449) );
  NAND U38566 ( .A(n28451), .B(n28452), .Z(c[192]) );
  NAND U38567 ( .A(n26658), .B(o[192]), .Z(n28452) );
  NAND U38568 ( .A(n26653), .B(creg[192]), .Z(n28451) );
  NAND U38569 ( .A(n28453), .B(n28454), .Z(c[191]) );
  NAND U38570 ( .A(n26658), .B(o[191]), .Z(n28454) );
  NAND U38571 ( .A(n26653), .B(creg[191]), .Z(n28453) );
  NAND U38572 ( .A(n28455), .B(n28456), .Z(c[190]) );
  NAND U38573 ( .A(n26658), .B(o[190]), .Z(n28456) );
  NAND U38574 ( .A(n26653), .B(creg[190]), .Z(n28455) );
  NAND U38575 ( .A(n28457), .B(n28458), .Z(c[18]) );
  NAND U38576 ( .A(n26658), .B(o[18]), .Z(n28458) );
  NAND U38577 ( .A(n26653), .B(creg[18]), .Z(n28457) );
  NAND U38578 ( .A(n28459), .B(n28460), .Z(c[189]) );
  NAND U38579 ( .A(n26658), .B(o[189]), .Z(n28460) );
  NAND U38580 ( .A(n26653), .B(creg[189]), .Z(n28459) );
  NAND U38581 ( .A(n28461), .B(n28462), .Z(c[188]) );
  NAND U38582 ( .A(n26658), .B(o[188]), .Z(n28462) );
  NAND U38583 ( .A(n26653), .B(creg[188]), .Z(n28461) );
  NAND U38584 ( .A(n28463), .B(n28464), .Z(c[187]) );
  NAND U38585 ( .A(n26658), .B(o[187]), .Z(n28464) );
  NAND U38586 ( .A(n26653), .B(creg[187]), .Z(n28463) );
  NAND U38587 ( .A(n28465), .B(n28466), .Z(c[186]) );
  NAND U38588 ( .A(n26658), .B(o[186]), .Z(n28466) );
  NAND U38589 ( .A(n26653), .B(creg[186]), .Z(n28465) );
  NAND U38590 ( .A(n28467), .B(n28468), .Z(c[185]) );
  NAND U38591 ( .A(n26658), .B(o[185]), .Z(n28468) );
  NAND U38592 ( .A(n26653), .B(creg[185]), .Z(n28467) );
  NAND U38593 ( .A(n28469), .B(n28470), .Z(c[184]) );
  NAND U38594 ( .A(n26658), .B(o[184]), .Z(n28470) );
  NAND U38595 ( .A(n26653), .B(creg[184]), .Z(n28469) );
  NAND U38596 ( .A(n28471), .B(n28472), .Z(c[183]) );
  NAND U38597 ( .A(n26658), .B(o[183]), .Z(n28472) );
  NAND U38598 ( .A(n26653), .B(creg[183]), .Z(n28471) );
  NAND U38599 ( .A(n28473), .B(n28474), .Z(c[182]) );
  NAND U38600 ( .A(n26658), .B(o[182]), .Z(n28474) );
  NAND U38601 ( .A(n26653), .B(creg[182]), .Z(n28473) );
  NAND U38602 ( .A(n28475), .B(n28476), .Z(c[181]) );
  NAND U38603 ( .A(n26658), .B(o[181]), .Z(n28476) );
  NAND U38604 ( .A(n26653), .B(creg[181]), .Z(n28475) );
  NAND U38605 ( .A(n28477), .B(n28478), .Z(c[180]) );
  NAND U38606 ( .A(n26658), .B(o[180]), .Z(n28478) );
  NAND U38607 ( .A(n26653), .B(creg[180]), .Z(n28477) );
  NAND U38608 ( .A(n28479), .B(n28480), .Z(c[17]) );
  NAND U38609 ( .A(n26658), .B(o[17]), .Z(n28480) );
  NAND U38610 ( .A(n26653), .B(creg[17]), .Z(n28479) );
  NAND U38611 ( .A(n28481), .B(n28482), .Z(c[179]) );
  NAND U38612 ( .A(n26658), .B(o[179]), .Z(n28482) );
  NAND U38613 ( .A(n26653), .B(creg[179]), .Z(n28481) );
  NAND U38614 ( .A(n28483), .B(n28484), .Z(c[178]) );
  NAND U38615 ( .A(n26658), .B(o[178]), .Z(n28484) );
  NAND U38616 ( .A(n26653), .B(creg[178]), .Z(n28483) );
  NAND U38617 ( .A(n28485), .B(n28486), .Z(c[177]) );
  NAND U38618 ( .A(n26658), .B(o[177]), .Z(n28486) );
  NAND U38619 ( .A(n26653), .B(creg[177]), .Z(n28485) );
  NAND U38620 ( .A(n28487), .B(n28488), .Z(c[176]) );
  NAND U38621 ( .A(n26658), .B(o[176]), .Z(n28488) );
  NAND U38622 ( .A(n26653), .B(creg[176]), .Z(n28487) );
  NAND U38623 ( .A(n28489), .B(n28490), .Z(c[175]) );
  NAND U38624 ( .A(n26658), .B(o[175]), .Z(n28490) );
  NAND U38625 ( .A(n26653), .B(creg[175]), .Z(n28489) );
  NAND U38626 ( .A(n28491), .B(n28492), .Z(c[174]) );
  NAND U38627 ( .A(n26658), .B(o[174]), .Z(n28492) );
  NAND U38628 ( .A(n26653), .B(creg[174]), .Z(n28491) );
  NAND U38629 ( .A(n28493), .B(n28494), .Z(c[173]) );
  NAND U38630 ( .A(n26658), .B(o[173]), .Z(n28494) );
  NAND U38631 ( .A(n26653), .B(creg[173]), .Z(n28493) );
  NAND U38632 ( .A(n28495), .B(n28496), .Z(c[172]) );
  NAND U38633 ( .A(n26658), .B(o[172]), .Z(n28496) );
  NAND U38634 ( .A(n26653), .B(creg[172]), .Z(n28495) );
  NAND U38635 ( .A(n28497), .B(n28498), .Z(c[171]) );
  NAND U38636 ( .A(n26658), .B(o[171]), .Z(n28498) );
  NAND U38637 ( .A(n26653), .B(creg[171]), .Z(n28497) );
  NAND U38638 ( .A(n28499), .B(n28500), .Z(c[170]) );
  NAND U38639 ( .A(n26658), .B(o[170]), .Z(n28500) );
  NAND U38640 ( .A(n26653), .B(creg[170]), .Z(n28499) );
  NAND U38641 ( .A(n28501), .B(n28502), .Z(c[16]) );
  NAND U38642 ( .A(n26658), .B(o[16]), .Z(n28502) );
  NAND U38643 ( .A(n26653), .B(creg[16]), .Z(n28501) );
  NAND U38644 ( .A(n28503), .B(n28504), .Z(c[169]) );
  NAND U38645 ( .A(n26658), .B(o[169]), .Z(n28504) );
  NAND U38646 ( .A(n26653), .B(creg[169]), .Z(n28503) );
  NAND U38647 ( .A(n28505), .B(n28506), .Z(c[168]) );
  NAND U38648 ( .A(n26658), .B(o[168]), .Z(n28506) );
  NAND U38649 ( .A(n26653), .B(creg[168]), .Z(n28505) );
  NAND U38650 ( .A(n28507), .B(n28508), .Z(c[167]) );
  NAND U38651 ( .A(n26658), .B(o[167]), .Z(n28508) );
  NAND U38652 ( .A(n26653), .B(creg[167]), .Z(n28507) );
  NAND U38653 ( .A(n28509), .B(n28510), .Z(c[166]) );
  NAND U38654 ( .A(n26658), .B(o[166]), .Z(n28510) );
  NAND U38655 ( .A(n26653), .B(creg[166]), .Z(n28509) );
  NAND U38656 ( .A(n28511), .B(n28512), .Z(c[165]) );
  NAND U38657 ( .A(n26658), .B(o[165]), .Z(n28512) );
  NAND U38658 ( .A(n26653), .B(creg[165]), .Z(n28511) );
  NAND U38659 ( .A(n28513), .B(n28514), .Z(c[164]) );
  NAND U38660 ( .A(n26658), .B(o[164]), .Z(n28514) );
  NAND U38661 ( .A(n26653), .B(creg[164]), .Z(n28513) );
  NAND U38662 ( .A(n28515), .B(n28516), .Z(c[163]) );
  NAND U38663 ( .A(n26658), .B(o[163]), .Z(n28516) );
  NAND U38664 ( .A(n26653), .B(creg[163]), .Z(n28515) );
  NAND U38665 ( .A(n28517), .B(n28518), .Z(c[162]) );
  NAND U38666 ( .A(n26658), .B(o[162]), .Z(n28518) );
  NAND U38667 ( .A(n26653), .B(creg[162]), .Z(n28517) );
  NAND U38668 ( .A(n28519), .B(n28520), .Z(c[161]) );
  NAND U38669 ( .A(n26658), .B(o[161]), .Z(n28520) );
  NAND U38670 ( .A(n26653), .B(creg[161]), .Z(n28519) );
  NAND U38671 ( .A(n28521), .B(n28522), .Z(c[160]) );
  NAND U38672 ( .A(n26658), .B(o[160]), .Z(n28522) );
  NAND U38673 ( .A(n26653), .B(creg[160]), .Z(n28521) );
  NAND U38674 ( .A(n28523), .B(n28524), .Z(c[15]) );
  NAND U38675 ( .A(n26658), .B(o[15]), .Z(n28524) );
  NAND U38676 ( .A(n26653), .B(creg[15]), .Z(n28523) );
  NAND U38677 ( .A(n28525), .B(n28526), .Z(c[159]) );
  NAND U38678 ( .A(n26658), .B(o[159]), .Z(n28526) );
  NAND U38679 ( .A(n26653), .B(creg[159]), .Z(n28525) );
  NAND U38680 ( .A(n28527), .B(n28528), .Z(c[158]) );
  NAND U38681 ( .A(n26658), .B(o[158]), .Z(n28528) );
  NAND U38682 ( .A(n26653), .B(creg[158]), .Z(n28527) );
  NAND U38683 ( .A(n28529), .B(n28530), .Z(c[157]) );
  NAND U38684 ( .A(n26658), .B(o[157]), .Z(n28530) );
  NAND U38685 ( .A(n26653), .B(creg[157]), .Z(n28529) );
  NAND U38686 ( .A(n28531), .B(n28532), .Z(c[156]) );
  NAND U38687 ( .A(n26658), .B(o[156]), .Z(n28532) );
  NAND U38688 ( .A(n26653), .B(creg[156]), .Z(n28531) );
  NAND U38689 ( .A(n28533), .B(n28534), .Z(c[155]) );
  NAND U38690 ( .A(n26658), .B(o[155]), .Z(n28534) );
  NAND U38691 ( .A(n26653), .B(creg[155]), .Z(n28533) );
  NAND U38692 ( .A(n28535), .B(n28536), .Z(c[154]) );
  NAND U38693 ( .A(n26658), .B(o[154]), .Z(n28536) );
  NAND U38694 ( .A(n26653), .B(creg[154]), .Z(n28535) );
  NAND U38695 ( .A(n28537), .B(n28538), .Z(c[153]) );
  NAND U38696 ( .A(n26658), .B(o[153]), .Z(n28538) );
  NAND U38697 ( .A(n26653), .B(creg[153]), .Z(n28537) );
  NAND U38698 ( .A(n28539), .B(n28540), .Z(c[152]) );
  NAND U38699 ( .A(n26658), .B(o[152]), .Z(n28540) );
  NAND U38700 ( .A(n26653), .B(creg[152]), .Z(n28539) );
  NAND U38701 ( .A(n28541), .B(n28542), .Z(c[151]) );
  NAND U38702 ( .A(n26658), .B(o[151]), .Z(n28542) );
  NAND U38703 ( .A(n26653), .B(creg[151]), .Z(n28541) );
  NAND U38704 ( .A(n28543), .B(n28544), .Z(c[150]) );
  NAND U38705 ( .A(n26658), .B(o[150]), .Z(n28544) );
  NAND U38706 ( .A(n26653), .B(creg[150]), .Z(n28543) );
  NAND U38707 ( .A(n28545), .B(n28546), .Z(c[14]) );
  NAND U38708 ( .A(n26658), .B(o[14]), .Z(n28546) );
  NAND U38709 ( .A(n26653), .B(creg[14]), .Z(n28545) );
  NAND U38710 ( .A(n28547), .B(n28548), .Z(c[149]) );
  NAND U38711 ( .A(n26658), .B(o[149]), .Z(n28548) );
  NAND U38712 ( .A(n26653), .B(creg[149]), .Z(n28547) );
  NAND U38713 ( .A(n28549), .B(n28550), .Z(c[148]) );
  NAND U38714 ( .A(n26658), .B(o[148]), .Z(n28550) );
  NAND U38715 ( .A(n26653), .B(creg[148]), .Z(n28549) );
  NAND U38716 ( .A(n28551), .B(n28552), .Z(c[147]) );
  NAND U38717 ( .A(n26658), .B(o[147]), .Z(n28552) );
  NAND U38718 ( .A(n26653), .B(creg[147]), .Z(n28551) );
  NAND U38719 ( .A(n28553), .B(n28554), .Z(c[146]) );
  NAND U38720 ( .A(n26658), .B(o[146]), .Z(n28554) );
  NAND U38721 ( .A(n26653), .B(creg[146]), .Z(n28553) );
  NAND U38722 ( .A(n28555), .B(n28556), .Z(c[145]) );
  NAND U38723 ( .A(n26658), .B(o[145]), .Z(n28556) );
  NAND U38724 ( .A(n26653), .B(creg[145]), .Z(n28555) );
  NAND U38725 ( .A(n28557), .B(n28558), .Z(c[144]) );
  NAND U38726 ( .A(n26658), .B(o[144]), .Z(n28558) );
  NAND U38727 ( .A(n26653), .B(creg[144]), .Z(n28557) );
  NAND U38728 ( .A(n28559), .B(n28560), .Z(c[143]) );
  NAND U38729 ( .A(n26658), .B(o[143]), .Z(n28560) );
  NAND U38730 ( .A(n26653), .B(creg[143]), .Z(n28559) );
  NAND U38731 ( .A(n28561), .B(n28562), .Z(c[142]) );
  NAND U38732 ( .A(n26658), .B(o[142]), .Z(n28562) );
  NAND U38733 ( .A(n26653), .B(creg[142]), .Z(n28561) );
  NAND U38734 ( .A(n28563), .B(n28564), .Z(c[141]) );
  NAND U38735 ( .A(n26658), .B(o[141]), .Z(n28564) );
  NAND U38736 ( .A(n26653), .B(creg[141]), .Z(n28563) );
  NAND U38737 ( .A(n28565), .B(n28566), .Z(c[140]) );
  NAND U38738 ( .A(n26658), .B(o[140]), .Z(n28566) );
  NAND U38739 ( .A(n26653), .B(creg[140]), .Z(n28565) );
  NAND U38740 ( .A(n28567), .B(n28568), .Z(c[13]) );
  NAND U38741 ( .A(n26658), .B(o[13]), .Z(n28568) );
  NAND U38742 ( .A(n26653), .B(creg[13]), .Z(n28567) );
  NAND U38743 ( .A(n28569), .B(n28570), .Z(c[139]) );
  NAND U38744 ( .A(n26658), .B(o[139]), .Z(n28570) );
  NAND U38745 ( .A(n26653), .B(creg[139]), .Z(n28569) );
  NAND U38746 ( .A(n28571), .B(n28572), .Z(c[138]) );
  NAND U38747 ( .A(n26658), .B(o[138]), .Z(n28572) );
  NAND U38748 ( .A(n26653), .B(creg[138]), .Z(n28571) );
  NAND U38749 ( .A(n28573), .B(n28574), .Z(c[137]) );
  NAND U38750 ( .A(n26658), .B(o[137]), .Z(n28574) );
  NAND U38751 ( .A(n26653), .B(creg[137]), .Z(n28573) );
  NAND U38752 ( .A(n28575), .B(n28576), .Z(c[136]) );
  NAND U38753 ( .A(n26658), .B(o[136]), .Z(n28576) );
  NAND U38754 ( .A(n26653), .B(creg[136]), .Z(n28575) );
  NAND U38755 ( .A(n28577), .B(n28578), .Z(c[135]) );
  NAND U38756 ( .A(n26658), .B(o[135]), .Z(n28578) );
  NAND U38757 ( .A(n26653), .B(creg[135]), .Z(n28577) );
  NAND U38758 ( .A(n28579), .B(n28580), .Z(c[134]) );
  NAND U38759 ( .A(n26658), .B(o[134]), .Z(n28580) );
  NAND U38760 ( .A(n26653), .B(creg[134]), .Z(n28579) );
  NAND U38761 ( .A(n28581), .B(n28582), .Z(c[133]) );
  NAND U38762 ( .A(n26658), .B(o[133]), .Z(n28582) );
  NAND U38763 ( .A(n26653), .B(creg[133]), .Z(n28581) );
  NAND U38764 ( .A(n28583), .B(n28584), .Z(c[132]) );
  NAND U38765 ( .A(n26658), .B(o[132]), .Z(n28584) );
  NAND U38766 ( .A(n26653), .B(creg[132]), .Z(n28583) );
  NAND U38767 ( .A(n28585), .B(n28586), .Z(c[131]) );
  NAND U38768 ( .A(n26658), .B(o[131]), .Z(n28586) );
  NAND U38769 ( .A(n26653), .B(creg[131]), .Z(n28585) );
  NAND U38770 ( .A(n28587), .B(n28588), .Z(c[130]) );
  NAND U38771 ( .A(n26658), .B(o[130]), .Z(n28588) );
  NAND U38772 ( .A(n26653), .B(creg[130]), .Z(n28587) );
  NAND U38773 ( .A(n28589), .B(n28590), .Z(c[12]) );
  NAND U38774 ( .A(n26658), .B(o[12]), .Z(n28590) );
  NAND U38775 ( .A(n26653), .B(creg[12]), .Z(n28589) );
  NAND U38776 ( .A(n28591), .B(n28592), .Z(c[129]) );
  NAND U38777 ( .A(n26658), .B(o[129]), .Z(n28592) );
  NAND U38778 ( .A(n26653), .B(creg[129]), .Z(n28591) );
  NAND U38779 ( .A(n28593), .B(n28594), .Z(c[128]) );
  NAND U38780 ( .A(n26658), .B(o[128]), .Z(n28594) );
  NAND U38781 ( .A(n26653), .B(creg[128]), .Z(n28593) );
  NAND U38782 ( .A(n28595), .B(n28596), .Z(c[127]) );
  NAND U38783 ( .A(n26658), .B(o[127]), .Z(n28596) );
  NAND U38784 ( .A(n26653), .B(creg[127]), .Z(n28595) );
  NAND U38785 ( .A(n28597), .B(n28598), .Z(c[126]) );
  NAND U38786 ( .A(n26658), .B(o[126]), .Z(n28598) );
  NAND U38787 ( .A(n26653), .B(creg[126]), .Z(n28597) );
  NAND U38788 ( .A(n28599), .B(n28600), .Z(c[125]) );
  NAND U38789 ( .A(n26658), .B(o[125]), .Z(n28600) );
  NAND U38790 ( .A(n26653), .B(creg[125]), .Z(n28599) );
  NAND U38791 ( .A(n28601), .B(n28602), .Z(c[124]) );
  NAND U38792 ( .A(n26658), .B(o[124]), .Z(n28602) );
  NAND U38793 ( .A(n26653), .B(creg[124]), .Z(n28601) );
  NAND U38794 ( .A(n28603), .B(n28604), .Z(c[123]) );
  NAND U38795 ( .A(n26658), .B(o[123]), .Z(n28604) );
  NAND U38796 ( .A(n26653), .B(creg[123]), .Z(n28603) );
  NAND U38797 ( .A(n28605), .B(n28606), .Z(c[122]) );
  NAND U38798 ( .A(n26658), .B(o[122]), .Z(n28606) );
  NAND U38799 ( .A(n26653), .B(creg[122]), .Z(n28605) );
  NAND U38800 ( .A(n28607), .B(n28608), .Z(c[121]) );
  NAND U38801 ( .A(n26658), .B(o[121]), .Z(n28608) );
  NAND U38802 ( .A(n26653), .B(creg[121]), .Z(n28607) );
  NAND U38803 ( .A(n28609), .B(n28610), .Z(c[120]) );
  NAND U38804 ( .A(n26658), .B(o[120]), .Z(n28610) );
  NAND U38805 ( .A(n26653), .B(creg[120]), .Z(n28609) );
  NAND U38806 ( .A(n28611), .B(n28612), .Z(c[11]) );
  NAND U38807 ( .A(n26658), .B(o[11]), .Z(n28612) );
  NAND U38808 ( .A(n26653), .B(creg[11]), .Z(n28611) );
  NAND U38809 ( .A(n28613), .B(n28614), .Z(c[119]) );
  NAND U38810 ( .A(n26658), .B(o[119]), .Z(n28614) );
  NAND U38811 ( .A(n26653), .B(creg[119]), .Z(n28613) );
  NAND U38812 ( .A(n28615), .B(n28616), .Z(c[118]) );
  NAND U38813 ( .A(n26658), .B(o[118]), .Z(n28616) );
  NAND U38814 ( .A(n26653), .B(creg[118]), .Z(n28615) );
  NAND U38815 ( .A(n28617), .B(n28618), .Z(c[117]) );
  NAND U38816 ( .A(n26658), .B(o[117]), .Z(n28618) );
  NAND U38817 ( .A(n26653), .B(creg[117]), .Z(n28617) );
  NAND U38818 ( .A(n28619), .B(n28620), .Z(c[116]) );
  NAND U38819 ( .A(n26658), .B(o[116]), .Z(n28620) );
  NAND U38820 ( .A(n26653), .B(creg[116]), .Z(n28619) );
  NAND U38821 ( .A(n28621), .B(n28622), .Z(c[115]) );
  NAND U38822 ( .A(n26658), .B(o[115]), .Z(n28622) );
  NAND U38823 ( .A(n26653), .B(creg[115]), .Z(n28621) );
  NAND U38824 ( .A(n28623), .B(n28624), .Z(c[114]) );
  NAND U38825 ( .A(n26658), .B(o[114]), .Z(n28624) );
  NAND U38826 ( .A(n26653), .B(creg[114]), .Z(n28623) );
  NAND U38827 ( .A(n28625), .B(n28626), .Z(c[113]) );
  NAND U38828 ( .A(n26658), .B(o[113]), .Z(n28626) );
  NAND U38829 ( .A(n26653), .B(creg[113]), .Z(n28625) );
  NAND U38830 ( .A(n28627), .B(n28628), .Z(c[112]) );
  NAND U38831 ( .A(n26658), .B(o[112]), .Z(n28628) );
  NAND U38832 ( .A(n26653), .B(creg[112]), .Z(n28627) );
  NAND U38833 ( .A(n28629), .B(n28630), .Z(c[111]) );
  NAND U38834 ( .A(n26658), .B(o[111]), .Z(n28630) );
  NAND U38835 ( .A(n26653), .B(creg[111]), .Z(n28629) );
  NAND U38836 ( .A(n28631), .B(n28632), .Z(c[110]) );
  NAND U38837 ( .A(n26658), .B(o[110]), .Z(n28632) );
  NAND U38838 ( .A(n26653), .B(creg[110]), .Z(n28631) );
  NAND U38839 ( .A(n28633), .B(n28634), .Z(c[10]) );
  NAND U38840 ( .A(n26658), .B(o[10]), .Z(n28634) );
  NAND U38841 ( .A(n26653), .B(creg[10]), .Z(n28633) );
  NAND U38842 ( .A(n28635), .B(n28636), .Z(c[109]) );
  NAND U38843 ( .A(n26658), .B(o[109]), .Z(n28636) );
  NAND U38844 ( .A(n26653), .B(creg[109]), .Z(n28635) );
  NAND U38845 ( .A(n28637), .B(n28638), .Z(c[108]) );
  NAND U38846 ( .A(n26658), .B(o[108]), .Z(n28638) );
  NAND U38847 ( .A(n26653), .B(creg[108]), .Z(n28637) );
  NAND U38848 ( .A(n28639), .B(n28640), .Z(c[107]) );
  NAND U38849 ( .A(n26658), .B(o[107]), .Z(n28640) );
  NAND U38850 ( .A(n26653), .B(creg[107]), .Z(n28639) );
  NAND U38851 ( .A(n28641), .B(n28642), .Z(c[106]) );
  NAND U38852 ( .A(n26658), .B(o[106]), .Z(n28642) );
  NAND U38853 ( .A(n26653), .B(creg[106]), .Z(n28641) );
  NAND U38854 ( .A(n28643), .B(n28644), .Z(c[105]) );
  NAND U38855 ( .A(n26658), .B(o[105]), .Z(n28644) );
  NAND U38856 ( .A(n26653), .B(creg[105]), .Z(n28643) );
  NAND U38857 ( .A(n28645), .B(n28646), .Z(c[104]) );
  NAND U38858 ( .A(n26658), .B(o[104]), .Z(n28646) );
  NAND U38859 ( .A(n26653), .B(creg[104]), .Z(n28645) );
  NAND U38860 ( .A(n28647), .B(n28648), .Z(c[103]) );
  NAND U38861 ( .A(n26658), .B(o[103]), .Z(n28648) );
  NAND U38862 ( .A(n26653), .B(creg[103]), .Z(n28647) );
  NAND U38863 ( .A(n28649), .B(n28650), .Z(c[102]) );
  NAND U38864 ( .A(n26658), .B(o[102]), .Z(n28650) );
  NAND U38865 ( .A(n26653), .B(creg[102]), .Z(n28649) );
  NAND U38866 ( .A(n28651), .B(n28652), .Z(c[1023]) );
  NAND U38867 ( .A(n26658), .B(o[1023]), .Z(n28652) );
  NAND U38868 ( .A(n26653), .B(creg[1023]), .Z(n28651) );
  NAND U38869 ( .A(n28653), .B(n28654), .Z(c[1022]) );
  NAND U38870 ( .A(n26658), .B(o[1022]), .Z(n28654) );
  NAND U38871 ( .A(n26653), .B(creg[1022]), .Z(n28653) );
  NAND U38872 ( .A(n28655), .B(n28656), .Z(c[1021]) );
  NAND U38873 ( .A(n26658), .B(o[1021]), .Z(n28656) );
  NAND U38874 ( .A(n26653), .B(creg[1021]), .Z(n28655) );
  NAND U38875 ( .A(n28657), .B(n28658), .Z(c[1020]) );
  NAND U38876 ( .A(n26658), .B(o[1020]), .Z(n28658) );
  NAND U38877 ( .A(n26653), .B(creg[1020]), .Z(n28657) );
  NAND U38878 ( .A(n28659), .B(n28660), .Z(c[101]) );
  NAND U38879 ( .A(n26658), .B(o[101]), .Z(n28660) );
  NAND U38880 ( .A(n26653), .B(creg[101]), .Z(n28659) );
  NAND U38881 ( .A(n28661), .B(n28662), .Z(c[1019]) );
  NAND U38882 ( .A(n26658), .B(o[1019]), .Z(n28662) );
  NAND U38883 ( .A(n26653), .B(creg[1019]), .Z(n28661) );
  NAND U38884 ( .A(n28663), .B(n28664), .Z(c[1018]) );
  NAND U38885 ( .A(n26658), .B(o[1018]), .Z(n28664) );
  NAND U38886 ( .A(n26653), .B(creg[1018]), .Z(n28663) );
  NAND U38887 ( .A(n28665), .B(n28666), .Z(c[1017]) );
  NAND U38888 ( .A(n26658), .B(o[1017]), .Z(n28666) );
  NAND U38889 ( .A(n26653), .B(creg[1017]), .Z(n28665) );
  NAND U38890 ( .A(n28667), .B(n28668), .Z(c[1016]) );
  NAND U38891 ( .A(n26658), .B(o[1016]), .Z(n28668) );
  NAND U38892 ( .A(n26653), .B(creg[1016]), .Z(n28667) );
  NAND U38893 ( .A(n28669), .B(n28670), .Z(c[1015]) );
  NAND U38894 ( .A(n26658), .B(o[1015]), .Z(n28670) );
  NAND U38895 ( .A(n26653), .B(creg[1015]), .Z(n28669) );
  NAND U38896 ( .A(n28671), .B(n28672), .Z(c[1014]) );
  NAND U38897 ( .A(n26658), .B(o[1014]), .Z(n28672) );
  NAND U38898 ( .A(n26653), .B(creg[1014]), .Z(n28671) );
  NAND U38899 ( .A(n28673), .B(n28674), .Z(c[1013]) );
  NAND U38900 ( .A(n26658), .B(o[1013]), .Z(n28674) );
  NAND U38901 ( .A(n26653), .B(creg[1013]), .Z(n28673) );
  NAND U38902 ( .A(n28675), .B(n28676), .Z(c[1012]) );
  NAND U38903 ( .A(n26658), .B(o[1012]), .Z(n28676) );
  NAND U38904 ( .A(n26653), .B(creg[1012]), .Z(n28675) );
  NAND U38905 ( .A(n28677), .B(n28678), .Z(c[1011]) );
  NAND U38906 ( .A(n26658), .B(o[1011]), .Z(n28678) );
  NAND U38907 ( .A(n26653), .B(creg[1011]), .Z(n28677) );
  NAND U38908 ( .A(n28679), .B(n28680), .Z(c[1010]) );
  NAND U38909 ( .A(n26658), .B(o[1010]), .Z(n28680) );
  NAND U38910 ( .A(n26653), .B(creg[1010]), .Z(n28679) );
  NAND U38911 ( .A(n28681), .B(n28682), .Z(c[100]) );
  NAND U38912 ( .A(n26658), .B(o[100]), .Z(n28682) );
  NAND U38913 ( .A(n26653), .B(creg[100]), .Z(n28681) );
  NAND U38914 ( .A(n28683), .B(n28684), .Z(c[1009]) );
  NAND U38915 ( .A(n26658), .B(o[1009]), .Z(n28684) );
  NAND U38916 ( .A(n26653), .B(creg[1009]), .Z(n28683) );
  NAND U38917 ( .A(n28685), .B(n28686), .Z(c[1008]) );
  NAND U38918 ( .A(n26658), .B(o[1008]), .Z(n28686) );
  NAND U38919 ( .A(n26653), .B(creg[1008]), .Z(n28685) );
  NAND U38920 ( .A(n28687), .B(n28688), .Z(c[1007]) );
  NAND U38921 ( .A(n26658), .B(o[1007]), .Z(n28688) );
  NAND U38922 ( .A(n26653), .B(creg[1007]), .Z(n28687) );
  NAND U38923 ( .A(n28689), .B(n28690), .Z(c[1006]) );
  NAND U38924 ( .A(n26658), .B(o[1006]), .Z(n28690) );
  NAND U38925 ( .A(n26653), .B(creg[1006]), .Z(n28689) );
  NAND U38926 ( .A(n28691), .B(n28692), .Z(c[1005]) );
  NAND U38927 ( .A(n26658), .B(o[1005]), .Z(n28692) );
  NAND U38928 ( .A(n26653), .B(creg[1005]), .Z(n28691) );
  NAND U38929 ( .A(n28693), .B(n28694), .Z(c[1004]) );
  NAND U38930 ( .A(n26658), .B(o[1004]), .Z(n28694) );
  NAND U38931 ( .A(n26653), .B(creg[1004]), .Z(n28693) );
  NAND U38932 ( .A(n28695), .B(n28696), .Z(c[1003]) );
  NAND U38933 ( .A(n26658), .B(o[1003]), .Z(n28696) );
  NAND U38934 ( .A(n26653), .B(creg[1003]), .Z(n28695) );
  NAND U38935 ( .A(n28697), .B(n28698), .Z(c[1002]) );
  NAND U38936 ( .A(n26658), .B(o[1002]), .Z(n28698) );
  NAND U38937 ( .A(n26653), .B(creg[1002]), .Z(n28697) );
  NAND U38938 ( .A(n28699), .B(n28700), .Z(c[1001]) );
  NAND U38939 ( .A(n26658), .B(o[1001]), .Z(n28700) );
  NAND U38940 ( .A(n26653), .B(creg[1001]), .Z(n28699) );
  NAND U38941 ( .A(n28701), .B(n28702), .Z(c[1000]) );
  NAND U38942 ( .A(n26658), .B(o[1000]), .Z(n28702) );
  NAND U38943 ( .A(n26653), .B(creg[1000]), .Z(n28701) );
  NAND U38944 ( .A(n28703), .B(n28704), .Z(c[0]) );
  NAND U38945 ( .A(n26658), .B(o[0]), .Z(n28704) );
  IV U38946 ( .A(n26653), .Z(n26658) );
  NAND U38947 ( .A(n26653), .B(creg[0]), .Z(n28703) );
  NAND U38948 ( .A(n28705), .B(n28706), .Z(n26653) );
  NANDN U38949 ( .A(ereg[1023]), .B(init), .Z(n28706) );
  OR U38950 ( .A(init), .B(e[1023]), .Z(n28705) );
endmodule

