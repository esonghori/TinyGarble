
module sum_N1024_CC2 ( clk, rst, a, b, c );
  input [511:0] a;
  input [511:0] b;
  output [511:0] c;
  input clk, rst;
  wire   carry_on, carry_on_d, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
         n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
         n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
         n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
         n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
         n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
         n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
         n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
         n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
         n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
         n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
         n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
         n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
         n2049, n2050;

  DFF carry_on_reg ( .D(carry_on_d), .CLK(clk), .RST(rst), .Q(carry_on) );
  NAND U3 ( .A(carry_on), .B(a[0]), .Z(n1) );
  XOR U4 ( .A(a[0]), .B(carry_on), .Z(n2) );
  NAND U5 ( .A(n2), .B(b[0]), .Z(n3) );
  NAND U6 ( .A(n1), .B(n3), .Z(n11) );
  NAND U7 ( .A(n1552), .B(b[386]), .Z(n4) );
  XOR U8 ( .A(b[386]), .B(n1552), .Z(n5) );
  NAND U9 ( .A(n5), .B(a[386]), .Z(n6) );
  NAND U10 ( .A(n4), .B(n6), .Z(n1553) );
  NAND U11 ( .A(n2050), .B(b[511]), .Z(n7) );
  XOR U12 ( .A(b[511]), .B(n2050), .Z(n8) );
  NAND U13 ( .A(n8), .B(a[511]), .Z(n9) );
  NAND U14 ( .A(n7), .B(n9), .Z(carry_on_d) );
  XNOR U15 ( .A(b[0]), .B(a[0]), .Z(n10) );
  XNOR U16 ( .A(carry_on), .B(n10), .Z(c[0]) );
  XOR U17 ( .A(a[1]), .B(b[1]), .Z(n12) );
  XOR U18 ( .A(n11), .B(n12), .Z(c[1]) );
  XOR U19 ( .A(a[2]), .B(b[2]), .Z(n15) );
  NAND U20 ( .A(b[1]), .B(a[1]), .Z(n14) );
  NAND U21 ( .A(n12), .B(n11), .Z(n13) );
  AND U22 ( .A(n14), .B(n13), .Z(n16) );
  XNOR U23 ( .A(n15), .B(n16), .Z(c[2]) );
  XOR U24 ( .A(a[3]), .B(b[3]), .Z(n19) );
  NAND U25 ( .A(b[2]), .B(a[2]), .Z(n18) );
  NANDN U26 ( .A(n16), .B(n15), .Z(n17) );
  AND U27 ( .A(n18), .B(n17), .Z(n20) );
  XNOR U28 ( .A(n19), .B(n20), .Z(c[3]) );
  XOR U29 ( .A(a[4]), .B(b[4]), .Z(n23) );
  NAND U30 ( .A(b[3]), .B(a[3]), .Z(n22) );
  NANDN U31 ( .A(n20), .B(n19), .Z(n21) );
  AND U32 ( .A(n22), .B(n21), .Z(n24) );
  XNOR U33 ( .A(n23), .B(n24), .Z(c[4]) );
  XOR U34 ( .A(a[5]), .B(b[5]), .Z(n27) );
  NAND U35 ( .A(b[4]), .B(a[4]), .Z(n26) );
  NANDN U36 ( .A(n24), .B(n23), .Z(n25) );
  AND U37 ( .A(n26), .B(n25), .Z(n28) );
  XNOR U38 ( .A(n27), .B(n28), .Z(c[5]) );
  NAND U39 ( .A(b[5]), .B(a[5]), .Z(n30) );
  NANDN U40 ( .A(n28), .B(n27), .Z(n29) );
  NAND U41 ( .A(n30), .B(n29), .Z(n32) );
  XNOR U42 ( .A(b[6]), .B(a[6]), .Z(n31) );
  XNOR U43 ( .A(n32), .B(n31), .Z(c[6]) );
  XOR U44 ( .A(a[7]), .B(b[7]), .Z(n35) );
  OR U45 ( .A(b[6]), .B(a[6]), .Z(n34) );
  OR U46 ( .A(n32), .B(n31), .Z(n33) );
  NAND U47 ( .A(n34), .B(n33), .Z(n36) );
  XNOR U48 ( .A(n35), .B(n36), .Z(c[7]) );
  NAND U49 ( .A(b[7]), .B(a[7]), .Z(n38) );
  NANDN U50 ( .A(n36), .B(n35), .Z(n37) );
  NAND U51 ( .A(n38), .B(n37), .Z(n40) );
  XNOR U52 ( .A(b[8]), .B(a[8]), .Z(n39) );
  XNOR U53 ( .A(n40), .B(n39), .Z(c[8]) );
  XNOR U54 ( .A(b[9]), .B(a[9]), .Z(n44) );
  OR U55 ( .A(b[8]), .B(a[8]), .Z(n42) );
  OR U56 ( .A(n40), .B(n39), .Z(n41) );
  AND U57 ( .A(n42), .B(n41), .Z(n43) );
  XNOR U58 ( .A(n44), .B(n43), .Z(c[9]) );
  XNOR U59 ( .A(b[10]), .B(a[10]), .Z(n48) );
  OR U60 ( .A(b[9]), .B(a[9]), .Z(n46) );
  OR U61 ( .A(n44), .B(n43), .Z(n45) );
  AND U62 ( .A(n46), .B(n45), .Z(n47) );
  XNOR U63 ( .A(n48), .B(n47), .Z(c[10]) );
  XNOR U64 ( .A(b[11]), .B(a[11]), .Z(n52) );
  OR U65 ( .A(b[10]), .B(a[10]), .Z(n50) );
  OR U66 ( .A(n48), .B(n47), .Z(n49) );
  AND U67 ( .A(n50), .B(n49), .Z(n51) );
  XNOR U68 ( .A(n52), .B(n51), .Z(c[11]) );
  XNOR U69 ( .A(b[12]), .B(a[12]), .Z(n56) );
  OR U70 ( .A(b[11]), .B(a[11]), .Z(n54) );
  OR U71 ( .A(n52), .B(n51), .Z(n53) );
  AND U72 ( .A(n54), .B(n53), .Z(n55) );
  XNOR U73 ( .A(n56), .B(n55), .Z(c[12]) );
  XNOR U74 ( .A(b[13]), .B(a[13]), .Z(n60) );
  OR U75 ( .A(b[12]), .B(a[12]), .Z(n58) );
  OR U76 ( .A(n56), .B(n55), .Z(n57) );
  AND U77 ( .A(n58), .B(n57), .Z(n59) );
  XNOR U78 ( .A(n60), .B(n59), .Z(c[13]) );
  XNOR U79 ( .A(b[14]), .B(a[14]), .Z(n64) );
  OR U80 ( .A(b[13]), .B(a[13]), .Z(n62) );
  OR U81 ( .A(n60), .B(n59), .Z(n61) );
  AND U82 ( .A(n62), .B(n61), .Z(n63) );
  XNOR U83 ( .A(n64), .B(n63), .Z(c[14]) );
  OR U84 ( .A(b[14]), .B(a[14]), .Z(n66) );
  OR U85 ( .A(n64), .B(n63), .Z(n65) );
  NAND U86 ( .A(n66), .B(n65), .Z(n68) );
  XOR U87 ( .A(a[15]), .B(b[15]), .Z(n67) );
  XNOR U88 ( .A(n68), .B(n67), .Z(c[15]) );
  XOR U89 ( .A(a[16]), .B(b[16]), .Z(n71) );
  NAND U90 ( .A(b[15]), .B(a[15]), .Z(n70) );
  NANDN U91 ( .A(n68), .B(n67), .Z(n69) );
  AND U92 ( .A(n70), .B(n69), .Z(n72) );
  XNOR U93 ( .A(n71), .B(n72), .Z(c[16]) );
  XOR U94 ( .A(a[17]), .B(b[17]), .Z(n75) );
  NAND U95 ( .A(b[16]), .B(a[16]), .Z(n74) );
  NANDN U96 ( .A(n72), .B(n71), .Z(n73) );
  AND U97 ( .A(n74), .B(n73), .Z(n76) );
  XNOR U98 ( .A(n75), .B(n76), .Z(c[17]) );
  XOR U99 ( .A(a[18]), .B(b[18]), .Z(n79) );
  NAND U100 ( .A(b[17]), .B(a[17]), .Z(n78) );
  NANDN U101 ( .A(n76), .B(n75), .Z(n77) );
  AND U102 ( .A(n78), .B(n77), .Z(n80) );
  XNOR U103 ( .A(n79), .B(n80), .Z(c[18]) );
  XOR U104 ( .A(a[19]), .B(b[19]), .Z(n83) );
  NAND U105 ( .A(b[18]), .B(a[18]), .Z(n82) );
  NANDN U106 ( .A(n80), .B(n79), .Z(n81) );
  AND U107 ( .A(n82), .B(n81), .Z(n84) );
  XNOR U108 ( .A(n83), .B(n84), .Z(c[19]) );
  XOR U109 ( .A(a[20]), .B(b[20]), .Z(n87) );
  NAND U110 ( .A(b[19]), .B(a[19]), .Z(n86) );
  NANDN U111 ( .A(n84), .B(n83), .Z(n85) );
  AND U112 ( .A(n86), .B(n85), .Z(n88) );
  XNOR U113 ( .A(n87), .B(n88), .Z(c[20]) );
  XOR U114 ( .A(a[21]), .B(b[21]), .Z(n91) );
  NAND U115 ( .A(b[20]), .B(a[20]), .Z(n90) );
  NANDN U116 ( .A(n88), .B(n87), .Z(n89) );
  AND U117 ( .A(n90), .B(n89), .Z(n92) );
  XNOR U118 ( .A(n91), .B(n92), .Z(c[21]) );
  XOR U119 ( .A(a[22]), .B(b[22]), .Z(n95) );
  NAND U120 ( .A(b[21]), .B(a[21]), .Z(n94) );
  NANDN U121 ( .A(n92), .B(n91), .Z(n93) );
  AND U122 ( .A(n94), .B(n93), .Z(n96) );
  XNOR U123 ( .A(n95), .B(n96), .Z(c[22]) );
  XOR U124 ( .A(a[23]), .B(b[23]), .Z(n99) );
  NAND U125 ( .A(b[22]), .B(a[22]), .Z(n98) );
  NANDN U126 ( .A(n96), .B(n95), .Z(n97) );
  AND U127 ( .A(n98), .B(n97), .Z(n100) );
  XNOR U128 ( .A(n99), .B(n100), .Z(c[23]) );
  XOR U129 ( .A(a[24]), .B(b[24]), .Z(n103) );
  NAND U130 ( .A(b[23]), .B(a[23]), .Z(n102) );
  NANDN U131 ( .A(n100), .B(n99), .Z(n101) );
  AND U132 ( .A(n102), .B(n101), .Z(n104) );
  XNOR U133 ( .A(n103), .B(n104), .Z(c[24]) );
  XOR U134 ( .A(a[25]), .B(b[25]), .Z(n107) );
  NAND U135 ( .A(b[24]), .B(a[24]), .Z(n106) );
  NANDN U136 ( .A(n104), .B(n103), .Z(n105) );
  AND U137 ( .A(n106), .B(n105), .Z(n108) );
  XNOR U138 ( .A(n107), .B(n108), .Z(c[25]) );
  NAND U139 ( .A(b[25]), .B(a[25]), .Z(n110) );
  NANDN U140 ( .A(n108), .B(n107), .Z(n109) );
  NAND U141 ( .A(n110), .B(n109), .Z(n112) );
  XNOR U142 ( .A(b[26]), .B(a[26]), .Z(n111) );
  XNOR U143 ( .A(n112), .B(n111), .Z(c[26]) );
  OR U144 ( .A(b[26]), .B(a[26]), .Z(n114) );
  OR U145 ( .A(n112), .B(n111), .Z(n113) );
  NAND U146 ( .A(n114), .B(n113), .Z(n116) );
  XOR U147 ( .A(a[27]), .B(b[27]), .Z(n115) );
  XNOR U148 ( .A(n116), .B(n115), .Z(c[27]) );
  XOR U149 ( .A(a[28]), .B(b[28]), .Z(n119) );
  NAND U150 ( .A(b[27]), .B(a[27]), .Z(n118) );
  NANDN U151 ( .A(n116), .B(n115), .Z(n117) );
  AND U152 ( .A(n118), .B(n117), .Z(n120) );
  XNOR U153 ( .A(n119), .B(n120), .Z(c[28]) );
  XOR U154 ( .A(a[29]), .B(b[29]), .Z(n123) );
  NAND U155 ( .A(b[28]), .B(a[28]), .Z(n122) );
  NANDN U156 ( .A(n120), .B(n119), .Z(n121) );
  AND U157 ( .A(n122), .B(n121), .Z(n124) );
  XNOR U158 ( .A(n123), .B(n124), .Z(c[29]) );
  XOR U159 ( .A(a[30]), .B(b[30]), .Z(n127) );
  NAND U160 ( .A(b[29]), .B(a[29]), .Z(n126) );
  NANDN U161 ( .A(n124), .B(n123), .Z(n125) );
  AND U162 ( .A(n126), .B(n125), .Z(n128) );
  XNOR U163 ( .A(n127), .B(n128), .Z(c[30]) );
  XOR U164 ( .A(a[31]), .B(b[31]), .Z(n131) );
  NAND U165 ( .A(b[30]), .B(a[30]), .Z(n130) );
  NANDN U166 ( .A(n128), .B(n127), .Z(n129) );
  AND U167 ( .A(n130), .B(n129), .Z(n132) );
  XNOR U168 ( .A(n131), .B(n132), .Z(c[31]) );
  XOR U169 ( .A(a[32]), .B(b[32]), .Z(n135) );
  NAND U170 ( .A(b[31]), .B(a[31]), .Z(n134) );
  NANDN U171 ( .A(n132), .B(n131), .Z(n133) );
  AND U172 ( .A(n134), .B(n133), .Z(n136) );
  XNOR U173 ( .A(n135), .B(n136), .Z(c[32]) );
  XOR U174 ( .A(a[33]), .B(b[33]), .Z(n139) );
  NAND U175 ( .A(b[32]), .B(a[32]), .Z(n138) );
  NANDN U176 ( .A(n136), .B(n135), .Z(n137) );
  AND U177 ( .A(n138), .B(n137), .Z(n140) );
  XNOR U178 ( .A(n139), .B(n140), .Z(c[33]) );
  XOR U179 ( .A(a[34]), .B(b[34]), .Z(n143) );
  NAND U180 ( .A(b[33]), .B(a[33]), .Z(n142) );
  NANDN U181 ( .A(n140), .B(n139), .Z(n141) );
  AND U182 ( .A(n142), .B(n141), .Z(n144) );
  XNOR U183 ( .A(n143), .B(n144), .Z(c[34]) );
  XOR U184 ( .A(a[35]), .B(b[35]), .Z(n147) );
  NAND U185 ( .A(b[34]), .B(a[34]), .Z(n146) );
  NANDN U186 ( .A(n144), .B(n143), .Z(n145) );
  AND U187 ( .A(n146), .B(n145), .Z(n148) );
  XNOR U188 ( .A(n147), .B(n148), .Z(c[35]) );
  XOR U189 ( .A(a[36]), .B(b[36]), .Z(n151) );
  NAND U190 ( .A(b[35]), .B(a[35]), .Z(n150) );
  NANDN U191 ( .A(n148), .B(n147), .Z(n149) );
  AND U192 ( .A(n150), .B(n149), .Z(n152) );
  XNOR U193 ( .A(n151), .B(n152), .Z(c[36]) );
  XOR U194 ( .A(a[37]), .B(b[37]), .Z(n155) );
  NAND U195 ( .A(b[36]), .B(a[36]), .Z(n154) );
  NANDN U196 ( .A(n152), .B(n151), .Z(n153) );
  AND U197 ( .A(n154), .B(n153), .Z(n156) );
  XNOR U198 ( .A(n155), .B(n156), .Z(c[37]) );
  XOR U199 ( .A(a[38]), .B(b[38]), .Z(n159) );
  NAND U200 ( .A(b[37]), .B(a[37]), .Z(n158) );
  NANDN U201 ( .A(n156), .B(n155), .Z(n157) );
  AND U202 ( .A(n158), .B(n157), .Z(n160) );
  XNOR U203 ( .A(n159), .B(n160), .Z(c[38]) );
  XOR U204 ( .A(a[39]), .B(b[39]), .Z(n163) );
  NAND U205 ( .A(b[38]), .B(a[38]), .Z(n162) );
  NANDN U206 ( .A(n160), .B(n159), .Z(n161) );
  AND U207 ( .A(n162), .B(n161), .Z(n164) );
  XNOR U208 ( .A(n163), .B(n164), .Z(c[39]) );
  XOR U209 ( .A(a[40]), .B(b[40]), .Z(n167) );
  NAND U210 ( .A(b[39]), .B(a[39]), .Z(n166) );
  NANDN U211 ( .A(n164), .B(n163), .Z(n165) );
  AND U212 ( .A(n166), .B(n165), .Z(n168) );
  XNOR U213 ( .A(n167), .B(n168), .Z(c[40]) );
  XOR U214 ( .A(a[41]), .B(b[41]), .Z(n171) );
  NAND U215 ( .A(b[40]), .B(a[40]), .Z(n170) );
  NANDN U216 ( .A(n168), .B(n167), .Z(n169) );
  AND U217 ( .A(n170), .B(n169), .Z(n172) );
  XNOR U218 ( .A(n171), .B(n172), .Z(c[41]) );
  XOR U219 ( .A(a[42]), .B(b[42]), .Z(n175) );
  NAND U220 ( .A(b[41]), .B(a[41]), .Z(n174) );
  NANDN U221 ( .A(n172), .B(n171), .Z(n173) );
  AND U222 ( .A(n174), .B(n173), .Z(n176) );
  XNOR U223 ( .A(n175), .B(n176), .Z(c[42]) );
  XOR U224 ( .A(a[43]), .B(b[43]), .Z(n179) );
  NAND U225 ( .A(b[42]), .B(a[42]), .Z(n178) );
  NANDN U226 ( .A(n176), .B(n175), .Z(n177) );
  AND U227 ( .A(n178), .B(n177), .Z(n180) );
  XNOR U228 ( .A(n179), .B(n180), .Z(c[43]) );
  XOR U229 ( .A(a[44]), .B(b[44]), .Z(n183) );
  NAND U230 ( .A(b[43]), .B(a[43]), .Z(n182) );
  NANDN U231 ( .A(n180), .B(n179), .Z(n181) );
  AND U232 ( .A(n182), .B(n181), .Z(n184) );
  XNOR U233 ( .A(n183), .B(n184), .Z(c[44]) );
  XOR U234 ( .A(a[45]), .B(b[45]), .Z(n187) );
  NAND U235 ( .A(b[44]), .B(a[44]), .Z(n186) );
  NANDN U236 ( .A(n184), .B(n183), .Z(n185) );
  AND U237 ( .A(n186), .B(n185), .Z(n188) );
  XNOR U238 ( .A(n187), .B(n188), .Z(c[45]) );
  XOR U239 ( .A(a[46]), .B(b[46]), .Z(n191) );
  NAND U240 ( .A(b[45]), .B(a[45]), .Z(n190) );
  NANDN U241 ( .A(n188), .B(n187), .Z(n189) );
  AND U242 ( .A(n190), .B(n189), .Z(n192) );
  XNOR U243 ( .A(n191), .B(n192), .Z(c[46]) );
  XOR U244 ( .A(a[47]), .B(b[47]), .Z(n195) );
  NAND U245 ( .A(b[46]), .B(a[46]), .Z(n194) );
  NANDN U246 ( .A(n192), .B(n191), .Z(n193) );
  AND U247 ( .A(n194), .B(n193), .Z(n196) );
  XNOR U248 ( .A(n195), .B(n196), .Z(c[47]) );
  XOR U249 ( .A(a[48]), .B(b[48]), .Z(n199) );
  NAND U250 ( .A(b[47]), .B(a[47]), .Z(n198) );
  NANDN U251 ( .A(n196), .B(n195), .Z(n197) );
  AND U252 ( .A(n198), .B(n197), .Z(n200) );
  XNOR U253 ( .A(n199), .B(n200), .Z(c[48]) );
  XOR U254 ( .A(a[49]), .B(b[49]), .Z(n203) );
  NAND U255 ( .A(b[48]), .B(a[48]), .Z(n202) );
  NANDN U256 ( .A(n200), .B(n199), .Z(n201) );
  AND U257 ( .A(n202), .B(n201), .Z(n204) );
  XNOR U258 ( .A(n203), .B(n204), .Z(c[49]) );
  XOR U259 ( .A(a[50]), .B(b[50]), .Z(n207) );
  NAND U260 ( .A(b[49]), .B(a[49]), .Z(n206) );
  NANDN U261 ( .A(n204), .B(n203), .Z(n205) );
  AND U262 ( .A(n206), .B(n205), .Z(n208) );
  XNOR U263 ( .A(n207), .B(n208), .Z(c[50]) );
  XOR U264 ( .A(a[51]), .B(b[51]), .Z(n211) );
  NAND U265 ( .A(b[50]), .B(a[50]), .Z(n210) );
  NANDN U266 ( .A(n208), .B(n207), .Z(n209) );
  AND U267 ( .A(n210), .B(n209), .Z(n212) );
  XNOR U268 ( .A(n211), .B(n212), .Z(c[51]) );
  XOR U269 ( .A(a[52]), .B(b[52]), .Z(n215) );
  NAND U270 ( .A(b[51]), .B(a[51]), .Z(n214) );
  NANDN U271 ( .A(n212), .B(n211), .Z(n213) );
  AND U272 ( .A(n214), .B(n213), .Z(n216) );
  XNOR U273 ( .A(n215), .B(n216), .Z(c[52]) );
  XOR U274 ( .A(a[53]), .B(b[53]), .Z(n219) );
  NAND U275 ( .A(b[52]), .B(a[52]), .Z(n218) );
  NANDN U276 ( .A(n216), .B(n215), .Z(n217) );
  AND U277 ( .A(n218), .B(n217), .Z(n220) );
  XNOR U278 ( .A(n219), .B(n220), .Z(c[53]) );
  NAND U279 ( .A(b[53]), .B(a[53]), .Z(n222) );
  NANDN U280 ( .A(n220), .B(n219), .Z(n221) );
  NAND U281 ( .A(n222), .B(n221), .Z(n224) );
  XNOR U282 ( .A(b[54]), .B(a[54]), .Z(n223) );
  XNOR U283 ( .A(n224), .B(n223), .Z(c[54]) );
  XNOR U284 ( .A(b[55]), .B(a[55]), .Z(n228) );
  OR U285 ( .A(b[54]), .B(a[54]), .Z(n226) );
  OR U286 ( .A(n224), .B(n223), .Z(n225) );
  AND U287 ( .A(n226), .B(n225), .Z(n227) );
  XNOR U288 ( .A(n228), .B(n227), .Z(c[55]) );
  XNOR U289 ( .A(b[56]), .B(a[56]), .Z(n232) );
  OR U290 ( .A(b[55]), .B(a[55]), .Z(n230) );
  OR U291 ( .A(n228), .B(n227), .Z(n229) );
  AND U292 ( .A(n230), .B(n229), .Z(n231) );
  XNOR U293 ( .A(n232), .B(n231), .Z(c[56]) );
  XNOR U294 ( .A(b[57]), .B(a[57]), .Z(n236) );
  OR U295 ( .A(b[56]), .B(a[56]), .Z(n234) );
  OR U296 ( .A(n232), .B(n231), .Z(n233) );
  AND U297 ( .A(n234), .B(n233), .Z(n235) );
  XNOR U298 ( .A(n236), .B(n235), .Z(c[57]) );
  XNOR U299 ( .A(b[58]), .B(a[58]), .Z(n240) );
  OR U300 ( .A(b[57]), .B(a[57]), .Z(n238) );
  OR U301 ( .A(n236), .B(n235), .Z(n237) );
  AND U302 ( .A(n238), .B(n237), .Z(n239) );
  XNOR U303 ( .A(n240), .B(n239), .Z(c[58]) );
  XNOR U304 ( .A(b[59]), .B(a[59]), .Z(n244) );
  OR U305 ( .A(b[58]), .B(a[58]), .Z(n242) );
  OR U306 ( .A(n240), .B(n239), .Z(n241) );
  AND U307 ( .A(n242), .B(n241), .Z(n243) );
  XNOR U308 ( .A(n244), .B(n243), .Z(c[59]) );
  XNOR U309 ( .A(b[60]), .B(a[60]), .Z(n248) );
  OR U310 ( .A(b[59]), .B(a[59]), .Z(n246) );
  OR U311 ( .A(n244), .B(n243), .Z(n245) );
  AND U312 ( .A(n246), .B(n245), .Z(n247) );
  XNOR U313 ( .A(n248), .B(n247), .Z(c[60]) );
  XNOR U314 ( .A(b[61]), .B(a[61]), .Z(n252) );
  OR U315 ( .A(b[60]), .B(a[60]), .Z(n250) );
  OR U316 ( .A(n248), .B(n247), .Z(n249) );
  AND U317 ( .A(n250), .B(n249), .Z(n251) );
  XNOR U318 ( .A(n252), .B(n251), .Z(c[61]) );
  XNOR U319 ( .A(b[62]), .B(a[62]), .Z(n256) );
  OR U320 ( .A(b[61]), .B(a[61]), .Z(n254) );
  OR U321 ( .A(n252), .B(n251), .Z(n253) );
  AND U322 ( .A(n254), .B(n253), .Z(n255) );
  XNOR U323 ( .A(n256), .B(n255), .Z(c[62]) );
  XNOR U324 ( .A(b[63]), .B(a[63]), .Z(n260) );
  OR U325 ( .A(b[62]), .B(a[62]), .Z(n258) );
  OR U326 ( .A(n256), .B(n255), .Z(n257) );
  AND U327 ( .A(n258), .B(n257), .Z(n259) );
  XNOR U328 ( .A(n260), .B(n259), .Z(c[63]) );
  XNOR U329 ( .A(b[64]), .B(a[64]), .Z(n264) );
  OR U330 ( .A(b[63]), .B(a[63]), .Z(n262) );
  OR U331 ( .A(n260), .B(n259), .Z(n261) );
  AND U332 ( .A(n262), .B(n261), .Z(n263) );
  XNOR U333 ( .A(n264), .B(n263), .Z(c[64]) );
  XNOR U334 ( .A(b[65]), .B(a[65]), .Z(n268) );
  OR U335 ( .A(b[64]), .B(a[64]), .Z(n266) );
  OR U336 ( .A(n264), .B(n263), .Z(n265) );
  AND U337 ( .A(n266), .B(n265), .Z(n267) );
  XNOR U338 ( .A(n268), .B(n267), .Z(c[65]) );
  XNOR U339 ( .A(b[66]), .B(a[66]), .Z(n272) );
  OR U340 ( .A(b[65]), .B(a[65]), .Z(n270) );
  OR U341 ( .A(n268), .B(n267), .Z(n269) );
  AND U342 ( .A(n270), .B(n269), .Z(n271) );
  XNOR U343 ( .A(n272), .B(n271), .Z(c[66]) );
  XNOR U344 ( .A(b[67]), .B(a[67]), .Z(n276) );
  OR U345 ( .A(b[66]), .B(a[66]), .Z(n274) );
  OR U346 ( .A(n272), .B(n271), .Z(n273) );
  AND U347 ( .A(n274), .B(n273), .Z(n275) );
  XNOR U348 ( .A(n276), .B(n275), .Z(c[67]) );
  XNOR U349 ( .A(b[68]), .B(a[68]), .Z(n280) );
  OR U350 ( .A(b[67]), .B(a[67]), .Z(n278) );
  OR U351 ( .A(n276), .B(n275), .Z(n277) );
  AND U352 ( .A(n278), .B(n277), .Z(n279) );
  XNOR U353 ( .A(n280), .B(n279), .Z(c[68]) );
  XNOR U354 ( .A(b[69]), .B(a[69]), .Z(n284) );
  OR U355 ( .A(b[68]), .B(a[68]), .Z(n282) );
  OR U356 ( .A(n280), .B(n279), .Z(n281) );
  AND U357 ( .A(n282), .B(n281), .Z(n283) );
  XNOR U358 ( .A(n284), .B(n283), .Z(c[69]) );
  XNOR U359 ( .A(b[70]), .B(a[70]), .Z(n288) );
  OR U360 ( .A(b[69]), .B(a[69]), .Z(n286) );
  OR U361 ( .A(n284), .B(n283), .Z(n285) );
  AND U362 ( .A(n286), .B(n285), .Z(n287) );
  XNOR U363 ( .A(n288), .B(n287), .Z(c[70]) );
  XNOR U364 ( .A(b[71]), .B(a[71]), .Z(n292) );
  OR U365 ( .A(b[70]), .B(a[70]), .Z(n290) );
  OR U366 ( .A(n288), .B(n287), .Z(n289) );
  AND U367 ( .A(n290), .B(n289), .Z(n291) );
  XNOR U368 ( .A(n292), .B(n291), .Z(c[71]) );
  XNOR U369 ( .A(b[72]), .B(a[72]), .Z(n296) );
  OR U370 ( .A(b[71]), .B(a[71]), .Z(n294) );
  OR U371 ( .A(n292), .B(n291), .Z(n293) );
  AND U372 ( .A(n294), .B(n293), .Z(n295) );
  XNOR U373 ( .A(n296), .B(n295), .Z(c[72]) );
  XNOR U374 ( .A(b[73]), .B(a[73]), .Z(n300) );
  OR U375 ( .A(b[72]), .B(a[72]), .Z(n298) );
  OR U376 ( .A(n296), .B(n295), .Z(n297) );
  AND U377 ( .A(n298), .B(n297), .Z(n299) );
  XNOR U378 ( .A(n300), .B(n299), .Z(c[73]) );
  XNOR U379 ( .A(b[74]), .B(a[74]), .Z(n304) );
  OR U380 ( .A(b[73]), .B(a[73]), .Z(n302) );
  OR U381 ( .A(n300), .B(n299), .Z(n301) );
  AND U382 ( .A(n302), .B(n301), .Z(n303) );
  XNOR U383 ( .A(n304), .B(n303), .Z(c[74]) );
  XNOR U384 ( .A(b[75]), .B(a[75]), .Z(n308) );
  OR U385 ( .A(b[74]), .B(a[74]), .Z(n306) );
  OR U386 ( .A(n304), .B(n303), .Z(n305) );
  AND U387 ( .A(n306), .B(n305), .Z(n307) );
  XNOR U388 ( .A(n308), .B(n307), .Z(c[75]) );
  XNOR U389 ( .A(b[76]), .B(a[76]), .Z(n312) );
  OR U390 ( .A(b[75]), .B(a[75]), .Z(n310) );
  OR U391 ( .A(n308), .B(n307), .Z(n309) );
  AND U392 ( .A(n310), .B(n309), .Z(n311) );
  XNOR U393 ( .A(n312), .B(n311), .Z(c[76]) );
  XNOR U394 ( .A(b[77]), .B(a[77]), .Z(n316) );
  OR U395 ( .A(b[76]), .B(a[76]), .Z(n314) );
  OR U396 ( .A(n312), .B(n311), .Z(n313) );
  AND U397 ( .A(n314), .B(n313), .Z(n315) );
  XNOR U398 ( .A(n316), .B(n315), .Z(c[77]) );
  XNOR U399 ( .A(b[78]), .B(a[78]), .Z(n320) );
  OR U400 ( .A(b[77]), .B(a[77]), .Z(n318) );
  OR U401 ( .A(n316), .B(n315), .Z(n317) );
  AND U402 ( .A(n318), .B(n317), .Z(n319) );
  XNOR U403 ( .A(n320), .B(n319), .Z(c[78]) );
  XNOR U404 ( .A(b[79]), .B(a[79]), .Z(n324) );
  OR U405 ( .A(b[78]), .B(a[78]), .Z(n322) );
  OR U406 ( .A(n320), .B(n319), .Z(n321) );
  AND U407 ( .A(n322), .B(n321), .Z(n323) );
  XNOR U408 ( .A(n324), .B(n323), .Z(c[79]) );
  XNOR U409 ( .A(b[80]), .B(a[80]), .Z(n328) );
  OR U410 ( .A(b[79]), .B(a[79]), .Z(n326) );
  OR U411 ( .A(n324), .B(n323), .Z(n325) );
  AND U412 ( .A(n326), .B(n325), .Z(n327) );
  XNOR U413 ( .A(n328), .B(n327), .Z(c[80]) );
  OR U414 ( .A(b[80]), .B(a[80]), .Z(n330) );
  OR U415 ( .A(n328), .B(n327), .Z(n329) );
  NAND U416 ( .A(n330), .B(n329), .Z(n332) );
  XOR U417 ( .A(a[81]), .B(b[81]), .Z(n331) );
  XNOR U418 ( .A(n332), .B(n331), .Z(c[81]) );
  XOR U419 ( .A(a[82]), .B(b[82]), .Z(n335) );
  NAND U420 ( .A(b[81]), .B(a[81]), .Z(n334) );
  NANDN U421 ( .A(n332), .B(n331), .Z(n333) );
  AND U422 ( .A(n334), .B(n333), .Z(n336) );
  XNOR U423 ( .A(n335), .B(n336), .Z(c[82]) );
  XOR U424 ( .A(a[83]), .B(b[83]), .Z(n339) );
  NAND U425 ( .A(b[82]), .B(a[82]), .Z(n338) );
  NANDN U426 ( .A(n336), .B(n335), .Z(n337) );
  AND U427 ( .A(n338), .B(n337), .Z(n340) );
  XNOR U428 ( .A(n339), .B(n340), .Z(c[83]) );
  XOR U429 ( .A(a[84]), .B(b[84]), .Z(n343) );
  NAND U430 ( .A(b[83]), .B(a[83]), .Z(n342) );
  NANDN U431 ( .A(n340), .B(n339), .Z(n341) );
  AND U432 ( .A(n342), .B(n341), .Z(n344) );
  XNOR U433 ( .A(n343), .B(n344), .Z(c[84]) );
  XOR U434 ( .A(a[85]), .B(b[85]), .Z(n347) );
  NAND U435 ( .A(b[84]), .B(a[84]), .Z(n346) );
  NANDN U436 ( .A(n344), .B(n343), .Z(n345) );
  AND U437 ( .A(n346), .B(n345), .Z(n348) );
  XNOR U438 ( .A(n347), .B(n348), .Z(c[85]) );
  XOR U439 ( .A(a[86]), .B(b[86]), .Z(n351) );
  NAND U440 ( .A(b[85]), .B(a[85]), .Z(n350) );
  NANDN U441 ( .A(n348), .B(n347), .Z(n349) );
  AND U442 ( .A(n350), .B(n349), .Z(n352) );
  XNOR U443 ( .A(n351), .B(n352), .Z(c[86]) );
  XOR U444 ( .A(a[87]), .B(b[87]), .Z(n355) );
  NAND U445 ( .A(b[86]), .B(a[86]), .Z(n354) );
  NANDN U446 ( .A(n352), .B(n351), .Z(n353) );
  AND U447 ( .A(n354), .B(n353), .Z(n356) );
  XNOR U448 ( .A(n355), .B(n356), .Z(c[87]) );
  XOR U449 ( .A(a[88]), .B(b[88]), .Z(n359) );
  NAND U450 ( .A(b[87]), .B(a[87]), .Z(n358) );
  NANDN U451 ( .A(n356), .B(n355), .Z(n357) );
  AND U452 ( .A(n358), .B(n357), .Z(n360) );
  XNOR U453 ( .A(n359), .B(n360), .Z(c[88]) );
  XOR U454 ( .A(a[89]), .B(b[89]), .Z(n363) );
  NAND U455 ( .A(b[88]), .B(a[88]), .Z(n362) );
  NANDN U456 ( .A(n360), .B(n359), .Z(n361) );
  AND U457 ( .A(n362), .B(n361), .Z(n364) );
  XNOR U458 ( .A(n363), .B(n364), .Z(c[89]) );
  XOR U459 ( .A(a[90]), .B(b[90]), .Z(n367) );
  NAND U460 ( .A(b[89]), .B(a[89]), .Z(n366) );
  NANDN U461 ( .A(n364), .B(n363), .Z(n365) );
  AND U462 ( .A(n366), .B(n365), .Z(n368) );
  XNOR U463 ( .A(n367), .B(n368), .Z(c[90]) );
  XOR U464 ( .A(a[91]), .B(b[91]), .Z(n371) );
  NAND U465 ( .A(b[90]), .B(a[90]), .Z(n370) );
  NANDN U466 ( .A(n368), .B(n367), .Z(n369) );
  AND U467 ( .A(n370), .B(n369), .Z(n372) );
  XNOR U468 ( .A(n371), .B(n372), .Z(c[91]) );
  XOR U469 ( .A(a[92]), .B(b[92]), .Z(n375) );
  NAND U470 ( .A(b[91]), .B(a[91]), .Z(n374) );
  NANDN U471 ( .A(n372), .B(n371), .Z(n373) );
  AND U472 ( .A(n374), .B(n373), .Z(n376) );
  XNOR U473 ( .A(n375), .B(n376), .Z(c[92]) );
  XOR U474 ( .A(a[93]), .B(b[93]), .Z(n379) );
  NAND U475 ( .A(b[92]), .B(a[92]), .Z(n378) );
  NANDN U476 ( .A(n376), .B(n375), .Z(n377) );
  AND U477 ( .A(n378), .B(n377), .Z(n380) );
  XNOR U478 ( .A(n379), .B(n380), .Z(c[93]) );
  XOR U479 ( .A(a[94]), .B(b[94]), .Z(n383) );
  NAND U480 ( .A(b[93]), .B(a[93]), .Z(n382) );
  NANDN U481 ( .A(n380), .B(n379), .Z(n381) );
  AND U482 ( .A(n382), .B(n381), .Z(n384) );
  XNOR U483 ( .A(n383), .B(n384), .Z(c[94]) );
  XOR U484 ( .A(a[95]), .B(b[95]), .Z(n387) );
  NAND U485 ( .A(b[94]), .B(a[94]), .Z(n386) );
  NANDN U486 ( .A(n384), .B(n383), .Z(n385) );
  AND U487 ( .A(n386), .B(n385), .Z(n388) );
  XNOR U488 ( .A(n387), .B(n388), .Z(c[95]) );
  XOR U489 ( .A(a[96]), .B(b[96]), .Z(n391) );
  NAND U490 ( .A(b[95]), .B(a[95]), .Z(n390) );
  NANDN U491 ( .A(n388), .B(n387), .Z(n389) );
  AND U492 ( .A(n390), .B(n389), .Z(n392) );
  XNOR U493 ( .A(n391), .B(n392), .Z(c[96]) );
  XOR U494 ( .A(a[97]), .B(b[97]), .Z(n395) );
  NAND U495 ( .A(b[96]), .B(a[96]), .Z(n394) );
  NANDN U496 ( .A(n392), .B(n391), .Z(n393) );
  AND U497 ( .A(n394), .B(n393), .Z(n396) );
  XNOR U498 ( .A(n395), .B(n396), .Z(c[97]) );
  XOR U499 ( .A(a[98]), .B(b[98]), .Z(n399) );
  NAND U500 ( .A(b[97]), .B(a[97]), .Z(n398) );
  NANDN U501 ( .A(n396), .B(n395), .Z(n397) );
  AND U502 ( .A(n398), .B(n397), .Z(n400) );
  XNOR U503 ( .A(n399), .B(n400), .Z(c[98]) );
  XOR U504 ( .A(a[99]), .B(b[99]), .Z(n403) );
  NAND U505 ( .A(b[98]), .B(a[98]), .Z(n402) );
  NANDN U506 ( .A(n400), .B(n399), .Z(n401) );
  AND U507 ( .A(n402), .B(n401), .Z(n404) );
  XNOR U508 ( .A(n403), .B(n404), .Z(c[99]) );
  XOR U509 ( .A(a[100]), .B(b[100]), .Z(n407) );
  NAND U510 ( .A(b[99]), .B(a[99]), .Z(n406) );
  NANDN U511 ( .A(n404), .B(n403), .Z(n405) );
  AND U512 ( .A(n406), .B(n405), .Z(n408) );
  XNOR U513 ( .A(n407), .B(n408), .Z(c[100]) );
  NAND U514 ( .A(b[100]), .B(a[100]), .Z(n410) );
  NANDN U515 ( .A(n408), .B(n407), .Z(n409) );
  NAND U516 ( .A(n410), .B(n409), .Z(n412) );
  XNOR U517 ( .A(b[101]), .B(a[101]), .Z(n411) );
  XNOR U518 ( .A(n412), .B(n411), .Z(c[101]) );
  XNOR U519 ( .A(b[102]), .B(a[102]), .Z(n416) );
  OR U520 ( .A(b[101]), .B(a[101]), .Z(n414) );
  OR U521 ( .A(n412), .B(n411), .Z(n413) );
  AND U522 ( .A(n414), .B(n413), .Z(n415) );
  XNOR U523 ( .A(n416), .B(n415), .Z(c[102]) );
  XNOR U524 ( .A(b[103]), .B(a[103]), .Z(n420) );
  OR U525 ( .A(b[102]), .B(a[102]), .Z(n418) );
  OR U526 ( .A(n416), .B(n415), .Z(n417) );
  AND U527 ( .A(n418), .B(n417), .Z(n419) );
  XNOR U528 ( .A(n420), .B(n419), .Z(c[103]) );
  XNOR U529 ( .A(b[104]), .B(a[104]), .Z(n424) );
  OR U530 ( .A(b[103]), .B(a[103]), .Z(n422) );
  OR U531 ( .A(n420), .B(n419), .Z(n421) );
  AND U532 ( .A(n422), .B(n421), .Z(n423) );
  XNOR U533 ( .A(n424), .B(n423), .Z(c[104]) );
  XNOR U534 ( .A(b[105]), .B(a[105]), .Z(n428) );
  OR U535 ( .A(b[104]), .B(a[104]), .Z(n426) );
  OR U536 ( .A(n424), .B(n423), .Z(n425) );
  AND U537 ( .A(n426), .B(n425), .Z(n427) );
  XNOR U538 ( .A(n428), .B(n427), .Z(c[105]) );
  XNOR U539 ( .A(b[106]), .B(a[106]), .Z(n432) );
  OR U540 ( .A(b[105]), .B(a[105]), .Z(n430) );
  OR U541 ( .A(n428), .B(n427), .Z(n429) );
  AND U542 ( .A(n430), .B(n429), .Z(n431) );
  XNOR U543 ( .A(n432), .B(n431), .Z(c[106]) );
  XNOR U544 ( .A(b[107]), .B(a[107]), .Z(n436) );
  OR U545 ( .A(b[106]), .B(a[106]), .Z(n434) );
  OR U546 ( .A(n432), .B(n431), .Z(n433) );
  AND U547 ( .A(n434), .B(n433), .Z(n435) );
  XNOR U548 ( .A(n436), .B(n435), .Z(c[107]) );
  XNOR U549 ( .A(b[108]), .B(a[108]), .Z(n440) );
  OR U550 ( .A(b[107]), .B(a[107]), .Z(n438) );
  OR U551 ( .A(n436), .B(n435), .Z(n437) );
  AND U552 ( .A(n438), .B(n437), .Z(n439) );
  XNOR U553 ( .A(n440), .B(n439), .Z(c[108]) );
  XNOR U554 ( .A(b[109]), .B(a[109]), .Z(n444) );
  OR U555 ( .A(b[108]), .B(a[108]), .Z(n442) );
  OR U556 ( .A(n440), .B(n439), .Z(n441) );
  AND U557 ( .A(n442), .B(n441), .Z(n443) );
  XNOR U558 ( .A(n444), .B(n443), .Z(c[109]) );
  XNOR U559 ( .A(b[110]), .B(a[110]), .Z(n448) );
  OR U560 ( .A(b[109]), .B(a[109]), .Z(n446) );
  OR U561 ( .A(n444), .B(n443), .Z(n445) );
  AND U562 ( .A(n446), .B(n445), .Z(n447) );
  XNOR U563 ( .A(n448), .B(n447), .Z(c[110]) );
  XNOR U564 ( .A(b[111]), .B(a[111]), .Z(n452) );
  OR U565 ( .A(b[110]), .B(a[110]), .Z(n450) );
  OR U566 ( .A(n448), .B(n447), .Z(n449) );
  AND U567 ( .A(n450), .B(n449), .Z(n451) );
  XNOR U568 ( .A(n452), .B(n451), .Z(c[111]) );
  XNOR U569 ( .A(b[112]), .B(a[112]), .Z(n456) );
  OR U570 ( .A(b[111]), .B(a[111]), .Z(n454) );
  OR U571 ( .A(n452), .B(n451), .Z(n453) );
  AND U572 ( .A(n454), .B(n453), .Z(n455) );
  XNOR U573 ( .A(n456), .B(n455), .Z(c[112]) );
  XNOR U574 ( .A(b[113]), .B(a[113]), .Z(n460) );
  OR U575 ( .A(b[112]), .B(a[112]), .Z(n458) );
  OR U576 ( .A(n456), .B(n455), .Z(n457) );
  AND U577 ( .A(n458), .B(n457), .Z(n459) );
  XNOR U578 ( .A(n460), .B(n459), .Z(c[113]) );
  XNOR U579 ( .A(b[114]), .B(a[114]), .Z(n464) );
  OR U580 ( .A(b[113]), .B(a[113]), .Z(n462) );
  OR U581 ( .A(n460), .B(n459), .Z(n461) );
  AND U582 ( .A(n462), .B(n461), .Z(n463) );
  XNOR U583 ( .A(n464), .B(n463), .Z(c[114]) );
  XNOR U584 ( .A(b[115]), .B(a[115]), .Z(n468) );
  OR U585 ( .A(b[114]), .B(a[114]), .Z(n466) );
  OR U586 ( .A(n464), .B(n463), .Z(n465) );
  AND U587 ( .A(n466), .B(n465), .Z(n467) );
  XNOR U588 ( .A(n468), .B(n467), .Z(c[115]) );
  OR U589 ( .A(b[115]), .B(a[115]), .Z(n470) );
  OR U590 ( .A(n468), .B(n467), .Z(n469) );
  NAND U591 ( .A(n470), .B(n469), .Z(n472) );
  XOR U592 ( .A(a[116]), .B(b[116]), .Z(n471) );
  XNOR U593 ( .A(n472), .B(n471), .Z(c[116]) );
  XOR U594 ( .A(a[117]), .B(b[117]), .Z(n475) );
  NAND U595 ( .A(b[116]), .B(a[116]), .Z(n474) );
  NANDN U596 ( .A(n472), .B(n471), .Z(n473) );
  AND U597 ( .A(n474), .B(n473), .Z(n476) );
  XNOR U598 ( .A(n475), .B(n476), .Z(c[117]) );
  XOR U599 ( .A(a[118]), .B(b[118]), .Z(n479) );
  NAND U600 ( .A(b[117]), .B(a[117]), .Z(n478) );
  NANDN U601 ( .A(n476), .B(n475), .Z(n477) );
  AND U602 ( .A(n478), .B(n477), .Z(n480) );
  XNOR U603 ( .A(n479), .B(n480), .Z(c[118]) );
  XOR U604 ( .A(a[119]), .B(b[119]), .Z(n483) );
  NAND U605 ( .A(b[118]), .B(a[118]), .Z(n482) );
  NANDN U606 ( .A(n480), .B(n479), .Z(n481) );
  AND U607 ( .A(n482), .B(n481), .Z(n484) );
  XNOR U608 ( .A(n483), .B(n484), .Z(c[119]) );
  XOR U609 ( .A(a[120]), .B(b[120]), .Z(n487) );
  NAND U610 ( .A(b[119]), .B(a[119]), .Z(n486) );
  NANDN U611 ( .A(n484), .B(n483), .Z(n485) );
  AND U612 ( .A(n486), .B(n485), .Z(n488) );
  XNOR U613 ( .A(n487), .B(n488), .Z(c[120]) );
  XOR U614 ( .A(a[121]), .B(b[121]), .Z(n491) );
  NAND U615 ( .A(b[120]), .B(a[120]), .Z(n490) );
  NANDN U616 ( .A(n488), .B(n487), .Z(n489) );
  AND U617 ( .A(n490), .B(n489), .Z(n492) );
  XNOR U618 ( .A(n491), .B(n492), .Z(c[121]) );
  XOR U619 ( .A(a[122]), .B(b[122]), .Z(n495) );
  NAND U620 ( .A(b[121]), .B(a[121]), .Z(n494) );
  NANDN U621 ( .A(n492), .B(n491), .Z(n493) );
  AND U622 ( .A(n494), .B(n493), .Z(n496) );
  XNOR U623 ( .A(n495), .B(n496), .Z(c[122]) );
  XOR U624 ( .A(a[123]), .B(b[123]), .Z(n499) );
  NAND U625 ( .A(b[122]), .B(a[122]), .Z(n498) );
  NANDN U626 ( .A(n496), .B(n495), .Z(n497) );
  AND U627 ( .A(n498), .B(n497), .Z(n500) );
  XNOR U628 ( .A(n499), .B(n500), .Z(c[123]) );
  XOR U629 ( .A(a[124]), .B(b[124]), .Z(n503) );
  NAND U630 ( .A(b[123]), .B(a[123]), .Z(n502) );
  NANDN U631 ( .A(n500), .B(n499), .Z(n501) );
  AND U632 ( .A(n502), .B(n501), .Z(n504) );
  XNOR U633 ( .A(n503), .B(n504), .Z(c[124]) );
  XOR U634 ( .A(a[125]), .B(b[125]), .Z(n507) );
  NAND U635 ( .A(b[124]), .B(a[124]), .Z(n506) );
  NANDN U636 ( .A(n504), .B(n503), .Z(n505) );
  AND U637 ( .A(n506), .B(n505), .Z(n508) );
  XNOR U638 ( .A(n507), .B(n508), .Z(c[125]) );
  XOR U639 ( .A(a[126]), .B(b[126]), .Z(n511) );
  NAND U640 ( .A(b[125]), .B(a[125]), .Z(n510) );
  NANDN U641 ( .A(n508), .B(n507), .Z(n509) );
  AND U642 ( .A(n510), .B(n509), .Z(n512) );
  XNOR U643 ( .A(n511), .B(n512), .Z(c[126]) );
  XOR U644 ( .A(a[127]), .B(b[127]), .Z(n515) );
  NAND U645 ( .A(b[126]), .B(a[126]), .Z(n514) );
  NANDN U646 ( .A(n512), .B(n511), .Z(n513) );
  AND U647 ( .A(n514), .B(n513), .Z(n516) );
  XNOR U648 ( .A(n515), .B(n516), .Z(c[127]) );
  XOR U649 ( .A(a[128]), .B(b[128]), .Z(n519) );
  NAND U650 ( .A(b[127]), .B(a[127]), .Z(n518) );
  NANDN U651 ( .A(n516), .B(n515), .Z(n517) );
  AND U652 ( .A(n518), .B(n517), .Z(n520) );
  XNOR U653 ( .A(n519), .B(n520), .Z(c[128]) );
  XOR U654 ( .A(a[129]), .B(b[129]), .Z(n523) );
  NAND U655 ( .A(b[128]), .B(a[128]), .Z(n522) );
  NANDN U656 ( .A(n520), .B(n519), .Z(n521) );
  AND U657 ( .A(n522), .B(n521), .Z(n524) );
  XNOR U658 ( .A(n523), .B(n524), .Z(c[129]) );
  XOR U659 ( .A(a[130]), .B(b[130]), .Z(n527) );
  NAND U660 ( .A(b[129]), .B(a[129]), .Z(n526) );
  NANDN U661 ( .A(n524), .B(n523), .Z(n525) );
  AND U662 ( .A(n526), .B(n525), .Z(n528) );
  XNOR U663 ( .A(n527), .B(n528), .Z(c[130]) );
  XOR U664 ( .A(a[131]), .B(b[131]), .Z(n531) );
  NAND U665 ( .A(b[130]), .B(a[130]), .Z(n530) );
  NANDN U666 ( .A(n528), .B(n527), .Z(n529) );
  AND U667 ( .A(n530), .B(n529), .Z(n532) );
  XNOR U668 ( .A(n531), .B(n532), .Z(c[131]) );
  XOR U669 ( .A(a[132]), .B(b[132]), .Z(n535) );
  NAND U670 ( .A(b[131]), .B(a[131]), .Z(n534) );
  NANDN U671 ( .A(n532), .B(n531), .Z(n533) );
  AND U672 ( .A(n534), .B(n533), .Z(n536) );
  XNOR U673 ( .A(n535), .B(n536), .Z(c[132]) );
  XOR U674 ( .A(a[133]), .B(b[133]), .Z(n539) );
  NAND U675 ( .A(b[132]), .B(a[132]), .Z(n538) );
  NANDN U676 ( .A(n536), .B(n535), .Z(n537) );
  AND U677 ( .A(n538), .B(n537), .Z(n540) );
  XNOR U678 ( .A(n539), .B(n540), .Z(c[133]) );
  XOR U679 ( .A(a[134]), .B(b[134]), .Z(n543) );
  NAND U680 ( .A(b[133]), .B(a[133]), .Z(n542) );
  NANDN U681 ( .A(n540), .B(n539), .Z(n541) );
  AND U682 ( .A(n542), .B(n541), .Z(n544) );
  XNOR U683 ( .A(n543), .B(n544), .Z(c[134]) );
  XOR U684 ( .A(a[135]), .B(b[135]), .Z(n547) );
  NAND U685 ( .A(b[134]), .B(a[134]), .Z(n546) );
  NANDN U686 ( .A(n544), .B(n543), .Z(n545) );
  AND U687 ( .A(n546), .B(n545), .Z(n548) );
  XNOR U688 ( .A(n547), .B(n548), .Z(c[135]) );
  XOR U689 ( .A(a[136]), .B(b[136]), .Z(n551) );
  NAND U690 ( .A(b[135]), .B(a[135]), .Z(n550) );
  NANDN U691 ( .A(n548), .B(n547), .Z(n549) );
  AND U692 ( .A(n550), .B(n549), .Z(n552) );
  XNOR U693 ( .A(n551), .B(n552), .Z(c[136]) );
  XOR U694 ( .A(a[137]), .B(b[137]), .Z(n555) );
  NAND U695 ( .A(b[136]), .B(a[136]), .Z(n554) );
  NANDN U696 ( .A(n552), .B(n551), .Z(n553) );
  AND U697 ( .A(n554), .B(n553), .Z(n556) );
  XNOR U698 ( .A(n555), .B(n556), .Z(c[137]) );
  XOR U699 ( .A(a[138]), .B(b[138]), .Z(n559) );
  NAND U700 ( .A(b[137]), .B(a[137]), .Z(n558) );
  NANDN U701 ( .A(n556), .B(n555), .Z(n557) );
  AND U702 ( .A(n558), .B(n557), .Z(n560) );
  XNOR U703 ( .A(n559), .B(n560), .Z(c[138]) );
  XOR U704 ( .A(a[139]), .B(b[139]), .Z(n563) );
  NAND U705 ( .A(b[138]), .B(a[138]), .Z(n562) );
  NANDN U706 ( .A(n560), .B(n559), .Z(n561) );
  AND U707 ( .A(n562), .B(n561), .Z(n564) );
  XNOR U708 ( .A(n563), .B(n564), .Z(c[139]) );
  XOR U709 ( .A(a[140]), .B(b[140]), .Z(n567) );
  NAND U710 ( .A(b[139]), .B(a[139]), .Z(n566) );
  NANDN U711 ( .A(n564), .B(n563), .Z(n565) );
  AND U712 ( .A(n566), .B(n565), .Z(n568) );
  XNOR U713 ( .A(n567), .B(n568), .Z(c[140]) );
  XOR U714 ( .A(a[141]), .B(b[141]), .Z(n571) );
  NAND U715 ( .A(b[140]), .B(a[140]), .Z(n570) );
  NANDN U716 ( .A(n568), .B(n567), .Z(n569) );
  AND U717 ( .A(n570), .B(n569), .Z(n572) );
  XNOR U718 ( .A(n571), .B(n572), .Z(c[141]) );
  XOR U719 ( .A(a[142]), .B(b[142]), .Z(n575) );
  NAND U720 ( .A(b[141]), .B(a[141]), .Z(n574) );
  NANDN U721 ( .A(n572), .B(n571), .Z(n573) );
  AND U722 ( .A(n574), .B(n573), .Z(n576) );
  XNOR U723 ( .A(n575), .B(n576), .Z(c[142]) );
  XOR U724 ( .A(a[143]), .B(b[143]), .Z(n579) );
  NAND U725 ( .A(b[142]), .B(a[142]), .Z(n578) );
  NANDN U726 ( .A(n576), .B(n575), .Z(n577) );
  AND U727 ( .A(n578), .B(n577), .Z(n580) );
  XNOR U728 ( .A(n579), .B(n580), .Z(c[143]) );
  XOR U729 ( .A(a[144]), .B(b[144]), .Z(n583) );
  NAND U730 ( .A(b[143]), .B(a[143]), .Z(n582) );
  NANDN U731 ( .A(n580), .B(n579), .Z(n581) );
  AND U732 ( .A(n582), .B(n581), .Z(n584) );
  XNOR U733 ( .A(n583), .B(n584), .Z(c[144]) );
  XOR U734 ( .A(a[145]), .B(b[145]), .Z(n587) );
  NAND U735 ( .A(b[144]), .B(a[144]), .Z(n586) );
  NANDN U736 ( .A(n584), .B(n583), .Z(n585) );
  AND U737 ( .A(n586), .B(n585), .Z(n588) );
  XNOR U738 ( .A(n587), .B(n588), .Z(c[145]) );
  XOR U739 ( .A(a[146]), .B(b[146]), .Z(n591) );
  NAND U740 ( .A(b[145]), .B(a[145]), .Z(n590) );
  NANDN U741 ( .A(n588), .B(n587), .Z(n589) );
  AND U742 ( .A(n590), .B(n589), .Z(n592) );
  XNOR U743 ( .A(n591), .B(n592), .Z(c[146]) );
  XOR U744 ( .A(a[147]), .B(b[147]), .Z(n595) );
  NAND U745 ( .A(b[146]), .B(a[146]), .Z(n594) );
  NANDN U746 ( .A(n592), .B(n591), .Z(n593) );
  AND U747 ( .A(n594), .B(n593), .Z(n596) );
  XNOR U748 ( .A(n595), .B(n596), .Z(c[147]) );
  XOR U749 ( .A(a[148]), .B(b[148]), .Z(n599) );
  NAND U750 ( .A(b[147]), .B(a[147]), .Z(n598) );
  NANDN U751 ( .A(n596), .B(n595), .Z(n597) );
  AND U752 ( .A(n598), .B(n597), .Z(n600) );
  XNOR U753 ( .A(n599), .B(n600), .Z(c[148]) );
  XOR U754 ( .A(a[149]), .B(b[149]), .Z(n603) );
  NAND U755 ( .A(b[148]), .B(a[148]), .Z(n602) );
  NANDN U756 ( .A(n600), .B(n599), .Z(n601) );
  AND U757 ( .A(n602), .B(n601), .Z(n604) );
  XNOR U758 ( .A(n603), .B(n604), .Z(c[149]) );
  XOR U759 ( .A(a[150]), .B(b[150]), .Z(n607) );
  NAND U760 ( .A(b[149]), .B(a[149]), .Z(n606) );
  NANDN U761 ( .A(n604), .B(n603), .Z(n605) );
  AND U762 ( .A(n606), .B(n605), .Z(n608) );
  XNOR U763 ( .A(n607), .B(n608), .Z(c[150]) );
  XOR U764 ( .A(a[151]), .B(b[151]), .Z(n611) );
  NAND U765 ( .A(b[150]), .B(a[150]), .Z(n610) );
  NANDN U766 ( .A(n608), .B(n607), .Z(n609) );
  AND U767 ( .A(n610), .B(n609), .Z(n612) );
  XNOR U768 ( .A(n611), .B(n612), .Z(c[151]) );
  NAND U769 ( .A(b[151]), .B(a[151]), .Z(n614) );
  NANDN U770 ( .A(n612), .B(n611), .Z(n613) );
  NAND U771 ( .A(n614), .B(n613), .Z(n616) );
  XNOR U772 ( .A(b[152]), .B(a[152]), .Z(n615) );
  XNOR U773 ( .A(n616), .B(n615), .Z(c[152]) );
  XNOR U774 ( .A(b[153]), .B(a[153]), .Z(n620) );
  OR U775 ( .A(b[152]), .B(a[152]), .Z(n618) );
  OR U776 ( .A(n616), .B(n615), .Z(n617) );
  AND U777 ( .A(n618), .B(n617), .Z(n619) );
  XNOR U778 ( .A(n620), .B(n619), .Z(c[153]) );
  XNOR U779 ( .A(b[154]), .B(a[154]), .Z(n624) );
  OR U780 ( .A(b[153]), .B(a[153]), .Z(n622) );
  OR U781 ( .A(n620), .B(n619), .Z(n621) );
  AND U782 ( .A(n622), .B(n621), .Z(n623) );
  XNOR U783 ( .A(n624), .B(n623), .Z(c[154]) );
  XNOR U784 ( .A(b[155]), .B(a[155]), .Z(n628) );
  OR U785 ( .A(b[154]), .B(a[154]), .Z(n626) );
  OR U786 ( .A(n624), .B(n623), .Z(n625) );
  AND U787 ( .A(n626), .B(n625), .Z(n627) );
  XNOR U788 ( .A(n628), .B(n627), .Z(c[155]) );
  XNOR U789 ( .A(b[156]), .B(a[156]), .Z(n632) );
  OR U790 ( .A(b[155]), .B(a[155]), .Z(n630) );
  OR U791 ( .A(n628), .B(n627), .Z(n629) );
  AND U792 ( .A(n630), .B(n629), .Z(n631) );
  XNOR U793 ( .A(n632), .B(n631), .Z(c[156]) );
  XNOR U794 ( .A(b[157]), .B(a[157]), .Z(n636) );
  OR U795 ( .A(b[156]), .B(a[156]), .Z(n634) );
  OR U796 ( .A(n632), .B(n631), .Z(n633) );
  AND U797 ( .A(n634), .B(n633), .Z(n635) );
  XNOR U798 ( .A(n636), .B(n635), .Z(c[157]) );
  XNOR U799 ( .A(b[158]), .B(a[158]), .Z(n640) );
  OR U800 ( .A(b[157]), .B(a[157]), .Z(n638) );
  OR U801 ( .A(n636), .B(n635), .Z(n637) );
  AND U802 ( .A(n638), .B(n637), .Z(n639) );
  XNOR U803 ( .A(n640), .B(n639), .Z(c[158]) );
  OR U804 ( .A(b[158]), .B(a[158]), .Z(n642) );
  OR U805 ( .A(n640), .B(n639), .Z(n641) );
  NAND U806 ( .A(n642), .B(n641), .Z(n644) );
  XOR U807 ( .A(a[159]), .B(b[159]), .Z(n643) );
  XNOR U808 ( .A(n644), .B(n643), .Z(c[159]) );
  XOR U809 ( .A(a[160]), .B(b[160]), .Z(n647) );
  NAND U810 ( .A(b[159]), .B(a[159]), .Z(n646) );
  NANDN U811 ( .A(n644), .B(n643), .Z(n645) );
  AND U812 ( .A(n646), .B(n645), .Z(n648) );
  XNOR U813 ( .A(n647), .B(n648), .Z(c[160]) );
  XOR U814 ( .A(a[161]), .B(b[161]), .Z(n651) );
  NAND U815 ( .A(b[160]), .B(a[160]), .Z(n650) );
  NANDN U816 ( .A(n648), .B(n647), .Z(n649) );
  AND U817 ( .A(n650), .B(n649), .Z(n652) );
  XNOR U818 ( .A(n651), .B(n652), .Z(c[161]) );
  XOR U819 ( .A(a[162]), .B(b[162]), .Z(n655) );
  NAND U820 ( .A(b[161]), .B(a[161]), .Z(n654) );
  NANDN U821 ( .A(n652), .B(n651), .Z(n653) );
  AND U822 ( .A(n654), .B(n653), .Z(n656) );
  XNOR U823 ( .A(n655), .B(n656), .Z(c[162]) );
  XOR U824 ( .A(a[163]), .B(b[163]), .Z(n659) );
  NAND U825 ( .A(b[162]), .B(a[162]), .Z(n658) );
  NANDN U826 ( .A(n656), .B(n655), .Z(n657) );
  AND U827 ( .A(n658), .B(n657), .Z(n660) );
  XNOR U828 ( .A(n659), .B(n660), .Z(c[163]) );
  XOR U829 ( .A(a[164]), .B(b[164]), .Z(n663) );
  NAND U830 ( .A(b[163]), .B(a[163]), .Z(n662) );
  NANDN U831 ( .A(n660), .B(n659), .Z(n661) );
  AND U832 ( .A(n662), .B(n661), .Z(n664) );
  XNOR U833 ( .A(n663), .B(n664), .Z(c[164]) );
  XOR U834 ( .A(a[165]), .B(b[165]), .Z(n667) );
  NAND U835 ( .A(b[164]), .B(a[164]), .Z(n666) );
  NANDN U836 ( .A(n664), .B(n663), .Z(n665) );
  AND U837 ( .A(n666), .B(n665), .Z(n668) );
  XNOR U838 ( .A(n667), .B(n668), .Z(c[165]) );
  XOR U839 ( .A(a[166]), .B(b[166]), .Z(n671) );
  NAND U840 ( .A(b[165]), .B(a[165]), .Z(n670) );
  NANDN U841 ( .A(n668), .B(n667), .Z(n669) );
  AND U842 ( .A(n670), .B(n669), .Z(n672) );
  XNOR U843 ( .A(n671), .B(n672), .Z(c[166]) );
  XOR U844 ( .A(a[167]), .B(b[167]), .Z(n675) );
  NAND U845 ( .A(b[166]), .B(a[166]), .Z(n674) );
  NANDN U846 ( .A(n672), .B(n671), .Z(n673) );
  AND U847 ( .A(n674), .B(n673), .Z(n676) );
  XNOR U848 ( .A(n675), .B(n676), .Z(c[167]) );
  XOR U849 ( .A(a[168]), .B(b[168]), .Z(n679) );
  NAND U850 ( .A(b[167]), .B(a[167]), .Z(n678) );
  NANDN U851 ( .A(n676), .B(n675), .Z(n677) );
  AND U852 ( .A(n678), .B(n677), .Z(n680) );
  XNOR U853 ( .A(n679), .B(n680), .Z(c[168]) );
  XOR U854 ( .A(a[169]), .B(b[169]), .Z(n683) );
  NAND U855 ( .A(b[168]), .B(a[168]), .Z(n682) );
  NANDN U856 ( .A(n680), .B(n679), .Z(n681) );
  AND U857 ( .A(n682), .B(n681), .Z(n684) );
  XNOR U858 ( .A(n683), .B(n684), .Z(c[169]) );
  XOR U859 ( .A(a[170]), .B(b[170]), .Z(n687) );
  NAND U860 ( .A(b[169]), .B(a[169]), .Z(n686) );
  NANDN U861 ( .A(n684), .B(n683), .Z(n685) );
  AND U862 ( .A(n686), .B(n685), .Z(n688) );
  XNOR U863 ( .A(n687), .B(n688), .Z(c[170]) );
  XOR U864 ( .A(a[171]), .B(b[171]), .Z(n691) );
  NAND U865 ( .A(b[170]), .B(a[170]), .Z(n690) );
  NANDN U866 ( .A(n688), .B(n687), .Z(n689) );
  AND U867 ( .A(n690), .B(n689), .Z(n692) );
  XNOR U868 ( .A(n691), .B(n692), .Z(c[171]) );
  XOR U869 ( .A(a[172]), .B(b[172]), .Z(n695) );
  NAND U870 ( .A(b[171]), .B(a[171]), .Z(n694) );
  NANDN U871 ( .A(n692), .B(n691), .Z(n693) );
  AND U872 ( .A(n694), .B(n693), .Z(n696) );
  XNOR U873 ( .A(n695), .B(n696), .Z(c[172]) );
  XOR U874 ( .A(a[173]), .B(b[173]), .Z(n699) );
  NAND U875 ( .A(b[172]), .B(a[172]), .Z(n698) );
  NANDN U876 ( .A(n696), .B(n695), .Z(n697) );
  AND U877 ( .A(n698), .B(n697), .Z(n700) );
  XNOR U878 ( .A(n699), .B(n700), .Z(c[173]) );
  XOR U879 ( .A(a[174]), .B(b[174]), .Z(n703) );
  NAND U880 ( .A(b[173]), .B(a[173]), .Z(n702) );
  NANDN U881 ( .A(n700), .B(n699), .Z(n701) );
  AND U882 ( .A(n702), .B(n701), .Z(n704) );
  XNOR U883 ( .A(n703), .B(n704), .Z(c[174]) );
  XOR U884 ( .A(a[175]), .B(b[175]), .Z(n707) );
  NAND U885 ( .A(b[174]), .B(a[174]), .Z(n706) );
  NANDN U886 ( .A(n704), .B(n703), .Z(n705) );
  AND U887 ( .A(n706), .B(n705), .Z(n708) );
  XNOR U888 ( .A(n707), .B(n708), .Z(c[175]) );
  XOR U889 ( .A(a[176]), .B(b[176]), .Z(n711) );
  NAND U890 ( .A(b[175]), .B(a[175]), .Z(n710) );
  NANDN U891 ( .A(n708), .B(n707), .Z(n709) );
  AND U892 ( .A(n710), .B(n709), .Z(n712) );
  XNOR U893 ( .A(n711), .B(n712), .Z(c[176]) );
  XOR U894 ( .A(a[177]), .B(b[177]), .Z(n715) );
  NAND U895 ( .A(b[176]), .B(a[176]), .Z(n714) );
  NANDN U896 ( .A(n712), .B(n711), .Z(n713) );
  AND U897 ( .A(n714), .B(n713), .Z(n716) );
  XNOR U898 ( .A(n715), .B(n716), .Z(c[177]) );
  XOR U899 ( .A(a[178]), .B(b[178]), .Z(n719) );
  NAND U900 ( .A(b[177]), .B(a[177]), .Z(n718) );
  NANDN U901 ( .A(n716), .B(n715), .Z(n717) );
  AND U902 ( .A(n718), .B(n717), .Z(n720) );
  XNOR U903 ( .A(n719), .B(n720), .Z(c[178]) );
  XOR U904 ( .A(a[179]), .B(b[179]), .Z(n723) );
  NAND U905 ( .A(b[178]), .B(a[178]), .Z(n722) );
  NANDN U906 ( .A(n720), .B(n719), .Z(n721) );
  AND U907 ( .A(n722), .B(n721), .Z(n724) );
  XNOR U908 ( .A(n723), .B(n724), .Z(c[179]) );
  XOR U909 ( .A(a[180]), .B(b[180]), .Z(n727) );
  NAND U910 ( .A(b[179]), .B(a[179]), .Z(n726) );
  NANDN U911 ( .A(n724), .B(n723), .Z(n725) );
  AND U912 ( .A(n726), .B(n725), .Z(n728) );
  XNOR U913 ( .A(n727), .B(n728), .Z(c[180]) );
  XOR U914 ( .A(a[181]), .B(b[181]), .Z(n731) );
  NAND U915 ( .A(b[180]), .B(a[180]), .Z(n730) );
  NANDN U916 ( .A(n728), .B(n727), .Z(n729) );
  AND U917 ( .A(n730), .B(n729), .Z(n732) );
  XNOR U918 ( .A(n731), .B(n732), .Z(c[181]) );
  XOR U919 ( .A(a[182]), .B(b[182]), .Z(n735) );
  NAND U920 ( .A(b[181]), .B(a[181]), .Z(n734) );
  NANDN U921 ( .A(n732), .B(n731), .Z(n733) );
  AND U922 ( .A(n734), .B(n733), .Z(n736) );
  XNOR U923 ( .A(n735), .B(n736), .Z(c[182]) );
  XOR U924 ( .A(a[183]), .B(b[183]), .Z(n739) );
  NAND U925 ( .A(b[182]), .B(a[182]), .Z(n738) );
  NANDN U926 ( .A(n736), .B(n735), .Z(n737) );
  AND U927 ( .A(n738), .B(n737), .Z(n740) );
  XNOR U928 ( .A(n739), .B(n740), .Z(c[183]) );
  NAND U929 ( .A(b[183]), .B(a[183]), .Z(n742) );
  NANDN U930 ( .A(n740), .B(n739), .Z(n741) );
  NAND U931 ( .A(n742), .B(n741), .Z(n744) );
  XNOR U932 ( .A(b[184]), .B(a[184]), .Z(n743) );
  XNOR U933 ( .A(n744), .B(n743), .Z(c[184]) );
  XOR U934 ( .A(a[185]), .B(b[185]), .Z(n747) );
  OR U935 ( .A(b[184]), .B(a[184]), .Z(n746) );
  OR U936 ( .A(n744), .B(n743), .Z(n745) );
  NAND U937 ( .A(n746), .B(n745), .Z(n748) );
  XNOR U938 ( .A(n747), .B(n748), .Z(c[185]) );
  NAND U939 ( .A(b[185]), .B(a[185]), .Z(n750) );
  NANDN U940 ( .A(n748), .B(n747), .Z(n749) );
  NAND U941 ( .A(n750), .B(n749), .Z(n752) );
  XNOR U942 ( .A(b[186]), .B(a[186]), .Z(n751) );
  XNOR U943 ( .A(n752), .B(n751), .Z(c[186]) );
  XNOR U944 ( .A(b[187]), .B(a[187]), .Z(n756) );
  OR U945 ( .A(b[186]), .B(a[186]), .Z(n754) );
  OR U946 ( .A(n752), .B(n751), .Z(n753) );
  AND U947 ( .A(n754), .B(n753), .Z(n755) );
  XNOR U948 ( .A(n756), .B(n755), .Z(c[187]) );
  XNOR U949 ( .A(b[188]), .B(a[188]), .Z(n760) );
  OR U950 ( .A(b[187]), .B(a[187]), .Z(n758) );
  OR U951 ( .A(n756), .B(n755), .Z(n757) );
  AND U952 ( .A(n758), .B(n757), .Z(n759) );
  XNOR U953 ( .A(n760), .B(n759), .Z(c[188]) );
  XNOR U954 ( .A(b[189]), .B(a[189]), .Z(n764) );
  OR U955 ( .A(b[188]), .B(a[188]), .Z(n762) );
  OR U956 ( .A(n760), .B(n759), .Z(n761) );
  AND U957 ( .A(n762), .B(n761), .Z(n763) );
  XNOR U958 ( .A(n764), .B(n763), .Z(c[189]) );
  XNOR U959 ( .A(b[190]), .B(a[190]), .Z(n768) );
  OR U960 ( .A(b[189]), .B(a[189]), .Z(n766) );
  OR U961 ( .A(n764), .B(n763), .Z(n765) );
  AND U962 ( .A(n766), .B(n765), .Z(n767) );
  XNOR U963 ( .A(n768), .B(n767), .Z(c[190]) );
  XNOR U964 ( .A(b[191]), .B(a[191]), .Z(n772) );
  OR U965 ( .A(b[190]), .B(a[190]), .Z(n770) );
  OR U966 ( .A(n768), .B(n767), .Z(n769) );
  AND U967 ( .A(n770), .B(n769), .Z(n771) );
  XNOR U968 ( .A(n772), .B(n771), .Z(c[191]) );
  XNOR U969 ( .A(b[192]), .B(a[192]), .Z(n776) );
  OR U970 ( .A(b[191]), .B(a[191]), .Z(n774) );
  OR U971 ( .A(n772), .B(n771), .Z(n773) );
  AND U972 ( .A(n774), .B(n773), .Z(n775) );
  XNOR U973 ( .A(n776), .B(n775), .Z(c[192]) );
  XNOR U974 ( .A(b[193]), .B(a[193]), .Z(n780) );
  OR U975 ( .A(b[192]), .B(a[192]), .Z(n778) );
  OR U976 ( .A(n776), .B(n775), .Z(n777) );
  AND U977 ( .A(n778), .B(n777), .Z(n779) );
  XNOR U978 ( .A(n780), .B(n779), .Z(c[193]) );
  XNOR U979 ( .A(b[194]), .B(a[194]), .Z(n784) );
  OR U980 ( .A(b[193]), .B(a[193]), .Z(n782) );
  OR U981 ( .A(n780), .B(n779), .Z(n781) );
  AND U982 ( .A(n782), .B(n781), .Z(n783) );
  XNOR U983 ( .A(n784), .B(n783), .Z(c[194]) );
  XNOR U984 ( .A(b[195]), .B(a[195]), .Z(n788) );
  OR U985 ( .A(b[194]), .B(a[194]), .Z(n786) );
  OR U986 ( .A(n784), .B(n783), .Z(n785) );
  AND U987 ( .A(n786), .B(n785), .Z(n787) );
  XNOR U988 ( .A(n788), .B(n787), .Z(c[195]) );
  XNOR U989 ( .A(b[196]), .B(a[196]), .Z(n792) );
  OR U990 ( .A(b[195]), .B(a[195]), .Z(n790) );
  OR U991 ( .A(n788), .B(n787), .Z(n789) );
  AND U992 ( .A(n790), .B(n789), .Z(n791) );
  XNOR U993 ( .A(n792), .B(n791), .Z(c[196]) );
  XNOR U994 ( .A(b[197]), .B(a[197]), .Z(n796) );
  OR U995 ( .A(b[196]), .B(a[196]), .Z(n794) );
  OR U996 ( .A(n792), .B(n791), .Z(n793) );
  AND U997 ( .A(n794), .B(n793), .Z(n795) );
  XNOR U998 ( .A(n796), .B(n795), .Z(c[197]) );
  XNOR U999 ( .A(b[198]), .B(a[198]), .Z(n800) );
  OR U1000 ( .A(b[197]), .B(a[197]), .Z(n798) );
  OR U1001 ( .A(n796), .B(n795), .Z(n797) );
  AND U1002 ( .A(n798), .B(n797), .Z(n799) );
  XNOR U1003 ( .A(n800), .B(n799), .Z(c[198]) );
  XNOR U1004 ( .A(b[199]), .B(a[199]), .Z(n804) );
  OR U1005 ( .A(b[198]), .B(a[198]), .Z(n802) );
  OR U1006 ( .A(n800), .B(n799), .Z(n801) );
  AND U1007 ( .A(n802), .B(n801), .Z(n803) );
  XNOR U1008 ( .A(n804), .B(n803), .Z(c[199]) );
  XNOR U1009 ( .A(b[200]), .B(a[200]), .Z(n808) );
  OR U1010 ( .A(b[199]), .B(a[199]), .Z(n806) );
  OR U1011 ( .A(n804), .B(n803), .Z(n805) );
  AND U1012 ( .A(n806), .B(n805), .Z(n807) );
  XNOR U1013 ( .A(n808), .B(n807), .Z(c[200]) );
  XNOR U1014 ( .A(b[201]), .B(a[201]), .Z(n812) );
  OR U1015 ( .A(b[200]), .B(a[200]), .Z(n810) );
  OR U1016 ( .A(n808), .B(n807), .Z(n809) );
  AND U1017 ( .A(n810), .B(n809), .Z(n811) );
  XNOR U1018 ( .A(n812), .B(n811), .Z(c[201]) );
  XNOR U1019 ( .A(b[202]), .B(a[202]), .Z(n816) );
  OR U1020 ( .A(b[201]), .B(a[201]), .Z(n814) );
  OR U1021 ( .A(n812), .B(n811), .Z(n813) );
  AND U1022 ( .A(n814), .B(n813), .Z(n815) );
  XNOR U1023 ( .A(n816), .B(n815), .Z(c[202]) );
  XNOR U1024 ( .A(b[203]), .B(a[203]), .Z(n820) );
  OR U1025 ( .A(b[202]), .B(a[202]), .Z(n818) );
  OR U1026 ( .A(n816), .B(n815), .Z(n817) );
  AND U1027 ( .A(n818), .B(n817), .Z(n819) );
  XNOR U1028 ( .A(n820), .B(n819), .Z(c[203]) );
  XNOR U1029 ( .A(b[204]), .B(a[204]), .Z(n824) );
  OR U1030 ( .A(b[203]), .B(a[203]), .Z(n822) );
  OR U1031 ( .A(n820), .B(n819), .Z(n821) );
  AND U1032 ( .A(n822), .B(n821), .Z(n823) );
  XNOR U1033 ( .A(n824), .B(n823), .Z(c[204]) );
  XNOR U1034 ( .A(b[205]), .B(a[205]), .Z(n828) );
  OR U1035 ( .A(b[204]), .B(a[204]), .Z(n826) );
  OR U1036 ( .A(n824), .B(n823), .Z(n825) );
  AND U1037 ( .A(n826), .B(n825), .Z(n827) );
  XNOR U1038 ( .A(n828), .B(n827), .Z(c[205]) );
  XOR U1039 ( .A(a[206]), .B(b[206]), .Z(n831) );
  OR U1040 ( .A(b[205]), .B(a[205]), .Z(n830) );
  OR U1041 ( .A(n828), .B(n827), .Z(n829) );
  NAND U1042 ( .A(n830), .B(n829), .Z(n832) );
  XNOR U1043 ( .A(n831), .B(n832), .Z(c[206]) );
  NAND U1044 ( .A(b[206]), .B(a[206]), .Z(n834) );
  NANDN U1045 ( .A(n832), .B(n831), .Z(n833) );
  NAND U1046 ( .A(n834), .B(n833), .Z(n836) );
  XNOR U1047 ( .A(b[207]), .B(a[207]), .Z(n835) );
  XNOR U1048 ( .A(n836), .B(n835), .Z(c[207]) );
  XNOR U1049 ( .A(b[208]), .B(a[208]), .Z(n840) );
  OR U1050 ( .A(b[207]), .B(a[207]), .Z(n838) );
  OR U1051 ( .A(n836), .B(n835), .Z(n837) );
  AND U1052 ( .A(n838), .B(n837), .Z(n839) );
  XNOR U1053 ( .A(n840), .B(n839), .Z(c[208]) );
  XNOR U1054 ( .A(b[209]), .B(a[209]), .Z(n844) );
  OR U1055 ( .A(b[208]), .B(a[208]), .Z(n842) );
  OR U1056 ( .A(n840), .B(n839), .Z(n841) );
  AND U1057 ( .A(n842), .B(n841), .Z(n843) );
  XNOR U1058 ( .A(n844), .B(n843), .Z(c[209]) );
  XNOR U1059 ( .A(b[210]), .B(a[210]), .Z(n848) );
  OR U1060 ( .A(b[209]), .B(a[209]), .Z(n846) );
  OR U1061 ( .A(n844), .B(n843), .Z(n845) );
  AND U1062 ( .A(n846), .B(n845), .Z(n847) );
  XNOR U1063 ( .A(n848), .B(n847), .Z(c[210]) );
  XNOR U1064 ( .A(b[211]), .B(a[211]), .Z(n852) );
  OR U1065 ( .A(b[210]), .B(a[210]), .Z(n850) );
  OR U1066 ( .A(n848), .B(n847), .Z(n849) );
  AND U1067 ( .A(n850), .B(n849), .Z(n851) );
  XNOR U1068 ( .A(n852), .B(n851), .Z(c[211]) );
  XNOR U1069 ( .A(b[212]), .B(a[212]), .Z(n856) );
  OR U1070 ( .A(b[211]), .B(a[211]), .Z(n854) );
  OR U1071 ( .A(n852), .B(n851), .Z(n853) );
  AND U1072 ( .A(n854), .B(n853), .Z(n855) );
  XNOR U1073 ( .A(n856), .B(n855), .Z(c[212]) );
  OR U1074 ( .A(b[212]), .B(a[212]), .Z(n858) );
  OR U1075 ( .A(n856), .B(n855), .Z(n857) );
  NAND U1076 ( .A(n858), .B(n857), .Z(n860) );
  XOR U1077 ( .A(a[213]), .B(b[213]), .Z(n859) );
  XNOR U1078 ( .A(n860), .B(n859), .Z(c[213]) );
  XOR U1079 ( .A(a[214]), .B(b[214]), .Z(n863) );
  NAND U1080 ( .A(b[213]), .B(a[213]), .Z(n862) );
  NANDN U1081 ( .A(n860), .B(n859), .Z(n861) );
  AND U1082 ( .A(n862), .B(n861), .Z(n864) );
  XNOR U1083 ( .A(n863), .B(n864), .Z(c[214]) );
  XOR U1084 ( .A(a[215]), .B(b[215]), .Z(n867) );
  NAND U1085 ( .A(b[214]), .B(a[214]), .Z(n866) );
  NANDN U1086 ( .A(n864), .B(n863), .Z(n865) );
  AND U1087 ( .A(n866), .B(n865), .Z(n868) );
  XNOR U1088 ( .A(n867), .B(n868), .Z(c[215]) );
  XOR U1089 ( .A(a[216]), .B(b[216]), .Z(n871) );
  NAND U1090 ( .A(b[215]), .B(a[215]), .Z(n870) );
  NANDN U1091 ( .A(n868), .B(n867), .Z(n869) );
  AND U1092 ( .A(n870), .B(n869), .Z(n872) );
  XNOR U1093 ( .A(n871), .B(n872), .Z(c[216]) );
  XOR U1094 ( .A(a[217]), .B(b[217]), .Z(n875) );
  NAND U1095 ( .A(b[216]), .B(a[216]), .Z(n874) );
  NANDN U1096 ( .A(n872), .B(n871), .Z(n873) );
  AND U1097 ( .A(n874), .B(n873), .Z(n876) );
  XNOR U1098 ( .A(n875), .B(n876), .Z(c[217]) );
  XOR U1099 ( .A(a[218]), .B(b[218]), .Z(n879) );
  NAND U1100 ( .A(b[217]), .B(a[217]), .Z(n878) );
  NANDN U1101 ( .A(n876), .B(n875), .Z(n877) );
  AND U1102 ( .A(n878), .B(n877), .Z(n880) );
  XNOR U1103 ( .A(n879), .B(n880), .Z(c[218]) );
  XOR U1104 ( .A(a[219]), .B(b[219]), .Z(n883) );
  NAND U1105 ( .A(b[218]), .B(a[218]), .Z(n882) );
  NANDN U1106 ( .A(n880), .B(n879), .Z(n881) );
  AND U1107 ( .A(n882), .B(n881), .Z(n884) );
  XNOR U1108 ( .A(n883), .B(n884), .Z(c[219]) );
  XOR U1109 ( .A(a[220]), .B(b[220]), .Z(n887) );
  NAND U1110 ( .A(b[219]), .B(a[219]), .Z(n886) );
  NANDN U1111 ( .A(n884), .B(n883), .Z(n885) );
  AND U1112 ( .A(n886), .B(n885), .Z(n888) );
  XNOR U1113 ( .A(n887), .B(n888), .Z(c[220]) );
  XOR U1114 ( .A(a[221]), .B(b[221]), .Z(n891) );
  NAND U1115 ( .A(b[220]), .B(a[220]), .Z(n890) );
  NANDN U1116 ( .A(n888), .B(n887), .Z(n889) );
  AND U1117 ( .A(n890), .B(n889), .Z(n892) );
  XNOR U1118 ( .A(n891), .B(n892), .Z(c[221]) );
  XOR U1119 ( .A(a[222]), .B(b[222]), .Z(n895) );
  NAND U1120 ( .A(b[221]), .B(a[221]), .Z(n894) );
  NANDN U1121 ( .A(n892), .B(n891), .Z(n893) );
  AND U1122 ( .A(n894), .B(n893), .Z(n896) );
  XNOR U1123 ( .A(n895), .B(n896), .Z(c[222]) );
  XOR U1124 ( .A(a[223]), .B(b[223]), .Z(n899) );
  NAND U1125 ( .A(b[222]), .B(a[222]), .Z(n898) );
  NANDN U1126 ( .A(n896), .B(n895), .Z(n897) );
  AND U1127 ( .A(n898), .B(n897), .Z(n900) );
  XNOR U1128 ( .A(n899), .B(n900), .Z(c[223]) );
  XOR U1129 ( .A(a[224]), .B(b[224]), .Z(n903) );
  NAND U1130 ( .A(b[223]), .B(a[223]), .Z(n902) );
  NANDN U1131 ( .A(n900), .B(n899), .Z(n901) );
  AND U1132 ( .A(n902), .B(n901), .Z(n904) );
  XNOR U1133 ( .A(n903), .B(n904), .Z(c[224]) );
  XOR U1134 ( .A(a[225]), .B(b[225]), .Z(n907) );
  NAND U1135 ( .A(b[224]), .B(a[224]), .Z(n906) );
  NANDN U1136 ( .A(n904), .B(n903), .Z(n905) );
  AND U1137 ( .A(n906), .B(n905), .Z(n908) );
  XNOR U1138 ( .A(n907), .B(n908), .Z(c[225]) );
  XOR U1139 ( .A(a[226]), .B(b[226]), .Z(n911) );
  NAND U1140 ( .A(b[225]), .B(a[225]), .Z(n910) );
  NANDN U1141 ( .A(n908), .B(n907), .Z(n909) );
  AND U1142 ( .A(n910), .B(n909), .Z(n912) );
  XNOR U1143 ( .A(n911), .B(n912), .Z(c[226]) );
  XOR U1144 ( .A(a[227]), .B(b[227]), .Z(n915) );
  NAND U1145 ( .A(b[226]), .B(a[226]), .Z(n914) );
  NANDN U1146 ( .A(n912), .B(n911), .Z(n913) );
  AND U1147 ( .A(n914), .B(n913), .Z(n916) );
  XNOR U1148 ( .A(n915), .B(n916), .Z(c[227]) );
  XOR U1149 ( .A(a[228]), .B(b[228]), .Z(n919) );
  NAND U1150 ( .A(b[227]), .B(a[227]), .Z(n918) );
  NANDN U1151 ( .A(n916), .B(n915), .Z(n917) );
  AND U1152 ( .A(n918), .B(n917), .Z(n920) );
  XNOR U1153 ( .A(n919), .B(n920), .Z(c[228]) );
  XOR U1154 ( .A(a[229]), .B(b[229]), .Z(n923) );
  NAND U1155 ( .A(b[228]), .B(a[228]), .Z(n922) );
  NANDN U1156 ( .A(n920), .B(n919), .Z(n921) );
  AND U1157 ( .A(n922), .B(n921), .Z(n924) );
  XNOR U1158 ( .A(n923), .B(n924), .Z(c[229]) );
  XOR U1159 ( .A(a[230]), .B(b[230]), .Z(n927) );
  NAND U1160 ( .A(b[229]), .B(a[229]), .Z(n926) );
  NANDN U1161 ( .A(n924), .B(n923), .Z(n925) );
  AND U1162 ( .A(n926), .B(n925), .Z(n928) );
  XNOR U1163 ( .A(n927), .B(n928), .Z(c[230]) );
  XOR U1164 ( .A(a[231]), .B(b[231]), .Z(n931) );
  NAND U1165 ( .A(b[230]), .B(a[230]), .Z(n930) );
  NANDN U1166 ( .A(n928), .B(n927), .Z(n929) );
  AND U1167 ( .A(n930), .B(n929), .Z(n932) );
  XNOR U1168 ( .A(n931), .B(n932), .Z(c[231]) );
  NAND U1169 ( .A(b[231]), .B(a[231]), .Z(n934) );
  NANDN U1170 ( .A(n932), .B(n931), .Z(n933) );
  NAND U1171 ( .A(n934), .B(n933), .Z(n936) );
  XNOR U1172 ( .A(b[232]), .B(a[232]), .Z(n935) );
  XNOR U1173 ( .A(n936), .B(n935), .Z(c[232]) );
  XNOR U1174 ( .A(b[233]), .B(a[233]), .Z(n940) );
  OR U1175 ( .A(b[232]), .B(a[232]), .Z(n938) );
  OR U1176 ( .A(n936), .B(n935), .Z(n937) );
  AND U1177 ( .A(n938), .B(n937), .Z(n939) );
  XNOR U1178 ( .A(n940), .B(n939), .Z(c[233]) );
  XOR U1179 ( .A(a[234]), .B(b[234]), .Z(n943) );
  OR U1180 ( .A(b[233]), .B(a[233]), .Z(n942) );
  OR U1181 ( .A(n940), .B(n939), .Z(n941) );
  NAND U1182 ( .A(n942), .B(n941), .Z(n944) );
  XNOR U1183 ( .A(n943), .B(n944), .Z(c[234]) );
  NAND U1184 ( .A(b[234]), .B(a[234]), .Z(n946) );
  NANDN U1185 ( .A(n944), .B(n943), .Z(n945) );
  NAND U1186 ( .A(n946), .B(n945), .Z(n948) );
  XNOR U1187 ( .A(b[235]), .B(a[235]), .Z(n947) );
  XNOR U1188 ( .A(n948), .B(n947), .Z(c[235]) );
  XNOR U1189 ( .A(b[236]), .B(a[236]), .Z(n952) );
  OR U1190 ( .A(b[235]), .B(a[235]), .Z(n950) );
  OR U1191 ( .A(n948), .B(n947), .Z(n949) );
  AND U1192 ( .A(n950), .B(n949), .Z(n951) );
  XNOR U1193 ( .A(n952), .B(n951), .Z(c[236]) );
  OR U1194 ( .A(b[236]), .B(a[236]), .Z(n954) );
  OR U1195 ( .A(n952), .B(n951), .Z(n953) );
  NAND U1196 ( .A(n954), .B(n953), .Z(n956) );
  XOR U1197 ( .A(a[237]), .B(b[237]), .Z(n955) );
  XNOR U1198 ( .A(n956), .B(n955), .Z(c[237]) );
  XOR U1199 ( .A(a[238]), .B(b[238]), .Z(n959) );
  NAND U1200 ( .A(b[237]), .B(a[237]), .Z(n958) );
  NANDN U1201 ( .A(n956), .B(n955), .Z(n957) );
  AND U1202 ( .A(n958), .B(n957), .Z(n960) );
  XNOR U1203 ( .A(n959), .B(n960), .Z(c[238]) );
  XOR U1204 ( .A(a[239]), .B(b[239]), .Z(n963) );
  NAND U1205 ( .A(b[238]), .B(a[238]), .Z(n962) );
  NANDN U1206 ( .A(n960), .B(n959), .Z(n961) );
  AND U1207 ( .A(n962), .B(n961), .Z(n964) );
  XNOR U1208 ( .A(n963), .B(n964), .Z(c[239]) );
  XOR U1209 ( .A(a[240]), .B(b[240]), .Z(n967) );
  NAND U1210 ( .A(b[239]), .B(a[239]), .Z(n966) );
  NANDN U1211 ( .A(n964), .B(n963), .Z(n965) );
  AND U1212 ( .A(n966), .B(n965), .Z(n968) );
  XNOR U1213 ( .A(n967), .B(n968), .Z(c[240]) );
  XOR U1214 ( .A(a[241]), .B(b[241]), .Z(n971) );
  NAND U1215 ( .A(b[240]), .B(a[240]), .Z(n970) );
  NANDN U1216 ( .A(n968), .B(n967), .Z(n969) );
  AND U1217 ( .A(n970), .B(n969), .Z(n972) );
  XNOR U1218 ( .A(n971), .B(n972), .Z(c[241]) );
  XOR U1219 ( .A(a[242]), .B(b[242]), .Z(n975) );
  NAND U1220 ( .A(b[241]), .B(a[241]), .Z(n974) );
  NANDN U1221 ( .A(n972), .B(n971), .Z(n973) );
  AND U1222 ( .A(n974), .B(n973), .Z(n976) );
  XNOR U1223 ( .A(n975), .B(n976), .Z(c[242]) );
  NAND U1224 ( .A(b[242]), .B(a[242]), .Z(n978) );
  NANDN U1225 ( .A(n976), .B(n975), .Z(n977) );
  NAND U1226 ( .A(n978), .B(n977), .Z(n980) );
  XNOR U1227 ( .A(b[243]), .B(a[243]), .Z(n979) );
  XNOR U1228 ( .A(n980), .B(n979), .Z(c[243]) );
  XOR U1229 ( .A(a[244]), .B(b[244]), .Z(n983) );
  OR U1230 ( .A(b[243]), .B(a[243]), .Z(n982) );
  OR U1231 ( .A(n980), .B(n979), .Z(n981) );
  NAND U1232 ( .A(n982), .B(n981), .Z(n984) );
  XNOR U1233 ( .A(n983), .B(n984), .Z(c[244]) );
  NAND U1234 ( .A(b[244]), .B(a[244]), .Z(n986) );
  NANDN U1235 ( .A(n984), .B(n983), .Z(n985) );
  NAND U1236 ( .A(n986), .B(n985), .Z(n988) );
  XNOR U1237 ( .A(b[245]), .B(a[245]), .Z(n987) );
  XNOR U1238 ( .A(n988), .B(n987), .Z(c[245]) );
  XNOR U1239 ( .A(b[246]), .B(a[246]), .Z(n992) );
  OR U1240 ( .A(b[245]), .B(a[245]), .Z(n990) );
  OR U1241 ( .A(n988), .B(n987), .Z(n989) );
  AND U1242 ( .A(n990), .B(n989), .Z(n991) );
  XNOR U1243 ( .A(n992), .B(n991), .Z(c[246]) );
  XNOR U1244 ( .A(b[247]), .B(a[247]), .Z(n996) );
  OR U1245 ( .A(b[246]), .B(a[246]), .Z(n994) );
  OR U1246 ( .A(n992), .B(n991), .Z(n993) );
  AND U1247 ( .A(n994), .B(n993), .Z(n995) );
  XNOR U1248 ( .A(n996), .B(n995), .Z(c[247]) );
  XNOR U1249 ( .A(b[248]), .B(a[248]), .Z(n1000) );
  OR U1250 ( .A(b[247]), .B(a[247]), .Z(n998) );
  OR U1251 ( .A(n996), .B(n995), .Z(n997) );
  AND U1252 ( .A(n998), .B(n997), .Z(n999) );
  XNOR U1253 ( .A(n1000), .B(n999), .Z(c[248]) );
  XNOR U1254 ( .A(b[249]), .B(a[249]), .Z(n1004) );
  OR U1255 ( .A(b[248]), .B(a[248]), .Z(n1002) );
  OR U1256 ( .A(n1000), .B(n999), .Z(n1001) );
  AND U1257 ( .A(n1002), .B(n1001), .Z(n1003) );
  XNOR U1258 ( .A(n1004), .B(n1003), .Z(c[249]) );
  XNOR U1259 ( .A(b[250]), .B(a[250]), .Z(n1008) );
  OR U1260 ( .A(b[249]), .B(a[249]), .Z(n1006) );
  OR U1261 ( .A(n1004), .B(n1003), .Z(n1005) );
  AND U1262 ( .A(n1006), .B(n1005), .Z(n1007) );
  XNOR U1263 ( .A(n1008), .B(n1007), .Z(c[250]) );
  XNOR U1264 ( .A(b[251]), .B(a[251]), .Z(n1012) );
  OR U1265 ( .A(b[250]), .B(a[250]), .Z(n1010) );
  OR U1266 ( .A(n1008), .B(n1007), .Z(n1009) );
  AND U1267 ( .A(n1010), .B(n1009), .Z(n1011) );
  XNOR U1268 ( .A(n1012), .B(n1011), .Z(c[251]) );
  XNOR U1269 ( .A(b[252]), .B(a[252]), .Z(n1016) );
  OR U1270 ( .A(b[251]), .B(a[251]), .Z(n1014) );
  OR U1271 ( .A(n1012), .B(n1011), .Z(n1013) );
  AND U1272 ( .A(n1014), .B(n1013), .Z(n1015) );
  XNOR U1273 ( .A(n1016), .B(n1015), .Z(c[252]) );
  XNOR U1274 ( .A(b[253]), .B(a[253]), .Z(n1020) );
  OR U1275 ( .A(b[252]), .B(a[252]), .Z(n1018) );
  OR U1276 ( .A(n1016), .B(n1015), .Z(n1017) );
  AND U1277 ( .A(n1018), .B(n1017), .Z(n1019) );
  XNOR U1278 ( .A(n1020), .B(n1019), .Z(c[253]) );
  XNOR U1279 ( .A(b[254]), .B(a[254]), .Z(n1024) );
  OR U1280 ( .A(b[253]), .B(a[253]), .Z(n1022) );
  OR U1281 ( .A(n1020), .B(n1019), .Z(n1021) );
  AND U1282 ( .A(n1022), .B(n1021), .Z(n1023) );
  XNOR U1283 ( .A(n1024), .B(n1023), .Z(c[254]) );
  XNOR U1284 ( .A(b[255]), .B(a[255]), .Z(n1028) );
  OR U1285 ( .A(b[254]), .B(a[254]), .Z(n1026) );
  OR U1286 ( .A(n1024), .B(n1023), .Z(n1025) );
  AND U1287 ( .A(n1026), .B(n1025), .Z(n1027) );
  XNOR U1288 ( .A(n1028), .B(n1027), .Z(c[255]) );
  XNOR U1289 ( .A(b[256]), .B(a[256]), .Z(n1032) );
  OR U1290 ( .A(b[255]), .B(a[255]), .Z(n1030) );
  OR U1291 ( .A(n1028), .B(n1027), .Z(n1029) );
  AND U1292 ( .A(n1030), .B(n1029), .Z(n1031) );
  XNOR U1293 ( .A(n1032), .B(n1031), .Z(c[256]) );
  XNOR U1294 ( .A(b[257]), .B(a[257]), .Z(n1036) );
  OR U1295 ( .A(b[256]), .B(a[256]), .Z(n1034) );
  OR U1296 ( .A(n1032), .B(n1031), .Z(n1033) );
  AND U1297 ( .A(n1034), .B(n1033), .Z(n1035) );
  XNOR U1298 ( .A(n1036), .B(n1035), .Z(c[257]) );
  XNOR U1299 ( .A(b[258]), .B(a[258]), .Z(n1040) );
  OR U1300 ( .A(b[257]), .B(a[257]), .Z(n1038) );
  OR U1301 ( .A(n1036), .B(n1035), .Z(n1037) );
  AND U1302 ( .A(n1038), .B(n1037), .Z(n1039) );
  XNOR U1303 ( .A(n1040), .B(n1039), .Z(c[258]) );
  XNOR U1304 ( .A(b[259]), .B(a[259]), .Z(n1044) );
  OR U1305 ( .A(b[258]), .B(a[258]), .Z(n1042) );
  OR U1306 ( .A(n1040), .B(n1039), .Z(n1041) );
  AND U1307 ( .A(n1042), .B(n1041), .Z(n1043) );
  XNOR U1308 ( .A(n1044), .B(n1043), .Z(c[259]) );
  XNOR U1309 ( .A(b[260]), .B(a[260]), .Z(n1048) );
  OR U1310 ( .A(b[259]), .B(a[259]), .Z(n1046) );
  OR U1311 ( .A(n1044), .B(n1043), .Z(n1045) );
  AND U1312 ( .A(n1046), .B(n1045), .Z(n1047) );
  XNOR U1313 ( .A(n1048), .B(n1047), .Z(c[260]) );
  XNOR U1314 ( .A(b[261]), .B(a[261]), .Z(n1052) );
  OR U1315 ( .A(b[260]), .B(a[260]), .Z(n1050) );
  OR U1316 ( .A(n1048), .B(n1047), .Z(n1049) );
  AND U1317 ( .A(n1050), .B(n1049), .Z(n1051) );
  XNOR U1318 ( .A(n1052), .B(n1051), .Z(c[261]) );
  OR U1319 ( .A(b[261]), .B(a[261]), .Z(n1054) );
  OR U1320 ( .A(n1052), .B(n1051), .Z(n1053) );
  NAND U1321 ( .A(n1054), .B(n1053), .Z(n1056) );
  XOR U1322 ( .A(a[262]), .B(b[262]), .Z(n1055) );
  XNOR U1323 ( .A(n1056), .B(n1055), .Z(c[262]) );
  NAND U1324 ( .A(b[262]), .B(a[262]), .Z(n1058) );
  NANDN U1325 ( .A(n1056), .B(n1055), .Z(n1057) );
  NAND U1326 ( .A(n1058), .B(n1057), .Z(n1060) );
  XNOR U1327 ( .A(b[263]), .B(a[263]), .Z(n1059) );
  XNOR U1328 ( .A(n1060), .B(n1059), .Z(c[263]) );
  XNOR U1329 ( .A(b[264]), .B(a[264]), .Z(n1064) );
  OR U1330 ( .A(b[263]), .B(a[263]), .Z(n1062) );
  OR U1331 ( .A(n1060), .B(n1059), .Z(n1061) );
  AND U1332 ( .A(n1062), .B(n1061), .Z(n1063) );
  XNOR U1333 ( .A(n1064), .B(n1063), .Z(c[264]) );
  XOR U1334 ( .A(a[265]), .B(b[265]), .Z(n1067) );
  OR U1335 ( .A(b[264]), .B(a[264]), .Z(n1066) );
  OR U1336 ( .A(n1064), .B(n1063), .Z(n1065) );
  NAND U1337 ( .A(n1066), .B(n1065), .Z(n1068) );
  XNOR U1338 ( .A(n1067), .B(n1068), .Z(c[265]) );
  NAND U1339 ( .A(b[265]), .B(a[265]), .Z(n1070) );
  NANDN U1340 ( .A(n1068), .B(n1067), .Z(n1069) );
  NAND U1341 ( .A(n1070), .B(n1069), .Z(n1072) );
  XNOR U1342 ( .A(b[266]), .B(a[266]), .Z(n1071) );
  XNOR U1343 ( .A(n1072), .B(n1071), .Z(c[266]) );
  XNOR U1344 ( .A(b[267]), .B(a[267]), .Z(n1076) );
  OR U1345 ( .A(b[266]), .B(a[266]), .Z(n1074) );
  OR U1346 ( .A(n1072), .B(n1071), .Z(n1073) );
  AND U1347 ( .A(n1074), .B(n1073), .Z(n1075) );
  XNOR U1348 ( .A(n1076), .B(n1075), .Z(c[267]) );
  XNOR U1349 ( .A(b[268]), .B(a[268]), .Z(n1080) );
  OR U1350 ( .A(b[267]), .B(a[267]), .Z(n1078) );
  OR U1351 ( .A(n1076), .B(n1075), .Z(n1077) );
  AND U1352 ( .A(n1078), .B(n1077), .Z(n1079) );
  XNOR U1353 ( .A(n1080), .B(n1079), .Z(c[268]) );
  XNOR U1354 ( .A(b[269]), .B(a[269]), .Z(n1084) );
  OR U1355 ( .A(b[268]), .B(a[268]), .Z(n1082) );
  OR U1356 ( .A(n1080), .B(n1079), .Z(n1081) );
  AND U1357 ( .A(n1082), .B(n1081), .Z(n1083) );
  XNOR U1358 ( .A(n1084), .B(n1083), .Z(c[269]) );
  XNOR U1359 ( .A(b[270]), .B(a[270]), .Z(n1088) );
  OR U1360 ( .A(b[269]), .B(a[269]), .Z(n1086) );
  OR U1361 ( .A(n1084), .B(n1083), .Z(n1085) );
  AND U1362 ( .A(n1086), .B(n1085), .Z(n1087) );
  XNOR U1363 ( .A(n1088), .B(n1087), .Z(c[270]) );
  XNOR U1364 ( .A(b[271]), .B(a[271]), .Z(n1092) );
  OR U1365 ( .A(b[270]), .B(a[270]), .Z(n1090) );
  OR U1366 ( .A(n1088), .B(n1087), .Z(n1089) );
  AND U1367 ( .A(n1090), .B(n1089), .Z(n1091) );
  XNOR U1368 ( .A(n1092), .B(n1091), .Z(c[271]) );
  XNOR U1369 ( .A(b[272]), .B(a[272]), .Z(n1096) );
  OR U1370 ( .A(b[271]), .B(a[271]), .Z(n1094) );
  OR U1371 ( .A(n1092), .B(n1091), .Z(n1093) );
  AND U1372 ( .A(n1094), .B(n1093), .Z(n1095) );
  XNOR U1373 ( .A(n1096), .B(n1095), .Z(c[272]) );
  XNOR U1374 ( .A(b[273]), .B(a[273]), .Z(n1100) );
  OR U1375 ( .A(b[272]), .B(a[272]), .Z(n1098) );
  OR U1376 ( .A(n1096), .B(n1095), .Z(n1097) );
  AND U1377 ( .A(n1098), .B(n1097), .Z(n1099) );
  XNOR U1378 ( .A(n1100), .B(n1099), .Z(c[273]) );
  XNOR U1379 ( .A(b[274]), .B(a[274]), .Z(n1104) );
  OR U1380 ( .A(b[273]), .B(a[273]), .Z(n1102) );
  OR U1381 ( .A(n1100), .B(n1099), .Z(n1101) );
  AND U1382 ( .A(n1102), .B(n1101), .Z(n1103) );
  XNOR U1383 ( .A(n1104), .B(n1103), .Z(c[274]) );
  XNOR U1384 ( .A(b[275]), .B(a[275]), .Z(n1108) );
  OR U1385 ( .A(b[274]), .B(a[274]), .Z(n1106) );
  OR U1386 ( .A(n1104), .B(n1103), .Z(n1105) );
  AND U1387 ( .A(n1106), .B(n1105), .Z(n1107) );
  XNOR U1388 ( .A(n1108), .B(n1107), .Z(c[275]) );
  XNOR U1389 ( .A(b[276]), .B(a[276]), .Z(n1112) );
  OR U1390 ( .A(b[275]), .B(a[275]), .Z(n1110) );
  OR U1391 ( .A(n1108), .B(n1107), .Z(n1109) );
  AND U1392 ( .A(n1110), .B(n1109), .Z(n1111) );
  XNOR U1393 ( .A(n1112), .B(n1111), .Z(c[276]) );
  XNOR U1394 ( .A(b[277]), .B(a[277]), .Z(n1116) );
  OR U1395 ( .A(b[276]), .B(a[276]), .Z(n1114) );
  OR U1396 ( .A(n1112), .B(n1111), .Z(n1113) );
  AND U1397 ( .A(n1114), .B(n1113), .Z(n1115) );
  XNOR U1398 ( .A(n1116), .B(n1115), .Z(c[277]) );
  XNOR U1399 ( .A(b[278]), .B(a[278]), .Z(n1120) );
  OR U1400 ( .A(b[277]), .B(a[277]), .Z(n1118) );
  OR U1401 ( .A(n1116), .B(n1115), .Z(n1117) );
  AND U1402 ( .A(n1118), .B(n1117), .Z(n1119) );
  XNOR U1403 ( .A(n1120), .B(n1119), .Z(c[278]) );
  XNOR U1404 ( .A(b[279]), .B(a[279]), .Z(n1124) );
  OR U1405 ( .A(b[278]), .B(a[278]), .Z(n1122) );
  OR U1406 ( .A(n1120), .B(n1119), .Z(n1121) );
  AND U1407 ( .A(n1122), .B(n1121), .Z(n1123) );
  XNOR U1408 ( .A(n1124), .B(n1123), .Z(c[279]) );
  XNOR U1409 ( .A(b[280]), .B(a[280]), .Z(n1128) );
  OR U1410 ( .A(b[279]), .B(a[279]), .Z(n1126) );
  OR U1411 ( .A(n1124), .B(n1123), .Z(n1125) );
  AND U1412 ( .A(n1126), .B(n1125), .Z(n1127) );
  XNOR U1413 ( .A(n1128), .B(n1127), .Z(c[280]) );
  XNOR U1414 ( .A(b[281]), .B(a[281]), .Z(n1132) );
  OR U1415 ( .A(b[280]), .B(a[280]), .Z(n1130) );
  OR U1416 ( .A(n1128), .B(n1127), .Z(n1129) );
  AND U1417 ( .A(n1130), .B(n1129), .Z(n1131) );
  XNOR U1418 ( .A(n1132), .B(n1131), .Z(c[281]) );
  XNOR U1419 ( .A(b[282]), .B(a[282]), .Z(n1136) );
  OR U1420 ( .A(b[281]), .B(a[281]), .Z(n1134) );
  OR U1421 ( .A(n1132), .B(n1131), .Z(n1133) );
  AND U1422 ( .A(n1134), .B(n1133), .Z(n1135) );
  XNOR U1423 ( .A(n1136), .B(n1135), .Z(c[282]) );
  XNOR U1424 ( .A(b[283]), .B(a[283]), .Z(n1140) );
  OR U1425 ( .A(b[282]), .B(a[282]), .Z(n1138) );
  OR U1426 ( .A(n1136), .B(n1135), .Z(n1137) );
  AND U1427 ( .A(n1138), .B(n1137), .Z(n1139) );
  XNOR U1428 ( .A(n1140), .B(n1139), .Z(c[283]) );
  XNOR U1429 ( .A(b[284]), .B(a[284]), .Z(n1144) );
  OR U1430 ( .A(b[283]), .B(a[283]), .Z(n1142) );
  OR U1431 ( .A(n1140), .B(n1139), .Z(n1141) );
  AND U1432 ( .A(n1142), .B(n1141), .Z(n1143) );
  XNOR U1433 ( .A(n1144), .B(n1143), .Z(c[284]) );
  XNOR U1434 ( .A(b[285]), .B(a[285]), .Z(n1148) );
  OR U1435 ( .A(b[284]), .B(a[284]), .Z(n1146) );
  OR U1436 ( .A(n1144), .B(n1143), .Z(n1145) );
  AND U1437 ( .A(n1146), .B(n1145), .Z(n1147) );
  XNOR U1438 ( .A(n1148), .B(n1147), .Z(c[285]) );
  OR U1439 ( .A(b[285]), .B(a[285]), .Z(n1150) );
  OR U1440 ( .A(n1148), .B(n1147), .Z(n1149) );
  NAND U1441 ( .A(n1150), .B(n1149), .Z(n1152) );
  XOR U1442 ( .A(a[286]), .B(b[286]), .Z(n1151) );
  XNOR U1443 ( .A(n1152), .B(n1151), .Z(c[286]) );
  XOR U1444 ( .A(a[287]), .B(b[287]), .Z(n1155) );
  NAND U1445 ( .A(b[286]), .B(a[286]), .Z(n1154) );
  NANDN U1446 ( .A(n1152), .B(n1151), .Z(n1153) );
  AND U1447 ( .A(n1154), .B(n1153), .Z(n1156) );
  XNOR U1448 ( .A(n1155), .B(n1156), .Z(c[287]) );
  XNOR U1449 ( .A(b[288]), .B(a[288]), .Z(n1160) );
  NAND U1450 ( .A(b[287]), .B(a[287]), .Z(n1158) );
  NANDN U1451 ( .A(n1156), .B(n1155), .Z(n1157) );
  NAND U1452 ( .A(n1158), .B(n1157), .Z(n1159) );
  XNOR U1453 ( .A(n1160), .B(n1159), .Z(c[288]) );
  OR U1454 ( .A(b[288]), .B(a[288]), .Z(n1162) );
  OR U1455 ( .A(n1160), .B(n1159), .Z(n1161) );
  NAND U1456 ( .A(n1162), .B(n1161), .Z(n1164) );
  XOR U1457 ( .A(a[289]), .B(b[289]), .Z(n1163) );
  XNOR U1458 ( .A(n1164), .B(n1163), .Z(c[289]) );
  XOR U1459 ( .A(a[290]), .B(b[290]), .Z(n1167) );
  NAND U1460 ( .A(b[289]), .B(a[289]), .Z(n1166) );
  NANDN U1461 ( .A(n1164), .B(n1163), .Z(n1165) );
  AND U1462 ( .A(n1166), .B(n1165), .Z(n1168) );
  XNOR U1463 ( .A(n1167), .B(n1168), .Z(c[290]) );
  XOR U1464 ( .A(a[291]), .B(b[291]), .Z(n1171) );
  NAND U1465 ( .A(b[290]), .B(a[290]), .Z(n1170) );
  NANDN U1466 ( .A(n1168), .B(n1167), .Z(n1169) );
  AND U1467 ( .A(n1170), .B(n1169), .Z(n1172) );
  XNOR U1468 ( .A(n1171), .B(n1172), .Z(c[291]) );
  XOR U1469 ( .A(a[292]), .B(b[292]), .Z(n1175) );
  NAND U1470 ( .A(b[291]), .B(a[291]), .Z(n1174) );
  NANDN U1471 ( .A(n1172), .B(n1171), .Z(n1173) );
  AND U1472 ( .A(n1174), .B(n1173), .Z(n1176) );
  XNOR U1473 ( .A(n1175), .B(n1176), .Z(c[292]) );
  XOR U1474 ( .A(a[293]), .B(b[293]), .Z(n1179) );
  NAND U1475 ( .A(b[292]), .B(a[292]), .Z(n1178) );
  NANDN U1476 ( .A(n1176), .B(n1175), .Z(n1177) );
  AND U1477 ( .A(n1178), .B(n1177), .Z(n1180) );
  XNOR U1478 ( .A(n1179), .B(n1180), .Z(c[293]) );
  XOR U1479 ( .A(a[294]), .B(b[294]), .Z(n1183) );
  NAND U1480 ( .A(b[293]), .B(a[293]), .Z(n1182) );
  NANDN U1481 ( .A(n1180), .B(n1179), .Z(n1181) );
  AND U1482 ( .A(n1182), .B(n1181), .Z(n1184) );
  XNOR U1483 ( .A(n1183), .B(n1184), .Z(c[294]) );
  XOR U1484 ( .A(a[295]), .B(b[295]), .Z(n1187) );
  NAND U1485 ( .A(b[294]), .B(a[294]), .Z(n1186) );
  NANDN U1486 ( .A(n1184), .B(n1183), .Z(n1185) );
  AND U1487 ( .A(n1186), .B(n1185), .Z(n1188) );
  XNOR U1488 ( .A(n1187), .B(n1188), .Z(c[295]) );
  XOR U1489 ( .A(a[296]), .B(b[296]), .Z(n1191) );
  NAND U1490 ( .A(b[295]), .B(a[295]), .Z(n1190) );
  NANDN U1491 ( .A(n1188), .B(n1187), .Z(n1189) );
  AND U1492 ( .A(n1190), .B(n1189), .Z(n1192) );
  XNOR U1493 ( .A(n1191), .B(n1192), .Z(c[296]) );
  XOR U1494 ( .A(a[297]), .B(b[297]), .Z(n1195) );
  NAND U1495 ( .A(b[296]), .B(a[296]), .Z(n1194) );
  NANDN U1496 ( .A(n1192), .B(n1191), .Z(n1193) );
  AND U1497 ( .A(n1194), .B(n1193), .Z(n1196) );
  XNOR U1498 ( .A(n1195), .B(n1196), .Z(c[297]) );
  XOR U1499 ( .A(a[298]), .B(b[298]), .Z(n1199) );
  NAND U1500 ( .A(b[297]), .B(a[297]), .Z(n1198) );
  NANDN U1501 ( .A(n1196), .B(n1195), .Z(n1197) );
  AND U1502 ( .A(n1198), .B(n1197), .Z(n1200) );
  XNOR U1503 ( .A(n1199), .B(n1200), .Z(c[298]) );
  XOR U1504 ( .A(a[299]), .B(b[299]), .Z(n1203) );
  NAND U1505 ( .A(b[298]), .B(a[298]), .Z(n1202) );
  NANDN U1506 ( .A(n1200), .B(n1199), .Z(n1201) );
  AND U1507 ( .A(n1202), .B(n1201), .Z(n1204) );
  XNOR U1508 ( .A(n1203), .B(n1204), .Z(c[299]) );
  NAND U1509 ( .A(b[299]), .B(a[299]), .Z(n1206) );
  NANDN U1510 ( .A(n1204), .B(n1203), .Z(n1205) );
  NAND U1511 ( .A(n1206), .B(n1205), .Z(n1208) );
  XNOR U1512 ( .A(b[300]), .B(a[300]), .Z(n1207) );
  XNOR U1513 ( .A(n1208), .B(n1207), .Z(c[300]) );
  XNOR U1514 ( .A(b[301]), .B(a[301]), .Z(n1212) );
  OR U1515 ( .A(b[300]), .B(a[300]), .Z(n1210) );
  OR U1516 ( .A(n1208), .B(n1207), .Z(n1209) );
  AND U1517 ( .A(n1210), .B(n1209), .Z(n1211) );
  XNOR U1518 ( .A(n1212), .B(n1211), .Z(c[301]) );
  OR U1519 ( .A(b[301]), .B(a[301]), .Z(n1214) );
  OR U1520 ( .A(n1212), .B(n1211), .Z(n1213) );
  NAND U1521 ( .A(n1214), .B(n1213), .Z(n1216) );
  XOR U1522 ( .A(a[302]), .B(b[302]), .Z(n1215) );
  XNOR U1523 ( .A(n1216), .B(n1215), .Z(c[302]) );
  NAND U1524 ( .A(b[302]), .B(a[302]), .Z(n1218) );
  NANDN U1525 ( .A(n1216), .B(n1215), .Z(n1217) );
  NAND U1526 ( .A(n1218), .B(n1217), .Z(n1220) );
  XNOR U1527 ( .A(b[303]), .B(a[303]), .Z(n1219) );
  XNOR U1528 ( .A(n1220), .B(n1219), .Z(c[303]) );
  XNOR U1529 ( .A(b[304]), .B(a[304]), .Z(n1224) );
  OR U1530 ( .A(b[303]), .B(a[303]), .Z(n1222) );
  OR U1531 ( .A(n1220), .B(n1219), .Z(n1221) );
  AND U1532 ( .A(n1222), .B(n1221), .Z(n1223) );
  XNOR U1533 ( .A(n1224), .B(n1223), .Z(c[304]) );
  XNOR U1534 ( .A(b[305]), .B(a[305]), .Z(n1228) );
  OR U1535 ( .A(b[304]), .B(a[304]), .Z(n1226) );
  OR U1536 ( .A(n1224), .B(n1223), .Z(n1225) );
  AND U1537 ( .A(n1226), .B(n1225), .Z(n1227) );
  XNOR U1538 ( .A(n1228), .B(n1227), .Z(c[305]) );
  XNOR U1539 ( .A(b[306]), .B(a[306]), .Z(n1232) );
  OR U1540 ( .A(b[305]), .B(a[305]), .Z(n1230) );
  OR U1541 ( .A(n1228), .B(n1227), .Z(n1229) );
  AND U1542 ( .A(n1230), .B(n1229), .Z(n1231) );
  XNOR U1543 ( .A(n1232), .B(n1231), .Z(c[306]) );
  XNOR U1544 ( .A(b[307]), .B(a[307]), .Z(n1236) );
  OR U1545 ( .A(b[306]), .B(a[306]), .Z(n1234) );
  OR U1546 ( .A(n1232), .B(n1231), .Z(n1233) );
  AND U1547 ( .A(n1234), .B(n1233), .Z(n1235) );
  XNOR U1548 ( .A(n1236), .B(n1235), .Z(c[307]) );
  XNOR U1549 ( .A(b[308]), .B(a[308]), .Z(n1240) );
  OR U1550 ( .A(b[307]), .B(a[307]), .Z(n1238) );
  OR U1551 ( .A(n1236), .B(n1235), .Z(n1237) );
  AND U1552 ( .A(n1238), .B(n1237), .Z(n1239) );
  XNOR U1553 ( .A(n1240), .B(n1239), .Z(c[308]) );
  XNOR U1554 ( .A(b[309]), .B(a[309]), .Z(n1244) );
  OR U1555 ( .A(b[308]), .B(a[308]), .Z(n1242) );
  OR U1556 ( .A(n1240), .B(n1239), .Z(n1241) );
  AND U1557 ( .A(n1242), .B(n1241), .Z(n1243) );
  XNOR U1558 ( .A(n1244), .B(n1243), .Z(c[309]) );
  XNOR U1559 ( .A(b[310]), .B(a[310]), .Z(n1248) );
  OR U1560 ( .A(b[309]), .B(a[309]), .Z(n1246) );
  OR U1561 ( .A(n1244), .B(n1243), .Z(n1245) );
  AND U1562 ( .A(n1246), .B(n1245), .Z(n1247) );
  XNOR U1563 ( .A(n1248), .B(n1247), .Z(c[310]) );
  OR U1564 ( .A(b[310]), .B(a[310]), .Z(n1250) );
  OR U1565 ( .A(n1248), .B(n1247), .Z(n1249) );
  NAND U1566 ( .A(n1250), .B(n1249), .Z(n1252) );
  XOR U1567 ( .A(a[311]), .B(b[311]), .Z(n1251) );
  XNOR U1568 ( .A(n1252), .B(n1251), .Z(c[311]) );
  XOR U1569 ( .A(a[312]), .B(b[312]), .Z(n1255) );
  NAND U1570 ( .A(b[311]), .B(a[311]), .Z(n1254) );
  NANDN U1571 ( .A(n1252), .B(n1251), .Z(n1253) );
  AND U1572 ( .A(n1254), .B(n1253), .Z(n1256) );
  XNOR U1573 ( .A(n1255), .B(n1256), .Z(c[312]) );
  XNOR U1574 ( .A(b[313]), .B(a[313]), .Z(n1260) );
  NAND U1575 ( .A(b[312]), .B(a[312]), .Z(n1258) );
  NANDN U1576 ( .A(n1256), .B(n1255), .Z(n1257) );
  NAND U1577 ( .A(n1258), .B(n1257), .Z(n1259) );
  XNOR U1578 ( .A(n1260), .B(n1259), .Z(c[313]) );
  OR U1579 ( .A(b[313]), .B(a[313]), .Z(n1262) );
  OR U1580 ( .A(n1260), .B(n1259), .Z(n1261) );
  NAND U1581 ( .A(n1262), .B(n1261), .Z(n1264) );
  XOR U1582 ( .A(a[314]), .B(b[314]), .Z(n1263) );
  XNOR U1583 ( .A(n1264), .B(n1263), .Z(c[314]) );
  XOR U1584 ( .A(a[315]), .B(b[315]), .Z(n1267) );
  NAND U1585 ( .A(b[314]), .B(a[314]), .Z(n1266) );
  NANDN U1586 ( .A(n1264), .B(n1263), .Z(n1265) );
  AND U1587 ( .A(n1266), .B(n1265), .Z(n1268) );
  XNOR U1588 ( .A(n1267), .B(n1268), .Z(c[315]) );
  NAND U1589 ( .A(b[315]), .B(a[315]), .Z(n1270) );
  NANDN U1590 ( .A(n1268), .B(n1267), .Z(n1269) );
  NAND U1591 ( .A(n1270), .B(n1269), .Z(n1272) );
  XNOR U1592 ( .A(b[316]), .B(a[316]), .Z(n1271) );
  XNOR U1593 ( .A(n1272), .B(n1271), .Z(c[316]) );
  XNOR U1594 ( .A(b[317]), .B(a[317]), .Z(n1276) );
  OR U1595 ( .A(b[316]), .B(a[316]), .Z(n1274) );
  OR U1596 ( .A(n1272), .B(n1271), .Z(n1273) );
  AND U1597 ( .A(n1274), .B(n1273), .Z(n1275) );
  XNOR U1598 ( .A(n1276), .B(n1275), .Z(c[317]) );
  XOR U1599 ( .A(a[318]), .B(b[318]), .Z(n1279) );
  OR U1600 ( .A(b[317]), .B(a[317]), .Z(n1278) );
  OR U1601 ( .A(n1276), .B(n1275), .Z(n1277) );
  NAND U1602 ( .A(n1278), .B(n1277), .Z(n1280) );
  XNOR U1603 ( .A(n1279), .B(n1280), .Z(c[318]) );
  XNOR U1604 ( .A(b[319]), .B(a[319]), .Z(n1284) );
  NAND U1605 ( .A(b[318]), .B(a[318]), .Z(n1282) );
  NANDN U1606 ( .A(n1280), .B(n1279), .Z(n1281) );
  NAND U1607 ( .A(n1282), .B(n1281), .Z(n1283) );
  XNOR U1608 ( .A(n1284), .B(n1283), .Z(c[319]) );
  XNOR U1609 ( .A(b[320]), .B(a[320]), .Z(n1288) );
  OR U1610 ( .A(b[319]), .B(a[319]), .Z(n1286) );
  OR U1611 ( .A(n1284), .B(n1283), .Z(n1285) );
  AND U1612 ( .A(n1286), .B(n1285), .Z(n1287) );
  XNOR U1613 ( .A(n1288), .B(n1287), .Z(c[320]) );
  XOR U1614 ( .A(a[321]), .B(b[321]), .Z(n1291) );
  OR U1615 ( .A(b[320]), .B(a[320]), .Z(n1290) );
  OR U1616 ( .A(n1288), .B(n1287), .Z(n1289) );
  NAND U1617 ( .A(n1290), .B(n1289), .Z(n1292) );
  XNOR U1618 ( .A(n1291), .B(n1292), .Z(c[321]) );
  XOR U1619 ( .A(a[322]), .B(b[322]), .Z(n1295) );
  NAND U1620 ( .A(b[321]), .B(a[321]), .Z(n1294) );
  NANDN U1621 ( .A(n1292), .B(n1291), .Z(n1293) );
  AND U1622 ( .A(n1294), .B(n1293), .Z(n1296) );
  XNOR U1623 ( .A(n1295), .B(n1296), .Z(c[322]) );
  XOR U1624 ( .A(a[323]), .B(b[323]), .Z(n1299) );
  NAND U1625 ( .A(b[322]), .B(a[322]), .Z(n1298) );
  NANDN U1626 ( .A(n1296), .B(n1295), .Z(n1297) );
  AND U1627 ( .A(n1298), .B(n1297), .Z(n1300) );
  XNOR U1628 ( .A(n1299), .B(n1300), .Z(c[323]) );
  XOR U1629 ( .A(a[324]), .B(b[324]), .Z(n1303) );
  NAND U1630 ( .A(b[323]), .B(a[323]), .Z(n1302) );
  NANDN U1631 ( .A(n1300), .B(n1299), .Z(n1301) );
  AND U1632 ( .A(n1302), .B(n1301), .Z(n1304) );
  XNOR U1633 ( .A(n1303), .B(n1304), .Z(c[324]) );
  XOR U1634 ( .A(a[325]), .B(b[325]), .Z(n1307) );
  NAND U1635 ( .A(b[324]), .B(a[324]), .Z(n1306) );
  NANDN U1636 ( .A(n1304), .B(n1303), .Z(n1305) );
  AND U1637 ( .A(n1306), .B(n1305), .Z(n1308) );
  XNOR U1638 ( .A(n1307), .B(n1308), .Z(c[325]) );
  XOR U1639 ( .A(a[326]), .B(b[326]), .Z(n1311) );
  NAND U1640 ( .A(b[325]), .B(a[325]), .Z(n1310) );
  NANDN U1641 ( .A(n1308), .B(n1307), .Z(n1309) );
  AND U1642 ( .A(n1310), .B(n1309), .Z(n1312) );
  XNOR U1643 ( .A(n1311), .B(n1312), .Z(c[326]) );
  XOR U1644 ( .A(a[327]), .B(b[327]), .Z(n1315) );
  NAND U1645 ( .A(b[326]), .B(a[326]), .Z(n1314) );
  NANDN U1646 ( .A(n1312), .B(n1311), .Z(n1313) );
  AND U1647 ( .A(n1314), .B(n1313), .Z(n1316) );
  XNOR U1648 ( .A(n1315), .B(n1316), .Z(c[327]) );
  XOR U1649 ( .A(a[328]), .B(b[328]), .Z(n1319) );
  NAND U1650 ( .A(b[327]), .B(a[327]), .Z(n1318) );
  NANDN U1651 ( .A(n1316), .B(n1315), .Z(n1317) );
  AND U1652 ( .A(n1318), .B(n1317), .Z(n1320) );
  XNOR U1653 ( .A(n1319), .B(n1320), .Z(c[328]) );
  XOR U1654 ( .A(a[329]), .B(b[329]), .Z(n1323) );
  NAND U1655 ( .A(b[328]), .B(a[328]), .Z(n1322) );
  NANDN U1656 ( .A(n1320), .B(n1319), .Z(n1321) );
  AND U1657 ( .A(n1322), .B(n1321), .Z(n1324) );
  XNOR U1658 ( .A(n1323), .B(n1324), .Z(c[329]) );
  XOR U1659 ( .A(a[330]), .B(b[330]), .Z(n1327) );
  NAND U1660 ( .A(b[329]), .B(a[329]), .Z(n1326) );
  NANDN U1661 ( .A(n1324), .B(n1323), .Z(n1325) );
  AND U1662 ( .A(n1326), .B(n1325), .Z(n1328) );
  XNOR U1663 ( .A(n1327), .B(n1328), .Z(c[330]) );
  XOR U1664 ( .A(a[331]), .B(b[331]), .Z(n1331) );
  NAND U1665 ( .A(b[330]), .B(a[330]), .Z(n1330) );
  NANDN U1666 ( .A(n1328), .B(n1327), .Z(n1329) );
  AND U1667 ( .A(n1330), .B(n1329), .Z(n1332) );
  XNOR U1668 ( .A(n1331), .B(n1332), .Z(c[331]) );
  XOR U1669 ( .A(a[332]), .B(b[332]), .Z(n1335) );
  NAND U1670 ( .A(b[331]), .B(a[331]), .Z(n1334) );
  NANDN U1671 ( .A(n1332), .B(n1331), .Z(n1333) );
  AND U1672 ( .A(n1334), .B(n1333), .Z(n1336) );
  XNOR U1673 ( .A(n1335), .B(n1336), .Z(c[332]) );
  NAND U1674 ( .A(b[332]), .B(a[332]), .Z(n1338) );
  NANDN U1675 ( .A(n1336), .B(n1335), .Z(n1337) );
  NAND U1676 ( .A(n1338), .B(n1337), .Z(n1340) );
  XNOR U1677 ( .A(b[333]), .B(a[333]), .Z(n1339) );
  XNOR U1678 ( .A(n1340), .B(n1339), .Z(c[333]) );
  XOR U1679 ( .A(a[334]), .B(b[334]), .Z(n1343) );
  OR U1680 ( .A(b[333]), .B(a[333]), .Z(n1342) );
  OR U1681 ( .A(n1340), .B(n1339), .Z(n1341) );
  NAND U1682 ( .A(n1342), .B(n1341), .Z(n1344) );
  XNOR U1683 ( .A(n1343), .B(n1344), .Z(c[334]) );
  NAND U1684 ( .A(b[334]), .B(a[334]), .Z(n1346) );
  NANDN U1685 ( .A(n1344), .B(n1343), .Z(n1345) );
  NAND U1686 ( .A(n1346), .B(n1345), .Z(n1348) );
  XNOR U1687 ( .A(b[335]), .B(a[335]), .Z(n1347) );
  XNOR U1688 ( .A(n1348), .B(n1347), .Z(c[335]) );
  XNOR U1689 ( .A(b[336]), .B(a[336]), .Z(n1352) );
  OR U1690 ( .A(b[335]), .B(a[335]), .Z(n1350) );
  OR U1691 ( .A(n1348), .B(n1347), .Z(n1349) );
  AND U1692 ( .A(n1350), .B(n1349), .Z(n1351) );
  XNOR U1693 ( .A(n1352), .B(n1351), .Z(c[336]) );
  XNOR U1694 ( .A(b[337]), .B(a[337]), .Z(n1356) );
  OR U1695 ( .A(b[336]), .B(a[336]), .Z(n1354) );
  OR U1696 ( .A(n1352), .B(n1351), .Z(n1353) );
  AND U1697 ( .A(n1354), .B(n1353), .Z(n1355) );
  XNOR U1698 ( .A(n1356), .B(n1355), .Z(c[337]) );
  XNOR U1699 ( .A(b[338]), .B(a[338]), .Z(n1360) );
  OR U1700 ( .A(b[337]), .B(a[337]), .Z(n1358) );
  OR U1701 ( .A(n1356), .B(n1355), .Z(n1357) );
  AND U1702 ( .A(n1358), .B(n1357), .Z(n1359) );
  XNOR U1703 ( .A(n1360), .B(n1359), .Z(c[338]) );
  XNOR U1704 ( .A(b[339]), .B(a[339]), .Z(n1364) );
  OR U1705 ( .A(b[338]), .B(a[338]), .Z(n1362) );
  OR U1706 ( .A(n1360), .B(n1359), .Z(n1361) );
  AND U1707 ( .A(n1362), .B(n1361), .Z(n1363) );
  XNOR U1708 ( .A(n1364), .B(n1363), .Z(c[339]) );
  XNOR U1709 ( .A(b[340]), .B(a[340]), .Z(n1368) );
  OR U1710 ( .A(b[339]), .B(a[339]), .Z(n1366) );
  OR U1711 ( .A(n1364), .B(n1363), .Z(n1365) );
  AND U1712 ( .A(n1366), .B(n1365), .Z(n1367) );
  XNOR U1713 ( .A(n1368), .B(n1367), .Z(c[340]) );
  XNOR U1714 ( .A(b[341]), .B(a[341]), .Z(n1372) );
  OR U1715 ( .A(b[340]), .B(a[340]), .Z(n1370) );
  OR U1716 ( .A(n1368), .B(n1367), .Z(n1369) );
  AND U1717 ( .A(n1370), .B(n1369), .Z(n1371) );
  XNOR U1718 ( .A(n1372), .B(n1371), .Z(c[341]) );
  XNOR U1719 ( .A(b[342]), .B(a[342]), .Z(n1376) );
  OR U1720 ( .A(b[341]), .B(a[341]), .Z(n1374) );
  OR U1721 ( .A(n1372), .B(n1371), .Z(n1373) );
  AND U1722 ( .A(n1374), .B(n1373), .Z(n1375) );
  XNOR U1723 ( .A(n1376), .B(n1375), .Z(c[342]) );
  XNOR U1724 ( .A(b[343]), .B(a[343]), .Z(n1380) );
  OR U1725 ( .A(b[342]), .B(a[342]), .Z(n1378) );
  OR U1726 ( .A(n1376), .B(n1375), .Z(n1377) );
  AND U1727 ( .A(n1378), .B(n1377), .Z(n1379) );
  XNOR U1728 ( .A(n1380), .B(n1379), .Z(c[343]) );
  XNOR U1729 ( .A(b[344]), .B(a[344]), .Z(n1384) );
  OR U1730 ( .A(b[343]), .B(a[343]), .Z(n1382) );
  OR U1731 ( .A(n1380), .B(n1379), .Z(n1381) );
  AND U1732 ( .A(n1382), .B(n1381), .Z(n1383) );
  XNOR U1733 ( .A(n1384), .B(n1383), .Z(c[344]) );
  XNOR U1734 ( .A(b[345]), .B(a[345]), .Z(n1388) );
  OR U1735 ( .A(b[344]), .B(a[344]), .Z(n1386) );
  OR U1736 ( .A(n1384), .B(n1383), .Z(n1385) );
  AND U1737 ( .A(n1386), .B(n1385), .Z(n1387) );
  XNOR U1738 ( .A(n1388), .B(n1387), .Z(c[345]) );
  XNOR U1739 ( .A(b[346]), .B(a[346]), .Z(n1392) );
  OR U1740 ( .A(b[345]), .B(a[345]), .Z(n1390) );
  OR U1741 ( .A(n1388), .B(n1387), .Z(n1389) );
  AND U1742 ( .A(n1390), .B(n1389), .Z(n1391) );
  XNOR U1743 ( .A(n1392), .B(n1391), .Z(c[346]) );
  XNOR U1744 ( .A(b[347]), .B(a[347]), .Z(n1396) );
  OR U1745 ( .A(b[346]), .B(a[346]), .Z(n1394) );
  OR U1746 ( .A(n1392), .B(n1391), .Z(n1393) );
  AND U1747 ( .A(n1394), .B(n1393), .Z(n1395) );
  XNOR U1748 ( .A(n1396), .B(n1395), .Z(c[347]) );
  XNOR U1749 ( .A(b[348]), .B(a[348]), .Z(n1400) );
  OR U1750 ( .A(b[347]), .B(a[347]), .Z(n1398) );
  OR U1751 ( .A(n1396), .B(n1395), .Z(n1397) );
  AND U1752 ( .A(n1398), .B(n1397), .Z(n1399) );
  XNOR U1753 ( .A(n1400), .B(n1399), .Z(c[348]) );
  XNOR U1754 ( .A(b[349]), .B(a[349]), .Z(n1404) );
  OR U1755 ( .A(b[348]), .B(a[348]), .Z(n1402) );
  OR U1756 ( .A(n1400), .B(n1399), .Z(n1401) );
  AND U1757 ( .A(n1402), .B(n1401), .Z(n1403) );
  XNOR U1758 ( .A(n1404), .B(n1403), .Z(c[349]) );
  XNOR U1759 ( .A(b[350]), .B(a[350]), .Z(n1408) );
  OR U1760 ( .A(b[349]), .B(a[349]), .Z(n1406) );
  OR U1761 ( .A(n1404), .B(n1403), .Z(n1405) );
  AND U1762 ( .A(n1406), .B(n1405), .Z(n1407) );
  XNOR U1763 ( .A(n1408), .B(n1407), .Z(c[350]) );
  XNOR U1764 ( .A(b[351]), .B(a[351]), .Z(n1412) );
  OR U1765 ( .A(b[350]), .B(a[350]), .Z(n1410) );
  OR U1766 ( .A(n1408), .B(n1407), .Z(n1409) );
  AND U1767 ( .A(n1410), .B(n1409), .Z(n1411) );
  XNOR U1768 ( .A(n1412), .B(n1411), .Z(c[351]) );
  XNOR U1769 ( .A(b[352]), .B(a[352]), .Z(n1416) );
  OR U1770 ( .A(b[351]), .B(a[351]), .Z(n1414) );
  OR U1771 ( .A(n1412), .B(n1411), .Z(n1413) );
  AND U1772 ( .A(n1414), .B(n1413), .Z(n1415) );
  XNOR U1773 ( .A(n1416), .B(n1415), .Z(c[352]) );
  XNOR U1774 ( .A(b[353]), .B(a[353]), .Z(n1420) );
  OR U1775 ( .A(b[352]), .B(a[352]), .Z(n1418) );
  OR U1776 ( .A(n1416), .B(n1415), .Z(n1417) );
  AND U1777 ( .A(n1418), .B(n1417), .Z(n1419) );
  XNOR U1778 ( .A(n1420), .B(n1419), .Z(c[353]) );
  OR U1779 ( .A(b[353]), .B(a[353]), .Z(n1422) );
  OR U1780 ( .A(n1420), .B(n1419), .Z(n1421) );
  NAND U1781 ( .A(n1422), .B(n1421), .Z(n1424) );
  XOR U1782 ( .A(a[354]), .B(b[354]), .Z(n1423) );
  XNOR U1783 ( .A(n1424), .B(n1423), .Z(c[354]) );
  XNOR U1784 ( .A(b[355]), .B(a[355]), .Z(n1428) );
  NAND U1785 ( .A(b[354]), .B(a[354]), .Z(n1426) );
  NANDN U1786 ( .A(n1424), .B(n1423), .Z(n1425) );
  NAND U1787 ( .A(n1426), .B(n1425), .Z(n1427) );
  XNOR U1788 ( .A(n1428), .B(n1427), .Z(c[355]) );
  XNOR U1789 ( .A(b[356]), .B(a[356]), .Z(n1432) );
  OR U1790 ( .A(b[355]), .B(a[355]), .Z(n1430) );
  OR U1791 ( .A(n1428), .B(n1427), .Z(n1429) );
  AND U1792 ( .A(n1430), .B(n1429), .Z(n1431) );
  XNOR U1793 ( .A(n1432), .B(n1431), .Z(c[356]) );
  OR U1794 ( .A(b[356]), .B(a[356]), .Z(n1434) );
  OR U1795 ( .A(n1432), .B(n1431), .Z(n1433) );
  NAND U1796 ( .A(n1434), .B(n1433), .Z(n1436) );
  XOR U1797 ( .A(a[357]), .B(b[357]), .Z(n1435) );
  XNOR U1798 ( .A(n1436), .B(n1435), .Z(c[357]) );
  XNOR U1799 ( .A(b[358]), .B(a[358]), .Z(n1440) );
  NAND U1800 ( .A(b[357]), .B(a[357]), .Z(n1438) );
  NANDN U1801 ( .A(n1436), .B(n1435), .Z(n1437) );
  NAND U1802 ( .A(n1438), .B(n1437), .Z(n1439) );
  XNOR U1803 ( .A(n1440), .B(n1439), .Z(c[358]) );
  OR U1804 ( .A(b[358]), .B(a[358]), .Z(n1442) );
  OR U1805 ( .A(n1440), .B(n1439), .Z(n1441) );
  NAND U1806 ( .A(n1442), .B(n1441), .Z(n1444) );
  XOR U1807 ( .A(a[359]), .B(b[359]), .Z(n1443) );
  XNOR U1808 ( .A(n1444), .B(n1443), .Z(c[359]) );
  XOR U1809 ( .A(a[360]), .B(b[360]), .Z(n1447) );
  NAND U1810 ( .A(b[359]), .B(a[359]), .Z(n1446) );
  NANDN U1811 ( .A(n1444), .B(n1443), .Z(n1445) );
  AND U1812 ( .A(n1446), .B(n1445), .Z(n1448) );
  XNOR U1813 ( .A(n1447), .B(n1448), .Z(c[360]) );
  XNOR U1814 ( .A(b[361]), .B(a[361]), .Z(n1452) );
  NAND U1815 ( .A(b[360]), .B(a[360]), .Z(n1450) );
  NANDN U1816 ( .A(n1448), .B(n1447), .Z(n1449) );
  NAND U1817 ( .A(n1450), .B(n1449), .Z(n1451) );
  XNOR U1818 ( .A(n1452), .B(n1451), .Z(c[361]) );
  OR U1819 ( .A(b[361]), .B(a[361]), .Z(n1454) );
  OR U1820 ( .A(n1452), .B(n1451), .Z(n1453) );
  NAND U1821 ( .A(n1454), .B(n1453), .Z(n1456) );
  XOR U1822 ( .A(a[362]), .B(b[362]), .Z(n1455) );
  XNOR U1823 ( .A(n1456), .B(n1455), .Z(c[362]) );
  XOR U1824 ( .A(a[363]), .B(b[363]), .Z(n1459) );
  NAND U1825 ( .A(b[362]), .B(a[362]), .Z(n1458) );
  NANDN U1826 ( .A(n1456), .B(n1455), .Z(n1457) );
  AND U1827 ( .A(n1458), .B(n1457), .Z(n1460) );
  XNOR U1828 ( .A(n1459), .B(n1460), .Z(c[363]) );
  XNOR U1829 ( .A(b[364]), .B(a[364]), .Z(n1464) );
  NAND U1830 ( .A(b[363]), .B(a[363]), .Z(n1462) );
  NANDN U1831 ( .A(n1460), .B(n1459), .Z(n1461) );
  NAND U1832 ( .A(n1462), .B(n1461), .Z(n1463) );
  XNOR U1833 ( .A(n1464), .B(n1463), .Z(c[364]) );
  OR U1834 ( .A(b[364]), .B(a[364]), .Z(n1466) );
  OR U1835 ( .A(n1464), .B(n1463), .Z(n1465) );
  NAND U1836 ( .A(n1466), .B(n1465), .Z(n1468) );
  XOR U1837 ( .A(a[365]), .B(b[365]), .Z(n1467) );
  XNOR U1838 ( .A(n1468), .B(n1467), .Z(c[365]) );
  XOR U1839 ( .A(a[366]), .B(b[366]), .Z(n1471) );
  NAND U1840 ( .A(b[365]), .B(a[365]), .Z(n1470) );
  NANDN U1841 ( .A(n1468), .B(n1467), .Z(n1469) );
  AND U1842 ( .A(n1470), .B(n1469), .Z(n1472) );
  XNOR U1843 ( .A(n1471), .B(n1472), .Z(c[366]) );
  NAND U1844 ( .A(b[366]), .B(a[366]), .Z(n1474) );
  NANDN U1845 ( .A(n1472), .B(n1471), .Z(n1473) );
  NAND U1846 ( .A(n1474), .B(n1473), .Z(n1476) );
  XNOR U1847 ( .A(b[367]), .B(a[367]), .Z(n1475) );
  XNOR U1848 ( .A(n1476), .B(n1475), .Z(c[367]) );
  XNOR U1849 ( .A(b[368]), .B(a[368]), .Z(n1480) );
  OR U1850 ( .A(b[367]), .B(a[367]), .Z(n1478) );
  OR U1851 ( .A(n1476), .B(n1475), .Z(n1477) );
  AND U1852 ( .A(n1478), .B(n1477), .Z(n1479) );
  XNOR U1853 ( .A(n1480), .B(n1479), .Z(c[368]) );
  XNOR U1854 ( .A(b[369]), .B(a[369]), .Z(n1484) );
  OR U1855 ( .A(b[368]), .B(a[368]), .Z(n1482) );
  OR U1856 ( .A(n1480), .B(n1479), .Z(n1481) );
  AND U1857 ( .A(n1482), .B(n1481), .Z(n1483) );
  XNOR U1858 ( .A(n1484), .B(n1483), .Z(c[369]) );
  XNOR U1859 ( .A(b[370]), .B(a[370]), .Z(n1488) );
  OR U1860 ( .A(b[369]), .B(a[369]), .Z(n1486) );
  OR U1861 ( .A(n1484), .B(n1483), .Z(n1485) );
  AND U1862 ( .A(n1486), .B(n1485), .Z(n1487) );
  XNOR U1863 ( .A(n1488), .B(n1487), .Z(c[370]) );
  XNOR U1864 ( .A(b[371]), .B(a[371]), .Z(n1492) );
  OR U1865 ( .A(b[370]), .B(a[370]), .Z(n1490) );
  OR U1866 ( .A(n1488), .B(n1487), .Z(n1489) );
  AND U1867 ( .A(n1490), .B(n1489), .Z(n1491) );
  XNOR U1868 ( .A(n1492), .B(n1491), .Z(c[371]) );
  XNOR U1869 ( .A(b[372]), .B(a[372]), .Z(n1496) );
  OR U1870 ( .A(b[371]), .B(a[371]), .Z(n1494) );
  OR U1871 ( .A(n1492), .B(n1491), .Z(n1493) );
  AND U1872 ( .A(n1494), .B(n1493), .Z(n1495) );
  XNOR U1873 ( .A(n1496), .B(n1495), .Z(c[372]) );
  XNOR U1874 ( .A(b[373]), .B(a[373]), .Z(n1500) );
  OR U1875 ( .A(b[372]), .B(a[372]), .Z(n1498) );
  OR U1876 ( .A(n1496), .B(n1495), .Z(n1497) );
  AND U1877 ( .A(n1498), .B(n1497), .Z(n1499) );
  XNOR U1878 ( .A(n1500), .B(n1499), .Z(c[373]) );
  XNOR U1879 ( .A(b[374]), .B(a[374]), .Z(n1504) );
  OR U1880 ( .A(b[373]), .B(a[373]), .Z(n1502) );
  OR U1881 ( .A(n1500), .B(n1499), .Z(n1501) );
  AND U1882 ( .A(n1502), .B(n1501), .Z(n1503) );
  XNOR U1883 ( .A(n1504), .B(n1503), .Z(c[374]) );
  XNOR U1884 ( .A(b[375]), .B(a[375]), .Z(n1508) );
  OR U1885 ( .A(b[374]), .B(a[374]), .Z(n1506) );
  OR U1886 ( .A(n1504), .B(n1503), .Z(n1505) );
  AND U1887 ( .A(n1506), .B(n1505), .Z(n1507) );
  XNOR U1888 ( .A(n1508), .B(n1507), .Z(c[375]) );
  XNOR U1889 ( .A(b[376]), .B(a[376]), .Z(n1512) );
  OR U1890 ( .A(b[375]), .B(a[375]), .Z(n1510) );
  OR U1891 ( .A(n1508), .B(n1507), .Z(n1509) );
  AND U1892 ( .A(n1510), .B(n1509), .Z(n1511) );
  XNOR U1893 ( .A(n1512), .B(n1511), .Z(c[376]) );
  XNOR U1894 ( .A(b[377]), .B(a[377]), .Z(n1516) );
  OR U1895 ( .A(b[376]), .B(a[376]), .Z(n1514) );
  OR U1896 ( .A(n1512), .B(n1511), .Z(n1513) );
  AND U1897 ( .A(n1514), .B(n1513), .Z(n1515) );
  XNOR U1898 ( .A(n1516), .B(n1515), .Z(c[377]) );
  XNOR U1899 ( .A(b[378]), .B(a[378]), .Z(n1520) );
  OR U1900 ( .A(b[377]), .B(a[377]), .Z(n1518) );
  OR U1901 ( .A(n1516), .B(n1515), .Z(n1517) );
  AND U1902 ( .A(n1518), .B(n1517), .Z(n1519) );
  XNOR U1903 ( .A(n1520), .B(n1519), .Z(c[378]) );
  XNOR U1904 ( .A(b[379]), .B(a[379]), .Z(n1524) );
  OR U1905 ( .A(b[378]), .B(a[378]), .Z(n1522) );
  OR U1906 ( .A(n1520), .B(n1519), .Z(n1521) );
  AND U1907 ( .A(n1522), .B(n1521), .Z(n1523) );
  XNOR U1908 ( .A(n1524), .B(n1523), .Z(c[379]) );
  XNOR U1909 ( .A(b[380]), .B(a[380]), .Z(n1528) );
  OR U1910 ( .A(b[379]), .B(a[379]), .Z(n1526) );
  OR U1911 ( .A(n1524), .B(n1523), .Z(n1525) );
  AND U1912 ( .A(n1526), .B(n1525), .Z(n1527) );
  XNOR U1913 ( .A(n1528), .B(n1527), .Z(c[380]) );
  OR U1914 ( .A(b[380]), .B(a[380]), .Z(n1530) );
  OR U1915 ( .A(n1528), .B(n1527), .Z(n1529) );
  NAND U1916 ( .A(n1530), .B(n1529), .Z(n1532) );
  XOR U1917 ( .A(a[381]), .B(b[381]), .Z(n1531) );
  XNOR U1918 ( .A(n1532), .B(n1531), .Z(c[381]) );
  XOR U1919 ( .A(a[382]), .B(b[382]), .Z(n1535) );
  NAND U1920 ( .A(b[381]), .B(a[381]), .Z(n1534) );
  NANDN U1921 ( .A(n1532), .B(n1531), .Z(n1533) );
  AND U1922 ( .A(n1534), .B(n1533), .Z(n1536) );
  XNOR U1923 ( .A(n1535), .B(n1536), .Z(c[382]) );
  XNOR U1924 ( .A(b[383]), .B(a[383]), .Z(n1540) );
  NAND U1925 ( .A(b[382]), .B(a[382]), .Z(n1538) );
  NANDN U1926 ( .A(n1536), .B(n1535), .Z(n1537) );
  NAND U1927 ( .A(n1538), .B(n1537), .Z(n1539) );
  XNOR U1928 ( .A(n1540), .B(n1539), .Z(c[383]) );
  OR U1929 ( .A(b[383]), .B(a[383]), .Z(n1542) );
  OR U1930 ( .A(n1540), .B(n1539), .Z(n1541) );
  NAND U1931 ( .A(n1542), .B(n1541), .Z(n1544) );
  XOR U1932 ( .A(a[384]), .B(b[384]), .Z(n1543) );
  XNOR U1933 ( .A(n1544), .B(n1543), .Z(c[384]) );
  XOR U1934 ( .A(a[385]), .B(b[385]), .Z(n1547) );
  NAND U1935 ( .A(b[384]), .B(a[384]), .Z(n1546) );
  NANDN U1936 ( .A(n1544), .B(n1543), .Z(n1545) );
  AND U1937 ( .A(n1546), .B(n1545), .Z(n1548) );
  XNOR U1938 ( .A(n1547), .B(n1548), .Z(c[385]) );
  NAND U1939 ( .A(b[385]), .B(a[385]), .Z(n1550) );
  NANDN U1940 ( .A(n1548), .B(n1547), .Z(n1549) );
  NAND U1941 ( .A(n1550), .B(n1549), .Z(n1552) );
  XOR U1942 ( .A(a[386]), .B(b[386]), .Z(n1551) );
  XOR U1943 ( .A(n1552), .B(n1551), .Z(c[386]) );
  XOR U1944 ( .A(a[387]), .B(b[387]), .Z(n1554) );
  XOR U1945 ( .A(n1553), .B(n1554), .Z(c[387]) );
  XOR U1946 ( .A(a[388]), .B(b[388]), .Z(n1557) );
  NAND U1947 ( .A(b[387]), .B(a[387]), .Z(n1556) );
  NAND U1948 ( .A(n1554), .B(n1553), .Z(n1555) );
  AND U1949 ( .A(n1556), .B(n1555), .Z(n1558) );
  XNOR U1950 ( .A(n1557), .B(n1558), .Z(c[388]) );
  NAND U1951 ( .A(b[388]), .B(a[388]), .Z(n1560) );
  NANDN U1952 ( .A(n1558), .B(n1557), .Z(n1559) );
  NAND U1953 ( .A(n1560), .B(n1559), .Z(n1562) );
  XNOR U1954 ( .A(b[389]), .B(a[389]), .Z(n1561) );
  XNOR U1955 ( .A(n1562), .B(n1561), .Z(c[389]) );
  OR U1956 ( .A(b[389]), .B(a[389]), .Z(n1564) );
  OR U1957 ( .A(n1562), .B(n1561), .Z(n1563) );
  NAND U1958 ( .A(n1564), .B(n1563), .Z(n1566) );
  XOR U1959 ( .A(a[390]), .B(b[390]), .Z(n1565) );
  XNOR U1960 ( .A(n1566), .B(n1565), .Z(c[390]) );
  XOR U1961 ( .A(a[391]), .B(b[391]), .Z(n1569) );
  NAND U1962 ( .A(b[390]), .B(a[390]), .Z(n1568) );
  NANDN U1963 ( .A(n1566), .B(n1565), .Z(n1567) );
  AND U1964 ( .A(n1568), .B(n1567), .Z(n1570) );
  XNOR U1965 ( .A(n1569), .B(n1570), .Z(c[391]) );
  XOR U1966 ( .A(a[392]), .B(b[392]), .Z(n1573) );
  NAND U1967 ( .A(b[391]), .B(a[391]), .Z(n1572) );
  NANDN U1968 ( .A(n1570), .B(n1569), .Z(n1571) );
  AND U1969 ( .A(n1572), .B(n1571), .Z(n1574) );
  XNOR U1970 ( .A(n1573), .B(n1574), .Z(c[392]) );
  XOR U1971 ( .A(a[393]), .B(b[393]), .Z(n1577) );
  NAND U1972 ( .A(b[392]), .B(a[392]), .Z(n1576) );
  NANDN U1973 ( .A(n1574), .B(n1573), .Z(n1575) );
  AND U1974 ( .A(n1576), .B(n1575), .Z(n1578) );
  XNOR U1975 ( .A(n1577), .B(n1578), .Z(c[393]) );
  XOR U1976 ( .A(a[394]), .B(b[394]), .Z(n1581) );
  NAND U1977 ( .A(b[393]), .B(a[393]), .Z(n1580) );
  NANDN U1978 ( .A(n1578), .B(n1577), .Z(n1579) );
  AND U1979 ( .A(n1580), .B(n1579), .Z(n1582) );
  XNOR U1980 ( .A(n1581), .B(n1582), .Z(c[394]) );
  XOR U1981 ( .A(a[395]), .B(b[395]), .Z(n1585) );
  NAND U1982 ( .A(b[394]), .B(a[394]), .Z(n1584) );
  NANDN U1983 ( .A(n1582), .B(n1581), .Z(n1583) );
  AND U1984 ( .A(n1584), .B(n1583), .Z(n1586) );
  XNOR U1985 ( .A(n1585), .B(n1586), .Z(c[395]) );
  XOR U1986 ( .A(a[396]), .B(b[396]), .Z(n1589) );
  NAND U1987 ( .A(b[395]), .B(a[395]), .Z(n1588) );
  NANDN U1988 ( .A(n1586), .B(n1585), .Z(n1587) );
  AND U1989 ( .A(n1588), .B(n1587), .Z(n1590) );
  XNOR U1990 ( .A(n1589), .B(n1590), .Z(c[396]) );
  XOR U1991 ( .A(a[397]), .B(b[397]), .Z(n1593) );
  NAND U1992 ( .A(b[396]), .B(a[396]), .Z(n1592) );
  NANDN U1993 ( .A(n1590), .B(n1589), .Z(n1591) );
  AND U1994 ( .A(n1592), .B(n1591), .Z(n1594) );
  XNOR U1995 ( .A(n1593), .B(n1594), .Z(c[397]) );
  XOR U1996 ( .A(a[398]), .B(b[398]), .Z(n1597) );
  NAND U1997 ( .A(b[397]), .B(a[397]), .Z(n1596) );
  NANDN U1998 ( .A(n1594), .B(n1593), .Z(n1595) );
  AND U1999 ( .A(n1596), .B(n1595), .Z(n1598) );
  XNOR U2000 ( .A(n1597), .B(n1598), .Z(c[398]) );
  NAND U2001 ( .A(b[398]), .B(a[398]), .Z(n1600) );
  NANDN U2002 ( .A(n1598), .B(n1597), .Z(n1599) );
  NAND U2003 ( .A(n1600), .B(n1599), .Z(n1602) );
  XNOR U2004 ( .A(b[399]), .B(a[399]), .Z(n1601) );
  XNOR U2005 ( .A(n1602), .B(n1601), .Z(c[399]) );
  XOR U2006 ( .A(a[400]), .B(b[400]), .Z(n1605) );
  OR U2007 ( .A(b[399]), .B(a[399]), .Z(n1604) );
  OR U2008 ( .A(n1602), .B(n1601), .Z(n1603) );
  NAND U2009 ( .A(n1604), .B(n1603), .Z(n1606) );
  XNOR U2010 ( .A(n1605), .B(n1606), .Z(c[400]) );
  NAND U2011 ( .A(b[400]), .B(a[400]), .Z(n1608) );
  NANDN U2012 ( .A(n1606), .B(n1605), .Z(n1607) );
  NAND U2013 ( .A(n1608), .B(n1607), .Z(n1610) );
  XNOR U2014 ( .A(b[401]), .B(a[401]), .Z(n1609) );
  XNOR U2015 ( .A(n1610), .B(n1609), .Z(c[401]) );
  XNOR U2016 ( .A(b[402]), .B(a[402]), .Z(n1614) );
  OR U2017 ( .A(b[401]), .B(a[401]), .Z(n1612) );
  OR U2018 ( .A(n1610), .B(n1609), .Z(n1611) );
  AND U2019 ( .A(n1612), .B(n1611), .Z(n1613) );
  XNOR U2020 ( .A(n1614), .B(n1613), .Z(c[402]) );
  XNOR U2021 ( .A(b[403]), .B(a[403]), .Z(n1618) );
  OR U2022 ( .A(b[402]), .B(a[402]), .Z(n1616) );
  OR U2023 ( .A(n1614), .B(n1613), .Z(n1615) );
  AND U2024 ( .A(n1616), .B(n1615), .Z(n1617) );
  XNOR U2025 ( .A(n1618), .B(n1617), .Z(c[403]) );
  XNOR U2026 ( .A(b[404]), .B(a[404]), .Z(n1622) );
  OR U2027 ( .A(b[403]), .B(a[403]), .Z(n1620) );
  OR U2028 ( .A(n1618), .B(n1617), .Z(n1619) );
  AND U2029 ( .A(n1620), .B(n1619), .Z(n1621) );
  XNOR U2030 ( .A(n1622), .B(n1621), .Z(c[404]) );
  XNOR U2031 ( .A(b[405]), .B(a[405]), .Z(n1626) );
  OR U2032 ( .A(b[404]), .B(a[404]), .Z(n1624) );
  OR U2033 ( .A(n1622), .B(n1621), .Z(n1623) );
  AND U2034 ( .A(n1624), .B(n1623), .Z(n1625) );
  XNOR U2035 ( .A(n1626), .B(n1625), .Z(c[405]) );
  XNOR U2036 ( .A(b[406]), .B(a[406]), .Z(n1630) );
  OR U2037 ( .A(b[405]), .B(a[405]), .Z(n1628) );
  OR U2038 ( .A(n1626), .B(n1625), .Z(n1627) );
  AND U2039 ( .A(n1628), .B(n1627), .Z(n1629) );
  XNOR U2040 ( .A(n1630), .B(n1629), .Z(c[406]) );
  XNOR U2041 ( .A(b[407]), .B(a[407]), .Z(n1634) );
  OR U2042 ( .A(b[406]), .B(a[406]), .Z(n1632) );
  OR U2043 ( .A(n1630), .B(n1629), .Z(n1631) );
  AND U2044 ( .A(n1632), .B(n1631), .Z(n1633) );
  XNOR U2045 ( .A(n1634), .B(n1633), .Z(c[407]) );
  XNOR U2046 ( .A(b[408]), .B(a[408]), .Z(n1638) );
  OR U2047 ( .A(b[407]), .B(a[407]), .Z(n1636) );
  OR U2048 ( .A(n1634), .B(n1633), .Z(n1635) );
  AND U2049 ( .A(n1636), .B(n1635), .Z(n1637) );
  XNOR U2050 ( .A(n1638), .B(n1637), .Z(c[408]) );
  XNOR U2051 ( .A(b[409]), .B(a[409]), .Z(n1642) );
  OR U2052 ( .A(b[408]), .B(a[408]), .Z(n1640) );
  OR U2053 ( .A(n1638), .B(n1637), .Z(n1639) );
  AND U2054 ( .A(n1640), .B(n1639), .Z(n1641) );
  XNOR U2055 ( .A(n1642), .B(n1641), .Z(c[409]) );
  XNOR U2056 ( .A(b[410]), .B(a[410]), .Z(n1646) );
  OR U2057 ( .A(b[409]), .B(a[409]), .Z(n1644) );
  OR U2058 ( .A(n1642), .B(n1641), .Z(n1643) );
  AND U2059 ( .A(n1644), .B(n1643), .Z(n1645) );
  XNOR U2060 ( .A(n1646), .B(n1645), .Z(c[410]) );
  XNOR U2061 ( .A(b[411]), .B(a[411]), .Z(n1650) );
  OR U2062 ( .A(b[410]), .B(a[410]), .Z(n1648) );
  OR U2063 ( .A(n1646), .B(n1645), .Z(n1647) );
  AND U2064 ( .A(n1648), .B(n1647), .Z(n1649) );
  XNOR U2065 ( .A(n1650), .B(n1649), .Z(c[411]) );
  XNOR U2066 ( .A(b[412]), .B(a[412]), .Z(n1654) );
  OR U2067 ( .A(b[411]), .B(a[411]), .Z(n1652) );
  OR U2068 ( .A(n1650), .B(n1649), .Z(n1651) );
  AND U2069 ( .A(n1652), .B(n1651), .Z(n1653) );
  XNOR U2070 ( .A(n1654), .B(n1653), .Z(c[412]) );
  XNOR U2071 ( .A(b[413]), .B(a[413]), .Z(n1658) );
  OR U2072 ( .A(b[412]), .B(a[412]), .Z(n1656) );
  OR U2073 ( .A(n1654), .B(n1653), .Z(n1655) );
  AND U2074 ( .A(n1656), .B(n1655), .Z(n1657) );
  XNOR U2075 ( .A(n1658), .B(n1657), .Z(c[413]) );
  XNOR U2076 ( .A(b[414]), .B(a[414]), .Z(n1662) );
  OR U2077 ( .A(b[413]), .B(a[413]), .Z(n1660) );
  OR U2078 ( .A(n1658), .B(n1657), .Z(n1659) );
  AND U2079 ( .A(n1660), .B(n1659), .Z(n1661) );
  XNOR U2080 ( .A(n1662), .B(n1661), .Z(c[414]) );
  XNOR U2081 ( .A(b[415]), .B(a[415]), .Z(n1666) );
  OR U2082 ( .A(b[414]), .B(a[414]), .Z(n1664) );
  OR U2083 ( .A(n1662), .B(n1661), .Z(n1663) );
  AND U2084 ( .A(n1664), .B(n1663), .Z(n1665) );
  XNOR U2085 ( .A(n1666), .B(n1665), .Z(c[415]) );
  OR U2086 ( .A(b[415]), .B(a[415]), .Z(n1668) );
  OR U2087 ( .A(n1666), .B(n1665), .Z(n1667) );
  NAND U2088 ( .A(n1668), .B(n1667), .Z(n1670) );
  XOR U2089 ( .A(a[416]), .B(b[416]), .Z(n1669) );
  XNOR U2090 ( .A(n1670), .B(n1669), .Z(c[416]) );
  XOR U2091 ( .A(a[417]), .B(b[417]), .Z(n1673) );
  NAND U2092 ( .A(b[416]), .B(a[416]), .Z(n1672) );
  NANDN U2093 ( .A(n1670), .B(n1669), .Z(n1671) );
  AND U2094 ( .A(n1672), .B(n1671), .Z(n1674) );
  XNOR U2095 ( .A(n1673), .B(n1674), .Z(c[417]) );
  XNOR U2096 ( .A(b[418]), .B(a[418]), .Z(n1678) );
  NAND U2097 ( .A(b[417]), .B(a[417]), .Z(n1676) );
  NANDN U2098 ( .A(n1674), .B(n1673), .Z(n1675) );
  NAND U2099 ( .A(n1676), .B(n1675), .Z(n1677) );
  XNOR U2100 ( .A(n1678), .B(n1677), .Z(c[418]) );
  OR U2101 ( .A(b[418]), .B(a[418]), .Z(n1680) );
  OR U2102 ( .A(n1678), .B(n1677), .Z(n1679) );
  NAND U2103 ( .A(n1680), .B(n1679), .Z(n1682) );
  XOR U2104 ( .A(a[419]), .B(b[419]), .Z(n1681) );
  XNOR U2105 ( .A(n1682), .B(n1681), .Z(c[419]) );
  XOR U2106 ( .A(a[420]), .B(b[420]), .Z(n1685) );
  NAND U2107 ( .A(b[419]), .B(a[419]), .Z(n1684) );
  NANDN U2108 ( .A(n1682), .B(n1681), .Z(n1683) );
  AND U2109 ( .A(n1684), .B(n1683), .Z(n1686) );
  XNOR U2110 ( .A(n1685), .B(n1686), .Z(c[420]) );
  NAND U2111 ( .A(b[420]), .B(a[420]), .Z(n1688) );
  NANDN U2112 ( .A(n1686), .B(n1685), .Z(n1687) );
  NAND U2113 ( .A(n1688), .B(n1687), .Z(n1690) );
  XNOR U2114 ( .A(b[421]), .B(a[421]), .Z(n1689) );
  XNOR U2115 ( .A(n1690), .B(n1689), .Z(c[421]) );
  XNOR U2116 ( .A(b[422]), .B(a[422]), .Z(n1694) );
  OR U2117 ( .A(b[421]), .B(a[421]), .Z(n1692) );
  OR U2118 ( .A(n1690), .B(n1689), .Z(n1691) );
  AND U2119 ( .A(n1692), .B(n1691), .Z(n1693) );
  XNOR U2120 ( .A(n1694), .B(n1693), .Z(c[422]) );
  XNOR U2121 ( .A(b[423]), .B(a[423]), .Z(n1698) );
  OR U2122 ( .A(b[422]), .B(a[422]), .Z(n1696) );
  OR U2123 ( .A(n1694), .B(n1693), .Z(n1695) );
  AND U2124 ( .A(n1696), .B(n1695), .Z(n1697) );
  XNOR U2125 ( .A(n1698), .B(n1697), .Z(c[423]) );
  XNOR U2126 ( .A(b[424]), .B(a[424]), .Z(n1702) );
  OR U2127 ( .A(b[423]), .B(a[423]), .Z(n1700) );
  OR U2128 ( .A(n1698), .B(n1697), .Z(n1699) );
  AND U2129 ( .A(n1700), .B(n1699), .Z(n1701) );
  XNOR U2130 ( .A(n1702), .B(n1701), .Z(c[424]) );
  XNOR U2131 ( .A(b[425]), .B(a[425]), .Z(n1706) );
  OR U2132 ( .A(b[424]), .B(a[424]), .Z(n1704) );
  OR U2133 ( .A(n1702), .B(n1701), .Z(n1703) );
  AND U2134 ( .A(n1704), .B(n1703), .Z(n1705) );
  XNOR U2135 ( .A(n1706), .B(n1705), .Z(c[425]) );
  XNOR U2136 ( .A(b[426]), .B(a[426]), .Z(n1710) );
  OR U2137 ( .A(b[425]), .B(a[425]), .Z(n1708) );
  OR U2138 ( .A(n1706), .B(n1705), .Z(n1707) );
  AND U2139 ( .A(n1708), .B(n1707), .Z(n1709) );
  XNOR U2140 ( .A(n1710), .B(n1709), .Z(c[426]) );
  OR U2141 ( .A(b[426]), .B(a[426]), .Z(n1712) );
  OR U2142 ( .A(n1710), .B(n1709), .Z(n1711) );
  NAND U2143 ( .A(n1712), .B(n1711), .Z(n1714) );
  XOR U2144 ( .A(a[427]), .B(b[427]), .Z(n1713) );
  XNOR U2145 ( .A(n1714), .B(n1713), .Z(c[427]) );
  XOR U2146 ( .A(a[428]), .B(b[428]), .Z(n1717) );
  NAND U2147 ( .A(b[427]), .B(a[427]), .Z(n1716) );
  NANDN U2148 ( .A(n1714), .B(n1713), .Z(n1715) );
  AND U2149 ( .A(n1716), .B(n1715), .Z(n1718) );
  XNOR U2150 ( .A(n1717), .B(n1718), .Z(c[428]) );
  XOR U2151 ( .A(a[429]), .B(b[429]), .Z(n1721) );
  NAND U2152 ( .A(b[428]), .B(a[428]), .Z(n1720) );
  NANDN U2153 ( .A(n1718), .B(n1717), .Z(n1719) );
  AND U2154 ( .A(n1720), .B(n1719), .Z(n1722) );
  XNOR U2155 ( .A(n1721), .B(n1722), .Z(c[429]) );
  XOR U2156 ( .A(a[430]), .B(b[430]), .Z(n1725) );
  NAND U2157 ( .A(b[429]), .B(a[429]), .Z(n1724) );
  NANDN U2158 ( .A(n1722), .B(n1721), .Z(n1723) );
  AND U2159 ( .A(n1724), .B(n1723), .Z(n1726) );
  XNOR U2160 ( .A(n1725), .B(n1726), .Z(c[430]) );
  XOR U2161 ( .A(a[431]), .B(b[431]), .Z(n1729) );
  NAND U2162 ( .A(b[430]), .B(a[430]), .Z(n1728) );
  NANDN U2163 ( .A(n1726), .B(n1725), .Z(n1727) );
  AND U2164 ( .A(n1728), .B(n1727), .Z(n1730) );
  XNOR U2165 ( .A(n1729), .B(n1730), .Z(c[431]) );
  XOR U2166 ( .A(a[432]), .B(b[432]), .Z(n1733) );
  NAND U2167 ( .A(b[431]), .B(a[431]), .Z(n1732) );
  NANDN U2168 ( .A(n1730), .B(n1729), .Z(n1731) );
  AND U2169 ( .A(n1732), .B(n1731), .Z(n1734) );
  XNOR U2170 ( .A(n1733), .B(n1734), .Z(c[432]) );
  XOR U2171 ( .A(a[433]), .B(b[433]), .Z(n1737) );
  NAND U2172 ( .A(b[432]), .B(a[432]), .Z(n1736) );
  NANDN U2173 ( .A(n1734), .B(n1733), .Z(n1735) );
  AND U2174 ( .A(n1736), .B(n1735), .Z(n1738) );
  XNOR U2175 ( .A(n1737), .B(n1738), .Z(c[433]) );
  XOR U2176 ( .A(a[434]), .B(b[434]), .Z(n1741) );
  NAND U2177 ( .A(b[433]), .B(a[433]), .Z(n1740) );
  NANDN U2178 ( .A(n1738), .B(n1737), .Z(n1739) );
  AND U2179 ( .A(n1740), .B(n1739), .Z(n1742) );
  XNOR U2180 ( .A(n1741), .B(n1742), .Z(c[434]) );
  XOR U2181 ( .A(a[435]), .B(b[435]), .Z(n1745) );
  NAND U2182 ( .A(b[434]), .B(a[434]), .Z(n1744) );
  NANDN U2183 ( .A(n1742), .B(n1741), .Z(n1743) );
  AND U2184 ( .A(n1744), .B(n1743), .Z(n1746) );
  XNOR U2185 ( .A(n1745), .B(n1746), .Z(c[435]) );
  XOR U2186 ( .A(a[436]), .B(b[436]), .Z(n1749) );
  NAND U2187 ( .A(b[435]), .B(a[435]), .Z(n1748) );
  NANDN U2188 ( .A(n1746), .B(n1745), .Z(n1747) );
  AND U2189 ( .A(n1748), .B(n1747), .Z(n1750) );
  XNOR U2190 ( .A(n1749), .B(n1750), .Z(c[436]) );
  XOR U2191 ( .A(a[437]), .B(b[437]), .Z(n1753) );
  NAND U2192 ( .A(b[436]), .B(a[436]), .Z(n1752) );
  NANDN U2193 ( .A(n1750), .B(n1749), .Z(n1751) );
  AND U2194 ( .A(n1752), .B(n1751), .Z(n1754) );
  XNOR U2195 ( .A(n1753), .B(n1754), .Z(c[437]) );
  XOR U2196 ( .A(a[438]), .B(b[438]), .Z(n1757) );
  NAND U2197 ( .A(b[437]), .B(a[437]), .Z(n1756) );
  NANDN U2198 ( .A(n1754), .B(n1753), .Z(n1755) );
  AND U2199 ( .A(n1756), .B(n1755), .Z(n1758) );
  XNOR U2200 ( .A(n1757), .B(n1758), .Z(c[438]) );
  XOR U2201 ( .A(a[439]), .B(b[439]), .Z(n1761) );
  NAND U2202 ( .A(b[438]), .B(a[438]), .Z(n1760) );
  NANDN U2203 ( .A(n1758), .B(n1757), .Z(n1759) );
  AND U2204 ( .A(n1760), .B(n1759), .Z(n1762) );
  XNOR U2205 ( .A(n1761), .B(n1762), .Z(c[439]) );
  XOR U2206 ( .A(a[440]), .B(b[440]), .Z(n1765) );
  NAND U2207 ( .A(b[439]), .B(a[439]), .Z(n1764) );
  NANDN U2208 ( .A(n1762), .B(n1761), .Z(n1763) );
  AND U2209 ( .A(n1764), .B(n1763), .Z(n1766) );
  XNOR U2210 ( .A(n1765), .B(n1766), .Z(c[440]) );
  XOR U2211 ( .A(a[441]), .B(b[441]), .Z(n1769) );
  NAND U2212 ( .A(b[440]), .B(a[440]), .Z(n1768) );
  NANDN U2213 ( .A(n1766), .B(n1765), .Z(n1767) );
  AND U2214 ( .A(n1768), .B(n1767), .Z(n1770) );
  XNOR U2215 ( .A(n1769), .B(n1770), .Z(c[441]) );
  XOR U2216 ( .A(a[442]), .B(b[442]), .Z(n1773) );
  NAND U2217 ( .A(b[441]), .B(a[441]), .Z(n1772) );
  NANDN U2218 ( .A(n1770), .B(n1769), .Z(n1771) );
  AND U2219 ( .A(n1772), .B(n1771), .Z(n1774) );
  XNOR U2220 ( .A(n1773), .B(n1774), .Z(c[442]) );
  XOR U2221 ( .A(a[443]), .B(b[443]), .Z(n1777) );
  NAND U2222 ( .A(b[442]), .B(a[442]), .Z(n1776) );
  NANDN U2223 ( .A(n1774), .B(n1773), .Z(n1775) );
  AND U2224 ( .A(n1776), .B(n1775), .Z(n1778) );
  XNOR U2225 ( .A(n1777), .B(n1778), .Z(c[443]) );
  XOR U2226 ( .A(a[444]), .B(b[444]), .Z(n1781) );
  NAND U2227 ( .A(b[443]), .B(a[443]), .Z(n1780) );
  NANDN U2228 ( .A(n1778), .B(n1777), .Z(n1779) );
  AND U2229 ( .A(n1780), .B(n1779), .Z(n1782) );
  XNOR U2230 ( .A(n1781), .B(n1782), .Z(c[444]) );
  NAND U2231 ( .A(b[444]), .B(a[444]), .Z(n1784) );
  NANDN U2232 ( .A(n1782), .B(n1781), .Z(n1783) );
  NAND U2233 ( .A(n1784), .B(n1783), .Z(n1786) );
  XNOR U2234 ( .A(b[445]), .B(a[445]), .Z(n1785) );
  XNOR U2235 ( .A(n1786), .B(n1785), .Z(c[445]) );
  XNOR U2236 ( .A(b[446]), .B(a[446]), .Z(n1790) );
  OR U2237 ( .A(b[445]), .B(a[445]), .Z(n1788) );
  OR U2238 ( .A(n1786), .B(n1785), .Z(n1787) );
  AND U2239 ( .A(n1788), .B(n1787), .Z(n1789) );
  XNOR U2240 ( .A(n1790), .B(n1789), .Z(c[446]) );
  XOR U2241 ( .A(a[447]), .B(b[447]), .Z(n1793) );
  OR U2242 ( .A(b[446]), .B(a[446]), .Z(n1792) );
  OR U2243 ( .A(n1790), .B(n1789), .Z(n1791) );
  NAND U2244 ( .A(n1792), .B(n1791), .Z(n1794) );
  XNOR U2245 ( .A(n1793), .B(n1794), .Z(c[447]) );
  NAND U2246 ( .A(b[447]), .B(a[447]), .Z(n1796) );
  NANDN U2247 ( .A(n1794), .B(n1793), .Z(n1795) );
  NAND U2248 ( .A(n1796), .B(n1795), .Z(n1798) );
  XNOR U2249 ( .A(b[448]), .B(a[448]), .Z(n1797) );
  XNOR U2250 ( .A(n1798), .B(n1797), .Z(c[448]) );
  XNOR U2251 ( .A(b[449]), .B(a[449]), .Z(n1802) );
  OR U2252 ( .A(b[448]), .B(a[448]), .Z(n1800) );
  OR U2253 ( .A(n1798), .B(n1797), .Z(n1799) );
  AND U2254 ( .A(n1800), .B(n1799), .Z(n1801) );
  XNOR U2255 ( .A(n1802), .B(n1801), .Z(c[449]) );
  XOR U2256 ( .A(a[450]), .B(b[450]), .Z(n1805) );
  OR U2257 ( .A(b[449]), .B(a[449]), .Z(n1804) );
  OR U2258 ( .A(n1802), .B(n1801), .Z(n1803) );
  NAND U2259 ( .A(n1804), .B(n1803), .Z(n1806) );
  XNOR U2260 ( .A(n1805), .B(n1806), .Z(c[450]) );
  NAND U2261 ( .A(b[450]), .B(a[450]), .Z(n1808) );
  NANDN U2262 ( .A(n1806), .B(n1805), .Z(n1807) );
  NAND U2263 ( .A(n1808), .B(n1807), .Z(n1810) );
  XNOR U2264 ( .A(b[451]), .B(a[451]), .Z(n1809) );
  XNOR U2265 ( .A(n1810), .B(n1809), .Z(c[451]) );
  XNOR U2266 ( .A(b[452]), .B(a[452]), .Z(n1814) );
  OR U2267 ( .A(b[451]), .B(a[451]), .Z(n1812) );
  OR U2268 ( .A(n1810), .B(n1809), .Z(n1811) );
  AND U2269 ( .A(n1812), .B(n1811), .Z(n1813) );
  XNOR U2270 ( .A(n1814), .B(n1813), .Z(c[452]) );
  XNOR U2271 ( .A(b[453]), .B(a[453]), .Z(n1818) );
  OR U2272 ( .A(b[452]), .B(a[452]), .Z(n1816) );
  OR U2273 ( .A(n1814), .B(n1813), .Z(n1815) );
  AND U2274 ( .A(n1816), .B(n1815), .Z(n1817) );
  XNOR U2275 ( .A(n1818), .B(n1817), .Z(c[453]) );
  XNOR U2276 ( .A(b[454]), .B(a[454]), .Z(n1822) );
  OR U2277 ( .A(b[453]), .B(a[453]), .Z(n1820) );
  OR U2278 ( .A(n1818), .B(n1817), .Z(n1819) );
  AND U2279 ( .A(n1820), .B(n1819), .Z(n1821) );
  XNOR U2280 ( .A(n1822), .B(n1821), .Z(c[454]) );
  XNOR U2281 ( .A(b[455]), .B(a[455]), .Z(n1826) );
  OR U2282 ( .A(b[454]), .B(a[454]), .Z(n1824) );
  OR U2283 ( .A(n1822), .B(n1821), .Z(n1823) );
  AND U2284 ( .A(n1824), .B(n1823), .Z(n1825) );
  XNOR U2285 ( .A(n1826), .B(n1825), .Z(c[455]) );
  XNOR U2286 ( .A(b[456]), .B(a[456]), .Z(n1830) );
  OR U2287 ( .A(b[455]), .B(a[455]), .Z(n1828) );
  OR U2288 ( .A(n1826), .B(n1825), .Z(n1827) );
  AND U2289 ( .A(n1828), .B(n1827), .Z(n1829) );
  XNOR U2290 ( .A(n1830), .B(n1829), .Z(c[456]) );
  XNOR U2291 ( .A(b[457]), .B(a[457]), .Z(n1834) );
  OR U2292 ( .A(b[456]), .B(a[456]), .Z(n1832) );
  OR U2293 ( .A(n1830), .B(n1829), .Z(n1831) );
  AND U2294 ( .A(n1832), .B(n1831), .Z(n1833) );
  XNOR U2295 ( .A(n1834), .B(n1833), .Z(c[457]) );
  XNOR U2296 ( .A(b[458]), .B(a[458]), .Z(n1838) );
  OR U2297 ( .A(b[457]), .B(a[457]), .Z(n1836) );
  OR U2298 ( .A(n1834), .B(n1833), .Z(n1835) );
  AND U2299 ( .A(n1836), .B(n1835), .Z(n1837) );
  XNOR U2300 ( .A(n1838), .B(n1837), .Z(c[458]) );
  XNOR U2301 ( .A(b[459]), .B(a[459]), .Z(n1842) );
  OR U2302 ( .A(b[458]), .B(a[458]), .Z(n1840) );
  OR U2303 ( .A(n1838), .B(n1837), .Z(n1839) );
  AND U2304 ( .A(n1840), .B(n1839), .Z(n1841) );
  XNOR U2305 ( .A(n1842), .B(n1841), .Z(c[459]) );
  XNOR U2306 ( .A(b[460]), .B(a[460]), .Z(n1846) );
  OR U2307 ( .A(b[459]), .B(a[459]), .Z(n1844) );
  OR U2308 ( .A(n1842), .B(n1841), .Z(n1843) );
  AND U2309 ( .A(n1844), .B(n1843), .Z(n1845) );
  XNOR U2310 ( .A(n1846), .B(n1845), .Z(c[460]) );
  XNOR U2311 ( .A(b[461]), .B(a[461]), .Z(n1850) );
  OR U2312 ( .A(b[460]), .B(a[460]), .Z(n1848) );
  OR U2313 ( .A(n1846), .B(n1845), .Z(n1847) );
  AND U2314 ( .A(n1848), .B(n1847), .Z(n1849) );
  XNOR U2315 ( .A(n1850), .B(n1849), .Z(c[461]) );
  XNOR U2316 ( .A(b[462]), .B(a[462]), .Z(n1854) );
  OR U2317 ( .A(b[461]), .B(a[461]), .Z(n1852) );
  OR U2318 ( .A(n1850), .B(n1849), .Z(n1851) );
  AND U2319 ( .A(n1852), .B(n1851), .Z(n1853) );
  XNOR U2320 ( .A(n1854), .B(n1853), .Z(c[462]) );
  XNOR U2321 ( .A(b[463]), .B(a[463]), .Z(n1858) );
  OR U2322 ( .A(b[462]), .B(a[462]), .Z(n1856) );
  OR U2323 ( .A(n1854), .B(n1853), .Z(n1855) );
  AND U2324 ( .A(n1856), .B(n1855), .Z(n1857) );
  XNOR U2325 ( .A(n1858), .B(n1857), .Z(c[463]) );
  OR U2326 ( .A(b[463]), .B(a[463]), .Z(n1860) );
  OR U2327 ( .A(n1858), .B(n1857), .Z(n1859) );
  NAND U2328 ( .A(n1860), .B(n1859), .Z(n1862) );
  XOR U2329 ( .A(a[464]), .B(b[464]), .Z(n1861) );
  XNOR U2330 ( .A(n1862), .B(n1861), .Z(c[464]) );
  XOR U2331 ( .A(a[465]), .B(b[465]), .Z(n1865) );
  NAND U2332 ( .A(b[464]), .B(a[464]), .Z(n1864) );
  NANDN U2333 ( .A(n1862), .B(n1861), .Z(n1863) );
  AND U2334 ( .A(n1864), .B(n1863), .Z(n1866) );
  XNOR U2335 ( .A(n1865), .B(n1866), .Z(c[465]) );
  XOR U2336 ( .A(a[466]), .B(b[466]), .Z(n1869) );
  NAND U2337 ( .A(b[465]), .B(a[465]), .Z(n1868) );
  NANDN U2338 ( .A(n1866), .B(n1865), .Z(n1867) );
  AND U2339 ( .A(n1868), .B(n1867), .Z(n1870) );
  XNOR U2340 ( .A(n1869), .B(n1870), .Z(c[466]) );
  XOR U2341 ( .A(a[467]), .B(b[467]), .Z(n1873) );
  NAND U2342 ( .A(b[466]), .B(a[466]), .Z(n1872) );
  NANDN U2343 ( .A(n1870), .B(n1869), .Z(n1871) );
  AND U2344 ( .A(n1872), .B(n1871), .Z(n1874) );
  XNOR U2345 ( .A(n1873), .B(n1874), .Z(c[467]) );
  XOR U2346 ( .A(a[468]), .B(b[468]), .Z(n1877) );
  NAND U2347 ( .A(b[467]), .B(a[467]), .Z(n1876) );
  NANDN U2348 ( .A(n1874), .B(n1873), .Z(n1875) );
  AND U2349 ( .A(n1876), .B(n1875), .Z(n1878) );
  XNOR U2350 ( .A(n1877), .B(n1878), .Z(c[468]) );
  XOR U2351 ( .A(a[469]), .B(b[469]), .Z(n1881) );
  NAND U2352 ( .A(b[468]), .B(a[468]), .Z(n1880) );
  NANDN U2353 ( .A(n1878), .B(n1877), .Z(n1879) );
  AND U2354 ( .A(n1880), .B(n1879), .Z(n1882) );
  XNOR U2355 ( .A(n1881), .B(n1882), .Z(c[469]) );
  XOR U2356 ( .A(a[470]), .B(b[470]), .Z(n1885) );
  NAND U2357 ( .A(b[469]), .B(a[469]), .Z(n1884) );
  NANDN U2358 ( .A(n1882), .B(n1881), .Z(n1883) );
  AND U2359 ( .A(n1884), .B(n1883), .Z(n1886) );
  XNOR U2360 ( .A(n1885), .B(n1886), .Z(c[470]) );
  XOR U2361 ( .A(a[471]), .B(b[471]), .Z(n1889) );
  NAND U2362 ( .A(b[470]), .B(a[470]), .Z(n1888) );
  NANDN U2363 ( .A(n1886), .B(n1885), .Z(n1887) );
  AND U2364 ( .A(n1888), .B(n1887), .Z(n1890) );
  XNOR U2365 ( .A(n1889), .B(n1890), .Z(c[471]) );
  XOR U2366 ( .A(a[472]), .B(b[472]), .Z(n1893) );
  NAND U2367 ( .A(b[471]), .B(a[471]), .Z(n1892) );
  NANDN U2368 ( .A(n1890), .B(n1889), .Z(n1891) );
  AND U2369 ( .A(n1892), .B(n1891), .Z(n1894) );
  XNOR U2370 ( .A(n1893), .B(n1894), .Z(c[472]) );
  XOR U2371 ( .A(a[473]), .B(b[473]), .Z(n1897) );
  NAND U2372 ( .A(b[472]), .B(a[472]), .Z(n1896) );
  NANDN U2373 ( .A(n1894), .B(n1893), .Z(n1895) );
  AND U2374 ( .A(n1896), .B(n1895), .Z(n1898) );
  XNOR U2375 ( .A(n1897), .B(n1898), .Z(c[473]) );
  XOR U2376 ( .A(a[474]), .B(b[474]), .Z(n1901) );
  NAND U2377 ( .A(b[473]), .B(a[473]), .Z(n1900) );
  NANDN U2378 ( .A(n1898), .B(n1897), .Z(n1899) );
  AND U2379 ( .A(n1900), .B(n1899), .Z(n1902) );
  XNOR U2380 ( .A(n1901), .B(n1902), .Z(c[474]) );
  XOR U2381 ( .A(a[475]), .B(b[475]), .Z(n1905) );
  NAND U2382 ( .A(b[474]), .B(a[474]), .Z(n1904) );
  NANDN U2383 ( .A(n1902), .B(n1901), .Z(n1903) );
  AND U2384 ( .A(n1904), .B(n1903), .Z(n1906) );
  XNOR U2385 ( .A(n1905), .B(n1906), .Z(c[475]) );
  XOR U2386 ( .A(a[476]), .B(b[476]), .Z(n1909) );
  NAND U2387 ( .A(b[475]), .B(a[475]), .Z(n1908) );
  NANDN U2388 ( .A(n1906), .B(n1905), .Z(n1907) );
  AND U2389 ( .A(n1908), .B(n1907), .Z(n1910) );
  XNOR U2390 ( .A(n1909), .B(n1910), .Z(c[476]) );
  XOR U2391 ( .A(a[477]), .B(b[477]), .Z(n1913) );
  NAND U2392 ( .A(b[476]), .B(a[476]), .Z(n1912) );
  NANDN U2393 ( .A(n1910), .B(n1909), .Z(n1911) );
  AND U2394 ( .A(n1912), .B(n1911), .Z(n1914) );
  XNOR U2395 ( .A(n1913), .B(n1914), .Z(c[477]) );
  XOR U2396 ( .A(a[478]), .B(b[478]), .Z(n1917) );
  NAND U2397 ( .A(b[477]), .B(a[477]), .Z(n1916) );
  NANDN U2398 ( .A(n1914), .B(n1913), .Z(n1915) );
  AND U2399 ( .A(n1916), .B(n1915), .Z(n1918) );
  XNOR U2400 ( .A(n1917), .B(n1918), .Z(c[478]) );
  XOR U2401 ( .A(a[479]), .B(b[479]), .Z(n1921) );
  NAND U2402 ( .A(b[478]), .B(a[478]), .Z(n1920) );
  NANDN U2403 ( .A(n1918), .B(n1917), .Z(n1919) );
  AND U2404 ( .A(n1920), .B(n1919), .Z(n1922) );
  XNOR U2405 ( .A(n1921), .B(n1922), .Z(c[479]) );
  XOR U2406 ( .A(a[480]), .B(b[480]), .Z(n1925) );
  NAND U2407 ( .A(b[479]), .B(a[479]), .Z(n1924) );
  NANDN U2408 ( .A(n1922), .B(n1921), .Z(n1923) );
  AND U2409 ( .A(n1924), .B(n1923), .Z(n1926) );
  XNOR U2410 ( .A(n1925), .B(n1926), .Z(c[480]) );
  XOR U2411 ( .A(a[481]), .B(b[481]), .Z(n1929) );
  NAND U2412 ( .A(b[480]), .B(a[480]), .Z(n1928) );
  NANDN U2413 ( .A(n1926), .B(n1925), .Z(n1927) );
  AND U2414 ( .A(n1928), .B(n1927), .Z(n1930) );
  XNOR U2415 ( .A(n1929), .B(n1930), .Z(c[481]) );
  XOR U2416 ( .A(a[482]), .B(b[482]), .Z(n1933) );
  NAND U2417 ( .A(b[481]), .B(a[481]), .Z(n1932) );
  NANDN U2418 ( .A(n1930), .B(n1929), .Z(n1931) );
  AND U2419 ( .A(n1932), .B(n1931), .Z(n1934) );
  XNOR U2420 ( .A(n1933), .B(n1934), .Z(c[482]) );
  XOR U2421 ( .A(a[483]), .B(b[483]), .Z(n1937) );
  NAND U2422 ( .A(b[482]), .B(a[482]), .Z(n1936) );
  NANDN U2423 ( .A(n1934), .B(n1933), .Z(n1935) );
  AND U2424 ( .A(n1936), .B(n1935), .Z(n1938) );
  XNOR U2425 ( .A(n1937), .B(n1938), .Z(c[483]) );
  XOR U2426 ( .A(a[484]), .B(b[484]), .Z(n1941) );
  NAND U2427 ( .A(b[483]), .B(a[483]), .Z(n1940) );
  NANDN U2428 ( .A(n1938), .B(n1937), .Z(n1939) );
  AND U2429 ( .A(n1940), .B(n1939), .Z(n1942) );
  XNOR U2430 ( .A(n1941), .B(n1942), .Z(c[484]) );
  XOR U2431 ( .A(a[485]), .B(b[485]), .Z(n1945) );
  NAND U2432 ( .A(b[484]), .B(a[484]), .Z(n1944) );
  NANDN U2433 ( .A(n1942), .B(n1941), .Z(n1943) );
  AND U2434 ( .A(n1944), .B(n1943), .Z(n1946) );
  XNOR U2435 ( .A(n1945), .B(n1946), .Z(c[485]) );
  XOR U2436 ( .A(a[486]), .B(b[486]), .Z(n1949) );
  NAND U2437 ( .A(b[485]), .B(a[485]), .Z(n1948) );
  NANDN U2438 ( .A(n1946), .B(n1945), .Z(n1947) );
  AND U2439 ( .A(n1948), .B(n1947), .Z(n1950) );
  XNOR U2440 ( .A(n1949), .B(n1950), .Z(c[486]) );
  XOR U2441 ( .A(a[487]), .B(b[487]), .Z(n1953) );
  NAND U2442 ( .A(b[486]), .B(a[486]), .Z(n1952) );
  NANDN U2443 ( .A(n1950), .B(n1949), .Z(n1951) );
  AND U2444 ( .A(n1952), .B(n1951), .Z(n1954) );
  XNOR U2445 ( .A(n1953), .B(n1954), .Z(c[487]) );
  XOR U2446 ( .A(a[488]), .B(b[488]), .Z(n1957) );
  NAND U2447 ( .A(b[487]), .B(a[487]), .Z(n1956) );
  NANDN U2448 ( .A(n1954), .B(n1953), .Z(n1955) );
  AND U2449 ( .A(n1956), .B(n1955), .Z(n1958) );
  XNOR U2450 ( .A(n1957), .B(n1958), .Z(c[488]) );
  XOR U2451 ( .A(a[489]), .B(b[489]), .Z(n1961) );
  NAND U2452 ( .A(b[488]), .B(a[488]), .Z(n1960) );
  NANDN U2453 ( .A(n1958), .B(n1957), .Z(n1959) );
  AND U2454 ( .A(n1960), .B(n1959), .Z(n1962) );
  XNOR U2455 ( .A(n1961), .B(n1962), .Z(c[489]) );
  XOR U2456 ( .A(a[490]), .B(b[490]), .Z(n1965) );
  NAND U2457 ( .A(b[489]), .B(a[489]), .Z(n1964) );
  NANDN U2458 ( .A(n1962), .B(n1961), .Z(n1963) );
  AND U2459 ( .A(n1964), .B(n1963), .Z(n1966) );
  XNOR U2460 ( .A(n1965), .B(n1966), .Z(c[490]) );
  XOR U2461 ( .A(a[491]), .B(b[491]), .Z(n1969) );
  NAND U2462 ( .A(b[490]), .B(a[490]), .Z(n1968) );
  NANDN U2463 ( .A(n1966), .B(n1965), .Z(n1967) );
  AND U2464 ( .A(n1968), .B(n1967), .Z(n1970) );
  XNOR U2465 ( .A(n1969), .B(n1970), .Z(c[491]) );
  XOR U2466 ( .A(a[492]), .B(b[492]), .Z(n1973) );
  NAND U2467 ( .A(b[491]), .B(a[491]), .Z(n1972) );
  NANDN U2468 ( .A(n1970), .B(n1969), .Z(n1971) );
  AND U2469 ( .A(n1972), .B(n1971), .Z(n1974) );
  XNOR U2470 ( .A(n1973), .B(n1974), .Z(c[492]) );
  NAND U2471 ( .A(b[492]), .B(a[492]), .Z(n1976) );
  NANDN U2472 ( .A(n1974), .B(n1973), .Z(n1975) );
  NAND U2473 ( .A(n1976), .B(n1975), .Z(n1978) );
  XNOR U2474 ( .A(b[493]), .B(a[493]), .Z(n1977) );
  XNOR U2475 ( .A(n1978), .B(n1977), .Z(c[493]) );
  XOR U2476 ( .A(a[494]), .B(b[494]), .Z(n1981) );
  OR U2477 ( .A(b[493]), .B(a[493]), .Z(n1980) );
  OR U2478 ( .A(n1978), .B(n1977), .Z(n1979) );
  NAND U2479 ( .A(n1980), .B(n1979), .Z(n1982) );
  XNOR U2480 ( .A(n1981), .B(n1982), .Z(c[494]) );
  XOR U2481 ( .A(a[495]), .B(b[495]), .Z(n1985) );
  NAND U2482 ( .A(b[494]), .B(a[494]), .Z(n1984) );
  NANDN U2483 ( .A(n1982), .B(n1981), .Z(n1983) );
  AND U2484 ( .A(n1984), .B(n1983), .Z(n1986) );
  XNOR U2485 ( .A(n1985), .B(n1986), .Z(c[495]) );
  NAND U2486 ( .A(b[495]), .B(a[495]), .Z(n1988) );
  NANDN U2487 ( .A(n1986), .B(n1985), .Z(n1987) );
  NAND U2488 ( .A(n1988), .B(n1987), .Z(n1990) );
  XNOR U2489 ( .A(b[496]), .B(a[496]), .Z(n1989) );
  XNOR U2490 ( .A(n1990), .B(n1989), .Z(c[496]) );
  XOR U2491 ( .A(a[497]), .B(b[497]), .Z(n1993) );
  OR U2492 ( .A(b[496]), .B(a[496]), .Z(n1992) );
  OR U2493 ( .A(n1990), .B(n1989), .Z(n1991) );
  NAND U2494 ( .A(n1992), .B(n1991), .Z(n1994) );
  XNOR U2495 ( .A(n1993), .B(n1994), .Z(c[497]) );
  NAND U2496 ( .A(b[497]), .B(a[497]), .Z(n1996) );
  NANDN U2497 ( .A(n1994), .B(n1993), .Z(n1995) );
  NAND U2498 ( .A(n1996), .B(n1995), .Z(n1998) );
  XNOR U2499 ( .A(b[498]), .B(a[498]), .Z(n1997) );
  XNOR U2500 ( .A(n1998), .B(n1997), .Z(c[498]) );
  XNOR U2501 ( .A(b[499]), .B(a[499]), .Z(n2002) );
  OR U2502 ( .A(b[498]), .B(a[498]), .Z(n2000) );
  OR U2503 ( .A(n1998), .B(n1997), .Z(n1999) );
  AND U2504 ( .A(n2000), .B(n1999), .Z(n2001) );
  XNOR U2505 ( .A(n2002), .B(n2001), .Z(c[499]) );
  XOR U2506 ( .A(a[500]), .B(b[500]), .Z(n2005) );
  OR U2507 ( .A(b[499]), .B(a[499]), .Z(n2004) );
  OR U2508 ( .A(n2002), .B(n2001), .Z(n2003) );
  NAND U2509 ( .A(n2004), .B(n2003), .Z(n2006) );
  XNOR U2510 ( .A(n2005), .B(n2006), .Z(c[500]) );
  NAND U2511 ( .A(b[500]), .B(a[500]), .Z(n2008) );
  NANDN U2512 ( .A(n2006), .B(n2005), .Z(n2007) );
  NAND U2513 ( .A(n2008), .B(n2007), .Z(n2010) );
  XNOR U2514 ( .A(b[501]), .B(a[501]), .Z(n2009) );
  XNOR U2515 ( .A(n2010), .B(n2009), .Z(c[501]) );
  XNOR U2516 ( .A(b[502]), .B(a[502]), .Z(n2014) );
  OR U2517 ( .A(b[501]), .B(a[501]), .Z(n2012) );
  OR U2518 ( .A(n2010), .B(n2009), .Z(n2011) );
  AND U2519 ( .A(n2012), .B(n2011), .Z(n2013) );
  XNOR U2520 ( .A(n2014), .B(n2013), .Z(c[502]) );
  XNOR U2521 ( .A(b[503]), .B(a[503]), .Z(n2018) );
  OR U2522 ( .A(b[502]), .B(a[502]), .Z(n2016) );
  OR U2523 ( .A(n2014), .B(n2013), .Z(n2015) );
  AND U2524 ( .A(n2016), .B(n2015), .Z(n2017) );
  XNOR U2525 ( .A(n2018), .B(n2017), .Z(c[503]) );
  XNOR U2526 ( .A(b[504]), .B(a[504]), .Z(n2022) );
  OR U2527 ( .A(b[503]), .B(a[503]), .Z(n2020) );
  OR U2528 ( .A(n2018), .B(n2017), .Z(n2019) );
  AND U2529 ( .A(n2020), .B(n2019), .Z(n2021) );
  XNOR U2530 ( .A(n2022), .B(n2021), .Z(c[504]) );
  XNOR U2531 ( .A(b[505]), .B(a[505]), .Z(n2026) );
  OR U2532 ( .A(b[504]), .B(a[504]), .Z(n2024) );
  OR U2533 ( .A(n2022), .B(n2021), .Z(n2023) );
  AND U2534 ( .A(n2024), .B(n2023), .Z(n2025) );
  XNOR U2535 ( .A(n2026), .B(n2025), .Z(c[505]) );
  XNOR U2536 ( .A(b[506]), .B(a[506]), .Z(n2030) );
  OR U2537 ( .A(b[505]), .B(a[505]), .Z(n2028) );
  OR U2538 ( .A(n2026), .B(n2025), .Z(n2027) );
  AND U2539 ( .A(n2028), .B(n2027), .Z(n2029) );
  XNOR U2540 ( .A(n2030), .B(n2029), .Z(c[506]) );
  XNOR U2541 ( .A(b[507]), .B(a[507]), .Z(n2034) );
  OR U2542 ( .A(b[506]), .B(a[506]), .Z(n2032) );
  OR U2543 ( .A(n2030), .B(n2029), .Z(n2031) );
  AND U2544 ( .A(n2032), .B(n2031), .Z(n2033) );
  XNOR U2545 ( .A(n2034), .B(n2033), .Z(c[507]) );
  XNOR U2546 ( .A(b[508]), .B(a[508]), .Z(n2038) );
  OR U2547 ( .A(b[507]), .B(a[507]), .Z(n2036) );
  OR U2548 ( .A(n2034), .B(n2033), .Z(n2035) );
  AND U2549 ( .A(n2036), .B(n2035), .Z(n2037) );
  XNOR U2550 ( .A(n2038), .B(n2037), .Z(c[508]) );
  XNOR U2551 ( .A(b[509]), .B(a[509]), .Z(n2042) );
  OR U2552 ( .A(b[508]), .B(a[508]), .Z(n2040) );
  OR U2553 ( .A(n2038), .B(n2037), .Z(n2039) );
  AND U2554 ( .A(n2040), .B(n2039), .Z(n2041) );
  XNOR U2555 ( .A(n2042), .B(n2041), .Z(c[509]) );
  XNOR U2556 ( .A(b[510]), .B(a[510]), .Z(n2046) );
  OR U2557 ( .A(b[509]), .B(a[509]), .Z(n2044) );
  OR U2558 ( .A(n2042), .B(n2041), .Z(n2043) );
  AND U2559 ( .A(n2044), .B(n2043), .Z(n2045) );
  XNOR U2560 ( .A(n2046), .B(n2045), .Z(c[510]) );
  OR U2561 ( .A(b[510]), .B(a[510]), .Z(n2048) );
  OR U2562 ( .A(n2046), .B(n2045), .Z(n2047) );
  AND U2563 ( .A(n2048), .B(n2047), .Z(n2050) );
  XOR U2564 ( .A(a[511]), .B(b[511]), .Z(n2049) );
  XOR U2565 ( .A(n2050), .B(n2049), .Z(c[511]) );
endmodule

