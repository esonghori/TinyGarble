
module compare_N16384_CC8 ( clk, rst, x, y, g, e );
  input [2047:0] x;
  input [2047:0] y;
  input clk, rst;
  output g, e;
  wire   ebreg, n4, n5, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
         n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
         n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
         n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
         n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303,
         n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
         n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323,
         n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333,
         n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343,
         n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353,
         n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363,
         n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373,
         n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383,
         n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393,
         n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
         n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
         n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423,
         n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433,
         n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443,
         n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453,
         n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463,
         n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
         n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
         n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493,
         n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503,
         n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513,
         n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523,
         n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533,
         n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543,
         n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553,
         n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563,
         n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
         n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583,
         n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
         n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603,
         n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
         n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
         n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
         n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
         n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
         n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
         n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
         n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
         n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
         n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
         n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743,
         n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753,
         n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763,
         n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773,
         n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783,
         n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793,
         n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
         n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
         n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
         n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
         n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843,
         n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853,
         n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863,
         n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873,
         n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883,
         n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893,
         n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903,
         n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913,
         n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923,
         n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933,
         n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943,
         n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
         n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963,
         n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973,
         n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
         n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
         n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
         n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
         n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
         n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
         n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
         n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
         n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063,
         n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
         n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
         n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
         n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
         n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
         n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
         n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
         n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
         n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
         n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
         n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
         n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
         n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
         n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
         n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
         n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
         n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
         n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
         n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
         n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
         n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
         n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
         n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
         n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
         n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
         n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
         n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
         n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
         n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
         n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
         n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
         n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
         n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
         n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,
         n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
         n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,
         n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,
         n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
         n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
         n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
         n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,
         n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,
         n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,
         n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770,
         n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778,
         n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786,
         n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,
         n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802,
         n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
         n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,
         n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
         n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834,
         n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842,
         n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,
         n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858,
         n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866,
         n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874,
         n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
         n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890,
         n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
         n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906,
         n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,
         n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922,
         n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
         n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938,
         n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946,
         n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954,
         n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,
         n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
         n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
         n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986,
         n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,
         n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
         n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010,
         n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
         n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026,
         n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034,
         n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
         n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
         n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,
         n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
         n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
         n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
         n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
         n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
         n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
         n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122,
         n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130,
         n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138,
         n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146,
         n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154,
         n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162,
         n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,
         n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178,
         n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
         n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
         n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
         n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,
         n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
         n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
         n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
         n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
         n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,
         n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
         n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
         n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
         n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
         n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
         n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
         n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
         n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
         n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
         n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
         n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
         n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
         n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
         n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
         n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
         n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
         n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,
         n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
         n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
         n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,
         n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
         n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
         n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
         n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
         n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
         n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
         n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
         n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
         n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
         n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
         n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
         n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898,
         n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
         n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
         n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
         n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
         n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
         n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
         n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
         n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
         n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970,
         n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
         n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986,
         n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
         n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
         n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
         n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
         n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
         n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
         n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
         n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
         n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162,
         n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
         n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
         n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186,
         n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
         n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
         n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
         n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,
         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,
         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
         n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
         n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
         n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
         n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
         n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,
         n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,
         n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,
         n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522,
         n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
         n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,
         n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546,
         n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
         n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
         n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570,
         n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578,
         n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586,
         n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594,
         n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602,
         n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,
         n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618,
         n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
         n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634,
         n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642,
         n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650,
         n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658,
         n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666,
         n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674,
         n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682,
         n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690,
         n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
         n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,
         n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714,
         n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722,
         n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,
         n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738,
         n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746,
         n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
         n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762,
         n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
         n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,
         n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786,
         n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794,
         n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
         n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,
         n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
         n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,
         n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834,
         n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
         n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850,
         n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858,
         n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,
         n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
         n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882,
         n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890,
         n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
         n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
         n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
         n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
         n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930,
         n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,
         n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,
         n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954,
         n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,
         n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
         n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,
         n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
         n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
         n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
         n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,
         n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
         n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
         n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
         n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042,
         n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
         n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
         n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
         n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074,
         n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082,
         n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,
         n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
         n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
         n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,
         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
         n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,
         n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
         n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234,
         n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
         n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,
         n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
         n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
         n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
         n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079;

  DFF ebreg_reg ( .D(n5), .CLK(clk), .RST(rst), .Q(ebreg) );
  DFF greg_reg ( .D(n4), .CLK(clk), .RST(rst), .Q(g) );
  NANDN U10 ( .A(x[475]), .B(y[475]), .Z(n8) );
  NANDN U11 ( .A(x[476]), .B(y[476]), .Z(n9) );
  NANDN U12 ( .A(x[477]), .B(y[477]), .Z(n10) );
  NAND U13 ( .A(n9), .B(n10), .Z(n11) );
  ANDN U14 ( .B(n8), .A(n11), .Z(n12) );
  NANDN U15 ( .A(x[474]), .B(y[474]), .Z(n13) );
  XNOR U16 ( .A(y[475]), .B(x[475]), .Z(n14) );
  NANDN U17 ( .A(n13), .B(n14), .Z(n15) );
  NAND U18 ( .A(n12), .B(n15), .Z(n10826) );
  NANDN U19 ( .A(y[563]), .B(x[563]), .Z(n16) );
  NANDN U20 ( .A(y[564]), .B(x[564]), .Z(n17) );
  NANDN U21 ( .A(y[565]), .B(x[565]), .Z(n18) );
  NAND U22 ( .A(n17), .B(n18), .Z(n19) );
  ANDN U23 ( .B(n16), .A(n19), .Z(n20) );
  NANDN U24 ( .A(y[562]), .B(x[562]), .Z(n21) );
  XNOR U25 ( .A(x[563]), .B(y[563]), .Z(n22) );
  NANDN U26 ( .A(n21), .B(n22), .Z(n23) );
  NAND U27 ( .A(n20), .B(n23), .Z(n10965) );
  NANDN U28 ( .A(y[620]), .B(x[620]), .Z(n24) );
  NANDN U29 ( .A(n6514), .B(n24), .Z(n11068) );
  NANDN U30 ( .A(y[685]), .B(x[685]), .Z(n25) );
  XNOR U31 ( .A(y[685]), .B(x[685]), .Z(n26) );
  NANDN U32 ( .A(x[684]), .B(y[684]), .Z(n27) );
  NAND U33 ( .A(n26), .B(n27), .Z(n28) );
  NAND U34 ( .A(n25), .B(n28), .Z(n11135) );
  NANDN U35 ( .A(y[1096]), .B(x[1096]), .Z(n29) );
  AND U36 ( .A(n4132), .B(n29), .Z(n30) );
  ANDN U37 ( .B(x[1094]), .A(y[1094]), .Z(n31) );
  NAND U38 ( .A(n31), .B(x[1095]), .Z(n32) );
  AND U39 ( .A(n30), .B(n32), .Z(n33) );
  XOR U40 ( .A(x[1095]), .B(n31), .Z(n34) );
  NANDN U41 ( .A(y[1095]), .B(n34), .Z(n35) );
  NAND U42 ( .A(n33), .B(n35), .Z(n12053) );
  NANDN U43 ( .A(y[196]), .B(x[196]), .Z(n36) );
  AND U44 ( .A(n6565), .B(n36), .Z(n10352) );
  NANDN U45 ( .A(x[350]), .B(y[350]), .Z(n37) );
  NAND U46 ( .A(n37), .B(n2677), .Z(n10632) );
  NANDN U47 ( .A(x[386]), .B(y[386]), .Z(n38) );
  AND U48 ( .A(n2766), .B(n38), .Z(n10683) );
  NANDN U49 ( .A(x[456]), .B(y[456]), .Z(n39) );
  NAND U50 ( .A(n39), .B(n2894), .Z(n10800) );
  NANDN U51 ( .A(x[489]), .B(y[489]), .Z(n40) );
  XNOR U52 ( .A(x[489]), .B(y[489]), .Z(n41) );
  NANDN U53 ( .A(y[488]), .B(x[488]), .Z(n42) );
  NAND U54 ( .A(n41), .B(n42), .Z(n43) );
  NAND U55 ( .A(n40), .B(n43), .Z(n10847) );
  NANDN U56 ( .A(y[527]), .B(x[527]), .Z(n44) );
  NANDN U57 ( .A(y[528]), .B(x[528]), .Z(n45) );
  NANDN U58 ( .A(y[529]), .B(x[529]), .Z(n46) );
  NAND U59 ( .A(n45), .B(n46), .Z(n47) );
  ANDN U60 ( .B(n44), .A(n47), .Z(n48) );
  NANDN U61 ( .A(y[526]), .B(x[526]), .Z(n49) );
  XNOR U62 ( .A(x[527]), .B(y[527]), .Z(n50) );
  NANDN U63 ( .A(n49), .B(n50), .Z(n51) );
  NAND U64 ( .A(n48), .B(n51), .Z(n10924) );
  NANDN U65 ( .A(x[575]), .B(y[575]), .Z(n52) );
  NANDN U66 ( .A(x[576]), .B(y[576]), .Z(n53) );
  NANDN U67 ( .A(x[577]), .B(y[577]), .Z(n54) );
  NAND U68 ( .A(n53), .B(n54), .Z(n55) );
  ANDN U69 ( .B(n52), .A(n55), .Z(n56) );
  NANDN U70 ( .A(x[574]), .B(y[574]), .Z(n57) );
  XNOR U71 ( .A(y[575]), .B(x[575]), .Z(n58) );
  NANDN U72 ( .A(n57), .B(n58), .Z(n59) );
  NAND U73 ( .A(n56), .B(n59), .Z(n10983) );
  ANDN U74 ( .B(x[622]), .A(y[622]), .Z(n60) );
  NANDN U75 ( .A(y[625]), .B(x[625]), .Z(n61) );
  NANDN U76 ( .A(y[624]), .B(x[624]), .Z(n62) );
  AND U77 ( .A(n61), .B(n62), .Z(n63) );
  OR U78 ( .A(x[623]), .B(n60), .Z(n64) );
  XOR U79 ( .A(x[623]), .B(n60), .Z(n65) );
  NAND U80 ( .A(n65), .B(y[623]), .Z(n66) );
  NAND U81 ( .A(n64), .B(n66), .Z(n67) );
  AND U82 ( .A(n63), .B(n67), .Z(n11071) );
  NANDN U83 ( .A(x[653]), .B(y[653]), .Z(n68) );
  NANDN U84 ( .A(x[654]), .B(y[654]), .Z(n69) );
  NANDN U85 ( .A(x[655]), .B(y[655]), .Z(n70) );
  NAND U86 ( .A(n69), .B(n70), .Z(n71) );
  ANDN U87 ( .B(n68), .A(n71), .Z(n72) );
  NANDN U88 ( .A(x[652]), .B(y[652]), .Z(n73) );
  XNOR U89 ( .A(y[653]), .B(x[653]), .Z(n74) );
  NANDN U90 ( .A(n73), .B(n74), .Z(n75) );
  NAND U91 ( .A(n72), .B(n75), .Z(n11101) );
  NANDN U92 ( .A(x[672]), .B(y[672]), .Z(n76) );
  AND U93 ( .A(n3286), .B(n76), .Z(n11122) );
  NANDN U94 ( .A(y[1091]), .B(x[1091]), .Z(n77) );
  ANDN U95 ( .B(n77), .A(n8078), .Z(n12046) );
  NANDN U96 ( .A(x[1240]), .B(y[1240]), .Z(n78) );
  NAND U97 ( .A(n78), .B(n4459), .Z(n12350) );
  NANDN U98 ( .A(x[134]), .B(y[134]), .Z(n79) );
  AND U99 ( .A(n2278), .B(n79), .Z(n10252) );
  NANDN U100 ( .A(x[204]), .B(y[204]), .Z(n80) );
  NAND U101 ( .A(n80), .B(n2415), .Z(n10377) );
  NANDN U102 ( .A(y[237]), .B(x[237]), .Z(n81) );
  NANDN U103 ( .A(y[238]), .B(x[238]), .Z(n82) );
  NANDN U104 ( .A(y[239]), .B(x[239]), .Z(n83) );
  NAND U105 ( .A(n82), .B(n83), .Z(n84) );
  ANDN U106 ( .B(n81), .A(n84), .Z(n85) );
  NANDN U107 ( .A(y[236]), .B(x[236]), .Z(n86) );
  XNOR U108 ( .A(x[237]), .B(y[237]), .Z(n87) );
  NANDN U109 ( .A(n86), .B(n87), .Z(n88) );
  NAND U110 ( .A(n85), .B(n88), .Z(n10411) );
  NANDN U111 ( .A(y[319]), .B(x[319]), .Z(n89) );
  XNOR U112 ( .A(y[319]), .B(x[319]), .Z(n90) );
  NANDN U113 ( .A(x[318]), .B(y[318]), .Z(n91) );
  NAND U114 ( .A(n90), .B(n91), .Z(n92) );
  NAND U115 ( .A(n89), .B(n92), .Z(n10571) );
  NANDN U116 ( .A(y[355]), .B(x[355]), .Z(n93) );
  NANDN U117 ( .A(y[356]), .B(x[356]), .Z(n94) );
  NANDN U118 ( .A(y[357]), .B(x[357]), .Z(n95) );
  NAND U119 ( .A(n94), .B(n95), .Z(n96) );
  ANDN U120 ( .B(n93), .A(n96), .Z(n97) );
  NANDN U121 ( .A(y[354]), .B(x[354]), .Z(n98) );
  XNOR U122 ( .A(x[355]), .B(y[355]), .Z(n99) );
  NANDN U123 ( .A(n98), .B(n99), .Z(n100) );
  NAND U124 ( .A(n97), .B(n100), .Z(n10639) );
  NANDN U125 ( .A(x[401]), .B(y[401]), .Z(n101) );
  NANDN U126 ( .A(x[402]), .B(y[402]), .Z(n102) );
  NANDN U127 ( .A(x[403]), .B(y[403]), .Z(n103) );
  NAND U128 ( .A(n102), .B(n103), .Z(n104) );
  ANDN U129 ( .B(n101), .A(n104), .Z(n105) );
  NANDN U130 ( .A(x[400]), .B(y[400]), .Z(n106) );
  XNOR U131 ( .A(y[401]), .B(x[401]), .Z(n107) );
  NANDN U132 ( .A(n106), .B(n107), .Z(n108) );
  NAND U133 ( .A(n105), .B(n108), .Z(n10709) );
  NANDN U134 ( .A(y[462]), .B(x[462]), .Z(n109) );
  AND U135 ( .A(n1542), .B(n109), .Z(n110) );
  ANDN U136 ( .B(x[460]), .A(y[460]), .Z(n111) );
  NAND U137 ( .A(n111), .B(x[461]), .Z(n112) );
  AND U138 ( .A(n110), .B(n112), .Z(n113) );
  XOR U139 ( .A(x[461]), .B(n111), .Z(n114) );
  NANDN U140 ( .A(y[461]), .B(n114), .Z(n115) );
  NAND U141 ( .A(n113), .B(n115), .Z(n10807) );
  NANDN U142 ( .A(x[493]), .B(y[493]), .Z(n116) );
  NANDN U143 ( .A(x[494]), .B(y[494]), .Z(n117) );
  NANDN U144 ( .A(x[495]), .B(y[495]), .Z(n118) );
  NAND U145 ( .A(n117), .B(n118), .Z(n119) );
  ANDN U146 ( .B(n116), .A(n119), .Z(n120) );
  NANDN U147 ( .A(x[492]), .B(y[492]), .Z(n121) );
  XNOR U148 ( .A(y[493]), .B(x[493]), .Z(n122) );
  NANDN U149 ( .A(n121), .B(n122), .Z(n123) );
  NAND U150 ( .A(n120), .B(n123), .Z(n10853) );
  NANDN U151 ( .A(x[531]), .B(y[531]), .Z(n124) );
  XNOR U152 ( .A(x[531]), .B(y[531]), .Z(n125) );
  NANDN U153 ( .A(y[530]), .B(x[530]), .Z(n126) );
  NAND U154 ( .A(n125), .B(n126), .Z(n127) );
  NAND U155 ( .A(n124), .B(n127), .Z(n10927) );
  NANDN U156 ( .A(y[565]), .B(x[565]), .Z(n128) );
  XNOR U157 ( .A(y[565]), .B(x[565]), .Z(n129) );
  NANDN U158 ( .A(x[564]), .B(y[564]), .Z(n130) );
  NAND U159 ( .A(n129), .B(n130), .Z(n131) );
  NAND U160 ( .A(n128), .B(n131), .Z(n10966) );
  NANDN U161 ( .A(x[582]), .B(y[582]), .Z(n132) );
  AND U162 ( .A(n3104), .B(n132), .Z(n10999) );
  NANDN U163 ( .A(x[592]), .B(y[592]), .Z(n133) );
  NAND U164 ( .A(n133), .B(n3123), .Z(n11026) );
  NANDN U165 ( .A(x[627]), .B(y[627]), .Z(n134) );
  XNOR U166 ( .A(x[627]), .B(y[627]), .Z(n135) );
  NANDN U167 ( .A(y[626]), .B(x[626]), .Z(n136) );
  NAND U168 ( .A(n135), .B(n136), .Z(n137) );
  NAND U169 ( .A(n134), .B(n137), .Z(n11075) );
  NANDN U170 ( .A(n11098), .B(n11097), .Z(n138) );
  NAND U171 ( .A(n138), .B(n11099), .Z(n139) );
  NANDN U172 ( .A(n11100), .B(n139), .Z(n140) );
  NANDN U173 ( .A(n11101), .B(n140), .Z(n141) );
  NAND U174 ( .A(n141), .B(n11102), .Z(n142) );
  ANDN U175 ( .B(n142), .A(n11103), .Z(n143) );
  NOR U176 ( .A(n143), .B(n11104), .Z(n144) );
  NAND U177 ( .A(n144), .B(n11105), .Z(n145) );
  NAND U178 ( .A(n145), .B(n11106), .Z(n146) );
  NOR U179 ( .A(n11108), .B(n11107), .Z(n147) );
  NAND U180 ( .A(n147), .B(n146), .Z(n148) );
  NAND U181 ( .A(n148), .B(n11109), .Z(n149) );
  NANDN U182 ( .A(n11110), .B(n149), .Z(n150) );
  NAND U183 ( .A(n150), .B(n11111), .Z(n151) );
  ANDN U184 ( .B(n151), .A(n11112), .Z(n152) );
  NAND U185 ( .A(n152), .B(n11113), .Z(n153) );
  NAND U186 ( .A(n153), .B(n11114), .Z(n154) );
  ANDN U187 ( .B(n154), .A(n11115), .Z(n155) );
  NAND U188 ( .A(n155), .B(n10015), .Z(n11117) );
  NANDN U189 ( .A(y[686]), .B(x[686]), .Z(n156) );
  AND U190 ( .A(n7475), .B(n156), .Z(n11136) );
  NANDN U191 ( .A(y[712]), .B(x[712]), .Z(n157) );
  AND U192 ( .A(n6506), .B(n157), .Z(n11177) );
  NANDN U193 ( .A(x[836]), .B(y[836]), .Z(n158) );
  ANDN U194 ( .B(n158), .A(n7691), .Z(n11425) );
  NANDN U195 ( .A(y[1103]), .B(x[1103]), .Z(n159) );
  NAND U196 ( .A(n159), .B(n6440), .Z(n12069) );
  NANDN U197 ( .A(y[1235]), .B(x[1235]), .Z(n160) );
  ANDN U198 ( .B(n160), .A(n8341), .Z(n12332) );
  NANDN U199 ( .A(x[1736]), .B(y[1736]), .Z(n161) );
  NANDN U200 ( .A(x[1737]), .B(y[1737]), .Z(n162) );
  NAND U201 ( .A(n161), .B(n162), .Z(n13430) );
  NANDN U202 ( .A(y[46]), .B(x[46]), .Z(n163) );
  AND U203 ( .A(n2106), .B(n163), .Z(n10057) );
  NANDN U204 ( .A(x[86]), .B(y[86]), .Z(n164) );
  NAND U205 ( .A(n164), .B(n1950), .Z(n10152) );
  NANDN U206 ( .A(y[143]), .B(x[143]), .Z(n165) );
  XNOR U207 ( .A(y[143]), .B(x[143]), .Z(n166) );
  NANDN U208 ( .A(x[142]), .B(y[142]), .Z(n167) );
  NAND U209 ( .A(n166), .B(n167), .Z(n168) );
  NAND U210 ( .A(n165), .B(n168), .Z(n10266) );
  NANDN U211 ( .A(y[167]), .B(x[167]), .Z(n169) );
  XNOR U212 ( .A(y[167]), .B(x[167]), .Z(n170) );
  NANDN U213 ( .A(x[166]), .B(y[166]), .Z(n171) );
  NAND U214 ( .A(n170), .B(n171), .Z(n172) );
  NAND U215 ( .A(n169), .B(n172), .Z(n10299) );
  NANDN U216 ( .A(y[208]), .B(x[208]), .Z(n173) );
  NAND U217 ( .A(n173), .B(n6911), .Z(n10383) );
  NANDN U218 ( .A(y[227]), .B(x[227]), .Z(n174) );
  NANDN U219 ( .A(y[228]), .B(x[228]), .Z(n175) );
  NANDN U220 ( .A(y[229]), .B(x[229]), .Z(n176) );
  NAND U221 ( .A(n175), .B(n176), .Z(n177) );
  ANDN U222 ( .B(n174), .A(n177), .Z(n178) );
  NANDN U223 ( .A(y[226]), .B(x[226]), .Z(n179) );
  XNOR U224 ( .A(x[227]), .B(y[227]), .Z(n180) );
  NANDN U225 ( .A(n179), .B(n180), .Z(n181) );
  NAND U226 ( .A(n178), .B(n181), .Z(n10399) );
  NANDN U227 ( .A(x[262]), .B(y[262]), .Z(n182) );
  AND U228 ( .A(n2512), .B(n182), .Z(n10449) );
  NANDN U229 ( .A(x[298]), .B(y[298]), .Z(n183) );
  AND U230 ( .A(n2575), .B(n183), .Z(n10533) );
  OR U231 ( .A(n10589), .B(n10590), .Z(n184) );
  AND U232 ( .A(n10591), .B(n184), .Z(n185) );
  NAND U233 ( .A(n10592), .B(n10595), .Z(n186) );
  NANDN U234 ( .A(n185), .B(n186), .Z(n187) );
  ANDN U235 ( .B(n187), .A(n10596), .Z(n188) );
  ANDN U236 ( .B(n10034), .A(n188), .Z(n189) );
  NAND U237 ( .A(n189), .B(n10035), .Z(n190) );
  ANDN U238 ( .B(n190), .A(n10597), .Z(n191) );
  NAND U239 ( .A(n191), .B(n10598), .Z(n192) );
  NAND U240 ( .A(n192), .B(n10599), .Z(n193) );
  ANDN U241 ( .B(n193), .A(n10600), .Z(n194) );
  NAND U242 ( .A(n194), .B(n10601), .Z(n195) );
  NAND U243 ( .A(n195), .B(n10602), .Z(n196) );
  ANDN U244 ( .B(n196), .A(n10603), .Z(n197) );
  NANDN U245 ( .A(n10604), .B(n197), .Z(n198) );
  NAND U246 ( .A(n198), .B(n10605), .Z(n199) );
  ANDN U247 ( .B(n199), .A(n10606), .Z(n200) );
  OR U248 ( .A(n10607), .B(n200), .Z(n201) );
  AND U249 ( .A(n10608), .B(n201), .Z(n10609) );
  NANDN U250 ( .A(x[372]), .B(y[372]), .Z(n202) );
  NAND U251 ( .A(n202), .B(n1635), .Z(n10658) );
  NANDN U252 ( .A(y[392]), .B(x[392]), .Z(n203) );
  NANDN U253 ( .A(n6554), .B(n203), .Z(n10696) );
  NANDN U254 ( .A(x[410]), .B(y[410]), .Z(n204) );
  AND U255 ( .A(n2814), .B(n204), .Z(n10725) );
  NANDN U256 ( .A(y[451]), .B(x[451]), .Z(n205) );
  NANDN U257 ( .A(y[452]), .B(x[452]), .Z(n206) );
  NANDN U258 ( .A(y[453]), .B(x[453]), .Z(n207) );
  NAND U259 ( .A(n206), .B(n207), .Z(n208) );
  ANDN U260 ( .B(n205), .A(n208), .Z(n209) );
  NANDN U261 ( .A(y[450]), .B(x[450]), .Z(n210) );
  XNOR U262 ( .A(x[451]), .B(y[451]), .Z(n211) );
  NANDN U263 ( .A(n210), .B(n211), .Z(n212) );
  NAND U264 ( .A(n209), .B(n212), .Z(n10791) );
  NANDN U265 ( .A(x[480]), .B(y[480]), .Z(n213) );
  NAND U266 ( .A(n213), .B(n1511), .Z(n10834) );
  NANDN U267 ( .A(x[499]), .B(y[499]), .Z(n214) );
  XNOR U268 ( .A(x[499]), .B(y[499]), .Z(n215) );
  NANDN U269 ( .A(y[498]), .B(x[498]), .Z(n216) );
  NAND U270 ( .A(n215), .B(n216), .Z(n217) );
  NAND U271 ( .A(n214), .B(n217), .Z(n10861) );
  NANDN U272 ( .A(x[532]), .B(y[532]), .Z(n218) );
  NAND U273 ( .A(n218), .B(n1457), .Z(n10932) );
  NANDN U274 ( .A(y[745]), .B(x[745]), .Z(n219) );
  NAND U275 ( .A(n219), .B(n11249), .Z(n7548) );
  NANDN U276 ( .A(x[580]), .B(y[580]), .Z(n220) );
  AND U277 ( .A(n3099), .B(n220), .Z(n10993) );
  NANDN U278 ( .A(y[599]), .B(x[599]), .Z(n221) );
  NANDN U279 ( .A(y[600]), .B(x[600]), .Z(n222) );
  NANDN U280 ( .A(y[601]), .B(x[601]), .Z(n223) );
  NAND U281 ( .A(n222), .B(n223), .Z(n224) );
  ANDN U282 ( .B(n221), .A(n224), .Z(n225) );
  NANDN U283 ( .A(y[598]), .B(x[598]), .Z(n226) );
  XNOR U284 ( .A(x[599]), .B(y[599]), .Z(n227) );
  NANDN U285 ( .A(n226), .B(n227), .Z(n228) );
  NAND U286 ( .A(n225), .B(n228), .Z(n11036) );
  NANDN U287 ( .A(x[628]), .B(y[628]), .Z(n229) );
  NAND U288 ( .A(n229), .B(n3201), .Z(n11080) );
  NAND U289 ( .A(n11117), .B(n11116), .Z(n230) );
  NAND U290 ( .A(n230), .B(n11118), .Z(n231) );
  ANDN U291 ( .B(n231), .A(n11119), .Z(n232) );
  NOR U292 ( .A(n232), .B(n11121), .Z(n233) );
  NAND U293 ( .A(n233), .B(n11120), .Z(n234) );
  AND U294 ( .A(n11122), .B(n234), .Z(n235) );
  OR U295 ( .A(n11123), .B(n235), .Z(n236) );
  NANDN U296 ( .A(n11124), .B(n236), .Z(n237) );
  NAND U297 ( .A(n237), .B(n11125), .Z(n238) );
  AND U298 ( .A(n11127), .B(n11128), .Z(n239) );
  NANDN U299 ( .A(n11126), .B(n238), .Z(n240) );
  NAND U300 ( .A(n239), .B(n240), .Z(n241) );
  NANDN U301 ( .A(n11129), .B(n241), .Z(n242) );
  NANDN U302 ( .A(n11130), .B(n242), .Z(n243) );
  ANDN U303 ( .B(n243), .A(n11131), .Z(n244) );
  OR U304 ( .A(n11132), .B(n244), .Z(n245) );
  NANDN U305 ( .A(n11133), .B(n245), .Z(n246) );
  NANDN U306 ( .A(n11134), .B(n246), .Z(n247) );
  NAND U307 ( .A(n247), .B(n11135), .Z(n11137) );
  NANDN U308 ( .A(x[724]), .B(y[724]), .Z(n248) );
  NAND U309 ( .A(n248), .B(n1286), .Z(n11210) );
  NANDN U310 ( .A(x[769]), .B(y[769]), .Z(n249) );
  XNOR U311 ( .A(x[769]), .B(y[769]), .Z(n250) );
  NANDN U312 ( .A(y[768]), .B(x[768]), .Z(n251) );
  NAND U313 ( .A(n250), .B(n251), .Z(n252) );
  NAND U314 ( .A(n249), .B(n252), .Z(n11297) );
  NANDN U315 ( .A(x[828]), .B(y[828]), .Z(n253) );
  NANDN U316 ( .A(n7669), .B(n253), .Z(n7661) );
  NANDN U317 ( .A(n11382), .B(n11381), .Z(n254) );
  NAND U318 ( .A(n254), .B(n11383), .Z(n255) );
  ANDN U319 ( .B(n255), .A(n11384), .Z(n256) );
  NANDN U320 ( .A(n256), .B(n11385), .Z(n257) );
  ANDN U321 ( .B(n257), .A(n11386), .Z(n258) );
  ANDN U322 ( .B(n11389), .A(n11388), .Z(n259) );
  OR U323 ( .A(n11387), .B(n258), .Z(n260) );
  NAND U324 ( .A(n259), .B(n260), .Z(n261) );
  NANDN U325 ( .A(n10010), .B(n10009), .Z(n262) );
  NAND U326 ( .A(n262), .B(n261), .Z(n263) );
  NANDN U327 ( .A(n11390), .B(n263), .Z(n264) );
  NAND U328 ( .A(n264), .B(n11391), .Z(n265) );
  NANDN U329 ( .A(n11392), .B(n265), .Z(n266) );
  AND U330 ( .A(n11393), .B(n266), .Z(n267) );
  NANDN U331 ( .A(n267), .B(n11394), .Z(n268) );
  ANDN U332 ( .B(n268), .A(n11395), .Z(n269) );
  NOR U333 ( .A(n269), .B(n11396), .Z(n270) );
  NAND U334 ( .A(n270), .B(n11397), .Z(n271) );
  AND U335 ( .A(n11398), .B(n271), .Z(n11399) );
  NANDN U336 ( .A(y[1105]), .B(x[1105]), .Z(n272) );
  NANDN U337 ( .A(y[1104]), .B(x[1104]), .Z(n273) );
  NAND U338 ( .A(n272), .B(n273), .Z(n12074) );
  NAND U339 ( .A(n8142), .B(n8141), .Z(n12124) );
  NANDN U340 ( .A(x[1152]), .B(y[1152]), .Z(n274) );
  NANDN U341 ( .A(x[1151]), .B(y[1151]), .Z(n275) );
  NAND U342 ( .A(n274), .B(n275), .Z(n12158) );
  NAND U343 ( .A(n12312), .B(n12311), .Z(n276) );
  NANDN U344 ( .A(n12313), .B(n276), .Z(n277) );
  NANDN U345 ( .A(n12314), .B(n277), .Z(n278) );
  NAND U346 ( .A(n12316), .B(n12315), .Z(n279) );
  NANDN U347 ( .A(n278), .B(n279), .Z(n280) );
  ANDN U348 ( .B(n280), .A(n12317), .Z(n281) );
  OR U349 ( .A(n12318), .B(n281), .Z(n282) );
  NAND U350 ( .A(n282), .B(n12319), .Z(n283) );
  AND U351 ( .A(n12320), .B(n283), .Z(n284) );
  NANDN U352 ( .A(n284), .B(n12321), .Z(n285) );
  NANDN U353 ( .A(n12322), .B(n285), .Z(n286) );
  NAND U354 ( .A(n286), .B(n12323), .Z(n287) );
  NAND U355 ( .A(n287), .B(n12324), .Z(n288) );
  NAND U356 ( .A(n288), .B(n12325), .Z(n289) );
  ANDN U357 ( .B(n289), .A(n12326), .Z(n290) );
  NANDN U358 ( .A(n290), .B(n12327), .Z(n291) );
  NAND U359 ( .A(n291), .B(n12328), .Z(n292) );
  NAND U360 ( .A(n292), .B(n12329), .Z(n293) );
  NAND U361 ( .A(n293), .B(n12330), .Z(n12331) );
  NANDN U362 ( .A(x[1552]), .B(y[1552]), .Z(n294) );
  AND U363 ( .A(n5169), .B(n294), .Z(n9996) );
  NANDN U364 ( .A(y[1740]), .B(x[1740]), .Z(n295) );
  AND U365 ( .A(n9336), .B(n295), .Z(n13433) );
  NANDN U366 ( .A(y[1790]), .B(x[1790]), .Z(n296) );
  ANDN U367 ( .B(n296), .A(n9470), .Z(n13548) );
  NANDN U368 ( .A(y[1796]), .B(x[1796]), .Z(n297) );
  NAND U369 ( .A(n297), .B(n5639), .Z(n13560) );
  XNOR U370 ( .A(y[1851]), .B(x[1851]), .Z(n13691) );
  NANDN U371 ( .A(n9695), .B(n9694), .Z(n298) );
  NANDN U372 ( .A(n9696), .B(n298), .Z(n299) );
  ANDN U373 ( .B(n299), .A(n9697), .Z(n300) );
  NAND U374 ( .A(n300), .B(n9698), .Z(n13774) );
  NANDN U375 ( .A(n13901), .B(n13900), .Z(n301) );
  NANDN U376 ( .A(n13902), .B(n301), .Z(n302) );
  ANDN U377 ( .B(n302), .A(n13903), .Z(n303) );
  OR U378 ( .A(n13904), .B(n303), .Z(n304) );
  NAND U379 ( .A(n304), .B(n13905), .Z(n305) );
  NANDN U380 ( .A(n13906), .B(n305), .Z(n306) );
  ANDN U381 ( .B(n13908), .A(n13909), .Z(n307) );
  NANDN U382 ( .A(n13907), .B(n306), .Z(n308) );
  NAND U383 ( .A(n307), .B(n308), .Z(n309) );
  NOR U384 ( .A(n13911), .B(n13910), .Z(n310) );
  NAND U385 ( .A(n310), .B(n309), .Z(n311) );
  NANDN U386 ( .A(n13912), .B(n311), .Z(n312) );
  NANDN U387 ( .A(n13913), .B(n312), .Z(n313) );
  NAND U388 ( .A(n313), .B(n13914), .Z(n314) );
  ANDN U389 ( .B(n314), .A(n13915), .Z(n315) );
  NANDN U390 ( .A(n315), .B(n13916), .Z(n316) );
  NANDN U391 ( .A(n13917), .B(n316), .Z(n317) );
  NAND U392 ( .A(n317), .B(n13918), .Z(n318) );
  NANDN U393 ( .A(n13919), .B(n318), .Z(n13921) );
  NAND U394 ( .A(n6093), .B(n6092), .Z(n14030) );
  ANDN U395 ( .B(y[2040]), .A(x[2040]), .Z(n9973) );
  NAND U396 ( .A(n10052), .B(n10051), .Z(n10053) );
  NANDN U397 ( .A(x[76]), .B(y[76]), .Z(n319) );
  NAND U398 ( .A(n319), .B(n2168), .Z(n10128) );
  OR U399 ( .A(y[104]), .B(n1927), .Z(n6787) );
  NANDN U400 ( .A(x[104]), .B(y[104]), .Z(n320) );
  NANDN U401 ( .A(x[105]), .B(y[105]), .Z(n321) );
  NAND U402 ( .A(n320), .B(n321), .Z(n10196) );
  NAND U403 ( .A(n10283), .B(n10282), .Z(n322) );
  NANDN U404 ( .A(n10284), .B(n322), .Z(n323) );
  AND U405 ( .A(n10285), .B(n323), .Z(n324) );
  ANDN U406 ( .B(n10044), .A(n324), .Z(n325) );
  NAND U407 ( .A(n325), .B(n10045), .Z(n326) );
  ANDN U408 ( .B(n326), .A(n10286), .Z(n327) );
  OR U409 ( .A(n10287), .B(n327), .Z(n328) );
  NAND U410 ( .A(n328), .B(n10288), .Z(n329) );
  NANDN U411 ( .A(n10289), .B(n329), .Z(n330) );
  NAND U412 ( .A(n330), .B(n10290), .Z(n331) );
  AND U413 ( .A(n10292), .B(n331), .Z(n332) );
  NANDN U414 ( .A(n10291), .B(n332), .Z(n333) );
  NAND U415 ( .A(n333), .B(n10293), .Z(n334) );
  NANDN U416 ( .A(n10294), .B(n334), .Z(n335) );
  AND U417 ( .A(n10295), .B(n335), .Z(n336) );
  OR U418 ( .A(n10296), .B(n336), .Z(n337) );
  NAND U419 ( .A(n337), .B(n10297), .Z(n338) );
  NANDN U420 ( .A(n10298), .B(n338), .Z(n339) );
  NAND U421 ( .A(n339), .B(n10299), .Z(n10301) );
  NANDN U422 ( .A(n10381), .B(n10380), .Z(n340) );
  NAND U423 ( .A(n340), .B(n10382), .Z(n341) );
  ANDN U424 ( .B(n341), .A(n10383), .Z(n342) );
  AND U425 ( .A(n10043), .B(n10042), .Z(n343) );
  OR U426 ( .A(n10384), .B(n342), .Z(n344) );
  AND U427 ( .A(n343), .B(n344), .Z(n345) );
  OR U428 ( .A(n10385), .B(n345), .Z(n346) );
  NANDN U429 ( .A(n10386), .B(n346), .Z(n347) );
  NAND U430 ( .A(n347), .B(n10387), .Z(n348) );
  NANDN U431 ( .A(n10388), .B(n348), .Z(n349) );
  NAND U432 ( .A(n349), .B(n10389), .Z(n350) );
  ANDN U433 ( .B(n350), .A(n10390), .Z(n351) );
  AND U434 ( .A(n10041), .B(n10040), .Z(n352) );
  NANDN U435 ( .A(n351), .B(n10391), .Z(n353) );
  AND U436 ( .A(n352), .B(n353), .Z(n354) );
  OR U437 ( .A(n10392), .B(n354), .Z(n355) );
  NANDN U438 ( .A(n10393), .B(n355), .Z(n356) );
  NANDN U439 ( .A(n10394), .B(n356), .Z(n10396) );
  NANDN U440 ( .A(x[267]), .B(y[267]), .Z(n357) );
  NANDN U441 ( .A(x[268]), .B(y[268]), .Z(n358) );
  NANDN U442 ( .A(x[269]), .B(y[269]), .Z(n359) );
  NAND U443 ( .A(n358), .B(n359), .Z(n360) );
  ANDN U444 ( .B(n357), .A(n360), .Z(n361) );
  NANDN U445 ( .A(x[266]), .B(y[266]), .Z(n362) );
  XNOR U446 ( .A(y[267]), .B(x[267]), .Z(n363) );
  NANDN U447 ( .A(n362), .B(n363), .Z(n364) );
  NAND U448 ( .A(n361), .B(n364), .Z(n10460) );
  NANDN U449 ( .A(x[278]), .B(y[278]), .Z(n365) );
  AND U450 ( .A(n2538), .B(n365), .Z(n10485) );
  NANDN U451 ( .A(x[306]), .B(y[306]), .Z(n366) );
  AND U452 ( .A(n2589), .B(n366), .Z(n10553) );
  NAND U453 ( .A(n10594), .B(n10593), .Z(n10595) );
  NANDN U454 ( .A(y[416]), .B(x[416]), .Z(n367) );
  NAND U455 ( .A(n367), .B(n6538), .Z(n7154) );
  NANDN U456 ( .A(n10648), .B(n10647), .Z(n368) );
  NANDN U457 ( .A(n10649), .B(n368), .Z(n369) );
  NANDN U458 ( .A(n10650), .B(n369), .Z(n370) );
  NANDN U459 ( .A(n370), .B(n10651), .Z(n371) );
  NANDN U460 ( .A(n10033), .B(n10032), .Z(n372) );
  AND U461 ( .A(n371), .B(n372), .Z(n373) );
  OR U462 ( .A(n10652), .B(n373), .Z(n374) );
  NANDN U463 ( .A(n10653), .B(n374), .Z(n375) );
  ANDN U464 ( .B(n375), .A(n10654), .Z(n376) );
  NAND U465 ( .A(n376), .B(n10655), .Z(n377) );
  NAND U466 ( .A(n377), .B(n10656), .Z(n378) );
  NANDN U467 ( .A(n10657), .B(n378), .Z(n379) );
  NANDN U468 ( .A(y[372]), .B(x[372]), .Z(n380) );
  NANDN U469 ( .A(n379), .B(n380), .Z(n381) );
  ANDN U470 ( .B(n381), .A(n10658), .Z(n382) );
  NOR U471 ( .A(n382), .B(n10659), .Z(n383) );
  NANDN U472 ( .A(n10660), .B(n383), .Z(n384) );
  NANDN U473 ( .A(n10661), .B(n384), .Z(n385) );
  NANDN U474 ( .A(n10662), .B(n385), .Z(n10664) );
  NANDN U475 ( .A(n10026), .B(n10027), .Z(n386) );
  NAND U476 ( .A(n10741), .B(n10742), .Z(n387) );
  NAND U477 ( .A(n387), .B(n10743), .Z(n388) );
  NANDN U478 ( .A(n10744), .B(n388), .Z(n389) );
  NAND U479 ( .A(n389), .B(n10745), .Z(n390) );
  NANDN U480 ( .A(n10746), .B(n390), .Z(n391) );
  AND U481 ( .A(n10747), .B(n391), .Z(n392) );
  OR U482 ( .A(n10748), .B(n392), .Z(n393) );
  NAND U483 ( .A(n393), .B(n10749), .Z(n394) );
  NAND U484 ( .A(n394), .B(n10750), .Z(n395) );
  NAND U485 ( .A(n395), .B(n10751), .Z(n396) );
  AND U486 ( .A(n10028), .B(n396), .Z(n397) );
  NAND U487 ( .A(n397), .B(n10029), .Z(n398) );
  NAND U488 ( .A(n398), .B(n10752), .Z(n399) );
  NANDN U489 ( .A(n10753), .B(n399), .Z(n400) );
  AND U490 ( .A(n10754), .B(n400), .Z(n401) );
  AND U491 ( .A(n10024), .B(n10025), .Z(n402) );
  OR U492 ( .A(n386), .B(n401), .Z(n403) );
  AND U493 ( .A(n402), .B(n403), .Z(n10755) );
  NANDN U494 ( .A(y[469]), .B(x[469]), .Z(n404) );
  NANDN U495 ( .A(y[470]), .B(x[470]), .Z(n405) );
  NANDN U496 ( .A(y[471]), .B(x[471]), .Z(n406) );
  NAND U497 ( .A(n405), .B(n406), .Z(n407) );
  ANDN U498 ( .B(n404), .A(n407), .Z(n408) );
  NANDN U499 ( .A(y[468]), .B(x[468]), .Z(n409) );
  XNOR U500 ( .A(x[469]), .B(y[469]), .Z(n410) );
  NANDN U501 ( .A(n409), .B(n410), .Z(n411) );
  NAND U502 ( .A(n408), .B(n411), .Z(n10819) );
  NANDN U503 ( .A(x[506]), .B(y[506]), .Z(n412) );
  NAND U504 ( .A(n412), .B(n1478), .Z(n10880) );
  NANDN U505 ( .A(y[522]), .B(x[522]), .Z(n413) );
  NANDN U506 ( .A(n1460), .B(n413), .Z(n7269) );
  NANDN U507 ( .A(n10951), .B(n10952), .Z(n414) );
  NANDN U508 ( .A(n10953), .B(n414), .Z(n415) );
  NAND U509 ( .A(n415), .B(n10954), .Z(n416) );
  ANDN U510 ( .B(n10023), .A(n10022), .Z(n417) );
  NANDN U511 ( .A(n10955), .B(n416), .Z(n418) );
  NAND U512 ( .A(n417), .B(n418), .Z(n419) );
  NAND U513 ( .A(n10020), .B(n10021), .Z(n420) );
  NAND U514 ( .A(n420), .B(n419), .Z(n421) );
  NANDN U515 ( .A(n10956), .B(n421), .Z(n422) );
  ANDN U516 ( .B(n10959), .A(n10958), .Z(n423) );
  NANDN U517 ( .A(n10957), .B(n422), .Z(n424) );
  NAND U518 ( .A(n423), .B(n424), .Z(n425) );
  NAND U519 ( .A(n425), .B(n10960), .Z(n426) );
  NANDN U520 ( .A(n10961), .B(n426), .Z(n427) );
  AND U521 ( .A(n10962), .B(n427), .Z(n428) );
  OR U522 ( .A(n10963), .B(n428), .Z(n429) );
  NAND U523 ( .A(n429), .B(n10964), .Z(n430) );
  NANDN U524 ( .A(n10965), .B(n430), .Z(n431) );
  NAND U525 ( .A(n431), .B(n10966), .Z(n10968) );
  NANDN U526 ( .A(n10019), .B(n10018), .Z(n11006) );
  NOR U527 ( .A(n11081), .B(n11082), .Z(n432) );
  NANDN U528 ( .A(n11080), .B(n11079), .Z(n433) );
  AND U529 ( .A(n432), .B(n433), .Z(n434) );
  OR U530 ( .A(n11083), .B(n434), .Z(n435) );
  NAND U531 ( .A(n435), .B(n11084), .Z(n436) );
  NANDN U532 ( .A(n11085), .B(n436), .Z(n437) );
  NANDN U533 ( .A(n11086), .B(n437), .Z(n438) );
  NANDN U534 ( .A(n11087), .B(n438), .Z(n439) );
  ANDN U535 ( .B(n439), .A(n11088), .Z(n440) );
  ANDN U536 ( .B(n11091), .A(n11090), .Z(n441) );
  OR U537 ( .A(n11089), .B(n440), .Z(n442) );
  AND U538 ( .A(n441), .B(n442), .Z(n443) );
  NANDN U539 ( .A(n443), .B(n11092), .Z(n444) );
  NANDN U540 ( .A(n11093), .B(n444), .Z(n445) );
  NANDN U541 ( .A(n11094), .B(n445), .Z(n446) );
  AND U542 ( .A(n10016), .B(n10017), .Z(n447) );
  NAND U543 ( .A(n447), .B(n446), .Z(n448) );
  NANDN U544 ( .A(n11095), .B(n448), .Z(n449) );
  ANDN U545 ( .B(n449), .A(n11096), .Z(n11097) );
  NAND U546 ( .A(n11137), .B(n11136), .Z(n450) );
  NANDN U547 ( .A(n11138), .B(n450), .Z(n451) );
  AND U548 ( .A(n11139), .B(n451), .Z(n452) );
  OR U549 ( .A(n11140), .B(n452), .Z(n453) );
  NAND U550 ( .A(n453), .B(n11141), .Z(n454) );
  NANDN U551 ( .A(n11142), .B(n454), .Z(n455) );
  NAND U552 ( .A(n455), .B(n11143), .Z(n456) );
  NANDN U553 ( .A(n11144), .B(n456), .Z(n457) );
  AND U554 ( .A(n11145), .B(n457), .Z(n458) );
  NAND U555 ( .A(n458), .B(n11146), .Z(n459) );
  NAND U556 ( .A(n459), .B(n11147), .Z(n460) );
  ANDN U557 ( .B(n460), .A(n11148), .Z(n461) );
  ANDN U558 ( .B(n10013), .A(n10014), .Z(n462) );
  OR U559 ( .A(n11149), .B(n461), .Z(n463) );
  AND U560 ( .A(n462), .B(n463), .Z(n464) );
  OR U561 ( .A(n11150), .B(n464), .Z(n465) );
  NANDN U562 ( .A(n11151), .B(n465), .Z(n466) );
  ANDN U563 ( .B(n466), .A(n11152), .Z(n11154) );
  ANDN U564 ( .B(y[734]), .A(x[734]), .Z(n467) );
  NANDN U565 ( .A(x[736]), .B(y[736]), .Z(n468) );
  AND U566 ( .A(n1269), .B(n468), .Z(n469) );
  OR U567 ( .A(y[735]), .B(n467), .Z(n470) );
  XOR U568 ( .A(y[735]), .B(n467), .Z(n471) );
  NAND U569 ( .A(n471), .B(x[735]), .Z(n472) );
  NAND U570 ( .A(n470), .B(n472), .Z(n473) );
  AND U571 ( .A(n469), .B(n473), .Z(n11230) );
  NANDN U572 ( .A(y[752]), .B(x[752]), .Z(n474) );
  NANDN U573 ( .A(n7563), .B(n474), .Z(n6501) );
  NANDN U574 ( .A(x[770]), .B(y[770]), .Z(n475) );
  AND U575 ( .A(n3477), .B(n475), .Z(n11301) );
  NANDN U576 ( .A(x[792]), .B(y[792]), .Z(n476) );
  AND U577 ( .A(n3521), .B(n476), .Z(n11350) );
  NANDN U578 ( .A(y[823]), .B(x[823]), .Z(n477) );
  XNOR U579 ( .A(y[823]), .B(x[823]), .Z(n478) );
  NANDN U580 ( .A(x[822]), .B(y[822]), .Z(n479) );
  NAND U581 ( .A(n478), .B(n479), .Z(n480) );
  NAND U582 ( .A(n477), .B(n480), .Z(n11401) );
  OR U583 ( .A(y[922]), .B(n6481), .Z(n6480) );
  NANDN U584 ( .A(y[1055]), .B(x[1055]), .Z(n481) );
  ANDN U585 ( .B(n481), .A(n8012), .Z(n11963) );
  OR U586 ( .A(x[1062]), .B(n1034), .Z(n8021) );
  NANDN U587 ( .A(x[1071]), .B(y[1071]), .Z(n482) );
  XNOR U588 ( .A(x[1071]), .B(y[1071]), .Z(n483) );
  NANDN U589 ( .A(y[1070]), .B(x[1070]), .Z(n484) );
  NAND U590 ( .A(n483), .B(n484), .Z(n485) );
  NAND U591 ( .A(n482), .B(n485), .Z(n12001) );
  OR U592 ( .A(x[1127]), .B(n1004), .Z(n6435) );
  OR U593 ( .A(x[1134]), .B(n1001), .Z(n8148) );
  NANDN U594 ( .A(x[1098]), .B(y[1098]), .Z(n486) );
  NANDN U595 ( .A(n6443), .B(n486), .Z(n12056) );
  NAND U596 ( .A(n12135), .B(n12136), .Z(n487) );
  NAND U597 ( .A(n487), .B(n12137), .Z(n488) );
  ANDN U598 ( .B(n488), .A(n12138), .Z(n489) );
  NANDN U599 ( .A(n489), .B(n12139), .Z(n490) );
  NAND U600 ( .A(n490), .B(n12140), .Z(n491) );
  NANDN U601 ( .A(n12141), .B(n491), .Z(n492) );
  NANDN U602 ( .A(n12142), .B(n492), .Z(n493) );
  NAND U603 ( .A(n493), .B(n12143), .Z(n494) );
  AND U604 ( .A(n12144), .B(n494), .Z(n495) );
  OR U605 ( .A(n12145), .B(n495), .Z(n496) );
  NANDN U606 ( .A(n12146), .B(n496), .Z(n497) );
  NANDN U607 ( .A(n12147), .B(n497), .Z(n498) );
  NANDN U608 ( .A(n498), .B(n12148), .Z(n499) );
  NANDN U609 ( .A(n10003), .B(n10002), .Z(n500) );
  AND U610 ( .A(n499), .B(n500), .Z(n501) );
  NAND U611 ( .A(n501), .B(n12149), .Z(n502) );
  NANDN U612 ( .A(n12150), .B(n502), .Z(n503) );
  NAND U613 ( .A(n503), .B(n12151), .Z(n504) );
  NANDN U614 ( .A(n12152), .B(n504), .Z(n12153) );
  NANDN U615 ( .A(x[1170]), .B(y[1170]), .Z(n505) );
  ANDN U616 ( .B(n505), .A(n8225), .Z(n12199) );
  NANDN U617 ( .A(x[1205]), .B(y[1205]), .Z(n506) );
  XNOR U618 ( .A(x[1205]), .B(y[1205]), .Z(n507) );
  NANDN U619 ( .A(y[1204]), .B(x[1204]), .Z(n508) );
  NAND U620 ( .A(n507), .B(n508), .Z(n509) );
  NAND U621 ( .A(n506), .B(n509), .Z(n12277) );
  NANDN U622 ( .A(x[1224]), .B(y[1224]), .Z(n510) );
  NANDN U623 ( .A(x[1223]), .B(y[1223]), .Z(n511) );
  NAND U624 ( .A(n510), .B(n511), .Z(n12318) );
  NANDN U625 ( .A(n12370), .B(n12369), .Z(n512) );
  NANDN U626 ( .A(n12371), .B(n512), .Z(n513) );
  ANDN U627 ( .B(n513), .A(n12372), .Z(n514) );
  NANDN U628 ( .A(n514), .B(n12373), .Z(n515) );
  NAND U629 ( .A(n515), .B(n12374), .Z(n516) );
  NAND U630 ( .A(n516), .B(n12375), .Z(n517) );
  NAND U631 ( .A(n517), .B(n12376), .Z(n518) );
  NAND U632 ( .A(n518), .B(n12377), .Z(n519) );
  AND U633 ( .A(n12378), .B(n519), .Z(n520) );
  ANDN U634 ( .B(n12379), .A(n520), .Z(n521) );
  NANDN U635 ( .A(n12381), .B(n12380), .Z(n522) );
  NAND U636 ( .A(n521), .B(n522), .Z(n523) );
  NAND U637 ( .A(n523), .B(n12382), .Z(n524) );
  NAND U638 ( .A(n524), .B(n12383), .Z(n525) );
  ANDN U639 ( .B(n525), .A(n12384), .Z(n526) );
  NANDN U640 ( .A(n526), .B(n12385), .Z(n527) );
  NANDN U641 ( .A(n12386), .B(n527), .Z(n528) );
  NANDN U642 ( .A(n12387), .B(n528), .Z(n529) );
  NANDN U643 ( .A(n12388), .B(n529), .Z(n12390) );
  NANDN U644 ( .A(y[1367]), .B(x[1367]), .Z(n530) );
  ANDN U645 ( .B(n530), .A(n8588), .Z(n12606) );
  NANDN U646 ( .A(x[1382]), .B(y[1382]), .Z(n531) );
  NANDN U647 ( .A(x[1381]), .B(y[1381]), .Z(n532) );
  NAND U648 ( .A(n531), .B(n532), .Z(n12632) );
  NANDN U649 ( .A(y[1406]), .B(x[1406]), .Z(n533) );
  NANDN U650 ( .A(y[1408]), .B(x[1408]), .Z(n534) );
  NANDN U651 ( .A(y[1409]), .B(x[1409]), .Z(n535) );
  NAND U652 ( .A(n534), .B(n535), .Z(n536) );
  NANDN U653 ( .A(y[1407]), .B(x[1407]), .Z(n537) );
  ANDN U654 ( .B(n537), .A(n536), .Z(n538) );
  XNOR U655 ( .A(x[1407]), .B(y[1407]), .Z(n539) );
  NANDN U656 ( .A(n533), .B(n539), .Z(n540) );
  NAND U657 ( .A(n538), .B(n540), .Z(n12689) );
  NANDN U658 ( .A(y[1463]), .B(x[1463]), .Z(n541) );
  ANDN U659 ( .B(n541), .A(n8771), .Z(n12816) );
  NANDN U660 ( .A(n6300), .B(n6299), .Z(n12866) );
  NANDN U661 ( .A(y[1540]), .B(x[1540]), .Z(n542) );
  NANDN U662 ( .A(x[1541]), .B(y[1541]), .Z(n543) );
  XNOR U663 ( .A(x[1541]), .B(y[1541]), .Z(n544) );
  NAND U664 ( .A(n544), .B(n542), .Z(n545) );
  NAND U665 ( .A(n543), .B(n545), .Z(n12961) );
  NANDN U666 ( .A(x[1560]), .B(y[1560]), .Z(n546) );
  NANDN U667 ( .A(x[1559]), .B(y[1559]), .Z(n547) );
  NAND U668 ( .A(n546), .B(n547), .Z(n13011) );
  OR U669 ( .A(y[1620]), .B(n833), .Z(n6259) );
  NANDN U670 ( .A(x[1634]), .B(y[1634]), .Z(n548) );
  NAND U671 ( .A(n548), .B(n9086), .Z(n9082) );
  ANDN U672 ( .B(n5335), .A(n9078), .Z(n13190) );
  OR U673 ( .A(x[1666]), .B(n6242), .Z(n9156) );
  NANDN U674 ( .A(y[1652]), .B(x[1652]), .Z(n549) );
  NAND U675 ( .A(n549), .B(n6243), .Z(n13235) );
  OR U676 ( .A(x[1673]), .B(n6234), .Z(n6233) );
  OR U677 ( .A(y[1701]), .B(n6212), .Z(n9251) );
  NAND U678 ( .A(n13421), .B(n13420), .Z(n550) );
  NAND U679 ( .A(n550), .B(n13422), .Z(n551) );
  AND U680 ( .A(n13423), .B(n551), .Z(n552) );
  OR U681 ( .A(n13424), .B(n552), .Z(n553) );
  NANDN U682 ( .A(n13425), .B(n553), .Z(n554) );
  NANDN U683 ( .A(n13426), .B(n554), .Z(n555) );
  NAND U684 ( .A(n555), .B(n13427), .Z(n556) );
  NAND U685 ( .A(n556), .B(n13428), .Z(n557) );
  ANDN U686 ( .B(n557), .A(n13429), .Z(n558) );
  OR U687 ( .A(n13430), .B(n558), .Z(n559) );
  NANDN U688 ( .A(n13431), .B(n559), .Z(n560) );
  NAND U689 ( .A(n560), .B(n13432), .Z(n561) );
  XNOR U690 ( .A(x[1739]), .B(y[1739]), .Z(n562) );
  NANDN U691 ( .A(n561), .B(n562), .Z(n563) );
  AND U692 ( .A(n13433), .B(n563), .Z(n564) );
  NANDN U693 ( .A(n564), .B(n13434), .Z(n565) );
  NAND U694 ( .A(n565), .B(n13435), .Z(n566) );
  NANDN U695 ( .A(n13436), .B(n566), .Z(n567) );
  NANDN U696 ( .A(n13437), .B(n567), .Z(n13438) );
  OR U697 ( .A(y[1813]), .B(n6155), .Z(n9521) );
  OR U698 ( .A(n13558), .B(n13559), .Z(n568) );
  NANDN U699 ( .A(n13560), .B(n568), .Z(n569) );
  ANDN U700 ( .B(n569), .A(n13561), .Z(n570) );
  NANDN U701 ( .A(x[1798]), .B(y[1798]), .Z(n571) );
  AND U702 ( .A(n13562), .B(n571), .Z(n572) );
  XNOR U703 ( .A(y[1798]), .B(x[1798]), .Z(n573) );
  NANDN U704 ( .A(n570), .B(n573), .Z(n574) );
  NAND U705 ( .A(n572), .B(n574), .Z(n575) );
  AND U706 ( .A(n9990), .B(n9991), .Z(n576) );
  NAND U707 ( .A(n576), .B(n575), .Z(n577) );
  NAND U708 ( .A(n577), .B(n13563), .Z(n578) );
  NAND U709 ( .A(n578), .B(n13564), .Z(n579) );
  NAND U710 ( .A(n579), .B(n13565), .Z(n580) );
  ANDN U711 ( .B(n580), .A(n13566), .Z(n581) );
  NANDN U712 ( .A(n581), .B(n13567), .Z(n582) );
  AND U713 ( .A(n13568), .B(n582), .Z(n583) );
  OR U714 ( .A(n13569), .B(n583), .Z(n584) );
  NANDN U715 ( .A(n13570), .B(n584), .Z(n585) );
  NANDN U716 ( .A(n13571), .B(n585), .Z(n13573) );
  ANDN U717 ( .B(x[1868]), .A(y[1868]), .Z(n13729) );
  OR U718 ( .A(x[1876]), .B(n6138), .Z(n9675) );
  NANDN U719 ( .A(n13806), .B(n13807), .Z(n586) );
  NANDN U720 ( .A(n13808), .B(n586), .Z(n587) );
  ANDN U721 ( .B(n587), .A(n13809), .Z(n588) );
  NANDN U722 ( .A(n588), .B(n13810), .Z(n589) );
  NANDN U723 ( .A(n13811), .B(n589), .Z(n590) );
  NAND U724 ( .A(n590), .B(n13812), .Z(n591) );
  NANDN U725 ( .A(n13813), .B(n591), .Z(n592) );
  NAND U726 ( .A(n592), .B(n13814), .Z(n593) );
  ANDN U727 ( .B(n593), .A(n13815), .Z(n594) );
  NANDN U728 ( .A(n594), .B(n13816), .Z(n595) );
  NANDN U729 ( .A(n13817), .B(n595), .Z(n596) );
  NANDN U730 ( .A(n13818), .B(n596), .Z(n597) );
  ANDN U731 ( .B(n13820), .A(n13819), .Z(n598) );
  NAND U732 ( .A(n598), .B(n597), .Z(n599) );
  NANDN U733 ( .A(n13821), .B(n599), .Z(n600) );
  NAND U734 ( .A(n600), .B(n13822), .Z(n601) );
  AND U735 ( .A(n9981), .B(n601), .Z(n602) );
  NAND U736 ( .A(n602), .B(n9982), .Z(n603) );
  NANDN U737 ( .A(n13823), .B(n603), .Z(n13824) );
  NANDN U738 ( .A(x[1954]), .B(y[1954]), .Z(n604) );
  NAND U739 ( .A(n604), .B(n9809), .Z(n13904) );
  NAND U740 ( .A(n13957), .B(n13956), .Z(n605) );
  NANDN U741 ( .A(n13958), .B(n605), .Z(n606) );
  NAND U742 ( .A(n606), .B(n13959), .Z(n607) );
  NAND U743 ( .A(n607), .B(n13960), .Z(n608) );
  NAND U744 ( .A(n608), .B(n13961), .Z(n609) );
  ANDN U745 ( .B(n609), .A(n13962), .Z(n610) );
  ANDN U746 ( .B(n9977), .A(n610), .Z(n611) );
  NAND U747 ( .A(n611), .B(n9978), .Z(n612) );
  AND U748 ( .A(n13963), .B(n612), .Z(n613) );
  OR U749 ( .A(n13964), .B(n613), .Z(n614) );
  NANDN U750 ( .A(n13965), .B(n614), .Z(n615) );
  NAND U751 ( .A(n615), .B(n13966), .Z(n616) );
  NAND U752 ( .A(n616), .B(n13967), .Z(n617) );
  NAND U753 ( .A(n617), .B(n13968), .Z(n618) );
  ANDN U754 ( .B(n618), .A(n13969), .Z(n619) );
  OR U755 ( .A(n13970), .B(n619), .Z(n620) );
  NANDN U756 ( .A(n13971), .B(n620), .Z(n621) );
  NAND U757 ( .A(n621), .B(n13972), .Z(n622) );
  NAND U758 ( .A(n622), .B(n13973), .Z(n13975) );
  NANDN U759 ( .A(y[2028]), .B(x[2028]), .Z(n14035) );
  NANDN U760 ( .A(y[2041]), .B(x[2041]), .Z(n9971) );
  IV U761 ( .A(ebreg), .Z(e) );
  NANDN U762 ( .A(y[2044]), .B(x[2044]), .Z(n624) );
  NANDN U763 ( .A(y[2043]), .B(x[2043]), .Z(n623) );
  AND U764 ( .A(n624), .B(n623), .Z(n14067) );
  NANDN U765 ( .A(x[2046]), .B(y[2046]), .Z(n626) );
  NANDN U766 ( .A(x[2047]), .B(y[2047]), .Z(n625) );
  NAND U767 ( .A(n626), .B(n625), .Z(n14073) );
  ANDN U768 ( .B(n14067), .A(n14073), .Z(n627) );
  ANDN U769 ( .B(y[2038]), .A(x[2038]), .Z(n14055) );
  ANDN U770 ( .B(n627), .A(n14055), .Z(n630) );
  XNOR U771 ( .A(y[2041]), .B(x[2041]), .Z(n628) );
  NANDN U772 ( .A(y[2039]), .B(x[2039]), .Z(n9974) );
  NAND U773 ( .A(n628), .B(n9974), .Z(n629) );
  ANDN U774 ( .B(n630), .A(n629), .Z(n633) );
  NANDN U775 ( .A(y[2038]), .B(x[2038]), .Z(n632) );
  NANDN U776 ( .A(y[2037]), .B(x[2037]), .Z(n631) );
  NAND U777 ( .A(n632), .B(n631), .Z(n14053) );
  ANDN U778 ( .B(n633), .A(n14053), .Z(n640) );
  ANDN U779 ( .B(x[2047]), .A(y[2047]), .Z(n14074) );
  ANDN U780 ( .B(x[2042]), .A(y[2042]), .Z(n14062) );
  NOR U781 ( .A(n14074), .B(n14062), .Z(n635) );
  NANDN U782 ( .A(y[2036]), .B(x[2036]), .Z(n643) );
  NANDN U783 ( .A(x[2037]), .B(y[2037]), .Z(n642) );
  NANDN U784 ( .A(n643), .B(n642), .Z(n634) );
  AND U785 ( .A(n635), .B(n634), .Z(n638) );
  NANDN U786 ( .A(y[2046]), .B(x[2046]), .Z(n637) );
  NANDN U787 ( .A(y[2045]), .B(x[2045]), .Z(n636) );
  NAND U788 ( .A(n637), .B(n636), .Z(n14068) );
  ANDN U789 ( .B(n638), .A(n14068), .Z(n639) );
  AND U790 ( .A(n640), .B(n639), .Z(n647) );
  NANDN U791 ( .A(x[2036]), .B(y[2036]), .Z(n641) );
  NAND U792 ( .A(n642), .B(n641), .Z(n9962) );
  ANDN U793 ( .B(x[2035]), .A(y[2035]), .Z(n658) );
  ANDN U794 ( .B(y[2035]), .A(x[2035]), .Z(n9964) );
  NANDN U795 ( .A(x[2034]), .B(y[2034]), .Z(n9956) );
  NANDN U796 ( .A(n9964), .B(n9956), .Z(n644) );
  IV U797 ( .A(n643), .Z(n660) );
  ANDN U798 ( .B(n644), .A(n660), .Z(n645) );
  NANDN U799 ( .A(n658), .B(n645), .Z(n646) );
  NANDN U800 ( .A(n9962), .B(n646), .Z(n14051) );
  ANDN U801 ( .B(n647), .A(n14051), .Z(n656) );
  NANDN U802 ( .A(x[2043]), .B(y[2043]), .Z(n649) );
  NANDN U803 ( .A(x[2042]), .B(y[2042]), .Z(n648) );
  AND U804 ( .A(n649), .B(n648), .Z(n652) );
  NANDN U805 ( .A(x[2045]), .B(y[2045]), .Z(n651) );
  NANDN U806 ( .A(x[2044]), .B(y[2044]), .Z(n650) );
  AND U807 ( .A(n651), .B(n650), .Z(n14066) );
  NAND U808 ( .A(n652), .B(n14066), .Z(n14065) );
  XNOR U809 ( .A(y[2040]), .B(x[2040]), .Z(n654) );
  NANDN U810 ( .A(x[2039]), .B(y[2039]), .Z(n653) );
  NAND U811 ( .A(n654), .B(n653), .Z(n14057) );
  NOR U812 ( .A(n14065), .B(n14057), .Z(n655) );
  AND U813 ( .A(n656), .B(n655), .Z(n9969) );
  NANDN U814 ( .A(y[2034]), .B(x[2034]), .Z(n657) );
  NANDN U815 ( .A(n658), .B(n657), .Z(n9961) );
  ANDN U816 ( .B(x[2033]), .A(y[2033]), .Z(n9955) );
  NOR U817 ( .A(n9961), .B(n9955), .Z(n659) );
  NANDN U818 ( .A(n660), .B(n659), .Z(n14048) );
  NANDN U819 ( .A(x[2030]), .B(y[2030]), .Z(n662) );
  NANDN U820 ( .A(x[2031]), .B(y[2031]), .Z(n661) );
  NAND U821 ( .A(n662), .B(n661), .Z(n14043) );
  NANDN U822 ( .A(x[2029]), .B(y[2029]), .Z(n14036) );
  NANDN U823 ( .A(x[2028]), .B(y[2028]), .Z(n14037) );
  NANDN U824 ( .A(y[2027]), .B(x[2027]), .Z(n6092) );
  ANDN U825 ( .B(n14037), .A(n6092), .Z(n6084) );
  NANDN U826 ( .A(x[2026]), .B(y[2026]), .Z(n14028) );
  ANDN U827 ( .B(y[2027]), .A(x[2027]), .Z(n14033) );
  XNOR U828 ( .A(x[2028]), .B(y[2028]), .Z(n663) );
  NANDN U829 ( .A(n14033), .B(n663), .Z(n9939) );
  ANDN U830 ( .B(n14028), .A(n9939), .Z(n6081) );
  NANDN U831 ( .A(y[2026]), .B(x[2026]), .Z(n6093) );
  NANDN U832 ( .A(y[2025]), .B(x[2025]), .Z(n14027) );
  NAND U833 ( .A(n6093), .B(n14027), .Z(n6079) );
  NANDN U834 ( .A(y[2023]), .B(x[2023]), .Z(n9927) );
  NANDN U835 ( .A(y[2024]), .B(x[2024]), .Z(n664) );
  NAND U836 ( .A(n9927), .B(n664), .Z(n14022) );
  NANDN U837 ( .A(x[2021]), .B(y[2021]), .Z(n14016) );
  NANDN U838 ( .A(x[2020]), .B(y[2020]), .Z(n6094) );
  AND U839 ( .A(n14016), .B(n6094), .Z(n6070) );
  NANDN U840 ( .A(y[2019]), .B(x[2019]), .Z(n666) );
  NANDN U841 ( .A(y[2018]), .B(x[2018]), .Z(n665) );
  NAND U842 ( .A(n666), .B(n665), .Z(n14011) );
  NANDN U843 ( .A(y[2017]), .B(x[2017]), .Z(n672) );
  ANDN U844 ( .B(x[2015]), .A(y[2015]), .Z(n667) );
  OR U845 ( .A(n667), .B(x[2016]), .Z(n670) );
  XOR U846 ( .A(x[2016]), .B(n667), .Z(n668) );
  NAND U847 ( .A(n668), .B(y[2016]), .Z(n669) );
  NAND U848 ( .A(n670), .B(n669), .Z(n671) );
  NAND U849 ( .A(n672), .B(n671), .Z(n14007) );
  NANDN U850 ( .A(x[2015]), .B(y[2015]), .Z(n674) );
  NANDN U851 ( .A(x[2014]), .B(y[2014]), .Z(n673) );
  AND U852 ( .A(n674), .B(n673), .Z(n676) );
  NANDN U853 ( .A(x[2016]), .B(y[2016]), .Z(n675) );
  NAND U854 ( .A(n676), .B(n675), .Z(n14005) );
  NANDN U855 ( .A(y[2011]), .B(x[2011]), .Z(n678) );
  NANDN U856 ( .A(y[2012]), .B(x[2012]), .Z(n677) );
  AND U857 ( .A(n678), .B(n677), .Z(n13998) );
  NANDN U858 ( .A(y[2010]), .B(x[2010]), .Z(n679) );
  ANDN U859 ( .B(x[2009]), .A(y[2009]), .Z(n9906) );
  ANDN U860 ( .B(n679), .A(n9906), .Z(n13994) );
  NANDN U861 ( .A(y[2007]), .B(x[2007]), .Z(n681) );
  NANDN U862 ( .A(y[2008]), .B(x[2008]), .Z(n680) );
  AND U863 ( .A(n681), .B(n680), .Z(n13990) );
  NANDN U864 ( .A(y[2005]), .B(x[2005]), .Z(n683) );
  NANDN U865 ( .A(y[2006]), .B(x[2006]), .Z(n682) );
  AND U866 ( .A(n683), .B(n682), .Z(n13986) );
  NANDN U867 ( .A(x[2004]), .B(y[2004]), .Z(n685) );
  NANDN U868 ( .A(x[2005]), .B(y[2005]), .Z(n684) );
  NAND U869 ( .A(n685), .B(n684), .Z(n13984) );
  NANDN U870 ( .A(y[2004]), .B(x[2004]), .Z(n687) );
  NANDN U871 ( .A(y[2003]), .B(x[2003]), .Z(n686) );
  NAND U872 ( .A(n687), .B(n686), .Z(n13983) );
  NANDN U873 ( .A(y[2001]), .B(x[2001]), .Z(n6096) );
  NANDN U874 ( .A(y[2002]), .B(x[2002]), .Z(n688) );
  NAND U875 ( .A(n6096), .B(n688), .Z(n6037) );
  ANDN U876 ( .B(x[1999]), .A(y[1999]), .Z(n6105) );
  NANDN U877 ( .A(y[2000]), .B(x[2000]), .Z(n6099) );
  NANDN U878 ( .A(x[1998]), .B(y[1998]), .Z(n13973) );
  NANDN U879 ( .A(y[1997]), .B(x[1997]), .Z(n13972) );
  ANDN U880 ( .B(x[1998]), .A(y[1998]), .Z(n6104) );
  ANDN U881 ( .B(n13972), .A(n6104), .Z(n6029) );
  NANDN U882 ( .A(x[1997]), .B(y[1997]), .Z(n9894) );
  NANDN U883 ( .A(x[1996]), .B(y[1996]), .Z(n9888) );
  NAND U884 ( .A(n9894), .B(n9888), .Z(n13971) );
  NANDN U885 ( .A(y[1996]), .B(x[1996]), .Z(n9891) );
  NANDN U886 ( .A(y[1995]), .B(x[1995]), .Z(n6107) );
  NAND U887 ( .A(n9891), .B(n6107), .Z(n13970) );
  NANDN U888 ( .A(x[1994]), .B(y[1994]), .Z(n689) );
  NANDN U889 ( .A(x[1995]), .B(y[1995]), .Z(n9886) );
  NAND U890 ( .A(n689), .B(n9886), .Z(n13969) );
  NANDN U891 ( .A(x[1993]), .B(y[1993]), .Z(n13967) );
  NANDN U892 ( .A(x[1992]), .B(y[1992]), .Z(n6110) );
  AND U893 ( .A(n13967), .B(n6110), .Z(n6022) );
  NANDN U894 ( .A(x[1991]), .B(y[1991]), .Z(n6111) );
  NANDN U895 ( .A(x[1990]), .B(y[1990]), .Z(n13963) );
  XNOR U896 ( .A(y[1987]), .B(x[1987]), .Z(n13960) );
  NANDN U897 ( .A(x[1985]), .B(y[1985]), .Z(n691) );
  NANDN U898 ( .A(x[1986]), .B(y[1986]), .Z(n690) );
  NAND U899 ( .A(n691), .B(n690), .Z(n13958) );
  ANDN U900 ( .B(x[1985]), .A(y[1985]), .Z(n9865) );
  NANDN U901 ( .A(x[1984]), .B(y[1984]), .Z(n13954) );
  NANDN U902 ( .A(y[1981]), .B(x[1981]), .Z(n692) );
  NANDN U903 ( .A(y[1982]), .B(x[1982]), .Z(n9859) );
  NAND U904 ( .A(n692), .B(n9859), .Z(n13949) );
  XOR U905 ( .A(x[1980]), .B(y[1980]), .Z(n9847) );
  NANDN U906 ( .A(y[1979]), .B(x[1979]), .Z(n694) );
  NANDN U907 ( .A(y[1978]), .B(x[1978]), .Z(n693) );
  AND U908 ( .A(n694), .B(n693), .Z(n9845) );
  NANDN U909 ( .A(x[1979]), .B(y[1979]), .Z(n5995) );
  IV U910 ( .A(n5995), .Z(n9849) );
  OR U911 ( .A(n9845), .B(n9849), .Z(n695) );
  NANDN U912 ( .A(n9847), .B(n695), .Z(n13944) );
  NANDN U913 ( .A(y[1976]), .B(x[1976]), .Z(n697) );
  NANDN U914 ( .A(y[1977]), .B(x[1977]), .Z(n696) );
  AND U915 ( .A(n697), .B(n696), .Z(n13941) );
  NANDN U916 ( .A(y[1975]), .B(x[1975]), .Z(n698) );
  ANDN U917 ( .B(x[1974]), .A(y[1974]), .Z(n13934) );
  ANDN U918 ( .B(n698), .A(n13934), .Z(n9838) );
  NANDN U919 ( .A(x[1974]), .B(y[1974]), .Z(n700) );
  NANDN U920 ( .A(x[1973]), .B(y[1973]), .Z(n699) );
  NAND U921 ( .A(n700), .B(n699), .Z(n13933) );
  NANDN U922 ( .A(y[1971]), .B(x[1971]), .Z(n5984) );
  IV U923 ( .A(x[1971]), .Z(n9829) );
  IV U924 ( .A(y[1971]), .Z(n9828) );
  XNOR U925 ( .A(n9829), .B(n9828), .Z(n5982) );
  NANDN U926 ( .A(x[1970]), .B(y[1970]), .Z(n13924) );
  NANDN U927 ( .A(y[1968]), .B(x[1968]), .Z(n702) );
  NANDN U928 ( .A(y[1967]), .B(x[1967]), .Z(n701) );
  NAND U929 ( .A(n702), .B(n701), .Z(n13919) );
  NANDN U930 ( .A(y[1966]), .B(x[1966]), .Z(n704) );
  NANDN U931 ( .A(y[1965]), .B(x[1965]), .Z(n703) );
  NAND U932 ( .A(n704), .B(n703), .Z(n13917) );
  NANDN U933 ( .A(y[1962]), .B(x[1962]), .Z(n706) );
  NANDN U934 ( .A(y[1961]), .B(x[1961]), .Z(n705) );
  NAND U935 ( .A(n706), .B(n705), .Z(n13913) );
  ANDN U936 ( .B(y[1961]), .A(x[1961]), .Z(n5958) );
  ANDN U937 ( .B(x[1960]), .A(y[1960]), .Z(n13910) );
  NANDN U938 ( .A(n5958), .B(n13910), .Z(n707) );
  NANDN U939 ( .A(n13913), .B(n707), .Z(n9818) );
  NANDN U940 ( .A(y[1957]), .B(x[1957]), .Z(n5952) );
  XNOR U941 ( .A(y[1957]), .B(x[1957]), .Z(n709) );
  NANDN U942 ( .A(x[1956]), .B(y[1956]), .Z(n708) );
  NAND U943 ( .A(n709), .B(n708), .Z(n710) );
  AND U944 ( .A(n5952), .B(n710), .Z(n13906) );
  ANDN U945 ( .B(y[1958]), .A(x[1958]), .Z(n13909) );
  OR U946 ( .A(n13906), .B(n13909), .Z(n9812) );
  NANDN U947 ( .A(x[1955]), .B(y[1955]), .Z(n9809) );
  NANDN U948 ( .A(y[1954]), .B(x[1954]), .Z(n711) );
  NANDN U949 ( .A(y[1953]), .B(x[1953]), .Z(n9802) );
  NAND U950 ( .A(n711), .B(n9802), .Z(n13903) );
  NANDN U951 ( .A(y[1951]), .B(x[1951]), .Z(n9796) );
  XOR U952 ( .A(x[1952]), .B(y[1952]), .Z(n9800) );
  ANDN U953 ( .B(n9796), .A(n9800), .Z(n13900) );
  NANDN U954 ( .A(x[1951]), .B(y[1951]), .Z(n13893) );
  NANDN U955 ( .A(y[1950]), .B(x[1950]), .Z(n713) );
  NANDN U956 ( .A(y[1949]), .B(x[1949]), .Z(n712) );
  NAND U957 ( .A(n713), .B(n712), .Z(n13891) );
  NANDN U958 ( .A(x[1949]), .B(y[1949]), .Z(n13894) );
  NANDN U959 ( .A(y[1943]), .B(x[1943]), .Z(n715) );
  NANDN U960 ( .A(y[1944]), .B(x[1944]), .Z(n714) );
  AND U961 ( .A(n715), .B(n714), .Z(n13878) );
  NANDN U962 ( .A(y[1939]), .B(x[1939]), .Z(n9780) );
  ANDN U963 ( .B(x[1940]), .A(y[1940]), .Z(n9783) );
  ANDN U964 ( .B(n9780), .A(n9783), .Z(n13870) );
  NANDN U965 ( .A(y[1937]), .B(x[1937]), .Z(n717) );
  NANDN U966 ( .A(y[1938]), .B(x[1938]), .Z(n716) );
  AND U967 ( .A(n717), .B(n716), .Z(n13866) );
  ANDN U968 ( .B(x[1930]), .A(y[1930]), .Z(n13851) );
  ANDN U969 ( .B(x[1929]), .A(y[1929]), .Z(n9765) );
  NOR U970 ( .A(n13851), .B(n9765), .Z(n5892) );
  ANDN U971 ( .B(y[1929]), .A(x[1929]), .Z(n13848) );
  NANDN U972 ( .A(x[1928]), .B(y[1928]), .Z(n13844) );
  NANDN U973 ( .A(n13848), .B(n13844), .Z(n5890) );
  ANDN U974 ( .B(x[1928]), .A(y[1928]), .Z(n9764) );
  NANDN U975 ( .A(y[1927]), .B(x[1927]), .Z(n13842) );
  NANDN U976 ( .A(y[1924]), .B(x[1924]), .Z(n719) );
  NANDN U977 ( .A(y[1925]), .B(x[1925]), .Z(n718) );
  NAND U978 ( .A(n719), .B(n718), .Z(n13835) );
  NANDN U979 ( .A(y[1923]), .B(x[1923]), .Z(n9755) );
  NANDN U980 ( .A(y[1921]), .B(x[1921]), .Z(n6112) );
  NANDN U981 ( .A(y[1920]), .B(x[1920]), .Z(n5868) );
  NANDN U982 ( .A(y[1919]), .B(x[1919]), .Z(n720) );
  NAND U983 ( .A(n5868), .B(n720), .Z(n13823) );
  NANDN U984 ( .A(x[1918]), .B(y[1918]), .Z(n9982) );
  ANDN U985 ( .B(y[1915]), .A(x[1915]), .Z(n9733) );
  NANDN U986 ( .A(x[1914]), .B(y[1914]), .Z(n721) );
  NANDN U987 ( .A(n9733), .B(n721), .Z(n13818) );
  ANDN U988 ( .B(x[1913]), .A(y[1913]), .Z(n13817) );
  NANDN U989 ( .A(y[1914]), .B(x[1914]), .Z(n9732) );
  NANDN U990 ( .A(n13817), .B(n9732), .Z(n5859) );
  NANDN U991 ( .A(x[1913]), .B(y[1913]), .Z(n723) );
  NANDN U992 ( .A(x[1912]), .B(y[1912]), .Z(n722) );
  AND U993 ( .A(n723), .B(n722), .Z(n13816) );
  NANDN U994 ( .A(y[1912]), .B(x[1912]), .Z(n725) );
  NANDN U995 ( .A(y[1911]), .B(x[1911]), .Z(n724) );
  NAND U996 ( .A(n725), .B(n724), .Z(n13815) );
  NANDN U997 ( .A(x[1905]), .B(y[1905]), .Z(n6116) );
  NANDN U998 ( .A(x[1904]), .B(y[1904]), .Z(n726) );
  NAND U999 ( .A(n6116), .B(n726), .Z(n6121) );
  NANDN U1000 ( .A(y[1904]), .B(x[1904]), .Z(n6117) );
  NANDN U1001 ( .A(y[1903]), .B(x[1903]), .Z(n6122) );
  AND U1002 ( .A(n6117), .B(n6122), .Z(n5836) );
  NANDN U1003 ( .A(x[1903]), .B(y[1903]), .Z(n6120) );
  ANDN U1004 ( .B(x[1901]), .A(y[1901]), .Z(n6127) );
  NANDN U1005 ( .A(y[1902]), .B(x[1902]), .Z(n6123) );
  NANDN U1006 ( .A(y[1899]), .B(x[1899]), .Z(n13798) );
  ANDN U1007 ( .B(x[1900]), .A(y[1900]), .Z(n6126) );
  ANDN U1008 ( .B(n13798), .A(n6126), .Z(n5828) );
  NANDN U1009 ( .A(y[1898]), .B(x[1898]), .Z(n728) );
  NANDN U1010 ( .A(y[1897]), .B(x[1897]), .Z(n727) );
  NAND U1011 ( .A(n728), .B(n727), .Z(n13795) );
  NANDN U1012 ( .A(y[1894]), .B(x[1894]), .Z(n6128) );
  NANDN U1013 ( .A(y[1893]), .B(x[1893]), .Z(n729) );
  NAND U1014 ( .A(n6128), .B(n729), .Z(n13786) );
  NANDN U1015 ( .A(y[1891]), .B(x[1891]), .Z(n730) );
  NANDN U1016 ( .A(y[1892]), .B(x[1892]), .Z(n9709) );
  NAND U1017 ( .A(n730), .B(n9709), .Z(n13782) );
  NANDN U1018 ( .A(x[1891]), .B(y[1891]), .Z(n6132) );
  NANDN U1019 ( .A(x[1890]), .B(y[1890]), .Z(n9700) );
  NAND U1020 ( .A(n6132), .B(n9700), .Z(n13781) );
  ANDN U1021 ( .B(x[1890]), .A(y[1890]), .Z(n13779) );
  ANDN U1022 ( .B(x[1889]), .A(y[1889]), .Z(n9697) );
  NOR U1023 ( .A(n13779), .B(n9697), .Z(n5808) );
  ANDN U1024 ( .B(x[1880]), .A(y[1880]), .Z(n9983) );
  ANDN U1025 ( .B(x[1879]), .A(y[1879]), .Z(n13754) );
  OR U1026 ( .A(n9983), .B(n13754), .Z(n9680) );
  ANDN U1027 ( .B(y[1879]), .A(x[1879]), .Z(n6133) );
  NANDN U1028 ( .A(x[1878]), .B(y[1878]), .Z(n13752) );
  NANDN U1029 ( .A(n6133), .B(n13752), .Z(n5783) );
  IV U1030 ( .A(y[1877]), .Z(n6137) );
  IV U1031 ( .A(x[1877]), .Z(n6136) );
  NANDN U1032 ( .A(n6137), .B(n6136), .Z(n731) );
  IV U1033 ( .A(y[1876]), .Z(n6138) );
  NAND U1034 ( .A(n731), .B(n9675), .Z(n13749) );
  NANDN U1035 ( .A(y[1876]), .B(x[1876]), .Z(n732) );
  NANDN U1036 ( .A(y[1875]), .B(x[1875]), .Z(n6139) );
  NAND U1037 ( .A(n732), .B(n6139), .Z(n13747) );
  NANDN U1038 ( .A(x[1875]), .B(y[1875]), .Z(n13745) );
  NANDN U1039 ( .A(y[1873]), .B(x[1873]), .Z(n734) );
  NANDN U1040 ( .A(y[1872]), .B(x[1872]), .Z(n733) );
  NAND U1041 ( .A(n734), .B(n733), .Z(n13739) );
  NANDN U1042 ( .A(y[1871]), .B(x[1871]), .Z(n5769) );
  ANDN U1043 ( .B(y[1870]), .A(x[1870]), .Z(n6140) );
  NAND U1044 ( .A(n5769), .B(n6140), .Z(n737) );
  NANDN U1045 ( .A(x[1871]), .B(y[1871]), .Z(n736) );
  NANDN U1046 ( .A(x[1872]), .B(y[1872]), .Z(n735) );
  AND U1047 ( .A(n736), .B(n735), .Z(n9665) );
  NAND U1048 ( .A(n737), .B(n9665), .Z(n13737) );
  NANDN U1049 ( .A(x[1869]), .B(y[1869]), .Z(n9985) );
  NANDN U1050 ( .A(y[1867]), .B(x[1867]), .Z(n13730) );
  NANDN U1051 ( .A(x[1865]), .B(y[1865]), .Z(n739) );
  NANDN U1052 ( .A(x[1864]), .B(y[1864]), .Z(n738) );
  NAND U1053 ( .A(n739), .B(n738), .Z(n13722) );
  ANDN U1054 ( .B(y[1858]), .A(x[1858]), .Z(n13707) );
  NANDN U1055 ( .A(x[1856]), .B(y[1856]), .Z(n741) );
  NANDN U1056 ( .A(x[1857]), .B(y[1857]), .Z(n740) );
  NAND U1057 ( .A(n741), .B(n740), .Z(n13703) );
  NANDN U1058 ( .A(y[1854]), .B(x[1854]), .Z(n9638) );
  NANDN U1059 ( .A(y[1853]), .B(x[1853]), .Z(n9630) );
  NAND U1060 ( .A(n9638), .B(n9630), .Z(n13697) );
  NANDN U1061 ( .A(y[1852]), .B(x[1852]), .Z(n9631) );
  NANDN U1062 ( .A(y[1851]), .B(x[1851]), .Z(n9623) );
  AND U1063 ( .A(n9631), .B(n9623), .Z(n13693) );
  NANDN U1064 ( .A(x[1850]), .B(y[1850]), .Z(n13689) );
  NANDN U1065 ( .A(y[1850]), .B(x[1850]), .Z(n9621) );
  NANDN U1066 ( .A(y[1849]), .B(x[1849]), .Z(n9616) );
  NAND U1067 ( .A(n9621), .B(n9616), .Z(n13687) );
  IV U1068 ( .A(x[1846]), .Z(n9987) );
  OR U1069 ( .A(y[1846]), .B(n9987), .Z(n742) );
  ANDN U1070 ( .B(x[1847]), .A(y[1847]), .Z(n13680) );
  ANDN U1071 ( .B(n742), .A(n13680), .Z(n9610) );
  ANDN U1072 ( .B(y[1845]), .A(x[1845]), .Z(n13673) );
  NANDN U1073 ( .A(x[1846]), .B(y[1846]), .Z(n13677) );
  NANDN U1074 ( .A(n13673), .B(n13677), .Z(n9609) );
  ANDN U1075 ( .B(x[1845]), .A(y[1845]), .Z(n9605) );
  ANDN U1076 ( .B(y[1843]), .A(x[1843]), .Z(n9604) );
  ANDN U1077 ( .B(y[1842]), .A(x[1842]), .Z(n9599) );
  NOR U1078 ( .A(n9604), .B(n9599), .Z(n13664) );
  NANDN U1079 ( .A(x[1841]), .B(y[1841]), .Z(n9988) );
  NANDN U1080 ( .A(x[1839]), .B(y[1839]), .Z(n9592) );
  NANDN U1081 ( .A(x[1838]), .B(y[1838]), .Z(n6147) );
  NAND U1082 ( .A(n9592), .B(n6147), .Z(n13653) );
  NANDN U1083 ( .A(x[1836]), .B(y[1836]), .Z(n6151) );
  IV U1084 ( .A(y[1837]), .Z(n6149) );
  IV U1085 ( .A(x[1837]), .Z(n6148) );
  NANDN U1086 ( .A(n6149), .B(n6148), .Z(n743) );
  NAND U1087 ( .A(n6151), .B(n743), .Z(n13649) );
  NANDN U1088 ( .A(x[1835]), .B(y[1835]), .Z(n6150) );
  NANDN U1089 ( .A(x[1834]), .B(y[1834]), .Z(n9575) );
  NAND U1090 ( .A(n6150), .B(n9575), .Z(n13644) );
  NANDN U1091 ( .A(x[1833]), .B(y[1833]), .Z(n13640) );
  ANDN U1092 ( .B(y[1832]), .A(x[1832]), .Z(n9568) );
  ANDN U1093 ( .B(n13640), .A(n9568), .Z(n5700) );
  XNOR U1094 ( .A(y[1831]), .B(x[1831]), .Z(n5696) );
  ANDN U1095 ( .B(x[1829]), .A(y[1829]), .Z(n13631) );
  ANDN U1096 ( .B(x[1830]), .A(y[1830]), .Z(n9565) );
  NOR U1097 ( .A(n13631), .B(n9565), .Z(n5693) );
  NANDN U1098 ( .A(x[1828]), .B(y[1828]), .Z(n745) );
  NANDN U1099 ( .A(x[1829]), .B(y[1829]), .Z(n744) );
  NAND U1100 ( .A(n745), .B(n744), .Z(n13629) );
  NANDN U1101 ( .A(y[1828]), .B(x[1828]), .Z(n747) );
  NANDN U1102 ( .A(y[1827]), .B(x[1827]), .Z(n746) );
  NAND U1103 ( .A(n747), .B(n746), .Z(n13627) );
  ANDN U1104 ( .B(y[1827]), .A(x[1827]), .Z(n5687) );
  ANDN U1105 ( .B(x[1826]), .A(y[1826]), .Z(n13621) );
  NANDN U1106 ( .A(n5687), .B(n13621), .Z(n748) );
  NANDN U1107 ( .A(n13627), .B(n748), .Z(n9561) );
  NANDN U1108 ( .A(y[1825]), .B(x[1825]), .Z(n13622) );
  NANDN U1109 ( .A(y[1824]), .B(x[1824]), .Z(n13617) );
  NANDN U1110 ( .A(y[1823]), .B(x[1823]), .Z(n9549) );
  AND U1111 ( .A(n13617), .B(n9549), .Z(n5684) );
  NANDN U1112 ( .A(x[1822]), .B(y[1822]), .Z(n13610) );
  NANDN U1113 ( .A(y[1821]), .B(x[1821]), .Z(n749) );
  XNOR U1114 ( .A(x[1822]), .B(y[1822]), .Z(n9543) );
  NAND U1115 ( .A(n749), .B(n9543), .Z(n13609) );
  NANDN U1116 ( .A(x[1820]), .B(y[1820]), .Z(n751) );
  NANDN U1117 ( .A(x[1821]), .B(y[1821]), .Z(n750) );
  NAND U1118 ( .A(n751), .B(n750), .Z(n13607) );
  IV U1119 ( .A(x[1820]), .Z(n9537) );
  OR U1120 ( .A(y[1820]), .B(n9537), .Z(n752) );
  NANDN U1121 ( .A(y[1819]), .B(x[1819]), .Z(n9534) );
  NAND U1122 ( .A(n752), .B(n9534), .Z(n13605) );
  NANDN U1123 ( .A(y[1815]), .B(x[1815]), .Z(n13592) );
  IV U1124 ( .A(x[1814]), .Z(n6154) );
  IV U1125 ( .A(y[1814]), .Z(n6153) );
  NANDN U1126 ( .A(n6154), .B(n6153), .Z(n753) );
  IV U1127 ( .A(x[1813]), .Z(n6155) );
  NAND U1128 ( .A(n753), .B(n9521), .Z(n13589) );
  NANDN U1129 ( .A(x[1813]), .B(y[1813]), .Z(n755) );
  IV U1130 ( .A(y[1812]), .Z(n6157) );
  IV U1131 ( .A(x[1812]), .Z(n6156) );
  NANDN U1132 ( .A(n6157), .B(n6156), .Z(n754) );
  NAND U1133 ( .A(n755), .B(n754), .Z(n13587) );
  NANDN U1134 ( .A(y[1812]), .B(x[1812]), .Z(n756) );
  NANDN U1135 ( .A(y[1811]), .B(x[1811]), .Z(n9511) );
  NAND U1136 ( .A(n756), .B(n9511), .Z(n13584) );
  NANDN U1137 ( .A(y[1809]), .B(x[1809]), .Z(n13576) );
  ANDN U1138 ( .B(x[1810]), .A(y[1810]), .Z(n13581) );
  ANDN U1139 ( .B(n13576), .A(n13581), .Z(n5661) );
  NANDN U1140 ( .A(x[1808]), .B(y[1808]), .Z(n13574) );
  NANDN U1141 ( .A(y[1807]), .B(x[1807]), .Z(n757) );
  NANDN U1142 ( .A(y[1808]), .B(x[1808]), .Z(n9506) );
  NAND U1143 ( .A(n757), .B(n9506), .Z(n13572) );
  NANDN U1144 ( .A(x[1806]), .B(y[1806]), .Z(n6162) );
  NANDN U1145 ( .A(x[1807]), .B(y[1807]), .Z(n6160) );
  NAND U1146 ( .A(n6162), .B(n6160), .Z(n13571) );
  NANDN U1147 ( .A(y[1805]), .B(x[1805]), .Z(n758) );
  NANDN U1148 ( .A(y[1806]), .B(x[1806]), .Z(n9501) );
  NAND U1149 ( .A(n758), .B(n9501), .Z(n13570) );
  NANDN U1150 ( .A(x[1804]), .B(y[1804]), .Z(n9492) );
  IV U1151 ( .A(y[1805]), .Z(n6164) );
  IV U1152 ( .A(x[1805]), .Z(n6163) );
  NANDN U1153 ( .A(n6164), .B(n6163), .Z(n759) );
  NAND U1154 ( .A(n9492), .B(n759), .Z(n13569) );
  NANDN U1155 ( .A(y[1804]), .B(x[1804]), .Z(n13568) );
  NANDN U1156 ( .A(y[1803]), .B(x[1803]), .Z(n9489) );
  AND U1157 ( .A(n13568), .B(n9489), .Z(n5653) );
  NANDN U1158 ( .A(y[1801]), .B(x[1801]), .Z(n13564) );
  NANDN U1159 ( .A(y[1802]), .B(x[1802]), .Z(n9490) );
  AND U1160 ( .A(n13564), .B(n9490), .Z(n5649) );
  NANDN U1161 ( .A(y[1798]), .B(x[1798]), .Z(n760) );
  NANDN U1162 ( .A(y[1799]), .B(x[1799]), .Z(n9990) );
  AND U1163 ( .A(n760), .B(n9990), .Z(n9479) );
  NANDN U1164 ( .A(y[1797]), .B(x[1797]), .Z(n5639) );
  ANDN U1165 ( .B(x[1795]), .A(y[1795]), .Z(n13556) );
  NOR U1166 ( .A(n13560), .B(n13556), .Z(n9475) );
  NANDN U1167 ( .A(x[1794]), .B(y[1794]), .Z(n762) );
  NANDN U1168 ( .A(x[1795]), .B(y[1795]), .Z(n761) );
  NAND U1169 ( .A(n762), .B(n761), .Z(n13555) );
  NANDN U1170 ( .A(x[1792]), .B(y[1792]), .Z(n764) );
  NANDN U1171 ( .A(x[1793]), .B(y[1793]), .Z(n763) );
  NAND U1172 ( .A(n764), .B(n763), .Z(n6168) );
  NANDN U1173 ( .A(x[1791]), .B(y[1791]), .Z(n6165) );
  ANDN U1174 ( .B(y[1788]), .A(x[1788]), .Z(n13543) );
  NANDN U1175 ( .A(y[1787]), .B(x[1787]), .Z(n13541) );
  ANDN U1176 ( .B(x[1788]), .A(y[1788]), .Z(n9466) );
  ANDN U1177 ( .B(n13541), .A(n9466), .Z(n5619) );
  NANDN U1178 ( .A(x[1787]), .B(y[1787]), .Z(n766) );
  NANDN U1179 ( .A(x[1786]), .B(y[1786]), .Z(n765) );
  NAND U1180 ( .A(n766), .B(n765), .Z(n13539) );
  NANDN U1181 ( .A(y[1786]), .B(x[1786]), .Z(n9457) );
  NANDN U1182 ( .A(y[1785]), .B(x[1785]), .Z(n767) );
  NAND U1183 ( .A(n9457), .B(n767), .Z(n13537) );
  NANDN U1184 ( .A(x[1785]), .B(y[1785]), .Z(n769) );
  NANDN U1185 ( .A(x[1784]), .B(y[1784]), .Z(n768) );
  NAND U1186 ( .A(n769), .B(n768), .Z(n13535) );
  ANDN U1187 ( .B(y[1782]), .A(x[1782]), .Z(n6172) );
  ANDN U1188 ( .B(y[1783]), .A(x[1783]), .Z(n13531) );
  OR U1189 ( .A(n6172), .B(n13531), .Z(n5612) );
  ANDN U1190 ( .B(x[1782]), .A(y[1782]), .Z(n13528) );
  NANDN U1191 ( .A(y[1781]), .B(x[1781]), .Z(n13524) );
  NANDN U1192 ( .A(n13528), .B(n13524), .Z(n5610) );
  NANDN U1193 ( .A(y[1780]), .B(x[1780]), .Z(n771) );
  NANDN U1194 ( .A(y[1779]), .B(x[1779]), .Z(n770) );
  NAND U1195 ( .A(n771), .B(n770), .Z(n13521) );
  NANDN U1196 ( .A(x[1778]), .B(y[1778]), .Z(n773) );
  NANDN U1197 ( .A(x[1779]), .B(y[1779]), .Z(n772) );
  AND U1198 ( .A(n773), .B(n772), .Z(n13518) );
  NANDN U1199 ( .A(y[1772]), .B(x[1772]), .Z(n6173) );
  NANDN U1200 ( .A(y[1771]), .B(x[1771]), .Z(n6175) );
  NAND U1201 ( .A(n6173), .B(n6175), .Z(n13508) );
  NANDN U1202 ( .A(x[1770]), .B(y[1770]), .Z(n774) );
  ANDN U1203 ( .B(y[1771]), .A(x[1771]), .Z(n9418) );
  ANDN U1204 ( .B(n774), .A(n9418), .Z(n13506) );
  NANDN U1205 ( .A(y[1769]), .B(x[1769]), .Z(n6179) );
  IV U1206 ( .A(x[1770]), .Z(n6177) );
  IV U1207 ( .A(y[1770]), .Z(n6176) );
  NANDN U1208 ( .A(n6177), .B(n6176), .Z(n775) );
  NAND U1209 ( .A(n6179), .B(n775), .Z(n13505) );
  NANDN U1210 ( .A(y[1767]), .B(x[1767]), .Z(n9401) );
  IV U1211 ( .A(x[1768]), .Z(n6181) );
  IV U1212 ( .A(y[1768]), .Z(n6180) );
  NANDN U1213 ( .A(n6181), .B(n6180), .Z(n776) );
  NAND U1214 ( .A(n9401), .B(n776), .Z(n13501) );
  NANDN U1215 ( .A(y[1765]), .B(x[1765]), .Z(n778) );
  NANDN U1216 ( .A(y[1766]), .B(x[1766]), .Z(n777) );
  NAND U1217 ( .A(n778), .B(n777), .Z(n13496) );
  IV U1218 ( .A(y[1765]), .Z(n9395) );
  OR U1219 ( .A(x[1765]), .B(n9395), .Z(n779) );
  ANDN U1220 ( .B(y[1764]), .A(x[1764]), .Z(n6182) );
  ANDN U1221 ( .B(n779), .A(n6182), .Z(n13494) );
  NANDN U1222 ( .A(y[1762]), .B(x[1762]), .Z(n13488) );
  ANDN U1223 ( .B(x[1761]), .A(y[1761]), .Z(n6187) );
  ANDN U1224 ( .B(n13488), .A(n6187), .Z(n5577) );
  NANDN U1225 ( .A(x[1761]), .B(y[1761]), .Z(n6185) );
  NANDN U1226 ( .A(y[1757]), .B(x[1757]), .Z(n780) );
  ANDN U1227 ( .B(x[1758]), .A(y[1758]), .Z(n9383) );
  ANDN U1228 ( .B(n780), .A(n9383), .Z(n13476) );
  NANDN U1229 ( .A(y[1753]), .B(x[1753]), .Z(n9367) );
  IV U1230 ( .A(n9367), .Z(n13465) );
  ANDN U1231 ( .B(x[1752]), .A(y[1752]), .Z(n9366) );
  NANDN U1232 ( .A(y[1751]), .B(x[1751]), .Z(n13459) );
  NANDN U1233 ( .A(x[1749]), .B(y[1749]), .Z(n13451) );
  NANDN U1234 ( .A(x[1748]), .B(y[1748]), .Z(n6196) );
  AND U1235 ( .A(n13451), .B(n6196), .Z(n5553) );
  NANDN U1236 ( .A(y[1747]), .B(x[1747]), .Z(n9353) );
  NANDN U1237 ( .A(x[1747]), .B(y[1747]), .Z(n6197) );
  NANDN U1238 ( .A(y[1744]), .B(x[1744]), .Z(n782) );
  NANDN U1239 ( .A(y[1743]), .B(x[1743]), .Z(n781) );
  NAND U1240 ( .A(n782), .B(n781), .Z(n13437) );
  NANDN U1241 ( .A(x[1742]), .B(y[1742]), .Z(n784) );
  NANDN U1242 ( .A(x[1743]), .B(y[1743]), .Z(n783) );
  NAND U1243 ( .A(n784), .B(n783), .Z(n13436) );
  NANDN U1244 ( .A(y[1739]), .B(x[1739]), .Z(n9336) );
  ANDN U1245 ( .B(x[1738]), .A(y[1738]), .Z(n9335) );
  NANDN U1246 ( .A(y[1737]), .B(x[1737]), .Z(n785) );
  NANDN U1247 ( .A(n9335), .B(n785), .Z(n13431) );
  NANDN U1248 ( .A(x[1734]), .B(y[1734]), .Z(n9319) );
  ANDN U1249 ( .B(y[1732]), .A(x[1732]), .Z(n13424) );
  NANDN U1250 ( .A(y[1731]), .B(x[1731]), .Z(n13423) );
  NANDN U1251 ( .A(y[1728]), .B(x[1728]), .Z(n787) );
  NANDN U1252 ( .A(y[1727]), .B(x[1727]), .Z(n786) );
  NAND U1253 ( .A(n787), .B(n786), .Z(n13417) );
  NANDN U1254 ( .A(x[1726]), .B(y[1726]), .Z(n789) );
  NANDN U1255 ( .A(x[1727]), .B(y[1727]), .Z(n788) );
  AND U1256 ( .A(n789), .B(n788), .Z(n13414) );
  NANDN U1257 ( .A(y[1724]), .B(x[1724]), .Z(n791) );
  NANDN U1258 ( .A(y[1723]), .B(x[1723]), .Z(n790) );
  NAND U1259 ( .A(n791), .B(n790), .Z(n13409) );
  NANDN U1260 ( .A(x[1722]), .B(y[1722]), .Z(n793) );
  NANDN U1261 ( .A(x[1723]), .B(y[1723]), .Z(n792) );
  NAND U1262 ( .A(n793), .B(n792), .Z(n13407) );
  NANDN U1263 ( .A(y[1717]), .B(x[1717]), .Z(n13392) );
  NANDN U1264 ( .A(x[1716]), .B(y[1716]), .Z(n795) );
  NANDN U1265 ( .A(x[1717]), .B(y[1717]), .Z(n794) );
  AND U1266 ( .A(n795), .B(n794), .Z(n13390) );
  NANDN U1267 ( .A(x[1715]), .B(y[1715]), .Z(n13384) );
  ANDN U1268 ( .B(x[1714]), .A(y[1714]), .Z(n13383) );
  ANDN U1269 ( .B(x[1715]), .A(y[1715]), .Z(n13386) );
  OR U1270 ( .A(n13383), .B(n13386), .Z(n9282) );
  NANDN U1271 ( .A(x[1713]), .B(y[1713]), .Z(n797) );
  NANDN U1272 ( .A(x[1714]), .B(y[1714]), .Z(n796) );
  NAND U1273 ( .A(n797), .B(n796), .Z(n13381) );
  NANDN U1274 ( .A(x[1712]), .B(y[1712]), .Z(n799) );
  NANDN U1275 ( .A(x[1711]), .B(y[1711]), .Z(n798) );
  NAND U1276 ( .A(n799), .B(n798), .Z(n13377) );
  NANDN U1277 ( .A(y[1708]), .B(x[1708]), .Z(n9273) );
  NANDN U1278 ( .A(y[1707]), .B(x[1707]), .Z(n800) );
  NAND U1279 ( .A(n9273), .B(n800), .Z(n13365) );
  ANDN U1280 ( .B(x[1706]), .A(y[1706]), .Z(n13358) );
  ANDN U1281 ( .B(x[1705]), .A(y[1705]), .Z(n9261) );
  NOR U1282 ( .A(n13358), .B(n9261), .Z(n5474) );
  NANDN U1283 ( .A(y[1703]), .B(x[1703]), .Z(n13354) );
  ANDN U1284 ( .B(x[1704]), .A(y[1704]), .Z(n9260) );
  ANDN U1285 ( .B(n13354), .A(n9260), .Z(n5471) );
  IV U1286 ( .A(x[1702]), .Z(n6211) );
  IV U1287 ( .A(y[1702]), .Z(n6210) );
  NANDN U1288 ( .A(n6211), .B(n6210), .Z(n801) );
  IV U1289 ( .A(x[1701]), .Z(n6212) );
  NAND U1290 ( .A(n801), .B(n9251), .Z(n13351) );
  IV U1291 ( .A(y[1700]), .Z(n6214) );
  IV U1292 ( .A(x[1700]), .Z(n6213) );
  NANDN U1293 ( .A(n6214), .B(n6213), .Z(n803) );
  NANDN U1294 ( .A(x[1701]), .B(y[1701]), .Z(n802) );
  NAND U1295 ( .A(n803), .B(n802), .Z(n13349) );
  NANDN U1296 ( .A(x[1699]), .B(y[1699]), .Z(n13340) );
  NANDN U1297 ( .A(x[1696]), .B(y[1696]), .Z(n13336) );
  ANDN U1298 ( .B(y[1697]), .A(x[1697]), .Z(n9237) );
  ANDN U1299 ( .B(n13336), .A(n9237), .Z(n5460) );
  NANDN U1300 ( .A(x[1694]), .B(y[1694]), .Z(n9225) );
  NANDN U1301 ( .A(x[1695]), .B(y[1695]), .Z(n6215) );
  NAND U1302 ( .A(n9225), .B(n6215), .Z(n13333) );
  NANDN U1303 ( .A(x[1693]), .B(y[1693]), .Z(n13328) );
  ANDN U1304 ( .B(y[1692]), .A(x[1692]), .Z(n9218) );
  ANDN U1305 ( .B(n13328), .A(n9218), .Z(n5454) );
  ANDN U1306 ( .B(y[1690]), .A(x[1690]), .Z(n13321) );
  NANDN U1307 ( .A(y[1689]), .B(x[1689]), .Z(n13318) );
  NANDN U1308 ( .A(x[1688]), .B(y[1688]), .Z(n804) );
  NANDN U1309 ( .A(x[1689]), .B(y[1689]), .Z(n9214) );
  NAND U1310 ( .A(n804), .B(n9214), .Z(n13317) );
  NANDN U1311 ( .A(y[1687]), .B(x[1687]), .Z(n6223) );
  IV U1312 ( .A(x[1688]), .Z(n6221) );
  IV U1313 ( .A(y[1688]), .Z(n6220) );
  NANDN U1314 ( .A(n6221), .B(n6220), .Z(n805) );
  NAND U1315 ( .A(n6223), .B(n805), .Z(n13315) );
  NANDN U1316 ( .A(x[1686]), .B(y[1686]), .Z(n806) );
  NANDN U1317 ( .A(x[1687]), .B(y[1687]), .Z(n9209) );
  NAND U1318 ( .A(n806), .B(n9209), .Z(n13312) );
  NANDN U1319 ( .A(y[1686]), .B(x[1686]), .Z(n6222) );
  NANDN U1320 ( .A(y[1685]), .B(x[1685]), .Z(n6225) );
  NAND U1321 ( .A(n6222), .B(n6225), .Z(n13311) );
  IV U1322 ( .A(x[1684]), .Z(n6227) );
  IV U1323 ( .A(y[1684]), .Z(n6226) );
  NANDN U1324 ( .A(n6227), .B(n6226), .Z(n807) );
  NANDN U1325 ( .A(y[1683]), .B(x[1683]), .Z(n6229) );
  NAND U1326 ( .A(n807), .B(n6229), .Z(n13307) );
  NANDN U1327 ( .A(x[1677]), .B(y[1677]), .Z(n808) );
  ANDN U1328 ( .B(y[1678]), .A(x[1678]), .Z(n5427) );
  ANDN U1329 ( .B(n808), .A(n5427), .Z(n13290) );
  NANDN U1330 ( .A(y[1673]), .B(x[1673]), .Z(n809) );
  NANDN U1331 ( .A(y[1674]), .B(x[1674]), .Z(n9172) );
  NAND U1332 ( .A(n809), .B(n9172), .Z(n13280) );
  IV U1333 ( .A(x[1671]), .Z(n5414) );
  IV U1334 ( .A(y[1671]), .Z(n5412) );
  NANDN U1335 ( .A(n5414), .B(n5412), .Z(n811) );
  NANDN U1336 ( .A(y[1670]), .B(x[1670]), .Z(n810) );
  NAND U1337 ( .A(n811), .B(n810), .Z(n6238) );
  NANDN U1338 ( .A(y[1669]), .B(x[1669]), .Z(n812) );
  NANDN U1339 ( .A(n6238), .B(n812), .Z(n13273) );
  NANDN U1340 ( .A(x[1669]), .B(y[1669]), .Z(n6235) );
  IV U1341 ( .A(y[1666]), .Z(n6242) );
  NANDN U1342 ( .A(x[1667]), .B(y[1667]), .Z(n6241) );
  NAND U1343 ( .A(n9156), .B(n6241), .Z(n13267) );
  NANDN U1344 ( .A(y[1666]), .B(x[1666]), .Z(n816) );
  NANDN U1345 ( .A(x[1665]), .B(y[1665]), .Z(n5403) );
  IV U1346 ( .A(n5403), .Z(n9151) );
  NANDN U1347 ( .A(y[1664]), .B(x[1664]), .Z(n814) );
  NANDN U1348 ( .A(y[1665]), .B(x[1665]), .Z(n813) );
  NAND U1349 ( .A(n814), .B(n813), .Z(n9149) );
  NANDN U1350 ( .A(n9151), .B(n9149), .Z(n815) );
  NAND U1351 ( .A(n816), .B(n815), .Z(n13264) );
  ANDN U1352 ( .B(x[1663]), .A(y[1663]), .Z(n9144) );
  NANDN U1353 ( .A(y[1661]), .B(x[1661]), .Z(n13257) );
  ANDN U1354 ( .B(x[1662]), .A(y[1662]), .Z(n9145) );
  ANDN U1355 ( .B(n13257), .A(n9145), .Z(n5398) );
  NANDN U1356 ( .A(x[1660]), .B(y[1660]), .Z(n818) );
  NANDN U1357 ( .A(x[1661]), .B(y[1661]), .Z(n817) );
  NAND U1358 ( .A(n818), .B(n817), .Z(n13255) );
  NANDN U1359 ( .A(y[1657]), .B(x[1657]), .Z(n13248) );
  NANDN U1360 ( .A(y[1656]), .B(x[1656]), .Z(n820) );
  NANDN U1361 ( .A(y[1655]), .B(x[1655]), .Z(n819) );
  NAND U1362 ( .A(n820), .B(n819), .Z(n13243) );
  NANDN U1363 ( .A(x[1652]), .B(y[1652]), .Z(n9127) );
  NANDN U1364 ( .A(x[1653]), .B(y[1653]), .Z(n9131) );
  NAND U1365 ( .A(n9127), .B(n9131), .Z(n13236) );
  ANDN U1366 ( .B(x[1644]), .A(y[1644]), .Z(n13214) );
  ANDN U1367 ( .B(x[1643]), .A(y[1643]), .Z(n9102) );
  NOR U1368 ( .A(n13214), .B(n9102), .Z(n5361) );
  NANDN U1369 ( .A(x[1643]), .B(y[1643]), .Z(n13212) );
  NANDN U1370 ( .A(x[1642]), .B(y[1642]), .Z(n821) );
  AND U1371 ( .A(n13212), .B(n821), .Z(n5359) );
  IV U1372 ( .A(y[1642]), .Z(n9098) );
  IV U1373 ( .A(x[1642]), .Z(n9097) );
  XNOR U1374 ( .A(n9098), .B(n9097), .Z(n5357) );
  NANDN U1375 ( .A(y[1641]), .B(x[1641]), .Z(n13206) );
  ANDN U1376 ( .B(y[1637]), .A(x[1637]), .Z(n826) );
  NANDN U1377 ( .A(y[1636]), .B(x[1636]), .Z(n9088) );
  OR U1378 ( .A(n826), .B(n9088), .Z(n824) );
  NANDN U1379 ( .A(y[1637]), .B(x[1637]), .Z(n823) );
  NANDN U1380 ( .A(y[1638]), .B(x[1638]), .Z(n822) );
  AND U1381 ( .A(n823), .B(n822), .Z(n9091) );
  NAND U1382 ( .A(n824), .B(n9091), .Z(n13198) );
  NANDN U1383 ( .A(x[1636]), .B(y[1636]), .Z(n825) );
  NANDN U1384 ( .A(n826), .B(n825), .Z(n13197) );
  ANDN U1385 ( .B(y[1633]), .A(x[1633]), .Z(n9083) );
  NANDN U1386 ( .A(y[1633]), .B(x[1633]), .Z(n5335) );
  NANDN U1387 ( .A(x[1632]), .B(y[1632]), .Z(n9078) );
  NOR U1388 ( .A(n9083), .B(n13190), .Z(n5339) );
  ANDN U1389 ( .B(y[1631]), .A(x[1631]), .Z(n13187) );
  NANDN U1390 ( .A(y[1630]), .B(x[1630]), .Z(n828) );
  NANDN U1391 ( .A(y[1631]), .B(x[1631]), .Z(n827) );
  NAND U1392 ( .A(n828), .B(n827), .Z(n13185) );
  NANDN U1393 ( .A(x[1629]), .B(y[1629]), .Z(n830) );
  NANDN U1394 ( .A(x[1630]), .B(y[1630]), .Z(n829) );
  AND U1395 ( .A(n830), .B(n829), .Z(n13182) );
  NANDN U1396 ( .A(x[1628]), .B(y[1628]), .Z(n13178) );
  NANDN U1397 ( .A(y[1627]), .B(x[1627]), .Z(n13176) );
  ANDN U1398 ( .B(x[1626]), .A(y[1626]), .Z(n5325) );
  NANDN U1399 ( .A(y[1625]), .B(x[1625]), .Z(n831) );
  NANDN U1400 ( .A(n5325), .B(n831), .Z(n13173) );
  ANDN U1401 ( .B(x[1624]), .A(y[1624]), .Z(n13167) );
  OR U1402 ( .A(n13173), .B(n13167), .Z(n9069) );
  NANDN U1403 ( .A(x[1624]), .B(y[1624]), .Z(n13170) );
  NANDN U1404 ( .A(y[1623]), .B(x[1623]), .Z(n6254) );
  XNOR U1405 ( .A(x[1623]), .B(y[1623]), .Z(n5319) );
  NANDN U1406 ( .A(y[1622]), .B(x[1622]), .Z(n6255) );
  NANDN U1407 ( .A(y[1621]), .B(x[1621]), .Z(n832) );
  AND U1408 ( .A(n6255), .B(n832), .Z(n5316) );
  IV U1409 ( .A(x[1621]), .Z(n6257) );
  IV U1410 ( .A(y[1621]), .Z(n6256) );
  XNOR U1411 ( .A(n6257), .B(n6256), .Z(n5314) );
  IV U1412 ( .A(x[1620]), .Z(n833) );
  XOR U1413 ( .A(y[1620]), .B(n833), .Z(n5311) );
  ANDN U1414 ( .B(y[1618]), .A(x[1618]), .Z(n13153) );
  ANDN U1415 ( .B(x[1617]), .A(y[1617]), .Z(n13151) );
  ANDN U1416 ( .B(y[1617]), .A(x[1617]), .Z(n5300) );
  ANDN U1417 ( .B(x[1616]), .A(y[1616]), .Z(n13144) );
  NANDN U1418 ( .A(n5300), .B(n13144), .Z(n834) );
  NANDN U1419 ( .A(n13151), .B(n834), .Z(n9056) );
  NANDN U1420 ( .A(x[1613]), .B(y[1613]), .Z(n13139) );
  ANDN U1421 ( .B(y[1612]), .A(x[1612]), .Z(n13135) );
  ANDN U1422 ( .B(n13139), .A(n13135), .Z(n5295) );
  NANDN U1423 ( .A(x[1606]), .B(y[1606]), .Z(n836) );
  NANDN U1424 ( .A(x[1607]), .B(y[1607]), .Z(n835) );
  NAND U1425 ( .A(n836), .B(n835), .Z(n13119) );
  NANDN U1426 ( .A(y[1606]), .B(x[1606]), .Z(n838) );
  NANDN U1427 ( .A(y[1605]), .B(x[1605]), .Z(n837) );
  NAND U1428 ( .A(n838), .B(n837), .Z(n13117) );
  NANDN U1429 ( .A(x[1604]), .B(y[1604]), .Z(n840) );
  NANDN U1430 ( .A(x[1605]), .B(y[1605]), .Z(n839) );
  AND U1431 ( .A(n840), .B(n839), .Z(n13114) );
  NANDN U1432 ( .A(y[1600]), .B(x[1600]), .Z(n13104) );
  ANDN U1433 ( .B(x[1601]), .A(y[1601]), .Z(n13108) );
  ANDN U1434 ( .B(n13104), .A(n13108), .Z(n841) );
  ANDN U1435 ( .B(y[1601]), .A(x[1601]), .Z(n5272) );
  OR U1436 ( .A(n841), .B(n5272), .Z(n9027) );
  NANDN U1437 ( .A(y[1599]), .B(x[1599]), .Z(n843) );
  NANDN U1438 ( .A(y[1598]), .B(x[1598]), .Z(n842) );
  AND U1439 ( .A(n843), .B(n842), .Z(n13100) );
  NANDN U1440 ( .A(x[1598]), .B(y[1598]), .Z(n845) );
  NANDN U1441 ( .A(x[1597]), .B(y[1597]), .Z(n844) );
  NAND U1442 ( .A(n845), .B(n844), .Z(n13099) );
  NANDN U1443 ( .A(x[1588]), .B(y[1588]), .Z(n847) );
  NANDN U1444 ( .A(x[1589]), .B(y[1589]), .Z(n846) );
  NAND U1445 ( .A(n847), .B(n846), .Z(n13083) );
  NANDN U1446 ( .A(x[1587]), .B(y[1587]), .Z(n13078) );
  NANDN U1447 ( .A(y[1586]), .B(x[1586]), .Z(n849) );
  NANDN U1448 ( .A(y[1587]), .B(x[1587]), .Z(n848) );
  NAND U1449 ( .A(n849), .B(n848), .Z(n13077) );
  NANDN U1450 ( .A(y[1585]), .B(x[1585]), .Z(n6274) );
  XNOR U1451 ( .A(x[1585]), .B(y[1585]), .Z(n5242) );
  NANDN U1452 ( .A(y[1584]), .B(x[1584]), .Z(n6275) );
  NANDN U1453 ( .A(y[1583]), .B(x[1583]), .Z(n850) );
  AND U1454 ( .A(n6275), .B(n850), .Z(n5239) );
  IV U1455 ( .A(x[1583]), .Z(n8995) );
  IV U1456 ( .A(y[1583]), .Z(n8994) );
  XNOR U1457 ( .A(n8995), .B(n8994), .Z(n5237) );
  NANDN U1458 ( .A(x[1582]), .B(y[1582]), .Z(n13066) );
  NANDN U1459 ( .A(y[1581]), .B(x[1581]), .Z(n13065) );
  ANDN U1460 ( .B(y[1581]), .A(x[1581]), .Z(n6276) );
  ANDN U1461 ( .B(y[1580]), .A(x[1580]), .Z(n8987) );
  NOR U1462 ( .A(n6276), .B(n8987), .Z(n13062) );
  NANDN U1463 ( .A(x[1579]), .B(y[1579]), .Z(n13058) );
  NANDN U1464 ( .A(y[1578]), .B(x[1578]), .Z(n8985) );
  XNOR U1465 ( .A(x[1578]), .B(y[1578]), .Z(n5227) );
  NANDN U1466 ( .A(x[1577]), .B(y[1577]), .Z(n6277) );
  NANDN U1467 ( .A(x[1574]), .B(y[1574]), .Z(n8977) );
  NANDN U1468 ( .A(y[1573]), .B(x[1573]), .Z(n5214) );
  IV U1469 ( .A(x[1573]), .Z(n6280) );
  IV U1470 ( .A(y[1573]), .Z(n6279) );
  XNOR U1471 ( .A(n6280), .B(n6279), .Z(n5212) );
  NANDN U1472 ( .A(y[1572]), .B(x[1572]), .Z(n6282) );
  NANDN U1473 ( .A(y[1571]), .B(x[1571]), .Z(n8973) );
  AND U1474 ( .A(n6282), .B(n8973), .Z(n5209) );
  XNOR U1475 ( .A(x[1571]), .B(y[1571]), .Z(n5207) );
  NANDN U1476 ( .A(x[1570]), .B(y[1570]), .Z(n13038) );
  NANDN U1477 ( .A(y[1568]), .B(x[1568]), .Z(n13032) );
  ANDN U1478 ( .B(x[1567]), .A(y[1567]), .Z(n8962) );
  ANDN U1479 ( .B(n13032), .A(n8962), .Z(n5201) );
  ANDN U1480 ( .B(x[1566]), .A(y[1566]), .Z(n8961) );
  ANDN U1481 ( .B(x[1562]), .A(y[1562]), .Z(n13017) );
  ANDN U1482 ( .B(x[1563]), .A(y[1563]), .Z(n9994) );
  NOR U1483 ( .A(n13017), .B(n9994), .Z(n8953) );
  NANDN U1484 ( .A(x[1561]), .B(y[1561]), .Z(n13014) );
  ANDN U1485 ( .B(y[1558]), .A(x[1558]), .Z(n13007) );
  NANDN U1486 ( .A(y[1557]), .B(x[1557]), .Z(n13005) );
  ANDN U1487 ( .B(x[1558]), .A(y[1558]), .Z(n8943) );
  ANDN U1488 ( .B(n13005), .A(n8943), .Z(n5177) );
  NANDN U1489 ( .A(y[1556]), .B(x[1556]), .Z(n13000) );
  NANDN U1490 ( .A(y[1555]), .B(x[1555]), .Z(n8932) );
  AND U1491 ( .A(n13000), .B(n8932), .Z(n5174) );
  NANDN U1492 ( .A(x[1554]), .B(y[1554]), .Z(n12994) );
  NANDN U1493 ( .A(x[1555]), .B(y[1555]), .Z(n12998) );
  NAND U1494 ( .A(n12994), .B(n12998), .Z(n5172) );
  NANDN U1495 ( .A(y[1554]), .B(x[1554]), .Z(n8933) );
  NANDN U1496 ( .A(x[1550]), .B(y[1550]), .Z(n6285) );
  XNOR U1497 ( .A(y[1550]), .B(x[1550]), .Z(n5163) );
  NANDN U1498 ( .A(x[1549]), .B(y[1549]), .Z(n6286) );
  NANDN U1499 ( .A(x[1548]), .B(y[1548]), .Z(n8917) );
  AND U1500 ( .A(n6286), .B(n8917), .Z(n5160) );
  XNOR U1501 ( .A(y[1548]), .B(x[1548]), .Z(n5158) );
  NANDN U1502 ( .A(x[1547]), .B(y[1547]), .Z(n8918) );
  NANDN U1503 ( .A(x[1546]), .B(y[1546]), .Z(n851) );
  AND U1504 ( .A(n8918), .B(n851), .Z(n5155) );
  IV U1505 ( .A(y[1546]), .Z(n6288) );
  IV U1506 ( .A(x[1546]), .Z(n6287) );
  XNOR U1507 ( .A(n6288), .B(n6287), .Z(n5153) );
  NANDN U1508 ( .A(y[1545]), .B(x[1545]), .Z(n12970) );
  NANDN U1509 ( .A(x[1544]), .B(y[1544]), .Z(n8908) );
  IV U1510 ( .A(y[1544]), .Z(n12971) );
  NAND U1511 ( .A(n12971), .B(x[1544]), .Z(n8910) );
  ANDN U1512 ( .B(x[1543]), .A(y[1543]), .Z(n8905) );
  ANDN U1513 ( .B(n8910), .A(n8905), .Z(n5148) );
  ANDN U1514 ( .B(y[1542]), .A(x[1542]), .Z(n12964) );
  NANDN U1515 ( .A(x[1543]), .B(y[1543]), .Z(n12967) );
  NANDN U1516 ( .A(n12964), .B(n12967), .Z(n5146) );
  ANDN U1517 ( .B(x[1542]), .A(y[1542]), .Z(n8904) );
  ANDN U1518 ( .B(n12961), .A(n8904), .Z(n5144) );
  NANDN U1519 ( .A(x[1539]), .B(y[1539]), .Z(n853) );
  NANDN U1520 ( .A(x[1540]), .B(y[1540]), .Z(n852) );
  AND U1521 ( .A(n853), .B(n852), .Z(n855) );
  NANDN U1522 ( .A(x[1541]), .B(y[1541]), .Z(n854) );
  NAND U1523 ( .A(n855), .B(n854), .Z(n12960) );
  NANDN U1524 ( .A(x[1538]), .B(y[1538]), .Z(n857) );
  NANDN U1525 ( .A(x[1537]), .B(y[1537]), .Z(n856) );
  NAND U1526 ( .A(n857), .B(n856), .Z(n12956) );
  NANDN U1527 ( .A(y[1536]), .B(x[1536]), .Z(n859) );
  NANDN U1528 ( .A(y[1537]), .B(x[1537]), .Z(n858) );
  AND U1529 ( .A(n859), .B(n858), .Z(n12953) );
  ANDN U1530 ( .B(x[1532]), .A(y[1532]), .Z(n12942) );
  ANDN U1531 ( .B(x[1531]), .A(y[1531]), .Z(n8883) );
  NOR U1532 ( .A(n12942), .B(n8883), .Z(n5128) );
  NANDN U1533 ( .A(x[1531]), .B(y[1531]), .Z(n12940) );
  NANDN U1534 ( .A(y[1525]), .B(x[1525]), .Z(n861) );
  NANDN U1535 ( .A(y[1524]), .B(x[1524]), .Z(n860) );
  AND U1536 ( .A(n861), .B(n860), .Z(n8875) );
  NANDN U1537 ( .A(x[1524]), .B(y[1524]), .Z(n862) );
  ANDN U1538 ( .B(x[1523]), .A(y[1523]), .Z(n8872) );
  NAND U1539 ( .A(n862), .B(n8872), .Z(n5107) );
  NANDN U1540 ( .A(x[1522]), .B(y[1522]), .Z(n864) );
  NANDN U1541 ( .A(x[1523]), .B(y[1523]), .Z(n863) );
  NAND U1542 ( .A(n863), .B(n862), .Z(n8874) );
  ANDN U1543 ( .B(n864), .A(n8874), .Z(n12923) );
  NANDN U1544 ( .A(x[1521]), .B(y[1521]), .Z(n8869) );
  NANDN U1545 ( .A(x[1520]), .B(y[1520]), .Z(n8864) );
  NAND U1546 ( .A(n8869), .B(n8864), .Z(n12920) );
  NANDN U1547 ( .A(y[1520]), .B(x[1520]), .Z(n12917) );
  NANDN U1548 ( .A(y[1516]), .B(x[1516]), .Z(n865) );
  NANDN U1549 ( .A(y[1517]), .B(x[1517]), .Z(n5092) );
  AND U1550 ( .A(n865), .B(n5092), .Z(n12911) );
  NANDN U1551 ( .A(x[1514]), .B(y[1514]), .Z(n867) );
  NANDN U1552 ( .A(x[1513]), .B(y[1513]), .Z(n866) );
  NAND U1553 ( .A(n867), .B(n866), .Z(n12905) );
  NANDN U1554 ( .A(y[1511]), .B(x[1511]), .Z(n8847) );
  NANDN U1555 ( .A(x[1512]), .B(y[1512]), .Z(n5078) );
  NANDN U1556 ( .A(n8847), .B(n5078), .Z(n5085) );
  NANDN U1557 ( .A(y[1509]), .B(x[1509]), .Z(n12899) );
  NANDN U1558 ( .A(y[1510]), .B(x[1510]), .Z(n8846) );
  AND U1559 ( .A(n12899), .B(n8846), .Z(n5076) );
  NANDN U1560 ( .A(y[1508]), .B(x[1508]), .Z(n8841) );
  ANDN U1561 ( .B(y[1507]), .A(x[1507]), .Z(n8836) );
  NANDN U1562 ( .A(y[1507]), .B(x[1507]), .Z(n869) );
  NANDN U1563 ( .A(y[1506]), .B(x[1506]), .Z(n868) );
  AND U1564 ( .A(n869), .B(n868), .Z(n8834) );
  OR U1565 ( .A(n8836), .B(n8834), .Z(n870) );
  NAND U1566 ( .A(n8841), .B(n870), .Z(n12895) );
  NANDN U1567 ( .A(y[1504]), .B(x[1504]), .Z(n872) );
  NANDN U1568 ( .A(y[1505]), .B(x[1505]), .Z(n871) );
  AND U1569 ( .A(n872), .B(n871), .Z(n12891) );
  NANDN U1570 ( .A(x[1504]), .B(y[1504]), .Z(n874) );
  NANDN U1571 ( .A(x[1503]), .B(y[1503]), .Z(n873) );
  NAND U1572 ( .A(n874), .B(n873), .Z(n12890) );
  NANDN U1573 ( .A(y[1501]), .B(x[1501]), .Z(n6295) );
  NANDN U1574 ( .A(x[1502]), .B(y[1502]), .Z(n5059) );
  NANDN U1575 ( .A(n6295), .B(n5059), .Z(n5067) );
  NANDN U1576 ( .A(y[1502]), .B(x[1502]), .Z(n876) );
  NANDN U1577 ( .A(y[1503]), .B(x[1503]), .Z(n875) );
  AND U1578 ( .A(n876), .B(n875), .Z(n12887) );
  ANDN U1579 ( .B(x[1499]), .A(y[1499]), .Z(n8824) );
  NANDN U1580 ( .A(x[1499]), .B(y[1499]), .Z(n6298) );
  ANDN U1581 ( .B(x[1496]), .A(y[1496]), .Z(n12872) );
  ANDN U1582 ( .B(x[1495]), .A(y[1495]), .Z(n8813) );
  NOR U1583 ( .A(n12872), .B(n8813), .Z(n5051) );
  NANDN U1584 ( .A(x[1492]), .B(y[1492]), .Z(n6299) );
  ANDN U1585 ( .B(x[1493]), .A(y[1493]), .Z(n5042) );
  NOR U1586 ( .A(n6299), .B(n5042), .Z(n877) );
  NANDN U1587 ( .A(y[1494]), .B(x[1494]), .Z(n5045) );
  NAND U1588 ( .A(n877), .B(n5045), .Z(n878) );
  NANDN U1589 ( .A(x[1495]), .B(y[1495]), .Z(n12869) );
  NAND U1590 ( .A(n878), .B(n12869), .Z(n5049) );
  NANDN U1591 ( .A(x[1494]), .B(y[1494]), .Z(n880) );
  NANDN U1592 ( .A(x[1493]), .B(y[1493]), .Z(n879) );
  NAND U1593 ( .A(n880), .B(n879), .Z(n5044) );
  NANDN U1594 ( .A(x[1491]), .B(y[1491]), .Z(n881) );
  NANDN U1595 ( .A(n5044), .B(n881), .Z(n6300) );
  NANDN U1596 ( .A(x[1488]), .B(y[1488]), .Z(n8805) );
  NANDN U1597 ( .A(y[1482]), .B(x[1482]), .Z(n8799) );
  NANDN U1598 ( .A(x[1481]), .B(y[1481]), .Z(n5008) );
  XNOR U1599 ( .A(x[1481]), .B(y[1481]), .Z(n883) );
  NANDN U1600 ( .A(y[1480]), .B(x[1480]), .Z(n882) );
  NAND U1601 ( .A(n883), .B(n882), .Z(n884) );
  AND U1602 ( .A(n5008), .B(n884), .Z(n12848) );
  ANDN U1603 ( .B(n8799), .A(n12848), .Z(n5012) );
  NANDN U1604 ( .A(y[1479]), .B(x[1479]), .Z(n886) );
  NANDN U1605 ( .A(y[1478]), .B(x[1478]), .Z(n885) );
  NAND U1606 ( .A(n886), .B(n885), .Z(n12843) );
  NANDN U1607 ( .A(y[1477]), .B(x[1477]), .Z(n6307) );
  NANDN U1608 ( .A(y[1475]), .B(x[1475]), .Z(n888) );
  NANDN U1609 ( .A(y[1474]), .B(x[1474]), .Z(n887) );
  NAND U1610 ( .A(n888), .B(n887), .Z(n12836) );
  ANDN U1611 ( .B(y[1471]), .A(x[1471]), .Z(n6313) );
  NANDN U1612 ( .A(x[1470]), .B(y[1470]), .Z(n889) );
  NANDN U1613 ( .A(n6313), .B(n889), .Z(n12830) );
  NANDN U1614 ( .A(y[1470]), .B(x[1470]), .Z(n6312) );
  NANDN U1615 ( .A(y[1467]), .B(x[1467]), .Z(n891) );
  ANDN U1616 ( .B(x[1468]), .A(y[1468]), .Z(n890) );
  ANDN U1617 ( .B(n891), .A(n890), .Z(n895) );
  XNOR U1618 ( .A(x[1467]), .B(y[1467]), .Z(n893) );
  ANDN U1619 ( .B(x[1466]), .A(y[1466]), .Z(n892) );
  NAND U1620 ( .A(n893), .B(n892), .Z(n894) );
  AND U1621 ( .A(n895), .B(n894), .Z(n12823) );
  NANDN U1622 ( .A(x[1466]), .B(y[1466]), .Z(n897) );
  NANDN U1623 ( .A(x[1465]), .B(y[1465]), .Z(n896) );
  AND U1624 ( .A(n897), .B(n896), .Z(n899) );
  NANDN U1625 ( .A(x[1467]), .B(y[1467]), .Z(n898) );
  NAND U1626 ( .A(n899), .B(n898), .Z(n12822) );
  NANDN U1627 ( .A(x[1464]), .B(y[1464]), .Z(n4973) );
  IV U1628 ( .A(y[1464]), .Z(n8774) );
  IV U1629 ( .A(x[1464]), .Z(n8773) );
  XNOR U1630 ( .A(n8774), .B(n8773), .Z(n4971) );
  NANDN U1631 ( .A(x[1463]), .B(y[1463]), .Z(n8776) );
  XNOR U1632 ( .A(x[1463]), .B(y[1463]), .Z(n4968) );
  NANDN U1633 ( .A(y[1461]), .B(x[1461]), .Z(n12811) );
  ANDN U1634 ( .B(x[1462]), .A(y[1462]), .Z(n8771) );
  ANDN U1635 ( .B(n12811), .A(n8771), .Z(n4965) );
  ANDN U1636 ( .B(y[1459]), .A(x[1459]), .Z(n12806) );
  ANDN U1637 ( .B(y[1458]), .A(x[1458]), .Z(n8758) );
  NOR U1638 ( .A(n12806), .B(n8758), .Z(n4960) );
  ANDN U1639 ( .B(y[1457]), .A(x[1457]), .Z(n8757) );
  NANDN U1640 ( .A(x[1454]), .B(y[1454]), .Z(n901) );
  NANDN U1641 ( .A(x[1453]), .B(y[1453]), .Z(n900) );
  AND U1642 ( .A(n901), .B(n900), .Z(n12793) );
  ANDN U1643 ( .B(x[1453]), .A(y[1453]), .Z(n902) );
  ANDN U1644 ( .B(y[1452]), .A(x[1452]), .Z(n6317) );
  NANDN U1645 ( .A(n902), .B(n6317), .Z(n4946) );
  NANDN U1646 ( .A(y[1452]), .B(x[1452]), .Z(n903) );
  ANDN U1647 ( .B(n903), .A(n902), .Z(n12792) );
  ANDN U1648 ( .B(x[1451]), .A(y[1451]), .Z(n8749) );
  ANDN U1649 ( .B(n12792), .A(n8749), .Z(n4944) );
  NANDN U1650 ( .A(y[1448]), .B(x[1448]), .Z(n12775) );
  ANDN U1651 ( .B(x[1447]), .A(y[1447]), .Z(n6320) );
  ANDN U1652 ( .B(n12775), .A(n6320), .Z(n4937) );
  NANDN U1653 ( .A(y[1443]), .B(x[1443]), .Z(n905) );
  NANDN U1654 ( .A(y[1442]), .B(x[1442]), .Z(n904) );
  NAND U1655 ( .A(n905), .B(n904), .Z(n12758) );
  NANDN U1656 ( .A(y[1439]), .B(x[1439]), .Z(n8723) );
  NANDN U1657 ( .A(x[1440]), .B(y[1440]), .Z(n907) );
  NANDN U1658 ( .A(n8723), .B(n907), .Z(n4926) );
  NANDN U1659 ( .A(x[1438]), .B(y[1438]), .Z(n908) );
  NANDN U1660 ( .A(x[1439]), .B(y[1439]), .Z(n906) );
  NAND U1661 ( .A(n907), .B(n906), .Z(n8726) );
  ANDN U1662 ( .B(n908), .A(n8726), .Z(n12751) );
  ANDN U1663 ( .B(y[1437]), .A(x[1437]), .Z(n8720) );
  NANDN U1664 ( .A(x[1436]), .B(y[1436]), .Z(n8716) );
  NANDN U1665 ( .A(n8720), .B(n8716), .Z(n12747) );
  ANDN U1666 ( .B(x[1434]), .A(y[1434]), .Z(n8712) );
  NANDN U1667 ( .A(x[1432]), .B(y[1432]), .Z(n8707) );
  NANDN U1668 ( .A(y[1433]), .B(x[1433]), .Z(n913) );
  NANDN U1669 ( .A(n8707), .B(n913), .Z(n911) );
  NANDN U1670 ( .A(x[1433]), .B(y[1433]), .Z(n910) );
  NANDN U1671 ( .A(x[1434]), .B(y[1434]), .Z(n909) );
  AND U1672 ( .A(n910), .B(n909), .Z(n8710) );
  NAND U1673 ( .A(n911), .B(n8710), .Z(n12740) );
  NANDN U1674 ( .A(y[1432]), .B(x[1432]), .Z(n912) );
  NAND U1675 ( .A(n913), .B(n912), .Z(n12738) );
  NANDN U1676 ( .A(y[1429]), .B(x[1429]), .Z(n8701) );
  NANDN U1677 ( .A(x[1428]), .B(y[1428]), .Z(n4903) );
  IV U1678 ( .A(y[1428]), .Z(n6322) );
  IV U1679 ( .A(x[1428]), .Z(n6321) );
  XNOR U1680 ( .A(n6322), .B(n6321), .Z(n4901) );
  NANDN U1681 ( .A(x[1427]), .B(y[1427]), .Z(n6324) );
  ANDN U1682 ( .B(y[1426]), .A(x[1426]), .Z(n6327) );
  ANDN U1683 ( .B(n6324), .A(n6327), .Z(n4898) );
  NANDN U1684 ( .A(x[1425]), .B(y[1425]), .Z(n915) );
  NANDN U1685 ( .A(x[1424]), .B(y[1424]), .Z(n914) );
  NAND U1686 ( .A(n915), .B(n914), .Z(n6325) );
  NANDN U1687 ( .A(y[1417]), .B(x[1417]), .Z(n4873) );
  IV U1688 ( .A(x[1417]), .Z(n8678) );
  IV U1689 ( .A(y[1417]), .Z(n8677) );
  XNOR U1690 ( .A(n8678), .B(n8677), .Z(n4871) );
  NANDN U1691 ( .A(y[1416]), .B(x[1416]), .Z(n8680) );
  NANDN U1692 ( .A(y[1415]), .B(x[1415]), .Z(n6328) );
  AND U1693 ( .A(n8680), .B(n6328), .Z(n4868) );
  XNOR U1694 ( .A(x[1415]), .B(y[1415]), .Z(n4866) );
  NANDN U1695 ( .A(x[1414]), .B(y[1414]), .Z(n12699) );
  NANDN U1696 ( .A(y[1413]), .B(x[1413]), .Z(n8667) );
  IV U1697 ( .A(n8667), .Z(n12702) );
  NANDN U1698 ( .A(x[1411]), .B(y[1411]), .Z(n12695) );
  NANDN U1699 ( .A(x[1406]), .B(y[1406]), .Z(n917) );
  NANDN U1700 ( .A(x[1405]), .B(y[1405]), .Z(n916) );
  AND U1701 ( .A(n917), .B(n916), .Z(n919) );
  NANDN U1702 ( .A(x[1407]), .B(y[1407]), .Z(n918) );
  NAND U1703 ( .A(n919), .B(n918), .Z(n12688) );
  NANDN U1704 ( .A(y[1405]), .B(x[1405]), .Z(n6331) );
  ANDN U1705 ( .B(x[1403]), .A(y[1403]), .Z(n8654) );
  NANDN U1706 ( .A(x[1403]), .B(y[1403]), .Z(n8657) );
  NANDN U1707 ( .A(y[1400]), .B(x[1400]), .Z(n12673) );
  ANDN U1708 ( .B(x[1399]), .A(y[1399]), .Z(n8642) );
  ANDN U1709 ( .B(n12673), .A(n8642), .Z(n4835) );
  NANDN U1710 ( .A(x[1399]), .B(y[1399]), .Z(n12671) );
  NANDN U1711 ( .A(y[1397]), .B(x[1397]), .Z(n921) );
  NANDN U1712 ( .A(y[1396]), .B(x[1396]), .Z(n920) );
  NAND U1713 ( .A(n921), .B(n920), .Z(n12665) );
  NANDN U1714 ( .A(y[1393]), .B(x[1393]), .Z(n8634) );
  NANDN U1715 ( .A(x[1392]), .B(y[1392]), .Z(n8631) );
  XNOR U1716 ( .A(y[1392]), .B(x[1392]), .Z(n4815) );
  NANDN U1717 ( .A(y[1391]), .B(x[1391]), .Z(n8628) );
  NANDN U1718 ( .A(y[1389]), .B(x[1389]), .Z(n12649) );
  NANDN U1719 ( .A(y[1390]), .B(x[1390]), .Z(n8629) );
  AND U1720 ( .A(n12649), .B(n8629), .Z(n4810) );
  NANDN U1721 ( .A(x[1388]), .B(y[1388]), .Z(n8621) );
  NANDN U1722 ( .A(x[1389]), .B(y[1389]), .Z(n8625) );
  NAND U1723 ( .A(n8621), .B(n8625), .Z(n12648) );
  NANDN U1724 ( .A(y[1383]), .B(x[1383]), .Z(n8613) );
  ANDN U1725 ( .B(y[1380]), .A(x[1380]), .Z(n8608) );
  NANDN U1726 ( .A(y[1380]), .B(x[1380]), .Z(n6336) );
  NANDN U1727 ( .A(y[1379]), .B(x[1379]), .Z(n922) );
  AND U1728 ( .A(n6336), .B(n922), .Z(n4783) );
  IV U1729 ( .A(x[1379]), .Z(n6339) );
  IV U1730 ( .A(y[1379]), .Z(n6338) );
  XNOR U1731 ( .A(n6339), .B(n6338), .Z(n4781) );
  NANDN U1732 ( .A(y[1377]), .B(x[1377]), .Z(n4772) );
  XNOR U1733 ( .A(y[1377]), .B(x[1377]), .Z(n924) );
  NANDN U1734 ( .A(x[1376]), .B(y[1376]), .Z(n923) );
  NAND U1735 ( .A(n924), .B(n923), .Z(n925) );
  AND U1736 ( .A(n4772), .B(n925), .Z(n8605) );
  ANDN U1737 ( .B(y[1375]), .A(x[1375]), .Z(n6343) );
  NANDN U1738 ( .A(x[1374]), .B(y[1374]), .Z(n926) );
  NANDN U1739 ( .A(n6343), .B(n926), .Z(n12620) );
  NANDN U1740 ( .A(y[1374]), .B(x[1374]), .Z(n6342) );
  NANDN U1741 ( .A(x[1373]), .B(y[1373]), .Z(n4764) );
  XNOR U1742 ( .A(x[1373]), .B(y[1373]), .Z(n928) );
  NANDN U1743 ( .A(y[1372]), .B(x[1372]), .Z(n927) );
  NAND U1744 ( .A(n928), .B(n927), .Z(n929) );
  AND U1745 ( .A(n4764), .B(n929), .Z(n12617) );
  ANDN U1746 ( .B(n6342), .A(n12617), .Z(n4768) );
  NANDN U1747 ( .A(y[1370]), .B(x[1370]), .Z(n931) );
  NANDN U1748 ( .A(y[1371]), .B(x[1371]), .Z(n930) );
  AND U1749 ( .A(n931), .B(n930), .Z(n12613) );
  NANDN U1750 ( .A(x[1370]), .B(y[1370]), .Z(n933) );
  NANDN U1751 ( .A(x[1369]), .B(y[1369]), .Z(n932) );
  NAND U1752 ( .A(n933), .B(n932), .Z(n12612) );
  NANDN U1753 ( .A(x[1368]), .B(y[1368]), .Z(n4758) );
  IV U1754 ( .A(y[1368]), .Z(n8591) );
  IV U1755 ( .A(x[1368]), .Z(n8590) );
  XNOR U1756 ( .A(n8591), .B(n8590), .Z(n4756) );
  NANDN U1757 ( .A(x[1367]), .B(y[1367]), .Z(n8593) );
  XNOR U1758 ( .A(x[1367]), .B(y[1367]), .Z(n4753) );
  NANDN U1759 ( .A(y[1365]), .B(x[1365]), .Z(n12601) );
  ANDN U1760 ( .B(x[1366]), .A(y[1366]), .Z(n8588) );
  ANDN U1761 ( .B(n12601), .A(n8588), .Z(n4750) );
  NANDN U1762 ( .A(x[1364]), .B(y[1364]), .Z(n8580) );
  NANDN U1763 ( .A(x[1365]), .B(y[1365]), .Z(n8586) );
  NAND U1764 ( .A(n8580), .B(n8586), .Z(n12599) );
  NANDN U1765 ( .A(x[1360]), .B(y[1360]), .Z(n935) );
  NANDN U1766 ( .A(x[1359]), .B(y[1359]), .Z(n934) );
  NAND U1767 ( .A(n935), .B(n934), .Z(n12591) );
  NANDN U1768 ( .A(x[1354]), .B(y[1354]), .Z(n12579) );
  NANDN U1769 ( .A(y[1353]), .B(x[1353]), .Z(n12578) );
  ANDN U1770 ( .B(y[1352]), .A(x[1352]), .Z(n8559) );
  ANDN U1771 ( .B(y[1353]), .A(x[1353]), .Z(n8566) );
  NOR U1772 ( .A(n8559), .B(n8566), .Z(n12575) );
  NANDN U1773 ( .A(y[1352]), .B(x[1352]), .Z(n12573) );
  NANDN U1774 ( .A(y[1349]), .B(x[1349]), .Z(n12566) );
  NANDN U1775 ( .A(y[1350]), .B(x[1350]), .Z(n8556) );
  AND U1776 ( .A(n12566), .B(n8556), .Z(n4715) );
  NANDN U1777 ( .A(x[1348]), .B(y[1348]), .Z(n937) );
  NANDN U1778 ( .A(x[1349]), .B(y[1349]), .Z(n936) );
  NAND U1779 ( .A(n937), .B(n936), .Z(n12564) );
  NANDN U1780 ( .A(x[1346]), .B(y[1346]), .Z(n939) );
  NANDN U1781 ( .A(x[1345]), .B(y[1345]), .Z(n938) );
  AND U1782 ( .A(n939), .B(n938), .Z(n941) );
  NANDN U1783 ( .A(x[1347]), .B(y[1347]), .Z(n940) );
  NAND U1784 ( .A(n941), .B(n940), .Z(n12560) );
  NANDN U1785 ( .A(y[1345]), .B(x[1345]), .Z(n8549) );
  IV U1786 ( .A(y[1343]), .Z(n8544) );
  IV U1787 ( .A(x[1343]), .Z(n8543) );
  XNOR U1788 ( .A(n8544), .B(n8543), .Z(n4697) );
  ANDN U1789 ( .B(x[1341]), .A(y[1341]), .Z(n12549) );
  ANDN U1790 ( .B(x[1342]), .A(y[1342]), .Z(n8540) );
  NOR U1791 ( .A(n12549), .B(n8540), .Z(n4694) );
  NANDN U1792 ( .A(y[1336]), .B(x[1336]), .Z(n943) );
  NANDN U1793 ( .A(y[1337]), .B(x[1337]), .Z(n942) );
  AND U1794 ( .A(n943), .B(n942), .Z(n12537) );
  NANDN U1795 ( .A(x[1336]), .B(y[1336]), .Z(n945) );
  NANDN U1796 ( .A(x[1335]), .B(y[1335]), .Z(n944) );
  NAND U1797 ( .A(n945), .B(n944), .Z(n12535) );
  NANDN U1798 ( .A(x[1334]), .B(y[1334]), .Z(n947) );
  NANDN U1799 ( .A(x[1333]), .B(y[1333]), .Z(n946) );
  NAND U1800 ( .A(n947), .B(n946), .Z(n12531) );
  NANDN U1801 ( .A(y[1331]), .B(x[1331]), .Z(n8520) );
  NANDN U1802 ( .A(x[1332]), .B(y[1332]), .Z(n4670) );
  NANDN U1803 ( .A(n8520), .B(n4670), .Z(n4677) );
  NANDN U1804 ( .A(y[1326]), .B(x[1326]), .Z(n949) );
  NANDN U1805 ( .A(y[1327]), .B(x[1327]), .Z(n948) );
  NAND U1806 ( .A(n949), .B(n948), .Z(n12518) );
  NANDN U1807 ( .A(x[1326]), .B(y[1326]), .Z(n951) );
  NANDN U1808 ( .A(x[1325]), .B(y[1325]), .Z(n950) );
  NAND U1809 ( .A(n951), .B(n950), .Z(n12515) );
  NANDN U1810 ( .A(x[1324]), .B(y[1324]), .Z(n953) );
  NANDN U1811 ( .A(x[1323]), .B(y[1323]), .Z(n952) );
  NAND U1812 ( .A(n953), .B(n952), .Z(n12511) );
  NANDN U1813 ( .A(y[1321]), .B(x[1321]), .Z(n8504) );
  ANDN U1814 ( .B(y[1318]), .A(x[1318]), .Z(n12500) );
  NANDN U1815 ( .A(y[1317]), .B(x[1317]), .Z(n12498) );
  ANDN U1816 ( .B(y[1316]), .A(x[1316]), .Z(n8496) );
  ANDN U1817 ( .B(y[1317]), .A(x[1317]), .Z(n6354) );
  NOR U1818 ( .A(n8496), .B(n6354), .Z(n12495) );
  NANDN U1819 ( .A(x[1314]), .B(y[1314]), .Z(n955) );
  NANDN U1820 ( .A(x[1313]), .B(y[1313]), .Z(n954) );
  NAND U1821 ( .A(n955), .B(n954), .Z(n12488) );
  NANDN U1822 ( .A(y[1309]), .B(x[1309]), .Z(n4623) );
  IV U1823 ( .A(x[1309]), .Z(n6356) );
  IV U1824 ( .A(y[1309]), .Z(n6355) );
  XNOR U1825 ( .A(n6356), .B(n6355), .Z(n4621) );
  NANDN U1826 ( .A(y[1308]), .B(x[1308]), .Z(n6358) );
  NANDN U1827 ( .A(y[1307]), .B(x[1307]), .Z(n8478) );
  AND U1828 ( .A(n6358), .B(n8478), .Z(n4618) );
  XNOR U1829 ( .A(x[1307]), .B(y[1307]), .Z(n4616) );
  NANDN U1830 ( .A(x[1306]), .B(y[1306]), .Z(n12471) );
  NANDN U1831 ( .A(y[1304]), .B(x[1304]), .Z(n12465) );
  ANDN U1832 ( .B(x[1303]), .A(y[1303]), .Z(n8467) );
  ANDN U1833 ( .B(n12465), .A(n8467), .Z(n4610) );
  NANDN U1834 ( .A(x[1302]), .B(y[1302]), .Z(n12459) );
  NANDN U1835 ( .A(x[1299]), .B(y[1299]), .Z(n957) );
  NANDN U1836 ( .A(x[1300]), .B(y[1300]), .Z(n956) );
  AND U1837 ( .A(n957), .B(n956), .Z(n959) );
  NANDN U1838 ( .A(x[1301]), .B(y[1301]), .Z(n958) );
  NAND U1839 ( .A(n959), .B(n958), .Z(n12456) );
  NANDN U1840 ( .A(x[1298]), .B(y[1298]), .Z(n6360) );
  NANDN U1841 ( .A(y[1297]), .B(x[1297]), .Z(n8459) );
  XNOR U1842 ( .A(x[1297]), .B(y[1297]), .Z(n4594) );
  NANDN U1843 ( .A(y[1296]), .B(x[1296]), .Z(n8460) );
  NANDN U1844 ( .A(y[1295]), .B(x[1295]), .Z(n6362) );
  AND U1845 ( .A(n8460), .B(n6362), .Z(n4591) );
  XNOR U1846 ( .A(x[1295]), .B(y[1295]), .Z(n4589) );
  NANDN U1847 ( .A(x[1294]), .B(y[1294]), .Z(n12443) );
  NANDN U1848 ( .A(y[1293]), .B(x[1293]), .Z(n12441) );
  NANDN U1849 ( .A(x[1291]), .B(y[1291]), .Z(n12436) );
  NANDN U1850 ( .A(y[1290]), .B(x[1290]), .Z(n8445) );
  XNOR U1851 ( .A(x[1290]), .B(y[1290]), .Z(n4579) );
  NANDN U1852 ( .A(x[1289]), .B(y[1289]), .Z(n6364) );
  NANDN U1853 ( .A(x[1288]), .B(y[1288]), .Z(n961) );
  NANDN U1854 ( .A(x[1287]), .B(y[1287]), .Z(n960) );
  NAND U1855 ( .A(n961), .B(n960), .Z(n12427) );
  NANDN U1856 ( .A(y[1285]), .B(x[1285]), .Z(n6366) );
  NANDN U1857 ( .A(x[1286]), .B(y[1286]), .Z(n4564) );
  NANDN U1858 ( .A(n6366), .B(n4564), .Z(n4572) );
  NANDN U1859 ( .A(y[1286]), .B(x[1286]), .Z(n963) );
  NANDN U1860 ( .A(y[1287]), .B(x[1287]), .Z(n962) );
  AND U1861 ( .A(n963), .B(n962), .Z(n12425) );
  ANDN U1862 ( .B(x[1283]), .A(y[1283]), .Z(n8433) );
  NANDN U1863 ( .A(x[1283]), .B(y[1283]), .Z(n8436) );
  NANDN U1864 ( .A(x[1276]), .B(y[1276]), .Z(n8416) );
  IV U1865 ( .A(y[1275]), .Z(n8414) );
  ANDN U1866 ( .B(y[1274]), .A(x[1274]), .Z(n8410) );
  NANDN U1867 ( .A(y[1274]), .B(x[1274]), .Z(n6370) );
  NANDN U1868 ( .A(y[1273]), .B(x[1273]), .Z(n964) );
  AND U1869 ( .A(n6370), .B(n964), .Z(n4539) );
  IV U1870 ( .A(x[1273]), .Z(n6372) );
  IV U1871 ( .A(y[1273]), .Z(n6371) );
  XNOR U1872 ( .A(n6372), .B(n6371), .Z(n4537) );
  NANDN U1873 ( .A(y[1272]), .B(x[1272]), .Z(n6374) );
  NANDN U1874 ( .A(y[1269]), .B(x[1269]), .Z(n8401) );
  IV U1875 ( .A(n8401), .Z(n6379) );
  NANDN U1876 ( .A(x[1267]), .B(y[1267]), .Z(n4518) );
  NANDN U1877 ( .A(x[1266]), .B(y[1266]), .Z(n965) );
  AND U1878 ( .A(n4518), .B(n965), .Z(n971) );
  NANDN U1879 ( .A(x[1264]), .B(y[1264]), .Z(n966) );
  NANDN U1880 ( .A(y[1265]), .B(n966), .Z(n969) );
  XNOR U1881 ( .A(n966), .B(y[1265]), .Z(n967) );
  NAND U1882 ( .A(n967), .B(x[1265]), .Z(n968) );
  NAND U1883 ( .A(n969), .B(n968), .Z(n970) );
  NAND U1884 ( .A(n971), .B(n970), .Z(n12388) );
  NANDN U1885 ( .A(y[1257]), .B(x[1257]), .Z(n12383) );
  ANDN U1886 ( .B(x[1258]), .A(y[1258]), .Z(n8390) );
  ANDN U1887 ( .B(n12383), .A(n8390), .Z(n4490) );
  NANDN U1888 ( .A(y[1256]), .B(x[1256]), .Z(n12379) );
  ANDN U1889 ( .B(x[1255]), .A(y[1255]), .Z(n6384) );
  ANDN U1890 ( .B(n12379), .A(n6384), .Z(n4487) );
  NANDN U1891 ( .A(y[1253]), .B(x[1253]), .Z(n12377) );
  ANDN U1892 ( .B(x[1254]), .A(y[1254]), .Z(n6383) );
  ANDN U1893 ( .B(n12377), .A(n6383), .Z(n4484) );
  NANDN U1894 ( .A(y[1251]), .B(x[1251]), .Z(n973) );
  NANDN U1895 ( .A(y[1250]), .B(x[1250]), .Z(n972) );
  AND U1896 ( .A(n973), .B(n972), .Z(n12373) );
  NANDN U1897 ( .A(x[1250]), .B(y[1250]), .Z(n975) );
  NANDN U1898 ( .A(x[1249]), .B(y[1249]), .Z(n974) );
  NAND U1899 ( .A(n975), .B(n974), .Z(n12372) );
  NANDN U1900 ( .A(y[1249]), .B(x[1249]), .Z(n6385) );
  NANDN U1901 ( .A(x[1248]), .B(y[1248]), .Z(n4476) );
  IV U1902 ( .A(y[1248]), .Z(n6388) );
  IV U1903 ( .A(x[1248]), .Z(n6387) );
  XNOR U1904 ( .A(n6388), .B(n6387), .Z(n4474) );
  NANDN U1905 ( .A(x[1247]), .B(y[1247]), .Z(n6390) );
  ANDN U1906 ( .B(x[1243]), .A(y[1243]), .Z(n8356) );
  NANDN U1907 ( .A(y[1244]), .B(x[1244]), .Z(n12359) );
  NANDN U1908 ( .A(x[1241]), .B(y[1241]), .Z(n4459) );
  NANDN U1909 ( .A(y[1240]), .B(x[1240]), .Z(n12347) );
  ANDN U1910 ( .B(x[1241]), .A(y[1241]), .Z(n12351) );
  ANDN U1911 ( .B(n12347), .A(n12351), .Z(n976) );
  ANDN U1912 ( .B(n4459), .A(n976), .Z(n8353) );
  ANDN U1913 ( .B(x[1242]), .A(y[1242]), .Z(n8355) );
  NOR U1914 ( .A(n8353), .B(n8355), .Z(n4462) );
  NANDN U1915 ( .A(y[1239]), .B(x[1239]), .Z(n978) );
  NANDN U1916 ( .A(y[1238]), .B(x[1238]), .Z(n977) );
  NAND U1917 ( .A(n978), .B(n977), .Z(n12339) );
  NANDN U1918 ( .A(x[1236]), .B(y[1236]), .Z(n4455) );
  IV U1919 ( .A(y[1236]), .Z(n6392) );
  IV U1920 ( .A(x[1236]), .Z(n6391) );
  XNOR U1921 ( .A(n6392), .B(n6391), .Z(n4453) );
  NANDN U1922 ( .A(x[1235]), .B(y[1235]), .Z(n6394) );
  XNOR U1923 ( .A(x[1235]), .B(y[1235]), .Z(n4450) );
  NANDN U1924 ( .A(y[1233]), .B(x[1233]), .Z(n12329) );
  ANDN U1925 ( .B(x[1234]), .A(y[1234]), .Z(n8341) );
  ANDN U1926 ( .B(n12329), .A(n8341), .Z(n4447) );
  ANDN U1927 ( .B(y[1231]), .A(x[1231]), .Z(n12326) );
  ANDN U1928 ( .B(y[1230]), .A(x[1230]), .Z(n8329) );
  NOR U1929 ( .A(n12326), .B(n8329), .Z(n4442) );
  ANDN U1930 ( .B(y[1229]), .A(x[1229]), .Z(n8328) );
  NANDN U1931 ( .A(x[1225]), .B(y[1225]), .Z(n979) );
  ANDN U1932 ( .B(y[1226]), .A(x[1226]), .Z(n4429) );
  ANDN U1933 ( .B(n979), .A(n4429), .Z(n12320) );
  ANDN U1934 ( .B(y[1222]), .A(x[1222]), .Z(n12314) );
  NANDN U1935 ( .A(y[1221]), .B(x[1221]), .Z(n12316) );
  NANDN U1936 ( .A(x[1218]), .B(y[1218]), .Z(n981) );
  NANDN U1937 ( .A(x[1217]), .B(y[1217]), .Z(n980) );
  NAND U1938 ( .A(n981), .B(n980), .Z(n12307) );
  NANDN U1939 ( .A(x[1206]), .B(y[1206]), .Z(n12279) );
  ANDN U1940 ( .B(y[1207]), .A(x[1207]), .Z(n12284) );
  ANDN U1941 ( .B(n12279), .A(n12284), .Z(n4381) );
  NANDN U1942 ( .A(y[1206]), .B(x[1206]), .Z(n6403) );
  NANDN U1943 ( .A(x[1204]), .B(y[1204]), .Z(n983) );
  NANDN U1944 ( .A(x[1203]), .B(y[1203]), .Z(n982) );
  AND U1945 ( .A(n983), .B(n982), .Z(n985) );
  NANDN U1946 ( .A(x[1205]), .B(y[1205]), .Z(n984) );
  NAND U1947 ( .A(n985), .B(n984), .Z(n12276) );
  NANDN U1948 ( .A(x[1202]), .B(y[1202]), .Z(n987) );
  NANDN U1949 ( .A(x[1201]), .B(y[1201]), .Z(n986) );
  NAND U1950 ( .A(n987), .B(n986), .Z(n12272) );
  NANDN U1951 ( .A(x[1199]), .B(y[1199]), .Z(n988) );
  NANDN U1952 ( .A(x[1200]), .B(y[1200]), .Z(n4367) );
  NAND U1953 ( .A(n988), .B(n4367), .Z(n8288) );
  NANDN U1954 ( .A(x[1198]), .B(y[1198]), .Z(n989) );
  NANDN U1955 ( .A(n8288), .B(n989), .Z(n12268) );
  NANDN U1956 ( .A(y[1198]), .B(x[1198]), .Z(n8285) );
  NANDN U1957 ( .A(y[1196]), .B(x[1196]), .Z(n12261) );
  NANDN U1958 ( .A(y[1195]), .B(x[1195]), .Z(n8274) );
  AND U1959 ( .A(n12261), .B(n8274), .Z(n4362) );
  NANDN U1960 ( .A(x[1195]), .B(y[1195]), .Z(n12259) );
  NANDN U1961 ( .A(y[1193]), .B(x[1193]), .Z(n991) );
  NANDN U1962 ( .A(y[1192]), .B(x[1192]), .Z(n990) );
  NAND U1963 ( .A(n991), .B(n990), .Z(n12253) );
  NANDN U1964 ( .A(y[1189]), .B(x[1189]), .Z(n8264) );
  NANDN U1965 ( .A(x[1188]), .B(y[1188]), .Z(n6404) );
  XNOR U1966 ( .A(y[1188]), .B(x[1188]), .Z(n4342) );
  ANDN U1967 ( .B(y[1186]), .A(x[1186]), .Z(n12240) );
  NANDN U1968 ( .A(y[1185]), .B(x[1185]), .Z(n12238) );
  ANDN U1969 ( .B(y[1184]), .A(x[1184]), .Z(n8253) );
  ANDN U1970 ( .B(y[1185]), .A(x[1185]), .Z(n8259) );
  NOR U1971 ( .A(n8253), .B(n8259), .Z(n12235) );
  NANDN U1972 ( .A(x[1183]), .B(y[1183]), .Z(n8254) );
  NANDN U1973 ( .A(x[1182]), .B(y[1182]), .Z(n6409) );
  NANDN U1974 ( .A(y[1183]), .B(x[1183]), .Z(n4327) );
  NANDN U1975 ( .A(n6409), .B(n4327), .Z(n992) );
  NAND U1976 ( .A(n8254), .B(n992), .Z(n12232) );
  IV U1977 ( .A(y[1181]), .Z(n6411) );
  IV U1978 ( .A(x[1181]), .Z(n6410) );
  NANDN U1979 ( .A(n6411), .B(n6410), .Z(n993) );
  NANDN U1980 ( .A(x[1180]), .B(y[1180]), .Z(n8243) );
  NAND U1981 ( .A(n993), .B(n8243), .Z(n12228) );
  NANDN U1982 ( .A(y[1177]), .B(x[1177]), .Z(n995) );
  NANDN U1983 ( .A(y[1176]), .B(x[1176]), .Z(n994) );
  NAND U1984 ( .A(n995), .B(n994), .Z(n12217) );
  NANDN U1985 ( .A(x[1176]), .B(y[1176]), .Z(n6414) );
  NANDN U1986 ( .A(y[1173]), .B(x[1173]), .Z(n12209) );
  NANDN U1987 ( .A(x[1172]), .B(y[1172]), .Z(n8230) );
  NANDN U1988 ( .A(x[1173]), .B(y[1173]), .Z(n8236) );
  NAND U1989 ( .A(n8230), .B(n8236), .Z(n12208) );
  NANDN U1990 ( .A(y[1171]), .B(x[1171]), .Z(n8227) );
  ANDN U1991 ( .B(y[1171]), .A(x[1171]), .Z(n12204) );
  ANDN U1992 ( .B(y[1169]), .A(x[1169]), .Z(n8225) );
  NANDN U1993 ( .A(x[1166]), .B(y[1166]), .Z(n8219) );
  ANDN U1994 ( .B(x[1163]), .A(y[1163]), .Z(n8214) );
  NANDN U1995 ( .A(x[1163]), .B(y[1163]), .Z(n6421) );
  NANDN U1996 ( .A(y[1160]), .B(x[1160]), .Z(n12177) );
  NANDN U1997 ( .A(y[1159]), .B(x[1159]), .Z(n8202) );
  AND U1998 ( .A(n12177), .B(n8202), .Z(n4275) );
  NANDN U1999 ( .A(x[1159]), .B(y[1159]), .Z(n12175) );
  NANDN U2000 ( .A(x[1158]), .B(y[1158]), .Z(n996) );
  AND U2001 ( .A(n12175), .B(n996), .Z(n4273) );
  IV U2002 ( .A(y[1158]), .Z(n6423) );
  IV U2003 ( .A(x[1158]), .Z(n6422) );
  XNOR U2004 ( .A(n6423), .B(n6422), .Z(n4271) );
  NANDN U2005 ( .A(y[1157]), .B(x[1157]), .Z(n9999) );
  ANDN U2006 ( .B(y[1156]), .A(x[1156]), .Z(n12166) );
  NANDN U2007 ( .A(x[1157]), .B(y[1157]), .Z(n6425) );
  ANDN U2008 ( .B(x[1156]), .A(y[1156]), .Z(n9998) );
  NANDN U2009 ( .A(y[1155]), .B(x[1155]), .Z(n998) );
  NANDN U2010 ( .A(y[1154]), .B(x[1154]), .Z(n997) );
  NAND U2011 ( .A(n998), .B(n997), .Z(n12164) );
  NANDN U2012 ( .A(y[1153]), .B(x[1153]), .Z(n6427) );
  NANDN U2013 ( .A(x[1149]), .B(y[1149]), .Z(n8186) );
  ANDN U2014 ( .B(x[1149]), .A(y[1149]), .Z(n4247) );
  NANDN U2015 ( .A(x[1148]), .B(y[1148]), .Z(n8181) );
  OR U2016 ( .A(n4247), .B(n8181), .Z(n999) );
  NAND U2017 ( .A(n8186), .B(n999), .Z(n10000) );
  ANDN U2018 ( .B(y[1145]), .A(x[1145]), .Z(n4241) );
  NANDN U2019 ( .A(x[1144]), .B(y[1144]), .Z(n1000) );
  NANDN U2020 ( .A(n4241), .B(n1000), .Z(n10002) );
  NANDN U2021 ( .A(x[1143]), .B(y[1143]), .Z(n8174) );
  NANDN U2022 ( .A(x[1142]), .B(y[1142]), .Z(n8170) );
  NAND U2023 ( .A(n8174), .B(n8170), .Z(n12146) );
  ANDN U2024 ( .B(x[1142]), .A(y[1142]), .Z(n12145) );
  ANDN U2025 ( .B(x[1141]), .A(y[1141]), .Z(n8166) );
  NOR U2026 ( .A(n12145), .B(n8166), .Z(n4235) );
  NANDN U2027 ( .A(x[1141]), .B(y[1141]), .Z(n12144) );
  NANDN U2028 ( .A(y[1137]), .B(x[1137]), .Z(n12139) );
  NANDN U2029 ( .A(y[1136]), .B(x[1136]), .Z(n12137) );
  IV U2030 ( .A(y[1134]), .Z(n1001) );
  XOR U2031 ( .A(x[1134]), .B(n1001), .Z(n4216) );
  ANDN U2032 ( .B(y[1133]), .A(x[1133]), .Z(n8147) );
  NANDN U2033 ( .A(y[1131]), .B(x[1131]), .Z(n4205) );
  NANDN U2034 ( .A(y[1130]), .B(x[1130]), .Z(n1002) );
  AND U2035 ( .A(n4205), .B(n1002), .Z(n12125) );
  ANDN U2036 ( .B(x[1129]), .A(y[1129]), .Z(n8138) );
  ANDN U2037 ( .B(n12125), .A(n8138), .Z(n4204) );
  NANDN U2038 ( .A(x[1129]), .B(y[1129]), .Z(n8142) );
  NANDN U2039 ( .A(x[1128]), .B(y[1128]), .Z(n1003) );
  AND U2040 ( .A(n8142), .B(n1003), .Z(n4202) );
  IV U2041 ( .A(y[1128]), .Z(n6433) );
  IV U2042 ( .A(x[1128]), .Z(n6432) );
  XNOR U2043 ( .A(n6433), .B(n6432), .Z(n4200) );
  IV U2044 ( .A(y[1127]), .Z(n1004) );
  XOR U2045 ( .A(x[1127]), .B(n1004), .Z(n4197) );
  ANDN U2046 ( .B(x[1126]), .A(y[1126]), .Z(n8134) );
  ANDN U2047 ( .B(x[1125]), .A(y[1125]), .Z(n12114) );
  NOR U2048 ( .A(n8134), .B(n12114), .Z(n4194) );
  ANDN U2049 ( .B(x[1124]), .A(y[1124]), .Z(n8129) );
  NANDN U2050 ( .A(x[1122]), .B(y[1122]), .Z(n1006) );
  NANDN U2051 ( .A(x[1121]), .B(y[1121]), .Z(n1005) );
  NAND U2052 ( .A(n1006), .B(n1005), .Z(n12103) );
  NANDN U2053 ( .A(x[1120]), .B(y[1120]), .Z(n1008) );
  NANDN U2054 ( .A(x[1119]), .B(y[1119]), .Z(n1007) );
  NAND U2055 ( .A(n1008), .B(n1007), .Z(n12100) );
  NANDN U2056 ( .A(y[1118]), .B(x[1118]), .Z(n1010) );
  NANDN U2057 ( .A(y[1119]), .B(x[1119]), .Z(n1009) );
  AND U2058 ( .A(n1010), .B(n1009), .Z(n12097) );
  NANDN U2059 ( .A(y[1116]), .B(x[1116]), .Z(n1012) );
  NANDN U2060 ( .A(y[1117]), .B(x[1117]), .Z(n1011) );
  AND U2061 ( .A(n1012), .B(n1011), .Z(n12093) );
  NANDN U2062 ( .A(x[1116]), .B(y[1116]), .Z(n1013) );
  ANDN U2063 ( .B(x[1115]), .A(y[1115]), .Z(n8115) );
  NAND U2064 ( .A(n1013), .B(n8115), .Z(n4176) );
  NANDN U2065 ( .A(x[1115]), .B(y[1115]), .Z(n1014) );
  AND U2066 ( .A(n1014), .B(n1013), .Z(n12092) );
  NANDN U2067 ( .A(x[1114]), .B(y[1114]), .Z(n1016) );
  NANDN U2068 ( .A(x[1113]), .B(y[1113]), .Z(n1015) );
  NAND U2069 ( .A(n1016), .B(n1015), .Z(n8114) );
  NANDN U2070 ( .A(y[1113]), .B(x[1113]), .Z(n4169) );
  ANDN U2071 ( .B(y[1112]), .A(x[1112]), .Z(n6436) );
  NAND U2072 ( .A(n4169), .B(n6436), .Z(n1017) );
  NANDN U2073 ( .A(n8114), .B(n1017), .Z(n12087) );
  NANDN U2074 ( .A(x[1107]), .B(y[1107]), .Z(n1019) );
  NANDN U2075 ( .A(x[1108]), .B(y[1108]), .Z(n1018) );
  AND U2076 ( .A(n1019), .B(n1018), .Z(n12079) );
  NANDN U2077 ( .A(y[1107]), .B(x[1107]), .Z(n1021) );
  NANDN U2078 ( .A(y[1106]), .B(x[1106]), .Z(n1020) );
  NAND U2079 ( .A(n1021), .B(n1020), .Z(n12078) );
  NANDN U2080 ( .A(x[1103]), .B(y[1103]), .Z(n6439) );
  XNOR U2081 ( .A(x[1103]), .B(y[1103]), .Z(n4146) );
  NANDN U2082 ( .A(y[1101]), .B(x[1101]), .Z(n12065) );
  NANDN U2083 ( .A(x[1101]), .B(y[1101]), .Z(n8094) );
  NANDN U2084 ( .A(x[1100]), .B(y[1100]), .Z(n8089) );
  NAND U2085 ( .A(n8094), .B(n8089), .Z(n12064) );
  NANDN U2086 ( .A(y[1099]), .B(x[1099]), .Z(n6441) );
  NANDN U2087 ( .A(x[1092]), .B(y[1092]), .Z(n4121) );
  IV U2088 ( .A(y[1092]), .Z(n6445) );
  IV U2089 ( .A(x[1092]), .Z(n6444) );
  XNOR U2090 ( .A(n6445), .B(n6444), .Z(n4119) );
  NANDN U2091 ( .A(x[1091]), .B(y[1091]), .Z(n6447) );
  XNOR U2092 ( .A(x[1091]), .B(y[1091]), .Z(n4116) );
  NANDN U2093 ( .A(y[1089]), .B(x[1089]), .Z(n12041) );
  ANDN U2094 ( .B(x[1090]), .A(y[1090]), .Z(n8078) );
  ANDN U2095 ( .B(n12041), .A(n8078), .Z(n4113) );
  NANDN U2096 ( .A(y[1088]), .B(x[1088]), .Z(n12037) );
  ANDN U2097 ( .B(x[1087]), .A(y[1087]), .Z(n8069) );
  ANDN U2098 ( .B(n12037), .A(n8069), .Z(n4110) );
  NANDN U2099 ( .A(x[1086]), .B(y[1086]), .Z(n12031) );
  NANDN U2100 ( .A(y[1082]), .B(x[1082]), .Z(n1023) );
  NANDN U2101 ( .A(y[1083]), .B(x[1083]), .Z(n1022) );
  AND U2102 ( .A(n1023), .B(n1022), .Z(n12025) );
  NANDN U2103 ( .A(x[1082]), .B(y[1082]), .Z(n1025) );
  NANDN U2104 ( .A(x[1081]), .B(y[1081]), .Z(n1024) );
  NAND U2105 ( .A(n1025), .B(n1024), .Z(n12024) );
  NANDN U2106 ( .A(y[1079]), .B(x[1079]), .Z(n8057) );
  NANDN U2107 ( .A(x[1080]), .B(y[1080]), .Z(n1027) );
  NANDN U2108 ( .A(n8057), .B(n1027), .Z(n4093) );
  NANDN U2109 ( .A(x[1079]), .B(y[1079]), .Z(n1026) );
  NAND U2110 ( .A(n1027), .B(n1026), .Z(n8059) );
  NANDN U2111 ( .A(x[1078]), .B(y[1078]), .Z(n1028) );
  NANDN U2112 ( .A(n8059), .B(n1028), .Z(n12020) );
  NANDN U2113 ( .A(x[1076]), .B(y[1076]), .Z(n8048) );
  ANDN U2114 ( .B(y[1077]), .A(x[1077]), .Z(n8055) );
  ANDN U2115 ( .B(n8048), .A(n8055), .Z(n12016) );
  ANDN U2116 ( .B(y[1075]), .A(x[1075]), .Z(n12012) );
  NANDN U2117 ( .A(x[1074]), .B(y[1074]), .Z(n12003) );
  NANDN U2118 ( .A(y[1074]), .B(x[1074]), .Z(n8045) );
  ANDN U2119 ( .B(y[1073]), .A(x[1073]), .Z(n1031) );
  ANDN U2120 ( .B(x[1073]), .A(y[1073]), .Z(n12006) );
  NANDN U2121 ( .A(y[1072]), .B(x[1072]), .Z(n1029) );
  NANDN U2122 ( .A(n12006), .B(n1029), .Z(n11999) );
  NANDN U2123 ( .A(n1031), .B(n11999), .Z(n1033) );
  NANDN U2124 ( .A(x[1072]), .B(y[1072]), .Z(n1030) );
  NANDN U2125 ( .A(n1031), .B(n1030), .Z(n12005) );
  OR U2126 ( .A(n12001), .B(n12005), .Z(n1032) );
  NAND U2127 ( .A(n1033), .B(n1032), .Z(n8042) );
  ANDN U2128 ( .B(n8045), .A(n8042), .Z(n4080) );
  NANDN U2129 ( .A(y[1069]), .B(x[1069]), .Z(n8037) );
  NANDN U2130 ( .A(y[1065]), .B(x[1065]), .Z(n11988) );
  XOR U2131 ( .A(y[1064]), .B(x[1064]), .Z(n4059) );
  NANDN U2132 ( .A(y[1063]), .B(x[1063]), .Z(n8023) );
  IV U2133 ( .A(y[1062]), .Z(n1034) );
  XOR U2134 ( .A(x[1062]), .B(n1034), .Z(n4054) );
  ANDN U2135 ( .B(y[1061]), .A(x[1061]), .Z(n8020) );
  NANDN U2136 ( .A(y[1061]), .B(x[1061]), .Z(n1036) );
  NANDN U2137 ( .A(y[1060]), .B(x[1060]), .Z(n1035) );
  NAND U2138 ( .A(n1036), .B(n1035), .Z(n11976) );
  ANDN U2139 ( .B(y[1058]), .A(x[1058]), .Z(n1040) );
  ANDN U2140 ( .B(x[1057]), .A(y[1057]), .Z(n6454) );
  NANDN U2141 ( .A(n1040), .B(n6454), .Z(n1039) );
  NANDN U2142 ( .A(y[1059]), .B(x[1059]), .Z(n1038) );
  NANDN U2143 ( .A(y[1058]), .B(x[1058]), .Z(n1037) );
  NAND U2144 ( .A(n1038), .B(n1037), .Z(n11972) );
  ANDN U2145 ( .B(n1039), .A(n11972), .Z(n4047) );
  NANDN U2146 ( .A(x[1057]), .B(y[1057]), .Z(n1041) );
  ANDN U2147 ( .B(n1041), .A(n1040), .Z(n11970) );
  NANDN U2148 ( .A(x[1055]), .B(y[1055]), .Z(n6457) );
  XNOR U2149 ( .A(x[1055]), .B(y[1055]), .Z(n4039) );
  ANDN U2150 ( .B(x[1053]), .A(y[1053]), .Z(n11960) );
  ANDN U2151 ( .B(x[1054]), .A(y[1054]), .Z(n8012) );
  NOR U2152 ( .A(n11960), .B(n8012), .Z(n4036) );
  NANDN U2153 ( .A(x[1050]), .B(y[1050]), .Z(n6458) );
  NANDN U2154 ( .A(x[1051]), .B(y[1051]), .Z(n11954) );
  NAND U2155 ( .A(n6458), .B(n11954), .Z(n4031) );
  NANDN U2156 ( .A(x[1046]), .B(y[1046]), .Z(n6460) );
  NANDN U2157 ( .A(y[1045]), .B(x[1045]), .Z(n6462) );
  XNOR U2158 ( .A(x[1045]), .B(y[1045]), .Z(n4016) );
  NANDN U2159 ( .A(y[1044]), .B(x[1044]), .Z(n6463) );
  NANDN U2160 ( .A(y[1043]), .B(x[1043]), .Z(n7990) );
  AND U2161 ( .A(n6463), .B(n7990), .Z(n4013) );
  XNOR U2162 ( .A(x[1043]), .B(y[1043]), .Z(n4011) );
  NANDN U2163 ( .A(x[1042]), .B(y[1042]), .Z(n11933) );
  NANDN U2164 ( .A(x[1041]), .B(y[1041]), .Z(n1043) );
  NANDN U2165 ( .A(x[1040]), .B(y[1040]), .Z(n1042) );
  NAND U2166 ( .A(n1043), .B(n1042), .Z(n11930) );
  NANDN U2167 ( .A(x[1038]), .B(y[1038]), .Z(n1045) );
  NANDN U2168 ( .A(x[1037]), .B(y[1037]), .Z(n1044) );
  AND U2169 ( .A(n1045), .B(n1044), .Z(n1047) );
  NANDN U2170 ( .A(x[1039]), .B(y[1039]), .Z(n1046) );
  NAND U2171 ( .A(n1047), .B(n1046), .Z(n11925) );
  NANDN U2172 ( .A(x[1036]), .B(y[1036]), .Z(n1049) );
  NANDN U2173 ( .A(x[1035]), .B(y[1035]), .Z(n1048) );
  NAND U2174 ( .A(n1049), .B(n1048), .Z(n11922) );
  NANDN U2175 ( .A(y[1034]), .B(x[1034]), .Z(n1051) );
  NANDN U2176 ( .A(y[1035]), .B(x[1035]), .Z(n1050) );
  AND U2177 ( .A(n1051), .B(n1050), .Z(n11919) );
  NANDN U2178 ( .A(x[1034]), .B(y[1034]), .Z(n6465) );
  NANDN U2179 ( .A(y[1032]), .B(x[1032]), .Z(n6467) );
  NANDN U2180 ( .A(y[1031]), .B(x[1031]), .Z(n6468) );
  AND U2181 ( .A(n6467), .B(n6468), .Z(n3986) );
  XNOR U2182 ( .A(x[1031]), .B(y[1031]), .Z(n3984) );
  NANDN U2183 ( .A(x[1030]), .B(y[1030]), .Z(n11909) );
  NANDN U2184 ( .A(y[1029]), .B(x[1029]), .Z(n11908) );
  NANDN U2185 ( .A(x[1028]), .B(y[1028]), .Z(n7968) );
  ANDN U2186 ( .B(y[1029]), .A(x[1029]), .Z(n7974) );
  ANDN U2187 ( .B(n7968), .A(n7974), .Z(n11905) );
  NANDN U2188 ( .A(x[1027]), .B(y[1027]), .Z(n11901) );
  NANDN U2189 ( .A(y[1026]), .B(x[1026]), .Z(n6471) );
  XNOR U2190 ( .A(x[1026]), .B(y[1026]), .Z(n3974) );
  NANDN U2191 ( .A(y[1025]), .B(x[1025]), .Z(n1053) );
  NANDN U2192 ( .A(y[1024]), .B(x[1024]), .Z(n1052) );
  NAND U2193 ( .A(n1053), .B(n1052), .Z(n11896) );
  ANDN U2194 ( .B(x[1023]), .A(y[1023]), .Z(n11891) );
  IV U2195 ( .A(x[1022]), .Z(n11887) );
  OR U2196 ( .A(y[1022]), .B(n11887), .Z(n1054) );
  NANDN U2197 ( .A(n11891), .B(n1054), .Z(n7959) );
  NANDN U2198 ( .A(y[1019]), .B(x[1019]), .Z(n7951) );
  NANDN U2199 ( .A(x[1020]), .B(y[1020]), .Z(n3957) );
  NANDN U2200 ( .A(n7951), .B(n3957), .Z(n3961) );
  NANDN U2201 ( .A(y[1017]), .B(x[1017]), .Z(n11878) );
  NANDN U2202 ( .A(y[1018]), .B(x[1018]), .Z(n7950) );
  AND U2203 ( .A(n11878), .B(n7950), .Z(n3955) );
  NANDN U2204 ( .A(x[1016]), .B(y[1016]), .Z(n1056) );
  NANDN U2205 ( .A(x[1017]), .B(y[1017]), .Z(n1055) );
  NAND U2206 ( .A(n1056), .B(n1055), .Z(n11876) );
  NANDN U2207 ( .A(y[1015]), .B(x[1015]), .Z(n1058) );
  NANDN U2208 ( .A(y[1016]), .B(x[1016]), .Z(n1057) );
  AND U2209 ( .A(n1058), .B(n1057), .Z(n11874) );
  ANDN U2210 ( .B(y[1015]), .A(x[1015]), .Z(n11872) );
  ANDN U2211 ( .B(y[1014]), .A(x[1014]), .Z(n11866) );
  OR U2212 ( .A(n11872), .B(n11866), .Z(n7945) );
  NANDN U2213 ( .A(x[1012]), .B(y[1012]), .Z(n1060) );
  NANDN U2214 ( .A(x[1011]), .B(y[1011]), .Z(n1059) );
  NAND U2215 ( .A(n1060), .B(n1059), .Z(n11863) );
  NANDN U2216 ( .A(y[1010]), .B(x[1010]), .Z(n1062) );
  NANDN U2217 ( .A(y[1011]), .B(x[1011]), .Z(n1061) );
  AND U2218 ( .A(n1062), .B(n1061), .Z(n11860) );
  NANDN U2219 ( .A(x[1010]), .B(y[1010]), .Z(n1064) );
  NANDN U2220 ( .A(x[1009]), .B(y[1009]), .Z(n1063) );
  NAND U2221 ( .A(n1064), .B(n1063), .Z(n11859) );
  ANDN U2222 ( .B(x[1004]), .A(y[1004]), .Z(n11845) );
  NANDN U2223 ( .A(x[1003]), .B(y[1003]), .Z(n1066) );
  NANDN U2224 ( .A(x[1004]), .B(y[1004]), .Z(n1065) );
  NAND U2225 ( .A(n1066), .B(n1065), .Z(n11843) );
  ANDN U2226 ( .B(x[1003]), .A(y[1003]), .Z(n3928) );
  ANDN U2227 ( .B(y[1002]), .A(x[1002]), .Z(n11836) );
  NANDN U2228 ( .A(n3928), .B(n11836), .Z(n1067) );
  NANDN U2229 ( .A(n11843), .B(n1067), .Z(n7924) );
  NANDN U2230 ( .A(y[1000]), .B(x[1000]), .Z(n1069) );
  NANDN U2231 ( .A(y[1001]), .B(x[1001]), .Z(n1068) );
  AND U2232 ( .A(n1069), .B(n1068), .Z(n11834) );
  NANDN U2233 ( .A(x[1000]), .B(y[1000]), .Z(n1071) );
  NANDN U2234 ( .A(x[999]), .B(y[999]), .Z(n1070) );
  NAND U2235 ( .A(n1071), .B(n1070), .Z(n11833) );
  NANDN U2236 ( .A(x[994]), .B(y[994]), .Z(n1073) );
  NANDN U2237 ( .A(x[995]), .B(y[995]), .Z(n1072) );
  NAND U2238 ( .A(n1073), .B(n1072), .Z(n11821) );
  NANDN U2239 ( .A(y[993]), .B(x[993]), .Z(n1075) );
  NANDN U2240 ( .A(y[994]), .B(x[994]), .Z(n1074) );
  AND U2241 ( .A(n1075), .B(n1074), .Z(n11818) );
  NANDN U2242 ( .A(x[993]), .B(y[993]), .Z(n1077) );
  NANDN U2243 ( .A(x[992]), .B(y[992]), .Z(n1076) );
  NAND U2244 ( .A(n1077), .B(n1076), .Z(n11817) );
  NANDN U2245 ( .A(y[991]), .B(x[991]), .Z(n1078) );
  NANDN U2246 ( .A(y[992]), .B(x[992]), .Z(n10005) );
  NAND U2247 ( .A(n1078), .B(n10005), .Z(n1082) );
  ANDN U2248 ( .B(y[990]), .A(x[990]), .Z(n11808) );
  ANDN U2249 ( .B(y[991]), .A(x[991]), .Z(n10004) );
  OR U2250 ( .A(n11808), .B(n10004), .Z(n1079) );
  NANDN U2251 ( .A(n1082), .B(n1079), .Z(n1080) );
  NANDN U2252 ( .A(n11817), .B(n1080), .Z(n7911) );
  NANDN U2253 ( .A(y[990]), .B(x[990]), .Z(n1081) );
  NANDN U2254 ( .A(n1082), .B(n1081), .Z(n11812) );
  NANDN U2255 ( .A(x[988]), .B(y[988]), .Z(n1084) );
  NANDN U2256 ( .A(x[987]), .B(y[987]), .Z(n1083) );
  NAND U2257 ( .A(n1084), .B(n1083), .Z(n11805) );
  NANDN U2258 ( .A(x[986]), .B(y[986]), .Z(n1086) );
  NANDN U2259 ( .A(x[985]), .B(y[985]), .Z(n1085) );
  NAND U2260 ( .A(n1086), .B(n1085), .Z(n11801) );
  NANDN U2261 ( .A(x[984]), .B(y[984]), .Z(n11796) );
  NANDN U2262 ( .A(x[981]), .B(y[981]), .Z(n1088) );
  NANDN U2263 ( .A(x[980]), .B(y[980]), .Z(n1087) );
  NAND U2264 ( .A(n1088), .B(n1087), .Z(n11789) );
  NANDN U2265 ( .A(x[978]), .B(y[978]), .Z(n1090) );
  NANDN U2266 ( .A(x[977]), .B(y[977]), .Z(n1089) );
  AND U2267 ( .A(n1090), .B(n1089), .Z(n1092) );
  NANDN U2268 ( .A(x[979]), .B(y[979]), .Z(n1091) );
  NAND U2269 ( .A(n1092), .B(n1091), .Z(n11785) );
  NANDN U2270 ( .A(x[974]), .B(y[974]), .Z(n1094) );
  NANDN U2271 ( .A(x[973]), .B(y[973]), .Z(n1093) );
  NAND U2272 ( .A(n1094), .B(n1093), .Z(n11777) );
  ANDN U2273 ( .B(y[969]), .A(x[969]), .Z(n11759) );
  NANDN U2274 ( .A(x[968]), .B(y[968]), .Z(n1095) );
  NANDN U2275 ( .A(n11759), .B(n1095), .Z(n7886) );
  NANDN U2276 ( .A(x[966]), .B(y[966]), .Z(n11750) );
  NANDN U2277 ( .A(x[967]), .B(y[967]), .Z(n1096) );
  NAND U2278 ( .A(n11750), .B(n1096), .Z(n7883) );
  NANDN U2279 ( .A(x[965]), .B(y[965]), .Z(n11749) );
  NANDN U2280 ( .A(x[964]), .B(y[964]), .Z(n1098) );
  NANDN U2281 ( .A(x[963]), .B(y[963]), .Z(n1097) );
  NAND U2282 ( .A(n1098), .B(n1097), .Z(n11746) );
  NANDN U2283 ( .A(x[962]), .B(y[962]), .Z(n1100) );
  NANDN U2284 ( .A(x[961]), .B(y[961]), .Z(n1099) );
  NAND U2285 ( .A(n1100), .B(n1099), .Z(n11742) );
  NANDN U2286 ( .A(x[960]), .B(y[960]), .Z(n11737) );
  ANDN U2287 ( .B(y[957]), .A(x[957]), .Z(n11724) );
  NANDN U2288 ( .A(x[956]), .B(y[956]), .Z(n1101) );
  NANDN U2289 ( .A(n11724), .B(n1101), .Z(n7866) );
  NANDN U2290 ( .A(x[952]), .B(y[952]), .Z(n1103) );
  NANDN U2291 ( .A(x[951]), .B(y[951]), .Z(n1102) );
  NAND U2292 ( .A(n1103), .B(n1102), .Z(n11711) );
  IV U2293 ( .A(x[946]), .Z(n6477) );
  IV U2294 ( .A(y[946]), .Z(n6476) );
  NANDN U2295 ( .A(n6477), .B(n6476), .Z(n1104) );
  NANDN U2296 ( .A(y[945]), .B(x[945]), .Z(n7845) );
  NAND U2297 ( .A(n1104), .B(n7845), .Z(n11697) );
  ANDN U2298 ( .B(y[945]), .A(x[945]), .Z(n11695) );
  ANDN U2299 ( .B(y[944]), .A(x[944]), .Z(n6478) );
  NOR U2300 ( .A(n11695), .B(n6478), .Z(n3809) );
  NANDN U2301 ( .A(x[943]), .B(y[943]), .Z(n6479) );
  NANDN U2302 ( .A(x[940]), .B(y[940]), .Z(n1106) );
  NANDN U2303 ( .A(x[939]), .B(y[939]), .Z(n1105) );
  NAND U2304 ( .A(n1106), .B(n1105), .Z(n11681) );
  NANDN U2305 ( .A(x[938]), .B(y[938]), .Z(n1108) );
  NANDN U2306 ( .A(x[937]), .B(y[937]), .Z(n1107) );
  NAND U2307 ( .A(n1108), .B(n1107), .Z(n11677) );
  NANDN U2308 ( .A(x[936]), .B(y[936]), .Z(n11672) );
  NANDN U2309 ( .A(x[935]), .B(y[935]), .Z(n1110) );
  NANDN U2310 ( .A(x[934]), .B(y[934]), .Z(n1109) );
  AND U2311 ( .A(n1110), .B(n1109), .Z(n11668) );
  NANDN U2312 ( .A(y[934]), .B(x[934]), .Z(n1112) );
  NANDN U2313 ( .A(y[933]), .B(x[933]), .Z(n1111) );
  NAND U2314 ( .A(n1112), .B(n1111), .Z(n11667) );
  NANDN U2315 ( .A(y[931]), .B(x[931]), .Z(n1113) );
  NANDN U2316 ( .A(y[932]), .B(x[932]), .Z(n10006) );
  NAND U2317 ( .A(n1113), .B(n10006), .Z(n3781) );
  NANDN U2318 ( .A(y[930]), .B(x[930]), .Z(n1114) );
  NANDN U2319 ( .A(n3781), .B(n1114), .Z(n11660) );
  NANDN U2320 ( .A(y[929]), .B(x[929]), .Z(n1116) );
  NANDN U2321 ( .A(y[928]), .B(x[928]), .Z(n1115) );
  NAND U2322 ( .A(n1116), .B(n1115), .Z(n11654) );
  NANDN U2323 ( .A(x[927]), .B(y[927]), .Z(n1118) );
  NANDN U2324 ( .A(x[928]), .B(y[928]), .Z(n1117) );
  AND U2325 ( .A(n1118), .B(n1117), .Z(n11652) );
  NANDN U2326 ( .A(y[927]), .B(x[927]), .Z(n1120) );
  NANDN U2327 ( .A(y[926]), .B(x[926]), .Z(n1119) );
  NAND U2328 ( .A(n1120), .B(n1119), .Z(n11651) );
  NANDN U2329 ( .A(y[925]), .B(x[925]), .Z(n1122) );
  NANDN U2330 ( .A(y[924]), .B(x[924]), .Z(n1121) );
  NAND U2331 ( .A(n1122), .B(n1121), .Z(n11647) );
  ANDN U2332 ( .B(y[924]), .A(x[924]), .Z(n11645) );
  NANDN U2333 ( .A(y[921]), .B(x[921]), .Z(n7810) );
  IV U2334 ( .A(x[922]), .Z(n6481) );
  NAND U2335 ( .A(n7810), .B(n6480), .Z(n11639) );
  NANDN U2336 ( .A(x[919]), .B(y[919]), .Z(n1124) );
  NANDN U2337 ( .A(x[920]), .B(y[920]), .Z(n1123) );
  NAND U2338 ( .A(n1124), .B(n1123), .Z(n11633) );
  ANDN U2339 ( .B(x[919]), .A(y[919]), .Z(n3760) );
  ANDN U2340 ( .B(y[918]), .A(x[918]), .Z(n11626) );
  NANDN U2341 ( .A(n3760), .B(n11626), .Z(n1125) );
  NANDN U2342 ( .A(n11633), .B(n1125), .Z(n7808) );
  NANDN U2343 ( .A(x[917]), .B(y[917]), .Z(n11627) );
  NANDN U2344 ( .A(x[916]), .B(y[916]), .Z(n1127) );
  NANDN U2345 ( .A(x[915]), .B(y[915]), .Z(n1126) );
  NAND U2346 ( .A(n1127), .B(n1126), .Z(n11623) );
  NANDN U2347 ( .A(x[914]), .B(y[914]), .Z(n1129) );
  NANDN U2348 ( .A(x[913]), .B(y[913]), .Z(n1128) );
  NAND U2349 ( .A(n1129), .B(n1128), .Z(n11619) );
  NANDN U2350 ( .A(x[912]), .B(y[912]), .Z(n11614) );
  NANDN U2351 ( .A(x[910]), .B(y[910]), .Z(n1131) );
  NANDN U2352 ( .A(x[911]), .B(y[911]), .Z(n1130) );
  NAND U2353 ( .A(n1131), .B(n1130), .Z(n11611) );
  NANDN U2354 ( .A(y[910]), .B(x[910]), .Z(n1133) );
  NANDN U2355 ( .A(y[909]), .B(x[909]), .Z(n1132) );
  NAND U2356 ( .A(n1133), .B(n1132), .Z(n11609) );
  NANDN U2357 ( .A(x[905]), .B(y[905]), .Z(n11598) );
  NANDN U2358 ( .A(y[905]), .B(x[905]), .Z(n1135) );
  NANDN U2359 ( .A(y[904]), .B(x[904]), .Z(n1134) );
  NAND U2360 ( .A(n1135), .B(n1134), .Z(n11595) );
  NANDN U2361 ( .A(y[903]), .B(x[903]), .Z(n1137) );
  NANDN U2362 ( .A(y[902]), .B(x[902]), .Z(n1136) );
  NAND U2363 ( .A(n1137), .B(n1136), .Z(n11591) );
  NANDN U2364 ( .A(y[901]), .B(x[901]), .Z(n1139) );
  NANDN U2365 ( .A(y[900]), .B(x[900]), .Z(n1138) );
  NAND U2366 ( .A(n1139), .B(n1138), .Z(n11587) );
  NANDN U2367 ( .A(x[900]), .B(y[900]), .Z(n11584) );
  NANDN U2368 ( .A(x[898]), .B(y[898]), .Z(n1141) );
  NANDN U2369 ( .A(x[899]), .B(y[899]), .Z(n1140) );
  NAND U2370 ( .A(n1141), .B(n1140), .Z(n11581) );
  ANDN U2371 ( .B(y[897]), .A(x[897]), .Z(n11576) );
  IV U2372 ( .A(y[896]), .Z(n11571) );
  OR U2373 ( .A(x[896]), .B(n11571), .Z(n1142) );
  NANDN U2374 ( .A(n11576), .B(n1142), .Z(n7782) );
  NANDN U2375 ( .A(x[892]), .B(y[892]), .Z(n1144) );
  NANDN U2376 ( .A(x[891]), .B(y[891]), .Z(n1143) );
  NAND U2377 ( .A(n1144), .B(n1143), .Z(n11558) );
  NANDN U2378 ( .A(x[886]), .B(y[886]), .Z(n1146) );
  NANDN U2379 ( .A(x[887]), .B(y[887]), .Z(n1145) );
  NAND U2380 ( .A(n1146), .B(n1145), .Z(n11546) );
  NANDN U2381 ( .A(x[885]), .B(y[885]), .Z(n1148) );
  NANDN U2382 ( .A(x[884]), .B(y[884]), .Z(n1147) );
  NAND U2383 ( .A(n1148), .B(n1147), .Z(n11541) );
  NANDN U2384 ( .A(y[883]), .B(x[883]), .Z(n1149) );
  NANDN U2385 ( .A(y[884]), .B(x[884]), .Z(n11538) );
  NAND U2386 ( .A(n1149), .B(n11538), .Z(n1153) );
  ANDN U2387 ( .B(y[882]), .A(x[882]), .Z(n11534) );
  ANDN U2388 ( .B(y[883]), .A(x[883]), .Z(n11537) );
  OR U2389 ( .A(n11534), .B(n11537), .Z(n1150) );
  NANDN U2390 ( .A(n1153), .B(n1150), .Z(n1151) );
  NANDN U2391 ( .A(n11541), .B(n1151), .Z(n7766) );
  NANDN U2392 ( .A(y[882]), .B(x[882]), .Z(n1152) );
  NANDN U2393 ( .A(n1153), .B(n1152), .Z(n11536) );
  NANDN U2394 ( .A(y[880]), .B(x[880]), .Z(n1155) );
  NANDN U2395 ( .A(y[881]), .B(x[881]), .Z(n1154) );
  AND U2396 ( .A(n1155), .B(n1154), .Z(n11529) );
  NANDN U2397 ( .A(x[880]), .B(y[880]), .Z(n1157) );
  NANDN U2398 ( .A(x[879]), .B(y[879]), .Z(n1156) );
  NAND U2399 ( .A(n1157), .B(n1156), .Z(n11528) );
  NANDN U2400 ( .A(x[878]), .B(y[878]), .Z(n1159) );
  NANDN U2401 ( .A(x[877]), .B(y[877]), .Z(n1158) );
  NAND U2402 ( .A(n1159), .B(n1158), .Z(n11524) );
  NANDN U2403 ( .A(y[875]), .B(x[875]), .Z(n11517) );
  NANDN U2404 ( .A(y[873]), .B(x[873]), .Z(n7748) );
  IV U2405 ( .A(x[874]), .Z(n6484) );
  IV U2406 ( .A(y[874]), .Z(n6483) );
  NANDN U2407 ( .A(n6484), .B(n6483), .Z(n1160) );
  NAND U2408 ( .A(n7748), .B(n1160), .Z(n11514) );
  NANDN U2409 ( .A(y[870]), .B(x[870]), .Z(n1161) );
  ANDN U2410 ( .B(x[871]), .A(y[871]), .Z(n3671) );
  ANDN U2411 ( .B(n1161), .A(n3671), .Z(n11505) );
  NANDN U2412 ( .A(x[868]), .B(y[868]), .Z(n1163) );
  NANDN U2413 ( .A(x[867]), .B(y[867]), .Z(n1162) );
  NAND U2414 ( .A(n1163), .B(n1162), .Z(n11498) );
  NANDN U2415 ( .A(x[866]), .B(y[866]), .Z(n1165) );
  NANDN U2416 ( .A(x[865]), .B(y[865]), .Z(n1164) );
  NAND U2417 ( .A(n1165), .B(n1164), .Z(n11494) );
  NANDN U2418 ( .A(y[864]), .B(x[864]), .Z(n1167) );
  NANDN U2419 ( .A(y[865]), .B(x[865]), .Z(n1166) );
  AND U2420 ( .A(n1167), .B(n1166), .Z(n11492) );
  NANDN U2421 ( .A(y[861]), .B(x[861]), .Z(n7728) );
  IV U2422 ( .A(x[862]), .Z(n6487) );
  IV U2423 ( .A(y[862]), .Z(n6486) );
  NANDN U2424 ( .A(n6487), .B(n6486), .Z(n1168) );
  NAND U2425 ( .A(n7728), .B(n1168), .Z(n11484) );
  NANDN U2426 ( .A(y[860]), .B(x[860]), .Z(n11480) );
  NANDN U2427 ( .A(x[859]), .B(y[859]), .Z(n1170) );
  NANDN U2428 ( .A(x[860]), .B(y[860]), .Z(n1169) );
  NAND U2429 ( .A(n1170), .B(n1169), .Z(n11478) );
  ANDN U2430 ( .B(x[859]), .A(y[859]), .Z(n3647) );
  ANDN U2431 ( .B(y[858]), .A(x[858]), .Z(n11474) );
  NANDN U2432 ( .A(n3647), .B(n11474), .Z(n1171) );
  NANDN U2433 ( .A(n11478), .B(n1171), .Z(n7726) );
  NANDN U2434 ( .A(x[856]), .B(y[856]), .Z(n1173) );
  NANDN U2435 ( .A(x[855]), .B(y[855]), .Z(n1172) );
  NAND U2436 ( .A(n1173), .B(n1172), .Z(n11468) );
  NANDN U2437 ( .A(y[854]), .B(x[854]), .Z(n1175) );
  NANDN U2438 ( .A(y[855]), .B(x[855]), .Z(n1174) );
  AND U2439 ( .A(n1175), .B(n1174), .Z(n11465) );
  NANDN U2440 ( .A(x[854]), .B(y[854]), .Z(n1177) );
  NANDN U2441 ( .A(x[853]), .B(y[853]), .Z(n1176) );
  NAND U2442 ( .A(n1177), .B(n1176), .Z(n11464) );
  NANDN U2443 ( .A(x[846]), .B(y[846]), .Z(n1179) );
  NANDN U2444 ( .A(x[845]), .B(y[845]), .Z(n1178) );
  NAND U2445 ( .A(n1179), .B(n1178), .Z(n11448) );
  NANDN U2446 ( .A(x[844]), .B(y[844]), .Z(n1181) );
  NANDN U2447 ( .A(x[843]), .B(y[843]), .Z(n1180) );
  NAND U2448 ( .A(n1181), .B(n1180), .Z(n11444) );
  NANDN U2449 ( .A(y[842]), .B(x[842]), .Z(n1183) );
  NANDN U2450 ( .A(y[843]), .B(x[843]), .Z(n1182) );
  AND U2451 ( .A(n1183), .B(n1182), .Z(n11441) );
  ANDN U2452 ( .B(y[842]), .A(x[842]), .Z(n11440) );
  NANDN U2453 ( .A(x[841]), .B(y[841]), .Z(n11434) );
  NANDN U2454 ( .A(n11440), .B(n11434), .Z(n7698) );
  NANDN U2455 ( .A(x[839]), .B(y[839]), .Z(n1185) );
  NANDN U2456 ( .A(x[838]), .B(y[838]), .Z(n1184) );
  NAND U2457 ( .A(n1185), .B(n1184), .Z(n11430) );
  NANDN U2458 ( .A(y[837]), .B(x[837]), .Z(n1187) );
  NANDN U2459 ( .A(y[838]), .B(x[838]), .Z(n1186) );
  AND U2460 ( .A(n1187), .B(n1186), .Z(n11427) );
  NANDN U2461 ( .A(y[836]), .B(x[836]), .Z(n1188) );
  NANDN U2462 ( .A(y[835]), .B(x[835]), .Z(n7685) );
  NAND U2463 ( .A(n1188), .B(n7685), .Z(n11424) );
  NANDN U2464 ( .A(x[835]), .B(y[835]), .Z(n6492) );
  NANDN U2465 ( .A(x[834]), .B(y[834]), .Z(n6491) );
  NAND U2466 ( .A(n6492), .B(n6491), .Z(n11421) );
  NANDN U2467 ( .A(y[834]), .B(x[834]), .Z(n1189) );
  NANDN U2468 ( .A(y[833]), .B(x[833]), .Z(n7680) );
  NAND U2469 ( .A(n1189), .B(n7680), .Z(n11419) );
  ANDN U2470 ( .B(y[829]), .A(x[829]), .Z(n7669) );
  ANDN U2471 ( .B(x[827]), .A(y[827]), .Z(n7660) );
  NANDN U2472 ( .A(y[826]), .B(x[826]), .Z(n1190) );
  NANDN U2473 ( .A(n7660), .B(n1190), .Z(n11408) );
  NANDN U2474 ( .A(y[822]), .B(x[822]), .Z(n1192) );
  NANDN U2475 ( .A(y[821]), .B(x[821]), .Z(n1191) );
  AND U2476 ( .A(n1192), .B(n1191), .Z(n1194) );
  NANDN U2477 ( .A(y[823]), .B(x[823]), .Z(n1193) );
  NAND U2478 ( .A(n1194), .B(n1193), .Z(n11400) );
  ANDN U2479 ( .B(y[821]), .A(x[821]), .Z(n3578) );
  ANDN U2480 ( .B(x[820]), .A(y[820]), .Z(n11396) );
  NANDN U2481 ( .A(n3578), .B(n11396), .Z(n1195) );
  NANDN U2482 ( .A(n11400), .B(n1195), .Z(n7654) );
  NANDN U2483 ( .A(y[819]), .B(x[819]), .Z(n11397) );
  NANDN U2484 ( .A(x[818]), .B(y[818]), .Z(n7646) );
  NANDN U2485 ( .A(x[819]), .B(y[819]), .Z(n7650) );
  NAND U2486 ( .A(n7646), .B(n7650), .Z(n11395) );
  NANDN U2487 ( .A(y[816]), .B(x[816]), .Z(n1197) );
  NANDN U2488 ( .A(y[817]), .B(x[817]), .Z(n1196) );
  NAND U2489 ( .A(n1197), .B(n1196), .Z(n11392) );
  ANDN U2490 ( .B(y[813]), .A(x[813]), .Z(n3563) );
  NANDN U2491 ( .A(x[812]), .B(y[812]), .Z(n1198) );
  NANDN U2492 ( .A(n3563), .B(n1198), .Z(n10009) );
  NANDN U2493 ( .A(y[811]), .B(x[811]), .Z(n11389) );
  NANDN U2494 ( .A(x[810]), .B(y[810]), .Z(n6498) );
  XNOR U2495 ( .A(y[810]), .B(x[810]), .Z(n3555) );
  NANDN U2496 ( .A(y[809]), .B(x[809]), .Z(n6499) );
  NANDN U2497 ( .A(y[808]), .B(x[808]), .Z(n1200) );
  NANDN U2498 ( .A(y[807]), .B(x[807]), .Z(n1199) );
  NAND U2499 ( .A(n1200), .B(n1199), .Z(n11384) );
  NANDN U2500 ( .A(y[804]), .B(x[804]), .Z(n1202) );
  NANDN U2501 ( .A(y[803]), .B(x[803]), .Z(n1201) );
  NAND U2502 ( .A(n1202), .B(n1201), .Z(n11378) );
  NANDN U2503 ( .A(y[802]), .B(x[802]), .Z(n1204) );
  NANDN U2504 ( .A(y[801]), .B(x[801]), .Z(n1203) );
  NAND U2505 ( .A(n1204), .B(n1203), .Z(n11373) );
  ANDN U2506 ( .B(y[801]), .A(x[801]), .Z(n3532) );
  ANDN U2507 ( .B(x[800]), .A(y[800]), .Z(n11367) );
  NANDN U2508 ( .A(n3532), .B(n11367), .Z(n1205) );
  NANDN U2509 ( .A(n11373), .B(n1205), .Z(n7629) );
  NANDN U2510 ( .A(x[799]), .B(y[799]), .Z(n7623) );
  NANDN U2511 ( .A(x[798]), .B(y[798]), .Z(n1206) );
  NAND U2512 ( .A(n7623), .B(n1206), .Z(n11366) );
  ANDN U2513 ( .B(x[797]), .A(y[797]), .Z(n11361) );
  ANDN U2514 ( .B(y[797]), .A(x[797]), .Z(n3525) );
  ANDN U2515 ( .B(x[796]), .A(y[796]), .Z(n11355) );
  NANDN U2516 ( .A(n3525), .B(n11355), .Z(n1207) );
  NANDN U2517 ( .A(n11361), .B(n1207), .Z(n7621) );
  NANDN U2518 ( .A(x[794]), .B(y[794]), .Z(n1208) );
  ANDN U2519 ( .B(y[795]), .A(x[795]), .Z(n7618) );
  ANDN U2520 ( .B(n1208), .A(n7618), .Z(n11353) );
  NANDN U2521 ( .A(y[793]), .B(x[793]), .Z(n7609) );
  IV U2522 ( .A(x[794]), .Z(n7614) );
  OR U2523 ( .A(y[794]), .B(n7614), .Z(n1209) );
  NAND U2524 ( .A(n7609), .B(n1209), .Z(n11352) );
  NANDN U2525 ( .A(x[793]), .B(y[793]), .Z(n3521) );
  NANDN U2526 ( .A(x[791]), .B(y[791]), .Z(n1211) );
  NANDN U2527 ( .A(x[790]), .B(y[790]), .Z(n1210) );
  NAND U2528 ( .A(n1211), .B(n1210), .Z(n11343) );
  NANDN U2529 ( .A(y[784]), .B(x[784]), .Z(n1213) );
  NANDN U2530 ( .A(y[783]), .B(x[783]), .Z(n1212) );
  AND U2531 ( .A(n1213), .B(n1212), .Z(n1215) );
  NANDN U2532 ( .A(y[785]), .B(x[785]), .Z(n1214) );
  AND U2533 ( .A(n1215), .B(n1214), .Z(n11329) );
  NANDN U2534 ( .A(x[783]), .B(y[783]), .Z(n1217) );
  NANDN U2535 ( .A(x[782]), .B(y[782]), .Z(n1216) );
  NAND U2536 ( .A(n1217), .B(n1216), .Z(n11328) );
  NANDN U2537 ( .A(x[780]), .B(y[780]), .Z(n1218) );
  ANDN U2538 ( .B(y[781]), .A(x[781]), .Z(n3494) );
  ANDN U2539 ( .B(n1218), .A(n3494), .Z(n11323) );
  NANDN U2540 ( .A(x[777]), .B(y[777]), .Z(n1223) );
  XNOR U2541 ( .A(x[777]), .B(y[777]), .Z(n1220) );
  NANDN U2542 ( .A(y[776]), .B(x[776]), .Z(n1219) );
  NAND U2543 ( .A(n1220), .B(n1219), .Z(n1221) );
  AND U2544 ( .A(n1223), .B(n1221), .Z(n11313) );
  NANDN U2545 ( .A(x[776]), .B(y[776]), .Z(n1222) );
  AND U2546 ( .A(n1223), .B(n1222), .Z(n1229) );
  NANDN U2547 ( .A(x[774]), .B(y[774]), .Z(n1224) );
  NANDN U2548 ( .A(y[775]), .B(n1224), .Z(n1227) );
  XNOR U2549 ( .A(n1224), .B(y[775]), .Z(n1225) );
  NAND U2550 ( .A(n1225), .B(x[775]), .Z(n1226) );
  NAND U2551 ( .A(n1227), .B(n1226), .Z(n1228) );
  NAND U2552 ( .A(n1229), .B(n1228), .Z(n11312) );
  NANDN U2553 ( .A(y[774]), .B(x[774]), .Z(n1231) );
  NANDN U2554 ( .A(y[773]), .B(x[773]), .Z(n1230) );
  AND U2555 ( .A(n1231), .B(n1230), .Z(n1233) );
  NANDN U2556 ( .A(y[775]), .B(x[775]), .Z(n1232) );
  NAND U2557 ( .A(n1233), .B(n1232), .Z(n11309) );
  ANDN U2558 ( .B(y[773]), .A(x[773]), .Z(n3480) );
  ANDN U2559 ( .B(x[772]), .A(y[772]), .Z(n11306) );
  NANDN U2560 ( .A(n3480), .B(n11306), .Z(n1234) );
  NANDN U2561 ( .A(n11309), .B(n1234), .Z(n7587) );
  NANDN U2562 ( .A(x[768]), .B(y[768]), .Z(n1236) );
  NANDN U2563 ( .A(x[767]), .B(y[767]), .Z(n1235) );
  AND U2564 ( .A(n1236), .B(n1235), .Z(n1238) );
  NANDN U2565 ( .A(x[769]), .B(y[769]), .Z(n1237) );
  NAND U2566 ( .A(n1238), .B(n1237), .Z(n11296) );
  NANDN U2567 ( .A(y[767]), .B(x[767]), .Z(n1240) );
  NANDN U2568 ( .A(y[766]), .B(x[766]), .Z(n1239) );
  NAND U2569 ( .A(n1240), .B(n1239), .Z(n11294) );
  NANDN U2570 ( .A(y[765]), .B(x[765]), .Z(n1242) );
  NANDN U2571 ( .A(y[764]), .B(x[764]), .Z(n1241) );
  NAND U2572 ( .A(n1242), .B(n1241), .Z(n11290) );
  ANDN U2573 ( .B(x[760]), .A(y[760]), .Z(n11282) );
  ANDN U2574 ( .B(y[759]), .A(x[759]), .Z(n3449) );
  NANDN U2575 ( .A(y[758]), .B(x[758]), .Z(n1243) );
  NANDN U2576 ( .A(y[759]), .B(x[759]), .Z(n11277) );
  NAND U2577 ( .A(n1243), .B(n11277), .Z(n11273) );
  NANDN U2578 ( .A(n3449), .B(n11273), .Z(n1244) );
  NANDN U2579 ( .A(n11282), .B(n1244), .Z(n7572) );
  NANDN U2580 ( .A(x[757]), .B(y[757]), .Z(n1250) );
  XNOR U2581 ( .A(x[757]), .B(y[757]), .Z(n1246) );
  NANDN U2582 ( .A(y[756]), .B(x[756]), .Z(n1245) );
  NAND U2583 ( .A(n1246), .B(n1245), .Z(n1247) );
  AND U2584 ( .A(n1250), .B(n1247), .Z(n11276) );
  NANDN U2585 ( .A(x[754]), .B(y[754]), .Z(n7565) );
  NANDN U2586 ( .A(y[755]), .B(x[755]), .Z(n3445) );
  NANDN U2587 ( .A(n7565), .B(n3445), .Z(n1252) );
  NANDN U2588 ( .A(x[756]), .B(y[756]), .Z(n1249) );
  NANDN U2589 ( .A(x[755]), .B(y[755]), .Z(n1248) );
  AND U2590 ( .A(n1249), .B(n1248), .Z(n1251) );
  AND U2591 ( .A(n1251), .B(n1250), .Z(n7568) );
  NAND U2592 ( .A(n1252), .B(n7568), .Z(n11272) );
  ANDN U2593 ( .B(x[753]), .A(y[753]), .Z(n7563) );
  ANDN U2594 ( .B(x[749]), .A(y[749]), .Z(n1258) );
  NANDN U2595 ( .A(x[748]), .B(y[748]), .Z(n7553) );
  OR U2596 ( .A(n1258), .B(n7553), .Z(n1256) );
  NANDN U2597 ( .A(x[750]), .B(y[750]), .Z(n1254) );
  NANDN U2598 ( .A(x[749]), .B(y[749]), .Z(n1253) );
  AND U2599 ( .A(n1254), .B(n1253), .Z(n1255) );
  NANDN U2600 ( .A(x[751]), .B(y[751]), .Z(n3438) );
  AND U2601 ( .A(n1255), .B(n3438), .Z(n7557) );
  NAND U2602 ( .A(n1256), .B(n7557), .Z(n11263) );
  NANDN U2603 ( .A(y[748]), .B(x[748]), .Z(n1257) );
  NANDN U2604 ( .A(n1258), .B(n1257), .Z(n11262) );
  ANDN U2605 ( .B(x[747]), .A(y[747]), .Z(n10011) );
  NANDN U2606 ( .A(y[746]), .B(x[746]), .Z(n10012) );
  NANDN U2607 ( .A(n10011), .B(n10012), .Z(n7551) );
  NANDN U2608 ( .A(x[742]), .B(y[742]), .Z(n7542) );
  NANDN U2609 ( .A(y[743]), .B(x[743]), .Z(n1263) );
  NANDN U2610 ( .A(n7542), .B(n1263), .Z(n1261) );
  NANDN U2611 ( .A(x[743]), .B(y[743]), .Z(n1260) );
  NANDN U2612 ( .A(x[744]), .B(y[744]), .Z(n1259) );
  AND U2613 ( .A(n1260), .B(n1259), .Z(n7545) );
  NAND U2614 ( .A(n1261), .B(n7545), .Z(n11247) );
  NANDN U2615 ( .A(y[742]), .B(x[742]), .Z(n1262) );
  NAND U2616 ( .A(n1263), .B(n1262), .Z(n11245) );
  NANDN U2617 ( .A(y[740]), .B(x[740]), .Z(n1265) );
  NANDN U2618 ( .A(y[741]), .B(x[741]), .Z(n1264) );
  NAND U2619 ( .A(n1265), .B(n1264), .Z(n11242) );
  NANDN U2620 ( .A(x[737]), .B(y[737]), .Z(n1269) );
  XNOR U2621 ( .A(x[737]), .B(y[737]), .Z(n1267) );
  NANDN U2622 ( .A(y[736]), .B(x[736]), .Z(n1266) );
  NAND U2623 ( .A(n1267), .B(n1266), .Z(n1268) );
  AND U2624 ( .A(n1269), .B(n1268), .Z(n11231) );
  NANDN U2625 ( .A(y[734]), .B(x[734]), .Z(n1271) );
  NANDN U2626 ( .A(y[733]), .B(x[733]), .Z(n1270) );
  AND U2627 ( .A(n1271), .B(n1270), .Z(n1273) );
  NANDN U2628 ( .A(y[735]), .B(x[735]), .Z(n1272) );
  NAND U2629 ( .A(n1273), .B(n1272), .Z(n11228) );
  ANDN U2630 ( .B(y[733]), .A(x[733]), .Z(n3411) );
  ANDN U2631 ( .B(x[732]), .A(y[732]), .Z(n11224) );
  NANDN U2632 ( .A(n3411), .B(n11224), .Z(n1274) );
  NANDN U2633 ( .A(n11228), .B(n1274), .Z(n7533) );
  NANDN U2634 ( .A(y[730]), .B(x[730]), .Z(n1280) );
  ANDN U2635 ( .B(x[728]), .A(y[728]), .Z(n1275) );
  OR U2636 ( .A(n1275), .B(x[729]), .Z(n1278) );
  XOR U2637 ( .A(x[729]), .B(n1275), .Z(n1276) );
  NAND U2638 ( .A(n1276), .B(y[729]), .Z(n1277) );
  NAND U2639 ( .A(n1278), .B(n1277), .Z(n1279) );
  NAND U2640 ( .A(n1280), .B(n1279), .Z(n11218) );
  NANDN U2641 ( .A(y[727]), .B(x[727]), .Z(n1282) );
  NANDN U2642 ( .A(y[726]), .B(x[726]), .Z(n1281) );
  NAND U2643 ( .A(n1282), .B(n1281), .Z(n11213) );
  NANDN U2644 ( .A(y[724]), .B(x[724]), .Z(n1283) );
  ANDN U2645 ( .B(x[725]), .A(y[725]), .Z(n11212) );
  ANDN U2646 ( .B(n1283), .A(n11212), .Z(n1284) );
  NANDN U2647 ( .A(x[725]), .B(y[725]), .Z(n1286) );
  NANDN U2648 ( .A(n1284), .B(n1286), .Z(n1285) );
  NANDN U2649 ( .A(n11213), .B(n1285), .Z(n7526) );
  NANDN U2650 ( .A(x[723]), .B(y[723]), .Z(n1288) );
  NANDN U2651 ( .A(x[722]), .B(y[722]), .Z(n1287) );
  NAND U2652 ( .A(n1288), .B(n1287), .Z(n11204) );
  NANDN U2653 ( .A(y[722]), .B(x[722]), .Z(n1290) );
  NANDN U2654 ( .A(y[721]), .B(x[721]), .Z(n1289) );
  NAND U2655 ( .A(n1290), .B(n1289), .Z(n11202) );
  ANDN U2656 ( .B(y[721]), .A(x[721]), .Z(n3389) );
  ANDN U2657 ( .B(x[720]), .A(y[720]), .Z(n11198) );
  NANDN U2658 ( .A(n3389), .B(n11198), .Z(n1291) );
  NANDN U2659 ( .A(n11202), .B(n1291), .Z(n7521) );
  NANDN U2660 ( .A(y[717]), .B(x[717]), .Z(n11190) );
  NANDN U2661 ( .A(y[715]), .B(x[715]), .Z(n1293) );
  NANDN U2662 ( .A(y[716]), .B(x[716]), .Z(n1292) );
  AND U2663 ( .A(n1293), .B(n1292), .Z(n11185) );
  NANDN U2664 ( .A(x[715]), .B(y[715]), .Z(n1295) );
  NANDN U2665 ( .A(x[714]), .B(y[714]), .Z(n1294) );
  NAND U2666 ( .A(n1295), .B(n1294), .Z(n11184) );
  NANDN U2667 ( .A(y[711]), .B(x[711]), .Z(n11175) );
  NANDN U2668 ( .A(x[706]), .B(y[706]), .Z(n1296) );
  ANDN U2669 ( .B(y[707]), .A(x[707]), .Z(n3361) );
  ANDN U2670 ( .B(n1296), .A(n3361), .Z(n11161) );
  NANDN U2671 ( .A(x[705]), .B(y[705]), .Z(n1298) );
  NANDN U2672 ( .A(x[704]), .B(y[704]), .Z(n1297) );
  NAND U2673 ( .A(n1298), .B(n1297), .Z(n11156) );
  NANDN U2674 ( .A(x[703]), .B(y[703]), .Z(n1300) );
  NANDN U2675 ( .A(x[702]), .B(y[702]), .Z(n1299) );
  NAND U2676 ( .A(n1300), .B(n1299), .Z(n11152) );
  NANDN U2677 ( .A(x[695]), .B(y[695]), .Z(n1302) );
  NANDN U2678 ( .A(x[694]), .B(y[694]), .Z(n1301) );
  NAND U2679 ( .A(n1302), .B(n1301), .Z(n11144) );
  NANDN U2680 ( .A(x[691]), .B(y[691]), .Z(n1304) );
  NANDN U2681 ( .A(x[690]), .B(y[690]), .Z(n1303) );
  NAND U2682 ( .A(n1304), .B(n1303), .Z(n7483) );
  NANDN U2683 ( .A(x[688]), .B(y[688]), .Z(n7477) );
  ANDN U2684 ( .B(y[689]), .A(x[689]), .Z(n7480) );
  ANDN U2685 ( .B(n7477), .A(n7480), .Z(n1305) );
  NANDN U2686 ( .A(y[689]), .B(x[689]), .Z(n3315) );
  NANDN U2687 ( .A(n1305), .B(n3315), .Z(n1306) );
  NANDN U2688 ( .A(n7483), .B(n1306), .Z(n11140) );
  NANDN U2689 ( .A(x[686]), .B(y[686]), .Z(n1307) );
  ANDN U2690 ( .B(y[687]), .A(x[687]), .Z(n3316) );
  ANDN U2691 ( .B(n1307), .A(n3316), .Z(n7474) );
  AND U2692 ( .A(n7474), .B(n11135), .Z(n3313) );
  NANDN U2693 ( .A(y[684]), .B(x[684]), .Z(n1309) );
  NANDN U2694 ( .A(y[683]), .B(x[683]), .Z(n1308) );
  AND U2695 ( .A(n1309), .B(n1308), .Z(n1311) );
  NANDN U2696 ( .A(y[685]), .B(x[685]), .Z(n1310) );
  NAND U2697 ( .A(n1311), .B(n1310), .Z(n11134) );
  ANDN U2698 ( .B(y[683]), .A(x[683]), .Z(n3305) );
  ANDN U2699 ( .B(x[682]), .A(y[682]), .Z(n11132) );
  NANDN U2700 ( .A(n3305), .B(n11132), .Z(n1312) );
  NANDN U2701 ( .A(n11134), .B(n1312), .Z(n7471) );
  NANDN U2702 ( .A(x[677]), .B(y[677]), .Z(n1314) );
  NANDN U2703 ( .A(x[676]), .B(y[676]), .Z(n1313) );
  NAND U2704 ( .A(n1314), .B(n1313), .Z(n11126) );
  NANDN U2705 ( .A(x[674]), .B(y[674]), .Z(n1315) );
  NANDN U2706 ( .A(x[675]), .B(y[675]), .Z(n7461) );
  NAND U2707 ( .A(n1315), .B(n7461), .Z(n11124) );
  NANDN U2708 ( .A(x[669]), .B(y[669]), .Z(n1316) );
  NANDN U2709 ( .A(y[668]), .B(x[668]), .Z(n10015) );
  ANDN U2710 ( .B(n1316), .A(n10015), .Z(n6509) );
  NANDN U2711 ( .A(y[670]), .B(x[670]), .Z(n7446) );
  ANDN U2712 ( .B(x[669]), .A(y[669]), .Z(n6510) );
  ANDN U2713 ( .B(n7446), .A(n6510), .Z(n11118) );
  NANDN U2714 ( .A(x[668]), .B(y[668]), .Z(n1317) );
  AND U2715 ( .A(n1317), .B(n1316), .Z(n11116) );
  NANDN U2716 ( .A(x[665]), .B(y[665]), .Z(n3266) );
  XNOR U2717 ( .A(x[665]), .B(y[665]), .Z(n1319) );
  NANDN U2718 ( .A(y[664]), .B(x[664]), .Z(n1318) );
  NAND U2719 ( .A(n1319), .B(n1318), .Z(n1320) );
  AND U2720 ( .A(n3266), .B(n1320), .Z(n11112) );
  NANDN U2721 ( .A(x[660]), .B(y[660]), .Z(n1321) );
  ANDN U2722 ( .B(y[661]), .A(x[661]), .Z(n3262) );
  ANDN U2723 ( .B(n1321), .A(n3262), .Z(n11109) );
  ANDN U2724 ( .B(x[659]), .A(y[659]), .Z(n11108) );
  ANDN U2725 ( .B(y[659]), .A(x[659]), .Z(n3253) );
  ANDN U2726 ( .B(x[658]), .A(y[658]), .Z(n11104) );
  NANDN U2727 ( .A(n3253), .B(n11104), .Z(n1322) );
  NANDN U2728 ( .A(n11108), .B(n1322), .Z(n7432) );
  NANDN U2729 ( .A(x[657]), .B(y[657]), .Z(n1324) );
  NANDN U2730 ( .A(x[656]), .B(y[656]), .Z(n1323) );
  NAND U2731 ( .A(n1324), .B(n1323), .Z(n11103) );
  NANDN U2732 ( .A(y[652]), .B(x[652]), .Z(n1326) );
  NANDN U2733 ( .A(y[651]), .B(x[651]), .Z(n1325) );
  AND U2734 ( .A(n1326), .B(n1325), .Z(n1328) );
  NANDN U2735 ( .A(y[653]), .B(x[653]), .Z(n1327) );
  NAND U2736 ( .A(n1328), .B(n1327), .Z(n11100) );
  ANDN U2737 ( .B(y[651]), .A(x[651]), .Z(n3239) );
  ANDN U2738 ( .B(x[650]), .A(y[650]), .Z(n11096) );
  NANDN U2739 ( .A(n3239), .B(n11096), .Z(n1329) );
  NANDN U2740 ( .A(n11100), .B(n1329), .Z(n7425) );
  NANDN U2741 ( .A(x[649]), .B(y[649]), .Z(n3236) );
  NANDN U2742 ( .A(x[648]), .B(y[648]), .Z(n1330) );
  NAND U2743 ( .A(n3236), .B(n1330), .Z(n11095) );
  NANDN U2744 ( .A(x[647]), .B(y[647]), .Z(n1332) );
  NANDN U2745 ( .A(x[646]), .B(y[646]), .Z(n1331) );
  NAND U2746 ( .A(n1332), .B(n1331), .Z(n11094) );
  NANDN U2747 ( .A(y[646]), .B(x[646]), .Z(n1334) );
  NANDN U2748 ( .A(y[645]), .B(x[645]), .Z(n1333) );
  NAND U2749 ( .A(n1334), .B(n1333), .Z(n11093) );
  ANDN U2750 ( .B(y[645]), .A(x[645]), .Z(n3229) );
  ANDN U2751 ( .B(x[644]), .A(y[644]), .Z(n11090) );
  NANDN U2752 ( .A(n3229), .B(n11090), .Z(n1335) );
  NANDN U2753 ( .A(n11093), .B(n1335), .Z(n7417) );
  NANDN U2754 ( .A(x[643]), .B(y[643]), .Z(n7414) );
  NANDN U2755 ( .A(x[642]), .B(y[642]), .Z(n1336) );
  NAND U2756 ( .A(n7414), .B(n1336), .Z(n11089) );
  NANDN U2757 ( .A(x[641]), .B(y[641]), .Z(n3218) );
  XNOR U2758 ( .A(x[641]), .B(y[641]), .Z(n1338) );
  NANDN U2759 ( .A(y[640]), .B(x[640]), .Z(n1337) );
  NAND U2760 ( .A(n1338), .B(n1337), .Z(n1339) );
  AND U2761 ( .A(n3218), .B(n1339), .Z(n7407) );
  NANDN U2762 ( .A(y[642]), .B(x[642]), .Z(n1340) );
  NANDN U2763 ( .A(n7407), .B(n1340), .Z(n11088) );
  NANDN U2764 ( .A(y[639]), .B(x[639]), .Z(n1342) );
  NANDN U2765 ( .A(y[638]), .B(x[638]), .Z(n1341) );
  AND U2766 ( .A(n1342), .B(n1341), .Z(n1348) );
  NANDN U2767 ( .A(y[636]), .B(x[636]), .Z(n1343) );
  NANDN U2768 ( .A(x[637]), .B(n1343), .Z(n1346) );
  XNOR U2769 ( .A(n1343), .B(x[637]), .Z(n1344) );
  NAND U2770 ( .A(n1344), .B(y[637]), .Z(n1345) );
  NAND U2771 ( .A(n1346), .B(n1345), .Z(n1347) );
  NAND U2772 ( .A(n1348), .B(n1347), .Z(n11086) );
  NANDN U2773 ( .A(x[637]), .B(y[637]), .Z(n1350) );
  NANDN U2774 ( .A(x[636]), .B(y[636]), .Z(n1349) );
  AND U2775 ( .A(n1350), .B(n1349), .Z(n1356) );
  NANDN U2776 ( .A(x[634]), .B(y[634]), .Z(n1351) );
  NANDN U2777 ( .A(y[635]), .B(n1351), .Z(n1354) );
  XNOR U2778 ( .A(n1351), .B(y[635]), .Z(n1352) );
  NAND U2779 ( .A(n1352), .B(x[635]), .Z(n1353) );
  NAND U2780 ( .A(n1354), .B(n1353), .Z(n1355) );
  NAND U2781 ( .A(n1356), .B(n1355), .Z(n11085) );
  NANDN U2782 ( .A(x[633]), .B(y[633]), .Z(n3206) );
  NANDN U2783 ( .A(y[631]), .B(x[631]), .Z(n3198) );
  ANDN U2784 ( .B(n3198), .A(x[630]), .Z(n1357) );
  NAND U2785 ( .A(n1357), .B(y[630]), .Z(n1359) );
  NANDN U2786 ( .A(x[631]), .B(y[631]), .Z(n1358) );
  AND U2787 ( .A(n1359), .B(n1358), .Z(n1360) );
  AND U2788 ( .A(n3206), .B(n1360), .Z(n1362) );
  NANDN U2789 ( .A(x[632]), .B(y[632]), .Z(n1361) );
  NAND U2790 ( .A(n1362), .B(n1361), .Z(n11083) );
  NANDN U2791 ( .A(x[623]), .B(y[623]), .Z(n1364) );
  NANDN U2792 ( .A(x[622]), .B(y[622]), .Z(n1363) );
  NAND U2793 ( .A(n1364), .B(n1363), .Z(n6516) );
  ANDN U2794 ( .B(x[621]), .A(y[621]), .Z(n6514) );
  NANDN U2795 ( .A(y[619]), .B(x[619]), .Z(n1366) );
  NANDN U2796 ( .A(y[618]), .B(x[618]), .Z(n1365) );
  AND U2797 ( .A(n1366), .B(n1365), .Z(n1372) );
  NANDN U2798 ( .A(y[616]), .B(x[616]), .Z(n1367) );
  NANDN U2799 ( .A(x[617]), .B(n1367), .Z(n1370) );
  XNOR U2800 ( .A(n1367), .B(x[617]), .Z(n1368) );
  NAND U2801 ( .A(n1368), .B(y[617]), .Z(n1369) );
  NAND U2802 ( .A(n1370), .B(n1369), .Z(n1371) );
  NAND U2803 ( .A(n1372), .B(n1371), .Z(n11064) );
  NANDN U2804 ( .A(x[614]), .B(y[614]), .Z(n7386) );
  NANDN U2805 ( .A(y[615]), .B(x[615]), .Z(n1379) );
  NANDN U2806 ( .A(n7386), .B(n1379), .Z(n1377) );
  NANDN U2807 ( .A(x[616]), .B(y[616]), .Z(n1374) );
  NANDN U2808 ( .A(x[615]), .B(y[615]), .Z(n1373) );
  AND U2809 ( .A(n1374), .B(n1373), .Z(n1376) );
  NANDN U2810 ( .A(x[617]), .B(y[617]), .Z(n1375) );
  AND U2811 ( .A(n1376), .B(n1375), .Z(n7389) );
  NAND U2812 ( .A(n1377), .B(n7389), .Z(n11062) );
  NANDN U2813 ( .A(y[614]), .B(x[614]), .Z(n1378) );
  NAND U2814 ( .A(n1379), .B(n1378), .Z(n11060) );
  NANDN U2815 ( .A(x[610]), .B(y[610]), .Z(n1380) );
  ANDN U2816 ( .B(y[611]), .A(x[611]), .Z(n3164) );
  ANDN U2817 ( .B(n1380), .A(n3164), .Z(n11053) );
  NANDN U2818 ( .A(x[609]), .B(y[609]), .Z(n7381) );
  NANDN U2819 ( .A(x[608]), .B(y[608]), .Z(n7376) );
  NANDN U2820 ( .A(y[609]), .B(x[609]), .Z(n1383) );
  NANDN U2821 ( .A(n7376), .B(n1383), .Z(n1381) );
  NAND U2822 ( .A(n7381), .B(n1381), .Z(n11050) );
  ANDN U2823 ( .B(n11053), .A(n11050), .Z(n3159) );
  NANDN U2824 ( .A(y[608]), .B(x[608]), .Z(n1382) );
  NAND U2825 ( .A(n1383), .B(n1382), .Z(n11048) );
  NANDN U2826 ( .A(y[605]), .B(x[605]), .Z(n1385) );
  NANDN U2827 ( .A(y[604]), .B(x[604]), .Z(n1384) );
  AND U2828 ( .A(n1385), .B(n1384), .Z(n1391) );
  NANDN U2829 ( .A(y[602]), .B(x[602]), .Z(n1386) );
  NANDN U2830 ( .A(x[603]), .B(n1386), .Z(n1389) );
  XNOR U2831 ( .A(n1386), .B(x[603]), .Z(n1387) );
  NAND U2832 ( .A(n1387), .B(y[603]), .Z(n1388) );
  NAND U2833 ( .A(n1389), .B(n1388), .Z(n1390) );
  NAND U2834 ( .A(n1391), .B(n1390), .Z(n11040) );
  ANDN U2835 ( .B(x[597]), .A(y[597]), .Z(n3131) );
  NANDN U2836 ( .A(x[596]), .B(y[596]), .Z(n6518) );
  OR U2837 ( .A(n3131), .B(n6518), .Z(n1396) );
  NANDN U2838 ( .A(x[598]), .B(y[598]), .Z(n1393) );
  NANDN U2839 ( .A(x[597]), .B(y[597]), .Z(n1392) );
  AND U2840 ( .A(n1393), .B(n1392), .Z(n1395) );
  NANDN U2841 ( .A(x[599]), .B(y[599]), .Z(n1394) );
  AND U2842 ( .A(n1395), .B(n1394), .Z(n7369) );
  NAND U2843 ( .A(n1396), .B(n7369), .Z(n11033) );
  IV U2844 ( .A(y[595]), .Z(n6520) );
  IV U2845 ( .A(x[595]), .Z(n6519) );
  NANDN U2846 ( .A(n6520), .B(n6519), .Z(n1398) );
  NANDN U2847 ( .A(x[594]), .B(y[594]), .Z(n1397) );
  NAND U2848 ( .A(n1398), .B(n1397), .Z(n11030) );
  NANDN U2849 ( .A(x[593]), .B(y[593]), .Z(n3123) );
  ANDN U2850 ( .B(x[592]), .A(y[592]), .Z(n11024) );
  NAND U2851 ( .A(n3123), .B(n11024), .Z(n6522) );
  NANDN U2852 ( .A(y[591]), .B(x[591]), .Z(n1400) );
  NANDN U2853 ( .A(y[590]), .B(x[590]), .Z(n1399) );
  NAND U2854 ( .A(n1400), .B(n1399), .Z(n11016) );
  NANDN U2855 ( .A(y[589]), .B(x[589]), .Z(n1402) );
  NANDN U2856 ( .A(y[588]), .B(x[588]), .Z(n1401) );
  NAND U2857 ( .A(n1402), .B(n1401), .Z(n11012) );
  ANDN U2858 ( .B(y[585]), .A(x[585]), .Z(n3110) );
  NANDN U2859 ( .A(x[584]), .B(y[584]), .Z(n1403) );
  NANDN U2860 ( .A(n3110), .B(n1403), .Z(n10018) );
  NANDN U2861 ( .A(x[581]), .B(y[581]), .Z(n3099) );
  NANDN U2862 ( .A(y[580]), .B(x[580]), .Z(n1404) );
  ANDN U2863 ( .B(x[581]), .A(y[581]), .Z(n10996) );
  ANDN U2864 ( .B(n1404), .A(n10996), .Z(n1405) );
  ANDN U2865 ( .B(n3099), .A(n1405), .Z(n7342) );
  NANDN U2866 ( .A(y[579]), .B(x[579]), .Z(n10989) );
  NANDN U2867 ( .A(x[579]), .B(y[579]), .Z(n1407) );
  NANDN U2868 ( .A(x[578]), .B(y[578]), .Z(n1406) );
  NAND U2869 ( .A(n1407), .B(n1406), .Z(n10988) );
  NANDN U2870 ( .A(y[574]), .B(x[574]), .Z(n1409) );
  NANDN U2871 ( .A(y[573]), .B(x[573]), .Z(n1408) );
  AND U2872 ( .A(n1409), .B(n1408), .Z(n1411) );
  NANDN U2873 ( .A(y[575]), .B(x[575]), .Z(n1410) );
  NAND U2874 ( .A(n1411), .B(n1410), .Z(n10981) );
  ANDN U2875 ( .B(y[573]), .A(x[573]), .Z(n3085) );
  ANDN U2876 ( .B(x[572]), .A(y[572]), .Z(n10975) );
  NANDN U2877 ( .A(n3085), .B(n10975), .Z(n1412) );
  NANDN U2878 ( .A(n10981), .B(n1412), .Z(n7336) );
  NANDN U2879 ( .A(y[571]), .B(x[571]), .Z(n10976) );
  NANDN U2880 ( .A(x[569]), .B(y[569]), .Z(n1419) );
  XNOR U2881 ( .A(x[569]), .B(y[569]), .Z(n1414) );
  NANDN U2882 ( .A(y[568]), .B(x[568]), .Z(n1413) );
  NAND U2883 ( .A(n1414), .B(n1413), .Z(n1415) );
  AND U2884 ( .A(n1419), .B(n1415), .Z(n7326) );
  NANDN U2885 ( .A(y[570]), .B(x[570]), .Z(n1416) );
  NANDN U2886 ( .A(n7326), .B(n1416), .Z(n10972) );
  NANDN U2887 ( .A(x[566]), .B(y[566]), .Z(n7320) );
  NANDN U2888 ( .A(y[567]), .B(x[567]), .Z(n3077) );
  NANDN U2889 ( .A(n7320), .B(n3077), .Z(n1421) );
  NANDN U2890 ( .A(x[568]), .B(y[568]), .Z(n1418) );
  NANDN U2891 ( .A(x[567]), .B(y[567]), .Z(n1417) );
  AND U2892 ( .A(n1418), .B(n1417), .Z(n1420) );
  AND U2893 ( .A(n1420), .B(n1419), .Z(n7323) );
  NAND U2894 ( .A(n1421), .B(n7323), .Z(n10970) );
  NANDN U2895 ( .A(y[561]), .B(x[561]), .Z(n1423) );
  NANDN U2896 ( .A(y[560]), .B(x[560]), .Z(n1422) );
  AND U2897 ( .A(n1423), .B(n1422), .Z(n1429) );
  NANDN U2898 ( .A(y[558]), .B(x[558]), .Z(n1424) );
  NANDN U2899 ( .A(x[559]), .B(n1424), .Z(n1427) );
  XNOR U2900 ( .A(n1424), .B(x[559]), .Z(n1425) );
  NAND U2901 ( .A(n1425), .B(y[559]), .Z(n1426) );
  NAND U2902 ( .A(n1427), .B(n1426), .Z(n1428) );
  NAND U2903 ( .A(n1429), .B(n1428), .Z(n10963) );
  NANDN U2904 ( .A(y[556]), .B(x[556]), .Z(n1431) );
  NANDN U2905 ( .A(y[555]), .B(x[555]), .Z(n1430) );
  AND U2906 ( .A(n1431), .B(n1430), .Z(n1433) );
  NANDN U2907 ( .A(y[557]), .B(x[557]), .Z(n1432) );
  NAND U2908 ( .A(n1433), .B(n1432), .Z(n10961) );
  ANDN U2909 ( .B(y[555]), .A(x[555]), .Z(n3051) );
  ANDN U2910 ( .B(x[554]), .A(y[554]), .Z(n10958) );
  NANDN U2911 ( .A(n3051), .B(n10958), .Z(n1434) );
  NANDN U2912 ( .A(n10961), .B(n1434), .Z(n7314) );
  NANDN U2913 ( .A(y[553]), .B(x[553]), .Z(n10959) );
  NANDN U2914 ( .A(x[553]), .B(y[553]), .Z(n1436) );
  NANDN U2915 ( .A(x[552]), .B(y[552]), .Z(n1435) );
  NAND U2916 ( .A(n1436), .B(n1435), .Z(n10957) );
  ANDN U2917 ( .B(x[552]), .A(y[552]), .Z(n10956) );
  ANDN U2918 ( .B(y[551]), .A(x[551]), .Z(n1440) );
  NANDN U2919 ( .A(y[550]), .B(x[550]), .Z(n1437) );
  NANDN U2920 ( .A(y[551]), .B(x[551]), .Z(n10021) );
  NAND U2921 ( .A(n1437), .B(n10021), .Z(n10022) );
  NANDN U2922 ( .A(n1440), .B(n10022), .Z(n1438) );
  NANDN U2923 ( .A(n10956), .B(n1438), .Z(n7309) );
  NANDN U2924 ( .A(x[550]), .B(y[550]), .Z(n1439) );
  NANDN U2925 ( .A(n1440), .B(n1439), .Z(n10020) );
  NANDN U2926 ( .A(x[549]), .B(y[549]), .Z(n1442) );
  NANDN U2927 ( .A(x[548]), .B(y[548]), .Z(n1441) );
  NAND U2928 ( .A(n1442), .B(n1441), .Z(n10955) );
  NANDN U2929 ( .A(y[548]), .B(x[548]), .Z(n10954) );
  NANDN U2930 ( .A(x[547]), .B(y[547]), .Z(n7302) );
  NANDN U2931 ( .A(x[546]), .B(y[546]), .Z(n7296) );
  NANDN U2932 ( .A(y[547]), .B(x[547]), .Z(n3038) );
  NANDN U2933 ( .A(n7296), .B(n3038), .Z(n1443) );
  NAND U2934 ( .A(n7302), .B(n1443), .Z(n10953) );
  NANDN U2935 ( .A(y[542]), .B(x[542]), .Z(n1444) );
  NANDN U2936 ( .A(y[543]), .B(x[543]), .Z(n3031) );
  NAND U2937 ( .A(n1444), .B(n3031), .Z(n7291) );
  ANDN U2938 ( .B(y[541]), .A(x[541]), .Z(n6523) );
  NANDN U2939 ( .A(y[541]), .B(x[541]), .Z(n1446) );
  NANDN U2940 ( .A(y[540]), .B(x[540]), .Z(n1445) );
  AND U2941 ( .A(n1446), .B(n1445), .Z(n7286) );
  OR U2942 ( .A(n6523), .B(n7286), .Z(n1447) );
  NANDN U2943 ( .A(n7291), .B(n1447), .Z(n10948) );
  NANDN U2944 ( .A(x[537]), .B(y[537]), .Z(n1449) );
  NANDN U2945 ( .A(x[536]), .B(y[536]), .Z(n1448) );
  NAND U2946 ( .A(n1449), .B(n1448), .Z(n10942) );
  NANDN U2947 ( .A(y[535]), .B(x[535]), .Z(n1451) );
  NANDN U2948 ( .A(y[536]), .B(x[536]), .Z(n1450) );
  AND U2949 ( .A(n1451), .B(n1450), .Z(n10939) );
  NANDN U2950 ( .A(x[535]), .B(y[535]), .Z(n1453) );
  NANDN U2951 ( .A(x[534]), .B(y[534]), .Z(n1452) );
  NAND U2952 ( .A(n1453), .B(n1452), .Z(n10938) );
  ANDN U2953 ( .B(x[534]), .A(y[534]), .Z(n10936) );
  NANDN U2954 ( .A(y[532]), .B(x[532]), .Z(n1454) );
  ANDN U2955 ( .B(x[533]), .A(y[533]), .Z(n10934) );
  ANDN U2956 ( .B(n1454), .A(n10934), .Z(n1455) );
  NANDN U2957 ( .A(x[533]), .B(y[533]), .Z(n1457) );
  NANDN U2958 ( .A(n1455), .B(n1457), .Z(n1456) );
  NANDN U2959 ( .A(n10936), .B(n1456), .Z(n7279) );
  ANDN U2960 ( .B(x[523]), .A(y[523]), .Z(n1460) );
  NANDN U2961 ( .A(x[523]), .B(y[523]), .Z(n7270) );
  NANDN U2962 ( .A(x[522]), .B(y[522]), .Z(n1458) );
  AND U2963 ( .A(n7270), .B(n1458), .Z(n1459) );
  OR U2964 ( .A(n1460), .B(n1459), .Z(n10918) );
  ANDN U2965 ( .B(x[521]), .A(y[521]), .Z(n7264) );
  NOR U2966 ( .A(n7264), .B(n7269), .Z(n10915) );
  NANDN U2967 ( .A(y[520]), .B(x[520]), .Z(n1462) );
  NANDN U2968 ( .A(y[519]), .B(x[519]), .Z(n1461) );
  NAND U2969 ( .A(n1462), .B(n1461), .Z(n10912) );
  NANDN U2970 ( .A(y[518]), .B(x[518]), .Z(n1464) );
  NANDN U2971 ( .A(y[517]), .B(x[517]), .Z(n1463) );
  NAND U2972 ( .A(n1464), .B(n1463), .Z(n10908) );
  ANDN U2973 ( .B(y[517]), .A(x[517]), .Z(n2982) );
  ANDN U2974 ( .B(x[516]), .A(y[516]), .Z(n10901) );
  NANDN U2975 ( .A(n2982), .B(n10901), .Z(n1465) );
  NANDN U2976 ( .A(n10908), .B(n1465), .Z(n7260) );
  NANDN U2977 ( .A(x[515]), .B(y[515]), .Z(n2979) );
  NANDN U2978 ( .A(x[514]), .B(y[514]), .Z(n1466) );
  NAND U2979 ( .A(n2979), .B(n1466), .Z(n10899) );
  NANDN U2980 ( .A(x[513]), .B(y[513]), .Z(n6530) );
  NANDN U2981 ( .A(y[513]), .B(x[513]), .Z(n10896) );
  NANDN U2982 ( .A(y[512]), .B(x[512]), .Z(n10891) );
  AND U2983 ( .A(n10896), .B(n10891), .Z(n2976) );
  NANDN U2984 ( .A(x[512]), .B(y[512]), .Z(n6529) );
  NANDN U2985 ( .A(x[510]), .B(y[510]), .Z(n1472) );
  ANDN U2986 ( .B(y[508]), .A(x[508]), .Z(n1467) );
  OR U2987 ( .A(n1467), .B(y[509]), .Z(n1470) );
  XOR U2988 ( .A(y[509]), .B(n1467), .Z(n1468) );
  NAND U2989 ( .A(n1468), .B(x[509]), .Z(n1469) );
  NAND U2990 ( .A(n1470), .B(n1469), .Z(n1471) );
  NAND U2991 ( .A(n1472), .B(n1471), .Z(n10886) );
  NANDN U2992 ( .A(y[509]), .B(x[509]), .Z(n1474) );
  NANDN U2993 ( .A(y[508]), .B(x[508]), .Z(n1473) );
  NAND U2994 ( .A(n1474), .B(n1473), .Z(n10883) );
  NANDN U2995 ( .A(y[506]), .B(x[506]), .Z(n1475) );
  ANDN U2996 ( .B(x[507]), .A(y[507]), .Z(n10882) );
  ANDN U2997 ( .B(n1475), .A(n10882), .Z(n1476) );
  NANDN U2998 ( .A(x[507]), .B(y[507]), .Z(n1478) );
  NANDN U2999 ( .A(n1476), .B(n1478), .Z(n1477) );
  NANDN U3000 ( .A(n10883), .B(n1477), .Z(n7248) );
  NANDN U3001 ( .A(x[503]), .B(y[503]), .Z(n1480) );
  NANDN U3002 ( .A(x[502]), .B(y[502]), .Z(n1479) );
  NAND U3003 ( .A(n1480), .B(n1479), .Z(n10869) );
  ANDN U3004 ( .B(x[502]), .A(y[502]), .Z(n10868) );
  ANDN U3005 ( .B(y[501]), .A(x[501]), .Z(n2955) );
  NANDN U3006 ( .A(y[500]), .B(x[500]), .Z(n1481) );
  NANDN U3007 ( .A(y[501]), .B(x[501]), .Z(n10863) );
  NAND U3008 ( .A(n1481), .B(n10863), .Z(n10859) );
  NANDN U3009 ( .A(n2955), .B(n10859), .Z(n1482) );
  NANDN U3010 ( .A(n10868), .B(n1482), .Z(n7241) );
  NANDN U3011 ( .A(y[497]), .B(x[497]), .Z(n1484) );
  NANDN U3012 ( .A(y[496]), .B(x[496]), .Z(n1483) );
  AND U3013 ( .A(n1484), .B(n1483), .Z(n1490) );
  NANDN U3014 ( .A(y[494]), .B(x[494]), .Z(n1485) );
  NANDN U3015 ( .A(x[495]), .B(n1485), .Z(n1488) );
  XNOR U3016 ( .A(n1485), .B(x[495]), .Z(n1486) );
  NAND U3017 ( .A(n1486), .B(y[495]), .Z(n1487) );
  NAND U3018 ( .A(n1488), .B(n1487), .Z(n1489) );
  NAND U3019 ( .A(n1490), .B(n1489), .Z(n10856) );
  NANDN U3020 ( .A(y[492]), .B(x[492]), .Z(n1492) );
  NANDN U3021 ( .A(y[491]), .B(x[491]), .Z(n1491) );
  AND U3022 ( .A(n1492), .B(n1491), .Z(n1494) );
  NANDN U3023 ( .A(y[493]), .B(x[493]), .Z(n1493) );
  NAND U3024 ( .A(n1494), .B(n1493), .Z(n10852) );
  ANDN U3025 ( .B(y[491]), .A(x[491]), .Z(n2939) );
  ANDN U3026 ( .B(x[490]), .A(y[490]), .Z(n10845) );
  NANDN U3027 ( .A(n2939), .B(n10845), .Z(n1495) );
  NANDN U3028 ( .A(n10852), .B(n1495), .Z(n7234) );
  NANDN U3029 ( .A(x[485]), .B(y[485]), .Z(n1497) );
  NANDN U3030 ( .A(x[484]), .B(y[484]), .Z(n1496) );
  AND U3031 ( .A(n1497), .B(n1496), .Z(n1504) );
  NANDN U3032 ( .A(y[484]), .B(x[484]), .Z(n1506) );
  ANDN U3033 ( .B(y[482]), .A(x[482]), .Z(n1499) );
  OR U3034 ( .A(n1499), .B(y[483]), .Z(n1498) );
  AND U3035 ( .A(n1506), .B(n1498), .Z(n1502) );
  XOR U3036 ( .A(y[483]), .B(n1499), .Z(n1500) );
  NAND U3037 ( .A(n1500), .B(x[483]), .Z(n1501) );
  NAND U3038 ( .A(n1502), .B(n1501), .Z(n1503) );
  NAND U3039 ( .A(n1504), .B(n1503), .Z(n10840) );
  NANDN U3040 ( .A(y[483]), .B(x[483]), .Z(n1505) );
  AND U3041 ( .A(n1506), .B(n1505), .Z(n1508) );
  NANDN U3042 ( .A(y[482]), .B(x[482]), .Z(n1507) );
  NAND U3043 ( .A(n1508), .B(n1507), .Z(n10838) );
  NANDN U3044 ( .A(y[480]), .B(x[480]), .Z(n10831) );
  ANDN U3045 ( .B(x[481]), .A(y[481]), .Z(n10835) );
  ANDN U3046 ( .B(n10831), .A(n10835), .Z(n1509) );
  NANDN U3047 ( .A(x[481]), .B(y[481]), .Z(n1511) );
  NANDN U3048 ( .A(n1509), .B(n1511), .Z(n1510) );
  NANDN U3049 ( .A(n10838), .B(n1510), .Z(n7227) );
  NANDN U3050 ( .A(y[479]), .B(x[479]), .Z(n2913) );
  XNOR U3051 ( .A(y[479]), .B(x[479]), .Z(n1513) );
  NANDN U3052 ( .A(x[478]), .B(y[478]), .Z(n1512) );
  NAND U3053 ( .A(n1513), .B(n1512), .Z(n1514) );
  AND U3054 ( .A(n2913), .B(n1514), .Z(n10830) );
  OR U3055 ( .A(n10834), .B(n10830), .Z(n7225) );
  NANDN U3056 ( .A(y[475]), .B(x[475]), .Z(n1516) );
  NANDN U3057 ( .A(y[474]), .B(x[474]), .Z(n1515) );
  AND U3058 ( .A(n1516), .B(n1515), .Z(n1523) );
  NANDN U3059 ( .A(y[472]), .B(x[472]), .Z(n1518) );
  NANDN U3060 ( .A(x[473]), .B(n1518), .Z(n1521) );
  IV U3061 ( .A(x[473]), .Z(n1517) );
  XOR U3062 ( .A(n1518), .B(n1517), .Z(n1519) );
  NAND U3063 ( .A(n1519), .B(y[473]), .Z(n1520) );
  NAND U3064 ( .A(n1521), .B(n1520), .Z(n1522) );
  NAND U3065 ( .A(n1523), .B(n1522), .Z(n10823) );
  NANDN U3066 ( .A(x[473]), .B(y[473]), .Z(n1525) );
  NANDN U3067 ( .A(x[472]), .B(y[472]), .Z(n1524) );
  AND U3068 ( .A(n1525), .B(n1524), .Z(n1531) );
  NANDN U3069 ( .A(x[470]), .B(y[470]), .Z(n1526) );
  NANDN U3070 ( .A(y[471]), .B(n1526), .Z(n1529) );
  XNOR U3071 ( .A(n1526), .B(y[471]), .Z(n1527) );
  NAND U3072 ( .A(n1527), .B(x[471]), .Z(n1528) );
  NAND U3073 ( .A(n1529), .B(n1528), .Z(n1530) );
  NAND U3074 ( .A(n1531), .B(n1530), .Z(n10822) );
  NANDN U3075 ( .A(x[468]), .B(y[468]), .Z(n1533) );
  NANDN U3076 ( .A(x[467]), .B(y[467]), .Z(n1532) );
  AND U3077 ( .A(n1533), .B(n1532), .Z(n1535) );
  NANDN U3078 ( .A(x[469]), .B(y[469]), .Z(n1534) );
  NAND U3079 ( .A(n1535), .B(n1534), .Z(n10818) );
  NANDN U3080 ( .A(x[466]), .B(y[466]), .Z(n1537) );
  NANDN U3081 ( .A(x[465]), .B(y[465]), .Z(n1536) );
  NAND U3082 ( .A(n1537), .B(n1536), .Z(n7216) );
  NANDN U3083 ( .A(y[465]), .B(x[465]), .Z(n2901) );
  ANDN U3084 ( .B(y[464]), .A(x[464]), .Z(n6531) );
  NAND U3085 ( .A(n2901), .B(n6531), .Z(n1538) );
  NANDN U3086 ( .A(n7216), .B(n1538), .Z(n10814) );
  NANDN U3087 ( .A(y[463]), .B(x[463]), .Z(n1542) );
  XNOR U3088 ( .A(y[463]), .B(x[463]), .Z(n1540) );
  NANDN U3089 ( .A(x[462]), .B(y[462]), .Z(n1539) );
  NAND U3090 ( .A(n1540), .B(n1539), .Z(n1541) );
  AND U3091 ( .A(n1542), .B(n1541), .Z(n10810) );
  NANDN U3092 ( .A(x[461]), .B(y[461]), .Z(n1547) );
  NANDN U3093 ( .A(y[459]), .B(x[459]), .Z(n1550) );
  NAND U3094 ( .A(n1550), .B(y[458]), .Z(n1543) );
  OR U3095 ( .A(x[458]), .B(n1543), .Z(n1545) );
  NANDN U3096 ( .A(x[459]), .B(y[459]), .Z(n1544) );
  AND U3097 ( .A(n1545), .B(n1544), .Z(n1546) );
  AND U3098 ( .A(n1547), .B(n1546), .Z(n1549) );
  NANDN U3099 ( .A(x[460]), .B(y[460]), .Z(n1548) );
  NAND U3100 ( .A(n1549), .B(n1548), .Z(n10806) );
  NANDN U3101 ( .A(y[458]), .B(x[458]), .Z(n1551) );
  NAND U3102 ( .A(n1551), .B(n1550), .Z(n10804) );
  NANDN U3103 ( .A(y[456]), .B(x[456]), .Z(n10797) );
  ANDN U3104 ( .B(x[457]), .A(y[457]), .Z(n10801) );
  ANDN U3105 ( .B(n10797), .A(n10801), .Z(n1552) );
  NANDN U3106 ( .A(x[457]), .B(y[457]), .Z(n2894) );
  NANDN U3107 ( .A(n1552), .B(n2894), .Z(n1553) );
  NANDN U3108 ( .A(n10804), .B(n1553), .Z(n7209) );
  NANDN U3109 ( .A(y[454]), .B(x[454]), .Z(n1554) );
  NANDN U3110 ( .A(n1554), .B(x[455]), .Z(n1557) );
  XNOR U3111 ( .A(n1554), .B(x[455]), .Z(n1555) );
  NANDN U3112 ( .A(y[455]), .B(n1555), .Z(n1556) );
  AND U3113 ( .A(n1557), .B(n1556), .Z(n10796) );
  NANDN U3114 ( .A(x[455]), .B(y[455]), .Z(n1559) );
  NANDN U3115 ( .A(x[454]), .B(y[454]), .Z(n1558) );
  AND U3116 ( .A(n1559), .B(n1558), .Z(n1565) );
  NANDN U3117 ( .A(x[452]), .B(y[452]), .Z(n1560) );
  NANDN U3118 ( .A(y[453]), .B(n1560), .Z(n1563) );
  XNOR U3119 ( .A(n1560), .B(y[453]), .Z(n1561) );
  NAND U3120 ( .A(n1561), .B(x[453]), .Z(n1562) );
  NAND U3121 ( .A(n1563), .B(n1562), .Z(n1564) );
  NAND U3122 ( .A(n1565), .B(n1564), .Z(n10794) );
  NANDN U3123 ( .A(x[451]), .B(y[451]), .Z(n1567) );
  NANDN U3124 ( .A(x[450]), .B(y[450]), .Z(n1566) );
  AND U3125 ( .A(n1567), .B(n1566), .Z(n1573) );
  NANDN U3126 ( .A(x[448]), .B(y[448]), .Z(n1568) );
  NANDN U3127 ( .A(y[449]), .B(n1568), .Z(n1571) );
  XNOR U3128 ( .A(n1568), .B(y[449]), .Z(n1569) );
  NAND U3129 ( .A(n1569), .B(x[449]), .Z(n1570) );
  NAND U3130 ( .A(n1571), .B(n1570), .Z(n1572) );
  NAND U3131 ( .A(n1573), .B(n1572), .Z(n10790) );
  NANDN U3132 ( .A(y[449]), .B(x[449]), .Z(n1575) );
  NANDN U3133 ( .A(y[448]), .B(x[448]), .Z(n1574) );
  NAND U3134 ( .A(n1575), .B(n1574), .Z(n10788) );
  NANDN U3135 ( .A(y[446]), .B(x[446]), .Z(n10781) );
  ANDN U3136 ( .B(x[447]), .A(y[447]), .Z(n10785) );
  ANDN U3137 ( .B(n10781), .A(n10785), .Z(n1576) );
  NANDN U3138 ( .A(x[447]), .B(y[447]), .Z(n1580) );
  NANDN U3139 ( .A(n1576), .B(n1580), .Z(n1577) );
  NANDN U3140 ( .A(n10788), .B(n1577), .Z(n7202) );
  IV U3141 ( .A(y[446]), .Z(n1578) );
  OR U3142 ( .A(x[446]), .B(n1578), .Z(n1579) );
  NAND U3143 ( .A(n1580), .B(n1579), .Z(n10784) );
  NANDN U3144 ( .A(x[445]), .B(y[445]), .Z(n1582) );
  NANDN U3145 ( .A(x[444]), .B(y[444]), .Z(n1581) );
  AND U3146 ( .A(n1582), .B(n1581), .Z(n1588) );
  NANDN U3147 ( .A(x[442]), .B(y[442]), .Z(n1583) );
  NANDN U3148 ( .A(y[443]), .B(n1583), .Z(n1586) );
  XNOR U3149 ( .A(n1583), .B(y[443]), .Z(n1584) );
  NAND U3150 ( .A(n1584), .B(x[443]), .Z(n1585) );
  NAND U3151 ( .A(n1586), .B(n1585), .Z(n1587) );
  NAND U3152 ( .A(n1588), .B(n1587), .Z(n10778) );
  NANDN U3153 ( .A(x[438]), .B(y[438]), .Z(n1589) );
  ANDN U3154 ( .B(y[439]), .A(x[439]), .Z(n2871) );
  ANDN U3155 ( .B(n1589), .A(n2871), .Z(n10769) );
  ANDN U3156 ( .B(x[437]), .A(y[437]), .Z(n10768) );
  ANDN U3157 ( .B(y[437]), .A(x[437]), .Z(n2864) );
  ANDN U3158 ( .B(x[436]), .A(y[436]), .Z(n10760) );
  NANDN U3159 ( .A(n2864), .B(n10760), .Z(n1590) );
  NANDN U3160 ( .A(n10768), .B(n1590), .Z(n7192) );
  NANDN U3161 ( .A(x[434]), .B(y[434]), .Z(n1591) );
  NANDN U3162 ( .A(x[435]), .B(y[435]), .Z(n7189) );
  NAND U3163 ( .A(n1591), .B(n7189), .Z(n10758) );
  NANDN U3164 ( .A(x[433]), .B(y[433]), .Z(n10024) );
  NANDN U3165 ( .A(x[430]), .B(y[430]), .Z(n1593) );
  NANDN U3166 ( .A(x[431]), .B(y[431]), .Z(n1592) );
  AND U3167 ( .A(n1593), .B(n1592), .Z(n10754) );
  ANDN U3168 ( .B(x[431]), .A(y[431]), .Z(n10026) );
  OR U3169 ( .A(n10754), .B(n10026), .Z(n7178) );
  NANDN U3170 ( .A(x[428]), .B(y[428]), .Z(n1594) );
  NANDN U3171 ( .A(x[429]), .B(y[429]), .Z(n2850) );
  AND U3172 ( .A(n1594), .B(n2850), .Z(n10752) );
  NANDN U3173 ( .A(y[424]), .B(x[424]), .Z(n1596) );
  NANDN U3174 ( .A(y[423]), .B(x[423]), .Z(n1595) );
  NAND U3175 ( .A(n1596), .B(n1595), .Z(n10748) );
  NANDN U3176 ( .A(x[422]), .B(y[422]), .Z(n1598) );
  NANDN U3177 ( .A(x[423]), .B(y[423]), .Z(n1597) );
  AND U3178 ( .A(n1598), .B(n1597), .Z(n10747) );
  NANDN U3179 ( .A(y[422]), .B(x[422]), .Z(n1600) );
  NANDN U3180 ( .A(y[421]), .B(x[421]), .Z(n1599) );
  NAND U3181 ( .A(n1600), .B(n1599), .Z(n10746) );
  NANDN U3182 ( .A(y[420]), .B(x[420]), .Z(n1602) );
  NANDN U3183 ( .A(y[419]), .B(x[419]), .Z(n1601) );
  NAND U3184 ( .A(n1602), .B(n1601), .Z(n10744) );
  NANDN U3185 ( .A(y[417]), .B(x[417]), .Z(n6538) );
  NANDN U3186 ( .A(x[416]), .B(y[416]), .Z(n6536) );
  NANDN U3187 ( .A(x[412]), .B(y[412]), .Z(n1603) );
  ANDN U3188 ( .B(y[413]), .A(x[413]), .Z(n2820) );
  ANDN U3189 ( .B(n1603), .A(n2820), .Z(n10731) );
  NANDN U3190 ( .A(x[411]), .B(y[411]), .Z(n2814) );
  NANDN U3191 ( .A(y[410]), .B(x[410]), .Z(n10723) );
  ANDN U3192 ( .B(x[411]), .A(y[411]), .Z(n10727) );
  ANDN U3193 ( .B(n10723), .A(n10727), .Z(n1604) );
  ANDN U3194 ( .B(n2814), .A(n1604), .Z(n7148) );
  NANDN U3195 ( .A(x[409]), .B(y[409]), .Z(n1606) );
  NANDN U3196 ( .A(x[408]), .B(y[408]), .Z(n1605) );
  AND U3197 ( .A(n1606), .B(n1605), .Z(n1612) );
  NANDN U3198 ( .A(x[406]), .B(y[406]), .Z(n1607) );
  NANDN U3199 ( .A(y[407]), .B(n1607), .Z(n1610) );
  XNOR U3200 ( .A(n1607), .B(y[407]), .Z(n1608) );
  NAND U3201 ( .A(n1608), .B(x[407]), .Z(n1609) );
  NAND U3202 ( .A(n1610), .B(n1609), .Z(n1611) );
  NAND U3203 ( .A(n1612), .B(n1611), .Z(n10720) );
  NANDN U3204 ( .A(x[404]), .B(y[404]), .Z(n1613) );
  ANDN U3205 ( .B(y[405]), .A(x[405]), .Z(n2805) );
  ANDN U3206 ( .B(n1613), .A(n2805), .Z(n10716) );
  NANDN U3207 ( .A(x[399]), .B(y[399]), .Z(n6539) );
  NANDN U3208 ( .A(x[398]), .B(y[398]), .Z(n1614) );
  NAND U3209 ( .A(n6539), .B(n1614), .Z(n6548) );
  NANDN U3210 ( .A(y[396]), .B(x[396]), .Z(n1615) );
  NANDN U3211 ( .A(y[397]), .B(x[397]), .Z(n6545) );
  NAND U3212 ( .A(n1615), .B(n6545), .Z(n6550) );
  NANDN U3213 ( .A(x[396]), .B(y[396]), .Z(n6544) );
  NANDN U3214 ( .A(x[395]), .B(y[395]), .Z(n1617) );
  NANDN U3215 ( .A(x[394]), .B(y[394]), .Z(n1616) );
  NAND U3216 ( .A(n1617), .B(n1616), .Z(n10702) );
  ANDN U3217 ( .B(x[393]), .A(y[393]), .Z(n6554) );
  NANDN U3218 ( .A(y[390]), .B(x[390]), .Z(n1619) );
  NANDN U3219 ( .A(y[389]), .B(x[389]), .Z(n1618) );
  AND U3220 ( .A(n1619), .B(n1618), .Z(n1620) );
  NANDN U3221 ( .A(y[391]), .B(x[391]), .Z(n2776) );
  NAND U3222 ( .A(n1620), .B(n2776), .Z(n10692) );
  ANDN U3223 ( .B(y[389]), .A(x[389]), .Z(n2769) );
  ANDN U3224 ( .B(x[388]), .A(y[388]), .Z(n10688) );
  NANDN U3225 ( .A(n2769), .B(n10688), .Z(n1621) );
  NANDN U3226 ( .A(n10692), .B(n1621), .Z(n7130) );
  NANDN U3227 ( .A(y[382]), .B(x[382]), .Z(n1623) );
  NANDN U3228 ( .A(y[381]), .B(x[381]), .Z(n1622) );
  AND U3229 ( .A(n1623), .B(n1622), .Z(n1625) );
  NANDN U3230 ( .A(y[383]), .B(x[383]), .Z(n1624) );
  NAND U3231 ( .A(n1625), .B(n1624), .Z(n10676) );
  ANDN U3232 ( .B(y[381]), .A(x[381]), .Z(n2747) );
  ANDN U3233 ( .B(x[380]), .A(y[380]), .Z(n10030) );
  NANDN U3234 ( .A(n2747), .B(n10030), .Z(n1626) );
  NANDN U3235 ( .A(n10676), .B(n1626), .Z(n7122) );
  NANDN U3236 ( .A(x[379]), .B(y[379]), .Z(n1628) );
  NANDN U3237 ( .A(x[378]), .B(y[378]), .Z(n1627) );
  NAND U3238 ( .A(n1628), .B(n1627), .Z(n10670) );
  NANDN U3239 ( .A(x[376]), .B(y[376]), .Z(n1629) );
  ANDN U3240 ( .B(y[377]), .A(x[377]), .Z(n2742) );
  ANDN U3241 ( .B(n1629), .A(n2742), .Z(n10665) );
  NANDN U3242 ( .A(x[375]), .B(y[375]), .Z(n1631) );
  NANDN U3243 ( .A(x[374]), .B(y[374]), .Z(n1630) );
  NAND U3244 ( .A(n1631), .B(n1630), .Z(n10661) );
  ANDN U3245 ( .B(x[374]), .A(y[374]), .Z(n10660) );
  NANDN U3246 ( .A(y[372]), .B(x[372]), .Z(n1632) );
  ANDN U3247 ( .B(x[373]), .A(y[373]), .Z(n10659) );
  ANDN U3248 ( .B(n1632), .A(n10659), .Z(n1633) );
  NANDN U3249 ( .A(x[373]), .B(y[373]), .Z(n1635) );
  NANDN U3250 ( .A(n1633), .B(n1635), .Z(n1634) );
  NANDN U3251 ( .A(n10660), .B(n1634), .Z(n7112) );
  NANDN U3252 ( .A(x[370]), .B(y[370]), .Z(n1636) );
  ANDN U3253 ( .B(y[371]), .A(x[371]), .Z(n2732) );
  ANDN U3254 ( .B(n1636), .A(n2732), .Z(n10656) );
  NANDN U3255 ( .A(x[369]), .B(y[369]), .Z(n1638) );
  NANDN U3256 ( .A(x[368]), .B(y[368]), .Z(n1637) );
  NAND U3257 ( .A(n1638), .B(n1637), .Z(n10653) );
  ANDN U3258 ( .B(x[368]), .A(y[368]), .Z(n10652) );
  ANDN U3259 ( .B(y[367]), .A(x[367]), .Z(n1642) );
  ANDN U3260 ( .B(x[367]), .A(y[367]), .Z(n10033) );
  NANDN U3261 ( .A(y[366]), .B(x[366]), .Z(n1639) );
  NANDN U3262 ( .A(n10033), .B(n1639), .Z(n10650) );
  NANDN U3263 ( .A(n1642), .B(n10650), .Z(n1640) );
  NANDN U3264 ( .A(n10652), .B(n1640), .Z(n7104) );
  NANDN U3265 ( .A(x[366]), .B(y[366]), .Z(n1641) );
  NANDN U3266 ( .A(n1642), .B(n1641), .Z(n10032) );
  NANDN U3267 ( .A(y[359]), .B(x[359]), .Z(n2697) );
  NANDN U3268 ( .A(y[358]), .B(x[358]), .Z(n1643) );
  NAND U3269 ( .A(n2697), .B(n1643), .Z(n10644) );
  NANDN U3270 ( .A(x[349]), .B(y[349]), .Z(n1648) );
  XNOR U3271 ( .A(x[349]), .B(y[349]), .Z(n1645) );
  NANDN U3272 ( .A(y[348]), .B(x[348]), .Z(n1644) );
  NAND U3273 ( .A(n1645), .B(n1644), .Z(n1646) );
  AND U3274 ( .A(n1648), .B(n1646), .Z(n10628) );
  NANDN U3275 ( .A(x[348]), .B(y[348]), .Z(n1647) );
  AND U3276 ( .A(n1648), .B(n1647), .Z(n1654) );
  NANDN U3277 ( .A(x[346]), .B(y[346]), .Z(n1649) );
  NANDN U3278 ( .A(y[347]), .B(n1649), .Z(n1652) );
  XNOR U3279 ( .A(n1649), .B(y[347]), .Z(n1650) );
  NAND U3280 ( .A(n1650), .B(x[347]), .Z(n1651) );
  NAND U3281 ( .A(n1652), .B(n1651), .Z(n1653) );
  NAND U3282 ( .A(n1654), .B(n1653), .Z(n10626) );
  NANDN U3283 ( .A(y[346]), .B(x[346]), .Z(n1656) );
  NANDN U3284 ( .A(y[345]), .B(x[345]), .Z(n1655) );
  AND U3285 ( .A(n1656), .B(n1655), .Z(n1658) );
  NANDN U3286 ( .A(y[347]), .B(x[347]), .Z(n1657) );
  NAND U3287 ( .A(n1658), .B(n1657), .Z(n10624) );
  ANDN U3288 ( .B(y[345]), .A(x[345]), .Z(n2667) );
  ANDN U3289 ( .B(x[344]), .A(y[344]), .Z(n10617) );
  NANDN U3290 ( .A(n2667), .B(n10617), .Z(n1659) );
  NANDN U3291 ( .A(n10624), .B(n1659), .Z(n7085) );
  NANDN U3292 ( .A(x[342]), .B(y[342]), .Z(n1661) );
  NANDN U3293 ( .A(x[343]), .B(y[343]), .Z(n1660) );
  AND U3294 ( .A(n1661), .B(n1660), .Z(n10616) );
  NANDN U3295 ( .A(y[342]), .B(x[342]), .Z(n1663) );
  NANDN U3296 ( .A(y[341]), .B(x[341]), .Z(n1662) );
  NAND U3297 ( .A(n1663), .B(n1662), .Z(n10614) );
  ANDN U3298 ( .B(y[341]), .A(x[341]), .Z(n2661) );
  ANDN U3299 ( .B(x[340]), .A(y[340]), .Z(n10610) );
  NANDN U3300 ( .A(n2661), .B(n10610), .Z(n1664) );
  NANDN U3301 ( .A(n10614), .B(n1664), .Z(n7080) );
  NANDN U3302 ( .A(x[339]), .B(y[339]), .Z(n1666) );
  NANDN U3303 ( .A(x[338]), .B(y[338]), .Z(n1665) );
  NAND U3304 ( .A(n1666), .B(n1665), .Z(n10607) );
  NANDN U3305 ( .A(x[336]), .B(y[336]), .Z(n1667) );
  ANDN U3306 ( .B(y[337]), .A(x[337]), .Z(n2656) );
  ANDN U3307 ( .B(n1667), .A(n2656), .Z(n10605) );
  ANDN U3308 ( .B(x[335]), .A(y[335]), .Z(n10604) );
  ANDN U3309 ( .B(y[335]), .A(x[335]), .Z(n2649) );
  ANDN U3310 ( .B(x[334]), .A(y[334]), .Z(n10600) );
  NANDN U3311 ( .A(n2649), .B(n10600), .Z(n1668) );
  NANDN U3312 ( .A(n10604), .B(n1668), .Z(n7072) );
  NANDN U3313 ( .A(x[331]), .B(y[331]), .Z(n10035) );
  ANDN U3314 ( .B(x[330]), .A(y[330]), .Z(n10596) );
  ANDN U3315 ( .B(x[331]), .A(y[331]), .Z(n10597) );
  OR U3316 ( .A(n10596), .B(n10597), .Z(n7064) );
  NANDN U3317 ( .A(x[329]), .B(y[329]), .Z(n10594) );
  NANDN U3318 ( .A(y[327]), .B(x[327]), .Z(n2638) );
  NANDN U3319 ( .A(y[326]), .B(x[326]), .Z(n1669) );
  NAND U3320 ( .A(n2638), .B(n1669), .Z(n10587) );
  ANDN U3321 ( .B(y[325]), .A(x[325]), .Z(n2631) );
  ANDN U3322 ( .B(x[325]), .A(y[325]), .Z(n10584) );
  NANDN U3323 ( .A(y[324]), .B(x[324]), .Z(n1670) );
  NANDN U3324 ( .A(n10584), .B(n1670), .Z(n10036) );
  NANDN U3325 ( .A(n2631), .B(n10036), .Z(n1671) );
  NANDN U3326 ( .A(n10587), .B(n1671), .Z(n7057) );
  NANDN U3327 ( .A(x[322]), .B(y[322]), .Z(n1673) );
  NANDN U3328 ( .A(x[323]), .B(y[323]), .Z(n1672) );
  AND U3329 ( .A(n1673), .B(n1672), .Z(n10579) );
  NANDN U3330 ( .A(y[321]), .B(x[321]), .Z(n6558) );
  NANDN U3331 ( .A(y[320]), .B(x[320]), .Z(n1674) );
  NAND U3332 ( .A(n6558), .B(n1674), .Z(n10573) );
  ANDN U3333 ( .B(y[320]), .A(x[320]), .Z(n6557) );
  ANDN U3334 ( .B(n10571), .A(n6557), .Z(n2625) );
  NANDN U3335 ( .A(y[319]), .B(x[319]), .Z(n1676) );
  NANDN U3336 ( .A(y[318]), .B(x[318]), .Z(n1675) );
  AND U3337 ( .A(n1676), .B(n1675), .Z(n1682) );
  NANDN U3338 ( .A(y[316]), .B(x[316]), .Z(n1677) );
  NANDN U3339 ( .A(x[317]), .B(n1677), .Z(n1680) );
  XNOR U3340 ( .A(n1677), .B(x[317]), .Z(n1678) );
  NAND U3341 ( .A(n1678), .B(y[317]), .Z(n1679) );
  NAND U3342 ( .A(n1680), .B(n1679), .Z(n1681) );
  NAND U3343 ( .A(n1682), .B(n1681), .Z(n10570) );
  NANDN U3344 ( .A(y[310]), .B(x[310]), .Z(n1684) );
  NANDN U3345 ( .A(y[309]), .B(x[309]), .Z(n1683) );
  AND U3346 ( .A(n1684), .B(n1683), .Z(n1686) );
  NANDN U3347 ( .A(y[311]), .B(x[311]), .Z(n1685) );
  NAND U3348 ( .A(n1686), .B(n1685), .Z(n10561) );
  ANDN U3349 ( .B(y[309]), .A(x[309]), .Z(n2592) );
  ANDN U3350 ( .B(x[308]), .A(y[308]), .Z(n10558) );
  NANDN U3351 ( .A(n2592), .B(n10558), .Z(n1687) );
  NANDN U3352 ( .A(n10561), .B(n1687), .Z(n7044) );
  NANDN U3353 ( .A(x[304]), .B(y[304]), .Z(n1688) );
  ANDN U3354 ( .B(y[305]), .A(x[305]), .Z(n2585) );
  ANDN U3355 ( .B(n1688), .A(n2585), .Z(n10547) );
  NANDN U3356 ( .A(x[303]), .B(y[303]), .Z(n1690) );
  NANDN U3357 ( .A(x[302]), .B(y[302]), .Z(n1689) );
  NAND U3358 ( .A(n1690), .B(n1689), .Z(n10544) );
  NANDN U3359 ( .A(y[302]), .B(x[302]), .Z(n1692) );
  NANDN U3360 ( .A(y[301]), .B(x[301]), .Z(n1691) );
  NAND U3361 ( .A(n1692), .B(n1691), .Z(n10541) );
  ANDN U3362 ( .B(y[301]), .A(x[301]), .Z(n2578) );
  ANDN U3363 ( .B(x[300]), .A(y[300]), .Z(n10538) );
  NANDN U3364 ( .A(n2578), .B(n10538), .Z(n1693) );
  NANDN U3365 ( .A(n10541), .B(n1693), .Z(n7033) );
  NANDN U3366 ( .A(x[299]), .B(y[299]), .Z(n2575) );
  NANDN U3367 ( .A(x[297]), .B(y[297]), .Z(n1695) );
  NANDN U3368 ( .A(x[296]), .B(y[296]), .Z(n1694) );
  NAND U3369 ( .A(n1695), .B(n1694), .Z(n10528) );
  NANDN U3370 ( .A(y[296]), .B(x[296]), .Z(n1697) );
  NANDN U3371 ( .A(y[295]), .B(x[295]), .Z(n1696) );
  NAND U3372 ( .A(n1697), .B(n1696), .Z(n10526) );
  ANDN U3373 ( .B(y[295]), .A(x[295]), .Z(n2567) );
  ANDN U3374 ( .B(x[294]), .A(y[294]), .Z(n10519) );
  NANDN U3375 ( .A(n2567), .B(n10519), .Z(n1698) );
  NANDN U3376 ( .A(n10526), .B(n1698), .Z(n7025) );
  NANDN U3377 ( .A(x[291]), .B(y[291]), .Z(n1700) );
  NANDN U3378 ( .A(x[290]), .B(y[290]), .Z(n1699) );
  NAND U3379 ( .A(n1700), .B(n1699), .Z(n10514) );
  NANDN U3380 ( .A(x[289]), .B(y[289]), .Z(n1702) );
  NANDN U3381 ( .A(x[288]), .B(y[288]), .Z(n1701) );
  NAND U3382 ( .A(n1702), .B(n1701), .Z(n10510) );
  NANDN U3383 ( .A(x[286]), .B(y[286]), .Z(n1703) );
  ANDN U3384 ( .B(y[287]), .A(x[287]), .Z(n2552) );
  ANDN U3385 ( .B(n1703), .A(n2552), .Z(n10506) );
  NANDN U3386 ( .A(x[285]), .B(y[285]), .Z(n1705) );
  NANDN U3387 ( .A(x[284]), .B(y[284]), .Z(n1704) );
  NAND U3388 ( .A(n1705), .B(n1704), .Z(n10499) );
  NANDN U3389 ( .A(y[284]), .B(x[284]), .Z(n1707) );
  NANDN U3390 ( .A(y[283]), .B(x[283]), .Z(n1706) );
  NAND U3391 ( .A(n1707), .B(n1706), .Z(n10498) );
  ANDN U3392 ( .B(y[283]), .A(x[283]), .Z(n2543) );
  ANDN U3393 ( .B(x[282]), .A(y[282]), .Z(n10494) );
  NANDN U3394 ( .A(n2543), .B(n10494), .Z(n1708) );
  NANDN U3395 ( .A(n10498), .B(n1708), .Z(n7011) );
  NANDN U3396 ( .A(y[279]), .B(x[279]), .Z(n6999) );
  IV U3397 ( .A(x[280]), .Z(n7004) );
  OR U3398 ( .A(y[280]), .B(n7004), .Z(n1709) );
  NAND U3399 ( .A(n6999), .B(n1709), .Z(n10488) );
  NANDN U3400 ( .A(x[279]), .B(y[279]), .Z(n2538) );
  NANDN U3401 ( .A(x[276]), .B(y[276]), .Z(n6991) );
  NANDN U3402 ( .A(y[277]), .B(x[277]), .Z(n2533) );
  NANDN U3403 ( .A(n6991), .B(n2533), .Z(n1710) );
  NANDN U3404 ( .A(x[277]), .B(y[277]), .Z(n6995) );
  NAND U3405 ( .A(n1710), .B(n6995), .Z(n10482) );
  ANDN U3406 ( .B(n10485), .A(n10482), .Z(n2536) );
  NANDN U3407 ( .A(x[275]), .B(y[275]), .Z(n10474) );
  NANDN U3408 ( .A(y[271]), .B(x[271]), .Z(n2524) );
  NANDN U3409 ( .A(y[270]), .B(x[270]), .Z(n1711) );
  AND U3410 ( .A(n2524), .B(n1711), .Z(n1717) );
  NANDN U3411 ( .A(y[268]), .B(x[268]), .Z(n1712) );
  NANDN U3412 ( .A(x[269]), .B(n1712), .Z(n1715) );
  XNOR U3413 ( .A(n1712), .B(x[269]), .Z(n1713) );
  NAND U3414 ( .A(n1713), .B(y[269]), .Z(n1714) );
  NAND U3415 ( .A(n1715), .B(n1714), .Z(n1716) );
  NAND U3416 ( .A(n1717), .B(n1716), .Z(n10462) );
  NANDN U3417 ( .A(y[266]), .B(x[266]), .Z(n1719) );
  NANDN U3418 ( .A(y[265]), .B(x[265]), .Z(n1718) );
  AND U3419 ( .A(n1719), .B(n1718), .Z(n1721) );
  NANDN U3420 ( .A(y[267]), .B(x[267]), .Z(n1720) );
  NAND U3421 ( .A(n1721), .B(n1720), .Z(n10457) );
  ANDN U3422 ( .B(y[265]), .A(x[265]), .Z(n2515) );
  ANDN U3423 ( .B(x[264]), .A(y[264]), .Z(n10454) );
  NANDN U3424 ( .A(n2515), .B(n10454), .Z(n1722) );
  NANDN U3425 ( .A(n10457), .B(n1722), .Z(n6977) );
  NANDN U3426 ( .A(x[263]), .B(y[263]), .Z(n2512) );
  ANDN U3427 ( .B(x[261]), .A(y[261]), .Z(n10445) );
  ANDN U3428 ( .B(y[261]), .A(x[261]), .Z(n1725) );
  ANDN U3429 ( .B(x[260]), .A(y[260]), .Z(n10441) );
  NANDN U3430 ( .A(n1725), .B(n10441), .Z(n1723) );
  NANDN U3431 ( .A(n10445), .B(n1723), .Z(n6971) );
  NANDN U3432 ( .A(x[260]), .B(y[260]), .Z(n1724) );
  NANDN U3433 ( .A(n1725), .B(n1724), .Z(n10443) );
  NANDN U3434 ( .A(x[259]), .B(y[259]), .Z(n10438) );
  NANDN U3435 ( .A(n10443), .B(n10438), .Z(n6969) );
  ANDN U3436 ( .B(y[258]), .A(x[258]), .Z(n2507) );
  NANDN U3437 ( .A(x[257]), .B(y[257]), .Z(n1731) );
  ANDN U3438 ( .B(y[254]), .A(x[254]), .Z(n1726) );
  OR U3439 ( .A(n1726), .B(y[255]), .Z(n1729) );
  XOR U3440 ( .A(y[255]), .B(n1726), .Z(n1727) );
  NAND U3441 ( .A(n1727), .B(x[255]), .Z(n1728) );
  NAND U3442 ( .A(n1729), .B(n1728), .Z(n1730) );
  AND U3443 ( .A(n1731), .B(n1730), .Z(n1733) );
  NANDN U3444 ( .A(x[256]), .B(y[256]), .Z(n1732) );
  NAND U3445 ( .A(n1733), .B(n1732), .Z(n10434) );
  OR U3446 ( .A(n2507), .B(n10434), .Z(n6965) );
  NANDN U3447 ( .A(y[255]), .B(x[255]), .Z(n1735) );
  NANDN U3448 ( .A(y[254]), .B(x[254]), .Z(n1734) );
  AND U3449 ( .A(n1735), .B(n1734), .Z(n1741) );
  NANDN U3450 ( .A(y[252]), .B(x[252]), .Z(n1736) );
  NANDN U3451 ( .A(x[253]), .B(n1736), .Z(n1739) );
  XNOR U3452 ( .A(n1736), .B(x[253]), .Z(n1737) );
  NAND U3453 ( .A(n1737), .B(y[253]), .Z(n1738) );
  NAND U3454 ( .A(n1739), .B(n1738), .Z(n1740) );
  NAND U3455 ( .A(n1741), .B(n1740), .Z(n10432) );
  NANDN U3456 ( .A(y[251]), .B(x[251]), .Z(n1743) );
  NANDN U3457 ( .A(y[250]), .B(x[250]), .Z(n1742) );
  AND U3458 ( .A(n1743), .B(n1742), .Z(n1749) );
  NANDN U3459 ( .A(y[248]), .B(x[248]), .Z(n1744) );
  NANDN U3460 ( .A(x[249]), .B(n1744), .Z(n1747) );
  XNOR U3461 ( .A(n1744), .B(x[249]), .Z(n1745) );
  NAND U3462 ( .A(n1745), .B(y[249]), .Z(n1746) );
  NAND U3463 ( .A(n1747), .B(n1746), .Z(n1748) );
  NAND U3464 ( .A(n1749), .B(n1748), .Z(n10428) );
  NANDN U3465 ( .A(x[248]), .B(y[248]), .Z(n1751) );
  NANDN U3466 ( .A(x[247]), .B(y[247]), .Z(n1750) );
  AND U3467 ( .A(n1751), .B(n1750), .Z(n1753) );
  NANDN U3468 ( .A(x[249]), .B(y[249]), .Z(n1752) );
  NAND U3469 ( .A(n1753), .B(n1752), .Z(n6960) );
  NANDN U3470 ( .A(x[246]), .B(y[246]), .Z(n6954) );
  NANDN U3471 ( .A(y[247]), .B(x[247]), .Z(n1756) );
  NANDN U3472 ( .A(n6954), .B(n1756), .Z(n1754) );
  NANDN U3473 ( .A(n6960), .B(n1754), .Z(n10425) );
  NANDN U3474 ( .A(y[246]), .B(x[246]), .Z(n1755) );
  NAND U3475 ( .A(n1756), .B(n1755), .Z(n6958) );
  NANDN U3476 ( .A(y[245]), .B(x[245]), .Z(n1758) );
  NANDN U3477 ( .A(y[244]), .B(x[244]), .Z(n1757) );
  AND U3478 ( .A(n1758), .B(n1757), .Z(n6951) );
  NANDN U3479 ( .A(x[245]), .B(y[245]), .Z(n6955) );
  NANDN U3480 ( .A(n6951), .B(n6955), .Z(n1759) );
  NANDN U3481 ( .A(n6958), .B(n1759), .Z(n10423) );
  NANDN U3482 ( .A(x[244]), .B(y[244]), .Z(n1761) );
  NANDN U3483 ( .A(x[243]), .B(y[243]), .Z(n1760) );
  NAND U3484 ( .A(n1761), .B(n1760), .Z(n6950) );
  ANDN U3485 ( .B(n6955), .A(n6950), .Z(n1763) );
  NANDN U3486 ( .A(y[243]), .B(x[243]), .Z(n2481) );
  ANDN U3487 ( .B(y[242]), .A(x[242]), .Z(n6561) );
  NAND U3488 ( .A(n2481), .B(n6561), .Z(n1762) );
  NAND U3489 ( .A(n1763), .B(n1762), .Z(n10422) );
  NANDN U3490 ( .A(x[241]), .B(y[241]), .Z(n10417) );
  NANDN U3491 ( .A(x[240]), .B(y[240]), .Z(n1769) );
  ANDN U3492 ( .B(y[238]), .A(x[238]), .Z(n1764) );
  OR U3493 ( .A(n1764), .B(y[239]), .Z(n1767) );
  XOR U3494 ( .A(y[239]), .B(n1764), .Z(n1765) );
  NAND U3495 ( .A(n1765), .B(x[239]), .Z(n1766) );
  NAND U3496 ( .A(n1767), .B(n1766), .Z(n1768) );
  NAND U3497 ( .A(n1769), .B(n1768), .Z(n10414) );
  NANDN U3498 ( .A(x[236]), .B(y[236]), .Z(n1771) );
  NANDN U3499 ( .A(x[235]), .B(y[235]), .Z(n1770) );
  AND U3500 ( .A(n1771), .B(n1770), .Z(n1773) );
  NANDN U3501 ( .A(x[237]), .B(y[237]), .Z(n1772) );
  NAND U3502 ( .A(n1773), .B(n1772), .Z(n6942) );
  NANDN U3503 ( .A(x[234]), .B(y[234]), .Z(n6938) );
  NANDN U3504 ( .A(y[235]), .B(x[235]), .Z(n2472) );
  NANDN U3505 ( .A(n6938), .B(n2472), .Z(n1774) );
  NANDN U3506 ( .A(n6942), .B(n1774), .Z(n10410) );
  NANDN U3507 ( .A(y[233]), .B(x[233]), .Z(n2469) );
  NANDN U3508 ( .A(y[232]), .B(x[232]), .Z(n1775) );
  AND U3509 ( .A(n2469), .B(n1775), .Z(n1781) );
  NANDN U3510 ( .A(y[230]), .B(x[230]), .Z(n1776) );
  NANDN U3511 ( .A(x[231]), .B(n1776), .Z(n1779) );
  XNOR U3512 ( .A(n1776), .B(x[231]), .Z(n1777) );
  NAND U3513 ( .A(n1777), .B(y[231]), .Z(n1778) );
  NAND U3514 ( .A(n1779), .B(n1778), .Z(n1780) );
  NAND U3515 ( .A(n1781), .B(n1780), .Z(n10404) );
  NANDN U3516 ( .A(x[231]), .B(y[231]), .Z(n1783) );
  NANDN U3517 ( .A(x[230]), .B(y[230]), .Z(n1782) );
  AND U3518 ( .A(n1783), .B(n1782), .Z(n1789) );
  NANDN U3519 ( .A(x[228]), .B(y[228]), .Z(n1784) );
  NANDN U3520 ( .A(y[229]), .B(n1784), .Z(n1787) );
  XNOR U3521 ( .A(n1784), .B(y[229]), .Z(n1785) );
  NAND U3522 ( .A(n1785), .B(x[229]), .Z(n1786) );
  NAND U3523 ( .A(n1787), .B(n1786), .Z(n1788) );
  NAND U3524 ( .A(n1789), .B(n1788), .Z(n10402) );
  NANDN U3525 ( .A(x[227]), .B(y[227]), .Z(n1791) );
  NANDN U3526 ( .A(x[226]), .B(y[226]), .Z(n1790) );
  AND U3527 ( .A(n1791), .B(n1790), .Z(n1797) );
  NANDN U3528 ( .A(x[224]), .B(y[224]), .Z(n1792) );
  NANDN U3529 ( .A(y[225]), .B(n1792), .Z(n1795) );
  XNOR U3530 ( .A(n1792), .B(y[225]), .Z(n1793) );
  NAND U3531 ( .A(n1793), .B(x[225]), .Z(n1794) );
  NAND U3532 ( .A(n1795), .B(n1794), .Z(n1796) );
  NAND U3533 ( .A(n1797), .B(n1796), .Z(n10398) );
  NANDN U3534 ( .A(y[220]), .B(x[220]), .Z(n1799) );
  NANDN U3535 ( .A(y[219]), .B(x[219]), .Z(n1798) );
  AND U3536 ( .A(n1799), .B(n1798), .Z(n1801) );
  NANDN U3537 ( .A(y[221]), .B(x[221]), .Z(n1800) );
  NAND U3538 ( .A(n1801), .B(n1800), .Z(n10393) );
  NANDN U3539 ( .A(y[218]), .B(x[218]), .Z(n10040) );
  NANDN U3540 ( .A(x[219]), .B(y[219]), .Z(n1804) );
  NANDN U3541 ( .A(n10040), .B(n1804), .Z(n1802) );
  NANDN U3542 ( .A(n10393), .B(n1802), .Z(n6929) );
  NANDN U3543 ( .A(x[218]), .B(y[218]), .Z(n1803) );
  NAND U3544 ( .A(n1804), .B(n1803), .Z(n10392) );
  NANDN U3545 ( .A(y[216]), .B(x[216]), .Z(n1806) );
  NANDN U3546 ( .A(y[215]), .B(x[215]), .Z(n1805) );
  NAND U3547 ( .A(n1806), .B(n1805), .Z(n10390) );
  NANDN U3548 ( .A(y[214]), .B(x[214]), .Z(n1808) );
  NANDN U3549 ( .A(y[213]), .B(x[213]), .Z(n1807) );
  NAND U3550 ( .A(n1808), .B(n1807), .Z(n10388) );
  NANDN U3551 ( .A(x[211]), .B(y[211]), .Z(n2428) );
  NANDN U3552 ( .A(x[210]), .B(y[210]), .Z(n1809) );
  NAND U3553 ( .A(n2428), .B(n1809), .Z(n10385) );
  NANDN U3554 ( .A(x[209]), .B(y[209]), .Z(n6918) );
  NANDN U3555 ( .A(x[208]), .B(y[208]), .Z(n1810) );
  NAND U3556 ( .A(n6918), .B(n1810), .Z(n10384) );
  NANDN U3557 ( .A(y[207]), .B(x[207]), .Z(n6911) );
  NANDN U3558 ( .A(x[205]), .B(y[205]), .Z(n2415) );
  ANDN U3559 ( .B(x[203]), .A(y[203]), .Z(n10372) );
  ANDN U3560 ( .B(y[203]), .A(x[203]), .Z(n2410) );
  ANDN U3561 ( .B(x[202]), .A(y[202]), .Z(n10366) );
  NANDN U3562 ( .A(n2410), .B(n10366), .Z(n1811) );
  NANDN U3563 ( .A(n10372), .B(n1811), .Z(n6905) );
  ANDN U3564 ( .B(x[201]), .A(y[201]), .Z(n10369) );
  ANDN U3565 ( .B(y[201]), .A(x[201]), .Z(n2406) );
  ANDN U3566 ( .B(x[200]), .A(y[200]), .Z(n10360) );
  NANDN U3567 ( .A(n2406), .B(n10360), .Z(n1812) );
  NANDN U3568 ( .A(n10369), .B(n1812), .Z(n6901) );
  NANDN U3569 ( .A(y[199]), .B(x[199]), .Z(n10362) );
  NANDN U3570 ( .A(y[194]), .B(x[194]), .Z(n1814) );
  NANDN U3571 ( .A(y[193]), .B(x[193]), .Z(n1813) );
  AND U3572 ( .A(n1814), .B(n1813), .Z(n1816) );
  NANDN U3573 ( .A(y[195]), .B(x[195]), .Z(n1815) );
  NAND U3574 ( .A(n1816), .B(n1815), .Z(n10348) );
  ANDN U3575 ( .B(y[193]), .A(x[193]), .Z(n2388) );
  ANDN U3576 ( .B(x[192]), .A(y[192]), .Z(n10342) );
  NANDN U3577 ( .A(n2388), .B(n10342), .Z(n1817) );
  NANDN U3578 ( .A(n10348), .B(n1817), .Z(n6893) );
  NANDN U3579 ( .A(x[190]), .B(y[190]), .Z(n1819) );
  NANDN U3580 ( .A(x[191]), .B(y[191]), .Z(n1818) );
  AND U3581 ( .A(n1819), .B(n1818), .Z(n10340) );
  NANDN U3582 ( .A(y[190]), .B(x[190]), .Z(n1821) );
  NANDN U3583 ( .A(y[189]), .B(x[189]), .Z(n1820) );
  NAND U3584 ( .A(n1821), .B(n1820), .Z(n10339) );
  ANDN U3585 ( .B(y[189]), .A(x[189]), .Z(n2382) );
  ANDN U3586 ( .B(x[188]), .A(y[188]), .Z(n10335) );
  NANDN U3587 ( .A(n2382), .B(n10335), .Z(n1822) );
  NANDN U3588 ( .A(n10339), .B(n1822), .Z(n6887) );
  NANDN U3589 ( .A(x[187]), .B(y[187]), .Z(n1828) );
  XNOR U3590 ( .A(x[187]), .B(y[187]), .Z(n1824) );
  NANDN U3591 ( .A(y[186]), .B(x[186]), .Z(n1823) );
  NAND U3592 ( .A(n1824), .B(n1823), .Z(n1825) );
  AND U3593 ( .A(n1828), .B(n1825), .Z(n10332) );
  NANDN U3594 ( .A(x[186]), .B(y[186]), .Z(n1827) );
  NANDN U3595 ( .A(x[185]), .B(y[185]), .Z(n1826) );
  AND U3596 ( .A(n1827), .B(n1826), .Z(n1829) );
  NAND U3597 ( .A(n1829), .B(n1828), .Z(n10331) );
  NANDN U3598 ( .A(y[182]), .B(x[182]), .Z(n1831) );
  NANDN U3599 ( .A(y[181]), .B(x[181]), .Z(n1830) );
  AND U3600 ( .A(n1831), .B(n1830), .Z(n1833) );
  NANDN U3601 ( .A(y[183]), .B(x[183]), .Z(n1832) );
  NAND U3602 ( .A(n1833), .B(n1832), .Z(n10324) );
  ANDN U3603 ( .B(y[181]), .A(x[181]), .Z(n2366) );
  ANDN U3604 ( .B(x[180]), .A(y[180]), .Z(n10318) );
  NANDN U3605 ( .A(n2366), .B(n10318), .Z(n1834) );
  NANDN U3606 ( .A(n10324), .B(n1834), .Z(n6880) );
  NANDN U3607 ( .A(x[177]), .B(y[177]), .Z(n6875) );
  NANDN U3608 ( .A(x[176]), .B(y[176]), .Z(n1835) );
  NAND U3609 ( .A(n6875), .B(n1835), .Z(n10311) );
  NANDN U3610 ( .A(x[175]), .B(y[175]), .Z(n2350) );
  XNOR U3611 ( .A(x[175]), .B(y[175]), .Z(n1837) );
  NANDN U3612 ( .A(y[174]), .B(x[174]), .Z(n1836) );
  NAND U3613 ( .A(n1837), .B(n1836), .Z(n1838) );
  AND U3614 ( .A(n2350), .B(n1838), .Z(n6868) );
  NANDN U3615 ( .A(y[176]), .B(x[176]), .Z(n1839) );
  NANDN U3616 ( .A(n6868), .B(n1839), .Z(n10309) );
  NANDN U3617 ( .A(x[168]), .B(y[168]), .Z(n6859) );
  NANDN U3618 ( .A(y[169]), .B(x[169]), .Z(n1846) );
  NANDN U3619 ( .A(n6859), .B(n1846), .Z(n1844) );
  NANDN U3620 ( .A(x[170]), .B(y[170]), .Z(n1841) );
  NANDN U3621 ( .A(x[169]), .B(y[169]), .Z(n1840) );
  AND U3622 ( .A(n1841), .B(n1840), .Z(n1843) );
  NANDN U3623 ( .A(x[171]), .B(y[171]), .Z(n1842) );
  AND U3624 ( .A(n1843), .B(n1842), .Z(n6863) );
  NAND U3625 ( .A(n1844), .B(n6863), .Z(n10302) );
  NANDN U3626 ( .A(y[168]), .B(x[168]), .Z(n1845) );
  NAND U3627 ( .A(n1846), .B(n1845), .Z(n10300) );
  NANDN U3628 ( .A(y[167]), .B(x[167]), .Z(n1848) );
  NANDN U3629 ( .A(y[166]), .B(x[166]), .Z(n1847) );
  AND U3630 ( .A(n1848), .B(n1847), .Z(n1854) );
  NANDN U3631 ( .A(y[164]), .B(x[164]), .Z(n1849) );
  NANDN U3632 ( .A(x[165]), .B(n1849), .Z(n1852) );
  XNOR U3633 ( .A(n1849), .B(x[165]), .Z(n1850) );
  NAND U3634 ( .A(n1850), .B(y[165]), .Z(n1851) );
  NAND U3635 ( .A(n1852), .B(n1851), .Z(n1853) );
  NAND U3636 ( .A(n1854), .B(n1853), .Z(n10298) );
  NANDN U3637 ( .A(y[160]), .B(x[160]), .Z(n1856) );
  NANDN U3638 ( .A(y[159]), .B(x[159]), .Z(n1855) );
  AND U3639 ( .A(n1856), .B(n1855), .Z(n1858) );
  NANDN U3640 ( .A(y[161]), .B(x[161]), .Z(n1857) );
  NAND U3641 ( .A(n1858), .B(n1857), .Z(n10294) );
  ANDN U3642 ( .B(y[159]), .A(x[159]), .Z(n2317) );
  ANDN U3643 ( .B(x[158]), .A(y[158]), .Z(n10291) );
  NANDN U3644 ( .A(n2317), .B(n10291), .Z(n1859) );
  NANDN U3645 ( .A(n10294), .B(n1859), .Z(n6854) );
  NANDN U3646 ( .A(y[154]), .B(x[154]), .Z(n1861) );
  NANDN U3647 ( .A(y[153]), .B(x[153]), .Z(n1860) );
  NAND U3648 ( .A(n1861), .B(n1860), .Z(n10287) );
  NANDN U3649 ( .A(y[152]), .B(x[152]), .Z(n10044) );
  NANDN U3650 ( .A(x[153]), .B(y[153]), .Z(n1864) );
  NANDN U3651 ( .A(n10044), .B(n1864), .Z(n1862) );
  NANDN U3652 ( .A(n10287), .B(n1862), .Z(n6847) );
  NANDN U3653 ( .A(x[152]), .B(y[152]), .Z(n1863) );
  NAND U3654 ( .A(n1864), .B(n1863), .Z(n10286) );
  ANDN U3655 ( .B(x[147]), .A(y[147]), .Z(n10281) );
  ANDN U3656 ( .B(y[147]), .A(x[147]), .Z(n2290) );
  ANDN U3657 ( .B(x[146]), .A(y[146]), .Z(n10272) );
  NANDN U3658 ( .A(n2290), .B(n10272), .Z(n1865) );
  NANDN U3659 ( .A(n10281), .B(n1865), .Z(n6839) );
  NANDN U3660 ( .A(x[144]), .B(y[144]), .Z(n6831) );
  NANDN U3661 ( .A(x[145]), .B(y[145]), .Z(n6835) );
  NAND U3662 ( .A(n6831), .B(n6835), .Z(n10271) );
  NANDN U3663 ( .A(y[144]), .B(x[144]), .Z(n10268) );
  NANDN U3664 ( .A(y[143]), .B(x[143]), .Z(n1867) );
  NANDN U3665 ( .A(y[142]), .B(x[142]), .Z(n1866) );
  AND U3666 ( .A(n1867), .B(n1866), .Z(n1873) );
  NANDN U3667 ( .A(y[140]), .B(x[140]), .Z(n1868) );
  NANDN U3668 ( .A(x[141]), .B(n1868), .Z(n1871) );
  XNOR U3669 ( .A(n1868), .B(x[141]), .Z(n1869) );
  NAND U3670 ( .A(n1869), .B(y[141]), .Z(n1870) );
  NAND U3671 ( .A(n1871), .B(n1870), .Z(n1872) );
  NAND U3672 ( .A(n1873), .B(n1872), .Z(n10265) );
  NANDN U3673 ( .A(x[141]), .B(y[141]), .Z(n1875) );
  NANDN U3674 ( .A(x[140]), .B(y[140]), .Z(n1874) );
  AND U3675 ( .A(n1875), .B(n1874), .Z(n1881) );
  NANDN U3676 ( .A(x[138]), .B(y[138]), .Z(n1876) );
  NANDN U3677 ( .A(y[139]), .B(n1876), .Z(n1879) );
  XNOR U3678 ( .A(n1876), .B(y[139]), .Z(n1877) );
  NAND U3679 ( .A(n1877), .B(x[139]), .Z(n1878) );
  NAND U3680 ( .A(n1879), .B(n1878), .Z(n1880) );
  NAND U3681 ( .A(n1881), .B(n1880), .Z(n10263) );
  NANDN U3682 ( .A(y[138]), .B(x[138]), .Z(n1883) );
  NANDN U3683 ( .A(y[137]), .B(x[137]), .Z(n1882) );
  AND U3684 ( .A(n1883), .B(n1882), .Z(n1885) );
  NANDN U3685 ( .A(y[139]), .B(x[139]), .Z(n1884) );
  NAND U3686 ( .A(n1885), .B(n1884), .Z(n10260) );
  ANDN U3687 ( .B(y[137]), .A(x[137]), .Z(n2280) );
  ANDN U3688 ( .B(x[136]), .A(y[136]), .Z(n10257) );
  NANDN U3689 ( .A(n2280), .B(n10257), .Z(n1886) );
  NANDN U3690 ( .A(n10260), .B(n1886), .Z(n6827) );
  NANDN U3691 ( .A(x[133]), .B(y[133]), .Z(n1890) );
  XNOR U3692 ( .A(x[133]), .B(y[133]), .Z(n1888) );
  NANDN U3693 ( .A(y[132]), .B(x[132]), .Z(n1887) );
  NAND U3694 ( .A(n1888), .B(n1887), .Z(n1889) );
  AND U3695 ( .A(n1890), .B(n1889), .Z(n10248) );
  NANDN U3696 ( .A(y[131]), .B(x[131]), .Z(n2266) );
  NANDN U3697 ( .A(y[130]), .B(x[130]), .Z(n1891) );
  AND U3698 ( .A(n2266), .B(n1891), .Z(n1897) );
  ANDN U3699 ( .B(x[128]), .A(y[128]), .Z(n1892) );
  OR U3700 ( .A(n1892), .B(x[129]), .Z(n1895) );
  XOR U3701 ( .A(x[129]), .B(n1892), .Z(n1893) );
  NAND U3702 ( .A(n1893), .B(y[129]), .Z(n1894) );
  NAND U3703 ( .A(n1895), .B(n1894), .Z(n1896) );
  NAND U3704 ( .A(n1897), .B(n1896), .Z(n10244) );
  NANDN U3705 ( .A(x[123]), .B(y[123]), .Z(n6814) );
  IV U3706 ( .A(y[122]), .Z(n6567) );
  IV U3707 ( .A(x[122]), .Z(n6566) );
  NANDN U3708 ( .A(n6567), .B(n6566), .Z(n1898) );
  NAND U3709 ( .A(n6814), .B(n1898), .Z(n10232) );
  NANDN U3710 ( .A(x[119]), .B(y[119]), .Z(n1900) );
  NANDN U3711 ( .A(x[118]), .B(y[118]), .Z(n1899) );
  NAND U3712 ( .A(n1900), .B(n1899), .Z(n10225) );
  NANDN U3713 ( .A(y[118]), .B(x[118]), .Z(n1902) );
  NANDN U3714 ( .A(y[117]), .B(x[117]), .Z(n1901) );
  NAND U3715 ( .A(n1902), .B(n1901), .Z(n10223) );
  ANDN U3716 ( .B(y[117]), .A(x[117]), .Z(n2232) );
  ANDN U3717 ( .B(x[116]), .A(y[116]), .Z(n10216) );
  NANDN U3718 ( .A(n2232), .B(n10216), .Z(n1903) );
  NANDN U3719 ( .A(n10223), .B(n1903), .Z(n6802) );
  NANDN U3720 ( .A(x[115]), .B(y[115]), .Z(n1905) );
  NANDN U3721 ( .A(x[114]), .B(y[114]), .Z(n1904) );
  NAND U3722 ( .A(n1905), .B(n1904), .Z(n10214) );
  NANDN U3723 ( .A(y[113]), .B(x[113]), .Z(n1907) );
  ANDN U3724 ( .B(x[114]), .A(y[114]), .Z(n1906) );
  ANDN U3725 ( .B(n1907), .A(n1906), .Z(n1911) );
  XNOR U3726 ( .A(x[113]), .B(y[113]), .Z(n1909) );
  ANDN U3727 ( .B(x[112]), .A(y[112]), .Z(n1908) );
  NAND U3728 ( .A(n1909), .B(n1908), .Z(n1910) );
  AND U3729 ( .A(n1911), .B(n1910), .Z(n10212) );
  NANDN U3730 ( .A(x[113]), .B(y[113]), .Z(n1913) );
  NANDN U3731 ( .A(x[112]), .B(y[112]), .Z(n1912) );
  AND U3732 ( .A(n1913), .B(n1912), .Z(n1919) );
  NANDN U3733 ( .A(x[110]), .B(y[110]), .Z(n1914) );
  NANDN U3734 ( .A(y[111]), .B(n1914), .Z(n1917) );
  XNOR U3735 ( .A(n1914), .B(y[111]), .Z(n1915) );
  NAND U3736 ( .A(n1915), .B(x[111]), .Z(n1916) );
  NAND U3737 ( .A(n1917), .B(n1916), .Z(n1918) );
  NAND U3738 ( .A(n1919), .B(n1918), .Z(n10211) );
  NANDN U3739 ( .A(y[110]), .B(x[110]), .Z(n1921) );
  NANDN U3740 ( .A(y[109]), .B(x[109]), .Z(n1920) );
  AND U3741 ( .A(n1921), .B(n1920), .Z(n1923) );
  NANDN U3742 ( .A(y[111]), .B(x[111]), .Z(n1922) );
  NAND U3743 ( .A(n1923), .B(n1922), .Z(n10209) );
  ANDN U3744 ( .B(y[109]), .A(x[109]), .Z(n2224) );
  ANDN U3745 ( .B(x[108]), .A(y[108]), .Z(n10203) );
  NANDN U3746 ( .A(n2224), .B(n10203), .Z(n1924) );
  NANDN U3747 ( .A(n10209), .B(n1924), .Z(n6795) );
  NANDN U3748 ( .A(x[107]), .B(y[107]), .Z(n1926) );
  NANDN U3749 ( .A(x[106]), .B(y[106]), .Z(n1925) );
  NAND U3750 ( .A(n1926), .B(n1925), .Z(n10201) );
  NANDN U3751 ( .A(y[106]), .B(x[106]), .Z(n6569) );
  IV U3752 ( .A(x[104]), .Z(n1927) );
  XOR U3753 ( .A(y[104]), .B(n1927), .Z(n2215) );
  ANDN U3754 ( .B(x[103]), .A(y[103]), .Z(n6786) );
  NANDN U3755 ( .A(x[103]), .B(y[103]), .Z(n1929) );
  NANDN U3756 ( .A(x[102]), .B(y[102]), .Z(n1928) );
  NAND U3757 ( .A(n1929), .B(n1928), .Z(n10193) );
  NANDN U3758 ( .A(y[98]), .B(x[98]), .Z(n1931) );
  ANDN U3759 ( .B(x[100]), .A(y[100]), .Z(n2206) );
  NANDN U3760 ( .A(y[99]), .B(x[99]), .Z(n1930) );
  NANDN U3761 ( .A(n2206), .B(n1930), .Z(n10186) );
  ANDN U3762 ( .B(n1931), .A(n10186), .Z(n6780) );
  IV U3763 ( .A(y[97]), .Z(n10046) );
  OR U3764 ( .A(x[97]), .B(n10046), .Z(n1933) );
  IV U3765 ( .A(y[98]), .Z(n10180) );
  OR U3766 ( .A(x[98]), .B(n10180), .Z(n1932) );
  NAND U3767 ( .A(n1933), .B(n1932), .Z(n6779) );
  NANDN U3768 ( .A(x[96]), .B(y[96]), .Z(n1935) );
  NANDN U3769 ( .A(x[95]), .B(y[95]), .Z(n1934) );
  NAND U3770 ( .A(n1935), .B(n1934), .Z(n10172) );
  NANDN U3771 ( .A(x[94]), .B(y[94]), .Z(n1941) );
  ANDN U3772 ( .B(y[92]), .A(x[92]), .Z(n1936) );
  OR U3773 ( .A(n1936), .B(y[93]), .Z(n1939) );
  XOR U3774 ( .A(y[93]), .B(n1936), .Z(n1937) );
  NAND U3775 ( .A(n1937), .B(x[93]), .Z(n1938) );
  NAND U3776 ( .A(n1939), .B(n1938), .Z(n1940) );
  NAND U3777 ( .A(n1941), .B(n1940), .Z(n10168) );
  NANDN U3778 ( .A(y[92]), .B(x[92]), .Z(n1943) );
  NANDN U3779 ( .A(y[91]), .B(x[91]), .Z(n1942) );
  AND U3780 ( .A(n1943), .B(n1942), .Z(n1945) );
  NANDN U3781 ( .A(y[93]), .B(x[93]), .Z(n1944) );
  NAND U3782 ( .A(n1945), .B(n1944), .Z(n10165) );
  ANDN U3783 ( .B(y[91]), .A(x[91]), .Z(n2192) );
  ANDN U3784 ( .B(x[90]), .A(y[90]), .Z(n10160) );
  NANDN U3785 ( .A(n2192), .B(n10160), .Z(n1946) );
  NANDN U3786 ( .A(n10165), .B(n1946), .Z(n6772) );
  ANDN U3787 ( .B(x[88]), .A(y[88]), .Z(n10156) );
  NANDN U3788 ( .A(y[86]), .B(x[86]), .Z(n1947) );
  ANDN U3789 ( .B(x[87]), .A(y[87]), .Z(n10154) );
  ANDN U3790 ( .B(n1947), .A(n10154), .Z(n1948) );
  NANDN U3791 ( .A(x[87]), .B(y[87]), .Z(n1950) );
  NANDN U3792 ( .A(n1948), .B(n1950), .Z(n1949) );
  NANDN U3793 ( .A(n10156), .B(n1949), .Z(n6767) );
  NANDN U3794 ( .A(x[85]), .B(y[85]), .Z(n1952) );
  NANDN U3795 ( .A(x[84]), .B(y[84]), .Z(n1951) );
  NAND U3796 ( .A(n1952), .B(n1951), .Z(n10146) );
  NANDN U3797 ( .A(x[82]), .B(y[82]), .Z(n1953) );
  ANDN U3798 ( .B(y[83]), .A(x[83]), .Z(n2181) );
  ANDN U3799 ( .B(n1953), .A(n2181), .Z(n10141) );
  NANDN U3800 ( .A(x[81]), .B(y[81]), .Z(n1955) );
  NANDN U3801 ( .A(x[80]), .B(y[80]), .Z(n1954) );
  NAND U3802 ( .A(n1955), .B(n1954), .Z(n10138) );
  NANDN U3803 ( .A(x[79]), .B(y[79]), .Z(n1957) );
  NANDN U3804 ( .A(x[78]), .B(y[78]), .Z(n1956) );
  NAND U3805 ( .A(n1957), .B(n1956), .Z(n10134) );
  NANDN U3806 ( .A(x[75]), .B(y[75]), .Z(n1959) );
  NANDN U3807 ( .A(x[74]), .B(y[74]), .Z(n1958) );
  NAND U3808 ( .A(n1959), .B(n1958), .Z(n10122) );
  NANDN U3809 ( .A(x[73]), .B(y[73]), .Z(n1961) );
  NANDN U3810 ( .A(x[72]), .B(y[72]), .Z(n1960) );
  AND U3811 ( .A(n1961), .B(n1960), .Z(n1967) );
  NANDN U3812 ( .A(x[70]), .B(y[70]), .Z(n1962) );
  NANDN U3813 ( .A(y[71]), .B(n1962), .Z(n1965) );
  XNOR U3814 ( .A(n1962), .B(y[71]), .Z(n1963) );
  NAND U3815 ( .A(n1963), .B(x[71]), .Z(n1964) );
  NAND U3816 ( .A(n1965), .B(n1964), .Z(n1966) );
  NAND U3817 ( .A(n1967), .B(n1966), .Z(n10118) );
  ANDN U3818 ( .B(x[67]), .A(y[67]), .Z(n10112) );
  NANDN U3819 ( .A(y[66]), .B(x[66]), .Z(n1969) );
  NANDN U3820 ( .A(y[65]), .B(x[65]), .Z(n1968) );
  NAND U3821 ( .A(n1969), .B(n1968), .Z(n10106) );
  NOR U3822 ( .A(n10112), .B(n10106), .Z(n1971) );
  NANDN U3823 ( .A(y[64]), .B(x[64]), .Z(n10100) );
  NANDN U3824 ( .A(x[65]), .B(y[65]), .Z(n1973) );
  NANDN U3825 ( .A(n10100), .B(n1973), .Z(n1970) );
  NAND U3826 ( .A(n1971), .B(n1970), .Z(n6744) );
  NANDN U3827 ( .A(x[64]), .B(y[64]), .Z(n1972) );
  NAND U3828 ( .A(n1973), .B(n1972), .Z(n10104) );
  ANDN U3829 ( .B(x[63]), .A(y[63]), .Z(n10102) );
  ANDN U3830 ( .B(y[63]), .A(x[63]), .Z(n2139) );
  ANDN U3831 ( .B(x[62]), .A(y[62]), .Z(n10093) );
  NANDN U3832 ( .A(n2139), .B(n10093), .Z(n1974) );
  NANDN U3833 ( .A(n10102), .B(n1974), .Z(n6741) );
  NANDN U3834 ( .A(x[60]), .B(y[60]), .Z(n1976) );
  NANDN U3835 ( .A(x[61]), .B(y[61]), .Z(n1975) );
  AND U3836 ( .A(n1976), .B(n1975), .Z(n10091) );
  NANDN U3837 ( .A(y[60]), .B(x[60]), .Z(n1978) );
  NANDN U3838 ( .A(y[59]), .B(x[59]), .Z(n1977) );
  NAND U3839 ( .A(n1978), .B(n1977), .Z(n10090) );
  NANDN U3840 ( .A(y[58]), .B(x[58]), .Z(n1980) );
  NANDN U3841 ( .A(y[57]), .B(x[57]), .Z(n1979) );
  NAND U3842 ( .A(n1980), .B(n1979), .Z(n10085) );
  NANDN U3843 ( .A(x[54]), .B(y[54]), .Z(n1981) );
  ANDN U3844 ( .B(y[55]), .A(x[55]), .Z(n2126) );
  ANDN U3845 ( .B(n1981), .A(n2126), .Z(n10079) );
  ANDN U3846 ( .B(x[53]), .A(y[53]), .Z(n10078) );
  ANDN U3847 ( .B(y[53]), .A(x[53]), .Z(n2119) );
  ANDN U3848 ( .B(x[52]), .A(y[52]), .Z(n10069) );
  NANDN U3849 ( .A(n2119), .B(n10069), .Z(n1982) );
  NANDN U3850 ( .A(n10078), .B(n1982), .Z(n6728) );
  NANDN U3851 ( .A(x[48]), .B(y[48]), .Z(n1983) );
  ANDN U3852 ( .B(y[49]), .A(x[49]), .Z(n2112) );
  ANDN U3853 ( .B(n1983), .A(n2112), .Z(n10063) );
  ANDN U3854 ( .B(y[46]), .A(x[46]), .Z(n6716) );
  NANDN U3855 ( .A(x[47]), .B(y[47]), .Z(n6721) );
  NANDN U3856 ( .A(n6716), .B(n6721), .Z(n1984) );
  NANDN U3857 ( .A(y[47]), .B(x[47]), .Z(n2106) );
  AND U3858 ( .A(n1984), .B(n2106), .Z(n10060) );
  ANDN U3859 ( .B(n10063), .A(n10060), .Z(n2109) );
  NANDN U3860 ( .A(y[38]), .B(x[38]), .Z(n1986) );
  NANDN U3861 ( .A(y[37]), .B(x[37]), .Z(n1985) );
  AND U3862 ( .A(n1986), .B(n1985), .Z(n1987) );
  NANDN U3863 ( .A(y[39]), .B(x[39]), .Z(n2089) );
  NAND U3864 ( .A(n1987), .B(n2089), .Z(n6691) );
  NANDN U3865 ( .A(x[35]), .B(y[35]), .Z(n1989) );
  NANDN U3866 ( .A(x[34]), .B(y[34]), .Z(n1988) );
  NAND U3867 ( .A(n1989), .B(n1988), .Z(n6685) );
  ANDN U3868 ( .B(x[33]), .A(y[33]), .Z(n6683) );
  NANDN U3869 ( .A(y[31]), .B(x[31]), .Z(n1991) );
  ANDN U3870 ( .B(x[32]), .A(y[32]), .Z(n1990) );
  ANDN U3871 ( .B(n1991), .A(n1990), .Z(n1995) );
  XNOR U3872 ( .A(x[31]), .B(y[31]), .Z(n1993) );
  ANDN U3873 ( .B(x[30]), .A(y[30]), .Z(n1992) );
  NAND U3874 ( .A(n1993), .B(n1992), .Z(n1994) );
  NAND U3875 ( .A(n1995), .B(n1994), .Z(n6679) );
  NANDN U3876 ( .A(x[31]), .B(y[31]), .Z(n1997) );
  NANDN U3877 ( .A(x[30]), .B(y[30]), .Z(n1996) );
  NAND U3878 ( .A(n1997), .B(n1996), .Z(n6677) );
  ANDN U3879 ( .B(x[28]), .A(y[28]), .Z(n6671) );
  NANDN U3880 ( .A(y[27]), .B(x[27]), .Z(n1999) );
  NANDN U3881 ( .A(y[26]), .B(x[26]), .Z(n1998) );
  NAND U3882 ( .A(n1999), .B(n1998), .Z(n6667) );
  NANDN U3883 ( .A(y[24]), .B(x[24]), .Z(n2055) );
  NANDN U3884 ( .A(y[22]), .B(x[22]), .Z(n2001) );
  NANDN U3885 ( .A(y[23]), .B(x[23]), .Z(n2000) );
  NAND U3886 ( .A(n2001), .B(n2000), .Z(n6651) );
  NANDN U3887 ( .A(x[20]), .B(y[20]), .Z(n2047) );
  IV U3888 ( .A(y[20]), .Z(n6571) );
  IV U3889 ( .A(x[20]), .Z(n6570) );
  XNOR U3890 ( .A(n6571), .B(n6570), .Z(n2045) );
  NANDN U3891 ( .A(y[19]), .B(x[19]), .Z(n6637) );
  NANDN U3892 ( .A(x[18]), .B(y[18]), .Z(n6573) );
  ANDN U3893 ( .B(x[18]), .A(y[18]), .Z(n6636) );
  ANDN U3894 ( .B(x[17]), .A(y[17]), .Z(n6631) );
  NOR U3895 ( .A(n6636), .B(n6631), .Z(n2040) );
  ANDN U3896 ( .B(x[16]), .A(y[16]), .Z(n6633) );
  ANDN U3897 ( .B(x[15]), .A(y[15]), .Z(n6622) );
  NOR U3898 ( .A(n6633), .B(n6622), .Z(n2036) );
  NANDN U3899 ( .A(x[15]), .B(y[15]), .Z(n6628) );
  NANDN U3900 ( .A(x[12]), .B(y[12]), .Z(n6575) );
  ANDN U3901 ( .B(x[12]), .A(y[12]), .Z(n6614) );
  ANDN U3902 ( .B(x[11]), .A(y[11]), .Z(n6609) );
  NOR U3903 ( .A(n6614), .B(n6609), .Z(n2028) );
  ANDN U3904 ( .B(x[10]), .A(y[10]), .Z(n6611) );
  NANDN U3905 ( .A(x[7]), .B(y[7]), .Z(n6600) );
  ANDN U3906 ( .B(x[5]), .A(y[5]), .Z(n6593) );
  ANDN U3907 ( .B(x[6]), .A(y[6]), .Z(n6599) );
  NOR U3908 ( .A(n6593), .B(n6599), .Z(n2012) );
  ANDN U3909 ( .B(x[4]), .A(y[4]), .Z(n6595) );
  ANDN U3910 ( .B(x[3]), .A(y[3]), .Z(n6584) );
  NOR U3911 ( .A(n6595), .B(n6584), .Z(n2008) );
  NANDN U3912 ( .A(x[3]), .B(y[3]), .Z(n6590) );
  ANDN U3913 ( .B(x[1]), .A(y[1]), .Z(n6579) );
  NANDN U3914 ( .A(x[0]), .B(y[0]), .Z(n2002) );
  NANDN U3915 ( .A(x[1]), .B(y[1]), .Z(n6582) );
  NAND U3916 ( .A(n2002), .B(n6582), .Z(n2003) );
  ANDN U3917 ( .B(x[2]), .A(y[2]), .Z(n6587) );
  ANDN U3918 ( .B(n2003), .A(n6587), .Z(n2004) );
  NANDN U3919 ( .A(n6579), .B(n2004), .Z(n2005) );
  AND U3920 ( .A(n6590), .B(n2005), .Z(n2006) );
  NANDN U3921 ( .A(x[2]), .B(y[2]), .Z(n6581) );
  NAND U3922 ( .A(n2006), .B(n6581), .Z(n2007) );
  NAND U3923 ( .A(n2008), .B(n2007), .Z(n2009) );
  NANDN U3924 ( .A(x[5]), .B(y[5]), .Z(n6576) );
  NAND U3925 ( .A(n2009), .B(n6576), .Z(n2010) );
  NANDN U3926 ( .A(x[4]), .B(y[4]), .Z(n6588) );
  NANDN U3927 ( .A(n2010), .B(n6588), .Z(n2011) );
  AND U3928 ( .A(n2012), .B(n2011), .Z(n2013) );
  ANDN U3929 ( .B(n6600), .A(n2013), .Z(n2014) );
  NANDN U3930 ( .A(x[6]), .B(y[6]), .Z(n6577) );
  NAND U3931 ( .A(n2014), .B(n6577), .Z(n2018) );
  NANDN U3932 ( .A(y[8]), .B(x[8]), .Z(n2016) );
  NANDN U3933 ( .A(y[7]), .B(x[7]), .Z(n2015) );
  AND U3934 ( .A(n2016), .B(n2015), .Z(n2017) );
  NANDN U3935 ( .A(y[9]), .B(x[9]), .Z(n2022) );
  NAND U3936 ( .A(n2017), .B(n2022), .Z(n6603) );
  ANDN U3937 ( .B(n2018), .A(n6603), .Z(n2023) );
  XNOR U3938 ( .A(y[9]), .B(x[9]), .Z(n2020) );
  NANDN U3939 ( .A(x[8]), .B(y[8]), .Z(n2019) );
  NAND U3940 ( .A(n2020), .B(n2019), .Z(n2021) );
  NAND U3941 ( .A(n2022), .B(n2021), .Z(n6605) );
  NANDN U3942 ( .A(n2023), .B(n6605), .Z(n2024) );
  NANDN U3943 ( .A(n6611), .B(n2024), .Z(n2025) );
  NANDN U3944 ( .A(x[11]), .B(y[11]), .Z(n6574) );
  NAND U3945 ( .A(n2025), .B(n6574), .Z(n2026) );
  NANDN U3946 ( .A(x[10]), .B(y[10]), .Z(n6606) );
  NANDN U3947 ( .A(n2026), .B(n6606), .Z(n2027) );
  AND U3948 ( .A(n2028), .B(n2027), .Z(n2029) );
  ANDN U3949 ( .B(n6575), .A(n2029), .Z(n2030) );
  NANDN U3950 ( .A(x[13]), .B(y[13]), .Z(n6620) );
  NAND U3951 ( .A(n2030), .B(n6620), .Z(n2031) );
  ANDN U3952 ( .B(x[14]), .A(y[14]), .Z(n6625) );
  ANDN U3953 ( .B(n2031), .A(n6625), .Z(n2032) );
  NANDN U3954 ( .A(y[13]), .B(x[13]), .Z(n6615) );
  NAND U3955 ( .A(n2032), .B(n6615), .Z(n2033) );
  AND U3956 ( .A(n6628), .B(n2033), .Z(n2034) );
  NANDN U3957 ( .A(x[14]), .B(y[14]), .Z(n6619) );
  NAND U3958 ( .A(n2034), .B(n6619), .Z(n2035) );
  NAND U3959 ( .A(n2036), .B(n2035), .Z(n2037) );
  NANDN U3960 ( .A(x[17]), .B(y[17]), .Z(n6572) );
  NAND U3961 ( .A(n2037), .B(n6572), .Z(n2038) );
  NANDN U3962 ( .A(x[16]), .B(y[16]), .Z(n6626) );
  NANDN U3963 ( .A(n2038), .B(n6626), .Z(n2039) );
  AND U3964 ( .A(n2040), .B(n2039), .Z(n2041) );
  ANDN U3965 ( .B(n6573), .A(n2041), .Z(n2042) );
  NANDN U3966 ( .A(x[19]), .B(y[19]), .Z(n6642) );
  NAND U3967 ( .A(n2042), .B(n6642), .Z(n2043) );
  AND U3968 ( .A(n6637), .B(n2043), .Z(n2044) );
  NAND U3969 ( .A(n2045), .B(n2044), .Z(n2046) );
  NAND U3970 ( .A(n2047), .B(n2046), .Z(n2048) );
  ANDN U3971 ( .B(x[21]), .A(y[21]), .Z(n6644) );
  ANDN U3972 ( .B(n2048), .A(n6644), .Z(n2051) );
  NANDN U3973 ( .A(x[22]), .B(y[22]), .Z(n2050) );
  NANDN U3974 ( .A(x[21]), .B(y[21]), .Z(n2049) );
  AND U3975 ( .A(n2050), .B(n2049), .Z(n6649) );
  NANDN U3976 ( .A(n2051), .B(n6649), .Z(n2052) );
  NANDN U3977 ( .A(n6651), .B(n2052), .Z(n2053) );
  NANDN U3978 ( .A(x[23]), .B(y[23]), .Z(n6653) );
  NAND U3979 ( .A(n2053), .B(n6653), .Z(n2054) );
  NAND U3980 ( .A(n2055), .B(n2054), .Z(n2058) );
  IV U3981 ( .A(y[24]), .Z(n6656) );
  IV U3982 ( .A(x[24]), .Z(n6657) );
  NANDN U3983 ( .A(n6656), .B(n6657), .Z(n2056) );
  ANDN U3984 ( .B(y[25]), .A(x[25]), .Z(n6662) );
  ANDN U3985 ( .B(n2056), .A(n6662), .Z(n2057) );
  NAND U3986 ( .A(n2058), .B(n2057), .Z(n2059) );
  ANDN U3987 ( .B(x[25]), .A(y[25]), .Z(n6658) );
  ANDN U3988 ( .B(n2059), .A(n6658), .Z(n2060) );
  NANDN U3989 ( .A(x[26]), .B(y[26]), .Z(n6664) );
  NANDN U3990 ( .A(n2060), .B(n6664), .Z(n2061) );
  NANDN U3991 ( .A(n6667), .B(n2061), .Z(n2062) );
  NANDN U3992 ( .A(x[27]), .B(y[27]), .Z(n6669) );
  NAND U3993 ( .A(n2062), .B(n6669), .Z(n2063) );
  NANDN U3994 ( .A(n6671), .B(n2063), .Z(n2066) );
  NANDN U3995 ( .A(x[28]), .B(y[28]), .Z(n2065) );
  NANDN U3996 ( .A(x[29]), .B(y[29]), .Z(n2064) );
  AND U3997 ( .A(n2065), .B(n2064), .Z(n6672) );
  NAND U3998 ( .A(n2066), .B(n6672), .Z(n2067) );
  ANDN U3999 ( .B(x[29]), .A(y[29]), .Z(n6675) );
  ANDN U4000 ( .B(n2067), .A(n6675), .Z(n2068) );
  OR U4001 ( .A(n6677), .B(n2068), .Z(n2069) );
  NANDN U4002 ( .A(n6679), .B(n2069), .Z(n2072) );
  NANDN U4003 ( .A(x[32]), .B(y[32]), .Z(n2071) );
  NANDN U4004 ( .A(x[33]), .B(y[33]), .Z(n2070) );
  AND U4005 ( .A(n2071), .B(n2070), .Z(n6681) );
  NAND U4006 ( .A(n2072), .B(n6681), .Z(n2073) );
  NANDN U4007 ( .A(n6683), .B(n2073), .Z(n2074) );
  NANDN U4008 ( .A(n6685), .B(n2074), .Z(n2081) );
  NANDN U4009 ( .A(y[35]), .B(x[35]), .Z(n2076) );
  ANDN U4010 ( .B(x[36]), .A(y[36]), .Z(n2075) );
  ANDN U4011 ( .B(n2076), .A(n2075), .Z(n2080) );
  XNOR U4012 ( .A(x[35]), .B(y[35]), .Z(n2078) );
  ANDN U4013 ( .B(x[34]), .A(y[34]), .Z(n2077) );
  NAND U4014 ( .A(n2078), .B(n2077), .Z(n2079) );
  NAND U4015 ( .A(n2080), .B(n2079), .Z(n6687) );
  ANDN U4016 ( .B(n2081), .A(n6687), .Z(n2084) );
  NANDN U4017 ( .A(x[37]), .B(y[37]), .Z(n2083) );
  NANDN U4018 ( .A(x[36]), .B(y[36]), .Z(n2082) );
  AND U4019 ( .A(n2083), .B(n2082), .Z(n6688) );
  NANDN U4020 ( .A(n2084), .B(n6688), .Z(n2085) );
  NANDN U4021 ( .A(n6691), .B(n2085), .Z(n2090) );
  XNOR U4022 ( .A(y[39]), .B(x[39]), .Z(n2087) );
  NANDN U4023 ( .A(x[38]), .B(y[38]), .Z(n2086) );
  NAND U4024 ( .A(n2087), .B(n2086), .Z(n2088) );
  NAND U4025 ( .A(n2089), .B(n2088), .Z(n6693) );
  NAND U4026 ( .A(n2090), .B(n6693), .Z(n2092) );
  ANDN U4027 ( .B(y[40]), .A(x[40]), .Z(n2091) );
  OR U4028 ( .A(n2092), .B(n2091), .Z(n2095) );
  IV U4029 ( .A(x[40]), .Z(n6696) );
  IV U4030 ( .A(y[40]), .Z(n6697) );
  NANDN U4031 ( .A(n6696), .B(n6697), .Z(n2093) );
  ANDN U4032 ( .B(x[41]), .A(y[41]), .Z(n6703) );
  ANDN U4033 ( .B(n2093), .A(n6703), .Z(n2094) );
  NAND U4034 ( .A(n2095), .B(n2094), .Z(n2096) );
  NANDN U4035 ( .A(x[41]), .B(y[41]), .Z(n6699) );
  NAND U4036 ( .A(n2096), .B(n6699), .Z(n2098) );
  NANDN U4037 ( .A(y[42]), .B(x[42]), .Z(n2097) );
  NAND U4038 ( .A(n2098), .B(n2097), .Z(n2101) );
  IV U4039 ( .A(y[42]), .Z(n6706) );
  IV U4040 ( .A(x[42]), .Z(n6707) );
  NANDN U4041 ( .A(n6706), .B(n6707), .Z(n2099) );
  ANDN U4042 ( .B(y[43]), .A(x[43]), .Z(n6713) );
  ANDN U4043 ( .B(n2099), .A(n6713), .Z(n2100) );
  NAND U4044 ( .A(n2101), .B(n2100), .Z(n2102) );
  ANDN U4045 ( .B(x[43]), .A(y[43]), .Z(n6708) );
  ANDN U4046 ( .B(n2102), .A(n6708), .Z(n2103) );
  NANDN U4047 ( .A(x[44]), .B(y[44]), .Z(n10050) );
  NANDN U4048 ( .A(n2103), .B(n10050), .Z(n2104) );
  NANDN U4049 ( .A(y[44]), .B(x[44]), .Z(n10052) );
  ANDN U4050 ( .B(x[45]), .A(y[45]), .Z(n10055) );
  ANDN U4051 ( .B(n10052), .A(n10055), .Z(n6714) );
  NAND U4052 ( .A(n2104), .B(n6714), .Z(n2105) );
  NANDN U4053 ( .A(x[45]), .B(y[45]), .Z(n10049) );
  NAND U4054 ( .A(n2105), .B(n10049), .Z(n2107) );
  NAND U4055 ( .A(n2107), .B(n10057), .Z(n2108) );
  AND U4056 ( .A(n2109), .B(n2108), .Z(n2114) );
  NANDN U4057 ( .A(y[50]), .B(x[50]), .Z(n2111) );
  NANDN U4058 ( .A(y[49]), .B(x[49]), .Z(n2110) );
  NAND U4059 ( .A(n2111), .B(n2110), .Z(n10066) );
  ANDN U4060 ( .B(x[48]), .A(y[48]), .Z(n10061) );
  NANDN U4061 ( .A(n2112), .B(n10061), .Z(n2113) );
  NANDN U4062 ( .A(n10066), .B(n2113), .Z(n6724) );
  OR U4063 ( .A(n2114), .B(n6724), .Z(n2117) );
  NANDN U4064 ( .A(x[50]), .B(y[50]), .Z(n2116) );
  NANDN U4065 ( .A(x[51]), .B(y[51]), .Z(n2115) );
  AND U4066 ( .A(n2116), .B(n2115), .Z(n10067) );
  NAND U4067 ( .A(n2117), .B(n10067), .Z(n2118) );
  NANDN U4068 ( .A(y[51]), .B(x[51]), .Z(n10071) );
  NAND U4069 ( .A(n2118), .B(n10071), .Z(n2121) );
  NANDN U4070 ( .A(x[52]), .B(y[52]), .Z(n2120) );
  ANDN U4071 ( .B(n2120), .A(n2119), .Z(n10073) );
  NAND U4072 ( .A(n2121), .B(n10073), .Z(n2122) );
  NANDN U4073 ( .A(n6728), .B(n2122), .Z(n2123) );
  AND U4074 ( .A(n10079), .B(n2123), .Z(n2128) );
  NANDN U4075 ( .A(y[56]), .B(x[56]), .Z(n2125) );
  NANDN U4076 ( .A(y[55]), .B(x[55]), .Z(n2124) );
  NAND U4077 ( .A(n2125), .B(n2124), .Z(n10082) );
  ANDN U4078 ( .B(x[54]), .A(y[54]), .Z(n10075) );
  NANDN U4079 ( .A(n2126), .B(n10075), .Z(n2127) );
  NANDN U4080 ( .A(n10082), .B(n2127), .Z(n6732) );
  OR U4081 ( .A(n2128), .B(n6732), .Z(n2131) );
  NANDN U4082 ( .A(x[56]), .B(y[56]), .Z(n2130) );
  NANDN U4083 ( .A(x[57]), .B(y[57]), .Z(n2129) );
  AND U4084 ( .A(n2130), .B(n2129), .Z(n10083) );
  NAND U4085 ( .A(n2131), .B(n10083), .Z(n2132) );
  NANDN U4086 ( .A(n10085), .B(n2132), .Z(n2135) );
  NANDN U4087 ( .A(x[58]), .B(y[58]), .Z(n2134) );
  NANDN U4088 ( .A(x[59]), .B(y[59]), .Z(n2133) );
  AND U4089 ( .A(n2134), .B(n2133), .Z(n10087) );
  NAND U4090 ( .A(n2135), .B(n10087), .Z(n2136) );
  NANDN U4091 ( .A(n10090), .B(n2136), .Z(n2137) );
  AND U4092 ( .A(n10091), .B(n2137), .Z(n2138) );
  NANDN U4093 ( .A(y[61]), .B(x[61]), .Z(n10095) );
  NANDN U4094 ( .A(n2138), .B(n10095), .Z(n2141) );
  NANDN U4095 ( .A(x[62]), .B(y[62]), .Z(n2140) );
  ANDN U4096 ( .B(n2140), .A(n2139), .Z(n10097) );
  NAND U4097 ( .A(n2141), .B(n10097), .Z(n2142) );
  NANDN U4098 ( .A(n6741), .B(n2142), .Z(n2143) );
  NANDN U4099 ( .A(n10104), .B(n2143), .Z(n2144) );
  NANDN U4100 ( .A(n6744), .B(n2144), .Z(n2149) );
  ANDN U4101 ( .B(y[69]), .A(x[69]), .Z(n2154) );
  NANDN U4102 ( .A(x[68]), .B(y[68]), .Z(n2145) );
  NANDN U4103 ( .A(n2154), .B(n2145), .Z(n10114) );
  NANDN U4104 ( .A(x[67]), .B(y[67]), .Z(n2147) );
  NANDN U4105 ( .A(x[66]), .B(y[66]), .Z(n2146) );
  NAND U4106 ( .A(n2147), .B(n2146), .Z(n10108) );
  NANDN U4107 ( .A(n10112), .B(n10108), .Z(n2148) );
  NANDN U4108 ( .A(n10114), .B(n2148), .Z(n6746) );
  ANDN U4109 ( .B(n2149), .A(n6746), .Z(n2156) );
  NANDN U4110 ( .A(y[70]), .B(x[70]), .Z(n2151) );
  NANDN U4111 ( .A(y[69]), .B(x[69]), .Z(n2150) );
  AND U4112 ( .A(n2151), .B(n2150), .Z(n2153) );
  NANDN U4113 ( .A(y[71]), .B(x[71]), .Z(n2152) );
  NAND U4114 ( .A(n2153), .B(n2152), .Z(n10115) );
  ANDN U4115 ( .B(x[68]), .A(y[68]), .Z(n10109) );
  NANDN U4116 ( .A(n2154), .B(n10109), .Z(n2155) );
  NANDN U4117 ( .A(n10115), .B(n2155), .Z(n6748) );
  OR U4118 ( .A(n2156), .B(n6748), .Z(n2157) );
  NANDN U4119 ( .A(n10118), .B(n2157), .Z(n2164) );
  NANDN U4120 ( .A(y[73]), .B(x[73]), .Z(n2159) );
  ANDN U4121 ( .B(x[74]), .A(y[74]), .Z(n2158) );
  ANDN U4122 ( .B(n2159), .A(n2158), .Z(n2163) );
  XNOR U4123 ( .A(x[73]), .B(y[73]), .Z(n2161) );
  ANDN U4124 ( .B(x[72]), .A(y[72]), .Z(n2160) );
  NAND U4125 ( .A(n2161), .B(n2160), .Z(n2162) );
  AND U4126 ( .A(n2163), .B(n2162), .Z(n10120) );
  NAND U4127 ( .A(n2164), .B(n10120), .Z(n2165) );
  NANDN U4128 ( .A(n10122), .B(n2165), .Z(n2166) );
  NANDN U4129 ( .A(y[75]), .B(x[75]), .Z(n10124) );
  NAND U4130 ( .A(n2166), .B(n10124), .Z(n2167) );
  NANDN U4131 ( .A(x[77]), .B(y[77]), .Z(n2168) );
  ANDN U4132 ( .B(n2167), .A(n10128), .Z(n2171) );
  ANDN U4133 ( .B(x[78]), .A(y[78]), .Z(n10132) );
  NANDN U4134 ( .A(y[76]), .B(x[76]), .Z(n10125) );
  ANDN U4135 ( .B(x[77]), .A(y[77]), .Z(n10129) );
  ANDN U4136 ( .B(n10125), .A(n10129), .Z(n2169) );
  NANDN U4137 ( .A(n2169), .B(n2168), .Z(n2170) );
  NANDN U4138 ( .A(n10132), .B(n2170), .Z(n6755) );
  OR U4139 ( .A(n2171), .B(n6755), .Z(n2172) );
  NANDN U4140 ( .A(n10134), .B(n2172), .Z(n2175) );
  NANDN U4141 ( .A(y[79]), .B(x[79]), .Z(n2174) );
  NANDN U4142 ( .A(y[80]), .B(x[80]), .Z(n2173) );
  AND U4143 ( .A(n2174), .B(n2173), .Z(n10136) );
  NAND U4144 ( .A(n2175), .B(n10136), .Z(n2176) );
  NANDN U4145 ( .A(n10138), .B(n2176), .Z(n2177) );
  NANDN U4146 ( .A(y[81]), .B(x[81]), .Z(n10048) );
  NAND U4147 ( .A(n2177), .B(n10048), .Z(n2178) );
  AND U4148 ( .A(n10141), .B(n2178), .Z(n2183) );
  NANDN U4149 ( .A(y[84]), .B(x[84]), .Z(n2180) );
  NANDN U4150 ( .A(y[83]), .B(x[83]), .Z(n2179) );
  NAND U4151 ( .A(n2180), .B(n2179), .Z(n10144) );
  ANDN U4152 ( .B(x[82]), .A(y[82]), .Z(n10047) );
  NANDN U4153 ( .A(n2181), .B(n10047), .Z(n2182) );
  NANDN U4154 ( .A(n10144), .B(n2182), .Z(n6762) );
  OR U4155 ( .A(n2183), .B(n6762), .Z(n2184) );
  NANDN U4156 ( .A(n10146), .B(n2184), .Z(n2185) );
  NANDN U4157 ( .A(y[85]), .B(x[85]), .Z(n10148) );
  NAND U4158 ( .A(n2185), .B(n10148), .Z(n2186) );
  NANDN U4159 ( .A(n10152), .B(n2186), .Z(n2187) );
  NANDN U4160 ( .A(n6767), .B(n2187), .Z(n2190) );
  NANDN U4161 ( .A(x[89]), .B(y[89]), .Z(n2189) );
  NANDN U4162 ( .A(x[88]), .B(y[88]), .Z(n2188) );
  NAND U4163 ( .A(n2189), .B(n2188), .Z(n10158) );
  ANDN U4164 ( .B(n2190), .A(n10158), .Z(n2191) );
  NANDN U4165 ( .A(y[89]), .B(x[89]), .Z(n10161) );
  NANDN U4166 ( .A(n2191), .B(n10161), .Z(n2194) );
  NANDN U4167 ( .A(x[90]), .B(y[90]), .Z(n2193) );
  ANDN U4168 ( .B(n2193), .A(n2192), .Z(n10163) );
  NAND U4169 ( .A(n2194), .B(n10163), .Z(n2195) );
  NANDN U4170 ( .A(n6772), .B(n2195), .Z(n2196) );
  NANDN U4171 ( .A(n10168), .B(n2196), .Z(n2199) );
  NANDN U4172 ( .A(y[94]), .B(x[94]), .Z(n2198) );
  NANDN U4173 ( .A(y[95]), .B(x[95]), .Z(n2197) );
  AND U4174 ( .A(n2198), .B(n2197), .Z(n10169) );
  NAND U4175 ( .A(n2199), .B(n10169), .Z(n2200) );
  NANDN U4176 ( .A(n10172), .B(n2200), .Z(n2201) );
  NANDN U4177 ( .A(y[97]), .B(x[97]), .Z(n10178) );
  ANDN U4178 ( .B(x[96]), .A(y[96]), .Z(n10174) );
  ANDN U4179 ( .B(n10178), .A(n10174), .Z(n6776) );
  NAND U4180 ( .A(n2201), .B(n6776), .Z(n2202) );
  NANDN U4181 ( .A(n6779), .B(n2202), .Z(n2203) );
  AND U4182 ( .A(n6780), .B(n2203), .Z(n2208) );
  NANDN U4183 ( .A(x[101]), .B(y[101]), .Z(n2205) );
  NANDN U4184 ( .A(x[100]), .B(y[100]), .Z(n2204) );
  NAND U4185 ( .A(n2205), .B(n2204), .Z(n10189) );
  ANDN U4186 ( .B(y[99]), .A(x[99]), .Z(n10184) );
  NANDN U4187 ( .A(n2206), .B(n10184), .Z(n2207) );
  NANDN U4188 ( .A(n10189), .B(n2207), .Z(n6782) );
  OR U4189 ( .A(n2208), .B(n6782), .Z(n2211) );
  NANDN U4190 ( .A(y[101]), .B(x[101]), .Z(n2210) );
  NANDN U4191 ( .A(y[102]), .B(x[102]), .Z(n2209) );
  AND U4192 ( .A(n2210), .B(n2209), .Z(n10190) );
  NAND U4193 ( .A(n2211), .B(n10190), .Z(n2212) );
  NANDN U4194 ( .A(n10193), .B(n2212), .Z(n2213) );
  NANDN U4195 ( .A(n6786), .B(n2213), .Z(n2214) );
  NAND U4196 ( .A(n2215), .B(n2214), .Z(n2216) );
  AND U4197 ( .A(n6787), .B(n2216), .Z(n2218) );
  OR U4198 ( .A(n2218), .B(y[105]), .Z(n2217) );
  AND U4199 ( .A(n6569), .B(n2217), .Z(n2221) );
  XOR U4200 ( .A(y[105]), .B(n2218), .Z(n2219) );
  NAND U4201 ( .A(n2219), .B(x[105]), .Z(n2220) );
  NAND U4202 ( .A(n2221), .B(n2220), .Z(n2222) );
  NANDN U4203 ( .A(n10201), .B(n2222), .Z(n2223) );
  NANDN U4204 ( .A(y[107]), .B(x[107]), .Z(n10204) );
  NAND U4205 ( .A(n2223), .B(n10204), .Z(n2226) );
  NANDN U4206 ( .A(x[108]), .B(y[108]), .Z(n2225) );
  ANDN U4207 ( .B(n2225), .A(n2224), .Z(n10206) );
  NAND U4208 ( .A(n2226), .B(n10206), .Z(n2227) );
  NANDN U4209 ( .A(n6795), .B(n2227), .Z(n2228) );
  NANDN U4210 ( .A(n10211), .B(n2228), .Z(n2229) );
  AND U4211 ( .A(n10212), .B(n2229), .Z(n2230) );
  OR U4212 ( .A(n10214), .B(n2230), .Z(n2231) );
  NANDN U4213 ( .A(y[115]), .B(x[115]), .Z(n10217) );
  NAND U4214 ( .A(n2231), .B(n10217), .Z(n2234) );
  NANDN U4215 ( .A(x[116]), .B(y[116]), .Z(n2233) );
  ANDN U4216 ( .B(n2233), .A(n2232), .Z(n10221) );
  NAND U4217 ( .A(n2234), .B(n10221), .Z(n2235) );
  NANDN U4218 ( .A(n6802), .B(n2235), .Z(n2236) );
  NANDN U4219 ( .A(n10225), .B(n2236), .Z(n2239) );
  NANDN U4220 ( .A(y[120]), .B(x[120]), .Z(n2238) );
  NANDN U4221 ( .A(y[119]), .B(x[119]), .Z(n2237) );
  NAND U4222 ( .A(n2238), .B(n2237), .Z(n10227) );
  ANDN U4223 ( .B(n2239), .A(n10227), .Z(n2242) );
  NANDN U4224 ( .A(x[120]), .B(y[120]), .Z(n2241) );
  NANDN U4225 ( .A(x[121]), .B(y[121]), .Z(n2240) );
  AND U4226 ( .A(n2241), .B(n2240), .Z(n10228) );
  NANDN U4227 ( .A(n2242), .B(n10228), .Z(n2244) );
  NANDN U4228 ( .A(y[122]), .B(x[122]), .Z(n2243) );
  ANDN U4229 ( .B(x[121]), .A(y[121]), .Z(n6806) );
  ANDN U4230 ( .B(n2243), .A(n6806), .Z(n10230) );
  NAND U4231 ( .A(n2244), .B(n10230), .Z(n2245) );
  NANDN U4232 ( .A(n10232), .B(n2245), .Z(n2246) );
  NANDN U4233 ( .A(y[123]), .B(x[123]), .Z(n10235) );
  NAND U4234 ( .A(n2246), .B(n10235), .Z(n2248) );
  NANDN U4235 ( .A(x[124]), .B(y[124]), .Z(n2247) );
  ANDN U4236 ( .B(y[125]), .A(x[125]), .Z(n2253) );
  ANDN U4237 ( .B(n2247), .A(n2253), .Z(n10239) );
  NAND U4238 ( .A(n2248), .B(n10239), .Z(n2255) );
  NANDN U4239 ( .A(y[126]), .B(x[126]), .Z(n2250) );
  NANDN U4240 ( .A(y[125]), .B(x[125]), .Z(n2249) );
  AND U4241 ( .A(n2250), .B(n2249), .Z(n2252) );
  NANDN U4242 ( .A(y[127]), .B(x[127]), .Z(n2251) );
  NAND U4243 ( .A(n2252), .B(n2251), .Z(n10240) );
  ANDN U4244 ( .B(x[124]), .A(y[124]), .Z(n10234) );
  NANDN U4245 ( .A(n2253), .B(n10234), .Z(n2254) );
  NANDN U4246 ( .A(n10240), .B(n2254), .Z(n6816) );
  ANDN U4247 ( .B(n2255), .A(n6816), .Z(n2264) );
  NANDN U4248 ( .A(x[129]), .B(y[129]), .Z(n2257) );
  NANDN U4249 ( .A(x[128]), .B(y[128]), .Z(n2256) );
  AND U4250 ( .A(n2257), .B(n2256), .Z(n2263) );
  NANDN U4251 ( .A(x[126]), .B(y[126]), .Z(n2258) );
  NANDN U4252 ( .A(y[127]), .B(n2258), .Z(n2261) );
  XNOR U4253 ( .A(n2258), .B(y[127]), .Z(n2259) );
  NAND U4254 ( .A(n2259), .B(x[127]), .Z(n2260) );
  NAND U4255 ( .A(n2261), .B(n2260), .Z(n2262) );
  NAND U4256 ( .A(n2263), .B(n2262), .Z(n10243) );
  OR U4257 ( .A(n2264), .B(n10243), .Z(n2265) );
  NANDN U4258 ( .A(n10244), .B(n2265), .Z(n2274) );
  ANDN U4259 ( .B(y[133]), .A(x[133]), .Z(n2271) );
  NANDN U4260 ( .A(x[131]), .B(y[131]), .Z(n2269) );
  AND U4261 ( .A(y[130]), .B(n2266), .Z(n2267) );
  NANDN U4262 ( .A(x[130]), .B(n2267), .Z(n2268) );
  NAND U4263 ( .A(n2269), .B(n2268), .Z(n2270) );
  NOR U4264 ( .A(n2271), .B(n2270), .Z(n2273) );
  NANDN U4265 ( .A(x[132]), .B(y[132]), .Z(n2272) );
  AND U4266 ( .A(n2273), .B(n2272), .Z(n10246) );
  NAND U4267 ( .A(n2274), .B(n10246), .Z(n2275) );
  NANDN U4268 ( .A(n10248), .B(n2275), .Z(n2276) );
  NANDN U4269 ( .A(x[135]), .B(y[135]), .Z(n2278) );
  NAND U4270 ( .A(n2276), .B(n10252), .Z(n2279) );
  NANDN U4271 ( .A(y[134]), .B(x[134]), .Z(n10250) );
  ANDN U4272 ( .B(x[135]), .A(y[135]), .Z(n10254) );
  ANDN U4273 ( .B(n10250), .A(n10254), .Z(n2277) );
  ANDN U4274 ( .B(n2278), .A(n2277), .Z(n6823) );
  ANDN U4275 ( .B(n2279), .A(n6823), .Z(n2282) );
  NANDN U4276 ( .A(x[136]), .B(y[136]), .Z(n2281) );
  ANDN U4277 ( .B(n2281), .A(n2280), .Z(n10258) );
  NANDN U4278 ( .A(n2282), .B(n10258), .Z(n2283) );
  NANDN U4279 ( .A(n6827), .B(n2283), .Z(n2284) );
  NANDN U4280 ( .A(n10263), .B(n2284), .Z(n2285) );
  NANDN U4281 ( .A(n10265), .B(n2285), .Z(n2286) );
  NAND U4282 ( .A(n2286), .B(n10266), .Z(n2287) );
  AND U4283 ( .A(n10268), .B(n2287), .Z(n2288) );
  OR U4284 ( .A(n10271), .B(n2288), .Z(n2289) );
  NANDN U4285 ( .A(y[145]), .B(x[145]), .Z(n10274) );
  NAND U4286 ( .A(n2289), .B(n10274), .Z(n2292) );
  NANDN U4287 ( .A(x[146]), .B(y[146]), .Z(n2291) );
  ANDN U4288 ( .B(n2291), .A(n2290), .Z(n10276) );
  NAND U4289 ( .A(n2292), .B(n10276), .Z(n2293) );
  NANDN U4290 ( .A(n6839), .B(n2293), .Z(n2295) );
  NANDN U4291 ( .A(x[148]), .B(y[148]), .Z(n2294) );
  ANDN U4292 ( .B(y[149]), .A(x[149]), .Z(n2298) );
  ANDN U4293 ( .B(n2294), .A(n2298), .Z(n10282) );
  NAND U4294 ( .A(n2295), .B(n10282), .Z(n2300) );
  NANDN U4295 ( .A(y[150]), .B(x[150]), .Z(n2297) );
  NANDN U4296 ( .A(y[149]), .B(x[149]), .Z(n2296) );
  NAND U4297 ( .A(n2297), .B(n2296), .Z(n10284) );
  ANDN U4298 ( .B(x[148]), .A(y[148]), .Z(n10278) );
  NANDN U4299 ( .A(n2298), .B(n10278), .Z(n2299) );
  NANDN U4300 ( .A(n10284), .B(n2299), .Z(n6842) );
  ANDN U4301 ( .B(n2300), .A(n6842), .Z(n2303) );
  NANDN U4302 ( .A(x[150]), .B(y[150]), .Z(n2302) );
  NANDN U4303 ( .A(x[151]), .B(y[151]), .Z(n2301) );
  AND U4304 ( .A(n2302), .B(n2301), .Z(n10285) );
  NANDN U4305 ( .A(n2303), .B(n10285), .Z(n2304) );
  NANDN U4306 ( .A(y[151]), .B(x[151]), .Z(n10045) );
  NAND U4307 ( .A(n2304), .B(n10045), .Z(n2305) );
  NANDN U4308 ( .A(n10286), .B(n2305), .Z(n2306) );
  NANDN U4309 ( .A(n6847), .B(n2306), .Z(n2309) );
  NANDN U4310 ( .A(x[154]), .B(y[154]), .Z(n2308) );
  NANDN U4311 ( .A(x[155]), .B(y[155]), .Z(n2307) );
  AND U4312 ( .A(n2308), .B(n2307), .Z(n10288) );
  NAND U4313 ( .A(n2309), .B(n10288), .Z(n2312) );
  NANDN U4314 ( .A(y[156]), .B(x[156]), .Z(n2311) );
  NANDN U4315 ( .A(y[155]), .B(x[155]), .Z(n2310) );
  NAND U4316 ( .A(n2311), .B(n2310), .Z(n10289) );
  ANDN U4317 ( .B(n2312), .A(n10289), .Z(n2315) );
  NANDN U4318 ( .A(x[156]), .B(y[156]), .Z(n2314) );
  NANDN U4319 ( .A(x[157]), .B(y[157]), .Z(n2313) );
  AND U4320 ( .A(n2314), .B(n2313), .Z(n10290) );
  NANDN U4321 ( .A(n2315), .B(n10290), .Z(n2316) );
  NANDN U4322 ( .A(y[157]), .B(x[157]), .Z(n10292) );
  NAND U4323 ( .A(n2316), .B(n10292), .Z(n2319) );
  NANDN U4324 ( .A(x[158]), .B(y[158]), .Z(n2318) );
  ANDN U4325 ( .B(n2318), .A(n2317), .Z(n10293) );
  NAND U4326 ( .A(n2319), .B(n10293), .Z(n2320) );
  NANDN U4327 ( .A(n6854), .B(n2320), .Z(n2327) );
  NANDN U4328 ( .A(x[161]), .B(y[161]), .Z(n2322) );
  ANDN U4329 ( .B(y[162]), .A(x[162]), .Z(n2321) );
  ANDN U4330 ( .B(n2322), .A(n2321), .Z(n2326) );
  XNOR U4331 ( .A(y[161]), .B(x[161]), .Z(n2324) );
  ANDN U4332 ( .B(y[160]), .A(x[160]), .Z(n2323) );
  NAND U4333 ( .A(n2324), .B(n2323), .Z(n2325) );
  AND U4334 ( .A(n2326), .B(n2325), .Z(n10295) );
  NAND U4335 ( .A(n2327), .B(n10295), .Z(n2330) );
  NANDN U4336 ( .A(y[163]), .B(x[163]), .Z(n2329) );
  NANDN U4337 ( .A(y[162]), .B(x[162]), .Z(n2328) );
  NAND U4338 ( .A(n2329), .B(n2328), .Z(n10296) );
  ANDN U4339 ( .B(n2330), .A(n10296), .Z(n2335) );
  NANDN U4340 ( .A(x[164]), .B(y[164]), .Z(n2332) );
  NANDN U4341 ( .A(x[163]), .B(y[163]), .Z(n2331) );
  AND U4342 ( .A(n2332), .B(n2331), .Z(n2334) );
  NANDN U4343 ( .A(x[165]), .B(y[165]), .Z(n2333) );
  AND U4344 ( .A(n2334), .B(n2333), .Z(n10297) );
  NANDN U4345 ( .A(n2335), .B(n10297), .Z(n2336) );
  NANDN U4346 ( .A(n10298), .B(n2336), .Z(n2337) );
  NAND U4347 ( .A(n2337), .B(n10299), .Z(n2338) );
  NANDN U4348 ( .A(n10300), .B(n2338), .Z(n2339) );
  NANDN U4349 ( .A(n10302), .B(n2339), .Z(n2348) );
  NANDN U4350 ( .A(y[173]), .B(x[173]), .Z(n2341) );
  NANDN U4351 ( .A(y[172]), .B(x[172]), .Z(n2340) );
  AND U4352 ( .A(n2341), .B(n2340), .Z(n2347) );
  NANDN U4353 ( .A(y[170]), .B(x[170]), .Z(n2342) );
  NANDN U4354 ( .A(x[171]), .B(n2342), .Z(n2345) );
  XNOR U4355 ( .A(n2342), .B(x[171]), .Z(n2343) );
  NAND U4356 ( .A(n2343), .B(y[171]), .Z(n2344) );
  NAND U4357 ( .A(n2345), .B(n2344), .Z(n2346) );
  NAND U4358 ( .A(n2347), .B(n2346), .Z(n10305) );
  ANDN U4359 ( .B(n2348), .A(n10305), .Z(n2357) );
  NANDN U4360 ( .A(x[174]), .B(y[174]), .Z(n2349) );
  AND U4361 ( .A(n2350), .B(n2349), .Z(n2356) );
  NANDN U4362 ( .A(x[172]), .B(y[172]), .Z(n2351) );
  NANDN U4363 ( .A(y[173]), .B(n2351), .Z(n2354) );
  XNOR U4364 ( .A(n2351), .B(y[173]), .Z(n2352) );
  NAND U4365 ( .A(n2352), .B(x[173]), .Z(n2353) );
  NAND U4366 ( .A(n2354), .B(n2353), .Z(n2355) );
  NAND U4367 ( .A(n2356), .B(n2355), .Z(n10307) );
  OR U4368 ( .A(n2357), .B(n10307), .Z(n2358) );
  NANDN U4369 ( .A(n10309), .B(n2358), .Z(n2359) );
  NANDN U4370 ( .A(n10311), .B(n2359), .Z(n2360) );
  NANDN U4371 ( .A(y[177]), .B(x[177]), .Z(n10314) );
  NAND U4372 ( .A(n2360), .B(n10314), .Z(n2362) );
  NANDN U4373 ( .A(x[178]), .B(y[178]), .Z(n2361) );
  ANDN U4374 ( .B(y[179]), .A(x[179]), .Z(n2363) );
  ANDN U4375 ( .B(n2361), .A(n2363), .Z(n10316) );
  NAND U4376 ( .A(n2362), .B(n10316), .Z(n2365) );
  ANDN U4377 ( .B(x[179]), .A(y[179]), .Z(n10321) );
  ANDN U4378 ( .B(x[178]), .A(y[178]), .Z(n10312) );
  NANDN U4379 ( .A(n2363), .B(n10312), .Z(n2364) );
  NANDN U4380 ( .A(n10321), .B(n2364), .Z(n6878) );
  ANDN U4381 ( .B(n2365), .A(n6878), .Z(n2368) );
  NANDN U4382 ( .A(x[180]), .B(y[180]), .Z(n2367) );
  ANDN U4383 ( .B(n2367), .A(n2366), .Z(n10322) );
  NANDN U4384 ( .A(n2368), .B(n10322), .Z(n2369) );
  NANDN U4385 ( .A(n6880), .B(n2369), .Z(n2376) );
  NANDN U4386 ( .A(x[183]), .B(y[183]), .Z(n2371) );
  ANDN U4387 ( .B(y[184]), .A(x[184]), .Z(n2370) );
  ANDN U4388 ( .B(n2371), .A(n2370), .Z(n2375) );
  XNOR U4389 ( .A(y[183]), .B(x[183]), .Z(n2373) );
  ANDN U4390 ( .B(y[182]), .A(x[182]), .Z(n2372) );
  NAND U4391 ( .A(n2373), .B(n2372), .Z(n2374) );
  AND U4392 ( .A(n2375), .B(n2374), .Z(n10326) );
  NAND U4393 ( .A(n2376), .B(n10326), .Z(n2379) );
  NANDN U4394 ( .A(y[184]), .B(x[184]), .Z(n2378) );
  NANDN U4395 ( .A(y[185]), .B(x[185]), .Z(n2377) );
  AND U4396 ( .A(n2378), .B(n2377), .Z(n10328) );
  NAND U4397 ( .A(n2379), .B(n10328), .Z(n2380) );
  NANDN U4398 ( .A(n10331), .B(n2380), .Z(n2381) );
  NANDN U4399 ( .A(n10332), .B(n2381), .Z(n2384) );
  NANDN U4400 ( .A(x[188]), .B(y[188]), .Z(n2383) );
  ANDN U4401 ( .B(n2383), .A(n2382), .Z(n10336) );
  NAND U4402 ( .A(n2384), .B(n10336), .Z(n2385) );
  NANDN U4403 ( .A(n6887), .B(n2385), .Z(n2386) );
  AND U4404 ( .A(n10340), .B(n2386), .Z(n2387) );
  NANDN U4405 ( .A(y[191]), .B(x[191]), .Z(n10344) );
  NANDN U4406 ( .A(n2387), .B(n10344), .Z(n2390) );
  NANDN U4407 ( .A(x[192]), .B(y[192]), .Z(n2389) );
  ANDN U4408 ( .B(n2389), .A(n2388), .Z(n10346) );
  NAND U4409 ( .A(n2390), .B(n10346), .Z(n2391) );
  NANDN U4410 ( .A(n6893), .B(n2391), .Z(n2396) );
  NANDN U4411 ( .A(x[194]), .B(y[194]), .Z(n2392) );
  NANDN U4412 ( .A(n2392), .B(y[195]), .Z(n2395) );
  XNOR U4413 ( .A(n2392), .B(y[195]), .Z(n2393) );
  NANDN U4414 ( .A(x[195]), .B(n2393), .Z(n2394) );
  AND U4415 ( .A(n2395), .B(n2394), .Z(n10350) );
  NAND U4416 ( .A(n2396), .B(n10350), .Z(n2398) );
  ANDN U4417 ( .B(y[196]), .A(x[196]), .Z(n2397) );
  OR U4418 ( .A(n2398), .B(n2397), .Z(n2399) );
  NANDN U4419 ( .A(y[197]), .B(x[197]), .Z(n6565) );
  NAND U4420 ( .A(n2399), .B(n10352), .Z(n2400) );
  NANDN U4421 ( .A(x[197]), .B(y[197]), .Z(n6563) );
  NAND U4422 ( .A(n2400), .B(n6563), .Z(n2401) );
  NANDN U4423 ( .A(y[198]), .B(x[198]), .Z(n10356) );
  NAND U4424 ( .A(n2401), .B(n10356), .Z(n2404) );
  NANDN U4425 ( .A(x[198]), .B(y[198]), .Z(n2403) );
  NANDN U4426 ( .A(x[199]), .B(y[199]), .Z(n2402) );
  AND U4427 ( .A(n2403), .B(n2402), .Z(n10358) );
  NAND U4428 ( .A(n2404), .B(n10358), .Z(n2405) );
  AND U4429 ( .A(n10362), .B(n2405), .Z(n2408) );
  NANDN U4430 ( .A(x[200]), .B(y[200]), .Z(n2407) );
  ANDN U4431 ( .B(n2407), .A(n2406), .Z(n10364) );
  NANDN U4432 ( .A(n2408), .B(n10364), .Z(n2409) );
  NANDN U4433 ( .A(n6901), .B(n2409), .Z(n2412) );
  NANDN U4434 ( .A(x[202]), .B(y[202]), .Z(n2411) );
  ANDN U4435 ( .B(n2411), .A(n2410), .Z(n10370) );
  NAND U4436 ( .A(n2412), .B(n10370), .Z(n2413) );
  NANDN U4437 ( .A(n6905), .B(n2413), .Z(n2414) );
  NANDN U4438 ( .A(n10377), .B(n2414), .Z(n2418) );
  ANDN U4439 ( .B(x[206]), .A(y[206]), .Z(n10381) );
  NANDN U4440 ( .A(y[204]), .B(x[204]), .Z(n10374) );
  ANDN U4441 ( .B(x[205]), .A(y[205]), .Z(n10378) );
  ANDN U4442 ( .B(n10374), .A(n10378), .Z(n2416) );
  NANDN U4443 ( .A(n2416), .B(n2415), .Z(n2417) );
  NANDN U4444 ( .A(n10381), .B(n2417), .Z(n6908) );
  ANDN U4445 ( .B(n2418), .A(n6908), .Z(n2421) );
  NANDN U4446 ( .A(x[206]), .B(y[206]), .Z(n2420) );
  NANDN U4447 ( .A(x[207]), .B(y[207]), .Z(n2419) );
  AND U4448 ( .A(n2420), .B(n2419), .Z(n10382) );
  NANDN U4449 ( .A(n2421), .B(n10382), .Z(n2422) );
  NANDN U4450 ( .A(n10383), .B(n2422), .Z(n2423) );
  NANDN U4451 ( .A(n10384), .B(n2423), .Z(n2424) );
  NANDN U4452 ( .A(y[209]), .B(x[209]), .Z(n10043) );
  NAND U4453 ( .A(n2424), .B(n10043), .Z(n2425) );
  NANDN U4454 ( .A(n10385), .B(n2425), .Z(n2430) );
  NANDN U4455 ( .A(y[212]), .B(x[212]), .Z(n2427) );
  NANDN U4456 ( .A(y[211]), .B(x[211]), .Z(n2426) );
  NAND U4457 ( .A(n2427), .B(n2426), .Z(n10386) );
  NANDN U4458 ( .A(y[210]), .B(x[210]), .Z(n10042) );
  NANDN U4459 ( .A(n10042), .B(n2428), .Z(n2429) );
  NANDN U4460 ( .A(n10386), .B(n2429), .Z(n6921) );
  ANDN U4461 ( .B(n2430), .A(n6921), .Z(n2433) );
  NANDN U4462 ( .A(x[212]), .B(y[212]), .Z(n2432) );
  NANDN U4463 ( .A(x[213]), .B(y[213]), .Z(n2431) );
  AND U4464 ( .A(n2432), .B(n2431), .Z(n10387) );
  NANDN U4465 ( .A(n2433), .B(n10387), .Z(n2434) );
  NANDN U4466 ( .A(n10388), .B(n2434), .Z(n2437) );
  NANDN U4467 ( .A(x[214]), .B(y[214]), .Z(n2436) );
  NANDN U4468 ( .A(x[215]), .B(y[215]), .Z(n2435) );
  AND U4469 ( .A(n2436), .B(n2435), .Z(n10389) );
  NAND U4470 ( .A(n2437), .B(n10389), .Z(n2438) );
  NANDN U4471 ( .A(n10390), .B(n2438), .Z(n2441) );
  NANDN U4472 ( .A(x[216]), .B(y[216]), .Z(n2440) );
  NANDN U4473 ( .A(x[217]), .B(y[217]), .Z(n2439) );
  AND U4474 ( .A(n2440), .B(n2439), .Z(n10391) );
  NAND U4475 ( .A(n2441), .B(n10391), .Z(n2442) );
  NANDN U4476 ( .A(y[217]), .B(x[217]), .Z(n10041) );
  NAND U4477 ( .A(n2442), .B(n10041), .Z(n2443) );
  NANDN U4478 ( .A(n10392), .B(n2443), .Z(n2444) );
  NANDN U4479 ( .A(n6929), .B(n2444), .Z(n2452) );
  NANDN U4480 ( .A(x[223]), .B(y[223]), .Z(n2453) );
  NANDN U4481 ( .A(x[222]), .B(y[222]), .Z(n2445) );
  AND U4482 ( .A(n2453), .B(n2445), .Z(n2451) );
  ANDN U4483 ( .B(y[220]), .A(x[220]), .Z(n2446) );
  OR U4484 ( .A(n2446), .B(y[221]), .Z(n2449) );
  XOR U4485 ( .A(y[221]), .B(n2446), .Z(n2447) );
  NAND U4486 ( .A(n2447), .B(x[221]), .Z(n2448) );
  NAND U4487 ( .A(n2449), .B(n2448), .Z(n2450) );
  NAND U4488 ( .A(n2451), .B(n2450), .Z(n10394) );
  ANDN U4489 ( .B(n2452), .A(n10394), .Z(n2461) );
  ANDN U4490 ( .B(x[225]), .A(y[225]), .Z(n2458) );
  NANDN U4491 ( .A(y[223]), .B(x[223]), .Z(n2456) );
  AND U4492 ( .A(x[222]), .B(n2453), .Z(n2454) );
  NANDN U4493 ( .A(y[222]), .B(n2454), .Z(n2455) );
  NAND U4494 ( .A(n2456), .B(n2455), .Z(n2457) );
  NOR U4495 ( .A(n2458), .B(n2457), .Z(n2460) );
  NANDN U4496 ( .A(y[224]), .B(x[224]), .Z(n2459) );
  AND U4497 ( .A(n2460), .B(n2459), .Z(n10395) );
  NANDN U4498 ( .A(n2461), .B(n10395), .Z(n2462) );
  NANDN U4499 ( .A(n10398), .B(n2462), .Z(n2463) );
  NANDN U4500 ( .A(n10399), .B(n2463), .Z(n2464) );
  NANDN U4501 ( .A(n10402), .B(n2464), .Z(n2465) );
  NANDN U4502 ( .A(n10404), .B(n2465), .Z(n2470) );
  XNOR U4503 ( .A(y[233]), .B(x[233]), .Z(n2467) );
  NANDN U4504 ( .A(x[232]), .B(y[232]), .Z(n2466) );
  NAND U4505 ( .A(n2467), .B(n2466), .Z(n2468) );
  AND U4506 ( .A(n2469), .B(n2468), .Z(n10406) );
  ANDN U4507 ( .B(n2470), .A(n10406), .Z(n2473) );
  NANDN U4508 ( .A(y[234]), .B(x[234]), .Z(n2471) );
  NAND U4509 ( .A(n2472), .B(n2471), .Z(n10408) );
  OR U4510 ( .A(n2473), .B(n10408), .Z(n2474) );
  NANDN U4511 ( .A(n10410), .B(n2474), .Z(n2475) );
  NANDN U4512 ( .A(n10411), .B(n2475), .Z(n2476) );
  NANDN U4513 ( .A(n10414), .B(n2476), .Z(n2479) );
  NANDN U4514 ( .A(y[241]), .B(x[241]), .Z(n2478) );
  NANDN U4515 ( .A(y[240]), .B(x[240]), .Z(n2477) );
  AND U4516 ( .A(n2478), .B(n2477), .Z(n10415) );
  NAND U4517 ( .A(n2479), .B(n10415), .Z(n2480) );
  AND U4518 ( .A(n10417), .B(n2480), .Z(n2483) );
  NANDN U4519 ( .A(y[242]), .B(x[242]), .Z(n2482) );
  AND U4520 ( .A(n2482), .B(n2481), .Z(n10419) );
  NANDN U4521 ( .A(n2483), .B(n10419), .Z(n2484) );
  NANDN U4522 ( .A(n10422), .B(n2484), .Z(n2485) );
  NANDN U4523 ( .A(n10423), .B(n2485), .Z(n2486) );
  NANDN U4524 ( .A(n10425), .B(n2486), .Z(n2487) );
  NANDN U4525 ( .A(n10428), .B(n2487), .Z(n2496) );
  NANDN U4526 ( .A(x[253]), .B(y[253]), .Z(n2489) );
  NANDN U4527 ( .A(x[252]), .B(y[252]), .Z(n2488) );
  AND U4528 ( .A(n2489), .B(n2488), .Z(n2495) );
  NANDN U4529 ( .A(x[250]), .B(y[250]), .Z(n2490) );
  NANDN U4530 ( .A(y[251]), .B(n2490), .Z(n2493) );
  XNOR U4531 ( .A(n2490), .B(y[251]), .Z(n2491) );
  NAND U4532 ( .A(n2491), .B(x[251]), .Z(n2492) );
  NAND U4533 ( .A(n2493), .B(n2492), .Z(n2494) );
  NAND U4534 ( .A(n2495), .B(n2494), .Z(n10430) );
  ANDN U4535 ( .B(n2496), .A(n10430), .Z(n2497) );
  OR U4536 ( .A(n10432), .B(n2497), .Z(n2498) );
  NANDN U4537 ( .A(n6965), .B(n2498), .Z(n2508) );
  NANDN U4538 ( .A(y[256]), .B(x[256]), .Z(n2499) );
  NANDN U4539 ( .A(n2499), .B(x[257]), .Z(n2502) );
  XNOR U4540 ( .A(n2499), .B(x[257]), .Z(n2500) );
  NANDN U4541 ( .A(y[257]), .B(n2500), .Z(n2501) );
  NAND U4542 ( .A(n2502), .B(n2501), .Z(n2503) );
  ANDN U4543 ( .B(x[259]), .A(y[259]), .Z(n2506) );
  NOR U4544 ( .A(n2503), .B(n2506), .Z(n2505) );
  NANDN U4545 ( .A(y[258]), .B(x[258]), .Z(n2504) );
  AND U4546 ( .A(n2505), .B(n2504), .Z(n10436) );
  ANDN U4547 ( .B(n2507), .A(n2506), .Z(n10437) );
  OR U4548 ( .A(n10436), .B(n10437), .Z(n6966) );
  NAND U4549 ( .A(n2508), .B(n6966), .Z(n2509) );
  NANDN U4550 ( .A(n6969), .B(n2509), .Z(n2510) );
  NANDN U4551 ( .A(n6971), .B(n2510), .Z(n2511) );
  AND U4552 ( .A(n10449), .B(n2511), .Z(n2514) );
  NANDN U4553 ( .A(y[262]), .B(x[262]), .Z(n10447) );
  ANDN U4554 ( .B(x[263]), .A(y[263]), .Z(n10451) );
  ANDN U4555 ( .B(n10447), .A(n10451), .Z(n2513) );
  NANDN U4556 ( .A(n2513), .B(n2512), .Z(n6973) );
  NANDN U4557 ( .A(n2514), .B(n6973), .Z(n2517) );
  NANDN U4558 ( .A(x[264]), .B(y[264]), .Z(n2516) );
  ANDN U4559 ( .B(n2516), .A(n2515), .Z(n10455) );
  NAND U4560 ( .A(n2517), .B(n10455), .Z(n2518) );
  NANDN U4561 ( .A(n6977), .B(n2518), .Z(n2519) );
  NANDN U4562 ( .A(n10460), .B(n2519), .Z(n2520) );
  NANDN U4563 ( .A(n10462), .B(n2520), .Z(n2525) );
  XNOR U4564 ( .A(y[271]), .B(x[271]), .Z(n2522) );
  NANDN U4565 ( .A(x[270]), .B(y[270]), .Z(n2521) );
  NAND U4566 ( .A(n2522), .B(n2521), .Z(n2523) );
  AND U4567 ( .A(n2524), .B(n2523), .Z(n10464) );
  ANDN U4568 ( .B(n2525), .A(n10464), .Z(n2526) );
  NANDN U4569 ( .A(y[272]), .B(x[272]), .Z(n10465) );
  NANDN U4570 ( .A(n2526), .B(n10465), .Z(n2527) );
  ANDN U4571 ( .B(y[273]), .A(x[273]), .Z(n6985) );
  ANDN U4572 ( .B(y[272]), .A(x[272]), .Z(n6980) );
  NOR U4573 ( .A(n6985), .B(n6980), .Z(n10467) );
  NAND U4574 ( .A(n2527), .B(n10467), .Z(n2528) );
  NANDN U4575 ( .A(y[273]), .B(x[273]), .Z(n10471) );
  NAND U4576 ( .A(n2528), .B(n10471), .Z(n2529) );
  NANDN U4577 ( .A(x[274]), .B(y[274]), .Z(n10475) );
  NAND U4578 ( .A(n2529), .B(n10475), .Z(n2530) );
  ANDN U4579 ( .B(x[274]), .A(y[274]), .Z(n10469) );
  ANDN U4580 ( .B(x[275]), .A(y[275]), .Z(n10480) );
  NOR U4581 ( .A(n10469), .B(n10480), .Z(n6988) );
  NAND U4582 ( .A(n2530), .B(n6988), .Z(n2531) );
  AND U4583 ( .A(n10474), .B(n2531), .Z(n2534) );
  NANDN U4584 ( .A(y[276]), .B(x[276]), .Z(n2532) );
  AND U4585 ( .A(n2533), .B(n2532), .Z(n10478) );
  NANDN U4586 ( .A(n2534), .B(n10478), .Z(n2535) );
  AND U4587 ( .A(n2536), .B(n2535), .Z(n2537) );
  NOR U4588 ( .A(n10488), .B(n2537), .Z(n2539) );
  NANDN U4589 ( .A(y[278]), .B(x[278]), .Z(n10483) );
  NANDN U4590 ( .A(n10483), .B(n2538), .Z(n6998) );
  NAND U4591 ( .A(n2539), .B(n6998), .Z(n2541) );
  NANDN U4592 ( .A(x[280]), .B(y[280]), .Z(n2540) );
  NANDN U4593 ( .A(x[281]), .B(y[281]), .Z(n7008) );
  NAND U4594 ( .A(n2540), .B(n7008), .Z(n10490) );
  ANDN U4595 ( .B(n2541), .A(n10490), .Z(n2542) );
  NANDN U4596 ( .A(y[281]), .B(x[281]), .Z(n10492) );
  NANDN U4597 ( .A(n2542), .B(n10492), .Z(n2545) );
  NANDN U4598 ( .A(x[282]), .B(y[282]), .Z(n2544) );
  ANDN U4599 ( .B(n2544), .A(n2543), .Z(n10495) );
  NAND U4600 ( .A(n2545), .B(n10495), .Z(n2546) );
  NANDN U4601 ( .A(n7011), .B(n2546), .Z(n2547) );
  NANDN U4602 ( .A(n10499), .B(n2547), .Z(n2548) );
  NANDN U4603 ( .A(y[285]), .B(x[285]), .Z(n10502) );
  NAND U4604 ( .A(n2548), .B(n10502), .Z(n2549) );
  AND U4605 ( .A(n10506), .B(n2549), .Z(n2554) );
  NANDN U4606 ( .A(y[288]), .B(x[288]), .Z(n2551) );
  NANDN U4607 ( .A(y[287]), .B(x[287]), .Z(n2550) );
  NAND U4608 ( .A(n2551), .B(n2550), .Z(n10508) );
  ANDN U4609 ( .B(x[286]), .A(y[286]), .Z(n10501) );
  NANDN U4610 ( .A(n2552), .B(n10501), .Z(n2553) );
  NANDN U4611 ( .A(n10508), .B(n2553), .Z(n7016) );
  OR U4612 ( .A(n2554), .B(n7016), .Z(n2555) );
  NANDN U4613 ( .A(n10510), .B(n2555), .Z(n2558) );
  NANDN U4614 ( .A(y[289]), .B(x[289]), .Z(n2557) );
  NANDN U4615 ( .A(y[290]), .B(x[290]), .Z(n2556) );
  AND U4616 ( .A(n2557), .B(n2556), .Z(n10511) );
  NAND U4617 ( .A(n2558), .B(n10511), .Z(n2559) );
  NANDN U4618 ( .A(n10514), .B(n2559), .Z(n2562) );
  NANDN U4619 ( .A(y[291]), .B(x[291]), .Z(n2561) );
  NANDN U4620 ( .A(y[292]), .B(x[292]), .Z(n2560) );
  AND U4621 ( .A(n2561), .B(n2560), .Z(n10515) );
  NAND U4622 ( .A(n2562), .B(n10515), .Z(n2565) );
  NANDN U4623 ( .A(x[293]), .B(y[293]), .Z(n2564) );
  NANDN U4624 ( .A(x[292]), .B(y[292]), .Z(n2563) );
  NAND U4625 ( .A(n2564), .B(n2563), .Z(n10517) );
  ANDN U4626 ( .B(n2565), .A(n10517), .Z(n2566) );
  NANDN U4627 ( .A(y[293]), .B(x[293]), .Z(n10520) );
  NANDN U4628 ( .A(n2566), .B(n10520), .Z(n2569) );
  NANDN U4629 ( .A(x[294]), .B(y[294]), .Z(n2568) );
  ANDN U4630 ( .B(n2568), .A(n2567), .Z(n10524) );
  NAND U4631 ( .A(n2569), .B(n10524), .Z(n2570) );
  NANDN U4632 ( .A(n7025), .B(n2570), .Z(n2571) );
  NANDN U4633 ( .A(n10528), .B(n2571), .Z(n2572) );
  NANDN U4634 ( .A(y[297]), .B(x[297]), .Z(n10529) );
  NAND U4635 ( .A(n2572), .B(n10529), .Z(n2573) );
  AND U4636 ( .A(n10533), .B(n2573), .Z(n2577) );
  NANDN U4637 ( .A(y[298]), .B(x[298]), .Z(n2574) );
  ANDN U4638 ( .B(x[299]), .A(y[299]), .Z(n10536) );
  ANDN U4639 ( .B(n2574), .A(n10536), .Z(n2576) );
  NANDN U4640 ( .A(n2576), .B(n2575), .Z(n7029) );
  NANDN U4641 ( .A(n2577), .B(n7029), .Z(n2580) );
  NANDN U4642 ( .A(x[300]), .B(y[300]), .Z(n2579) );
  ANDN U4643 ( .B(n2579), .A(n2578), .Z(n10539) );
  NAND U4644 ( .A(n2580), .B(n10539), .Z(n2581) );
  NANDN U4645 ( .A(n7033), .B(n2581), .Z(n2582) );
  NANDN U4646 ( .A(n10544), .B(n2582), .Z(n2583) );
  NANDN U4647 ( .A(y[303]), .B(x[303]), .Z(n10039) );
  NAND U4648 ( .A(n2583), .B(n10039), .Z(n2584) );
  AND U4649 ( .A(n10547), .B(n2584), .Z(n2587) );
  ANDN U4650 ( .B(x[305]), .A(y[305]), .Z(n10549) );
  ANDN U4651 ( .B(x[304]), .A(y[304]), .Z(n10038) );
  NANDN U4652 ( .A(n2585), .B(n10038), .Z(n2586) );
  NANDN U4653 ( .A(n10549), .B(n2586), .Z(n7038) );
  OR U4654 ( .A(n2587), .B(n7038), .Z(n2588) );
  NANDN U4655 ( .A(x[307]), .B(y[307]), .Z(n2589) );
  NAND U4656 ( .A(n2588), .B(n10553), .Z(n2591) );
  NANDN U4657 ( .A(y[306]), .B(x[306]), .Z(n10551) );
  ANDN U4658 ( .B(x[307]), .A(y[307]), .Z(n10555) );
  ANDN U4659 ( .B(n10551), .A(n10555), .Z(n2590) );
  NANDN U4660 ( .A(n2590), .B(n2589), .Z(n7040) );
  NAND U4661 ( .A(n2591), .B(n7040), .Z(n2594) );
  NANDN U4662 ( .A(x[308]), .B(y[308]), .Z(n2593) );
  ANDN U4663 ( .B(n2593), .A(n2592), .Z(n10559) );
  NAND U4664 ( .A(n2594), .B(n10559), .Z(n2595) );
  NANDN U4665 ( .A(n7044), .B(n2595), .Z(n2604) );
  NANDN U4666 ( .A(x[313]), .B(y[313]), .Z(n2597) );
  NANDN U4667 ( .A(x[312]), .B(y[312]), .Z(n2596) );
  AND U4668 ( .A(n2597), .B(n2596), .Z(n2603) );
  NANDN U4669 ( .A(x[310]), .B(y[310]), .Z(n2598) );
  NANDN U4670 ( .A(y[311]), .B(n2598), .Z(n2601) );
  XNOR U4671 ( .A(n2598), .B(y[311]), .Z(n2599) );
  NAND U4672 ( .A(n2599), .B(x[311]), .Z(n2600) );
  NAND U4673 ( .A(n2601), .B(n2600), .Z(n2602) );
  NAND U4674 ( .A(n2603), .B(n2602), .Z(n10564) );
  ANDN U4675 ( .B(n2604), .A(n10564), .Z(n2613) );
  NANDN U4676 ( .A(y[315]), .B(x[315]), .Z(n2606) );
  NANDN U4677 ( .A(y[314]), .B(x[314]), .Z(n2605) );
  AND U4678 ( .A(n2606), .B(n2605), .Z(n2612) );
  NANDN U4679 ( .A(y[312]), .B(x[312]), .Z(n2607) );
  NANDN U4680 ( .A(x[313]), .B(n2607), .Z(n2610) );
  XNOR U4681 ( .A(n2607), .B(x[313]), .Z(n2608) );
  NAND U4682 ( .A(n2608), .B(y[313]), .Z(n2609) );
  NAND U4683 ( .A(n2610), .B(n2609), .Z(n2611) );
  NAND U4684 ( .A(n2612), .B(n2611), .Z(n10566) );
  OR U4685 ( .A(n2613), .B(n10566), .Z(n2622) );
  NANDN U4686 ( .A(x[317]), .B(y[317]), .Z(n2615) );
  NANDN U4687 ( .A(x[316]), .B(y[316]), .Z(n2614) );
  AND U4688 ( .A(n2615), .B(n2614), .Z(n2621) );
  NANDN U4689 ( .A(x[314]), .B(y[314]), .Z(n2616) );
  NANDN U4690 ( .A(y[315]), .B(n2616), .Z(n2619) );
  XNOR U4691 ( .A(n2616), .B(y[315]), .Z(n2617) );
  NAND U4692 ( .A(n2617), .B(x[315]), .Z(n2618) );
  NAND U4693 ( .A(n2619), .B(n2618), .Z(n2620) );
  AND U4694 ( .A(n2621), .B(n2620), .Z(n10567) );
  NAND U4695 ( .A(n2622), .B(n10567), .Z(n2623) );
  NANDN U4696 ( .A(n10570), .B(n2623), .Z(n2624) );
  NAND U4697 ( .A(n2625), .B(n2624), .Z(n2626) );
  NANDN U4698 ( .A(n10573), .B(n2626), .Z(n2627) );
  NANDN U4699 ( .A(x[321]), .B(y[321]), .Z(n6559) );
  NAND U4700 ( .A(n2627), .B(n6559), .Z(n2628) );
  NANDN U4701 ( .A(y[322]), .B(x[322]), .Z(n10578) );
  NAND U4702 ( .A(n2628), .B(n10578), .Z(n2629) );
  AND U4703 ( .A(n10579), .B(n2629), .Z(n2630) );
  NANDN U4704 ( .A(y[323]), .B(x[323]), .Z(n10037) );
  NANDN U4705 ( .A(n2630), .B(n10037), .Z(n2633) );
  NANDN U4706 ( .A(x[324]), .B(y[324]), .Z(n2632) );
  ANDN U4707 ( .B(n2632), .A(n2631), .Z(n10583) );
  NAND U4708 ( .A(n2633), .B(n10583), .Z(n2634) );
  NANDN U4709 ( .A(n7057), .B(n2634), .Z(n2639) );
  NANDN U4710 ( .A(x[328]), .B(y[328]), .Z(n10593) );
  XNOR U4711 ( .A(y[327]), .B(x[327]), .Z(n2636) );
  NANDN U4712 ( .A(x[326]), .B(y[326]), .Z(n2635) );
  NAND U4713 ( .A(n2636), .B(n2635), .Z(n2637) );
  AND U4714 ( .A(n2638), .B(n2637), .Z(n10589) );
  ANDN U4715 ( .B(n10593), .A(n10589), .Z(n7058) );
  NAND U4716 ( .A(n2639), .B(n7058), .Z(n2641) );
  NANDN U4717 ( .A(y[328]), .B(x[328]), .Z(n2640) );
  NANDN U4718 ( .A(y[329]), .B(x[329]), .Z(n10592) );
  AND U4719 ( .A(n2640), .B(n10592), .Z(n10591) );
  NAND U4720 ( .A(n2641), .B(n10591), .Z(n2642) );
  AND U4721 ( .A(n10594), .B(n2642), .Z(n2643) );
  NANDN U4722 ( .A(x[330]), .B(y[330]), .Z(n10034) );
  NAND U4723 ( .A(n2643), .B(n10034), .Z(n2644) );
  NANDN U4724 ( .A(n7064), .B(n2644), .Z(n2645) );
  AND U4725 ( .A(n10035), .B(n2645), .Z(n2646) );
  NANDN U4726 ( .A(y[332]), .B(x[332]), .Z(n10598) );
  NANDN U4727 ( .A(n2646), .B(n10598), .Z(n2647) );
  ANDN U4728 ( .B(y[333]), .A(x[333]), .Z(n6555) );
  ANDN U4729 ( .B(y[332]), .A(x[332]), .Z(n6556) );
  NOR U4730 ( .A(n6555), .B(n6556), .Z(n10599) );
  NAND U4731 ( .A(n2647), .B(n10599), .Z(n2648) );
  NANDN U4732 ( .A(y[333]), .B(x[333]), .Z(n10601) );
  NAND U4733 ( .A(n2648), .B(n10601), .Z(n2651) );
  NANDN U4734 ( .A(x[334]), .B(y[334]), .Z(n2650) );
  ANDN U4735 ( .B(n2650), .A(n2649), .Z(n10602) );
  NAND U4736 ( .A(n2651), .B(n10602), .Z(n2652) );
  NANDN U4737 ( .A(n7072), .B(n2652), .Z(n2653) );
  AND U4738 ( .A(n10605), .B(n2653), .Z(n2658) );
  NANDN U4739 ( .A(y[338]), .B(x[338]), .Z(n2655) );
  NANDN U4740 ( .A(y[337]), .B(x[337]), .Z(n2654) );
  NAND U4741 ( .A(n2655), .B(n2654), .Z(n10606) );
  ANDN U4742 ( .B(x[336]), .A(y[336]), .Z(n10603) );
  NANDN U4743 ( .A(n2656), .B(n10603), .Z(n2657) );
  NANDN U4744 ( .A(n10606), .B(n2657), .Z(n7075) );
  OR U4745 ( .A(n2658), .B(n7075), .Z(n2659) );
  NANDN U4746 ( .A(n10607), .B(n2659), .Z(n2660) );
  NANDN U4747 ( .A(y[339]), .B(x[339]), .Z(n10608) );
  NAND U4748 ( .A(n2660), .B(n10608), .Z(n2663) );
  NANDN U4749 ( .A(x[340]), .B(y[340]), .Z(n2662) );
  ANDN U4750 ( .B(n2662), .A(n2661), .Z(n10611) );
  NAND U4751 ( .A(n2663), .B(n10611), .Z(n2664) );
  NANDN U4752 ( .A(n7080), .B(n2664), .Z(n2665) );
  AND U4753 ( .A(n10616), .B(n2665), .Z(n2666) );
  NANDN U4754 ( .A(y[343]), .B(x[343]), .Z(n10618) );
  NANDN U4755 ( .A(n2666), .B(n10618), .Z(n2669) );
  NANDN U4756 ( .A(x[344]), .B(y[344]), .Z(n2668) );
  ANDN U4757 ( .B(n2668), .A(n2667), .Z(n10622) );
  NAND U4758 ( .A(n2669), .B(n10622), .Z(n2670) );
  NANDN U4759 ( .A(n7085), .B(n2670), .Z(n2671) );
  NANDN U4760 ( .A(n10626), .B(n2671), .Z(n2672) );
  NANDN U4761 ( .A(n10628), .B(n2672), .Z(n2673) );
  NANDN U4762 ( .A(x[351]), .B(y[351]), .Z(n2677) );
  ANDN U4763 ( .B(n2673), .A(n10632), .Z(n2680) );
  NANDN U4764 ( .A(y[353]), .B(x[353]), .Z(n2675) );
  NANDN U4765 ( .A(y[352]), .B(x[352]), .Z(n2674) );
  NAND U4766 ( .A(n2675), .B(n2674), .Z(n10635) );
  NANDN U4767 ( .A(y[350]), .B(x[350]), .Z(n2676) );
  ANDN U4768 ( .B(x[351]), .A(y[351]), .Z(n10634) );
  ANDN U4769 ( .B(n2676), .A(n10634), .Z(n2678) );
  NANDN U4770 ( .A(n2678), .B(n2677), .Z(n2679) );
  NANDN U4771 ( .A(n10635), .B(n2679), .Z(n7089) );
  OR U4772 ( .A(n2680), .B(n7089), .Z(n2689) );
  NANDN U4773 ( .A(x[355]), .B(y[355]), .Z(n2682) );
  NANDN U4774 ( .A(x[354]), .B(y[354]), .Z(n2681) );
  AND U4775 ( .A(n2682), .B(n2681), .Z(n2688) );
  NANDN U4776 ( .A(x[352]), .B(y[352]), .Z(n2683) );
  NANDN U4777 ( .A(y[353]), .B(n2683), .Z(n2686) );
  XNOR U4778 ( .A(n2683), .B(y[353]), .Z(n2684) );
  NAND U4779 ( .A(n2684), .B(x[353]), .Z(n2685) );
  NAND U4780 ( .A(n2686), .B(n2685), .Z(n2687) );
  AND U4781 ( .A(n2688), .B(n2687), .Z(n10637) );
  NAND U4782 ( .A(n2689), .B(n10637), .Z(n2690) );
  NANDN U4783 ( .A(n10639), .B(n2690), .Z(n2695) );
  NANDN U4784 ( .A(x[356]), .B(y[356]), .Z(n2691) );
  NANDN U4785 ( .A(n2691), .B(y[357]), .Z(n2694) );
  XNOR U4786 ( .A(n2691), .B(y[357]), .Z(n2692) );
  NANDN U4787 ( .A(x[357]), .B(n2692), .Z(n2693) );
  AND U4788 ( .A(n2694), .B(n2693), .Z(n10641) );
  NAND U4789 ( .A(n2695), .B(n10641), .Z(n2696) );
  NANDN U4790 ( .A(n10644), .B(n2696), .Z(n2703) );
  NANDN U4791 ( .A(x[358]), .B(y[358]), .Z(n7094) );
  NANDN U4792 ( .A(n7094), .B(n2697), .Z(n2702) );
  NANDN U4793 ( .A(x[360]), .B(y[360]), .Z(n2699) );
  NANDN U4794 ( .A(x[359]), .B(y[359]), .Z(n2698) );
  AND U4795 ( .A(n2699), .B(n2698), .Z(n2701) );
  NANDN U4796 ( .A(x[361]), .B(y[361]), .Z(n2700) );
  AND U4797 ( .A(n2701), .B(n2700), .Z(n7097) );
  NAND U4798 ( .A(n2702), .B(n7097), .Z(n10646) );
  ANDN U4799 ( .B(n2703), .A(n10646), .Z(n2712) );
  NANDN U4800 ( .A(y[363]), .B(x[363]), .Z(n2705) );
  NANDN U4801 ( .A(y[362]), .B(x[362]), .Z(n2704) );
  AND U4802 ( .A(n2705), .B(n2704), .Z(n2711) );
  NANDN U4803 ( .A(y[360]), .B(x[360]), .Z(n2706) );
  NANDN U4804 ( .A(x[361]), .B(n2706), .Z(n2709) );
  XNOR U4805 ( .A(n2706), .B(x[361]), .Z(n2707) );
  NAND U4806 ( .A(n2707), .B(y[361]), .Z(n2708) );
  NAND U4807 ( .A(n2709), .B(n2708), .Z(n2710) );
  NAND U4808 ( .A(n2711), .B(n2710), .Z(n10648) );
  OR U4809 ( .A(n2712), .B(n10648), .Z(n2721) );
  NANDN U4810 ( .A(x[365]), .B(y[365]), .Z(n2714) );
  NANDN U4811 ( .A(x[364]), .B(y[364]), .Z(n2713) );
  AND U4812 ( .A(n2714), .B(n2713), .Z(n2720) );
  NANDN U4813 ( .A(x[362]), .B(y[362]), .Z(n2715) );
  NANDN U4814 ( .A(y[363]), .B(n2715), .Z(n2718) );
  XNOR U4815 ( .A(n2715), .B(y[363]), .Z(n2716) );
  NAND U4816 ( .A(n2716), .B(x[363]), .Z(n2717) );
  NAND U4817 ( .A(n2718), .B(n2717), .Z(n2719) );
  NAND U4818 ( .A(n2720), .B(n2719), .Z(n10649) );
  ANDN U4819 ( .B(n2721), .A(n10649), .Z(n2726) );
  NANDN U4820 ( .A(y[364]), .B(x[364]), .Z(n2722) );
  NANDN U4821 ( .A(n2722), .B(x[365]), .Z(n2725) );
  XNOR U4822 ( .A(n2722), .B(x[365]), .Z(n2723) );
  NANDN U4823 ( .A(y[365]), .B(n2723), .Z(n2724) );
  AND U4824 ( .A(n2725), .B(n2724), .Z(n10651) );
  NANDN U4825 ( .A(n2726), .B(n10651), .Z(n2727) );
  NANDN U4826 ( .A(n10032), .B(n2727), .Z(n2728) );
  NANDN U4827 ( .A(n7104), .B(n2728), .Z(n2729) );
  NANDN U4828 ( .A(n10653), .B(n2729), .Z(n2730) );
  NANDN U4829 ( .A(y[369]), .B(x[369]), .Z(n10655) );
  NAND U4830 ( .A(n2730), .B(n10655), .Z(n2731) );
  AND U4831 ( .A(n10656), .B(n2731), .Z(n2734) );
  ANDN U4832 ( .B(x[371]), .A(y[371]), .Z(n10657) );
  ANDN U4833 ( .B(x[370]), .A(y[370]), .Z(n10654) );
  NANDN U4834 ( .A(n2732), .B(n10654), .Z(n2733) );
  NANDN U4835 ( .A(n10657), .B(n2733), .Z(n7109) );
  OR U4836 ( .A(n2734), .B(n7109), .Z(n2735) );
  NANDN U4837 ( .A(n10658), .B(n2735), .Z(n2736) );
  NANDN U4838 ( .A(n7112), .B(n2736), .Z(n2737) );
  NANDN U4839 ( .A(n10661), .B(n2737), .Z(n2738) );
  NANDN U4840 ( .A(y[375]), .B(x[375]), .Z(n10663) );
  NAND U4841 ( .A(n2738), .B(n10663), .Z(n2739) );
  AND U4842 ( .A(n10665), .B(n2739), .Z(n2744) );
  NANDN U4843 ( .A(y[378]), .B(x[378]), .Z(n2741) );
  NANDN U4844 ( .A(y[377]), .B(x[377]), .Z(n2740) );
  NAND U4845 ( .A(n2741), .B(n2740), .Z(n10667) );
  ANDN U4846 ( .B(x[376]), .A(y[376]), .Z(n10662) );
  NANDN U4847 ( .A(n2742), .B(n10662), .Z(n2743) );
  NANDN U4848 ( .A(n10667), .B(n2743), .Z(n7117) );
  OR U4849 ( .A(n2744), .B(n7117), .Z(n2745) );
  NANDN U4850 ( .A(n10670), .B(n2745), .Z(n2746) );
  NANDN U4851 ( .A(y[379]), .B(x[379]), .Z(n10031) );
  NAND U4852 ( .A(n2746), .B(n10031), .Z(n2749) );
  NANDN U4853 ( .A(x[380]), .B(y[380]), .Z(n2748) );
  ANDN U4854 ( .B(n2748), .A(n2747), .Z(n10673) );
  NAND U4855 ( .A(n2749), .B(n10673), .Z(n2750) );
  NANDN U4856 ( .A(n7122), .B(n2750), .Z(n2759) );
  NANDN U4857 ( .A(x[385]), .B(y[385]), .Z(n2752) );
  NANDN U4858 ( .A(x[384]), .B(y[384]), .Z(n2751) );
  AND U4859 ( .A(n2752), .B(n2751), .Z(n2758) );
  NANDN U4860 ( .A(x[382]), .B(y[382]), .Z(n2753) );
  NANDN U4861 ( .A(y[383]), .B(n2753), .Z(n2756) );
  XNOR U4862 ( .A(n2753), .B(y[383]), .Z(n2754) );
  NAND U4863 ( .A(n2754), .B(x[383]), .Z(n2755) );
  NAND U4864 ( .A(n2756), .B(n2755), .Z(n2757) );
  NAND U4865 ( .A(n2758), .B(n2757), .Z(n10678) );
  ANDN U4866 ( .B(n2759), .A(n10678), .Z(n2764) );
  NANDN U4867 ( .A(y[384]), .B(x[384]), .Z(n2760) );
  NANDN U4868 ( .A(n2760), .B(x[385]), .Z(n2763) );
  XNOR U4869 ( .A(n2760), .B(x[385]), .Z(n2761) );
  NANDN U4870 ( .A(y[385]), .B(n2761), .Z(n2762) );
  AND U4871 ( .A(n2763), .B(n2762), .Z(n10680) );
  NANDN U4872 ( .A(n2764), .B(n10680), .Z(n2765) );
  NANDN U4873 ( .A(x[387]), .B(y[387]), .Z(n2766) );
  NAND U4874 ( .A(n2765), .B(n10683), .Z(n2768) );
  NANDN U4875 ( .A(y[386]), .B(x[386]), .Z(n10681) );
  ANDN U4876 ( .B(x[387]), .A(y[387]), .Z(n10685) );
  ANDN U4877 ( .B(n10681), .A(n10685), .Z(n2767) );
  NANDN U4878 ( .A(n2767), .B(n2766), .Z(n7126) );
  NAND U4879 ( .A(n2768), .B(n7126), .Z(n2771) );
  NANDN U4880 ( .A(x[388]), .B(y[388]), .Z(n2770) );
  ANDN U4881 ( .B(n2770), .A(n2769), .Z(n10689) );
  NAND U4882 ( .A(n2771), .B(n10689), .Z(n2772) );
  NANDN U4883 ( .A(n7130), .B(n2772), .Z(n2777) );
  XNOR U4884 ( .A(y[391]), .B(x[391]), .Z(n2774) );
  NANDN U4885 ( .A(x[390]), .B(y[390]), .Z(n2773) );
  NAND U4886 ( .A(n2774), .B(n2773), .Z(n2775) );
  AND U4887 ( .A(n2776), .B(n2775), .Z(n10694) );
  ANDN U4888 ( .B(n2777), .A(n10694), .Z(n2778) );
  NANDN U4889 ( .A(x[392]), .B(y[392]), .Z(n6552) );
  NAND U4890 ( .A(n2778), .B(n6552), .Z(n2779) );
  NANDN U4891 ( .A(n10696), .B(n2779), .Z(n2780) );
  ANDN U4892 ( .B(y[393]), .A(x[393]), .Z(n6551) );
  ANDN U4893 ( .B(n2780), .A(n6551), .Z(n2781) );
  NANDN U4894 ( .A(y[394]), .B(x[394]), .Z(n10699) );
  NANDN U4895 ( .A(n2781), .B(n10699), .Z(n2782) );
  NANDN U4896 ( .A(n10702), .B(n2782), .Z(n2783) );
  NANDN U4897 ( .A(y[395]), .B(x[395]), .Z(n6549) );
  NAND U4898 ( .A(n2783), .B(n6549), .Z(n2784) );
  NAND U4899 ( .A(n6544), .B(n2784), .Z(n2785) );
  NANDN U4900 ( .A(n6550), .B(n2785), .Z(n2786) );
  ANDN U4901 ( .B(y[397]), .A(x[397]), .Z(n6543) );
  ANDN U4902 ( .B(n2786), .A(n6543), .Z(n2787) );
  NANDN U4903 ( .A(y[398]), .B(x[398]), .Z(n6540) );
  NANDN U4904 ( .A(n2787), .B(n6540), .Z(n2788) );
  NANDN U4905 ( .A(n6548), .B(n2788), .Z(n2793) );
  NANDN U4906 ( .A(y[400]), .B(x[400]), .Z(n2790) );
  NANDN U4907 ( .A(y[399]), .B(x[399]), .Z(n2789) );
  AND U4908 ( .A(n2790), .B(n2789), .Z(n2792) );
  NANDN U4909 ( .A(y[401]), .B(x[401]), .Z(n2791) );
  AND U4910 ( .A(n2792), .B(n2791), .Z(n6541) );
  NAND U4911 ( .A(n2793), .B(n6541), .Z(n2794) );
  NANDN U4912 ( .A(n10709), .B(n2794), .Z(n2799) );
  NANDN U4913 ( .A(y[402]), .B(x[402]), .Z(n2795) );
  NANDN U4914 ( .A(n2795), .B(x[403]), .Z(n2798) );
  XNOR U4915 ( .A(n2795), .B(x[403]), .Z(n2796) );
  NANDN U4916 ( .A(y[403]), .B(n2796), .Z(n2797) );
  AND U4917 ( .A(n2798), .B(n2797), .Z(n10712) );
  NAND U4918 ( .A(n2799), .B(n10712), .Z(n2800) );
  AND U4919 ( .A(n10716), .B(n2800), .Z(n2807) );
  NANDN U4920 ( .A(y[406]), .B(x[406]), .Z(n2802) );
  NANDN U4921 ( .A(y[405]), .B(x[405]), .Z(n2801) );
  AND U4922 ( .A(n2802), .B(n2801), .Z(n2804) );
  NANDN U4923 ( .A(y[407]), .B(x[407]), .Z(n2803) );
  NAND U4924 ( .A(n2804), .B(n2803), .Z(n10717) );
  ANDN U4925 ( .B(x[404]), .A(y[404]), .Z(n10711) );
  NANDN U4926 ( .A(n2805), .B(n10711), .Z(n2806) );
  NANDN U4927 ( .A(n10717), .B(n2806), .Z(n7143) );
  OR U4928 ( .A(n2807), .B(n7143), .Z(n2808) );
  NANDN U4929 ( .A(n10720), .B(n2808), .Z(n2813) );
  NANDN U4930 ( .A(y[408]), .B(x[408]), .Z(n2809) );
  NANDN U4931 ( .A(n2809), .B(x[409]), .Z(n2812) );
  XNOR U4932 ( .A(n2809), .B(x[409]), .Z(n2810) );
  NANDN U4933 ( .A(y[409]), .B(n2810), .Z(n2811) );
  AND U4934 ( .A(n2812), .B(n2811), .Z(n10722) );
  NAND U4935 ( .A(n2813), .B(n10722), .Z(n2815) );
  NAND U4936 ( .A(n2815), .B(n10725), .Z(n2816) );
  NANDN U4937 ( .A(n7148), .B(n2816), .Z(n2817) );
  AND U4938 ( .A(n10731), .B(n2817), .Z(n2822) );
  NANDN U4939 ( .A(y[414]), .B(x[414]), .Z(n2819) );
  NANDN U4940 ( .A(y[413]), .B(x[413]), .Z(n2818) );
  NAND U4941 ( .A(n2819), .B(n2818), .Z(n10733) );
  ANDN U4942 ( .B(x[412]), .A(y[412]), .Z(n10730) );
  NANDN U4943 ( .A(n2820), .B(n10730), .Z(n2821) );
  NANDN U4944 ( .A(n10733), .B(n2821), .Z(n7151) );
  OR U4945 ( .A(n2822), .B(n7151), .Z(n2825) );
  NANDN U4946 ( .A(x[414]), .B(y[414]), .Z(n2824) );
  NANDN U4947 ( .A(x[415]), .B(y[415]), .Z(n2823) );
  AND U4948 ( .A(n2824), .B(n2823), .Z(n10735) );
  NAND U4949 ( .A(n2825), .B(n10735), .Z(n2826) );
  NANDN U4950 ( .A(y[415]), .B(x[415]), .Z(n7153) );
  NAND U4951 ( .A(n2826), .B(n7153), .Z(n2827) );
  NAND U4952 ( .A(n6536), .B(n2827), .Z(n2828) );
  NANDN U4953 ( .A(n7154), .B(n2828), .Z(n2829) );
  ANDN U4954 ( .B(y[417]), .A(x[417]), .Z(n6535) );
  ANDN U4955 ( .B(n2829), .A(n6535), .Z(n2830) );
  NANDN U4956 ( .A(y[418]), .B(x[418]), .Z(n10741) );
  NANDN U4957 ( .A(n2830), .B(n10741), .Z(n2833) );
  NANDN U4958 ( .A(x[418]), .B(y[418]), .Z(n2832) );
  NANDN U4959 ( .A(x[419]), .B(y[419]), .Z(n2831) );
  AND U4960 ( .A(n2832), .B(n2831), .Z(n10743) );
  NAND U4961 ( .A(n2833), .B(n10743), .Z(n2834) );
  NANDN U4962 ( .A(n10744), .B(n2834), .Z(n2837) );
  NANDN U4963 ( .A(x[420]), .B(y[420]), .Z(n2836) );
  NANDN U4964 ( .A(x[421]), .B(y[421]), .Z(n2835) );
  AND U4965 ( .A(n2836), .B(n2835), .Z(n10745) );
  NAND U4966 ( .A(n2837), .B(n10745), .Z(n2838) );
  NANDN U4967 ( .A(n10746), .B(n2838), .Z(n2839) );
  AND U4968 ( .A(n10747), .B(n2839), .Z(n2840) );
  OR U4969 ( .A(n10748), .B(n2840), .Z(n2843) );
  NANDN U4970 ( .A(x[424]), .B(y[424]), .Z(n2842) );
  NANDN U4971 ( .A(x[425]), .B(y[425]), .Z(n2841) );
  AND U4972 ( .A(n2842), .B(n2841), .Z(n10749) );
  NAND U4973 ( .A(n2843), .B(n10749), .Z(n2845) );
  NANDN U4974 ( .A(y[426]), .B(x[426]), .Z(n2844) );
  ANDN U4975 ( .B(x[425]), .A(y[425]), .Z(n7166) );
  ANDN U4976 ( .B(n2844), .A(n7166), .Z(n10750) );
  NAND U4977 ( .A(n2845), .B(n10750), .Z(n2847) );
  NANDN U4978 ( .A(x[426]), .B(y[426]), .Z(n2846) );
  ANDN U4979 ( .B(y[427]), .A(x[427]), .Z(n7174) );
  ANDN U4980 ( .B(n2846), .A(n7174), .Z(n10751) );
  NAND U4981 ( .A(n2847), .B(n10751), .Z(n2848) );
  NANDN U4982 ( .A(y[427]), .B(x[427]), .Z(n10029) );
  NAND U4983 ( .A(n2848), .B(n10029), .Z(n2849) );
  AND U4984 ( .A(n10752), .B(n2849), .Z(n2855) );
  NANDN U4985 ( .A(y[428]), .B(x[428]), .Z(n10028) );
  NANDN U4986 ( .A(n10028), .B(n2850), .Z(n2851) );
  ANDN U4987 ( .B(n2851), .A(n10026), .Z(n2854) );
  NANDN U4988 ( .A(y[430]), .B(x[430]), .Z(n2853) );
  NANDN U4989 ( .A(y[429]), .B(x[429]), .Z(n2852) );
  NAND U4990 ( .A(n2853), .B(n2852), .Z(n10753) );
  ANDN U4991 ( .B(n2854), .A(n10753), .Z(n7175) );
  NANDN U4992 ( .A(n2855), .B(n7175), .Z(n2856) );
  AND U4993 ( .A(n7178), .B(n2856), .Z(n2857) );
  NANDN U4994 ( .A(x[432]), .B(y[432]), .Z(n10025) );
  NAND U4995 ( .A(n2857), .B(n10025), .Z(n2858) );
  NANDN U4996 ( .A(y[432]), .B(x[432]), .Z(n10027) );
  NAND U4997 ( .A(n2858), .B(n10027), .Z(n2859) );
  AND U4998 ( .A(n10024), .B(n2859), .Z(n2861) );
  IV U4999 ( .A(x[434]), .Z(n6534) );
  IV U5000 ( .A(y[434]), .Z(n6533) );
  NANDN U5001 ( .A(n6534), .B(n6533), .Z(n2860) );
  NANDN U5002 ( .A(y[433]), .B(x[433]), .Z(n7181) );
  NAND U5003 ( .A(n2860), .B(n7181), .Z(n10756) );
  OR U5004 ( .A(n2861), .B(n10756), .Z(n2862) );
  NANDN U5005 ( .A(n10758), .B(n2862), .Z(n2863) );
  NANDN U5006 ( .A(y[435]), .B(x[435]), .Z(n10761) );
  NAND U5007 ( .A(n2863), .B(n10761), .Z(n2866) );
  NANDN U5008 ( .A(x[436]), .B(y[436]), .Z(n2865) );
  ANDN U5009 ( .B(n2865), .A(n2864), .Z(n10763) );
  NAND U5010 ( .A(n2866), .B(n10763), .Z(n2867) );
  NANDN U5011 ( .A(n7192), .B(n2867), .Z(n2868) );
  AND U5012 ( .A(n10769), .B(n2868), .Z(n2873) );
  NANDN U5013 ( .A(y[440]), .B(x[440]), .Z(n2870) );
  NANDN U5014 ( .A(y[439]), .B(x[439]), .Z(n2869) );
  NAND U5015 ( .A(n2870), .B(n2869), .Z(n10771) );
  ANDN U5016 ( .B(x[438]), .A(y[438]), .Z(n10766) );
  NANDN U5017 ( .A(n2871), .B(n10766), .Z(n2872) );
  NANDN U5018 ( .A(n10771), .B(n2872), .Z(n7195) );
  OR U5019 ( .A(n2873), .B(n7195), .Z(n2876) );
  NANDN U5020 ( .A(x[441]), .B(y[441]), .Z(n2875) );
  NANDN U5021 ( .A(x[440]), .B(y[440]), .Z(n2874) );
  NAND U5022 ( .A(n2875), .B(n2874), .Z(n10774) );
  ANDN U5023 ( .B(n2876), .A(n10774), .Z(n2881) );
  NANDN U5024 ( .A(y[442]), .B(x[442]), .Z(n2878) );
  NANDN U5025 ( .A(y[441]), .B(x[441]), .Z(n2877) );
  AND U5026 ( .A(n2878), .B(n2877), .Z(n2880) );
  NANDN U5027 ( .A(y[443]), .B(x[443]), .Z(n2879) );
  AND U5028 ( .A(n2880), .B(n2879), .Z(n10775) );
  NANDN U5029 ( .A(n2881), .B(n10775), .Z(n2882) );
  NANDN U5030 ( .A(n10778), .B(n2882), .Z(n2887) );
  NANDN U5031 ( .A(y[444]), .B(x[444]), .Z(n2883) );
  NANDN U5032 ( .A(n2883), .B(x[445]), .Z(n2886) );
  XNOR U5033 ( .A(n2883), .B(x[445]), .Z(n2884) );
  NANDN U5034 ( .A(y[445]), .B(n2884), .Z(n2885) );
  AND U5035 ( .A(n2886), .B(n2885), .Z(n10780) );
  NAND U5036 ( .A(n2887), .B(n10780), .Z(n2888) );
  NANDN U5037 ( .A(n10784), .B(n2888), .Z(n2889) );
  NANDN U5038 ( .A(n7202), .B(n2889), .Z(n2890) );
  NANDN U5039 ( .A(n10790), .B(n2890), .Z(n2891) );
  NANDN U5040 ( .A(n10791), .B(n2891), .Z(n2892) );
  NANDN U5041 ( .A(n10794), .B(n2892), .Z(n2893) );
  AND U5042 ( .A(n10796), .B(n2893), .Z(n2895) );
  OR U5043 ( .A(n2895), .B(n10800), .Z(n2896) );
  NANDN U5044 ( .A(n7209), .B(n2896), .Z(n2897) );
  NANDN U5045 ( .A(n10806), .B(n2897), .Z(n2898) );
  NANDN U5046 ( .A(n10807), .B(n2898), .Z(n2899) );
  NANDN U5047 ( .A(n10810), .B(n2899), .Z(n2902) );
  NANDN U5048 ( .A(y[464]), .B(x[464]), .Z(n2900) );
  NAND U5049 ( .A(n2901), .B(n2900), .Z(n10812) );
  ANDN U5050 ( .B(n2902), .A(n10812), .Z(n2903) );
  OR U5051 ( .A(n10814), .B(n2903), .Z(n2906) );
  NANDN U5052 ( .A(y[466]), .B(x[466]), .Z(n2905) );
  NANDN U5053 ( .A(y[467]), .B(x[467]), .Z(n2904) );
  AND U5054 ( .A(n2905), .B(n2904), .Z(n10815) );
  NAND U5055 ( .A(n2906), .B(n10815), .Z(n2907) );
  NANDN U5056 ( .A(n10818), .B(n2907), .Z(n2908) );
  NANDN U5057 ( .A(n10819), .B(n2908), .Z(n2909) );
  NANDN U5058 ( .A(n10822), .B(n2909), .Z(n2910) );
  NANDN U5059 ( .A(n10823), .B(n2910), .Z(n2911) );
  ANDN U5060 ( .B(n2911), .A(n10826), .Z(n2920) );
  NANDN U5061 ( .A(y[478]), .B(x[478]), .Z(n2912) );
  AND U5062 ( .A(n2913), .B(n2912), .Z(n2919) );
  NANDN U5063 ( .A(y[476]), .B(x[476]), .Z(n2914) );
  NANDN U5064 ( .A(x[477]), .B(n2914), .Z(n2917) );
  XNOR U5065 ( .A(n2914), .B(x[477]), .Z(n2915) );
  NAND U5066 ( .A(n2915), .B(y[477]), .Z(n2916) );
  NAND U5067 ( .A(n2917), .B(n2916), .Z(n2918) );
  AND U5068 ( .A(n2919), .B(n2918), .Z(n10827) );
  NANDN U5069 ( .A(n2920), .B(n10827), .Z(n2921) );
  NANDN U5070 ( .A(n7225), .B(n2921), .Z(n2922) );
  NANDN U5071 ( .A(n7227), .B(n2922), .Z(n2923) );
  NANDN U5072 ( .A(n10840), .B(n2923), .Z(n2928) );
  NANDN U5073 ( .A(y[486]), .B(x[486]), .Z(n2925) );
  NANDN U5074 ( .A(y[485]), .B(x[485]), .Z(n2924) );
  AND U5075 ( .A(n2925), .B(n2924), .Z(n2927) );
  NANDN U5076 ( .A(y[487]), .B(x[487]), .Z(n2926) );
  AND U5077 ( .A(n2927), .B(n2926), .Z(n10841) );
  NAND U5078 ( .A(n2928), .B(n10841), .Z(n2937) );
  NANDN U5079 ( .A(x[489]), .B(y[489]), .Z(n2930) );
  NANDN U5080 ( .A(x[488]), .B(y[488]), .Z(n2929) );
  AND U5081 ( .A(n2930), .B(n2929), .Z(n2936) );
  NANDN U5082 ( .A(x[486]), .B(y[486]), .Z(n2931) );
  NANDN U5083 ( .A(y[487]), .B(n2931), .Z(n2934) );
  XNOR U5084 ( .A(n2931), .B(y[487]), .Z(n2932) );
  NAND U5085 ( .A(n2932), .B(x[487]), .Z(n2933) );
  NAND U5086 ( .A(n2934), .B(n2933), .Z(n2935) );
  NAND U5087 ( .A(n2936), .B(n2935), .Z(n10844) );
  ANDN U5088 ( .B(n2937), .A(n10844), .Z(n2938) );
  NANDN U5089 ( .A(n2938), .B(n10847), .Z(n2941) );
  NANDN U5090 ( .A(x[490]), .B(y[490]), .Z(n2940) );
  ANDN U5091 ( .B(n2940), .A(n2939), .Z(n10849) );
  NAND U5092 ( .A(n2941), .B(n10849), .Z(n2942) );
  NANDN U5093 ( .A(n7234), .B(n2942), .Z(n2943) );
  NANDN U5094 ( .A(n10853), .B(n2943), .Z(n2944) );
  NANDN U5095 ( .A(n10856), .B(n2944), .Z(n2953) );
  NANDN U5096 ( .A(x[499]), .B(y[499]), .Z(n2946) );
  NANDN U5097 ( .A(x[498]), .B(y[498]), .Z(n2945) );
  AND U5098 ( .A(n2946), .B(n2945), .Z(n2952) );
  NANDN U5099 ( .A(x[496]), .B(y[496]), .Z(n2947) );
  NANDN U5100 ( .A(y[497]), .B(n2947), .Z(n2950) );
  XNOR U5101 ( .A(n2947), .B(y[497]), .Z(n2948) );
  NAND U5102 ( .A(n2948), .B(x[497]), .Z(n2949) );
  NAND U5103 ( .A(n2950), .B(n2949), .Z(n2951) );
  NAND U5104 ( .A(n2952), .B(n2951), .Z(n10858) );
  ANDN U5105 ( .B(n2953), .A(n10858), .Z(n2954) );
  NANDN U5106 ( .A(n2954), .B(n10861), .Z(n2957) );
  NANDN U5107 ( .A(x[500]), .B(y[500]), .Z(n2956) );
  ANDN U5108 ( .B(n2956), .A(n2955), .Z(n10864) );
  NAND U5109 ( .A(n2957), .B(n10864), .Z(n2958) );
  NANDN U5110 ( .A(n7241), .B(n2958), .Z(n2959) );
  NANDN U5111 ( .A(n10869), .B(n2959), .Z(n2962) );
  NANDN U5112 ( .A(y[503]), .B(x[503]), .Z(n2961) );
  NANDN U5113 ( .A(y[504]), .B(x[504]), .Z(n2960) );
  AND U5114 ( .A(n2961), .B(n2960), .Z(n10871) );
  NAND U5115 ( .A(n2962), .B(n10871), .Z(n2965) );
  NANDN U5116 ( .A(x[505]), .B(y[505]), .Z(n2964) );
  NANDN U5117 ( .A(x[504]), .B(y[504]), .Z(n2963) );
  NAND U5118 ( .A(n2964), .B(n2963), .Z(n10874) );
  ANDN U5119 ( .B(n2965), .A(n10874), .Z(n2966) );
  NANDN U5120 ( .A(y[505]), .B(x[505]), .Z(n10875) );
  NANDN U5121 ( .A(n2966), .B(n10875), .Z(n2967) );
  NANDN U5122 ( .A(n10880), .B(n2967), .Z(n2968) );
  NANDN U5123 ( .A(n7248), .B(n2968), .Z(n2969) );
  NANDN U5124 ( .A(n10886), .B(n2969), .Z(n2972) );
  NANDN U5125 ( .A(y[511]), .B(x[511]), .Z(n2971) );
  NANDN U5126 ( .A(y[510]), .B(x[510]), .Z(n2970) );
  AND U5127 ( .A(n2971), .B(n2970), .Z(n10887) );
  NAND U5128 ( .A(n2972), .B(n10887), .Z(n2973) );
  AND U5129 ( .A(n6529), .B(n2973), .Z(n2974) );
  NANDN U5130 ( .A(x[511]), .B(y[511]), .Z(n10889) );
  NAND U5131 ( .A(n2974), .B(n10889), .Z(n2975) );
  AND U5132 ( .A(n2976), .B(n2975), .Z(n2977) );
  ANDN U5133 ( .B(n6530), .A(n2977), .Z(n2978) );
  NANDN U5134 ( .A(n10899), .B(n2978), .Z(n2981) );
  NANDN U5135 ( .A(y[515]), .B(x[515]), .Z(n10902) );
  ANDN U5136 ( .B(x[514]), .A(y[514]), .Z(n10895) );
  NAND U5137 ( .A(n2979), .B(n10895), .Z(n2980) );
  NAND U5138 ( .A(n10902), .B(n2980), .Z(n7257) );
  ANDN U5139 ( .B(n2981), .A(n7257), .Z(n2984) );
  NANDN U5140 ( .A(x[516]), .B(y[516]), .Z(n2983) );
  ANDN U5141 ( .B(n2983), .A(n2982), .Z(n10906) );
  NANDN U5142 ( .A(n2984), .B(n10906), .Z(n2985) );
  NANDN U5143 ( .A(n7260), .B(n2985), .Z(n2988) );
  NANDN U5144 ( .A(x[518]), .B(y[518]), .Z(n2987) );
  NANDN U5145 ( .A(x[519]), .B(y[519]), .Z(n2986) );
  AND U5146 ( .A(n2987), .B(n2986), .Z(n10909) );
  NAND U5147 ( .A(n2988), .B(n10909), .Z(n2989) );
  NANDN U5148 ( .A(n10912), .B(n2989), .Z(n2992) );
  NANDN U5149 ( .A(x[520]), .B(y[520]), .Z(n2991) );
  NANDN U5150 ( .A(x[521]), .B(y[521]), .Z(n2990) );
  AND U5151 ( .A(n2991), .B(n2990), .Z(n10913) );
  NAND U5152 ( .A(n2992), .B(n10913), .Z(n2993) );
  AND U5153 ( .A(n10915), .B(n2993), .Z(n2994) );
  ANDN U5154 ( .B(n10918), .A(n2994), .Z(n2995) );
  NANDN U5155 ( .A(x[524]), .B(y[524]), .Z(n6525) );
  NAND U5156 ( .A(n2995), .B(n6525), .Z(n2997) );
  ANDN U5157 ( .B(x[525]), .A(y[525]), .Z(n6526) );
  NANDN U5158 ( .A(y[524]), .B(x[524]), .Z(n2996) );
  NANDN U5159 ( .A(n6526), .B(n2996), .Z(n10920) );
  ANDN U5160 ( .B(n2997), .A(n10920), .Z(n3002) );
  NANDN U5161 ( .A(x[526]), .B(y[526]), .Z(n2999) );
  NANDN U5162 ( .A(x[525]), .B(y[525]), .Z(n2998) );
  AND U5163 ( .A(n2999), .B(n2998), .Z(n3001) );
  NANDN U5164 ( .A(x[527]), .B(y[527]), .Z(n3000) );
  AND U5165 ( .A(n3001), .B(n3000), .Z(n6527) );
  NANDN U5166 ( .A(n3002), .B(n6527), .Z(n3003) );
  ANDN U5167 ( .B(n3003), .A(n10924), .Z(n3012) );
  NANDN U5168 ( .A(x[531]), .B(y[531]), .Z(n3005) );
  NANDN U5169 ( .A(x[530]), .B(y[530]), .Z(n3004) );
  AND U5170 ( .A(n3005), .B(n3004), .Z(n3011) );
  NANDN U5171 ( .A(x[528]), .B(y[528]), .Z(n3006) );
  NANDN U5172 ( .A(y[529]), .B(n3006), .Z(n3009) );
  XNOR U5173 ( .A(n3006), .B(y[529]), .Z(n3007) );
  NAND U5174 ( .A(n3007), .B(x[529]), .Z(n3008) );
  NAND U5175 ( .A(n3009), .B(n3008), .Z(n3010) );
  NAND U5176 ( .A(n3011), .B(n3010), .Z(n10926) );
  OR U5177 ( .A(n3012), .B(n10926), .Z(n3013) );
  NAND U5178 ( .A(n3013), .B(n10927), .Z(n3014) );
  NANDN U5179 ( .A(n10932), .B(n3014), .Z(n3015) );
  NANDN U5180 ( .A(n7279), .B(n3015), .Z(n3016) );
  NANDN U5181 ( .A(n10938), .B(n3016), .Z(n3017) );
  AND U5182 ( .A(n10939), .B(n3017), .Z(n3018) );
  OR U5183 ( .A(n10942), .B(n3018), .Z(n3022) );
  NANDN U5184 ( .A(y[538]), .B(x[538]), .Z(n3020) );
  NANDN U5185 ( .A(y[537]), .B(x[537]), .Z(n3019) );
  AND U5186 ( .A(n3020), .B(n3019), .Z(n3021) );
  NANDN U5187 ( .A(y[539]), .B(x[539]), .Z(n3026) );
  AND U5188 ( .A(n3021), .B(n3026), .Z(n10943) );
  NAND U5189 ( .A(n3022), .B(n10943), .Z(n3029) );
  XNOR U5190 ( .A(y[539]), .B(x[539]), .Z(n3024) );
  NANDN U5191 ( .A(x[538]), .B(y[538]), .Z(n3023) );
  NAND U5192 ( .A(n3024), .B(n3023), .Z(n3025) );
  NAND U5193 ( .A(n3026), .B(n3025), .Z(n3028) );
  NANDN U5194 ( .A(x[540]), .B(y[540]), .Z(n3027) );
  NAND U5195 ( .A(n3028), .B(n3027), .Z(n7284) );
  NOR U5196 ( .A(n6523), .B(n7284), .Z(n10945) );
  NAND U5197 ( .A(n3029), .B(n10945), .Z(n3030) );
  NANDN U5198 ( .A(n10948), .B(n3030), .Z(n3036) );
  NANDN U5199 ( .A(x[545]), .B(y[545]), .Z(n7297) );
  ANDN U5200 ( .B(y[542]), .A(x[542]), .Z(n6524) );
  NAND U5201 ( .A(n3031), .B(n6524), .Z(n3032) );
  AND U5202 ( .A(n7297), .B(n3032), .Z(n3035) );
  NANDN U5203 ( .A(x[543]), .B(y[543]), .Z(n3034) );
  NANDN U5204 ( .A(x[544]), .B(y[544]), .Z(n3033) );
  NAND U5205 ( .A(n3034), .B(n3033), .Z(n7293) );
  ANDN U5206 ( .B(n3035), .A(n7293), .Z(n10949) );
  NAND U5207 ( .A(n3036), .B(n10949), .Z(n3042) );
  NANDN U5208 ( .A(y[546]), .B(x[546]), .Z(n3037) );
  NAND U5209 ( .A(n3038), .B(n3037), .Z(n7300) );
  NANDN U5210 ( .A(y[544]), .B(x[544]), .Z(n3040) );
  NANDN U5211 ( .A(y[545]), .B(x[545]), .Z(n3039) );
  NAND U5212 ( .A(n3040), .B(n3039), .Z(n7294) );
  NAND U5213 ( .A(n7294), .B(n7297), .Z(n3041) );
  NANDN U5214 ( .A(n7300), .B(n3041), .Z(n10951) );
  ANDN U5215 ( .B(n3042), .A(n10951), .Z(n3043) );
  OR U5216 ( .A(n10953), .B(n3043), .Z(n3044) );
  AND U5217 ( .A(n10954), .B(n3044), .Z(n3045) );
  OR U5218 ( .A(n10955), .B(n3045), .Z(n3046) );
  NANDN U5219 ( .A(y[549]), .B(x[549]), .Z(n10023) );
  NAND U5220 ( .A(n3046), .B(n10023), .Z(n3047) );
  NANDN U5221 ( .A(n10020), .B(n3047), .Z(n3048) );
  NANDN U5222 ( .A(n7309), .B(n3048), .Z(n3049) );
  NANDN U5223 ( .A(n10957), .B(n3049), .Z(n3050) );
  AND U5224 ( .A(n10959), .B(n3050), .Z(n3053) );
  NANDN U5225 ( .A(x[554]), .B(y[554]), .Z(n3052) );
  ANDN U5226 ( .B(n3052), .A(n3051), .Z(n10960) );
  NANDN U5227 ( .A(n3053), .B(n10960), .Z(n3054) );
  NANDN U5228 ( .A(n7314), .B(n3054), .Z(n3063) );
  NANDN U5229 ( .A(x[559]), .B(y[559]), .Z(n3056) );
  NANDN U5230 ( .A(x[558]), .B(y[558]), .Z(n3055) );
  AND U5231 ( .A(n3056), .B(n3055), .Z(n3062) );
  NANDN U5232 ( .A(x[556]), .B(y[556]), .Z(n3057) );
  NANDN U5233 ( .A(y[557]), .B(n3057), .Z(n3060) );
  XNOR U5234 ( .A(n3057), .B(y[557]), .Z(n3058) );
  NAND U5235 ( .A(n3058), .B(x[557]), .Z(n3059) );
  NAND U5236 ( .A(n3060), .B(n3059), .Z(n3061) );
  AND U5237 ( .A(n3062), .B(n3061), .Z(n10962) );
  NAND U5238 ( .A(n3063), .B(n10962), .Z(n3064) );
  NANDN U5239 ( .A(n10963), .B(n3064), .Z(n3074) );
  NANDN U5240 ( .A(x[563]), .B(y[563]), .Z(n3066) );
  NANDN U5241 ( .A(x[562]), .B(y[562]), .Z(n3065) );
  AND U5242 ( .A(n3066), .B(n3065), .Z(n3073) );
  NANDN U5243 ( .A(x[560]), .B(y[560]), .Z(n3068) );
  NANDN U5244 ( .A(y[561]), .B(n3068), .Z(n3071) );
  IV U5245 ( .A(y[561]), .Z(n3067) );
  XOR U5246 ( .A(n3068), .B(n3067), .Z(n3069) );
  NAND U5247 ( .A(n3069), .B(x[561]), .Z(n3070) );
  NAND U5248 ( .A(n3071), .B(n3070), .Z(n3072) );
  AND U5249 ( .A(n3073), .B(n3072), .Z(n10964) );
  NAND U5250 ( .A(n3074), .B(n10964), .Z(n3075) );
  ANDN U5251 ( .B(n3075), .A(n10965), .Z(n3076) );
  NANDN U5252 ( .A(n3076), .B(n10966), .Z(n3079) );
  NANDN U5253 ( .A(y[566]), .B(x[566]), .Z(n3078) );
  AND U5254 ( .A(n3078), .B(n3077), .Z(n10967) );
  NAND U5255 ( .A(n3079), .B(n10967), .Z(n3080) );
  NANDN U5256 ( .A(n10970), .B(n3080), .Z(n3081) );
  NANDN U5257 ( .A(n10972), .B(n3081), .Z(n3083) );
  NANDN U5258 ( .A(x[570]), .B(y[570]), .Z(n3082) );
  ANDN U5259 ( .B(y[571]), .A(x[571]), .Z(n7334) );
  ANDN U5260 ( .B(n3082), .A(n7334), .Z(n10974) );
  NAND U5261 ( .A(n3083), .B(n10974), .Z(n3084) );
  AND U5262 ( .A(n10976), .B(n3084), .Z(n3087) );
  NANDN U5263 ( .A(x[572]), .B(y[572]), .Z(n3086) );
  ANDN U5264 ( .B(n3086), .A(n3085), .Z(n10980) );
  NANDN U5265 ( .A(n3087), .B(n10980), .Z(n3088) );
  NANDN U5266 ( .A(n7336), .B(n3088), .Z(n3089) );
  NANDN U5267 ( .A(n10983), .B(n3089), .Z(n3096) );
  NANDN U5268 ( .A(y[577]), .B(x[577]), .Z(n3091) );
  ANDN U5269 ( .B(x[578]), .A(y[578]), .Z(n3090) );
  ANDN U5270 ( .B(n3091), .A(n3090), .Z(n3095) );
  XNOR U5271 ( .A(x[577]), .B(y[577]), .Z(n3093) );
  ANDN U5272 ( .B(x[576]), .A(y[576]), .Z(n3092) );
  NAND U5273 ( .A(n3093), .B(n3092), .Z(n3094) );
  AND U5274 ( .A(n3095), .B(n3094), .Z(n10985) );
  NAND U5275 ( .A(n3096), .B(n10985), .Z(n3097) );
  NANDN U5276 ( .A(n10988), .B(n3097), .Z(n3098) );
  AND U5277 ( .A(n10989), .B(n3098), .Z(n3100) );
  NANDN U5278 ( .A(n3100), .B(n10993), .Z(n3101) );
  NANDN U5279 ( .A(n7342), .B(n3101), .Z(n3102) );
  NANDN U5280 ( .A(x[583]), .B(y[583]), .Z(n3104) );
  NAND U5281 ( .A(n3102), .B(n10999), .Z(n3105) );
  ANDN U5282 ( .B(x[582]), .A(y[582]), .Z(n10998) );
  ANDN U5283 ( .B(x[583]), .A(y[583]), .Z(n11004) );
  OR U5284 ( .A(n10998), .B(n11004), .Z(n3103) );
  NAND U5285 ( .A(n3104), .B(n3103), .Z(n7345) );
  NAND U5286 ( .A(n3105), .B(n7345), .Z(n3106) );
  NANDN U5287 ( .A(n10018), .B(n3106), .Z(n3112) );
  NANDN U5288 ( .A(y[587]), .B(x[587]), .Z(n3108) );
  NANDN U5289 ( .A(y[586]), .B(x[586]), .Z(n3107) );
  NAND U5290 ( .A(n3108), .B(n3107), .Z(n11007) );
  ANDN U5291 ( .B(x[585]), .A(y[585]), .Z(n10019) );
  NANDN U5292 ( .A(y[584]), .B(x[584]), .Z(n3109) );
  NANDN U5293 ( .A(n10019), .B(n3109), .Z(n11002) );
  NANDN U5294 ( .A(n3110), .B(n11002), .Z(n3111) );
  NANDN U5295 ( .A(n11007), .B(n3111), .Z(n7349) );
  ANDN U5296 ( .B(n3112), .A(n7349), .Z(n3119) );
  NANDN U5297 ( .A(x[587]), .B(y[587]), .Z(n3114) );
  ANDN U5298 ( .B(y[588]), .A(x[588]), .Z(n3113) );
  ANDN U5299 ( .B(n3114), .A(n3113), .Z(n3118) );
  XNOR U5300 ( .A(y[587]), .B(x[587]), .Z(n3116) );
  ANDN U5301 ( .B(y[586]), .A(x[586]), .Z(n3115) );
  NAND U5302 ( .A(n3116), .B(n3115), .Z(n3117) );
  AND U5303 ( .A(n3118), .B(n3117), .Z(n11010) );
  NANDN U5304 ( .A(n3119), .B(n11010), .Z(n3120) );
  NANDN U5305 ( .A(n11012), .B(n3120), .Z(n3121) );
  NANDN U5306 ( .A(x[590]), .B(y[590]), .Z(n11017) );
  ANDN U5307 ( .B(y[589]), .A(x[589]), .Z(n11014) );
  ANDN U5308 ( .B(n11017), .A(n11014), .Z(n7352) );
  NAND U5309 ( .A(n3121), .B(n7352), .Z(n3122) );
  NANDN U5310 ( .A(n11016), .B(n3122), .Z(n3125) );
  NANDN U5311 ( .A(x[591]), .B(y[591]), .Z(n3124) );
  ANDN U5312 ( .B(n3124), .A(n11026), .Z(n7355) );
  NAND U5313 ( .A(n3125), .B(n7355), .Z(n3126) );
  AND U5314 ( .A(n6522), .B(n3126), .Z(n3128) );
  NANDN U5315 ( .A(y[594]), .B(x[594]), .Z(n3127) );
  ANDN U5316 ( .B(x[593]), .A(y[593]), .Z(n6521) );
  ANDN U5317 ( .B(n3127), .A(n6521), .Z(n11027) );
  NAND U5318 ( .A(n3128), .B(n11027), .Z(n3129) );
  NANDN U5319 ( .A(n11030), .B(n3129), .Z(n3133) );
  NANDN U5320 ( .A(y[596]), .B(x[596]), .Z(n3130) );
  NANDN U5321 ( .A(n3131), .B(n3130), .Z(n7368) );
  NANDN U5322 ( .A(y[595]), .B(x[595]), .Z(n3132) );
  NANDN U5323 ( .A(n7368), .B(n3132), .Z(n11032) );
  ANDN U5324 ( .B(n3133), .A(n11032), .Z(n3134) );
  OR U5325 ( .A(n11033), .B(n3134), .Z(n3135) );
  NANDN U5326 ( .A(n11036), .B(n3135), .Z(n3144) );
  NANDN U5327 ( .A(x[603]), .B(y[603]), .Z(n3137) );
  NANDN U5328 ( .A(x[602]), .B(y[602]), .Z(n3136) );
  AND U5329 ( .A(n3137), .B(n3136), .Z(n3143) );
  NANDN U5330 ( .A(x[600]), .B(y[600]), .Z(n3138) );
  NANDN U5331 ( .A(y[601]), .B(n3138), .Z(n3141) );
  XNOR U5332 ( .A(n3138), .B(y[601]), .Z(n3139) );
  NAND U5333 ( .A(n3139), .B(x[601]), .Z(n3140) );
  NAND U5334 ( .A(n3141), .B(n3140), .Z(n3142) );
  AND U5335 ( .A(n3143), .B(n3142), .Z(n11037) );
  NAND U5336 ( .A(n3144), .B(n11037), .Z(n3145) );
  NANDN U5337 ( .A(n11040), .B(n3145), .Z(n3152) );
  NANDN U5338 ( .A(x[605]), .B(y[605]), .Z(n3147) );
  ANDN U5339 ( .B(y[606]), .A(x[606]), .Z(n3146) );
  ANDN U5340 ( .B(n3147), .A(n3146), .Z(n3151) );
  XNOR U5341 ( .A(y[605]), .B(x[605]), .Z(n3149) );
  ANDN U5342 ( .B(y[604]), .A(x[604]), .Z(n3148) );
  NAND U5343 ( .A(n3149), .B(n3148), .Z(n3150) );
  AND U5344 ( .A(n3151), .B(n3150), .Z(n11041) );
  NAND U5345 ( .A(n3152), .B(n11041), .Z(n3155) );
  NANDN U5346 ( .A(y[606]), .B(x[606]), .Z(n3154) );
  NANDN U5347 ( .A(y[607]), .B(x[607]), .Z(n3153) );
  NAND U5348 ( .A(n3154), .B(n3153), .Z(n11044) );
  ANDN U5349 ( .B(n3155), .A(n11044), .Z(n3156) );
  NANDN U5350 ( .A(x[607]), .B(y[607]), .Z(n11046) );
  NANDN U5351 ( .A(n3156), .B(n11046), .Z(n3157) );
  NANDN U5352 ( .A(n11048), .B(n3157), .Z(n3158) );
  AND U5353 ( .A(n3159), .B(n3158), .Z(n3166) );
  NANDN U5354 ( .A(y[612]), .B(x[612]), .Z(n3161) );
  NANDN U5355 ( .A(y[611]), .B(x[611]), .Z(n3160) );
  AND U5356 ( .A(n3161), .B(n3160), .Z(n3163) );
  NANDN U5357 ( .A(y[613]), .B(x[613]), .Z(n3162) );
  NAND U5358 ( .A(n3163), .B(n3162), .Z(n11056) );
  ANDN U5359 ( .B(x[610]), .A(y[610]), .Z(n11052) );
  NANDN U5360 ( .A(n3164), .B(n11052), .Z(n3165) );
  NANDN U5361 ( .A(n11056), .B(n3165), .Z(n7384) );
  OR U5362 ( .A(n3166), .B(n7384), .Z(n3171) );
  NANDN U5363 ( .A(x[612]), .B(y[612]), .Z(n3167) );
  NANDN U5364 ( .A(n3167), .B(y[613]), .Z(n3170) );
  XNOR U5365 ( .A(n3167), .B(y[613]), .Z(n3168) );
  NANDN U5366 ( .A(x[613]), .B(n3168), .Z(n3169) );
  AND U5367 ( .A(n3170), .B(n3169), .Z(n11058) );
  NAND U5368 ( .A(n3171), .B(n11058), .Z(n3172) );
  NANDN U5369 ( .A(n11060), .B(n3172), .Z(n3173) );
  NANDN U5370 ( .A(n11062), .B(n3173), .Z(n3174) );
  NANDN U5371 ( .A(n11064), .B(n3174), .Z(n3180) );
  NANDN U5372 ( .A(x[618]), .B(y[618]), .Z(n3176) );
  IV U5373 ( .A(y[619]), .Z(n3175) );
  OR U5374 ( .A(n3176), .B(n3175), .Z(n3179) );
  XNOR U5375 ( .A(n3176), .B(y[619]), .Z(n3177) );
  NANDN U5376 ( .A(x[619]), .B(n3177), .Z(n3178) );
  AND U5377 ( .A(n3179), .B(n3178), .Z(n11065) );
  NAND U5378 ( .A(n3180), .B(n11065), .Z(n3182) );
  ANDN U5379 ( .B(y[620]), .A(x[620]), .Z(n3181) );
  OR U5380 ( .A(n3182), .B(n3181), .Z(n3183) );
  NANDN U5381 ( .A(n11068), .B(n3183), .Z(n3184) );
  NANDN U5382 ( .A(x[621]), .B(y[621]), .Z(n6512) );
  NAND U5383 ( .A(n3184), .B(n6512), .Z(n3185) );
  OR U5384 ( .A(n6516), .B(n3185), .Z(n3186) );
  AND U5385 ( .A(n11071), .B(n3186), .Z(n3195) );
  NANDN U5386 ( .A(x[627]), .B(y[627]), .Z(n3188) );
  NANDN U5387 ( .A(x[626]), .B(y[626]), .Z(n3187) );
  AND U5388 ( .A(n3188), .B(n3187), .Z(n3194) );
  NANDN U5389 ( .A(x[624]), .B(y[624]), .Z(n3189) );
  NANDN U5390 ( .A(y[625]), .B(n3189), .Z(n3192) );
  XNOR U5391 ( .A(n3189), .B(y[625]), .Z(n3190) );
  NAND U5392 ( .A(n3190), .B(x[625]), .Z(n3191) );
  NAND U5393 ( .A(n3192), .B(n3191), .Z(n3193) );
  NAND U5394 ( .A(n3194), .B(n3193), .Z(n11074) );
  OR U5395 ( .A(n3195), .B(n11074), .Z(n3196) );
  NAND U5396 ( .A(n3196), .B(n11075), .Z(n3197) );
  NANDN U5397 ( .A(x[629]), .B(y[629]), .Z(n3201) );
  ANDN U5398 ( .B(n3197), .A(n11080), .Z(n3204) );
  NANDN U5399 ( .A(y[630]), .B(x[630]), .Z(n3199) );
  NAND U5400 ( .A(n3199), .B(n3198), .Z(n11082) );
  NANDN U5401 ( .A(y[628]), .B(x[628]), .Z(n3200) );
  ANDN U5402 ( .B(x[629]), .A(y[629]), .Z(n11081) );
  ANDN U5403 ( .B(n3200), .A(n11081), .Z(n3202) );
  NANDN U5404 ( .A(n3202), .B(n3201), .Z(n3203) );
  NANDN U5405 ( .A(n11082), .B(n3203), .Z(n7400) );
  OR U5406 ( .A(n3204), .B(n7400), .Z(n3205) );
  NANDN U5407 ( .A(n11083), .B(n3205), .Z(n3214) );
  ANDN U5408 ( .B(x[635]), .A(y[635]), .Z(n3211) );
  NANDN U5409 ( .A(y[633]), .B(x[633]), .Z(n3209) );
  AND U5410 ( .A(x[632]), .B(n3206), .Z(n3207) );
  NANDN U5411 ( .A(y[632]), .B(n3207), .Z(n3208) );
  NAND U5412 ( .A(n3209), .B(n3208), .Z(n3210) );
  NOR U5413 ( .A(n3211), .B(n3210), .Z(n3213) );
  NANDN U5414 ( .A(y[634]), .B(x[634]), .Z(n3212) );
  AND U5415 ( .A(n3213), .B(n3212), .Z(n11084) );
  NAND U5416 ( .A(n3214), .B(n11084), .Z(n3215) );
  NANDN U5417 ( .A(n11085), .B(n3215), .Z(n3216) );
  NANDN U5418 ( .A(n11086), .B(n3216), .Z(n3225) );
  NANDN U5419 ( .A(x[640]), .B(y[640]), .Z(n3217) );
  AND U5420 ( .A(n3218), .B(n3217), .Z(n3224) );
  NANDN U5421 ( .A(x[638]), .B(y[638]), .Z(n3219) );
  NANDN U5422 ( .A(y[639]), .B(n3219), .Z(n3222) );
  XNOR U5423 ( .A(n3219), .B(y[639]), .Z(n3220) );
  NAND U5424 ( .A(n3220), .B(x[639]), .Z(n3221) );
  NAND U5425 ( .A(n3222), .B(n3221), .Z(n3223) );
  NAND U5426 ( .A(n3224), .B(n3223), .Z(n11087) );
  ANDN U5427 ( .B(n3225), .A(n11087), .Z(n3226) );
  OR U5428 ( .A(n11088), .B(n3226), .Z(n3227) );
  NANDN U5429 ( .A(n11089), .B(n3227), .Z(n3228) );
  NANDN U5430 ( .A(y[643]), .B(x[643]), .Z(n11091) );
  NAND U5431 ( .A(n3228), .B(n11091), .Z(n3231) );
  NANDN U5432 ( .A(x[644]), .B(y[644]), .Z(n3230) );
  ANDN U5433 ( .B(n3230), .A(n3229), .Z(n11092) );
  NAND U5434 ( .A(n3231), .B(n11092), .Z(n3232) );
  NANDN U5435 ( .A(n7417), .B(n3232), .Z(n3233) );
  NANDN U5436 ( .A(n11094), .B(n3233), .Z(n3234) );
  NANDN U5437 ( .A(y[647]), .B(x[647]), .Z(n10017) );
  NAND U5438 ( .A(n3234), .B(n10017), .Z(n3235) );
  NANDN U5439 ( .A(n11095), .B(n3235), .Z(n3238) );
  ANDN U5440 ( .B(x[649]), .A(y[649]), .Z(n11098) );
  NANDN U5441 ( .A(y[648]), .B(x[648]), .Z(n10016) );
  NANDN U5442 ( .A(n10016), .B(n3236), .Z(n3237) );
  NANDN U5443 ( .A(n11098), .B(n3237), .Z(n7422) );
  ANDN U5444 ( .B(n3238), .A(n7422), .Z(n3241) );
  NANDN U5445 ( .A(x[650]), .B(y[650]), .Z(n3240) );
  ANDN U5446 ( .B(n3240), .A(n3239), .Z(n11099) );
  NANDN U5447 ( .A(n3241), .B(n11099), .Z(n3242) );
  NANDN U5448 ( .A(n7425), .B(n3242), .Z(n3243) );
  NANDN U5449 ( .A(n11101), .B(n3243), .Z(n3250) );
  NANDN U5450 ( .A(y[655]), .B(x[655]), .Z(n3245) );
  ANDN U5451 ( .B(x[656]), .A(y[656]), .Z(n3244) );
  ANDN U5452 ( .B(n3245), .A(n3244), .Z(n3249) );
  XNOR U5453 ( .A(x[655]), .B(y[655]), .Z(n3247) );
  ANDN U5454 ( .B(x[654]), .A(y[654]), .Z(n3246) );
  NAND U5455 ( .A(n3247), .B(n3246), .Z(n3248) );
  AND U5456 ( .A(n3249), .B(n3248), .Z(n11102) );
  NAND U5457 ( .A(n3250), .B(n11102), .Z(n3251) );
  NANDN U5458 ( .A(n11103), .B(n3251), .Z(n3252) );
  NANDN U5459 ( .A(y[657]), .B(x[657]), .Z(n11105) );
  NAND U5460 ( .A(n3252), .B(n11105), .Z(n3255) );
  NANDN U5461 ( .A(x[658]), .B(y[658]), .Z(n3254) );
  ANDN U5462 ( .B(n3254), .A(n3253), .Z(n11106) );
  NAND U5463 ( .A(n3255), .B(n11106), .Z(n3256) );
  NANDN U5464 ( .A(n7432), .B(n3256), .Z(n3257) );
  AND U5465 ( .A(n11109), .B(n3257), .Z(n3264) );
  NANDN U5466 ( .A(y[662]), .B(x[662]), .Z(n3259) );
  NANDN U5467 ( .A(y[661]), .B(x[661]), .Z(n3258) );
  AND U5468 ( .A(n3259), .B(n3258), .Z(n3261) );
  NANDN U5469 ( .A(y[663]), .B(x[663]), .Z(n3260) );
  NAND U5470 ( .A(n3261), .B(n3260), .Z(n11110) );
  ANDN U5471 ( .B(x[660]), .A(y[660]), .Z(n11107) );
  NANDN U5472 ( .A(n3262), .B(n11107), .Z(n3263) );
  NANDN U5473 ( .A(n11110), .B(n3263), .Z(n7434) );
  OR U5474 ( .A(n3264), .B(n7434), .Z(n3273) );
  NANDN U5475 ( .A(x[664]), .B(y[664]), .Z(n3265) );
  AND U5476 ( .A(n3266), .B(n3265), .Z(n3272) );
  NANDN U5477 ( .A(x[662]), .B(y[662]), .Z(n3267) );
  NANDN U5478 ( .A(y[663]), .B(n3267), .Z(n3270) );
  XNOR U5479 ( .A(n3267), .B(y[663]), .Z(n3268) );
  NAND U5480 ( .A(n3268), .B(x[663]), .Z(n3269) );
  NAND U5481 ( .A(n3270), .B(n3269), .Z(n3271) );
  AND U5482 ( .A(n3272), .B(n3271), .Z(n11111) );
  NAND U5483 ( .A(n3273), .B(n11111), .Z(n3274) );
  NANDN U5484 ( .A(n11112), .B(n3274), .Z(n3276) );
  NANDN U5485 ( .A(x[666]), .B(y[666]), .Z(n3275) );
  ANDN U5486 ( .B(y[667]), .A(x[667]), .Z(n3278) );
  ANDN U5487 ( .B(n3275), .A(n3278), .Z(n11114) );
  NAND U5488 ( .A(n3276), .B(n11114), .Z(n3279) );
  NANDN U5489 ( .A(y[666]), .B(x[666]), .Z(n11113) );
  ANDN U5490 ( .B(x[667]), .A(y[667]), .Z(n11115) );
  ANDN U5491 ( .B(n11113), .A(n11115), .Z(n3277) );
  OR U5492 ( .A(n3278), .B(n3277), .Z(n7439) );
  NAND U5493 ( .A(n3279), .B(n7439), .Z(n3280) );
  AND U5494 ( .A(n11116), .B(n3280), .Z(n3281) );
  ANDN U5495 ( .B(n11118), .A(n3281), .Z(n3282) );
  NANDN U5496 ( .A(n6509), .B(n3282), .Z(n3283) );
  NANDN U5497 ( .A(x[671]), .B(y[671]), .Z(n7450) );
  NANDN U5498 ( .A(x[670]), .B(y[670]), .Z(n7445) );
  NAND U5499 ( .A(n7450), .B(n7445), .Z(n11119) );
  ANDN U5500 ( .B(n3283), .A(n11119), .Z(n3284) );
  NANDN U5501 ( .A(y[671]), .B(x[671]), .Z(n11120) );
  NANDN U5502 ( .A(n3284), .B(n11120), .Z(n3285) );
  NANDN U5503 ( .A(x[673]), .B(y[673]), .Z(n3286) );
  NAND U5504 ( .A(n3285), .B(n11122), .Z(n3287) );
  ANDN U5505 ( .B(x[672]), .A(y[672]), .Z(n11121) );
  NAND U5506 ( .A(n3286), .B(n11121), .Z(n7455) );
  NAND U5507 ( .A(n3287), .B(n7455), .Z(n3289) );
  NANDN U5508 ( .A(y[673]), .B(x[673]), .Z(n7453) );
  NANDN U5509 ( .A(y[674]), .B(x[674]), .Z(n3288) );
  NAND U5510 ( .A(n7453), .B(n3288), .Z(n11123) );
  OR U5511 ( .A(n3289), .B(n11123), .Z(n3290) );
  NANDN U5512 ( .A(n11124), .B(n3290), .Z(n3293) );
  NANDN U5513 ( .A(y[675]), .B(x[675]), .Z(n3292) );
  NANDN U5514 ( .A(y[676]), .B(x[676]), .Z(n3291) );
  AND U5515 ( .A(n3292), .B(n3291), .Z(n11125) );
  NAND U5516 ( .A(n3293), .B(n11125), .Z(n3294) );
  NANDN U5517 ( .A(n11126), .B(n3294), .Z(n3295) );
  NANDN U5518 ( .A(y[677]), .B(x[677]), .Z(n11128) );
  NAND U5519 ( .A(n3295), .B(n11128), .Z(n3297) );
  NANDN U5520 ( .A(x[679]), .B(y[679]), .Z(n3301) );
  NANDN U5521 ( .A(x[678]), .B(y[678]), .Z(n3296) );
  NAND U5522 ( .A(n3301), .B(n3296), .Z(n11129) );
  ANDN U5523 ( .B(n3297), .A(n11129), .Z(n3303) );
  NANDN U5524 ( .A(y[680]), .B(x[680]), .Z(n3299) );
  NANDN U5525 ( .A(y[679]), .B(x[679]), .Z(n3298) );
  AND U5526 ( .A(n3299), .B(n3298), .Z(n3300) );
  NANDN U5527 ( .A(y[681]), .B(x[681]), .Z(n3309) );
  NAND U5528 ( .A(n3300), .B(n3309), .Z(n11130) );
  NANDN U5529 ( .A(y[678]), .B(x[678]), .Z(n11127) );
  NANDN U5530 ( .A(n11127), .B(n3301), .Z(n3302) );
  NANDN U5531 ( .A(n11130), .B(n3302), .Z(n7467) );
  OR U5532 ( .A(n3303), .B(n7467), .Z(n3310) );
  NANDN U5533 ( .A(x[682]), .B(y[682]), .Z(n3304) );
  NANDN U5534 ( .A(n3305), .B(n3304), .Z(n11133) );
  XNOR U5535 ( .A(y[681]), .B(x[681]), .Z(n3307) );
  NANDN U5536 ( .A(x[680]), .B(y[680]), .Z(n3306) );
  NAND U5537 ( .A(n3307), .B(n3306), .Z(n3308) );
  AND U5538 ( .A(n3309), .B(n3308), .Z(n11131) );
  NOR U5539 ( .A(n11133), .B(n11131), .Z(n7468) );
  NAND U5540 ( .A(n3310), .B(n7468), .Z(n3311) );
  NANDN U5541 ( .A(n7471), .B(n3311), .Z(n3312) );
  NAND U5542 ( .A(n3313), .B(n3312), .Z(n3319) );
  NANDN U5543 ( .A(y[688]), .B(x[688]), .Z(n3314) );
  AND U5544 ( .A(n3315), .B(n3314), .Z(n11139) );
  NANDN U5545 ( .A(y[687]), .B(x[687]), .Z(n7475) );
  OR U5546 ( .A(n11136), .B(n3316), .Z(n3317) );
  AND U5547 ( .A(n11139), .B(n3317), .Z(n3318) );
  NAND U5548 ( .A(n3319), .B(n3318), .Z(n3320) );
  NANDN U5549 ( .A(n11140), .B(n3320), .Z(n3327) );
  NANDN U5550 ( .A(y[691]), .B(x[691]), .Z(n3322) );
  ANDN U5551 ( .B(x[692]), .A(y[692]), .Z(n3321) );
  ANDN U5552 ( .B(n3322), .A(n3321), .Z(n3326) );
  XNOR U5553 ( .A(x[691]), .B(y[691]), .Z(n3324) );
  ANDN U5554 ( .B(x[690]), .A(y[690]), .Z(n3323) );
  NAND U5555 ( .A(n3324), .B(n3323), .Z(n3325) );
  AND U5556 ( .A(n3326), .B(n3325), .Z(n11141) );
  NAND U5557 ( .A(n3327), .B(n11141), .Z(n3330) );
  NANDN U5558 ( .A(x[693]), .B(y[693]), .Z(n3329) );
  NANDN U5559 ( .A(x[692]), .B(y[692]), .Z(n3328) );
  NAND U5560 ( .A(n3329), .B(n3328), .Z(n11142) );
  ANDN U5561 ( .B(n3330), .A(n11142), .Z(n3333) );
  NANDN U5562 ( .A(y[693]), .B(x[693]), .Z(n3332) );
  NANDN U5563 ( .A(y[694]), .B(x[694]), .Z(n3331) );
  AND U5564 ( .A(n3332), .B(n3331), .Z(n11143) );
  NANDN U5565 ( .A(n3333), .B(n11143), .Z(n3334) );
  NANDN U5566 ( .A(n11144), .B(n3334), .Z(n3335) );
  NANDN U5567 ( .A(y[695]), .B(x[695]), .Z(n11146) );
  NAND U5568 ( .A(n3335), .B(n11146), .Z(n3337) );
  NANDN U5569 ( .A(x[696]), .B(y[696]), .Z(n3336) );
  NANDN U5570 ( .A(x[697]), .B(y[697]), .Z(n3338) );
  AND U5571 ( .A(n3336), .B(n3338), .Z(n11147) );
  NAND U5572 ( .A(n3337), .B(n11147), .Z(n3343) );
  NANDN U5573 ( .A(y[696]), .B(x[696]), .Z(n11145) );
  NANDN U5574 ( .A(n11145), .B(n3338), .Z(n3339) );
  ANDN U5575 ( .B(x[699]), .A(y[699]), .Z(n10014) );
  ANDN U5576 ( .B(n3339), .A(n10014), .Z(n3342) );
  NANDN U5577 ( .A(y[698]), .B(x[698]), .Z(n3341) );
  NANDN U5578 ( .A(y[697]), .B(x[697]), .Z(n3340) );
  NAND U5579 ( .A(n3341), .B(n3340), .Z(n11148) );
  ANDN U5580 ( .B(n3342), .A(n11148), .Z(n7490) );
  NAND U5581 ( .A(n3343), .B(n7490), .Z(n3348) );
  NANDN U5582 ( .A(x[701]), .B(y[701]), .Z(n3351) );
  NANDN U5583 ( .A(x[700]), .B(y[700]), .Z(n3344) );
  NAND U5584 ( .A(n3351), .B(n3344), .Z(n11150) );
  NANDN U5585 ( .A(x[699]), .B(y[699]), .Z(n3346) );
  NANDN U5586 ( .A(x[698]), .B(y[698]), .Z(n3345) );
  NAND U5587 ( .A(n3346), .B(n3345), .Z(n11149) );
  NANDN U5588 ( .A(n10014), .B(n11149), .Z(n3347) );
  NANDN U5589 ( .A(n11150), .B(n3347), .Z(n7492) );
  ANDN U5590 ( .B(n3348), .A(n7492), .Z(n3353) );
  NANDN U5591 ( .A(y[702]), .B(x[702]), .Z(n3350) );
  NANDN U5592 ( .A(y[701]), .B(x[701]), .Z(n3349) );
  NAND U5593 ( .A(n3350), .B(n3349), .Z(n11151) );
  NANDN U5594 ( .A(y[700]), .B(x[700]), .Z(n10013) );
  NANDN U5595 ( .A(n10013), .B(n3351), .Z(n3352) );
  NANDN U5596 ( .A(n11151), .B(n3352), .Z(n7495) );
  OR U5597 ( .A(n3353), .B(n7495), .Z(n3354) );
  NANDN U5598 ( .A(n11152), .B(n3354), .Z(n3357) );
  NANDN U5599 ( .A(y[703]), .B(x[703]), .Z(n3356) );
  NANDN U5600 ( .A(y[704]), .B(x[704]), .Z(n3355) );
  AND U5601 ( .A(n3356), .B(n3355), .Z(n11153) );
  NAND U5602 ( .A(n3357), .B(n11153), .Z(n3358) );
  NANDN U5603 ( .A(n11156), .B(n3358), .Z(n3359) );
  NANDN U5604 ( .A(y[705]), .B(x[705]), .Z(n11159) );
  NAND U5605 ( .A(n3359), .B(n11159), .Z(n3360) );
  AND U5606 ( .A(n11161), .B(n3360), .Z(n3363) );
  ANDN U5607 ( .B(x[707]), .A(y[707]), .Z(n11166) );
  ANDN U5608 ( .B(x[706]), .A(y[706]), .Z(n11158) );
  NANDN U5609 ( .A(n3361), .B(n11158), .Z(n3362) );
  NANDN U5610 ( .A(n11166), .B(n3362), .Z(n7502) );
  OR U5611 ( .A(n3363), .B(n7502), .Z(n3365) );
  NANDN U5612 ( .A(x[708]), .B(y[708]), .Z(n3364) );
  ANDN U5613 ( .B(y[709]), .A(x[709]), .Z(n3366) );
  ANDN U5614 ( .B(n3364), .A(n3366), .Z(n11167) );
  NAND U5615 ( .A(n3365), .B(n11167), .Z(n3368) );
  ANDN U5616 ( .B(x[709]), .A(y[709]), .Z(n11170) );
  ANDN U5617 ( .B(x[708]), .A(y[708]), .Z(n11164) );
  NANDN U5618 ( .A(n3366), .B(n11164), .Z(n3367) );
  NANDN U5619 ( .A(n11170), .B(n3367), .Z(n7505) );
  ANDN U5620 ( .B(n3368), .A(n7505), .Z(n3369) );
  NANDN U5621 ( .A(y[710]), .B(x[710]), .Z(n11171) );
  NAND U5622 ( .A(n3369), .B(n11171), .Z(n3371) );
  NANDN U5623 ( .A(x[710]), .B(y[710]), .Z(n3370) );
  ANDN U5624 ( .B(y[711]), .A(x[711]), .Z(n6508) );
  ANDN U5625 ( .B(n3370), .A(n6508), .Z(n11173) );
  NAND U5626 ( .A(n3371), .B(n11173), .Z(n3372) );
  AND U5627 ( .A(n11175), .B(n3372), .Z(n3374) );
  ANDN U5628 ( .B(y[712]), .A(x[712]), .Z(n3373) );
  OR U5629 ( .A(n3374), .B(n3373), .Z(n3375) );
  NANDN U5630 ( .A(y[713]), .B(x[713]), .Z(n6506) );
  NAND U5631 ( .A(n3375), .B(n11177), .Z(n3376) );
  NANDN U5632 ( .A(x[713]), .B(y[713]), .Z(n6504) );
  NAND U5633 ( .A(n3376), .B(n6504), .Z(n3377) );
  NANDN U5634 ( .A(y[714]), .B(x[714]), .Z(n11182) );
  NAND U5635 ( .A(n3377), .B(n11182), .Z(n3378) );
  NANDN U5636 ( .A(n11184), .B(n3378), .Z(n3379) );
  AND U5637 ( .A(n11185), .B(n3379), .Z(n3382) );
  NANDN U5638 ( .A(x[717]), .B(y[717]), .Z(n3381) );
  NANDN U5639 ( .A(x[716]), .B(y[716]), .Z(n3380) );
  NAND U5640 ( .A(n3381), .B(n3380), .Z(n11188) );
  OR U5641 ( .A(n3382), .B(n11188), .Z(n3383) );
  AND U5642 ( .A(n11190), .B(n3383), .Z(n3385) );
  NANDN U5643 ( .A(x[718]), .B(y[718]), .Z(n3384) );
  ANDN U5644 ( .B(y[719]), .A(x[719]), .Z(n3386) );
  ANDN U5645 ( .B(n3384), .A(n3386), .Z(n11193) );
  NANDN U5646 ( .A(n3385), .B(n11193), .Z(n3388) );
  NANDN U5647 ( .A(y[718]), .B(x[718]), .Z(n11191) );
  ANDN U5648 ( .B(x[719]), .A(y[719]), .Z(n11195) );
  ANDN U5649 ( .B(n11191), .A(n11195), .Z(n3387) );
  OR U5650 ( .A(n3387), .B(n3386), .Z(n7517) );
  NAND U5651 ( .A(n3388), .B(n7517), .Z(n3391) );
  NANDN U5652 ( .A(x[720]), .B(y[720]), .Z(n3390) );
  ANDN U5653 ( .B(n3390), .A(n3389), .Z(n11200) );
  NAND U5654 ( .A(n3391), .B(n11200), .Z(n3392) );
  NANDN U5655 ( .A(n7521), .B(n3392), .Z(n3393) );
  NANDN U5656 ( .A(n11204), .B(n3393), .Z(n3394) );
  NANDN U5657 ( .A(y[723]), .B(x[723]), .Z(n11205) );
  NAND U5658 ( .A(n3394), .B(n11205), .Z(n3395) );
  NANDN U5659 ( .A(n11210), .B(n3395), .Z(n3396) );
  NANDN U5660 ( .A(n7526), .B(n3396), .Z(n3405) );
  NANDN U5661 ( .A(x[729]), .B(y[729]), .Z(n3398) );
  NANDN U5662 ( .A(x[728]), .B(y[728]), .Z(n3397) );
  AND U5663 ( .A(n3398), .B(n3397), .Z(n3404) );
  NANDN U5664 ( .A(x[726]), .B(y[726]), .Z(n3399) );
  NANDN U5665 ( .A(y[727]), .B(n3399), .Z(n3402) );
  XNOR U5666 ( .A(n3399), .B(y[727]), .Z(n3400) );
  NAND U5667 ( .A(n3400), .B(x[727]), .Z(n3401) );
  NAND U5668 ( .A(n3402), .B(n3401), .Z(n3403) );
  NAND U5669 ( .A(n3404), .B(n3403), .Z(n11216) );
  ANDN U5670 ( .B(n3405), .A(n11216), .Z(n3406) );
  OR U5671 ( .A(n11218), .B(n3406), .Z(n3409) );
  NANDN U5672 ( .A(x[730]), .B(y[730]), .Z(n3408) );
  NANDN U5673 ( .A(x[731]), .B(y[731]), .Z(n3407) );
  AND U5674 ( .A(n3408), .B(n3407), .Z(n11219) );
  NAND U5675 ( .A(n3409), .B(n11219), .Z(n3410) );
  NANDN U5676 ( .A(y[731]), .B(x[731]), .Z(n11222) );
  NAND U5677 ( .A(n3410), .B(n11222), .Z(n3413) );
  NANDN U5678 ( .A(x[732]), .B(y[732]), .Z(n3412) );
  ANDN U5679 ( .B(n3412), .A(n3411), .Z(n11225) );
  NAND U5680 ( .A(n3413), .B(n11225), .Z(n3414) );
  NANDN U5681 ( .A(n7533), .B(n3414), .Z(n3415) );
  AND U5682 ( .A(n11230), .B(n3415), .Z(n3416) );
  OR U5683 ( .A(n11231), .B(n3416), .Z(n3418) );
  NANDN U5684 ( .A(x[738]), .B(y[738]), .Z(n3417) );
  ANDN U5685 ( .B(y[739]), .A(x[739]), .Z(n3420) );
  ANDN U5686 ( .B(n3417), .A(n3420), .Z(n11236) );
  NAND U5687 ( .A(n3418), .B(n11236), .Z(n3421) );
  NANDN U5688 ( .A(y[738]), .B(x[738]), .Z(n3419) );
  ANDN U5689 ( .B(x[739]), .A(y[739]), .Z(n11235) );
  ANDN U5690 ( .B(n3419), .A(n11235), .Z(n11233) );
  OR U5691 ( .A(n3420), .B(n11233), .Z(n7538) );
  NAND U5692 ( .A(n3421), .B(n7538), .Z(n3422) );
  NANDN U5693 ( .A(x[740]), .B(y[740]), .Z(n11238) );
  NAND U5694 ( .A(n3422), .B(n11238), .Z(n3423) );
  NANDN U5695 ( .A(n11242), .B(n3423), .Z(n3424) );
  NANDN U5696 ( .A(x[741]), .B(y[741]), .Z(n11243) );
  NAND U5697 ( .A(n3424), .B(n11243), .Z(n3425) );
  NANDN U5698 ( .A(n11245), .B(n3425), .Z(n3426) );
  NANDN U5699 ( .A(n11247), .B(n3426), .Z(n3427) );
  NANDN U5700 ( .A(y[744]), .B(x[744]), .Z(n11249) );
  ANDN U5701 ( .B(n3427), .A(n7548), .Z(n3430) );
  NANDN U5702 ( .A(x[745]), .B(y[745]), .Z(n3429) );
  NANDN U5703 ( .A(x[746]), .B(y[746]), .Z(n3428) );
  AND U5704 ( .A(n3429), .B(n3428), .Z(n7549) );
  NANDN U5705 ( .A(n3430), .B(n7549), .Z(n3431) );
  NANDN U5706 ( .A(n7551), .B(n3431), .Z(n3432) );
  NANDN U5707 ( .A(x[747]), .B(y[747]), .Z(n11259) );
  NAND U5708 ( .A(n3432), .B(n11259), .Z(n3433) );
  NANDN U5709 ( .A(n11262), .B(n3433), .Z(n3434) );
  NANDN U5710 ( .A(n11263), .B(n3434), .Z(n3439) );
  XNOR U5711 ( .A(x[751]), .B(y[751]), .Z(n3436) );
  NANDN U5712 ( .A(y[750]), .B(x[750]), .Z(n3435) );
  NAND U5713 ( .A(n3436), .B(n3435), .Z(n3437) );
  AND U5714 ( .A(n3438), .B(n3437), .Z(n6502) );
  ANDN U5715 ( .B(n3439), .A(n6502), .Z(n3441) );
  ANDN U5716 ( .B(y[752]), .A(x[752]), .Z(n3440) );
  OR U5717 ( .A(n3441), .B(n3440), .Z(n3442) );
  NANDN U5718 ( .A(n6501), .B(n3442), .Z(n3443) );
  NANDN U5719 ( .A(x[753]), .B(y[753]), .Z(n7561) );
  NAND U5720 ( .A(n3443), .B(n7561), .Z(n3446) );
  NANDN U5721 ( .A(y[754]), .B(x[754]), .Z(n3444) );
  NAND U5722 ( .A(n3445), .B(n3444), .Z(n11270) );
  ANDN U5723 ( .B(n3446), .A(n11270), .Z(n3447) );
  OR U5724 ( .A(n11272), .B(n3447), .Z(n3448) );
  NANDN U5725 ( .A(n11276), .B(n3448), .Z(n3451) );
  NANDN U5726 ( .A(x[758]), .B(y[758]), .Z(n3450) );
  ANDN U5727 ( .B(n3450), .A(n3449), .Z(n11278) );
  NAND U5728 ( .A(n3451), .B(n11278), .Z(n3452) );
  NANDN U5729 ( .A(n7572), .B(n3452), .Z(n3455) );
  NANDN U5730 ( .A(x[760]), .B(y[760]), .Z(n3454) );
  NANDN U5731 ( .A(x[761]), .B(y[761]), .Z(n3453) );
  AND U5732 ( .A(n3454), .B(n3453), .Z(n11283) );
  NAND U5733 ( .A(n3455), .B(n11283), .Z(n3460) );
  NANDN U5734 ( .A(y[762]), .B(x[762]), .Z(n3457) );
  NANDN U5735 ( .A(y[761]), .B(x[761]), .Z(n3456) );
  AND U5736 ( .A(n3457), .B(n3456), .Z(n3459) );
  NANDN U5737 ( .A(y[763]), .B(x[763]), .Z(n3458) );
  NAND U5738 ( .A(n3459), .B(n3458), .Z(n11286) );
  ANDN U5739 ( .B(n3460), .A(n11286), .Z(n3467) );
  NANDN U5740 ( .A(x[763]), .B(y[763]), .Z(n3462) );
  ANDN U5741 ( .B(y[764]), .A(x[764]), .Z(n3461) );
  ANDN U5742 ( .B(n3462), .A(n3461), .Z(n3466) );
  XNOR U5743 ( .A(y[763]), .B(x[763]), .Z(n3464) );
  ANDN U5744 ( .B(y[762]), .A(x[762]), .Z(n3463) );
  NAND U5745 ( .A(n3464), .B(n3463), .Z(n3465) );
  AND U5746 ( .A(n3466), .B(n3465), .Z(n11287) );
  NANDN U5747 ( .A(n3467), .B(n11287), .Z(n3468) );
  NANDN U5748 ( .A(n11290), .B(n3468), .Z(n3471) );
  NANDN U5749 ( .A(x[765]), .B(y[765]), .Z(n3470) );
  NANDN U5750 ( .A(x[766]), .B(y[766]), .Z(n3469) );
  AND U5751 ( .A(n3470), .B(n3469), .Z(n11292) );
  NAND U5752 ( .A(n3471), .B(n11292), .Z(n3472) );
  NANDN U5753 ( .A(n11294), .B(n3472), .Z(n3473) );
  NANDN U5754 ( .A(n11296), .B(n3473), .Z(n3474) );
  AND U5755 ( .A(n11297), .B(n3474), .Z(n3475) );
  NANDN U5756 ( .A(x[771]), .B(y[771]), .Z(n3477) );
  NANDN U5757 ( .A(n3475), .B(n11301), .Z(n3479) );
  NANDN U5758 ( .A(y[770]), .B(x[770]), .Z(n3476) );
  ANDN U5759 ( .B(x[771]), .A(y[771]), .Z(n11304) );
  ANDN U5760 ( .B(n3476), .A(n11304), .Z(n3478) );
  NANDN U5761 ( .A(n3478), .B(n3477), .Z(n7583) );
  NAND U5762 ( .A(n3479), .B(n7583), .Z(n3482) );
  NANDN U5763 ( .A(x[772]), .B(y[772]), .Z(n3481) );
  ANDN U5764 ( .B(n3481), .A(n3480), .Z(n11307) );
  NAND U5765 ( .A(n3482), .B(n11307), .Z(n3483) );
  NANDN U5766 ( .A(n7587), .B(n3483), .Z(n3484) );
  NANDN U5767 ( .A(n11312), .B(n3484), .Z(n3485) );
  NANDN U5768 ( .A(n11313), .B(n3485), .Z(n3487) );
  NANDN U5769 ( .A(x[778]), .B(y[778]), .Z(n3486) );
  ANDN U5770 ( .B(y[779]), .A(x[779]), .Z(n3489) );
  ANDN U5771 ( .B(n3486), .A(n3489), .Z(n11317) );
  NAND U5772 ( .A(n3487), .B(n11317), .Z(n3490) );
  NANDN U5773 ( .A(y[778]), .B(x[778]), .Z(n11315) );
  ANDN U5774 ( .B(x[779]), .A(y[779]), .Z(n11319) );
  ANDN U5775 ( .B(n11315), .A(n11319), .Z(n3488) );
  OR U5776 ( .A(n3489), .B(n3488), .Z(n7591) );
  NAND U5777 ( .A(n3490), .B(n7591), .Z(n3491) );
  AND U5778 ( .A(n11323), .B(n3491), .Z(n3496) );
  NANDN U5779 ( .A(y[782]), .B(x[782]), .Z(n3493) );
  NANDN U5780 ( .A(y[781]), .B(x[781]), .Z(n3492) );
  NAND U5781 ( .A(n3493), .B(n3492), .Z(n11326) );
  ANDN U5782 ( .B(x[780]), .A(y[780]), .Z(n11322) );
  NANDN U5783 ( .A(n3494), .B(n11322), .Z(n3495) );
  NANDN U5784 ( .A(n11326), .B(n3495), .Z(n7595) );
  OR U5785 ( .A(n3496), .B(n7595), .Z(n3497) );
  NANDN U5786 ( .A(n11328), .B(n3497), .Z(n3498) );
  AND U5787 ( .A(n11329), .B(n3498), .Z(n3505) );
  NANDN U5788 ( .A(x[786]), .B(y[786]), .Z(n3504) );
  ANDN U5789 ( .B(y[784]), .A(x[784]), .Z(n3499) );
  OR U5790 ( .A(n3499), .B(y[785]), .Z(n3502) );
  XOR U5791 ( .A(y[785]), .B(n3499), .Z(n3500) );
  NAND U5792 ( .A(n3500), .B(x[785]), .Z(n3501) );
  NAND U5793 ( .A(n3502), .B(n3501), .Z(n3503) );
  NAND U5794 ( .A(n3504), .B(n3503), .Z(n11331) );
  OR U5795 ( .A(n3505), .B(n11331), .Z(n3508) );
  NANDN U5796 ( .A(y[786]), .B(x[786]), .Z(n3507) );
  NANDN U5797 ( .A(y[787]), .B(x[787]), .Z(n3506) );
  AND U5798 ( .A(n3507), .B(n3506), .Z(n11333) );
  NAND U5799 ( .A(n3508), .B(n11333), .Z(n3511) );
  NANDN U5800 ( .A(x[788]), .B(y[788]), .Z(n3510) );
  NANDN U5801 ( .A(x[787]), .B(y[787]), .Z(n3509) );
  NAND U5802 ( .A(n3510), .B(n3509), .Z(n11336) );
  ANDN U5803 ( .B(n3511), .A(n11336), .Z(n3514) );
  NANDN U5804 ( .A(y[789]), .B(x[789]), .Z(n3513) );
  NANDN U5805 ( .A(y[788]), .B(x[788]), .Z(n3512) );
  AND U5806 ( .A(n3513), .B(n3512), .Z(n11337) );
  NANDN U5807 ( .A(n3514), .B(n11337), .Z(n3515) );
  NANDN U5808 ( .A(x[789]), .B(y[789]), .Z(n11339) );
  NAND U5809 ( .A(n3515), .B(n11339), .Z(n3516) );
  NANDN U5810 ( .A(y[790]), .B(x[790]), .Z(n11341) );
  NAND U5811 ( .A(n3516), .B(n11341), .Z(n3517) );
  NANDN U5812 ( .A(n11343), .B(n3517), .Z(n3518) );
  NANDN U5813 ( .A(y[791]), .B(x[791]), .Z(n11346) );
  NAND U5814 ( .A(n3518), .B(n11346), .Z(n3519) );
  AND U5815 ( .A(n11350), .B(n3519), .Z(n3520) );
  NOR U5816 ( .A(n11352), .B(n3520), .Z(n3522) );
  ANDN U5817 ( .B(x[792]), .A(y[792]), .Z(n11345) );
  NAND U5818 ( .A(n3521), .B(n11345), .Z(n7608) );
  NAND U5819 ( .A(n3522), .B(n7608), .Z(n3523) );
  AND U5820 ( .A(n11353), .B(n3523), .Z(n3524) );
  NANDN U5821 ( .A(y[795]), .B(x[795]), .Z(n11357) );
  NANDN U5822 ( .A(n3524), .B(n11357), .Z(n3527) );
  NANDN U5823 ( .A(x[796]), .B(y[796]), .Z(n3526) );
  ANDN U5824 ( .B(n3526), .A(n3525), .Z(n11359) );
  NAND U5825 ( .A(n3527), .B(n11359), .Z(n3528) );
  NANDN U5826 ( .A(n7621), .B(n3528), .Z(n3529) );
  NANDN U5827 ( .A(y[798]), .B(x[798]), .Z(n11363) );
  NANDN U5828 ( .A(n3529), .B(n11363), .Z(n3530) );
  NANDN U5829 ( .A(n11366), .B(n3530), .Z(n3531) );
  NANDN U5830 ( .A(y[799]), .B(x[799]), .Z(n11369) );
  NAND U5831 ( .A(n3531), .B(n11369), .Z(n3534) );
  NANDN U5832 ( .A(x[800]), .B(y[800]), .Z(n3533) );
  ANDN U5833 ( .B(n3533), .A(n3532), .Z(n11371) );
  NAND U5834 ( .A(n3534), .B(n11371), .Z(n3535) );
  NANDN U5835 ( .A(n7629), .B(n3535), .Z(n3538) );
  NANDN U5836 ( .A(x[802]), .B(y[802]), .Z(n3537) );
  NANDN U5837 ( .A(x[803]), .B(y[803]), .Z(n3536) );
  AND U5838 ( .A(n3537), .B(n3536), .Z(n11375) );
  NAND U5839 ( .A(n3538), .B(n11375), .Z(n3539) );
  NANDN U5840 ( .A(n11378), .B(n3539), .Z(n3542) );
  NANDN U5841 ( .A(x[804]), .B(y[804]), .Z(n3541) );
  NANDN U5842 ( .A(x[805]), .B(y[805]), .Z(n3540) );
  AND U5843 ( .A(n3541), .B(n3540), .Z(n11379) );
  NAND U5844 ( .A(n3542), .B(n11379), .Z(n3545) );
  NANDN U5845 ( .A(y[806]), .B(x[806]), .Z(n3544) );
  NANDN U5846 ( .A(y[805]), .B(x[805]), .Z(n3543) );
  NAND U5847 ( .A(n3544), .B(n3543), .Z(n11382) );
  ANDN U5848 ( .B(n3545), .A(n11382), .Z(n3548) );
  NANDN U5849 ( .A(x[806]), .B(y[806]), .Z(n3547) );
  NANDN U5850 ( .A(x[807]), .B(y[807]), .Z(n3546) );
  AND U5851 ( .A(n3547), .B(n3546), .Z(n11383) );
  NANDN U5852 ( .A(n3548), .B(n11383), .Z(n3549) );
  NANDN U5853 ( .A(n11384), .B(n3549), .Z(n3552) );
  NANDN U5854 ( .A(x[808]), .B(y[808]), .Z(n3551) );
  NANDN U5855 ( .A(x[809]), .B(y[809]), .Z(n3550) );
  AND U5856 ( .A(n3551), .B(n3550), .Z(n11385) );
  NAND U5857 ( .A(n3552), .B(n11385), .Z(n3553) );
  AND U5858 ( .A(n6499), .B(n3553), .Z(n3554) );
  NAND U5859 ( .A(n3555), .B(n3554), .Z(n3556) );
  NAND U5860 ( .A(n6498), .B(n3556), .Z(n3557) );
  AND U5861 ( .A(n11389), .B(n3557), .Z(n3558) );
  NOR U5862 ( .A(n10009), .B(n3558), .Z(n3559) );
  NANDN U5863 ( .A(x[811]), .B(y[811]), .Z(n6497) );
  NAND U5864 ( .A(n3559), .B(n6497), .Z(n3565) );
  NANDN U5865 ( .A(y[815]), .B(x[815]), .Z(n3561) );
  NANDN U5866 ( .A(y[814]), .B(x[814]), .Z(n3560) );
  NAND U5867 ( .A(n3561), .B(n3560), .Z(n11390) );
  ANDN U5868 ( .B(x[813]), .A(y[813]), .Z(n10010) );
  NANDN U5869 ( .A(y[812]), .B(x[812]), .Z(n3562) );
  NANDN U5870 ( .A(n10010), .B(n3562), .Z(n11388) );
  NANDN U5871 ( .A(n3563), .B(n11388), .Z(n3564) );
  NANDN U5872 ( .A(n11390), .B(n3564), .Z(n7642) );
  ANDN U5873 ( .B(n3565), .A(n7642), .Z(n3572) );
  NANDN U5874 ( .A(x[815]), .B(y[815]), .Z(n3567) );
  ANDN U5875 ( .B(y[816]), .A(x[816]), .Z(n3566) );
  ANDN U5876 ( .B(n3567), .A(n3566), .Z(n3571) );
  XNOR U5877 ( .A(y[815]), .B(x[815]), .Z(n3569) );
  ANDN U5878 ( .B(y[814]), .A(x[814]), .Z(n3568) );
  NAND U5879 ( .A(n3569), .B(n3568), .Z(n3570) );
  AND U5880 ( .A(n3571), .B(n3570), .Z(n11391) );
  NANDN U5881 ( .A(n3572), .B(n11391), .Z(n3573) );
  NANDN U5882 ( .A(n11392), .B(n3573), .Z(n3574) );
  NANDN U5883 ( .A(x[817]), .B(y[817]), .Z(n11393) );
  NAND U5884 ( .A(n3574), .B(n11393), .Z(n3575) );
  NANDN U5885 ( .A(y[818]), .B(x[818]), .Z(n11394) );
  NAND U5886 ( .A(n3575), .B(n11394), .Z(n3576) );
  NANDN U5887 ( .A(n11395), .B(n3576), .Z(n3577) );
  AND U5888 ( .A(n11397), .B(n3577), .Z(n3580) );
  NANDN U5889 ( .A(x[820]), .B(y[820]), .Z(n3579) );
  ANDN U5890 ( .B(n3579), .A(n3578), .Z(n11398) );
  NANDN U5891 ( .A(n3580), .B(n11398), .Z(n3581) );
  NANDN U5892 ( .A(n7654), .B(n3581), .Z(n3582) );
  NAND U5893 ( .A(n3582), .B(n11401), .Z(n3584) );
  ANDN U5894 ( .B(y[824]), .A(x[824]), .Z(n3583) );
  OR U5895 ( .A(n3584), .B(n3583), .Z(n3586) );
  NANDN U5896 ( .A(y[824]), .B(x[824]), .Z(n3585) );
  ANDN U5897 ( .B(x[825]), .A(y[825]), .Z(n6495) );
  ANDN U5898 ( .B(n3585), .A(n6495), .Z(n11403) );
  NAND U5899 ( .A(n3586), .B(n11403), .Z(n3587) );
  NANDN U5900 ( .A(x[825]), .B(y[825]), .Z(n6494) );
  NAND U5901 ( .A(n3587), .B(n6494), .Z(n3588) );
  NANDN U5902 ( .A(x[826]), .B(y[826]), .Z(n7659) );
  NANDN U5903 ( .A(n3588), .B(n7659), .Z(n3589) );
  NANDN U5904 ( .A(n11408), .B(n3589), .Z(n3590) );
  ANDN U5905 ( .B(y[827]), .A(x[827]), .Z(n7663) );
  ANDN U5906 ( .B(n3590), .A(n7663), .Z(n3592) );
  ANDN U5907 ( .B(x[828]), .A(y[828]), .Z(n3591) );
  OR U5908 ( .A(n3592), .B(n3591), .Z(n3593) );
  NANDN U5909 ( .A(n7661), .B(n3593), .Z(n3594) );
  NANDN U5910 ( .A(y[829]), .B(x[829]), .Z(n7667) );
  NAND U5911 ( .A(n3594), .B(n7667), .Z(n3596) );
  NANDN U5912 ( .A(x[831]), .B(y[831]), .Z(n3597) );
  NANDN U5913 ( .A(x[830]), .B(y[830]), .Z(n3595) );
  AND U5914 ( .A(n3597), .B(n3595), .Z(n11413) );
  NAND U5915 ( .A(n3596), .B(n11413), .Z(n3600) );
  NANDN U5916 ( .A(y[830]), .B(x[830]), .Z(n7671) );
  ANDN U5917 ( .B(x[831]), .A(y[831]), .Z(n7674) );
  ANDN U5918 ( .B(n7671), .A(n7674), .Z(n3598) );
  NANDN U5919 ( .A(n3598), .B(n3597), .Z(n3599) );
  NANDN U5920 ( .A(y[832]), .B(x[832]), .Z(n7676) );
  NAND U5921 ( .A(n3599), .B(n7676), .Z(n11416) );
  ANDN U5922 ( .B(n3600), .A(n11416), .Z(n3603) );
  NANDN U5923 ( .A(x[832]), .B(y[832]), .Z(n3602) );
  NANDN U5924 ( .A(x[833]), .B(y[833]), .Z(n3601) );
  AND U5925 ( .A(n3602), .B(n3601), .Z(n11417) );
  NANDN U5926 ( .A(n3603), .B(n11417), .Z(n3604) );
  NANDN U5927 ( .A(n11419), .B(n3604), .Z(n3605) );
  NANDN U5928 ( .A(n11421), .B(n3605), .Z(n3606) );
  NANDN U5929 ( .A(n11424), .B(n3606), .Z(n3607) );
  ANDN U5930 ( .B(y[837]), .A(x[837]), .Z(n7691) );
  NAND U5931 ( .A(n3607), .B(n11425), .Z(n3608) );
  AND U5932 ( .A(n11427), .B(n3608), .Z(n3609) );
  OR U5933 ( .A(n11430), .B(n3609), .Z(n3612) );
  NANDN U5934 ( .A(y[839]), .B(x[839]), .Z(n3611) );
  NANDN U5935 ( .A(y[840]), .B(x[840]), .Z(n3610) );
  AND U5936 ( .A(n3611), .B(n3610), .Z(n11432) );
  NAND U5937 ( .A(n3612), .B(n11432), .Z(n3613) );
  NANDN U5938 ( .A(x[840]), .B(y[840]), .Z(n11433) );
  NAND U5939 ( .A(n3613), .B(n11433), .Z(n3614) );
  NANDN U5940 ( .A(y[841]), .B(x[841]), .Z(n11438) );
  NAND U5941 ( .A(n3614), .B(n11438), .Z(n3615) );
  NANDN U5942 ( .A(n7698), .B(n3615), .Z(n3616) );
  AND U5943 ( .A(n11441), .B(n3616), .Z(n3617) );
  OR U5944 ( .A(n11444), .B(n3617), .Z(n3620) );
  NANDN U5945 ( .A(y[844]), .B(x[844]), .Z(n3619) );
  NANDN U5946 ( .A(y[845]), .B(x[845]), .Z(n3618) );
  AND U5947 ( .A(n3619), .B(n3618), .Z(n11445) );
  NAND U5948 ( .A(n3620), .B(n11445), .Z(n3621) );
  NANDN U5949 ( .A(n11448), .B(n3621), .Z(n3624) );
  NANDN U5950 ( .A(y[846]), .B(x[846]), .Z(n3623) );
  NANDN U5951 ( .A(y[847]), .B(x[847]), .Z(n3622) );
  AND U5952 ( .A(n3623), .B(n3622), .Z(n11450) );
  NAND U5953 ( .A(n3624), .B(n11450), .Z(n3627) );
  ANDN U5954 ( .B(y[849]), .A(x[849]), .Z(n7709) );
  NANDN U5955 ( .A(x[848]), .B(y[848]), .Z(n3626) );
  NANDN U5956 ( .A(x[847]), .B(y[847]), .Z(n3625) );
  NAND U5957 ( .A(n3626), .B(n3625), .Z(n7705) );
  NOR U5958 ( .A(n7709), .B(n7705), .Z(n11451) );
  NAND U5959 ( .A(n3627), .B(n11451), .Z(n3632) );
  IV U5960 ( .A(x[850]), .Z(n6490) );
  IV U5961 ( .A(y[850]), .Z(n6489) );
  NANDN U5962 ( .A(n6490), .B(n6489), .Z(n3631) );
  NANDN U5963 ( .A(y[849]), .B(x[849]), .Z(n3629) );
  NANDN U5964 ( .A(y[848]), .B(x[848]), .Z(n3628) );
  AND U5965 ( .A(n3629), .B(n3628), .Z(n7707) );
  OR U5966 ( .A(n7709), .B(n7707), .Z(n3630) );
  NAND U5967 ( .A(n3631), .B(n3630), .Z(n11454) );
  ANDN U5968 ( .B(n3632), .A(n11454), .Z(n3634) );
  NANDN U5969 ( .A(x[850]), .B(y[850]), .Z(n3633) );
  ANDN U5970 ( .B(y[851]), .A(x[851]), .Z(n7715) );
  ANDN U5971 ( .B(n3633), .A(n7715), .Z(n11455) );
  NANDN U5972 ( .A(n3634), .B(n11455), .Z(n3635) );
  NANDN U5973 ( .A(y[851]), .B(x[851]), .Z(n11457) );
  NAND U5974 ( .A(n3635), .B(n11457), .Z(n3636) );
  NANDN U5975 ( .A(x[852]), .B(y[852]), .Z(n11459) );
  NAND U5976 ( .A(n3636), .B(n11459), .Z(n3639) );
  NANDN U5977 ( .A(y[852]), .B(x[852]), .Z(n3638) );
  NANDN U5978 ( .A(y[853]), .B(x[853]), .Z(n3637) );
  AND U5979 ( .A(n3638), .B(n3637), .Z(n11462) );
  NAND U5980 ( .A(n3639), .B(n11462), .Z(n3640) );
  NANDN U5981 ( .A(n11464), .B(n3640), .Z(n3641) );
  AND U5982 ( .A(n11465), .B(n3641), .Z(n3642) );
  OR U5983 ( .A(n11468), .B(n3642), .Z(n3645) );
  NANDN U5984 ( .A(y[856]), .B(x[856]), .Z(n3644) );
  NANDN U5985 ( .A(y[857]), .B(x[857]), .Z(n3643) );
  AND U5986 ( .A(n3644), .B(n3643), .Z(n11469) );
  NAND U5987 ( .A(n3645), .B(n11469), .Z(n3646) );
  NANDN U5988 ( .A(x[857]), .B(y[857]), .Z(n11472) );
  NAND U5989 ( .A(n3646), .B(n11472), .Z(n3649) );
  NANDN U5990 ( .A(y[858]), .B(x[858]), .Z(n3648) );
  ANDN U5991 ( .B(n3648), .A(n3647), .Z(n11475) );
  NAND U5992 ( .A(n3649), .B(n11475), .Z(n3650) );
  NANDN U5993 ( .A(n7726), .B(n3650), .Z(n3651) );
  AND U5994 ( .A(n11480), .B(n3651), .Z(n3652) );
  NANDN U5995 ( .A(x[861]), .B(y[861]), .Z(n11481) );
  NANDN U5996 ( .A(n3652), .B(n11481), .Z(n3653) );
  NANDN U5997 ( .A(n11484), .B(n3653), .Z(n3655) );
  NANDN U5998 ( .A(x[862]), .B(y[862]), .Z(n3654) );
  ANDN U5999 ( .B(y[863]), .A(x[863]), .Z(n7735) );
  ANDN U6000 ( .B(n3654), .A(n7735), .Z(n11485) );
  NAND U6001 ( .A(n3655), .B(n11485), .Z(n3656) );
  NANDN U6002 ( .A(y[863]), .B(x[863]), .Z(n11487) );
  NAND U6003 ( .A(n3656), .B(n11487), .Z(n3657) );
  NANDN U6004 ( .A(x[864]), .B(y[864]), .Z(n11489) );
  NAND U6005 ( .A(n3657), .B(n11489), .Z(n3658) );
  AND U6006 ( .A(n11492), .B(n3658), .Z(n3659) );
  OR U6007 ( .A(n11494), .B(n3659), .Z(n3662) );
  NANDN U6008 ( .A(y[866]), .B(x[866]), .Z(n3661) );
  NANDN U6009 ( .A(y[867]), .B(x[867]), .Z(n3660) );
  AND U6010 ( .A(n3661), .B(n3660), .Z(n11495) );
  NAND U6011 ( .A(n3662), .B(n11495), .Z(n3663) );
  NANDN U6012 ( .A(n11498), .B(n3663), .Z(n3666) );
  NANDN U6013 ( .A(y[868]), .B(x[868]), .Z(n3665) );
  NANDN U6014 ( .A(y[869]), .B(x[869]), .Z(n3664) );
  AND U6015 ( .A(n3665), .B(n3664), .Z(n11499) );
  NAND U6016 ( .A(n3666), .B(n11499), .Z(n3667) );
  NANDN U6017 ( .A(x[869]), .B(y[869]), .Z(n11502) );
  NAND U6018 ( .A(n3667), .B(n11502), .Z(n3668) );
  AND U6019 ( .A(n11505), .B(n3668), .Z(n3673) );
  NANDN U6020 ( .A(x[871]), .B(y[871]), .Z(n3670) );
  NANDN U6021 ( .A(x[872]), .B(y[872]), .Z(n3669) );
  NAND U6022 ( .A(n3670), .B(n3669), .Z(n11508) );
  ANDN U6023 ( .B(y[870]), .A(x[870]), .Z(n11504) );
  NANDN U6024 ( .A(n3671), .B(n11504), .Z(n3672) );
  NANDN U6025 ( .A(n11508), .B(n3672), .Z(n7746) );
  OR U6026 ( .A(n3673), .B(n7746), .Z(n3674) );
  NANDN U6027 ( .A(y[872]), .B(x[872]), .Z(n11510) );
  NAND U6028 ( .A(n3674), .B(n11510), .Z(n3675) );
  NANDN U6029 ( .A(x[873]), .B(y[873]), .Z(n11511) );
  NAND U6030 ( .A(n3675), .B(n11511), .Z(n3676) );
  NANDN U6031 ( .A(n11514), .B(n3676), .Z(n3678) );
  NANDN U6032 ( .A(x[874]), .B(y[874]), .Z(n3677) );
  ANDN U6033 ( .B(y[875]), .A(x[875]), .Z(n7755) );
  ANDN U6034 ( .B(n3677), .A(n7755), .Z(n11515) );
  NAND U6035 ( .A(n3678), .B(n11515), .Z(n3679) );
  AND U6036 ( .A(n11517), .B(n3679), .Z(n3680) );
  NANDN U6037 ( .A(x[876]), .B(y[876]), .Z(n11519) );
  NANDN U6038 ( .A(n3680), .B(n11519), .Z(n3683) );
  NANDN U6039 ( .A(y[876]), .B(x[876]), .Z(n3682) );
  NANDN U6040 ( .A(y[877]), .B(x[877]), .Z(n3681) );
  AND U6041 ( .A(n3682), .B(n3681), .Z(n11522) );
  NAND U6042 ( .A(n3683), .B(n11522), .Z(n3684) );
  NANDN U6043 ( .A(n11524), .B(n3684), .Z(n3687) );
  NANDN U6044 ( .A(y[878]), .B(x[878]), .Z(n3686) );
  NANDN U6045 ( .A(y[879]), .B(x[879]), .Z(n3685) );
  AND U6046 ( .A(n3686), .B(n3685), .Z(n11525) );
  NAND U6047 ( .A(n3687), .B(n11525), .Z(n3688) );
  NANDN U6048 ( .A(n11528), .B(n3688), .Z(n3689) );
  AND U6049 ( .A(n11529), .B(n3689), .Z(n3690) );
  NANDN U6050 ( .A(x[881]), .B(y[881]), .Z(n11532) );
  NANDN U6051 ( .A(n3690), .B(n11532), .Z(n3691) );
  NANDN U6052 ( .A(n11536), .B(n3691), .Z(n3692) );
  NANDN U6053 ( .A(n7766), .B(n3692), .Z(n3695) );
  NANDN U6054 ( .A(y[885]), .B(x[885]), .Z(n3694) );
  NANDN U6055 ( .A(y[886]), .B(x[886]), .Z(n3693) );
  AND U6056 ( .A(n3694), .B(n3693), .Z(n11543) );
  NAND U6057 ( .A(n3695), .B(n11543), .Z(n3696) );
  NANDN U6058 ( .A(n11546), .B(n3696), .Z(n3697) );
  NANDN U6059 ( .A(y[887]), .B(x[887]), .Z(n11547) );
  NAND U6060 ( .A(n3697), .B(n11547), .Z(n3698) );
  NANDN U6061 ( .A(x[888]), .B(y[888]), .Z(n11549) );
  NAND U6062 ( .A(n3698), .B(n11549), .Z(n3701) );
  NANDN U6063 ( .A(y[888]), .B(x[888]), .Z(n3700) );
  NANDN U6064 ( .A(y[889]), .B(x[889]), .Z(n3699) );
  AND U6065 ( .A(n3700), .B(n3699), .Z(n11552) );
  NAND U6066 ( .A(n3701), .B(n11552), .Z(n3704) );
  NANDN U6067 ( .A(x[890]), .B(y[890]), .Z(n3703) );
  NANDN U6068 ( .A(x[889]), .B(y[889]), .Z(n3702) );
  NAND U6069 ( .A(n3703), .B(n3702), .Z(n11554) );
  ANDN U6070 ( .B(n3704), .A(n11554), .Z(n3707) );
  NANDN U6071 ( .A(y[890]), .B(x[890]), .Z(n3706) );
  NANDN U6072 ( .A(y[891]), .B(x[891]), .Z(n3705) );
  AND U6073 ( .A(n3706), .B(n3705), .Z(n11555) );
  NANDN U6074 ( .A(n3707), .B(n11555), .Z(n3708) );
  NANDN U6075 ( .A(n11558), .B(n3708), .Z(n3711) );
  NANDN U6076 ( .A(y[892]), .B(x[892]), .Z(n3710) );
  NANDN U6077 ( .A(y[893]), .B(x[893]), .Z(n3709) );
  AND U6078 ( .A(n3710), .B(n3709), .Z(n11559) );
  NAND U6079 ( .A(n3711), .B(n11559), .Z(n3712) );
  NANDN U6080 ( .A(x[893]), .B(y[893]), .Z(n11562) );
  NAND U6081 ( .A(n3712), .B(n11562), .Z(n3713) );
  NANDN U6082 ( .A(y[894]), .B(x[894]), .Z(n11566) );
  NAND U6083 ( .A(n3713), .B(n11566), .Z(n3715) );
  ANDN U6084 ( .B(y[894]), .A(x[894]), .Z(n11564) );
  IV U6085 ( .A(y[895]), .Z(n10008) );
  OR U6086 ( .A(x[895]), .B(n10008), .Z(n3714) );
  NANDN U6087 ( .A(n11564), .B(n3714), .Z(n7779) );
  ANDN U6088 ( .B(n3715), .A(n7779), .Z(n3717) );
  NANDN U6089 ( .A(y[895]), .B(x[895]), .Z(n11570) );
  NANDN U6090 ( .A(y[896]), .B(x[896]), .Z(n3716) );
  AND U6091 ( .A(n11570), .B(n3716), .Z(n7780) );
  NANDN U6092 ( .A(n3717), .B(n7780), .Z(n3718) );
  NANDN U6093 ( .A(n7782), .B(n3718), .Z(n3721) );
  NANDN U6094 ( .A(y[897]), .B(x[897]), .Z(n3720) );
  NANDN U6095 ( .A(y[898]), .B(x[898]), .Z(n3719) );
  AND U6096 ( .A(n3720), .B(n3719), .Z(n11578) );
  NAND U6097 ( .A(n3721), .B(n11578), .Z(n3722) );
  NANDN U6098 ( .A(n11581), .B(n3722), .Z(n3723) );
  NANDN U6099 ( .A(y[899]), .B(x[899]), .Z(n11582) );
  NAND U6100 ( .A(n3723), .B(n11582), .Z(n3724) );
  AND U6101 ( .A(n11584), .B(n3724), .Z(n3725) );
  OR U6102 ( .A(n11587), .B(n3725), .Z(n3728) );
  NANDN U6103 ( .A(x[901]), .B(y[901]), .Z(n3727) );
  NANDN U6104 ( .A(x[902]), .B(y[902]), .Z(n3726) );
  AND U6105 ( .A(n3727), .B(n3726), .Z(n11589) );
  NAND U6106 ( .A(n3728), .B(n11589), .Z(n3729) );
  NANDN U6107 ( .A(n11591), .B(n3729), .Z(n3732) );
  NANDN U6108 ( .A(x[903]), .B(y[903]), .Z(n3731) );
  NANDN U6109 ( .A(x[904]), .B(y[904]), .Z(n3730) );
  AND U6110 ( .A(n3731), .B(n3730), .Z(n11592) );
  NAND U6111 ( .A(n3732), .B(n11592), .Z(n3733) );
  NANDN U6112 ( .A(n11595), .B(n3733), .Z(n3734) );
  AND U6113 ( .A(n11598), .B(n3734), .Z(n3737) );
  NANDN U6114 ( .A(y[907]), .B(x[907]), .Z(n3735) );
  NANDN U6115 ( .A(y[908]), .B(x[908]), .Z(n11602) );
  NAND U6116 ( .A(n3735), .B(n11602), .Z(n3739) );
  NANDN U6117 ( .A(y[906]), .B(x[906]), .Z(n3736) );
  NANDN U6118 ( .A(n3739), .B(n3736), .Z(n11601) );
  OR U6119 ( .A(n3737), .B(n11601), .Z(n3743) );
  ANDN U6120 ( .B(y[906]), .A(x[906]), .Z(n11596) );
  NANDN U6121 ( .A(x[907]), .B(y[907]), .Z(n11603) );
  NANDN U6122 ( .A(n11596), .B(n11603), .Z(n3738) );
  NANDN U6123 ( .A(n3739), .B(n3738), .Z(n3742) );
  NANDN U6124 ( .A(x[908]), .B(y[908]), .Z(n3741) );
  NANDN U6125 ( .A(x[909]), .B(y[909]), .Z(n3740) );
  NAND U6126 ( .A(n3741), .B(n3740), .Z(n11607) );
  ANDN U6127 ( .B(n3742), .A(n11607), .Z(n7795) );
  NAND U6128 ( .A(n3743), .B(n7795), .Z(n3744) );
  NANDN U6129 ( .A(n11609), .B(n3744), .Z(n3745) );
  NANDN U6130 ( .A(n11611), .B(n3745), .Z(n3746) );
  NANDN U6131 ( .A(y[911]), .B(x[911]), .Z(n11613) );
  NAND U6132 ( .A(n3746), .B(n11613), .Z(n3747) );
  AND U6133 ( .A(n11614), .B(n3747), .Z(n3750) );
  NANDN U6134 ( .A(y[912]), .B(x[912]), .Z(n3749) );
  NANDN U6135 ( .A(y[913]), .B(x[913]), .Z(n3748) );
  AND U6136 ( .A(n3749), .B(n3748), .Z(n11616) );
  NANDN U6137 ( .A(n3750), .B(n11616), .Z(n3751) );
  NANDN U6138 ( .A(n11619), .B(n3751), .Z(n3754) );
  NANDN U6139 ( .A(y[914]), .B(x[914]), .Z(n3753) );
  NANDN U6140 ( .A(y[915]), .B(x[915]), .Z(n3752) );
  AND U6141 ( .A(n3753), .B(n3752), .Z(n11620) );
  NAND U6142 ( .A(n3754), .B(n11620), .Z(n3755) );
  NANDN U6143 ( .A(n11623), .B(n3755), .Z(n3758) );
  NANDN U6144 ( .A(y[916]), .B(x[916]), .Z(n3757) );
  NANDN U6145 ( .A(y[917]), .B(x[917]), .Z(n3756) );
  AND U6146 ( .A(n3757), .B(n3756), .Z(n11625) );
  NAND U6147 ( .A(n3758), .B(n11625), .Z(n3759) );
  AND U6148 ( .A(n11627), .B(n3759), .Z(n3762) );
  NANDN U6149 ( .A(y[918]), .B(x[918]), .Z(n3761) );
  ANDN U6150 ( .B(n3761), .A(n3760), .Z(n11631) );
  NANDN U6151 ( .A(n3762), .B(n11631), .Z(n3763) );
  NANDN U6152 ( .A(n7808), .B(n3763), .Z(n3764) );
  NANDN U6153 ( .A(y[920]), .B(x[920]), .Z(n11634) );
  NAND U6154 ( .A(n3764), .B(n11634), .Z(n3765) );
  NANDN U6155 ( .A(x[921]), .B(y[921]), .Z(n11636) );
  NAND U6156 ( .A(n3765), .B(n11636), .Z(n3766) );
  NANDN U6157 ( .A(n11639), .B(n3766), .Z(n3768) );
  NANDN U6158 ( .A(x[923]), .B(y[923]), .Z(n7818) );
  NANDN U6159 ( .A(x[922]), .B(y[922]), .Z(n3767) );
  NAND U6160 ( .A(n7818), .B(n3767), .Z(n11641) );
  ANDN U6161 ( .B(n3768), .A(n11641), .Z(n3769) );
  NANDN U6162 ( .A(y[923]), .B(x[923]), .Z(n11643) );
  NANDN U6163 ( .A(n3769), .B(n11643), .Z(n3770) );
  NANDN U6164 ( .A(n11645), .B(n3770), .Z(n3771) );
  NANDN U6165 ( .A(n11647), .B(n3771), .Z(n3774) );
  NANDN U6166 ( .A(x[925]), .B(y[925]), .Z(n3773) );
  NANDN U6167 ( .A(x[926]), .B(y[926]), .Z(n3772) );
  AND U6168 ( .A(n3773), .B(n3772), .Z(n11648) );
  NAND U6169 ( .A(n3774), .B(n11648), .Z(n3775) );
  NANDN U6170 ( .A(n11651), .B(n3775), .Z(n3776) );
  AND U6171 ( .A(n11652), .B(n3776), .Z(n3777) );
  OR U6172 ( .A(n11654), .B(n3777), .Z(n3778) );
  NANDN U6173 ( .A(x[929]), .B(y[929]), .Z(n11657) );
  NAND U6174 ( .A(n3778), .B(n11657), .Z(n3779) );
  NANDN U6175 ( .A(n11660), .B(n3779), .Z(n3785) );
  ANDN U6176 ( .B(y[930]), .A(x[930]), .Z(n11656) );
  NANDN U6177 ( .A(x[931]), .B(y[931]), .Z(n10007) );
  NANDN U6178 ( .A(n11656), .B(n10007), .Z(n3780) );
  NANDN U6179 ( .A(n3781), .B(n3780), .Z(n3784) );
  NANDN U6180 ( .A(x[932]), .B(y[932]), .Z(n3783) );
  NANDN U6181 ( .A(x[933]), .B(y[933]), .Z(n3782) );
  NAND U6182 ( .A(n3783), .B(n3782), .Z(n11665) );
  ANDN U6183 ( .B(n3784), .A(n11665), .Z(n7828) );
  NAND U6184 ( .A(n3785), .B(n7828), .Z(n3786) );
  NANDN U6185 ( .A(n11667), .B(n3786), .Z(n3787) );
  AND U6186 ( .A(n11668), .B(n3787), .Z(n3788) );
  NANDN U6187 ( .A(y[935]), .B(x[935]), .Z(n11671) );
  NANDN U6188 ( .A(n3788), .B(n11671), .Z(n3789) );
  AND U6189 ( .A(n11672), .B(n3789), .Z(n3792) );
  NANDN U6190 ( .A(y[936]), .B(x[936]), .Z(n3791) );
  NANDN U6191 ( .A(y[937]), .B(x[937]), .Z(n3790) );
  AND U6192 ( .A(n3791), .B(n3790), .Z(n11674) );
  NANDN U6193 ( .A(n3792), .B(n11674), .Z(n3793) );
  NANDN U6194 ( .A(n11677), .B(n3793), .Z(n3796) );
  NANDN U6195 ( .A(y[938]), .B(x[938]), .Z(n3795) );
  NANDN U6196 ( .A(y[939]), .B(x[939]), .Z(n3794) );
  AND U6197 ( .A(n3795), .B(n3794), .Z(n11678) );
  NAND U6198 ( .A(n3796), .B(n11678), .Z(n3797) );
  NANDN U6199 ( .A(n11681), .B(n3797), .Z(n3800) );
  NANDN U6200 ( .A(y[940]), .B(x[940]), .Z(n3799) );
  NANDN U6201 ( .A(y[941]), .B(x[941]), .Z(n3798) );
  AND U6202 ( .A(n3799), .B(n3798), .Z(n11683) );
  NAND U6203 ( .A(n3800), .B(n11683), .Z(n3801) );
  NANDN U6204 ( .A(x[941]), .B(y[941]), .Z(n11685) );
  NAND U6205 ( .A(n3801), .B(n11685), .Z(n3803) );
  NANDN U6206 ( .A(y[942]), .B(x[942]), .Z(n3802) );
  ANDN U6207 ( .B(x[943]), .A(y[943]), .Z(n3805) );
  ANDN U6208 ( .B(n3802), .A(n3805), .Z(n11689) );
  NAND U6209 ( .A(n3803), .B(n11689), .Z(n3804) );
  AND U6210 ( .A(n6479), .B(n3804), .Z(n3806) );
  ANDN U6211 ( .B(y[942]), .A(x[942]), .Z(n11684) );
  NANDN U6212 ( .A(n3805), .B(n11684), .Z(n7842) );
  NAND U6213 ( .A(n3806), .B(n7842), .Z(n3807) );
  NANDN U6214 ( .A(y[944]), .B(x[944]), .Z(n11692) );
  NAND U6215 ( .A(n3807), .B(n11692), .Z(n3808) );
  AND U6216 ( .A(n3809), .B(n3808), .Z(n3810) );
  OR U6217 ( .A(n11697), .B(n3810), .Z(n3812) );
  NANDN U6218 ( .A(x[946]), .B(y[946]), .Z(n3811) );
  ANDN U6219 ( .B(y[947]), .A(x[947]), .Z(n7852) );
  ANDN U6220 ( .B(n3811), .A(n7852), .Z(n11698) );
  NAND U6221 ( .A(n3812), .B(n11698), .Z(n3813) );
  NANDN U6222 ( .A(y[947]), .B(x[947]), .Z(n11701) );
  NAND U6223 ( .A(n3813), .B(n11701), .Z(n3814) );
  NANDN U6224 ( .A(x[948]), .B(y[948]), .Z(n11702) );
  NAND U6225 ( .A(n3814), .B(n11702), .Z(n3817) );
  NANDN U6226 ( .A(y[948]), .B(x[948]), .Z(n3816) );
  NANDN U6227 ( .A(y[949]), .B(x[949]), .Z(n3815) );
  AND U6228 ( .A(n3816), .B(n3815), .Z(n11704) );
  NAND U6229 ( .A(n3817), .B(n11704), .Z(n3820) );
  NANDN U6230 ( .A(x[950]), .B(y[950]), .Z(n3819) );
  NANDN U6231 ( .A(x[949]), .B(y[949]), .Z(n3818) );
  NAND U6232 ( .A(n3819), .B(n3818), .Z(n11707) );
  ANDN U6233 ( .B(n3820), .A(n11707), .Z(n3823) );
  NANDN U6234 ( .A(y[950]), .B(x[950]), .Z(n3822) );
  NANDN U6235 ( .A(y[951]), .B(x[951]), .Z(n3821) );
  AND U6236 ( .A(n3822), .B(n3821), .Z(n11708) );
  NANDN U6237 ( .A(n3823), .B(n11708), .Z(n3824) );
  NANDN U6238 ( .A(n11711), .B(n3824), .Z(n3827) );
  NANDN U6239 ( .A(y[952]), .B(x[952]), .Z(n3826) );
  NANDN U6240 ( .A(y[953]), .B(x[953]), .Z(n3825) );
  AND U6241 ( .A(n3826), .B(n3825), .Z(n11713) );
  NAND U6242 ( .A(n3827), .B(n11713), .Z(n3828) );
  NANDN U6243 ( .A(x[953]), .B(y[953]), .Z(n11714) );
  NAND U6244 ( .A(n3828), .B(n11714), .Z(n3829) );
  NANDN U6245 ( .A(y[954]), .B(x[954]), .Z(n11719) );
  NAND U6246 ( .A(n3829), .B(n11719), .Z(n3831) );
  NANDN U6247 ( .A(x[954]), .B(y[954]), .Z(n11715) );
  NANDN U6248 ( .A(x[955]), .B(y[955]), .Z(n3830) );
  NAND U6249 ( .A(n11715), .B(n3830), .Z(n7863) );
  ANDN U6250 ( .B(n3831), .A(n7863), .Z(n3834) );
  NANDN U6251 ( .A(y[955]), .B(x[955]), .Z(n3833) );
  IV U6252 ( .A(x[956]), .Z(n11727) );
  OR U6253 ( .A(y[956]), .B(n11727), .Z(n3832) );
  AND U6254 ( .A(n3833), .B(n3832), .Z(n7864) );
  NANDN U6255 ( .A(n3834), .B(n7864), .Z(n3835) );
  NANDN U6256 ( .A(n7866), .B(n3835), .Z(n3838) );
  NANDN U6257 ( .A(y[957]), .B(x[957]), .Z(n3837) );
  NANDN U6258 ( .A(y[958]), .B(x[958]), .Z(n3836) );
  AND U6259 ( .A(n3837), .B(n3836), .Z(n11731) );
  NAND U6260 ( .A(n3838), .B(n11731), .Z(n3839) );
  ANDN U6261 ( .B(y[959]), .A(x[959]), .Z(n7872) );
  ANDN U6262 ( .B(y[958]), .A(x[958]), .Z(n7870) );
  NOR U6263 ( .A(n7872), .B(n7870), .Z(n11733) );
  NAND U6264 ( .A(n3839), .B(n11733), .Z(n3840) );
  NANDN U6265 ( .A(y[959]), .B(x[959]), .Z(n11736) );
  NAND U6266 ( .A(n3840), .B(n11736), .Z(n3841) );
  AND U6267 ( .A(n11737), .B(n3841), .Z(n3844) );
  NANDN U6268 ( .A(y[960]), .B(x[960]), .Z(n3843) );
  NANDN U6269 ( .A(y[961]), .B(x[961]), .Z(n3842) );
  AND U6270 ( .A(n3843), .B(n3842), .Z(n11739) );
  NANDN U6271 ( .A(n3844), .B(n11739), .Z(n3845) );
  NANDN U6272 ( .A(n11742), .B(n3845), .Z(n3848) );
  NANDN U6273 ( .A(y[962]), .B(x[962]), .Z(n3847) );
  NANDN U6274 ( .A(y[963]), .B(x[963]), .Z(n3846) );
  AND U6275 ( .A(n3847), .B(n3846), .Z(n11743) );
  NAND U6276 ( .A(n3848), .B(n11743), .Z(n3849) );
  NANDN U6277 ( .A(n11746), .B(n3849), .Z(n3852) );
  NANDN U6278 ( .A(y[964]), .B(x[964]), .Z(n3851) );
  NANDN U6279 ( .A(y[965]), .B(x[965]), .Z(n3850) );
  AND U6280 ( .A(n3851), .B(n3850), .Z(n11748) );
  NAND U6281 ( .A(n3852), .B(n11748), .Z(n3853) );
  AND U6282 ( .A(n11749), .B(n3853), .Z(n3854) );
  NANDN U6283 ( .A(y[966]), .B(x[966]), .Z(n11754) );
  NANDN U6284 ( .A(n3854), .B(n11754), .Z(n3855) );
  NANDN U6285 ( .A(n7883), .B(n3855), .Z(n3858) );
  NANDN U6286 ( .A(y[967]), .B(x[967]), .Z(n3857) );
  IV U6287 ( .A(x[968]), .Z(n11761) );
  OR U6288 ( .A(y[968]), .B(n11761), .Z(n3856) );
  AND U6289 ( .A(n3857), .B(n3856), .Z(n7884) );
  NAND U6290 ( .A(n3858), .B(n7884), .Z(n3859) );
  NANDN U6291 ( .A(n7886), .B(n3859), .Z(n3862) );
  NANDN U6292 ( .A(y[969]), .B(x[969]), .Z(n3861) );
  NANDN U6293 ( .A(y[970]), .B(x[970]), .Z(n3860) );
  AND U6294 ( .A(n3861), .B(n3860), .Z(n11766) );
  NAND U6295 ( .A(n3862), .B(n11766), .Z(n3865) );
  NANDN U6296 ( .A(x[970]), .B(y[970]), .Z(n3864) );
  NANDN U6297 ( .A(x[971]), .B(y[971]), .Z(n3863) );
  NAND U6298 ( .A(n3864), .B(n3863), .Z(n11769) );
  ANDN U6299 ( .B(n3865), .A(n11769), .Z(n3866) );
  NANDN U6300 ( .A(y[971]), .B(x[971]), .Z(n11771) );
  NANDN U6301 ( .A(n3866), .B(n11771), .Z(n3867) );
  NANDN U6302 ( .A(x[972]), .B(y[972]), .Z(n11772) );
  NAND U6303 ( .A(n3867), .B(n11772), .Z(n3870) );
  NANDN U6304 ( .A(y[972]), .B(x[972]), .Z(n3869) );
  NANDN U6305 ( .A(y[973]), .B(x[973]), .Z(n3868) );
  AND U6306 ( .A(n3869), .B(n3868), .Z(n11774) );
  NAND U6307 ( .A(n3870), .B(n11774), .Z(n3871) );
  NANDN U6308 ( .A(n11777), .B(n3871), .Z(n3874) );
  NANDN U6309 ( .A(y[974]), .B(x[974]), .Z(n3873) );
  NANDN U6310 ( .A(y[975]), .B(x[975]), .Z(n3872) );
  AND U6311 ( .A(n3873), .B(n3872), .Z(n11778) );
  NAND U6312 ( .A(n3874), .B(n11778), .Z(n3877) );
  NANDN U6313 ( .A(x[976]), .B(y[976]), .Z(n3876) );
  NANDN U6314 ( .A(x[975]), .B(y[975]), .Z(n3875) );
  NAND U6315 ( .A(n3876), .B(n3875), .Z(n11781) );
  ANDN U6316 ( .B(n3877), .A(n11781), .Z(n3880) );
  NANDN U6317 ( .A(y[976]), .B(x[976]), .Z(n3879) );
  NANDN U6318 ( .A(y[977]), .B(x[977]), .Z(n3878) );
  AND U6319 ( .A(n3879), .B(n3878), .Z(n11783) );
  NANDN U6320 ( .A(n3880), .B(n11783), .Z(n3881) );
  NANDN U6321 ( .A(n11785), .B(n3881), .Z(n3888) );
  NANDN U6322 ( .A(y[979]), .B(x[979]), .Z(n3883) );
  ANDN U6323 ( .B(x[980]), .A(y[980]), .Z(n3882) );
  ANDN U6324 ( .B(n3883), .A(n3882), .Z(n3887) );
  XNOR U6325 ( .A(x[979]), .B(y[979]), .Z(n3885) );
  ANDN U6326 ( .B(x[978]), .A(y[978]), .Z(n3884) );
  NAND U6327 ( .A(n3885), .B(n3884), .Z(n3886) );
  AND U6328 ( .A(n3887), .B(n3886), .Z(n11786) );
  NAND U6329 ( .A(n3888), .B(n11786), .Z(n3889) );
  NANDN U6330 ( .A(n11789), .B(n3889), .Z(n3892) );
  NANDN U6331 ( .A(y[981]), .B(x[981]), .Z(n3891) );
  NANDN U6332 ( .A(y[982]), .B(x[982]), .Z(n3890) );
  AND U6333 ( .A(n3891), .B(n3890), .Z(n11790) );
  NAND U6334 ( .A(n3892), .B(n11790), .Z(n3895) );
  NANDN U6335 ( .A(x[982]), .B(y[982]), .Z(n3894) );
  NANDN U6336 ( .A(x[983]), .B(y[983]), .Z(n3893) );
  NAND U6337 ( .A(n3894), .B(n3893), .Z(n11793) );
  ANDN U6338 ( .B(n3895), .A(n11793), .Z(n3896) );
  NANDN U6339 ( .A(y[983]), .B(x[983]), .Z(n11795) );
  NANDN U6340 ( .A(n3896), .B(n11795), .Z(n3897) );
  AND U6341 ( .A(n11796), .B(n3897), .Z(n3900) );
  NANDN U6342 ( .A(y[984]), .B(x[984]), .Z(n3899) );
  NANDN U6343 ( .A(y[985]), .B(x[985]), .Z(n3898) );
  AND U6344 ( .A(n3899), .B(n3898), .Z(n11798) );
  NANDN U6345 ( .A(n3900), .B(n11798), .Z(n3901) );
  NANDN U6346 ( .A(n11801), .B(n3901), .Z(n3904) );
  NANDN U6347 ( .A(y[986]), .B(x[986]), .Z(n3903) );
  NANDN U6348 ( .A(y[987]), .B(x[987]), .Z(n3902) );
  AND U6349 ( .A(n3903), .B(n3902), .Z(n11802) );
  NAND U6350 ( .A(n3904), .B(n11802), .Z(n3905) );
  NANDN U6351 ( .A(n11805), .B(n3905), .Z(n3908) );
  NANDN U6352 ( .A(y[988]), .B(x[988]), .Z(n3907) );
  NANDN U6353 ( .A(y[989]), .B(x[989]), .Z(n3906) );
  AND U6354 ( .A(n3907), .B(n3906), .Z(n11807) );
  NAND U6355 ( .A(n3908), .B(n11807), .Z(n3909) );
  NANDN U6356 ( .A(x[989]), .B(y[989]), .Z(n11809) );
  NAND U6357 ( .A(n3909), .B(n11809), .Z(n3910) );
  NANDN U6358 ( .A(n11812), .B(n3910), .Z(n3911) );
  NANDN U6359 ( .A(n7911), .B(n3911), .Z(n3912) );
  AND U6360 ( .A(n11818), .B(n3912), .Z(n3913) );
  OR U6361 ( .A(n11821), .B(n3913), .Z(n3914) );
  NANDN U6362 ( .A(y[995]), .B(x[995]), .Z(n11823) );
  NAND U6363 ( .A(n3914), .B(n11823), .Z(n3915) );
  NANDN U6364 ( .A(x[996]), .B(y[996]), .Z(n11824) );
  NAND U6365 ( .A(n3915), .B(n11824), .Z(n3918) );
  NANDN U6366 ( .A(y[996]), .B(x[996]), .Z(n3917) );
  NANDN U6367 ( .A(y[997]), .B(x[997]), .Z(n3916) );
  AND U6368 ( .A(n3917), .B(n3916), .Z(n11827) );
  NAND U6369 ( .A(n3918), .B(n11827), .Z(n3921) );
  NANDN U6370 ( .A(x[998]), .B(y[998]), .Z(n3920) );
  NANDN U6371 ( .A(x[997]), .B(y[997]), .Z(n3919) );
  NAND U6372 ( .A(n3920), .B(n3919), .Z(n11829) );
  ANDN U6373 ( .B(n3921), .A(n11829), .Z(n3924) );
  NANDN U6374 ( .A(y[998]), .B(x[998]), .Z(n3923) );
  NANDN U6375 ( .A(y[999]), .B(x[999]), .Z(n3922) );
  AND U6376 ( .A(n3923), .B(n3922), .Z(n11830) );
  NANDN U6377 ( .A(n3924), .B(n11830), .Z(n3925) );
  NANDN U6378 ( .A(n11833), .B(n3925), .Z(n3926) );
  AND U6379 ( .A(n11834), .B(n3926), .Z(n3927) );
  NANDN U6380 ( .A(x[1001]), .B(y[1001]), .Z(n11838) );
  NANDN U6381 ( .A(n3927), .B(n11838), .Z(n3930) );
  NANDN U6382 ( .A(y[1002]), .B(x[1002]), .Z(n3929) );
  ANDN U6383 ( .B(n3929), .A(n3928), .Z(n11841) );
  NAND U6384 ( .A(n3930), .B(n11841), .Z(n3931) );
  NANDN U6385 ( .A(n7924), .B(n3931), .Z(n3932) );
  NANDN U6386 ( .A(n11845), .B(n3932), .Z(n3933) );
  NANDN U6387 ( .A(x[1005]), .B(y[1005]), .Z(n11846) );
  NAND U6388 ( .A(n3933), .B(n11846), .Z(n3935) );
  NANDN U6389 ( .A(y[1005]), .B(x[1005]), .Z(n7926) );
  IV U6390 ( .A(x[1006]), .Z(n6474) );
  IV U6391 ( .A(y[1006]), .Z(n6473) );
  NANDN U6392 ( .A(n6474), .B(n6473), .Z(n3934) );
  NAND U6393 ( .A(n7926), .B(n3934), .Z(n11849) );
  ANDN U6394 ( .B(n3935), .A(n11849), .Z(n3937) );
  NANDN U6395 ( .A(x[1006]), .B(y[1006]), .Z(n3936) );
  ANDN U6396 ( .B(y[1007]), .A(x[1007]), .Z(n7934) );
  ANDN U6397 ( .B(n3936), .A(n7934), .Z(n11850) );
  NANDN U6398 ( .A(n3937), .B(n11850), .Z(n3938) );
  NANDN U6399 ( .A(y[1007]), .B(x[1007]), .Z(n11853) );
  NAND U6400 ( .A(n3938), .B(n11853), .Z(n3939) );
  NANDN U6401 ( .A(x[1008]), .B(y[1008]), .Z(n11854) );
  NAND U6402 ( .A(n3939), .B(n11854), .Z(n3942) );
  NANDN U6403 ( .A(y[1008]), .B(x[1008]), .Z(n3941) );
  NANDN U6404 ( .A(y[1009]), .B(x[1009]), .Z(n3940) );
  AND U6405 ( .A(n3941), .B(n3940), .Z(n11857) );
  NAND U6406 ( .A(n3942), .B(n11857), .Z(n3943) );
  NANDN U6407 ( .A(n11859), .B(n3943), .Z(n3944) );
  AND U6408 ( .A(n11860), .B(n3944), .Z(n3945) );
  OR U6409 ( .A(n11863), .B(n3945), .Z(n3948) );
  NANDN U6410 ( .A(y[1012]), .B(x[1012]), .Z(n3947) );
  NANDN U6411 ( .A(y[1013]), .B(x[1013]), .Z(n3946) );
  AND U6412 ( .A(n3947), .B(n3946), .Z(n11864) );
  NAND U6413 ( .A(n3948), .B(n11864), .Z(n3949) );
  NANDN U6414 ( .A(x[1013]), .B(y[1013]), .Z(n11868) );
  NAND U6415 ( .A(n3949), .B(n11868), .Z(n3950) );
  NANDN U6416 ( .A(y[1014]), .B(x[1014]), .Z(n11870) );
  NAND U6417 ( .A(n3950), .B(n11870), .Z(n3951) );
  NANDN U6418 ( .A(n7945), .B(n3951), .Z(n3952) );
  AND U6419 ( .A(n11874), .B(n3952), .Z(n3953) );
  OR U6420 ( .A(n11876), .B(n3953), .Z(n3954) );
  AND U6421 ( .A(n3955), .B(n3954), .Z(n3959) );
  NANDN U6422 ( .A(x[1019]), .B(y[1019]), .Z(n3956) );
  NAND U6423 ( .A(n3957), .B(n3956), .Z(n7953) );
  NANDN U6424 ( .A(x[1018]), .B(y[1018]), .Z(n3958) );
  NANDN U6425 ( .A(n7953), .B(n3958), .Z(n11881) );
  OR U6426 ( .A(n3959), .B(n11881), .Z(n3960) );
  AND U6427 ( .A(n3961), .B(n3960), .Z(n3964) );
  NANDN U6428 ( .A(y[1020]), .B(x[1020]), .Z(n3963) );
  NANDN U6429 ( .A(y[1021]), .B(x[1021]), .Z(n3962) );
  NAND U6430 ( .A(n3963), .B(n3962), .Z(n7954) );
  ANDN U6431 ( .B(n3964), .A(n7954), .Z(n3966) );
  NANDN U6432 ( .A(x[1022]), .B(y[1022]), .Z(n3965) );
  ANDN U6433 ( .B(y[1021]), .A(x[1021]), .Z(n11884) );
  ANDN U6434 ( .B(n3965), .A(n11884), .Z(n7957) );
  NANDN U6435 ( .A(n3966), .B(n7957), .Z(n3967) );
  NANDN U6436 ( .A(n7959), .B(n3967), .Z(n3970) );
  NANDN U6437 ( .A(x[1023]), .B(y[1023]), .Z(n3969) );
  NANDN U6438 ( .A(x[1024]), .B(y[1024]), .Z(n3968) );
  AND U6439 ( .A(n3969), .B(n3968), .Z(n11893) );
  NAND U6440 ( .A(n3970), .B(n11893), .Z(n3971) );
  NANDN U6441 ( .A(n11896), .B(n3971), .Z(n3972) );
  ANDN U6442 ( .B(y[1025]), .A(x[1025]), .Z(n7963) );
  ANDN U6443 ( .B(n3972), .A(n7963), .Z(n3973) );
  NAND U6444 ( .A(n3974), .B(n3973), .Z(n3975) );
  NAND U6445 ( .A(n6471), .B(n3975), .Z(n3976) );
  AND U6446 ( .A(n11901), .B(n3976), .Z(n3978) );
  NANDN U6447 ( .A(y[1027]), .B(x[1027]), .Z(n6470) );
  NANDN U6448 ( .A(y[1028]), .B(x[1028]), .Z(n11904) );
  NAND U6449 ( .A(n6470), .B(n11904), .Z(n3977) );
  OR U6450 ( .A(n3978), .B(n3977), .Z(n3979) );
  AND U6451 ( .A(n11905), .B(n3979), .Z(n3980) );
  ANDN U6452 ( .B(n11908), .A(n3980), .Z(n3981) );
  NANDN U6453 ( .A(y[1030]), .B(x[1030]), .Z(n6469) );
  NAND U6454 ( .A(n3981), .B(n6469), .Z(n3982) );
  AND U6455 ( .A(n11909), .B(n3982), .Z(n3983) );
  NAND U6456 ( .A(n3984), .B(n3983), .Z(n3985) );
  NAND U6457 ( .A(n3986), .B(n3985), .Z(n3987) );
  NANDN U6458 ( .A(x[1032]), .B(y[1032]), .Z(n7976) );
  AND U6459 ( .A(n3987), .B(n7976), .Z(n3989) );
  OR U6460 ( .A(n3989), .B(x[1033]), .Z(n3988) );
  AND U6461 ( .A(n6465), .B(n3988), .Z(n3992) );
  XOR U6462 ( .A(n3989), .B(x[1033]), .Z(n3990) );
  NAND U6463 ( .A(n3990), .B(y[1033]), .Z(n3991) );
  NAND U6464 ( .A(n3992), .B(n3991), .Z(n3993) );
  AND U6465 ( .A(n11919), .B(n3993), .Z(n3994) );
  OR U6466 ( .A(n11922), .B(n3994), .Z(n3997) );
  NANDN U6467 ( .A(y[1036]), .B(x[1036]), .Z(n3996) );
  NANDN U6468 ( .A(y[1037]), .B(x[1037]), .Z(n3995) );
  AND U6469 ( .A(n3996), .B(n3995), .Z(n11923) );
  NAND U6470 ( .A(n3997), .B(n11923), .Z(n3998) );
  NANDN U6471 ( .A(n11925), .B(n3998), .Z(n4005) );
  NANDN U6472 ( .A(y[1039]), .B(x[1039]), .Z(n4000) );
  ANDN U6473 ( .B(x[1040]), .A(y[1040]), .Z(n3999) );
  ANDN U6474 ( .B(n4000), .A(n3999), .Z(n4004) );
  XNOR U6475 ( .A(x[1039]), .B(y[1039]), .Z(n4002) );
  ANDN U6476 ( .B(x[1038]), .A(y[1038]), .Z(n4001) );
  NAND U6477 ( .A(n4002), .B(n4001), .Z(n4003) );
  AND U6478 ( .A(n4004), .B(n4003), .Z(n11927) );
  NAND U6479 ( .A(n4005), .B(n11927), .Z(n4006) );
  NANDN U6480 ( .A(n11930), .B(n4006), .Z(n4007) );
  ANDN U6481 ( .B(x[1042]), .A(y[1042]), .Z(n7989) );
  ANDN U6482 ( .B(n4007), .A(n7989), .Z(n4008) );
  NANDN U6483 ( .A(y[1041]), .B(x[1041]), .Z(n11931) );
  NAND U6484 ( .A(n4008), .B(n11931), .Z(n4009) );
  AND U6485 ( .A(n11933), .B(n4009), .Z(n4010) );
  NAND U6486 ( .A(n4011), .B(n4010), .Z(n4012) );
  NAND U6487 ( .A(n4013), .B(n4012), .Z(n4014) );
  NANDN U6488 ( .A(x[1044]), .B(y[1044]), .Z(n7992) );
  AND U6489 ( .A(n4014), .B(n7992), .Z(n4015) );
  NAND U6490 ( .A(n4016), .B(n4015), .Z(n4017) );
  NAND U6491 ( .A(n6462), .B(n4017), .Z(n4018) );
  AND U6492 ( .A(n6460), .B(n4018), .Z(n4021) );
  NANDN U6493 ( .A(y[1046]), .B(x[1046]), .Z(n4020) );
  NANDN U6494 ( .A(y[1047]), .B(x[1047]), .Z(n4019) );
  AND U6495 ( .A(n4020), .B(n4019), .Z(n11943) );
  NANDN U6496 ( .A(n4021), .B(n11943), .Z(n4024) );
  NANDN U6497 ( .A(x[1048]), .B(y[1048]), .Z(n4023) );
  NANDN U6498 ( .A(x[1047]), .B(y[1047]), .Z(n4022) );
  NAND U6499 ( .A(n4023), .B(n4022), .Z(n11945) );
  ANDN U6500 ( .B(n4024), .A(n11945), .Z(n4027) );
  NANDN U6501 ( .A(y[1048]), .B(x[1048]), .Z(n4026) );
  NANDN U6502 ( .A(y[1049]), .B(x[1049]), .Z(n4025) );
  AND U6503 ( .A(n4026), .B(n4025), .Z(n11947) );
  NANDN U6504 ( .A(n4027), .B(n11947), .Z(n4028) );
  NANDN U6505 ( .A(x[1049]), .B(y[1049]), .Z(n6459) );
  NAND U6506 ( .A(n4028), .B(n6459), .Z(n4029) );
  ANDN U6507 ( .B(x[1050]), .A(y[1050]), .Z(n8001) );
  ANDN U6508 ( .B(n4029), .A(n8001), .Z(n4030) );
  OR U6509 ( .A(n4031), .B(n4030), .Z(n4033) );
  ANDN U6510 ( .B(x[1052]), .A(y[1052]), .Z(n11956) );
  ANDN U6511 ( .B(x[1051]), .A(y[1051]), .Z(n8002) );
  NOR U6512 ( .A(n11956), .B(n8002), .Z(n4032) );
  NAND U6513 ( .A(n4033), .B(n4032), .Z(n4034) );
  ANDN U6514 ( .B(y[1052]), .A(x[1052]), .Z(n8004) );
  ANDN U6515 ( .B(y[1053]), .A(x[1053]), .Z(n8009) );
  NOR U6516 ( .A(n8004), .B(n8009), .Z(n11957) );
  NAND U6517 ( .A(n4034), .B(n11957), .Z(n4035) );
  NAND U6518 ( .A(n4036), .B(n4035), .Z(n4037) );
  NANDN U6519 ( .A(x[1054]), .B(y[1054]), .Z(n11961) );
  NAND U6520 ( .A(n4037), .B(n11961), .Z(n4038) );
  NAND U6521 ( .A(n4039), .B(n4038), .Z(n4040) );
  AND U6522 ( .A(n6457), .B(n4040), .Z(n4042) );
  OR U6523 ( .A(n4042), .B(x[1056]), .Z(n4041) );
  AND U6524 ( .A(n11970), .B(n4041), .Z(n4045) );
  XOR U6525 ( .A(n4042), .B(x[1056]), .Z(n4043) );
  NAND U6526 ( .A(n4043), .B(y[1056]), .Z(n4044) );
  NAND U6527 ( .A(n4045), .B(n4044), .Z(n4046) );
  NAND U6528 ( .A(n4047), .B(n4046), .Z(n4050) );
  NANDN U6529 ( .A(x[1059]), .B(y[1059]), .Z(n4049) );
  NANDN U6530 ( .A(x[1060]), .B(y[1060]), .Z(n4048) );
  AND U6531 ( .A(n4049), .B(n4048), .Z(n11973) );
  NAND U6532 ( .A(n4050), .B(n11973), .Z(n4051) );
  NANDN U6533 ( .A(n11976), .B(n4051), .Z(n4052) );
  NANDN U6534 ( .A(n8020), .B(n4052), .Z(n4053) );
  NAND U6535 ( .A(n4054), .B(n4053), .Z(n4055) );
  NAND U6536 ( .A(n8021), .B(n4055), .Z(n4056) );
  NANDN U6537 ( .A(x[1063]), .B(y[1063]), .Z(n11981) );
  NANDN U6538 ( .A(n4056), .B(n11981), .Z(n4057) );
  AND U6539 ( .A(n8023), .B(n4057), .Z(n4058) );
  NANDN U6540 ( .A(n4059), .B(n4058), .Z(n4061) );
  NANDN U6541 ( .A(x[1064]), .B(y[1064]), .Z(n4060) );
  NANDN U6542 ( .A(x[1065]), .B(y[1065]), .Z(n8031) );
  NAND U6543 ( .A(n4060), .B(n8031), .Z(n11986) );
  ANDN U6544 ( .B(n4061), .A(n11986), .Z(n4062) );
  ANDN U6545 ( .B(n11988), .A(n4062), .Z(n4063) );
  NANDN U6546 ( .A(y[1066]), .B(x[1066]), .Z(n6453) );
  NAND U6547 ( .A(n4063), .B(n6453), .Z(n4064) );
  NANDN U6548 ( .A(x[1066]), .B(y[1066]), .Z(n11989) );
  NAND U6549 ( .A(n4064), .B(n11989), .Z(n4065) );
  IV U6550 ( .A(x[1067]), .Z(n6451) );
  OR U6551 ( .A(n4065), .B(n6451), .Z(n4068) );
  XNOR U6552 ( .A(n4065), .B(x[1067]), .Z(n4066) );
  NANDN U6553 ( .A(y[1067]), .B(n4066), .Z(n4067) );
  AND U6554 ( .A(n4068), .B(n4067), .Z(n4070) );
  IV U6555 ( .A(x[1068]), .Z(n8036) );
  OR U6556 ( .A(n4070), .B(n8036), .Z(n4069) );
  AND U6557 ( .A(n8037), .B(n4069), .Z(n4073) );
  XNOR U6558 ( .A(n4070), .B(x[1068]), .Z(n4071) );
  NANDN U6559 ( .A(y[1068]), .B(n4071), .Z(n4072) );
  AND U6560 ( .A(n4073), .B(n4072), .Z(n4078) );
  NANDN U6561 ( .A(x[1070]), .B(y[1070]), .Z(n4075) );
  NANDN U6562 ( .A(x[1069]), .B(y[1069]), .Z(n4074) );
  AND U6563 ( .A(n4075), .B(n4074), .Z(n4077) );
  NANDN U6564 ( .A(x[1071]), .B(y[1071]), .Z(n4076) );
  NAND U6565 ( .A(n4077), .B(n4076), .Z(n11998) );
  NOR U6566 ( .A(n11998), .B(n12005), .Z(n8040) );
  NANDN U6567 ( .A(n4078), .B(n8040), .Z(n4079) );
  AND U6568 ( .A(n4080), .B(n4079), .Z(n4081) );
  ANDN U6569 ( .B(n12003), .A(n4081), .Z(n4082) );
  NANDN U6570 ( .A(n12012), .B(n4082), .Z(n4083) );
  NANDN U6571 ( .A(y[1075]), .B(x[1075]), .Z(n8046) );
  NAND U6572 ( .A(n4083), .B(n8046), .Z(n4084) );
  NANDN U6573 ( .A(y[1076]), .B(x[1076]), .Z(n12013) );
  NANDN U6574 ( .A(n4084), .B(n12013), .Z(n4085) );
  AND U6575 ( .A(n12016), .B(n4085), .Z(n4087) );
  NANDN U6576 ( .A(y[1077]), .B(x[1077]), .Z(n12017) );
  NANDN U6577 ( .A(y[1078]), .B(x[1078]), .Z(n8056) );
  AND U6578 ( .A(n12017), .B(n8056), .Z(n4086) );
  NANDN U6579 ( .A(n4087), .B(n4086), .Z(n4088) );
  NANDN U6580 ( .A(n12020), .B(n4088), .Z(n4091) );
  NANDN U6581 ( .A(y[1080]), .B(x[1080]), .Z(n4090) );
  NANDN U6582 ( .A(y[1081]), .B(x[1081]), .Z(n4089) );
  NAND U6583 ( .A(n4090), .B(n4089), .Z(n8060) );
  ANDN U6584 ( .B(n4091), .A(n8060), .Z(n4092) );
  NAND U6585 ( .A(n4093), .B(n4092), .Z(n4094) );
  NANDN U6586 ( .A(n12024), .B(n4094), .Z(n4095) );
  AND U6587 ( .A(n12025), .B(n4095), .Z(n4100) );
  NANDN U6588 ( .A(x[1084]), .B(y[1084]), .Z(n4097) );
  NANDN U6589 ( .A(x[1083]), .B(y[1083]), .Z(n4096) );
  AND U6590 ( .A(n4097), .B(n4096), .Z(n4099) );
  NANDN U6591 ( .A(x[1085]), .B(y[1085]), .Z(n4098) );
  NAND U6592 ( .A(n4099), .B(n4098), .Z(n12028) );
  OR U6593 ( .A(n4100), .B(n12028), .Z(n4101) );
  ANDN U6594 ( .B(x[1086]), .A(y[1086]), .Z(n8068) );
  ANDN U6595 ( .B(n4101), .A(n8068), .Z(n4106) );
  NANDN U6596 ( .A(y[1084]), .B(x[1084]), .Z(n4102) );
  NANDN U6597 ( .A(n4102), .B(x[1085]), .Z(n4105) );
  XNOR U6598 ( .A(n4102), .B(x[1085]), .Z(n4103) );
  NANDN U6599 ( .A(y[1085]), .B(n4103), .Z(n4104) );
  AND U6600 ( .A(n4105), .B(n4104), .Z(n12030) );
  NAND U6601 ( .A(n4106), .B(n12030), .Z(n4107) );
  AND U6602 ( .A(n12031), .B(n4107), .Z(n4108) );
  NANDN U6603 ( .A(x[1087]), .B(y[1087]), .Z(n12035) );
  NAND U6604 ( .A(n4108), .B(n12035), .Z(n4109) );
  NAND U6605 ( .A(n4110), .B(n4109), .Z(n4111) );
  ANDN U6606 ( .B(y[1089]), .A(x[1089]), .Z(n6448) );
  ANDN U6607 ( .B(y[1088]), .A(x[1088]), .Z(n8073) );
  NOR U6608 ( .A(n6448), .B(n8073), .Z(n12039) );
  NAND U6609 ( .A(n4111), .B(n12039), .Z(n4112) );
  NAND U6610 ( .A(n4113), .B(n4112), .Z(n4114) );
  NANDN U6611 ( .A(x[1090]), .B(y[1090]), .Z(n12043) );
  NAND U6612 ( .A(n4114), .B(n12043), .Z(n4115) );
  NAND U6613 ( .A(n4116), .B(n4115), .Z(n4117) );
  NAND U6614 ( .A(n6447), .B(n4117), .Z(n4118) );
  NAND U6615 ( .A(n4119), .B(n4118), .Z(n4120) );
  NAND U6616 ( .A(n4121), .B(n4120), .Z(n4122) );
  ANDN U6617 ( .B(x[1093]), .A(y[1093]), .Z(n8082) );
  ANDN U6618 ( .B(n4122), .A(n8082), .Z(n4127) );
  NANDN U6619 ( .A(x[1094]), .B(y[1094]), .Z(n4124) );
  NANDN U6620 ( .A(x[1093]), .B(y[1093]), .Z(n4123) );
  AND U6621 ( .A(n4124), .B(n4123), .Z(n4126) );
  NANDN U6622 ( .A(x[1095]), .B(y[1095]), .Z(n4125) );
  AND U6623 ( .A(n4126), .B(n4125), .Z(n12051) );
  NANDN U6624 ( .A(n4127), .B(n12051), .Z(n4128) );
  NANDN U6625 ( .A(y[1097]), .B(x[1097]), .Z(n4132) );
  ANDN U6626 ( .B(n4128), .A(n12053), .Z(n4133) );
  XNOR U6627 ( .A(y[1097]), .B(x[1097]), .Z(n4130) );
  NANDN U6628 ( .A(x[1096]), .B(y[1096]), .Z(n4129) );
  NAND U6629 ( .A(n4130), .B(n4129), .Z(n4131) );
  AND U6630 ( .A(n4132), .B(n4131), .Z(n6443) );
  OR U6631 ( .A(n4133), .B(n6443), .Z(n4134) );
  NANDN U6632 ( .A(n4134), .B(x[1098]), .Z(n4137) );
  XNOR U6633 ( .A(n4134), .B(x[1098]), .Z(n4135) );
  NANDN U6634 ( .A(y[1098]), .B(n4135), .Z(n4136) );
  NAND U6635 ( .A(n4137), .B(n4136), .Z(n4138) );
  NANDN U6636 ( .A(x[1099]), .B(y[1099]), .Z(n12059) );
  NAND U6637 ( .A(n4138), .B(n12059), .Z(n4139) );
  AND U6638 ( .A(n6441), .B(n4139), .Z(n4140) );
  NANDN U6639 ( .A(y[1100]), .B(x[1100]), .Z(n12061) );
  NAND U6640 ( .A(n4140), .B(n12061), .Z(n4141) );
  NANDN U6641 ( .A(n12064), .B(n4141), .Z(n4142) );
  AND U6642 ( .A(n12065), .B(n4142), .Z(n4143) );
  NANDN U6643 ( .A(y[1102]), .B(x[1102]), .Z(n6440) );
  NAND U6644 ( .A(n4143), .B(n6440), .Z(n4144) );
  NANDN U6645 ( .A(x[1102]), .B(y[1102]), .Z(n12067) );
  NAND U6646 ( .A(n4144), .B(n12067), .Z(n4145) );
  NAND U6647 ( .A(n4146), .B(n4145), .Z(n4147) );
  AND U6648 ( .A(n6439), .B(n4147), .Z(n4148) );
  NANDN U6649 ( .A(n4148), .B(y[1104]), .Z(n4151) );
  XNOR U6650 ( .A(n4148), .B(y[1104]), .Z(n4149) );
  NANDN U6651 ( .A(x[1104]), .B(n4149), .Z(n4150) );
  AND U6652 ( .A(n4151), .B(n4150), .Z(n4153) );
  NANDN U6653 ( .A(n4153), .B(y[1105]), .Z(n4152) );
  ANDN U6654 ( .B(y[1106]), .A(x[1106]), .Z(n8099) );
  ANDN U6655 ( .B(n4152), .A(n8099), .Z(n4156) );
  XNOR U6656 ( .A(n4153), .B(y[1105]), .Z(n4154) );
  NANDN U6657 ( .A(x[1105]), .B(n4154), .Z(n4155) );
  AND U6658 ( .A(n4156), .B(n4155), .Z(n4157) );
  OR U6659 ( .A(n12078), .B(n4157), .Z(n4158) );
  AND U6660 ( .A(n12079), .B(n4158), .Z(n4161) );
  NANDN U6661 ( .A(y[1109]), .B(x[1109]), .Z(n4160) );
  NANDN U6662 ( .A(y[1108]), .B(x[1108]), .Z(n4159) );
  NAND U6663 ( .A(n4160), .B(n4159), .Z(n12081) );
  OR U6664 ( .A(n4161), .B(n12081), .Z(n4164) );
  NANDN U6665 ( .A(x[1111]), .B(y[1111]), .Z(n4165) );
  NANDN U6666 ( .A(x[1109]), .B(y[1109]), .Z(n4163) );
  NANDN U6667 ( .A(x[1110]), .B(y[1110]), .Z(n4162) );
  NAND U6668 ( .A(n4163), .B(n4162), .Z(n8106) );
  ANDN U6669 ( .B(n4165), .A(n8106), .Z(n12083) );
  NAND U6670 ( .A(n4164), .B(n12083), .Z(n4171) );
  IV U6671 ( .A(n4165), .Z(n6437) );
  NANDN U6672 ( .A(y[1110]), .B(x[1110]), .Z(n4167) );
  NANDN U6673 ( .A(y[1111]), .B(x[1111]), .Z(n4166) );
  NAND U6674 ( .A(n4167), .B(n4166), .Z(n8108) );
  NANDN U6675 ( .A(n6437), .B(n8108), .Z(n4170) );
  NANDN U6676 ( .A(y[1112]), .B(x[1112]), .Z(n4168) );
  AND U6677 ( .A(n4169), .B(n4168), .Z(n8111) );
  NAND U6678 ( .A(n4170), .B(n8111), .Z(n12085) );
  ANDN U6679 ( .B(n4171), .A(n12085), .Z(n4172) );
  OR U6680 ( .A(n12087), .B(n4172), .Z(n4173) );
  NANDN U6681 ( .A(y[1114]), .B(x[1114]), .Z(n8116) );
  NAND U6682 ( .A(n4173), .B(n8116), .Z(n4174) );
  AND U6683 ( .A(n12092), .B(n4174), .Z(n4175) );
  ANDN U6684 ( .B(n4176), .A(n4175), .Z(n4177) );
  AND U6685 ( .A(n12093), .B(n4177), .Z(n4180) );
  NANDN U6686 ( .A(x[1118]), .B(y[1118]), .Z(n4179) );
  NANDN U6687 ( .A(x[1117]), .B(y[1117]), .Z(n4178) );
  NAND U6688 ( .A(n4179), .B(n4178), .Z(n12096) );
  OR U6689 ( .A(n4180), .B(n12096), .Z(n4181) );
  AND U6690 ( .A(n12097), .B(n4181), .Z(n4182) );
  OR U6691 ( .A(n12100), .B(n4182), .Z(n4185) );
  NANDN U6692 ( .A(y[1120]), .B(x[1120]), .Z(n4184) );
  NANDN U6693 ( .A(y[1121]), .B(x[1121]), .Z(n4183) );
  AND U6694 ( .A(n4184), .B(n4183), .Z(n12101) );
  NAND U6695 ( .A(n4185), .B(n12101), .Z(n4186) );
  NANDN U6696 ( .A(n12103), .B(n4186), .Z(n4189) );
  NANDN U6697 ( .A(y[1122]), .B(x[1122]), .Z(n4188) );
  NANDN U6698 ( .A(y[1123]), .B(x[1123]), .Z(n4187) );
  NAND U6699 ( .A(n4188), .B(n4187), .Z(n12106) );
  ANDN U6700 ( .B(n4189), .A(n12106), .Z(n4190) );
  NANDN U6701 ( .A(x[1123]), .B(y[1123]), .Z(n12107) );
  NANDN U6702 ( .A(n4190), .B(n12107), .Z(n4191) );
  NANDN U6703 ( .A(n8129), .B(n4191), .Z(n4192) );
  NANDN U6704 ( .A(x[1124]), .B(y[1124]), .Z(n8126) );
  NANDN U6705 ( .A(x[1125]), .B(y[1125]), .Z(n8132) );
  AND U6706 ( .A(n8126), .B(n8132), .Z(n12113) );
  NAND U6707 ( .A(n4192), .B(n12113), .Z(n4193) );
  NAND U6708 ( .A(n4194), .B(n4193), .Z(n4195) );
  NANDN U6709 ( .A(x[1126]), .B(y[1126]), .Z(n12111) );
  NAND U6710 ( .A(n4195), .B(n12111), .Z(n4196) );
  NAND U6711 ( .A(n4197), .B(n4196), .Z(n4198) );
  NAND U6712 ( .A(n6435), .B(n4198), .Z(n4199) );
  NAND U6713 ( .A(n4200), .B(n4199), .Z(n4201) );
  NAND U6714 ( .A(n4202), .B(n4201), .Z(n4203) );
  NAND U6715 ( .A(n4204), .B(n4203), .Z(n4210) );
  NANDN U6716 ( .A(x[1130]), .B(y[1130]), .Z(n8141) );
  NANDN U6717 ( .A(n8141), .B(n4205), .Z(n4208) );
  NANDN U6718 ( .A(x[1132]), .B(y[1132]), .Z(n4207) );
  NANDN U6719 ( .A(x[1131]), .B(y[1131]), .Z(n4206) );
  NAND U6720 ( .A(n4207), .B(n4206), .Z(n12127) );
  ANDN U6721 ( .B(n4208), .A(n12127), .Z(n4209) );
  NAND U6722 ( .A(n4210), .B(n4209), .Z(n4213) );
  NANDN U6723 ( .A(y[1132]), .B(x[1132]), .Z(n4212) );
  NANDN U6724 ( .A(y[1133]), .B(x[1133]), .Z(n4211) );
  AND U6725 ( .A(n4212), .B(n4211), .Z(n12129) );
  NAND U6726 ( .A(n4213), .B(n12129), .Z(n4214) );
  NANDN U6727 ( .A(n8147), .B(n4214), .Z(n4215) );
  NAND U6728 ( .A(n4216), .B(n4215), .Z(n4217) );
  NAND U6729 ( .A(n8148), .B(n4217), .Z(n4218) );
  NANDN U6730 ( .A(x[1135]), .B(y[1135]), .Z(n12136) );
  NANDN U6731 ( .A(n4218), .B(n12136), .Z(n4219) );
  AND U6732 ( .A(n12137), .B(n4219), .Z(n4220) );
  NANDN U6733 ( .A(y[1135]), .B(x[1135]), .Z(n8150) );
  NAND U6734 ( .A(n4220), .B(n8150), .Z(n4221) );
  NANDN U6735 ( .A(x[1136]), .B(y[1136]), .Z(n8154) );
  NANDN U6736 ( .A(x[1137]), .B(y[1137]), .Z(n8158) );
  NAND U6737 ( .A(n8154), .B(n8158), .Z(n12138) );
  ANDN U6738 ( .B(n4221), .A(n12138), .Z(n4222) );
  ANDN U6739 ( .B(n12139), .A(n4222), .Z(n4223) );
  NANDN U6740 ( .A(y[1138]), .B(x[1138]), .Z(n8163) );
  NAND U6741 ( .A(n4223), .B(n8163), .Z(n4224) );
  NANDN U6742 ( .A(x[1138]), .B(y[1138]), .Z(n12140) );
  NAND U6743 ( .A(n4224), .B(n12140), .Z(n4225) );
  IV U6744 ( .A(x[1139]), .Z(n8161) );
  OR U6745 ( .A(n4225), .B(n8161), .Z(n4228) );
  XNOR U6746 ( .A(n4225), .B(x[1139]), .Z(n4226) );
  NANDN U6747 ( .A(y[1139]), .B(n4226), .Z(n4227) );
  AND U6748 ( .A(n4228), .B(n4227), .Z(n4230) );
  NANDN U6749 ( .A(x[1140]), .B(n4230), .Z(n4229) );
  AND U6750 ( .A(n12144), .B(n4229), .Z(n4233) );
  XNOR U6751 ( .A(n4230), .B(x[1140]), .Z(n4231) );
  NAND U6752 ( .A(n4231), .B(y[1140]), .Z(n4232) );
  NAND U6753 ( .A(n4233), .B(n4232), .Z(n4234) );
  NAND U6754 ( .A(n4235), .B(n4234), .Z(n4236) );
  NANDN U6755 ( .A(n12146), .B(n4236), .Z(n4237) );
  NANDN U6756 ( .A(y[1143]), .B(x[1143]), .Z(n12148) );
  NAND U6757 ( .A(n4237), .B(n12148), .Z(n4238) );
  NANDN U6758 ( .A(n10002), .B(n4238), .Z(n4239) );
  NANDN U6759 ( .A(y[1146]), .B(x[1146]), .Z(n6429) );
  NAND U6760 ( .A(n4239), .B(n6429), .Z(n4242) );
  ANDN U6761 ( .B(x[1145]), .A(y[1145]), .Z(n10003) );
  NANDN U6762 ( .A(y[1144]), .B(x[1144]), .Z(n4240) );
  NANDN U6763 ( .A(n10003), .B(n4240), .Z(n12147) );
  NANDN U6764 ( .A(n4241), .B(n12147), .Z(n8178) );
  NANDN U6765 ( .A(n4242), .B(n8178), .Z(n4244) );
  NANDN U6766 ( .A(x[1146]), .B(y[1146]), .Z(n12149) );
  NANDN U6767 ( .A(x[1147]), .B(y[1147]), .Z(n12151) );
  AND U6768 ( .A(n12149), .B(n12151), .Z(n4243) );
  NAND U6769 ( .A(n4244), .B(n4243), .Z(n4245) );
  NANDN U6770 ( .A(y[1147]), .B(x[1147]), .Z(n6428) );
  NAND U6771 ( .A(n4245), .B(n6428), .Z(n4248) );
  NANDN U6772 ( .A(y[1148]), .B(x[1148]), .Z(n4246) );
  NANDN U6773 ( .A(n4247), .B(n4246), .Z(n12152) );
  OR U6774 ( .A(n4248), .B(n12152), .Z(n4249) );
  NANDN U6775 ( .A(n10000), .B(n4249), .Z(n4250) );
  NANDN U6776 ( .A(y[1150]), .B(x[1150]), .Z(n8189) );
  NAND U6777 ( .A(n4250), .B(n8189), .Z(n4251) );
  NANDN U6778 ( .A(x[1150]), .B(y[1150]), .Z(n10001) );
  NAND U6779 ( .A(n4251), .B(n10001), .Z(n4252) );
  NANDN U6780 ( .A(n4252), .B(x[1151]), .Z(n4255) );
  XNOR U6781 ( .A(n4252), .B(x[1151]), .Z(n4253) );
  NANDN U6782 ( .A(y[1151]), .B(n4253), .Z(n4254) );
  AND U6783 ( .A(n4255), .B(n4254), .Z(n4257) );
  OR U6784 ( .A(n4257), .B(y[1152]), .Z(n4256) );
  AND U6785 ( .A(n6427), .B(n4256), .Z(n4260) );
  XOR U6786 ( .A(n4257), .B(y[1152]), .Z(n4258) );
  NAND U6787 ( .A(n4258), .B(x[1152]), .Z(n4259) );
  NAND U6788 ( .A(n4260), .B(n4259), .Z(n4263) );
  NANDN U6789 ( .A(x[1153]), .B(y[1153]), .Z(n4262) );
  NANDN U6790 ( .A(x[1154]), .B(y[1154]), .Z(n4261) );
  AND U6791 ( .A(n4262), .B(n4261), .Z(n12161) );
  NAND U6792 ( .A(n4263), .B(n12161), .Z(n4264) );
  NANDN U6793 ( .A(n12164), .B(n4264), .Z(n4265) );
  NANDN U6794 ( .A(x[1155]), .B(y[1155]), .Z(n12167) );
  NAND U6795 ( .A(n4265), .B(n12167), .Z(n4266) );
  NANDN U6796 ( .A(n9998), .B(n4266), .Z(n4267) );
  AND U6797 ( .A(n6425), .B(n4267), .Z(n4268) );
  NANDN U6798 ( .A(n12166), .B(n4268), .Z(n4269) );
  AND U6799 ( .A(n9999), .B(n4269), .Z(n4270) );
  NAND U6800 ( .A(n4271), .B(n4270), .Z(n4272) );
  NAND U6801 ( .A(n4273), .B(n4272), .Z(n4274) );
  NAND U6802 ( .A(n4275), .B(n4274), .Z(n4276) );
  NANDN U6803 ( .A(x[1160]), .B(y[1160]), .Z(n8205) );
  ANDN U6804 ( .B(y[1161]), .A(x[1161]), .Z(n8210) );
  ANDN U6805 ( .B(n8205), .A(n8210), .Z(n12179) );
  NAND U6806 ( .A(n4276), .B(n12179), .Z(n4277) );
  ANDN U6807 ( .B(x[1162]), .A(y[1162]), .Z(n8213) );
  ANDN U6808 ( .B(n4277), .A(n8213), .Z(n4278) );
  NANDN U6809 ( .A(y[1161]), .B(x[1161]), .Z(n12182) );
  NAND U6810 ( .A(n4278), .B(n12182), .Z(n4279) );
  AND U6811 ( .A(n6421), .B(n4279), .Z(n4280) );
  NANDN U6812 ( .A(x[1162]), .B(y[1162]), .Z(n12183) );
  NAND U6813 ( .A(n4280), .B(n12183), .Z(n4281) );
  NANDN U6814 ( .A(n8214), .B(n4281), .Z(n4282) );
  IV U6815 ( .A(y[1164]), .Z(n6419) );
  OR U6816 ( .A(n4282), .B(n6419), .Z(n4285) );
  XNOR U6817 ( .A(n4282), .B(y[1164]), .Z(n4283) );
  NANDN U6818 ( .A(x[1164]), .B(n4283), .Z(n4284) );
  AND U6819 ( .A(n4285), .B(n4284), .Z(n4287) );
  IV U6820 ( .A(y[1165]), .Z(n8218) );
  OR U6821 ( .A(n4287), .B(n8218), .Z(n4286) );
  AND U6822 ( .A(n8219), .B(n4286), .Z(n4290) );
  XNOR U6823 ( .A(n4287), .B(y[1165]), .Z(n4288) );
  NANDN U6824 ( .A(x[1165]), .B(n4288), .Z(n4289) );
  AND U6825 ( .A(n4290), .B(n4289), .Z(n4293) );
  NANDN U6826 ( .A(y[1166]), .B(x[1166]), .Z(n4292) );
  NANDN U6827 ( .A(y[1167]), .B(x[1167]), .Z(n4291) );
  AND U6828 ( .A(n4292), .B(n4291), .Z(n12193) );
  NANDN U6829 ( .A(n4293), .B(n12193), .Z(n4296) );
  NANDN U6830 ( .A(x[1168]), .B(y[1168]), .Z(n4295) );
  NANDN U6831 ( .A(x[1167]), .B(y[1167]), .Z(n4294) );
  NAND U6832 ( .A(n4295), .B(n4294), .Z(n12196) );
  ANDN U6833 ( .B(n4296), .A(n12196), .Z(n4299) );
  NANDN U6834 ( .A(y[1169]), .B(x[1169]), .Z(n4298) );
  NANDN U6835 ( .A(y[1168]), .B(x[1168]), .Z(n4297) );
  NAND U6836 ( .A(n4298), .B(n4297), .Z(n12198) );
  OR U6837 ( .A(n4299), .B(n12198), .Z(n4300) );
  NANDN U6838 ( .A(n8225), .B(n4300), .Z(n4301) );
  NANDN U6839 ( .A(n4301), .B(x[1170]), .Z(n4304) );
  XNOR U6840 ( .A(n4301), .B(x[1170]), .Z(n4302) );
  NANDN U6841 ( .A(y[1170]), .B(n4302), .Z(n4303) );
  NAND U6842 ( .A(n4304), .B(n4303), .Z(n4305) );
  NANDN U6843 ( .A(n12204), .B(n4305), .Z(n4306) );
  AND U6844 ( .A(n8227), .B(n4306), .Z(n4307) );
  NANDN U6845 ( .A(y[1172]), .B(x[1172]), .Z(n12205) );
  NAND U6846 ( .A(n4307), .B(n12205), .Z(n4308) );
  NANDN U6847 ( .A(n12208), .B(n4308), .Z(n4309) );
  AND U6848 ( .A(n12209), .B(n4309), .Z(n4310) );
  NANDN U6849 ( .A(y[1174]), .B(x[1174]), .Z(n6416) );
  NAND U6850 ( .A(n4310), .B(n6416), .Z(n4311) );
  NANDN U6851 ( .A(x[1174]), .B(y[1174]), .Z(n12211) );
  NAND U6852 ( .A(n4311), .B(n12211), .Z(n4313) );
  NANDN U6853 ( .A(x[1175]), .B(n4313), .Z(n4312) );
  AND U6854 ( .A(n6414), .B(n4312), .Z(n4316) );
  IV U6855 ( .A(y[1175]), .Z(n6412) );
  XNOR U6856 ( .A(n4313), .B(x[1175]), .Z(n4314) );
  NANDN U6857 ( .A(n6412), .B(n4314), .Z(n4315) );
  NAND U6858 ( .A(n4316), .B(n4315), .Z(n4317) );
  NANDN U6859 ( .A(n12217), .B(n4317), .Z(n4320) );
  NANDN U6860 ( .A(x[1177]), .B(y[1177]), .Z(n4319) );
  NANDN U6861 ( .A(x[1178]), .B(y[1178]), .Z(n4318) );
  AND U6862 ( .A(n4319), .B(n4318), .Z(n12219) );
  NAND U6863 ( .A(n4320), .B(n12219), .Z(n4323) );
  NANDN U6864 ( .A(y[1178]), .B(x[1178]), .Z(n4322) );
  NANDN U6865 ( .A(y[1179]), .B(x[1179]), .Z(n4321) );
  NAND U6866 ( .A(n4322), .B(n4321), .Z(n12221) );
  ANDN U6867 ( .B(n4323), .A(n12221), .Z(n4324) );
  NANDN U6868 ( .A(x[1179]), .B(y[1179]), .Z(n12223) );
  NANDN U6869 ( .A(n4324), .B(n12223), .Z(n4325) );
  NANDN U6870 ( .A(y[1180]), .B(x[1180]), .Z(n12225) );
  NAND U6871 ( .A(n4325), .B(n12225), .Z(n4326) );
  NANDN U6872 ( .A(n12228), .B(n4326), .Z(n4330) );
  NANDN U6873 ( .A(y[1182]), .B(x[1182]), .Z(n4328) );
  NAND U6874 ( .A(n4328), .B(n4327), .Z(n8251) );
  NANDN U6875 ( .A(y[1181]), .B(x[1181]), .Z(n4329) );
  NANDN U6876 ( .A(n8251), .B(n4329), .Z(n12230) );
  ANDN U6877 ( .B(n4330), .A(n12230), .Z(n4331) );
  OR U6878 ( .A(n12232), .B(n4331), .Z(n4332) );
  NANDN U6879 ( .A(y[1184]), .B(x[1184]), .Z(n12233) );
  NAND U6880 ( .A(n4332), .B(n12233), .Z(n4333) );
  AND U6881 ( .A(n12235), .B(n4333), .Z(n4334) );
  ANDN U6882 ( .B(n12238), .A(n4334), .Z(n4335) );
  NANDN U6883 ( .A(y[1186]), .B(x[1186]), .Z(n6407) );
  NAND U6884 ( .A(n4335), .B(n6407), .Z(n4336) );
  NANDN U6885 ( .A(n12240), .B(n4336), .Z(n4338) );
  XNOR U6886 ( .A(x[1187]), .B(n4338), .Z(n4337) );
  NANDN U6887 ( .A(y[1187]), .B(n4337), .Z(n4340) );
  NANDN U6888 ( .A(n4338), .B(x[1187]), .Z(n4339) );
  AND U6889 ( .A(n4340), .B(n4339), .Z(n4341) );
  NAND U6890 ( .A(n4342), .B(n4341), .Z(n4343) );
  NAND U6891 ( .A(n6404), .B(n4343), .Z(n4344) );
  AND U6892 ( .A(n8264), .B(n4344), .Z(n4347) );
  NANDN U6893 ( .A(x[1189]), .B(y[1189]), .Z(n4346) );
  NANDN U6894 ( .A(x[1190]), .B(y[1190]), .Z(n4345) );
  AND U6895 ( .A(n4346), .B(n4345), .Z(n12247) );
  NANDN U6896 ( .A(n4347), .B(n12247), .Z(n4350) );
  NANDN U6897 ( .A(y[1191]), .B(x[1191]), .Z(n4349) );
  NANDN U6898 ( .A(y[1190]), .B(x[1190]), .Z(n4348) );
  NAND U6899 ( .A(n4349), .B(n4348), .Z(n12250) );
  ANDN U6900 ( .B(n4350), .A(n12250), .Z(n4353) );
  NANDN U6901 ( .A(x[1191]), .B(y[1191]), .Z(n4352) );
  NANDN U6902 ( .A(x[1192]), .B(y[1192]), .Z(n4351) );
  AND U6903 ( .A(n4352), .B(n4351), .Z(n12251) );
  NANDN U6904 ( .A(n4353), .B(n12251), .Z(n4354) );
  NANDN U6905 ( .A(n12253), .B(n4354), .Z(n4355) );
  NANDN U6906 ( .A(x[1193]), .B(y[1193]), .Z(n8272) );
  NAND U6907 ( .A(n4355), .B(n8272), .Z(n4357) );
  NANDN U6908 ( .A(x[1194]), .B(n4357), .Z(n4356) );
  AND U6909 ( .A(n12259), .B(n4356), .Z(n4360) );
  XNOR U6910 ( .A(x[1194]), .B(n4357), .Z(n4358) );
  NAND U6911 ( .A(n4358), .B(y[1194]), .Z(n4359) );
  NAND U6912 ( .A(n4360), .B(n4359), .Z(n4361) );
  NAND U6913 ( .A(n4362), .B(n4361), .Z(n4363) );
  NANDN U6914 ( .A(x[1196]), .B(y[1196]), .Z(n8277) );
  ANDN U6915 ( .B(y[1197]), .A(x[1197]), .Z(n8284) );
  ANDN U6916 ( .B(n8277), .A(n8284), .Z(n12263) );
  NAND U6917 ( .A(n4363), .B(n12263), .Z(n4364) );
  AND U6918 ( .A(n8285), .B(n4364), .Z(n4365) );
  NANDN U6919 ( .A(y[1197]), .B(x[1197]), .Z(n12265) );
  NAND U6920 ( .A(n4365), .B(n12265), .Z(n4366) );
  NANDN U6921 ( .A(n12268), .B(n4366), .Z(n4369) );
  ANDN U6922 ( .B(x[1199]), .A(y[1199]), .Z(n8286) );
  NAND U6923 ( .A(n4367), .B(n8286), .Z(n4368) );
  NAND U6924 ( .A(n4369), .B(n4368), .Z(n4372) );
  NANDN U6925 ( .A(y[1200]), .B(x[1200]), .Z(n4371) );
  NANDN U6926 ( .A(y[1201]), .B(x[1201]), .Z(n4370) );
  NAND U6927 ( .A(n4371), .B(n4370), .Z(n8289) );
  OR U6928 ( .A(n4372), .B(n8289), .Z(n4373) );
  NANDN U6929 ( .A(n12272), .B(n4373), .Z(n4376) );
  NANDN U6930 ( .A(y[1202]), .B(x[1202]), .Z(n4375) );
  NANDN U6931 ( .A(y[1203]), .B(x[1203]), .Z(n4374) );
  AND U6932 ( .A(n4375), .B(n4374), .Z(n12273) );
  NAND U6933 ( .A(n4376), .B(n12273), .Z(n4377) );
  NANDN U6934 ( .A(n12276), .B(n4377), .Z(n4378) );
  AND U6935 ( .A(n6403), .B(n4378), .Z(n4379) );
  NAND U6936 ( .A(n4379), .B(n12277), .Z(n4380) );
  NAND U6937 ( .A(n4381), .B(n4380), .Z(n4382) );
  NANDN U6938 ( .A(y[1207]), .B(x[1207]), .Z(n6402) );
  NAND U6939 ( .A(n4382), .B(n6402), .Z(n4383) );
  NANDN U6940 ( .A(y[1208]), .B(x[1208]), .Z(n12285) );
  NANDN U6941 ( .A(n4383), .B(n12285), .Z(n4384) );
  ANDN U6942 ( .B(y[1208]), .A(x[1208]), .Z(n8300) );
  ANDN U6943 ( .B(y[1209]), .A(x[1209]), .Z(n6401) );
  NOR U6944 ( .A(n8300), .B(n6401), .Z(n12287) );
  NAND U6945 ( .A(n4384), .B(n12287), .Z(n4385) );
  NANDN U6946 ( .A(y[1209]), .B(x[1209]), .Z(n12289) );
  NAND U6947 ( .A(n4385), .B(n12289), .Z(n4386) );
  NANDN U6948 ( .A(x[1210]), .B(y[1210]), .Z(n12292) );
  NAND U6949 ( .A(n4386), .B(n12292), .Z(n4389) );
  NANDN U6950 ( .A(y[1210]), .B(x[1210]), .Z(n4388) );
  NANDN U6951 ( .A(y[1211]), .B(x[1211]), .Z(n4387) );
  AND U6952 ( .A(n4388), .B(n4387), .Z(n12293) );
  NAND U6953 ( .A(n4389), .B(n12293), .Z(n4392) );
  NANDN U6954 ( .A(x[1212]), .B(y[1212]), .Z(n4391) );
  NANDN U6955 ( .A(x[1211]), .B(y[1211]), .Z(n4390) );
  NAND U6956 ( .A(n4391), .B(n4390), .Z(n12295) );
  ANDN U6957 ( .B(n4392), .A(n12295), .Z(n4395) );
  NANDN U6958 ( .A(y[1212]), .B(x[1212]), .Z(n4394) );
  NANDN U6959 ( .A(y[1213]), .B(x[1213]), .Z(n4393) );
  AND U6960 ( .A(n4394), .B(n4393), .Z(n12297) );
  NANDN U6961 ( .A(n4395), .B(n12297), .Z(n4398) );
  NANDN U6962 ( .A(x[1214]), .B(y[1214]), .Z(n4397) );
  NANDN U6963 ( .A(x[1213]), .B(y[1213]), .Z(n4396) );
  NAND U6964 ( .A(n4397), .B(n4396), .Z(n12300) );
  ANDN U6965 ( .B(n4398), .A(n12300), .Z(n4401) );
  NANDN U6966 ( .A(y[1214]), .B(x[1214]), .Z(n4400) );
  NANDN U6967 ( .A(y[1215]), .B(x[1215]), .Z(n4399) );
  AND U6968 ( .A(n4400), .B(n4399), .Z(n12301) );
  NANDN U6969 ( .A(n4401), .B(n12301), .Z(n4404) );
  NANDN U6970 ( .A(x[1216]), .B(y[1216]), .Z(n4403) );
  NANDN U6971 ( .A(x[1215]), .B(y[1215]), .Z(n4402) );
  NAND U6972 ( .A(n4403), .B(n4402), .Z(n12304) );
  ANDN U6973 ( .B(n4404), .A(n12304), .Z(n4407) );
  NANDN U6974 ( .A(y[1216]), .B(x[1216]), .Z(n4406) );
  NANDN U6975 ( .A(y[1217]), .B(x[1217]), .Z(n4405) );
  AND U6976 ( .A(n4406), .B(n4405), .Z(n12305) );
  NANDN U6977 ( .A(n4407), .B(n12305), .Z(n4408) );
  NANDN U6978 ( .A(n12307), .B(n4408), .Z(n4411) );
  NANDN U6979 ( .A(y[1219]), .B(x[1219]), .Z(n4410) );
  NANDN U6980 ( .A(y[1218]), .B(x[1218]), .Z(n4409) );
  AND U6981 ( .A(n4410), .B(n4409), .Z(n12309) );
  NAND U6982 ( .A(n4411), .B(n12309), .Z(n4412) );
  NANDN U6983 ( .A(x[1219]), .B(y[1219]), .Z(n12311) );
  NAND U6984 ( .A(n4412), .B(n12311), .Z(n4413) );
  NANDN U6985 ( .A(y[1220]), .B(x[1220]), .Z(n6399) );
  NAND U6986 ( .A(n4413), .B(n6399), .Z(n4414) );
  ANDN U6987 ( .B(y[1220]), .A(x[1220]), .Z(n6400) );
  NANDN U6988 ( .A(x[1221]), .B(y[1221]), .Z(n6398) );
  NANDN U6989 ( .A(n6400), .B(n6398), .Z(n12315) );
  ANDN U6990 ( .B(n4414), .A(n12315), .Z(n4415) );
  ANDN U6991 ( .B(n12316), .A(n4415), .Z(n4416) );
  NANDN U6992 ( .A(y[1222]), .B(x[1222]), .Z(n6397) );
  NAND U6993 ( .A(n4416), .B(n6397), .Z(n4417) );
  NANDN U6994 ( .A(n12314), .B(n4417), .Z(n4418) );
  NANDN U6995 ( .A(n4418), .B(x[1223]), .Z(n4421) );
  XNOR U6996 ( .A(n4418), .B(x[1223]), .Z(n4419) );
  NANDN U6997 ( .A(y[1223]), .B(n4419), .Z(n4420) );
  AND U6998 ( .A(n4421), .B(n4420), .Z(n4422) );
  OR U6999 ( .A(n4422), .B(y[1224]), .Z(n4425) );
  XOR U7000 ( .A(y[1224]), .B(n4422), .Z(n4423) );
  NAND U7001 ( .A(n4423), .B(x[1224]), .Z(n4424) );
  NAND U7002 ( .A(n4425), .B(n4424), .Z(n4426) );
  AND U7003 ( .A(n12320), .B(n4426), .Z(n4432) );
  NANDN U7004 ( .A(y[1226]), .B(x[1226]), .Z(n4428) );
  NANDN U7005 ( .A(y[1227]), .B(x[1227]), .Z(n4427) );
  AND U7006 ( .A(n4428), .B(n4427), .Z(n12321) );
  ANDN U7007 ( .B(x[1225]), .A(y[1225]), .Z(n8321) );
  NANDN U7008 ( .A(n4429), .B(n8321), .Z(n4430) );
  AND U7009 ( .A(n12321), .B(n4430), .Z(n4431) );
  NANDN U7010 ( .A(n4432), .B(n4431), .Z(n4435) );
  NANDN U7011 ( .A(x[1228]), .B(y[1228]), .Z(n4434) );
  NANDN U7012 ( .A(x[1227]), .B(y[1227]), .Z(n4433) );
  NAND U7013 ( .A(n4434), .B(n4433), .Z(n12322) );
  ANDN U7014 ( .B(n4435), .A(n12322), .Z(n4438) );
  NANDN U7015 ( .A(y[1228]), .B(x[1228]), .Z(n4437) );
  NANDN U7016 ( .A(y[1229]), .B(x[1229]), .Z(n4436) );
  AND U7017 ( .A(n4437), .B(n4436), .Z(n12323) );
  NANDN U7018 ( .A(n4438), .B(n12323), .Z(n4439) );
  NANDN U7019 ( .A(n8328), .B(n4439), .Z(n4440) );
  NANDN U7020 ( .A(y[1230]), .B(x[1230]), .Z(n8332) );
  NAND U7021 ( .A(n4440), .B(n8332), .Z(n4441) );
  NAND U7022 ( .A(n4442), .B(n4441), .Z(n4444) );
  NANDN U7023 ( .A(y[1232]), .B(x[1232]), .Z(n12327) );
  ANDN U7024 ( .B(x[1231]), .A(y[1231]), .Z(n8331) );
  ANDN U7025 ( .B(n12327), .A(n8331), .Z(n4443) );
  NAND U7026 ( .A(n4444), .B(n4443), .Z(n4445) );
  ANDN U7027 ( .B(y[1232]), .A(x[1232]), .Z(n8336) );
  ANDN U7028 ( .B(y[1233]), .A(x[1233]), .Z(n6395) );
  NOR U7029 ( .A(n8336), .B(n6395), .Z(n12328) );
  NAND U7030 ( .A(n4445), .B(n12328), .Z(n4446) );
  NAND U7031 ( .A(n4447), .B(n4446), .Z(n4448) );
  NANDN U7032 ( .A(x[1234]), .B(y[1234]), .Z(n12330) );
  NAND U7033 ( .A(n4448), .B(n12330), .Z(n4449) );
  NAND U7034 ( .A(n4450), .B(n4449), .Z(n4451) );
  NAND U7035 ( .A(n6394), .B(n4451), .Z(n4452) );
  NAND U7036 ( .A(n4453), .B(n4452), .Z(n4454) );
  NAND U7037 ( .A(n4455), .B(n4454), .Z(n4456) );
  ANDN U7038 ( .B(x[1237]), .A(y[1237]), .Z(n8344) );
  ANDN U7039 ( .B(n4456), .A(n8344), .Z(n4457) );
  ANDN U7040 ( .B(y[1237]), .A(x[1237]), .Z(n12338) );
  ANDN U7041 ( .B(y[1238]), .A(x[1238]), .Z(n12343) );
  NOR U7042 ( .A(n12338), .B(n12343), .Z(n8347) );
  NANDN U7043 ( .A(n4457), .B(n8347), .Z(n4458) );
  NANDN U7044 ( .A(n12339), .B(n4458), .Z(n4460) );
  NANDN U7045 ( .A(x[1239]), .B(y[1239]), .Z(n12342) );
  ANDN U7046 ( .B(n12342), .A(n12350), .Z(n8350) );
  NAND U7047 ( .A(n4460), .B(n8350), .Z(n4461) );
  NAND U7048 ( .A(n4462), .B(n4461), .Z(n4463) );
  NANDN U7049 ( .A(x[1242]), .B(y[1242]), .Z(n12353) );
  NAND U7050 ( .A(n4463), .B(n12353), .Z(n4464) );
  NANDN U7051 ( .A(x[1243]), .B(y[1243]), .Z(n12357) );
  NANDN U7052 ( .A(n4464), .B(n12357), .Z(n4465) );
  AND U7053 ( .A(n12359), .B(n4465), .Z(n4466) );
  NANDN U7054 ( .A(n8356), .B(n4466), .Z(n4467) );
  ANDN U7055 ( .B(y[1245]), .A(x[1245]), .Z(n8363) );
  ANDN U7056 ( .B(y[1244]), .A(x[1244]), .Z(n8358) );
  NOR U7057 ( .A(n8363), .B(n8358), .Z(n12361) );
  NAND U7058 ( .A(n4467), .B(n12361), .Z(n4468) );
  ANDN U7059 ( .B(x[1246]), .A(y[1246]), .Z(n8366) );
  ANDN U7060 ( .B(n4468), .A(n8366), .Z(n4469) );
  NANDN U7061 ( .A(y[1245]), .B(x[1245]), .Z(n12364) );
  NAND U7062 ( .A(n4469), .B(n12364), .Z(n4470) );
  AND U7063 ( .A(n6390), .B(n4470), .Z(n4471) );
  NANDN U7064 ( .A(x[1246]), .B(y[1246]), .Z(n12365) );
  NAND U7065 ( .A(n4471), .B(n12365), .Z(n4472) );
  ANDN U7066 ( .B(x[1247]), .A(y[1247]), .Z(n8367) );
  ANDN U7067 ( .B(n4472), .A(n8367), .Z(n4473) );
  NAND U7068 ( .A(n4474), .B(n4473), .Z(n4475) );
  NAND U7069 ( .A(n4476), .B(n4475), .Z(n4477) );
  AND U7070 ( .A(n6385), .B(n4477), .Z(n4478) );
  OR U7071 ( .A(n12372), .B(n4478), .Z(n4479) );
  AND U7072 ( .A(n12373), .B(n4479), .Z(n4480) );
  NANDN U7073 ( .A(x[1251]), .B(y[1251]), .Z(n12374) );
  NANDN U7074 ( .A(n4480), .B(n12374), .Z(n4481) );
  NANDN U7075 ( .A(y[1252]), .B(x[1252]), .Z(n12375) );
  NAND U7076 ( .A(n4481), .B(n12375), .Z(n4482) );
  ANDN U7077 ( .B(y[1253]), .A(x[1253]), .Z(n8381) );
  ANDN U7078 ( .B(y[1252]), .A(x[1252]), .Z(n8375) );
  NOR U7079 ( .A(n8381), .B(n8375), .Z(n12376) );
  NAND U7080 ( .A(n4482), .B(n12376), .Z(n4483) );
  NAND U7081 ( .A(n4484), .B(n4483), .Z(n4485) );
  ANDN U7082 ( .B(y[1254]), .A(x[1254]), .Z(n8378) );
  ANDN U7083 ( .B(y[1255]), .A(x[1255]), .Z(n12381) );
  NOR U7084 ( .A(n8378), .B(n12381), .Z(n12378) );
  NAND U7085 ( .A(n4485), .B(n12378), .Z(n4486) );
  NAND U7086 ( .A(n4487), .B(n4486), .Z(n4488) );
  ANDN U7087 ( .B(y[1257]), .A(x[1257]), .Z(n6382) );
  ANDN U7088 ( .B(y[1256]), .A(x[1256]), .Z(n8385) );
  NOR U7089 ( .A(n6382), .B(n8385), .Z(n12382) );
  NAND U7090 ( .A(n4488), .B(n12382), .Z(n4489) );
  NAND U7091 ( .A(n4490), .B(n4489), .Z(n4493) );
  ANDN U7092 ( .B(y[1260]), .A(x[1260]), .Z(n4494) );
  NANDN U7093 ( .A(x[1259]), .B(y[1259]), .Z(n4491) );
  NANDN U7094 ( .A(n4494), .B(n4491), .Z(n8393) );
  NANDN U7095 ( .A(x[1258]), .B(y[1258]), .Z(n4492) );
  NANDN U7096 ( .A(n8393), .B(n4492), .Z(n12384) );
  ANDN U7097 ( .B(n4493), .A(n12384), .Z(n4499) );
  ANDN U7098 ( .B(x[1259]), .A(y[1259]), .Z(n8391) );
  NANDN U7099 ( .A(n4494), .B(n8391), .Z(n4497) );
  NANDN U7100 ( .A(y[1260]), .B(x[1260]), .Z(n4496) );
  NANDN U7101 ( .A(y[1261]), .B(x[1261]), .Z(n4495) );
  NAND U7102 ( .A(n4496), .B(n4495), .Z(n8394) );
  ANDN U7103 ( .B(n4497), .A(n8394), .Z(n4498) );
  NANDN U7104 ( .A(n4499), .B(n4498), .Z(n4504) );
  NANDN U7105 ( .A(x[1262]), .B(y[1262]), .Z(n4501) );
  NANDN U7106 ( .A(x[1261]), .B(y[1261]), .Z(n4500) );
  AND U7107 ( .A(n4501), .B(n4500), .Z(n4503) );
  NANDN U7108 ( .A(x[1263]), .B(y[1263]), .Z(n4502) );
  NAND U7109 ( .A(n4503), .B(n4502), .Z(n12386) );
  ANDN U7110 ( .B(n4504), .A(n12386), .Z(n4513) );
  NANDN U7111 ( .A(y[1265]), .B(x[1265]), .Z(n4506) );
  NANDN U7112 ( .A(y[1264]), .B(x[1264]), .Z(n4505) );
  AND U7113 ( .A(n4506), .B(n4505), .Z(n4512) );
  NANDN U7114 ( .A(y[1262]), .B(x[1262]), .Z(n4507) );
  NANDN U7115 ( .A(x[1263]), .B(n4507), .Z(n4510) );
  XNOR U7116 ( .A(n4507), .B(x[1263]), .Z(n4508) );
  NAND U7117 ( .A(n4508), .B(y[1263]), .Z(n4509) );
  NAND U7118 ( .A(n4510), .B(n4509), .Z(n4511) );
  NAND U7119 ( .A(n4512), .B(n4511), .Z(n12387) );
  OR U7120 ( .A(n4513), .B(n12387), .Z(n4514) );
  NANDN U7121 ( .A(n12388), .B(n4514), .Z(n4521) );
  XNOR U7122 ( .A(x[1267]), .B(y[1267]), .Z(n4516) );
  NANDN U7123 ( .A(y[1266]), .B(x[1266]), .Z(n4515) );
  NAND U7124 ( .A(n4516), .B(n4515), .Z(n4517) );
  NAND U7125 ( .A(n4518), .B(n4517), .Z(n4520) );
  NANDN U7126 ( .A(y[1268]), .B(x[1268]), .Z(n4519) );
  NAND U7127 ( .A(n4520), .B(n4519), .Z(n8400) );
  ANDN U7128 ( .B(n4521), .A(n8400), .Z(n4524) );
  NANDN U7129 ( .A(x[1269]), .B(y[1269]), .Z(n4523) );
  NANDN U7130 ( .A(x[1268]), .B(y[1268]), .Z(n4522) );
  NAND U7131 ( .A(n4523), .B(n4522), .Z(n6378) );
  OR U7132 ( .A(n4524), .B(n6378), .Z(n4525) );
  NANDN U7133 ( .A(n6379), .B(n4525), .Z(n4526) );
  IV U7134 ( .A(y[1270]), .Z(n6377) );
  OR U7135 ( .A(n4526), .B(n6377), .Z(n4529) );
  XNOR U7136 ( .A(n4526), .B(y[1270]), .Z(n4527) );
  NANDN U7137 ( .A(x[1270]), .B(n4527), .Z(n4528) );
  AND U7138 ( .A(n4529), .B(n4528), .Z(n4531) );
  NANDN U7139 ( .A(y[1271]), .B(n4531), .Z(n4530) );
  AND U7140 ( .A(n6374), .B(n4530), .Z(n4534) );
  IV U7141 ( .A(y[1271]), .Z(n8405) );
  XOR U7142 ( .A(n4531), .B(n8405), .Z(n4532) );
  NAND U7143 ( .A(n4532), .B(x[1271]), .Z(n4533) );
  NAND U7144 ( .A(n4534), .B(n4533), .Z(n4535) );
  NANDN U7145 ( .A(x[1272]), .B(y[1272]), .Z(n8406) );
  AND U7146 ( .A(n4535), .B(n8406), .Z(n4536) );
  NAND U7147 ( .A(n4537), .B(n4536), .Z(n4538) );
  NAND U7148 ( .A(n4539), .B(n4538), .Z(n4540) );
  NANDN U7149 ( .A(n8410), .B(n4540), .Z(n4542) );
  NANDN U7150 ( .A(n8414), .B(n4542), .Z(n4541) );
  AND U7151 ( .A(n8416), .B(n4541), .Z(n4545) );
  XOR U7152 ( .A(y[1275]), .B(n4542), .Z(n4543) );
  NANDN U7153 ( .A(x[1275]), .B(n4543), .Z(n4544) );
  NAND U7154 ( .A(n4545), .B(n4544), .Z(n4548) );
  NANDN U7155 ( .A(y[1276]), .B(x[1276]), .Z(n4547) );
  NANDN U7156 ( .A(y[1277]), .B(x[1277]), .Z(n4546) );
  AND U7157 ( .A(n4547), .B(n4546), .Z(n12405) );
  NAND U7158 ( .A(n4548), .B(n12405), .Z(n4551) );
  ANDN U7159 ( .B(y[1279]), .A(x[1279]), .Z(n8423) );
  NANDN U7160 ( .A(x[1278]), .B(y[1278]), .Z(n4550) );
  NANDN U7161 ( .A(x[1277]), .B(y[1277]), .Z(n4549) );
  NAND U7162 ( .A(n4550), .B(n4549), .Z(n8419) );
  NOR U7163 ( .A(n8423), .B(n8419), .Z(n12408) );
  NAND U7164 ( .A(n4551), .B(n12408), .Z(n4555) );
  NANDN U7165 ( .A(y[1280]), .B(x[1280]), .Z(n6368) );
  NANDN U7166 ( .A(y[1278]), .B(x[1278]), .Z(n4553) );
  NANDN U7167 ( .A(y[1279]), .B(x[1279]), .Z(n4552) );
  NAND U7168 ( .A(n4553), .B(n4552), .Z(n8422) );
  NANDN U7169 ( .A(n8423), .B(n8422), .Z(n4554) );
  NAND U7170 ( .A(n6368), .B(n4554), .Z(n12409) );
  ANDN U7171 ( .B(n4555), .A(n12409), .Z(n4557) );
  NANDN U7172 ( .A(x[1280]), .B(y[1280]), .Z(n4556) );
  ANDN U7173 ( .B(y[1281]), .A(x[1281]), .Z(n8429) );
  ANDN U7174 ( .B(n4556), .A(n8429), .Z(n12412) );
  NANDN U7175 ( .A(n4557), .B(n12412), .Z(n4558) );
  ANDN U7176 ( .B(x[1282]), .A(y[1282]), .Z(n8432) );
  ANDN U7177 ( .B(n4558), .A(n8432), .Z(n4559) );
  NANDN U7178 ( .A(y[1281]), .B(x[1281]), .Z(n12413) );
  NAND U7179 ( .A(n4559), .B(n12413), .Z(n4560) );
  AND U7180 ( .A(n8436), .B(n4560), .Z(n4561) );
  NANDN U7181 ( .A(x[1282]), .B(y[1282]), .Z(n12415) );
  NAND U7182 ( .A(n4561), .B(n12415), .Z(n4562) );
  NANDN U7183 ( .A(n8433), .B(n4562), .Z(n4566) );
  OR U7184 ( .A(n4566), .B(x[1284]), .Z(n4565) );
  NANDN U7185 ( .A(x[1285]), .B(y[1285]), .Z(n4563) );
  NAND U7186 ( .A(n4564), .B(n4563), .Z(n12424) );
  ANDN U7187 ( .B(n4565), .A(n12424), .Z(n4569) );
  XOR U7188 ( .A(n4566), .B(x[1284]), .Z(n4567) );
  NAND U7189 ( .A(n4567), .B(y[1284]), .Z(n4568) );
  NAND U7190 ( .A(n4569), .B(n4568), .Z(n4570) );
  AND U7191 ( .A(n12425), .B(n4570), .Z(n4571) );
  NAND U7192 ( .A(n4572), .B(n4571), .Z(n4573) );
  NANDN U7193 ( .A(n12427), .B(n4573), .Z(n4576) );
  NANDN U7194 ( .A(y[1288]), .B(x[1288]), .Z(n4575) );
  NANDN U7195 ( .A(y[1289]), .B(x[1289]), .Z(n4574) );
  AND U7196 ( .A(n4575), .B(n4574), .Z(n12429) );
  NAND U7197 ( .A(n4576), .B(n12429), .Z(n4577) );
  AND U7198 ( .A(n6364), .B(n4577), .Z(n4578) );
  NAND U7199 ( .A(n4579), .B(n4578), .Z(n4580) );
  NAND U7200 ( .A(n8445), .B(n4580), .Z(n4581) );
  AND U7201 ( .A(n12436), .B(n4581), .Z(n4583) );
  ANDN U7202 ( .B(x[1291]), .A(y[1291]), .Z(n8444) );
  ANDN U7203 ( .B(x[1292]), .A(y[1292]), .Z(n12438) );
  OR U7204 ( .A(n8444), .B(n12438), .Z(n4582) );
  OR U7205 ( .A(n4583), .B(n4582), .Z(n4584) );
  NANDN U7206 ( .A(x[1292]), .B(y[1292]), .Z(n8447) );
  NANDN U7207 ( .A(x[1293]), .B(y[1293]), .Z(n8452) );
  NAND U7208 ( .A(n8447), .B(n8452), .Z(n12440) );
  ANDN U7209 ( .B(n4584), .A(n12440), .Z(n4585) );
  ANDN U7210 ( .B(n12441), .A(n4585), .Z(n4586) );
  NANDN U7211 ( .A(y[1294]), .B(x[1294]), .Z(n6363) );
  NAND U7212 ( .A(n4586), .B(n6363), .Z(n4587) );
  AND U7213 ( .A(n12443), .B(n4587), .Z(n4588) );
  NAND U7214 ( .A(n4589), .B(n4588), .Z(n4590) );
  NAND U7215 ( .A(n4591), .B(n4590), .Z(n4592) );
  ANDN U7216 ( .B(y[1296]), .A(x[1296]), .Z(n8456) );
  ANDN U7217 ( .B(n4592), .A(n8456), .Z(n4593) );
  NAND U7218 ( .A(n4594), .B(n4593), .Z(n4595) );
  NAND U7219 ( .A(n8459), .B(n4595), .Z(n4596) );
  AND U7220 ( .A(n6360), .B(n4596), .Z(n4599) );
  NANDN U7221 ( .A(y[1298]), .B(x[1298]), .Z(n4598) );
  NANDN U7222 ( .A(y[1299]), .B(x[1299]), .Z(n4597) );
  AND U7223 ( .A(n4598), .B(n4597), .Z(n12453) );
  NANDN U7224 ( .A(n4599), .B(n12453), .Z(n4600) );
  NANDN U7225 ( .A(n12456), .B(n4600), .Z(n4601) );
  NANDN U7226 ( .A(y[1302]), .B(x[1302]), .Z(n8468) );
  NAND U7227 ( .A(n4601), .B(n8468), .Z(n4606) );
  NANDN U7228 ( .A(y[1300]), .B(x[1300]), .Z(n4602) );
  NANDN U7229 ( .A(n4602), .B(x[1301]), .Z(n4605) );
  XNOR U7230 ( .A(n4602), .B(x[1301]), .Z(n4603) );
  NANDN U7231 ( .A(y[1301]), .B(n4603), .Z(n4604) );
  AND U7232 ( .A(n4605), .B(n4604), .Z(n12458) );
  NANDN U7233 ( .A(n4606), .B(n12458), .Z(n4607) );
  AND U7234 ( .A(n12459), .B(n4607), .Z(n4608) );
  NANDN U7235 ( .A(x[1303]), .B(y[1303]), .Z(n12463) );
  NAND U7236 ( .A(n4608), .B(n12463), .Z(n4609) );
  AND U7237 ( .A(n4610), .B(n4609), .Z(n4611) );
  ANDN U7238 ( .B(y[1305]), .A(x[1305]), .Z(n6359) );
  ANDN U7239 ( .B(y[1304]), .A(x[1304]), .Z(n8472) );
  NOR U7240 ( .A(n6359), .B(n8472), .Z(n12467) );
  NANDN U7241 ( .A(n4611), .B(n12467), .Z(n4612) );
  ANDN U7242 ( .B(x[1306]), .A(y[1306]), .Z(n8477) );
  ANDN U7243 ( .B(n4612), .A(n8477), .Z(n4613) );
  NANDN U7244 ( .A(y[1305]), .B(x[1305]), .Z(n12469) );
  NAND U7245 ( .A(n4613), .B(n12469), .Z(n4614) );
  AND U7246 ( .A(n12471), .B(n4614), .Z(n4615) );
  NAND U7247 ( .A(n4616), .B(n4615), .Z(n4617) );
  NAND U7248 ( .A(n4618), .B(n4617), .Z(n4619) );
  ANDN U7249 ( .B(y[1308]), .A(x[1308]), .Z(n8480) );
  ANDN U7250 ( .B(n4619), .A(n8480), .Z(n4620) );
  NAND U7251 ( .A(n4621), .B(n4620), .Z(n4622) );
  NAND U7252 ( .A(n4623), .B(n4622), .Z(n4624) );
  ANDN U7253 ( .B(y[1310]), .A(x[1310]), .Z(n8484) );
  ANDN U7254 ( .B(n4624), .A(n8484), .Z(n4627) );
  NANDN U7255 ( .A(y[1310]), .B(x[1310]), .Z(n4626) );
  NANDN U7256 ( .A(y[1311]), .B(x[1311]), .Z(n4625) );
  AND U7257 ( .A(n4626), .B(n4625), .Z(n12481) );
  NANDN U7258 ( .A(n4627), .B(n12481), .Z(n4630) );
  NANDN U7259 ( .A(x[1312]), .B(y[1312]), .Z(n4629) );
  NANDN U7260 ( .A(x[1311]), .B(y[1311]), .Z(n4628) );
  NAND U7261 ( .A(n4629), .B(n4628), .Z(n12484) );
  ANDN U7262 ( .B(n4630), .A(n12484), .Z(n4633) );
  NANDN U7263 ( .A(y[1312]), .B(x[1312]), .Z(n4632) );
  NANDN U7264 ( .A(y[1313]), .B(x[1313]), .Z(n4631) );
  AND U7265 ( .A(n4632), .B(n4631), .Z(n12486) );
  NANDN U7266 ( .A(n4633), .B(n12486), .Z(n4634) );
  NANDN U7267 ( .A(n12488), .B(n4634), .Z(n4635) );
  ANDN U7268 ( .B(x[1314]), .A(y[1314]), .Z(n8491) );
  ANDN U7269 ( .B(n4635), .A(n8491), .Z(n4636) );
  NANDN U7270 ( .A(x[1315]), .B(y[1315]), .Z(n12491) );
  NANDN U7271 ( .A(n4636), .B(n12491), .Z(n4637) );
  ANDN U7272 ( .B(x[1315]), .A(y[1315]), .Z(n8492) );
  ANDN U7273 ( .B(n4637), .A(n8492), .Z(n4638) );
  NANDN U7274 ( .A(y[1316]), .B(x[1316]), .Z(n12493) );
  NAND U7275 ( .A(n4638), .B(n12493), .Z(n4639) );
  AND U7276 ( .A(n12495), .B(n4639), .Z(n4640) );
  ANDN U7277 ( .B(n12498), .A(n4640), .Z(n4641) );
  NANDN U7278 ( .A(y[1318]), .B(x[1318]), .Z(n6353) );
  NAND U7279 ( .A(n4641), .B(n6353), .Z(n4642) );
  NANDN U7280 ( .A(n12500), .B(n4642), .Z(n4643) );
  IV U7281 ( .A(x[1319]), .Z(n6351) );
  OR U7282 ( .A(n4643), .B(n6351), .Z(n4646) );
  XNOR U7283 ( .A(n4643), .B(x[1319]), .Z(n4644) );
  NANDN U7284 ( .A(y[1319]), .B(n4644), .Z(n4645) );
  AND U7285 ( .A(n4646), .B(n4645), .Z(n4648) );
  OR U7286 ( .A(n4648), .B(y[1320]), .Z(n4647) );
  AND U7287 ( .A(n8504), .B(n4647), .Z(n4651) );
  XOR U7288 ( .A(n4648), .B(y[1320]), .Z(n4649) );
  NAND U7289 ( .A(n4649), .B(x[1320]), .Z(n4650) );
  NAND U7290 ( .A(n4651), .B(n4650), .Z(n4654) );
  NANDN U7291 ( .A(x[1322]), .B(y[1322]), .Z(n4653) );
  NANDN U7292 ( .A(x[1321]), .B(y[1321]), .Z(n4652) );
  NAND U7293 ( .A(n4653), .B(n4652), .Z(n12507) );
  ANDN U7294 ( .B(n4654), .A(n12507), .Z(n4657) );
  NANDN U7295 ( .A(y[1322]), .B(x[1322]), .Z(n4656) );
  NANDN U7296 ( .A(y[1323]), .B(x[1323]), .Z(n4655) );
  AND U7297 ( .A(n4656), .B(n4655), .Z(n12509) );
  NANDN U7298 ( .A(n4657), .B(n12509), .Z(n4658) );
  NANDN U7299 ( .A(n12511), .B(n4658), .Z(n4661) );
  NANDN U7300 ( .A(y[1324]), .B(x[1324]), .Z(n4660) );
  NANDN U7301 ( .A(y[1325]), .B(x[1325]), .Z(n4659) );
  AND U7302 ( .A(n4660), .B(n4659), .Z(n12513) );
  NAND U7303 ( .A(n4661), .B(n12513), .Z(n4662) );
  NANDN U7304 ( .A(n12515), .B(n4662), .Z(n4663) );
  NANDN U7305 ( .A(n12518), .B(n4663), .Z(n4664) );
  ANDN U7306 ( .B(y[1327]), .A(x[1327]), .Z(n12520) );
  ANDN U7307 ( .B(n4664), .A(n12520), .Z(n4665) );
  NANDN U7308 ( .A(y[1328]), .B(x[1328]), .Z(n12521) );
  NANDN U7309 ( .A(n4665), .B(n12521), .Z(n4666) );
  NANDN U7310 ( .A(x[1328]), .B(y[1328]), .Z(n6348) );
  NANDN U7311 ( .A(x[1329]), .B(y[1329]), .Z(n8517) );
  NAND U7312 ( .A(n6348), .B(n8517), .Z(n12524) );
  ANDN U7313 ( .B(n4666), .A(n12524), .Z(n4668) );
  NANDN U7314 ( .A(y[1329]), .B(x[1329]), .Z(n12525) );
  NANDN U7315 ( .A(y[1330]), .B(x[1330]), .Z(n8519) );
  AND U7316 ( .A(n12525), .B(n8519), .Z(n4667) );
  NANDN U7317 ( .A(n4668), .B(n4667), .Z(n4672) );
  NANDN U7318 ( .A(x[1330]), .B(y[1330]), .Z(n4671) );
  NANDN U7319 ( .A(x[1331]), .B(y[1331]), .Z(n4669) );
  NAND U7320 ( .A(n4670), .B(n4669), .Z(n8522) );
  ANDN U7321 ( .B(n4671), .A(n8522), .Z(n12528) );
  NAND U7322 ( .A(n4672), .B(n12528), .Z(n4675) );
  NANDN U7323 ( .A(y[1332]), .B(x[1332]), .Z(n4674) );
  NANDN U7324 ( .A(y[1333]), .B(x[1333]), .Z(n4673) );
  NAND U7325 ( .A(n4674), .B(n4673), .Z(n8523) );
  ANDN U7326 ( .B(n4675), .A(n8523), .Z(n4676) );
  NAND U7327 ( .A(n4677), .B(n4676), .Z(n4678) );
  NANDN U7328 ( .A(n12531), .B(n4678), .Z(n4681) );
  NANDN U7329 ( .A(y[1334]), .B(x[1334]), .Z(n4680) );
  NANDN U7330 ( .A(y[1335]), .B(x[1335]), .Z(n4679) );
  AND U7331 ( .A(n4680), .B(n4679), .Z(n12533) );
  NAND U7332 ( .A(n4681), .B(n12533), .Z(n4682) );
  NANDN U7333 ( .A(n12535), .B(n4682), .Z(n4683) );
  AND U7334 ( .A(n12537), .B(n4683), .Z(n4686) );
  NANDN U7335 ( .A(x[1338]), .B(y[1338]), .Z(n4685) );
  NANDN U7336 ( .A(x[1337]), .B(y[1337]), .Z(n4684) );
  NAND U7337 ( .A(n4685), .B(n4684), .Z(n12540) );
  OR U7338 ( .A(n4686), .B(n12540), .Z(n4689) );
  NANDN U7339 ( .A(y[1338]), .B(x[1338]), .Z(n4688) );
  NANDN U7340 ( .A(y[1339]), .B(x[1339]), .Z(n4687) );
  NAND U7341 ( .A(n4688), .B(n4687), .Z(n12542) );
  ANDN U7342 ( .B(n4689), .A(n12542), .Z(n4690) );
  NANDN U7343 ( .A(x[1339]), .B(y[1339]), .Z(n12544) );
  NANDN U7344 ( .A(n4690), .B(n12544), .Z(n4691) );
  NANDN U7345 ( .A(y[1340]), .B(x[1340]), .Z(n12545) );
  NAND U7346 ( .A(n4691), .B(n12545), .Z(n4692) );
  NANDN U7347 ( .A(x[1340]), .B(y[1340]), .Z(n8533) );
  ANDN U7348 ( .B(y[1341]), .A(x[1341]), .Z(n8539) );
  ANDN U7349 ( .B(n8533), .A(n8539), .Z(n12547) );
  NAND U7350 ( .A(n4692), .B(n12547), .Z(n4693) );
  NAND U7351 ( .A(n4694), .B(n4693), .Z(n4695) );
  NANDN U7352 ( .A(x[1342]), .B(y[1342]), .Z(n12551) );
  NAND U7353 ( .A(n4695), .B(n12551), .Z(n4696) );
  NAND U7354 ( .A(n4697), .B(n4696), .Z(n4699) );
  NANDN U7355 ( .A(x[1343]), .B(y[1343]), .Z(n4698) );
  NAND U7356 ( .A(n4699), .B(n4698), .Z(n4701) );
  OR U7357 ( .A(n4701), .B(y[1344]), .Z(n4700) );
  AND U7358 ( .A(n8549), .B(n4700), .Z(n4704) );
  XOR U7359 ( .A(n4701), .B(y[1344]), .Z(n4702) );
  NAND U7360 ( .A(n4702), .B(x[1344]), .Z(n4703) );
  NAND U7361 ( .A(n4704), .B(n4703), .Z(n4705) );
  NANDN U7362 ( .A(n12560), .B(n4705), .Z(n4712) );
  NANDN U7363 ( .A(y[1347]), .B(x[1347]), .Z(n4707) );
  ANDN U7364 ( .B(x[1348]), .A(y[1348]), .Z(n4706) );
  ANDN U7365 ( .B(n4707), .A(n4706), .Z(n4711) );
  XNOR U7366 ( .A(x[1347]), .B(y[1347]), .Z(n4709) );
  ANDN U7367 ( .B(x[1346]), .A(y[1346]), .Z(n4708) );
  NAND U7368 ( .A(n4709), .B(n4708), .Z(n4710) );
  AND U7369 ( .A(n4711), .B(n4710), .Z(n12561) );
  NAND U7370 ( .A(n4712), .B(n12561), .Z(n4713) );
  NANDN U7371 ( .A(n12564), .B(n4713), .Z(n4714) );
  NAND U7372 ( .A(n4715), .B(n4714), .Z(n4716) );
  NANDN U7373 ( .A(x[1350]), .B(y[1350]), .Z(n12567) );
  NAND U7374 ( .A(n4716), .B(n12567), .Z(n4717) );
  NANDN U7375 ( .A(x[1351]), .B(y[1351]), .Z(n12571) );
  NANDN U7376 ( .A(n4717), .B(n12571), .Z(n4718) );
  AND U7377 ( .A(n12573), .B(n4718), .Z(n4719) );
  NANDN U7378 ( .A(y[1351]), .B(x[1351]), .Z(n8557) );
  NAND U7379 ( .A(n4719), .B(n8557), .Z(n4720) );
  AND U7380 ( .A(n12575), .B(n4720), .Z(n4721) );
  ANDN U7381 ( .B(n12578), .A(n4721), .Z(n4722) );
  NANDN U7382 ( .A(y[1354]), .B(x[1354]), .Z(n6346) );
  NAND U7383 ( .A(n4722), .B(n6346), .Z(n4723) );
  AND U7384 ( .A(n12579), .B(n4723), .Z(n4724) );
  NANDN U7385 ( .A(y[1355]), .B(x[1355]), .Z(n6347) );
  NANDN U7386 ( .A(n4724), .B(n6347), .Z(n4727) );
  NANDN U7387 ( .A(x[1356]), .B(y[1356]), .Z(n4726) );
  NANDN U7388 ( .A(x[1355]), .B(y[1355]), .Z(n4725) );
  NAND U7389 ( .A(n4726), .B(n4725), .Z(n12583) );
  ANDN U7390 ( .B(n4727), .A(n12583), .Z(n4730) );
  NANDN U7391 ( .A(y[1356]), .B(x[1356]), .Z(n4729) );
  NANDN U7392 ( .A(y[1357]), .B(x[1357]), .Z(n4728) );
  AND U7393 ( .A(n4729), .B(n4728), .Z(n12585) );
  NANDN U7394 ( .A(n4730), .B(n12585), .Z(n4733) );
  NANDN U7395 ( .A(x[1358]), .B(y[1358]), .Z(n4732) );
  NANDN U7396 ( .A(x[1357]), .B(y[1357]), .Z(n4731) );
  NAND U7397 ( .A(n4732), .B(n4731), .Z(n12587) );
  ANDN U7398 ( .B(n4733), .A(n12587), .Z(n4736) );
  NANDN U7399 ( .A(y[1358]), .B(x[1358]), .Z(n4735) );
  NANDN U7400 ( .A(y[1359]), .B(x[1359]), .Z(n4734) );
  AND U7401 ( .A(n4735), .B(n4734), .Z(n12589) );
  NANDN U7402 ( .A(n4736), .B(n12589), .Z(n4737) );
  NANDN U7403 ( .A(n12591), .B(n4737), .Z(n4740) );
  NANDN U7404 ( .A(y[1360]), .B(x[1360]), .Z(n4739) );
  NANDN U7405 ( .A(y[1361]), .B(x[1361]), .Z(n4738) );
  AND U7406 ( .A(n4739), .B(n4738), .Z(n12593) );
  NAND U7407 ( .A(n4740), .B(n12593), .Z(n4743) );
  ANDN U7408 ( .B(y[1363]), .A(x[1363]), .Z(n8578) );
  NANDN U7409 ( .A(x[1362]), .B(y[1362]), .Z(n4742) );
  NANDN U7410 ( .A(x[1361]), .B(y[1361]), .Z(n4741) );
  NAND U7411 ( .A(n4742), .B(n4741), .Z(n8575) );
  NOR U7412 ( .A(n8578), .B(n8575), .Z(n12596) );
  NAND U7413 ( .A(n4743), .B(n12596), .Z(n4747) );
  NANDN U7414 ( .A(y[1364]), .B(x[1364]), .Z(n8583) );
  NANDN U7415 ( .A(y[1363]), .B(x[1363]), .Z(n4745) );
  NANDN U7416 ( .A(y[1362]), .B(x[1362]), .Z(n4744) );
  AND U7417 ( .A(n4745), .B(n4744), .Z(n8576) );
  OR U7418 ( .A(n8578), .B(n8576), .Z(n4746) );
  NAND U7419 ( .A(n8583), .B(n4746), .Z(n12597) );
  ANDN U7420 ( .B(n4747), .A(n12597), .Z(n4748) );
  OR U7421 ( .A(n12599), .B(n4748), .Z(n4749) );
  NAND U7422 ( .A(n4750), .B(n4749), .Z(n4751) );
  NANDN U7423 ( .A(x[1366]), .B(y[1366]), .Z(n12603) );
  NAND U7424 ( .A(n4751), .B(n12603), .Z(n4752) );
  NAND U7425 ( .A(n4753), .B(n4752), .Z(n4754) );
  NAND U7426 ( .A(n8593), .B(n4754), .Z(n4755) );
  NAND U7427 ( .A(n4756), .B(n4755), .Z(n4757) );
  NAND U7428 ( .A(n4758), .B(n4757), .Z(n4759) );
  ANDN U7429 ( .B(x[1369]), .A(y[1369]), .Z(n8595) );
  ANDN U7430 ( .B(n4759), .A(n8595), .Z(n4760) );
  OR U7431 ( .A(n12612), .B(n4760), .Z(n4761) );
  AND U7432 ( .A(n12613), .B(n4761), .Z(n4766) );
  NANDN U7433 ( .A(x[1372]), .B(y[1372]), .Z(n4763) );
  NANDN U7434 ( .A(x[1371]), .B(y[1371]), .Z(n4762) );
  AND U7435 ( .A(n4763), .B(n4762), .Z(n4765) );
  AND U7436 ( .A(n4765), .B(n4764), .Z(n12615) );
  NANDN U7437 ( .A(n4766), .B(n12615), .Z(n4767) );
  NAND U7438 ( .A(n4768), .B(n4767), .Z(n4769) );
  NANDN U7439 ( .A(n12620), .B(n4769), .Z(n4774) );
  NANDN U7440 ( .A(y[1376]), .B(x[1376]), .Z(n4771) );
  NANDN U7441 ( .A(y[1375]), .B(x[1375]), .Z(n4770) );
  AND U7442 ( .A(n4771), .B(n4770), .Z(n4773) );
  AND U7443 ( .A(n4773), .B(n4772), .Z(n6344) );
  NAND U7444 ( .A(n4774), .B(n6344), .Z(n4775) );
  NANDN U7445 ( .A(n8605), .B(n4775), .Z(n4776) );
  IV U7446 ( .A(x[1378]), .Z(n6337) );
  OR U7447 ( .A(n4776), .B(n6337), .Z(n4779) );
  XNOR U7448 ( .A(n4776), .B(x[1378]), .Z(n4777) );
  NANDN U7449 ( .A(y[1378]), .B(n4777), .Z(n4778) );
  NAND U7450 ( .A(n4779), .B(n4778), .Z(n4780) );
  NAND U7451 ( .A(n4781), .B(n4780), .Z(n4782) );
  NAND U7452 ( .A(n4783), .B(n4782), .Z(n4784) );
  NANDN U7453 ( .A(n8608), .B(n4784), .Z(n4785) );
  IV U7454 ( .A(x[1381]), .Z(n6334) );
  OR U7455 ( .A(n4785), .B(n6334), .Z(n4788) );
  XNOR U7456 ( .A(n4785), .B(x[1381]), .Z(n4786) );
  NANDN U7457 ( .A(y[1381]), .B(n4786), .Z(n4787) );
  AND U7458 ( .A(n4788), .B(n4787), .Z(n4790) );
  NANDN U7459 ( .A(n4790), .B(x[1382]), .Z(n4789) );
  AND U7460 ( .A(n8613), .B(n4789), .Z(n4793) );
  XNOR U7461 ( .A(n4790), .B(x[1382]), .Z(n4791) );
  NANDN U7462 ( .A(y[1382]), .B(n4791), .Z(n4792) );
  AND U7463 ( .A(n4793), .B(n4792), .Z(n4796) );
  NANDN U7464 ( .A(x[1383]), .B(y[1383]), .Z(n4795) );
  NANDN U7465 ( .A(x[1384]), .B(y[1384]), .Z(n4794) );
  AND U7466 ( .A(n4795), .B(n4794), .Z(n12635) );
  NANDN U7467 ( .A(n4796), .B(n12635), .Z(n4799) );
  NANDN U7468 ( .A(y[1385]), .B(x[1385]), .Z(n4798) );
  NANDN U7469 ( .A(y[1384]), .B(x[1384]), .Z(n4797) );
  NAND U7470 ( .A(n4798), .B(n4797), .Z(n12637) );
  ANDN U7471 ( .B(n4799), .A(n12637), .Z(n4802) );
  NANDN U7472 ( .A(x[1385]), .B(y[1385]), .Z(n4801) );
  NANDN U7473 ( .A(x[1386]), .B(y[1386]), .Z(n4800) );
  AND U7474 ( .A(n4801), .B(n4800), .Z(n12639) );
  NANDN U7475 ( .A(n4802), .B(n12639), .Z(n4805) );
  NANDN U7476 ( .A(y[1386]), .B(x[1386]), .Z(n4804) );
  NANDN U7477 ( .A(y[1387]), .B(x[1387]), .Z(n4803) );
  NAND U7478 ( .A(n4804), .B(n4803), .Z(n12641) );
  ANDN U7479 ( .B(n4805), .A(n12641), .Z(n4806) );
  NANDN U7480 ( .A(x[1387]), .B(y[1387]), .Z(n12643) );
  NANDN U7481 ( .A(n4806), .B(n12643), .Z(n4807) );
  NANDN U7482 ( .A(y[1388]), .B(x[1388]), .Z(n12645) );
  NAND U7483 ( .A(n4807), .B(n12645), .Z(n4808) );
  NANDN U7484 ( .A(n12648), .B(n4808), .Z(n4809) );
  NAND U7485 ( .A(n4810), .B(n4809), .Z(n4811) );
  NANDN U7486 ( .A(x[1391]), .B(y[1391]), .Z(n8632) );
  NAND U7487 ( .A(n4811), .B(n8632), .Z(n4812) );
  NANDN U7488 ( .A(x[1390]), .B(y[1390]), .Z(n12651) );
  NANDN U7489 ( .A(n4812), .B(n12651), .Z(n4813) );
  AND U7490 ( .A(n8628), .B(n4813), .Z(n4814) );
  NAND U7491 ( .A(n4815), .B(n4814), .Z(n4816) );
  NAND U7492 ( .A(n8631), .B(n4816), .Z(n4817) );
  AND U7493 ( .A(n8634), .B(n4817), .Z(n4820) );
  NANDN U7494 ( .A(x[1393]), .B(y[1393]), .Z(n4819) );
  NANDN U7495 ( .A(x[1394]), .B(y[1394]), .Z(n4818) );
  AND U7496 ( .A(n4819), .B(n4818), .Z(n12659) );
  NANDN U7497 ( .A(n4820), .B(n12659), .Z(n4823) );
  NANDN U7498 ( .A(y[1395]), .B(x[1395]), .Z(n4822) );
  NANDN U7499 ( .A(y[1394]), .B(x[1394]), .Z(n4821) );
  NAND U7500 ( .A(n4822), .B(n4821), .Z(n12661) );
  ANDN U7501 ( .B(n4823), .A(n12661), .Z(n4826) );
  NANDN U7502 ( .A(x[1395]), .B(y[1395]), .Z(n4825) );
  NANDN U7503 ( .A(x[1396]), .B(y[1396]), .Z(n4824) );
  AND U7504 ( .A(n4825), .B(n4824), .Z(n12663) );
  NANDN U7505 ( .A(n4826), .B(n12663), .Z(n4827) );
  NANDN U7506 ( .A(n12665), .B(n4827), .Z(n4828) );
  NANDN U7507 ( .A(x[1397]), .B(y[1397]), .Z(n6333) );
  NAND U7508 ( .A(n4828), .B(n6333), .Z(n4830) );
  NANDN U7509 ( .A(x[1398]), .B(n4830), .Z(n4829) );
  AND U7510 ( .A(n12671), .B(n4829), .Z(n4833) );
  XNOR U7511 ( .A(x[1398]), .B(n4830), .Z(n4831) );
  NAND U7512 ( .A(n4831), .B(y[1398]), .Z(n4832) );
  NAND U7513 ( .A(n4833), .B(n4832), .Z(n4834) );
  NAND U7514 ( .A(n4835), .B(n4834), .Z(n4836) );
  ANDN U7515 ( .B(y[1400]), .A(x[1400]), .Z(n8645) );
  ANDN U7516 ( .B(y[1401]), .A(x[1401]), .Z(n8650) );
  NOR U7517 ( .A(n8645), .B(n8650), .Z(n12675) );
  NAND U7518 ( .A(n4836), .B(n12675), .Z(n4837) );
  ANDN U7519 ( .B(x[1402]), .A(y[1402]), .Z(n8653) );
  ANDN U7520 ( .B(n4837), .A(n8653), .Z(n4838) );
  NANDN U7521 ( .A(y[1401]), .B(x[1401]), .Z(n12677) );
  NAND U7522 ( .A(n4838), .B(n12677), .Z(n4839) );
  AND U7523 ( .A(n8657), .B(n4839), .Z(n4840) );
  NANDN U7524 ( .A(x[1402]), .B(y[1402]), .Z(n12679) );
  NAND U7525 ( .A(n4840), .B(n12679), .Z(n4841) );
  NANDN U7526 ( .A(n8654), .B(n4841), .Z(n4843) );
  NANDN U7527 ( .A(y[1404]), .B(n4843), .Z(n4842) );
  AND U7528 ( .A(n6331), .B(n4842), .Z(n4846) );
  XNOR U7529 ( .A(n4843), .B(y[1404]), .Z(n4844) );
  NAND U7530 ( .A(n4844), .B(x[1404]), .Z(n4845) );
  NAND U7531 ( .A(n4846), .B(n4845), .Z(n4847) );
  NANDN U7532 ( .A(n12688), .B(n4847), .Z(n4848) );
  NANDN U7533 ( .A(n12689), .B(n4848), .Z(n4855) );
  NANDN U7534 ( .A(x[1410]), .B(y[1410]), .Z(n4854) );
  ANDN U7535 ( .B(y[1408]), .A(x[1408]), .Z(n4849) );
  OR U7536 ( .A(n4849), .B(y[1409]), .Z(n4852) );
  XOR U7537 ( .A(y[1409]), .B(n4849), .Z(n4850) );
  NAND U7538 ( .A(n4850), .B(x[1409]), .Z(n4851) );
  NAND U7539 ( .A(n4852), .B(n4851), .Z(n4853) );
  NAND U7540 ( .A(n4854), .B(n4853), .Z(n12692) );
  ANDN U7541 ( .B(n4855), .A(n12692), .Z(n4858) );
  NANDN U7542 ( .A(y[1411]), .B(x[1411]), .Z(n4857) );
  NANDN U7543 ( .A(y[1410]), .B(x[1410]), .Z(n4856) );
  AND U7544 ( .A(n4857), .B(n4856), .Z(n12694) );
  NANDN U7545 ( .A(n4858), .B(n12694), .Z(n4859) );
  AND U7546 ( .A(n12695), .B(n4859), .Z(n4860) );
  NANDN U7547 ( .A(y[1412]), .B(x[1412]), .Z(n8668) );
  NANDN U7548 ( .A(n4860), .B(n8668), .Z(n4861) );
  ANDN U7549 ( .B(y[1413]), .A(x[1413]), .Z(n8670) );
  ANDN U7550 ( .B(y[1412]), .A(x[1412]), .Z(n8664) );
  OR U7551 ( .A(n8670), .B(n8664), .Z(n12701) );
  ANDN U7552 ( .B(n4861), .A(n12701), .Z(n4862) );
  NOR U7553 ( .A(n12702), .B(n4862), .Z(n4863) );
  NANDN U7554 ( .A(y[1414]), .B(x[1414]), .Z(n6329) );
  NAND U7555 ( .A(n4863), .B(n6329), .Z(n4864) );
  AND U7556 ( .A(n12699), .B(n4864), .Z(n4865) );
  NAND U7557 ( .A(n4866), .B(n4865), .Z(n4867) );
  NAND U7558 ( .A(n4868), .B(n4867), .Z(n4869) );
  ANDN U7559 ( .B(y[1416]), .A(x[1416]), .Z(n8674) );
  ANDN U7560 ( .B(n4869), .A(n8674), .Z(n4870) );
  NAND U7561 ( .A(n4871), .B(n4870), .Z(n4872) );
  NAND U7562 ( .A(n4873), .B(n4872), .Z(n4874) );
  ANDN U7563 ( .B(y[1418]), .A(x[1418]), .Z(n8682) );
  ANDN U7564 ( .B(n4874), .A(n8682), .Z(n4877) );
  NANDN U7565 ( .A(y[1419]), .B(x[1419]), .Z(n4876) );
  NANDN U7566 ( .A(y[1418]), .B(x[1418]), .Z(n4875) );
  NAND U7567 ( .A(n4876), .B(n4875), .Z(n12714) );
  OR U7568 ( .A(n4877), .B(n12714), .Z(n4882) );
  NANDN U7569 ( .A(x[1420]), .B(y[1420]), .Z(n4879) );
  NANDN U7570 ( .A(x[1419]), .B(y[1419]), .Z(n4878) );
  AND U7571 ( .A(n4879), .B(n4878), .Z(n4881) );
  NANDN U7572 ( .A(x[1421]), .B(y[1421]), .Z(n4880) );
  AND U7573 ( .A(n4881), .B(n4880), .Z(n12716) );
  NAND U7574 ( .A(n4882), .B(n12716), .Z(n4883) );
  NANDN U7575 ( .A(y[1422]), .B(x[1422]), .Z(n8689) );
  NAND U7576 ( .A(n4883), .B(n8689), .Z(n4888) );
  NANDN U7577 ( .A(y[1420]), .B(x[1420]), .Z(n4884) );
  NANDN U7578 ( .A(n4884), .B(x[1421]), .Z(n4887) );
  XNOR U7579 ( .A(n4884), .B(x[1421]), .Z(n4885) );
  NANDN U7580 ( .A(y[1421]), .B(n4885), .Z(n4886) );
  AND U7581 ( .A(n4887), .B(n4886), .Z(n12717) );
  NANDN U7582 ( .A(n4888), .B(n12717), .Z(n4890) );
  ANDN U7583 ( .B(y[1423]), .A(x[1423]), .Z(n8690) );
  NANDN U7584 ( .A(x[1422]), .B(y[1422]), .Z(n4889) );
  NANDN U7585 ( .A(n8690), .B(n4889), .Z(n12719) );
  ANDN U7586 ( .B(n4890), .A(n12719), .Z(n4893) );
  NANDN U7587 ( .A(y[1424]), .B(x[1424]), .Z(n4892) );
  NANDN U7588 ( .A(y[1423]), .B(x[1423]), .Z(n4891) );
  AND U7589 ( .A(n4892), .B(n4891), .Z(n8693) );
  NANDN U7590 ( .A(n4893), .B(n8693), .Z(n4894) );
  NANDN U7591 ( .A(n6325), .B(n4894), .Z(n4895) );
  NANDN U7592 ( .A(y[1426]), .B(x[1426]), .Z(n8698) );
  NAND U7593 ( .A(n4895), .B(n8698), .Z(n4896) );
  NANDN U7594 ( .A(y[1425]), .B(x[1425]), .Z(n8692) );
  NANDN U7595 ( .A(n4896), .B(n8692), .Z(n4897) );
  NAND U7596 ( .A(n4898), .B(n4897), .Z(n4899) );
  ANDN U7597 ( .B(x[1427]), .A(y[1427]), .Z(n8697) );
  ANDN U7598 ( .B(n4899), .A(n8697), .Z(n4900) );
  NAND U7599 ( .A(n4901), .B(n4900), .Z(n4902) );
  NAND U7600 ( .A(n4903), .B(n4902), .Z(n4904) );
  AND U7601 ( .A(n8701), .B(n4904), .Z(n4907) );
  NANDN U7602 ( .A(x[1429]), .B(y[1429]), .Z(n4906) );
  NANDN U7603 ( .A(x[1430]), .B(y[1430]), .Z(n4905) );
  AND U7604 ( .A(n4906), .B(n4905), .Z(n12731) );
  NANDN U7605 ( .A(n4907), .B(n12731), .Z(n4910) );
  NANDN U7606 ( .A(y[1430]), .B(x[1430]), .Z(n4909) );
  NANDN U7607 ( .A(y[1431]), .B(x[1431]), .Z(n4908) );
  NAND U7608 ( .A(n4909), .B(n4908), .Z(n12733) );
  ANDN U7609 ( .B(n4910), .A(n12733), .Z(n4911) );
  NANDN U7610 ( .A(x[1431]), .B(y[1431]), .Z(n12735) );
  NANDN U7611 ( .A(n4911), .B(n12735), .Z(n4912) );
  NANDN U7612 ( .A(n12738), .B(n4912), .Z(n4913) );
  NANDN U7613 ( .A(n12740), .B(n4913), .Z(n4914) );
  NANDN U7614 ( .A(n8712), .B(n4914), .Z(n4915) );
  NANDN U7615 ( .A(x[1435]), .B(y[1435]), .Z(n12744) );
  NAND U7616 ( .A(n4915), .B(n12744), .Z(n4916) );
  NANDN U7617 ( .A(y[1436]), .B(x[1436]), .Z(n12745) );
  NAND U7618 ( .A(n4916), .B(n12745), .Z(n4917) );
  NANDN U7619 ( .A(y[1435]), .B(x[1435]), .Z(n8713) );
  NANDN U7620 ( .A(n4917), .B(n8713), .Z(n4918) );
  NANDN U7621 ( .A(n12747), .B(n4918), .Z(n4919) );
  NANDN U7622 ( .A(y[1438]), .B(x[1438]), .Z(n8724) );
  NAND U7623 ( .A(n4919), .B(n8724), .Z(n4920) );
  NANDN U7624 ( .A(y[1437]), .B(x[1437]), .Z(n12749) );
  NANDN U7625 ( .A(n4920), .B(n12749), .Z(n4921) );
  AND U7626 ( .A(n12751), .B(n4921), .Z(n4924) );
  NANDN U7627 ( .A(y[1441]), .B(x[1441]), .Z(n4923) );
  NANDN U7628 ( .A(y[1440]), .B(x[1440]), .Z(n4922) );
  NAND U7629 ( .A(n4923), .B(n4922), .Z(n8728) );
  NOR U7630 ( .A(n4924), .B(n8728), .Z(n4925) );
  NAND U7631 ( .A(n4926), .B(n4925), .Z(n4927) );
  NANDN U7632 ( .A(x[1442]), .B(y[1442]), .Z(n12759) );
  ANDN U7633 ( .B(y[1441]), .A(x[1441]), .Z(n12756) );
  ANDN U7634 ( .B(n12759), .A(n12756), .Z(n8730) );
  NAND U7635 ( .A(n4927), .B(n8730), .Z(n4928) );
  NANDN U7636 ( .A(n12758), .B(n4928), .Z(n4930) );
  NANDN U7637 ( .A(x[1443]), .B(y[1443]), .Z(n4929) );
  ANDN U7638 ( .B(y[1444]), .A(x[1444]), .Z(n12768) );
  ANDN U7639 ( .B(n4929), .A(n12768), .Z(n8733) );
  NAND U7640 ( .A(n4930), .B(n8733), .Z(n4932) );
  NANDN U7641 ( .A(y[1445]), .B(x[1445]), .Z(n12769) );
  NANDN U7642 ( .A(y[1444]), .B(x[1444]), .Z(n4931) );
  NAND U7643 ( .A(n12769), .B(n4931), .Z(n12766) );
  ANDN U7644 ( .B(n4932), .A(n12766), .Z(n4933) );
  NANDN U7645 ( .A(x[1445]), .B(y[1445]), .Z(n12767) );
  NANDN U7646 ( .A(n4933), .B(n12767), .Z(n4934) );
  ANDN U7647 ( .B(x[1446]), .A(y[1446]), .Z(n6319) );
  ANDN U7648 ( .B(n4934), .A(n6319), .Z(n4935) );
  NANDN U7649 ( .A(x[1447]), .B(y[1447]), .Z(n8740) );
  ANDN U7650 ( .B(y[1446]), .A(x[1446]), .Z(n8736) );
  ANDN U7651 ( .B(n8740), .A(n8736), .Z(n12772) );
  NANDN U7652 ( .A(n4935), .B(n12772), .Z(n4936) );
  AND U7653 ( .A(n4937), .B(n4936), .Z(n4938) );
  ANDN U7654 ( .B(y[1448]), .A(x[1448]), .Z(n8743) );
  ANDN U7655 ( .B(y[1449]), .A(x[1449]), .Z(n6318) );
  NOR U7656 ( .A(n8743), .B(n6318), .Z(n12782) );
  NANDN U7657 ( .A(n4938), .B(n12782), .Z(n4940) );
  NANDN U7658 ( .A(y[1449]), .B(x[1449]), .Z(n12783) );
  ANDN U7659 ( .B(x[1450]), .A(y[1450]), .Z(n8748) );
  ANDN U7660 ( .B(n12783), .A(n8748), .Z(n4939) );
  NAND U7661 ( .A(n4940), .B(n4939), .Z(n4941) );
  NANDN U7662 ( .A(x[1451]), .B(y[1451]), .Z(n6316) );
  NAND U7663 ( .A(n4941), .B(n6316), .Z(n4942) );
  NANDN U7664 ( .A(x[1450]), .B(y[1450]), .Z(n12785) );
  NANDN U7665 ( .A(n4942), .B(n12785), .Z(n4943) );
  AND U7666 ( .A(n4944), .B(n4943), .Z(n4945) );
  ANDN U7667 ( .B(n4946), .A(n4945), .Z(n4947) );
  AND U7668 ( .A(n12793), .B(n4947), .Z(n4950) );
  NANDN U7669 ( .A(y[1454]), .B(x[1454]), .Z(n4949) );
  NANDN U7670 ( .A(y[1455]), .B(x[1455]), .Z(n4948) );
  AND U7671 ( .A(n4949), .B(n4948), .Z(n12795) );
  NANDN U7672 ( .A(n4950), .B(n12795), .Z(n4953) );
  NANDN U7673 ( .A(x[1456]), .B(y[1456]), .Z(n4952) );
  NANDN U7674 ( .A(x[1455]), .B(y[1455]), .Z(n4951) );
  NAND U7675 ( .A(n4952), .B(n4951), .Z(n12798) );
  ANDN U7676 ( .B(n4953), .A(n12798), .Z(n4956) );
  NANDN U7677 ( .A(y[1456]), .B(x[1456]), .Z(n4955) );
  NANDN U7678 ( .A(y[1457]), .B(x[1457]), .Z(n4954) );
  AND U7679 ( .A(n4955), .B(n4954), .Z(n12800) );
  NANDN U7680 ( .A(n4956), .B(n12800), .Z(n4957) );
  NANDN U7681 ( .A(n8757), .B(n4957), .Z(n4958) );
  NANDN U7682 ( .A(y[1458]), .B(x[1458]), .Z(n8761) );
  NAND U7683 ( .A(n4958), .B(n8761), .Z(n4959) );
  NAND U7684 ( .A(n4960), .B(n4959), .Z(n4962) );
  NANDN U7685 ( .A(y[1460]), .B(x[1460]), .Z(n12807) );
  ANDN U7686 ( .B(x[1459]), .A(y[1459]), .Z(n8760) );
  ANDN U7687 ( .B(n12807), .A(n8760), .Z(n4961) );
  NAND U7688 ( .A(n4962), .B(n4961), .Z(n4963) );
  ANDN U7689 ( .B(y[1461]), .A(x[1461]), .Z(n8770) );
  ANDN U7690 ( .B(y[1460]), .A(x[1460]), .Z(n8765) );
  NOR U7691 ( .A(n8770), .B(n8765), .Z(n12809) );
  NAND U7692 ( .A(n4963), .B(n12809), .Z(n4964) );
  NAND U7693 ( .A(n4965), .B(n4964), .Z(n4966) );
  NANDN U7694 ( .A(x[1462]), .B(y[1462]), .Z(n12813) );
  NAND U7695 ( .A(n4966), .B(n12813), .Z(n4967) );
  NAND U7696 ( .A(n4968), .B(n4967), .Z(n4969) );
  NAND U7697 ( .A(n8776), .B(n4969), .Z(n4970) );
  NAND U7698 ( .A(n4971), .B(n4970), .Z(n4972) );
  NAND U7699 ( .A(n4973), .B(n4972), .Z(n4974) );
  ANDN U7700 ( .B(x[1465]), .A(y[1465]), .Z(n8778) );
  ANDN U7701 ( .B(n4974), .A(n8778), .Z(n4975) );
  OR U7702 ( .A(n12822), .B(n4975), .Z(n4976) );
  AND U7703 ( .A(n12823), .B(n4976), .Z(n4979) );
  NANDN U7704 ( .A(x[1469]), .B(y[1469]), .Z(n4978) );
  NANDN U7705 ( .A(x[1468]), .B(y[1468]), .Z(n4977) );
  NAND U7706 ( .A(n4978), .B(n4977), .Z(n12826) );
  OR U7707 ( .A(n4979), .B(n12826), .Z(n4980) );
  AND U7708 ( .A(n6312), .B(n4980), .Z(n4981) );
  NANDN U7709 ( .A(y[1469]), .B(x[1469]), .Z(n12828) );
  NAND U7710 ( .A(n4981), .B(n12828), .Z(n4982) );
  NANDN U7711 ( .A(n12830), .B(n4982), .Z(n4987) );
  NANDN U7712 ( .A(y[1472]), .B(x[1472]), .Z(n4984) );
  NANDN U7713 ( .A(y[1471]), .B(x[1471]), .Z(n4983) );
  AND U7714 ( .A(n4984), .B(n4983), .Z(n4986) );
  NANDN U7715 ( .A(y[1473]), .B(x[1473]), .Z(n4985) );
  NAND U7716 ( .A(n4986), .B(n4985), .Z(n6315) );
  ANDN U7717 ( .B(n4987), .A(n6315), .Z(n4994) );
  NANDN U7718 ( .A(x[1473]), .B(y[1473]), .Z(n4989) );
  ANDN U7719 ( .B(y[1474]), .A(x[1474]), .Z(n4988) );
  ANDN U7720 ( .B(n4989), .A(n4988), .Z(n4993) );
  XNOR U7721 ( .A(y[1473]), .B(x[1473]), .Z(n4991) );
  ANDN U7722 ( .B(y[1472]), .A(x[1472]), .Z(n4990) );
  NAND U7723 ( .A(n4991), .B(n4990), .Z(n4992) );
  AND U7724 ( .A(n4993), .B(n4992), .Z(n12833) );
  NANDN U7725 ( .A(n4994), .B(n12833), .Z(n4995) );
  NANDN U7726 ( .A(n12836), .B(n4995), .Z(n4996) );
  NANDN U7727 ( .A(x[1475]), .B(y[1475]), .Z(n6311) );
  NAND U7728 ( .A(n4996), .B(n6311), .Z(n4997) );
  NANDN U7729 ( .A(x[1476]), .B(n4997), .Z(n5000) );
  IV U7730 ( .A(y[1476]), .Z(n6309) );
  XNOR U7731 ( .A(x[1476]), .B(n4997), .Z(n4998) );
  NANDN U7732 ( .A(n6309), .B(n4998), .Z(n4999) );
  NAND U7733 ( .A(n5000), .B(n4999), .Z(n5001) );
  AND U7734 ( .A(n6307), .B(n5001), .Z(n5004) );
  NANDN U7735 ( .A(x[1477]), .B(y[1477]), .Z(n5003) );
  NANDN U7736 ( .A(x[1478]), .B(y[1478]), .Z(n5002) );
  AND U7737 ( .A(n5003), .B(n5002), .Z(n12841) );
  NANDN U7738 ( .A(n5004), .B(n12841), .Z(n5005) );
  NANDN U7739 ( .A(n12843), .B(n5005), .Z(n5010) );
  NANDN U7740 ( .A(x[1480]), .B(y[1480]), .Z(n5007) );
  NANDN U7741 ( .A(x[1479]), .B(y[1479]), .Z(n5006) );
  AND U7742 ( .A(n5007), .B(n5006), .Z(n5009) );
  AND U7743 ( .A(n5009), .B(n5008), .Z(n12845) );
  NAND U7744 ( .A(n5010), .B(n12845), .Z(n5011) );
  NAND U7745 ( .A(n5012), .B(n5011), .Z(n5014) );
  NANDN U7746 ( .A(x[1482]), .B(y[1482]), .Z(n5013) );
  NANDN U7747 ( .A(x[1483]), .B(y[1483]), .Z(n8798) );
  AND U7748 ( .A(n5013), .B(n8798), .Z(n12849) );
  NAND U7749 ( .A(n5014), .B(n12849), .Z(n5017) );
  NANDN U7750 ( .A(y[1484]), .B(x[1484]), .Z(n5016) );
  NANDN U7751 ( .A(y[1483]), .B(x[1483]), .Z(n5015) );
  AND U7752 ( .A(n5016), .B(n5015), .Z(n8796) );
  NAND U7753 ( .A(n5017), .B(n8796), .Z(n5020) );
  NANDN U7754 ( .A(x[1484]), .B(y[1484]), .Z(n5019) );
  NANDN U7755 ( .A(x[1485]), .B(y[1485]), .Z(n5018) );
  NAND U7756 ( .A(n5019), .B(n5018), .Z(n6304) );
  ANDN U7757 ( .B(n5020), .A(n6304), .Z(n5021) );
  NANDN U7758 ( .A(y[1485]), .B(x[1485]), .Z(n8797) );
  NANDN U7759 ( .A(n5021), .B(n8797), .Z(n5022) );
  IV U7760 ( .A(y[1486]), .Z(n6303) );
  OR U7761 ( .A(n5022), .B(n6303), .Z(n5025) );
  XNOR U7762 ( .A(n5022), .B(y[1486]), .Z(n5023) );
  NANDN U7763 ( .A(x[1486]), .B(n5023), .Z(n5024) );
  AND U7764 ( .A(n5025), .B(n5024), .Z(n5027) );
  NANDN U7765 ( .A(n5027), .B(y[1487]), .Z(n5026) );
  AND U7766 ( .A(n8805), .B(n5026), .Z(n5030) );
  XNOR U7767 ( .A(n5027), .B(y[1487]), .Z(n5028) );
  NANDN U7768 ( .A(x[1487]), .B(n5028), .Z(n5029) );
  AND U7769 ( .A(n5030), .B(n5029), .Z(n5033) );
  NANDN U7770 ( .A(y[1488]), .B(x[1488]), .Z(n5032) );
  NANDN U7771 ( .A(y[1489]), .B(x[1489]), .Z(n5031) );
  AND U7772 ( .A(n5032), .B(n5031), .Z(n12859) );
  NANDN U7773 ( .A(n5033), .B(n12859), .Z(n5036) );
  NANDN U7774 ( .A(x[1490]), .B(y[1490]), .Z(n5035) );
  NANDN U7775 ( .A(x[1489]), .B(y[1489]), .Z(n5034) );
  NAND U7776 ( .A(n5035), .B(n5034), .Z(n12861) );
  ANDN U7777 ( .B(n5036), .A(n12861), .Z(n5039) );
  NANDN U7778 ( .A(y[1490]), .B(x[1490]), .Z(n5038) );
  NANDN U7779 ( .A(y[1491]), .B(x[1491]), .Z(n5037) );
  AND U7780 ( .A(n5038), .B(n5037), .Z(n12863) );
  NANDN U7781 ( .A(n5039), .B(n12863), .Z(n5040) );
  NANDN U7782 ( .A(n6300), .B(n5040), .Z(n5047) );
  NANDN U7783 ( .A(y[1492]), .B(x[1492]), .Z(n5041) );
  NANDN U7784 ( .A(n5042), .B(n5041), .Z(n5043) );
  NANDN U7785 ( .A(n5044), .B(n5043), .Z(n5046) );
  NAND U7786 ( .A(n5046), .B(n5045), .Z(n8812) );
  ANDN U7787 ( .B(n5047), .A(n8812), .Z(n5048) );
  OR U7788 ( .A(n5049), .B(n5048), .Z(n5050) );
  AND U7789 ( .A(n5051), .B(n5050), .Z(n5052) );
  ANDN U7790 ( .B(y[1497]), .A(x[1497]), .Z(n8820) );
  ANDN U7791 ( .B(y[1496]), .A(x[1496]), .Z(n8815) );
  NOR U7792 ( .A(n8820), .B(n8815), .Z(n12873) );
  NANDN U7793 ( .A(n5052), .B(n12873), .Z(n5053) );
  ANDN U7794 ( .B(x[1498]), .A(y[1498]), .Z(n8823) );
  ANDN U7795 ( .B(n5053), .A(n8823), .Z(n5054) );
  NANDN U7796 ( .A(y[1497]), .B(x[1497]), .Z(n12876) );
  NAND U7797 ( .A(n5054), .B(n12876), .Z(n5055) );
  AND U7798 ( .A(n6298), .B(n5055), .Z(n5056) );
  NANDN U7799 ( .A(x[1498]), .B(y[1498]), .Z(n12877) );
  NAND U7800 ( .A(n5056), .B(n12877), .Z(n5057) );
  NANDN U7801 ( .A(n8824), .B(n5057), .Z(n5061) );
  OR U7802 ( .A(n5061), .B(x[1500]), .Z(n5060) );
  NANDN U7803 ( .A(x[1501]), .B(y[1501]), .Z(n5058) );
  NAND U7804 ( .A(n5059), .B(n5058), .Z(n12886) );
  ANDN U7805 ( .B(n5060), .A(n12886), .Z(n5064) );
  XOR U7806 ( .A(n5061), .B(x[1500]), .Z(n5062) );
  NAND U7807 ( .A(n5062), .B(y[1500]), .Z(n5063) );
  NAND U7808 ( .A(n5064), .B(n5063), .Z(n5065) );
  AND U7809 ( .A(n12887), .B(n5065), .Z(n5066) );
  NAND U7810 ( .A(n5067), .B(n5066), .Z(n5068) );
  NANDN U7811 ( .A(n12890), .B(n5068), .Z(n5069) );
  AND U7812 ( .A(n12891), .B(n5069), .Z(n5072) );
  NANDN U7813 ( .A(x[1506]), .B(y[1506]), .Z(n5071) );
  NANDN U7814 ( .A(x[1505]), .B(y[1505]), .Z(n5070) );
  NAND U7815 ( .A(n5071), .B(n5070), .Z(n8833) );
  NOR U7816 ( .A(n8836), .B(n8833), .Z(n12894) );
  NANDN U7817 ( .A(n5072), .B(n12894), .Z(n5073) );
  NANDN U7818 ( .A(n12895), .B(n5073), .Z(n5074) );
  ANDN U7819 ( .B(y[1509]), .A(x[1509]), .Z(n8843) );
  ANDN U7820 ( .B(y[1508]), .A(x[1508]), .Z(n8839) );
  NOR U7821 ( .A(n8843), .B(n8839), .Z(n12897) );
  NAND U7822 ( .A(n5074), .B(n12897), .Z(n5075) );
  AND U7823 ( .A(n5076), .B(n5075), .Z(n5080) );
  NANDN U7824 ( .A(x[1511]), .B(y[1511]), .Z(n5077) );
  NAND U7825 ( .A(n5078), .B(n5077), .Z(n8849) );
  NANDN U7826 ( .A(x[1510]), .B(y[1510]), .Z(n5079) );
  NANDN U7827 ( .A(n8849), .B(n5079), .Z(n12902) );
  OR U7828 ( .A(n5080), .B(n12902), .Z(n5083) );
  NANDN U7829 ( .A(y[1512]), .B(x[1512]), .Z(n5082) );
  NANDN U7830 ( .A(y[1513]), .B(x[1513]), .Z(n5081) );
  NAND U7831 ( .A(n5082), .B(n5081), .Z(n8850) );
  ANDN U7832 ( .B(n5083), .A(n8850), .Z(n5084) );
  NAND U7833 ( .A(n5085), .B(n5084), .Z(n5086) );
  NANDN U7834 ( .A(n12905), .B(n5086), .Z(n5089) );
  NANDN U7835 ( .A(y[1515]), .B(x[1515]), .Z(n5088) );
  NANDN U7836 ( .A(y[1514]), .B(x[1514]), .Z(n5087) );
  AND U7837 ( .A(n5088), .B(n5087), .Z(n12907) );
  NAND U7838 ( .A(n5089), .B(n12907), .Z(n5090) );
  NANDN U7839 ( .A(x[1515]), .B(y[1515]), .Z(n12909) );
  NAND U7840 ( .A(n5090), .B(n12909), .Z(n5091) );
  AND U7841 ( .A(n12911), .B(n5091), .Z(n5097) );
  NANDN U7842 ( .A(x[1519]), .B(y[1519]), .Z(n8862) );
  ANDN U7843 ( .B(y[1516]), .A(x[1516]), .Z(n6294) );
  NAND U7844 ( .A(n5092), .B(n6294), .Z(n5093) );
  AND U7845 ( .A(n8862), .B(n5093), .Z(n5096) );
  NANDN U7846 ( .A(x[1517]), .B(y[1517]), .Z(n5095) );
  NANDN U7847 ( .A(x[1518]), .B(y[1518]), .Z(n5094) );
  NAND U7848 ( .A(n5095), .B(n5094), .Z(n8859) );
  ANDN U7849 ( .B(n5096), .A(n8859), .Z(n12913) );
  NANDN U7850 ( .A(n5097), .B(n12913), .Z(n5098) );
  AND U7851 ( .A(n12917), .B(n5098), .Z(n5101) );
  NANDN U7852 ( .A(y[1519]), .B(x[1519]), .Z(n5100) );
  NANDN U7853 ( .A(y[1518]), .B(x[1518]), .Z(n5099) );
  NAND U7854 ( .A(n5100), .B(n5099), .Z(n8861) );
  NAND U7855 ( .A(n8861), .B(n8862), .Z(n12916) );
  NAND U7856 ( .A(n5101), .B(n12916), .Z(n5102) );
  NANDN U7857 ( .A(n12920), .B(n5102), .Z(n5103) );
  NANDN U7858 ( .A(y[1522]), .B(x[1522]), .Z(n8871) );
  NAND U7859 ( .A(n5103), .B(n8871), .Z(n5104) );
  NANDN U7860 ( .A(y[1521]), .B(x[1521]), .Z(n12922) );
  NANDN U7861 ( .A(n5104), .B(n12922), .Z(n5105) );
  AND U7862 ( .A(n12923), .B(n5105), .Z(n5106) );
  ANDN U7863 ( .B(n5107), .A(n5106), .Z(n5108) );
  AND U7864 ( .A(n8875), .B(n5108), .Z(n5111) );
  NANDN U7865 ( .A(x[1525]), .B(y[1525]), .Z(n5110) );
  NANDN U7866 ( .A(x[1526]), .B(y[1526]), .Z(n5109) );
  AND U7867 ( .A(n5110), .B(n5109), .Z(n12927) );
  NANDN U7868 ( .A(n5111), .B(n12927), .Z(n5114) );
  NANDN U7869 ( .A(y[1527]), .B(x[1527]), .Z(n5113) );
  NANDN U7870 ( .A(y[1526]), .B(x[1526]), .Z(n5112) );
  NAND U7871 ( .A(n5113), .B(n5112), .Z(n12930) );
  ANDN U7872 ( .B(n5114), .A(n12930), .Z(n5117) );
  NANDN U7873 ( .A(x[1527]), .B(y[1527]), .Z(n5116) );
  NANDN U7874 ( .A(x[1528]), .B(y[1528]), .Z(n5115) );
  AND U7875 ( .A(n5116), .B(n5115), .Z(n12931) );
  NANDN U7876 ( .A(n5117), .B(n12931), .Z(n5120) );
  NANDN U7877 ( .A(y[1528]), .B(x[1528]), .Z(n5119) );
  NANDN U7878 ( .A(y[1529]), .B(x[1529]), .Z(n5118) );
  AND U7879 ( .A(n5119), .B(n5118), .Z(n12933) );
  NAND U7880 ( .A(n5120), .B(n12933), .Z(n5121) );
  NANDN U7881 ( .A(x[1529]), .B(y[1529]), .Z(n6293) );
  NAND U7882 ( .A(n5121), .B(n6293), .Z(n5123) );
  NANDN U7883 ( .A(x[1530]), .B(n5123), .Z(n5122) );
  AND U7884 ( .A(n12940), .B(n5122), .Z(n5126) );
  IV U7885 ( .A(y[1530]), .Z(n6291) );
  XNOR U7886 ( .A(x[1530]), .B(n5123), .Z(n5124) );
  NANDN U7887 ( .A(n6291), .B(n5124), .Z(n5125) );
  NAND U7888 ( .A(n5126), .B(n5125), .Z(n5127) );
  NAND U7889 ( .A(n5128), .B(n5127), .Z(n5129) );
  ANDN U7890 ( .B(y[1533]), .A(x[1533]), .Z(n8893) );
  ANDN U7891 ( .B(y[1532]), .A(x[1532]), .Z(n8886) );
  NOR U7892 ( .A(n8893), .B(n8886), .Z(n12943) );
  NAND U7893 ( .A(n5129), .B(n12943), .Z(n5130) );
  ANDN U7894 ( .B(x[1534]), .A(y[1534]), .Z(n8895) );
  ANDN U7895 ( .B(n5130), .A(n8895), .Z(n5131) );
  NANDN U7896 ( .A(y[1533]), .B(x[1533]), .Z(n12945) );
  NAND U7897 ( .A(n5131), .B(n12945), .Z(n5132) );
  NANDN U7898 ( .A(x[1534]), .B(y[1534]), .Z(n12948) );
  NAND U7899 ( .A(n5132), .B(n12948), .Z(n5133) );
  ANDN U7900 ( .B(x[1535]), .A(y[1535]), .Z(n8894) );
  ANDN U7901 ( .B(n5133), .A(n8894), .Z(n5136) );
  NANDN U7902 ( .A(x[1536]), .B(y[1536]), .Z(n5135) );
  NANDN U7903 ( .A(x[1535]), .B(y[1535]), .Z(n5134) );
  NAND U7904 ( .A(n5135), .B(n5134), .Z(n12951) );
  OR U7905 ( .A(n5136), .B(n12951), .Z(n5137) );
  AND U7906 ( .A(n12953), .B(n5137), .Z(n5138) );
  OR U7907 ( .A(n12956), .B(n5138), .Z(n5141) );
  NANDN U7908 ( .A(y[1538]), .B(x[1538]), .Z(n5140) );
  NANDN U7909 ( .A(y[1539]), .B(x[1539]), .Z(n5139) );
  AND U7910 ( .A(n5140), .B(n5139), .Z(n12957) );
  NAND U7911 ( .A(n5141), .B(n12957), .Z(n5142) );
  NANDN U7912 ( .A(n12960), .B(n5142), .Z(n5143) );
  NAND U7913 ( .A(n5144), .B(n5143), .Z(n5145) );
  NANDN U7914 ( .A(n5146), .B(n5145), .Z(n5147) );
  NAND U7915 ( .A(n5148), .B(n5147), .Z(n5149) );
  AND U7916 ( .A(n8908), .B(n5149), .Z(n5150) );
  NANDN U7917 ( .A(x[1545]), .B(y[1545]), .Z(n6289) );
  NAND U7918 ( .A(n5150), .B(n6289), .Z(n5151) );
  AND U7919 ( .A(n12970), .B(n5151), .Z(n5152) );
  NAND U7920 ( .A(n5153), .B(n5152), .Z(n5154) );
  NAND U7921 ( .A(n5155), .B(n5154), .Z(n5156) );
  ANDN U7922 ( .B(x[1547]), .A(y[1547]), .Z(n8914) );
  ANDN U7923 ( .B(n5156), .A(n8914), .Z(n5157) );
  NAND U7924 ( .A(n5158), .B(n5157), .Z(n5159) );
  NAND U7925 ( .A(n5160), .B(n5159), .Z(n5161) );
  ANDN U7926 ( .B(x[1549]), .A(y[1549]), .Z(n8920) );
  ANDN U7927 ( .B(n5161), .A(n8920), .Z(n5162) );
  NAND U7928 ( .A(n5163), .B(n5162), .Z(n5164) );
  NAND U7929 ( .A(n6285), .B(n5164), .Z(n5165) );
  ANDN U7930 ( .B(x[1551]), .A(y[1551]), .Z(n8924) );
  ANDN U7931 ( .B(n5165), .A(n8924), .Z(n5166) );
  NANDN U7932 ( .A(x[1553]), .B(y[1553]), .Z(n5169) );
  ANDN U7933 ( .B(y[1551]), .A(x[1551]), .Z(n12989) );
  ANDN U7934 ( .B(n9996), .A(n12989), .Z(n8927) );
  NANDN U7935 ( .A(n5166), .B(n8927), .Z(n5167) );
  AND U7936 ( .A(n8933), .B(n5167), .Z(n5170) );
  NANDN U7937 ( .A(y[1552]), .B(x[1552]), .Z(n5168) );
  NANDN U7938 ( .A(y[1553]), .B(x[1553]), .Z(n9997) );
  NAND U7939 ( .A(n5168), .B(n9997), .Z(n12991) );
  NAND U7940 ( .A(n5169), .B(n12991), .Z(n8929) );
  NAND U7941 ( .A(n5170), .B(n8929), .Z(n5171) );
  NANDN U7942 ( .A(n5172), .B(n5171), .Z(n5173) );
  AND U7943 ( .A(n5174), .B(n5173), .Z(n5175) );
  ANDN U7944 ( .B(y[1556]), .A(x[1556]), .Z(n8935) );
  ANDN U7945 ( .B(y[1557]), .A(x[1557]), .Z(n8940) );
  NOR U7946 ( .A(n8935), .B(n8940), .Z(n13002) );
  NANDN U7947 ( .A(n5175), .B(n13002), .Z(n5176) );
  NAND U7948 ( .A(n5177), .B(n5176), .Z(n5178) );
  NANDN U7949 ( .A(n13007), .B(n5178), .Z(n5179) );
  NANDN U7950 ( .A(n5179), .B(x[1559]), .Z(n5182) );
  XNOR U7951 ( .A(n5179), .B(x[1559]), .Z(n5180) );
  NANDN U7952 ( .A(y[1559]), .B(n5180), .Z(n5181) );
  AND U7953 ( .A(n5182), .B(n5181), .Z(n5183) );
  OR U7954 ( .A(n5183), .B(y[1560]), .Z(n5186) );
  XOR U7955 ( .A(y[1560]), .B(n5183), .Z(n5184) );
  NAND U7956 ( .A(n5184), .B(x[1560]), .Z(n5185) );
  NAND U7957 ( .A(n5186), .B(n5185), .Z(n5187) );
  AND U7958 ( .A(n13014), .B(n5187), .Z(n5188) );
  ANDN U7959 ( .B(n8953), .A(n5188), .Z(n5189) );
  NANDN U7960 ( .A(y[1561]), .B(x[1561]), .Z(n8947) );
  NAND U7961 ( .A(n5189), .B(n8947), .Z(n5191) );
  NANDN U7962 ( .A(x[1565]), .B(y[1565]), .Z(n5194) );
  NANDN U7963 ( .A(x[1564]), .B(y[1564]), .Z(n5190) );
  NAND U7964 ( .A(n5194), .B(n5190), .Z(n13022) );
  ANDN U7965 ( .B(n5191), .A(n13022), .Z(n5193) );
  ANDN U7966 ( .B(y[1563]), .A(x[1563]), .Z(n8955) );
  NANDN U7967 ( .A(x[1562]), .B(y[1562]), .Z(n8951) );
  NANDN U7968 ( .A(n8955), .B(n8951), .Z(n13019) );
  NANDN U7969 ( .A(n9994), .B(n13019), .Z(n5192) );
  AND U7970 ( .A(n5193), .B(n5192), .Z(n5196) );
  ANDN U7971 ( .B(x[1565]), .A(y[1565]), .Z(n13025) );
  ANDN U7972 ( .B(x[1564]), .A(y[1564]), .Z(n9995) );
  NAND U7973 ( .A(n5194), .B(n9995), .Z(n5195) );
  NANDN U7974 ( .A(n13025), .B(n5195), .Z(n8959) );
  NOR U7975 ( .A(n5196), .B(n8959), .Z(n5197) );
  NANDN U7976 ( .A(n8961), .B(n5197), .Z(n5198) );
  NANDN U7977 ( .A(x[1566]), .B(y[1566]), .Z(n13026) );
  NAND U7978 ( .A(n5198), .B(n13026), .Z(n5199) );
  NANDN U7979 ( .A(x[1567]), .B(y[1567]), .Z(n13030) );
  NANDN U7980 ( .A(n5199), .B(n13030), .Z(n5200) );
  AND U7981 ( .A(n5201), .B(n5200), .Z(n5202) );
  ANDN U7982 ( .B(y[1568]), .A(x[1568]), .Z(n8966) );
  ANDN U7983 ( .B(y[1569]), .A(x[1569]), .Z(n8969) );
  NOR U7984 ( .A(n8966), .B(n8969), .Z(n13035) );
  NANDN U7985 ( .A(n5202), .B(n13035), .Z(n5203) );
  ANDN U7986 ( .B(x[1570]), .A(y[1570]), .Z(n8972) );
  ANDN U7987 ( .B(n5203), .A(n8972), .Z(n5204) );
  NANDN U7988 ( .A(y[1569]), .B(x[1569]), .Z(n13036) );
  NAND U7989 ( .A(n5204), .B(n13036), .Z(n5205) );
  AND U7990 ( .A(n13038), .B(n5205), .Z(n5206) );
  NAND U7991 ( .A(n5207), .B(n5206), .Z(n5208) );
  NAND U7992 ( .A(n5209), .B(n5208), .Z(n5210) );
  NANDN U7993 ( .A(x[1572]), .B(y[1572]), .Z(n6283) );
  AND U7994 ( .A(n5210), .B(n6283), .Z(n5211) );
  NAND U7995 ( .A(n5212), .B(n5211), .Z(n5213) );
  NAND U7996 ( .A(n5214), .B(n5213), .Z(n5215) );
  AND U7997 ( .A(n8977), .B(n5215), .Z(n5218) );
  NANDN U7998 ( .A(y[1574]), .B(x[1574]), .Z(n5217) );
  NANDN U7999 ( .A(y[1575]), .B(x[1575]), .Z(n5216) );
  AND U8000 ( .A(n5217), .B(n5216), .Z(n13048) );
  NANDN U8001 ( .A(n5218), .B(n13048), .Z(n5221) );
  NANDN U8002 ( .A(x[1576]), .B(y[1576]), .Z(n5220) );
  NANDN U8003 ( .A(x[1575]), .B(y[1575]), .Z(n5219) );
  NAND U8004 ( .A(n5220), .B(n5219), .Z(n13050) );
  ANDN U8005 ( .B(n5221), .A(n13050), .Z(n5224) );
  NANDN U8006 ( .A(y[1576]), .B(x[1576]), .Z(n5223) );
  NANDN U8007 ( .A(y[1577]), .B(x[1577]), .Z(n5222) );
  AND U8008 ( .A(n5223), .B(n5222), .Z(n13052) );
  NANDN U8009 ( .A(n5224), .B(n13052), .Z(n5225) );
  AND U8010 ( .A(n6277), .B(n5225), .Z(n5226) );
  NAND U8011 ( .A(n5227), .B(n5226), .Z(n5228) );
  NAND U8012 ( .A(n8985), .B(n5228), .Z(n5229) );
  AND U8013 ( .A(n13058), .B(n5229), .Z(n5231) );
  ANDN U8014 ( .B(x[1579]), .A(y[1579]), .Z(n8984) );
  ANDN U8015 ( .B(x[1580]), .A(y[1580]), .Z(n13061) );
  OR U8016 ( .A(n8984), .B(n13061), .Z(n5230) );
  OR U8017 ( .A(n5231), .B(n5230), .Z(n5232) );
  AND U8018 ( .A(n13062), .B(n5232), .Z(n5233) );
  ANDN U8019 ( .B(n13065), .A(n5233), .Z(n5234) );
  NANDN U8020 ( .A(y[1582]), .B(x[1582]), .Z(n8997) );
  NAND U8021 ( .A(n5234), .B(n8997), .Z(n5235) );
  AND U8022 ( .A(n13066), .B(n5235), .Z(n5236) );
  NAND U8023 ( .A(n5237), .B(n5236), .Z(n5238) );
  NAND U8024 ( .A(n5239), .B(n5238), .Z(n5240) );
  ANDN U8025 ( .B(y[1584]), .A(x[1584]), .Z(n8999) );
  ANDN U8026 ( .B(n5240), .A(n8999), .Z(n5241) );
  NAND U8027 ( .A(n5242), .B(n5241), .Z(n5243) );
  NAND U8028 ( .A(n6274), .B(n5243), .Z(n5244) );
  ANDN U8029 ( .B(y[1586]), .A(x[1586]), .Z(n9003) );
  ANDN U8030 ( .B(n5244), .A(n9003), .Z(n5245) );
  OR U8031 ( .A(n13077), .B(n5245), .Z(n5246) );
  AND U8032 ( .A(n13078), .B(n5246), .Z(n5247) );
  NANDN U8033 ( .A(y[1588]), .B(x[1588]), .Z(n13081) );
  NANDN U8034 ( .A(n5247), .B(n13081), .Z(n5248) );
  NANDN U8035 ( .A(n13083), .B(n5248), .Z(n5249) );
  NANDN U8036 ( .A(y[1590]), .B(x[1590]), .Z(n6271) );
  NAND U8037 ( .A(n5249), .B(n6271), .Z(n5250) );
  NANDN U8038 ( .A(y[1589]), .B(x[1589]), .Z(n13085) );
  NANDN U8039 ( .A(n5250), .B(n13085), .Z(n5252) );
  NANDN U8040 ( .A(x[1591]), .B(y[1591]), .Z(n6270) );
  NANDN U8041 ( .A(x[1590]), .B(y[1590]), .Z(n5251) );
  NAND U8042 ( .A(n6270), .B(n5251), .Z(n13087) );
  ANDN U8043 ( .B(n5252), .A(n13087), .Z(n5255) );
  NANDN U8044 ( .A(y[1592]), .B(x[1592]), .Z(n5254) );
  NANDN U8045 ( .A(y[1591]), .B(x[1591]), .Z(n5253) );
  AND U8046 ( .A(n5254), .B(n5253), .Z(n6272) );
  NANDN U8047 ( .A(n5255), .B(n6272), .Z(n5258) );
  NANDN U8048 ( .A(x[1593]), .B(y[1593]), .Z(n5257) );
  NANDN U8049 ( .A(x[1592]), .B(y[1592]), .Z(n5256) );
  NAND U8050 ( .A(n5257), .B(n5256), .Z(n13091) );
  ANDN U8051 ( .B(n5258), .A(n13091), .Z(n5260) );
  NANDN U8052 ( .A(y[1594]), .B(x[1594]), .Z(n9016) );
  NANDN U8053 ( .A(y[1593]), .B(x[1593]), .Z(n13092) );
  NAND U8054 ( .A(n9016), .B(n13092), .Z(n5259) );
  OR U8055 ( .A(n5260), .B(n5259), .Z(n5263) );
  ANDN U8056 ( .B(y[1596]), .A(x[1596]), .Z(n5264) );
  NANDN U8057 ( .A(x[1595]), .B(y[1595]), .Z(n5261) );
  NANDN U8058 ( .A(n5264), .B(n5261), .Z(n9019) );
  NANDN U8059 ( .A(x[1594]), .B(y[1594]), .Z(n5262) );
  NANDN U8060 ( .A(n9019), .B(n5262), .Z(n13095) );
  ANDN U8061 ( .B(n5263), .A(n13095), .Z(n5269) );
  ANDN U8062 ( .B(x[1595]), .A(y[1595]), .Z(n9017) );
  NANDN U8063 ( .A(n5264), .B(n9017), .Z(n5267) );
  NANDN U8064 ( .A(y[1596]), .B(x[1596]), .Z(n5266) );
  NANDN U8065 ( .A(y[1597]), .B(x[1597]), .Z(n5265) );
  NAND U8066 ( .A(n5266), .B(n5265), .Z(n9020) );
  ANDN U8067 ( .B(n5267), .A(n9020), .Z(n5268) );
  NANDN U8068 ( .A(n5269), .B(n5268), .Z(n5270) );
  NANDN U8069 ( .A(n13099), .B(n5270), .Z(n5271) );
  AND U8070 ( .A(n13100), .B(n5271), .Z(n5274) );
  NANDN U8071 ( .A(x[1600]), .B(y[1600]), .Z(n5273) );
  ANDN U8072 ( .B(n5273), .A(n5272), .Z(n13106) );
  ANDN U8073 ( .B(y[1599]), .A(x[1599]), .Z(n13103) );
  ANDN U8074 ( .B(n13106), .A(n13103), .Z(n9025) );
  NANDN U8075 ( .A(n5274), .B(n9025), .Z(n5275) );
  AND U8076 ( .A(n9027), .B(n5275), .Z(n5276) );
  NANDN U8077 ( .A(y[1602]), .B(x[1602]), .Z(n6266) );
  NAND U8078 ( .A(n5276), .B(n6266), .Z(n5278) );
  ANDN U8079 ( .B(y[1603]), .A(x[1603]), .Z(n6267) );
  NANDN U8080 ( .A(x[1602]), .B(y[1602]), .Z(n5277) );
  NANDN U8081 ( .A(n6267), .B(n5277), .Z(n13111) );
  ANDN U8082 ( .B(n5278), .A(n13111), .Z(n5281) );
  NANDN U8083 ( .A(y[1604]), .B(x[1604]), .Z(n5280) );
  NANDN U8084 ( .A(y[1603]), .B(x[1603]), .Z(n5279) );
  AND U8085 ( .A(n5280), .B(n5279), .Z(n6268) );
  NANDN U8086 ( .A(n5281), .B(n6268), .Z(n5282) );
  AND U8087 ( .A(n13114), .B(n5282), .Z(n5283) );
  OR U8088 ( .A(n13117), .B(n5283), .Z(n5284) );
  NANDN U8089 ( .A(n13119), .B(n5284), .Z(n5285) );
  NANDN U8090 ( .A(y[1607]), .B(x[1607]), .Z(n13121) );
  NAND U8091 ( .A(n5285), .B(n13121), .Z(n5286) );
  NANDN U8092 ( .A(y[1608]), .B(x[1608]), .Z(n6265) );
  NANDN U8093 ( .A(n5286), .B(n6265), .Z(n5288) );
  NANDN U8094 ( .A(x[1609]), .B(y[1609]), .Z(n13126) );
  ANDN U8095 ( .B(y[1608]), .A(x[1608]), .Z(n13123) );
  ANDN U8096 ( .B(n13126), .A(n13123), .Z(n5287) );
  NAND U8097 ( .A(n5288), .B(n5287), .Z(n5289) );
  NANDN U8098 ( .A(y[1609]), .B(x[1609]), .Z(n6264) );
  NAND U8099 ( .A(n5289), .B(n6264), .Z(n5290) );
  NANDN U8100 ( .A(y[1610]), .B(x[1610]), .Z(n13128) );
  NANDN U8101 ( .A(n5290), .B(n13128), .Z(n5291) );
  NANDN U8102 ( .A(x[1610]), .B(y[1610]), .Z(n9038) );
  NANDN U8103 ( .A(x[1611]), .B(y[1611]), .Z(n9043) );
  NAND U8104 ( .A(n9038), .B(n9043), .Z(n13131) );
  ANDN U8105 ( .B(n5291), .A(n13131), .Z(n5293) );
  ANDN U8106 ( .B(x[1612]), .A(y[1612]), .Z(n9045) );
  NANDN U8107 ( .A(y[1611]), .B(x[1611]), .Z(n13132) );
  NANDN U8108 ( .A(n9045), .B(n13132), .Z(n5292) );
  OR U8109 ( .A(n5293), .B(n5292), .Z(n5294) );
  AND U8110 ( .A(n5295), .B(n5294), .Z(n5297) );
  ANDN U8111 ( .B(x[1613]), .A(y[1613]), .Z(n9046) );
  NANDN U8112 ( .A(y[1614]), .B(x[1614]), .Z(n13140) );
  NANDN U8113 ( .A(n9046), .B(n13140), .Z(n5296) );
  OR U8114 ( .A(n5297), .B(n5296), .Z(n5298) );
  ANDN U8115 ( .B(y[1615]), .A(x[1615]), .Z(n6263) );
  NANDN U8116 ( .A(x[1614]), .B(y[1614]), .Z(n9049) );
  NANDN U8117 ( .A(n6263), .B(n9049), .Z(n13142) );
  ANDN U8118 ( .B(n5298), .A(n13142), .Z(n5299) );
  NANDN U8119 ( .A(y[1615]), .B(x[1615]), .Z(n13145) );
  NANDN U8120 ( .A(n5299), .B(n13145), .Z(n5302) );
  NANDN U8121 ( .A(x[1616]), .B(y[1616]), .Z(n5301) );
  ANDN U8122 ( .B(n5301), .A(n5300), .Z(n13149) );
  NAND U8123 ( .A(n5302), .B(n13149), .Z(n5303) );
  NANDN U8124 ( .A(n9056), .B(n5303), .Z(n5304) );
  NANDN U8125 ( .A(y[1618]), .B(x[1618]), .Z(n6262) );
  NANDN U8126 ( .A(n5304), .B(n6262), .Z(n5305) );
  NANDN U8127 ( .A(n13153), .B(n5305), .Z(n5306) );
  IV U8128 ( .A(x[1619]), .Z(n6260) );
  OR U8129 ( .A(n5306), .B(n6260), .Z(n5309) );
  XNOR U8130 ( .A(n5306), .B(x[1619]), .Z(n5307) );
  NANDN U8131 ( .A(y[1619]), .B(n5307), .Z(n5308) );
  NAND U8132 ( .A(n5309), .B(n5308), .Z(n5310) );
  NAND U8133 ( .A(n5311), .B(n5310), .Z(n5312) );
  NAND U8134 ( .A(n6259), .B(n5312), .Z(n5313) );
  NAND U8135 ( .A(n5314), .B(n5313), .Z(n5315) );
  NAND U8136 ( .A(n5316), .B(n5315), .Z(n5317) );
  ANDN U8137 ( .B(y[1622]), .A(x[1622]), .Z(n9063) );
  ANDN U8138 ( .B(n5317), .A(n9063), .Z(n5318) );
  NAND U8139 ( .A(n5319), .B(n5318), .Z(n5320) );
  NAND U8140 ( .A(n6254), .B(n5320), .Z(n5321) );
  AND U8141 ( .A(n13170), .B(n5321), .Z(n5322) );
  OR U8142 ( .A(n9069), .B(n5322), .Z(n5327) );
  NANDN U8143 ( .A(x[1627]), .B(y[1627]), .Z(n5324) );
  NANDN U8144 ( .A(x[1626]), .B(y[1626]), .Z(n5323) );
  NAND U8145 ( .A(n5324), .B(n5323), .Z(n13174) );
  ANDN U8146 ( .B(y[1625]), .A(x[1625]), .Z(n13168) );
  NANDN U8147 ( .A(n5325), .B(n13168), .Z(n5326) );
  NANDN U8148 ( .A(n13174), .B(n5326), .Z(n9072) );
  ANDN U8149 ( .B(n5327), .A(n9072), .Z(n5328) );
  ANDN U8150 ( .B(n13176), .A(n5328), .Z(n5329) );
  NANDN U8151 ( .A(y[1628]), .B(x[1628]), .Z(n6252) );
  NAND U8152 ( .A(n5329), .B(n6252), .Z(n5330) );
  AND U8153 ( .A(n13178), .B(n5330), .Z(n5331) );
  NANDN U8154 ( .A(y[1629]), .B(x[1629]), .Z(n6253) );
  NANDN U8155 ( .A(n5331), .B(n6253), .Z(n5332) );
  AND U8156 ( .A(n13182), .B(n5332), .Z(n5333) );
  OR U8157 ( .A(n13185), .B(n5333), .Z(n5334) );
  NANDN U8158 ( .A(n13187), .B(n5334), .Z(n5337) );
  NANDN U8159 ( .A(y[1632]), .B(x[1632]), .Z(n5336) );
  AND U8160 ( .A(n5336), .B(n5335), .Z(n13188) );
  NAND U8161 ( .A(n5337), .B(n13188), .Z(n5338) );
  NAND U8162 ( .A(n5339), .B(n5338), .Z(n5341) );
  NANDN U8163 ( .A(y[1634]), .B(x[1634]), .Z(n5340) );
  ANDN U8164 ( .B(x[1635]), .A(y[1635]), .Z(n5342) );
  ANDN U8165 ( .B(n5340), .A(n5342), .Z(n9085) );
  NAND U8166 ( .A(n5341), .B(n9085), .Z(n5344) );
  NANDN U8167 ( .A(x[1635]), .B(y[1635]), .Z(n9086) );
  NANDN U8168 ( .A(n5342), .B(n9082), .Z(n5343) );
  AND U8169 ( .A(n5344), .B(n5343), .Z(n5345) );
  NANDN U8170 ( .A(n13197), .B(n5345), .Z(n5346) );
  NANDN U8171 ( .A(n13198), .B(n5346), .Z(n5349) );
  NANDN U8172 ( .A(x[1639]), .B(y[1639]), .Z(n5348) );
  NANDN U8173 ( .A(x[1638]), .B(y[1638]), .Z(n5347) );
  NAND U8174 ( .A(n5348), .B(n5347), .Z(n13201) );
  ANDN U8175 ( .B(n5349), .A(n13201), .Z(n5352) );
  NANDN U8176 ( .A(y[1639]), .B(x[1639]), .Z(n5351) );
  NANDN U8177 ( .A(y[1640]), .B(x[1640]), .Z(n5350) );
  AND U8178 ( .A(n5351), .B(n5350), .Z(n13203) );
  NANDN U8179 ( .A(n5352), .B(n13203), .Z(n5353) );
  ANDN U8180 ( .B(y[1641]), .A(x[1641]), .Z(n9099) );
  ANDN U8181 ( .B(n5353), .A(n9099), .Z(n5354) );
  NANDN U8182 ( .A(x[1640]), .B(y[1640]), .Z(n13204) );
  NAND U8183 ( .A(n5354), .B(n13204), .Z(n5355) );
  AND U8184 ( .A(n13206), .B(n5355), .Z(n5356) );
  NAND U8185 ( .A(n5357), .B(n5356), .Z(n5358) );
  NAND U8186 ( .A(n5359), .B(n5358), .Z(n5360) );
  NAND U8187 ( .A(n5361), .B(n5360), .Z(n5363) );
  IV U8188 ( .A(y[1645]), .Z(n6251) );
  IV U8189 ( .A(x[1645]), .Z(n6250) );
  NANDN U8190 ( .A(n6251), .B(n6250), .Z(n5362) );
  ANDN U8191 ( .B(y[1644]), .A(x[1644]), .Z(n9107) );
  ANDN U8192 ( .B(n5362), .A(n9107), .Z(n13216) );
  NAND U8193 ( .A(n5363), .B(n13216), .Z(n5365) );
  NANDN U8194 ( .A(y[1645]), .B(x[1645]), .Z(n5364) );
  NANDN U8195 ( .A(y[1646]), .B(x[1646]), .Z(n9114) );
  NAND U8196 ( .A(n5364), .B(n9114), .Z(n13219) );
  ANDN U8197 ( .B(n5365), .A(n13219), .Z(n5366) );
  NANDN U8198 ( .A(x[1647]), .B(y[1647]), .Z(n9117) );
  NANDN U8199 ( .A(x[1646]), .B(y[1646]), .Z(n6249) );
  NAND U8200 ( .A(n9117), .B(n6249), .Z(n13221) );
  OR U8201 ( .A(n5366), .B(n13221), .Z(n5367) );
  ANDN U8202 ( .B(x[1648]), .A(y[1648]), .Z(n6246) );
  ANDN U8203 ( .B(n5367), .A(n6246), .Z(n5368) );
  NANDN U8204 ( .A(y[1647]), .B(x[1647]), .Z(n13222) );
  NAND U8205 ( .A(n5368), .B(n13222), .Z(n5369) );
  NANDN U8206 ( .A(x[1648]), .B(y[1648]), .Z(n13225) );
  AND U8207 ( .A(n5369), .B(n13225), .Z(n5370) );
  OR U8208 ( .A(n5370), .B(x[1649]), .Z(n5373) );
  XOR U8209 ( .A(x[1649]), .B(n5370), .Z(n5371) );
  NAND U8210 ( .A(n5371), .B(y[1649]), .Z(n5372) );
  NAND U8211 ( .A(n5373), .B(n5372), .Z(n5374) );
  ANDN U8212 ( .B(x[1650]), .A(y[1650]), .Z(n13231) );
  ANDN U8213 ( .B(n5374), .A(n13231), .Z(n5376) );
  NANDN U8214 ( .A(x[1650]), .B(y[1650]), .Z(n6244) );
  NANDN U8215 ( .A(x[1651]), .B(y[1651]), .Z(n13232) );
  NAND U8216 ( .A(n6244), .B(n13232), .Z(n5375) );
  OR U8217 ( .A(n5376), .B(n5375), .Z(n5377) );
  NANDN U8218 ( .A(y[1651]), .B(x[1651]), .Z(n6243) );
  ANDN U8219 ( .B(n5377), .A(n13235), .Z(n5378) );
  OR U8220 ( .A(n13236), .B(n5378), .Z(n5380) );
  NANDN U8221 ( .A(y[1653]), .B(x[1653]), .Z(n5379) );
  ANDN U8222 ( .B(x[1654]), .A(y[1654]), .Z(n9132) );
  ANDN U8223 ( .B(n5379), .A(n9132), .Z(n13238) );
  NAND U8224 ( .A(n5380), .B(n13238), .Z(n5383) );
  NANDN U8225 ( .A(x[1654]), .B(y[1654]), .Z(n5382) );
  NANDN U8226 ( .A(x[1655]), .B(y[1655]), .Z(n5381) );
  AND U8227 ( .A(n5382), .B(n5381), .Z(n13241) );
  NAND U8228 ( .A(n5383), .B(n13241), .Z(n5384) );
  NANDN U8229 ( .A(n13243), .B(n5384), .Z(n5387) );
  NANDN U8230 ( .A(x[1656]), .B(y[1656]), .Z(n5386) );
  NANDN U8231 ( .A(x[1657]), .B(y[1657]), .Z(n5385) );
  AND U8232 ( .A(n5386), .B(n5385), .Z(n13244) );
  NAND U8233 ( .A(n5387), .B(n13244), .Z(n5388) );
  AND U8234 ( .A(n13248), .B(n5388), .Z(n5390) );
  NANDN U8235 ( .A(x[1658]), .B(y[1658]), .Z(n5389) );
  ANDN U8236 ( .B(y[1659]), .A(x[1659]), .Z(n5393) );
  ANDN U8237 ( .B(n5389), .A(n5393), .Z(n13250) );
  NANDN U8238 ( .A(n5390), .B(n13250), .Z(n5395) );
  NANDN U8239 ( .A(y[1660]), .B(x[1660]), .Z(n5392) );
  NANDN U8240 ( .A(y[1659]), .B(x[1659]), .Z(n5391) );
  NAND U8241 ( .A(n5392), .B(n5391), .Z(n13252) );
  ANDN U8242 ( .B(x[1658]), .A(y[1658]), .Z(n13247) );
  NANDN U8243 ( .A(n5393), .B(n13247), .Z(n5394) );
  NANDN U8244 ( .A(n13252), .B(n5394), .Z(n9140) );
  ANDN U8245 ( .B(n5395), .A(n9140), .Z(n5396) );
  OR U8246 ( .A(n13255), .B(n5396), .Z(n5397) );
  AND U8247 ( .A(n5398), .B(n5397), .Z(n5399) );
  NANDN U8248 ( .A(x[1662]), .B(y[1662]), .Z(n13258) );
  NANDN U8249 ( .A(n5399), .B(n13258), .Z(n5400) );
  NANDN U8250 ( .A(n9144), .B(n5400), .Z(n5404) );
  NANDN U8251 ( .A(x[1663]), .B(y[1663]), .Z(n5402) );
  NANDN U8252 ( .A(x[1664]), .B(y[1664]), .Z(n5401) );
  NAND U8253 ( .A(n5402), .B(n5401), .Z(n9148) );
  ANDN U8254 ( .B(n5403), .A(n9148), .Z(n13262) );
  NAND U8255 ( .A(n5404), .B(n13262), .Z(n5405) );
  NANDN U8256 ( .A(n13264), .B(n5405), .Z(n5406) );
  NANDN U8257 ( .A(n13267), .B(n5406), .Z(n5408) );
  NANDN U8258 ( .A(y[1667]), .B(x[1667]), .Z(n5407) );
  NANDN U8259 ( .A(y[1668]), .B(x[1668]), .Z(n9162) );
  NAND U8260 ( .A(n5407), .B(n9162), .Z(n13268) );
  ANDN U8261 ( .B(n5408), .A(n13268), .Z(n5409) );
  ANDN U8262 ( .B(n6235), .A(n5409), .Z(n5410) );
  NANDN U8263 ( .A(x[1668]), .B(y[1668]), .Z(n13270) );
  NAND U8264 ( .A(n5410), .B(n13270), .Z(n5411) );
  NANDN U8265 ( .A(n13273), .B(n5411), .Z(n5418) );
  ANDN U8266 ( .B(y[1670]), .A(x[1670]), .Z(n6236) );
  NANDN U8267 ( .A(n6236), .B(n5412), .Z(n5416) );
  XOR U8268 ( .A(y[1671]), .B(n6236), .Z(n5413) );
  NANDN U8269 ( .A(n5414), .B(n5413), .Z(n5415) );
  NAND U8270 ( .A(n5416), .B(n5415), .Z(n5417) );
  AND U8271 ( .A(n5418), .B(n5417), .Z(n5419) );
  NANDN U8272 ( .A(y[1672]), .B(x[1672]), .Z(n13276) );
  NANDN U8273 ( .A(n5419), .B(n13276), .Z(n5420) );
  IV U8274 ( .A(y[1673]), .Z(n6234) );
  NANDN U8275 ( .A(x[1672]), .B(y[1672]), .Z(n9165) );
  NAND U8276 ( .A(n6233), .B(n9165), .Z(n13279) );
  ANDN U8277 ( .B(n5420), .A(n13279), .Z(n5421) );
  OR U8278 ( .A(n13280), .B(n5421), .Z(n5422) );
  ANDN U8279 ( .B(y[1674]), .A(x[1674]), .Z(n6232) );
  ANDN U8280 ( .B(y[1675]), .A(x[1675]), .Z(n9177) );
  NOR U8281 ( .A(n6232), .B(n9177), .Z(n13282) );
  NAND U8282 ( .A(n5422), .B(n13282), .Z(n5423) );
  NANDN U8283 ( .A(y[1676]), .B(x[1676]), .Z(n9179) );
  NAND U8284 ( .A(n5423), .B(n9179), .Z(n5424) );
  NANDN U8285 ( .A(y[1675]), .B(x[1675]), .Z(n13285) );
  NANDN U8286 ( .A(n5424), .B(n13285), .Z(n5425) );
  AND U8287 ( .A(n13290), .B(n5425), .Z(n5426) );
  NANDN U8288 ( .A(x[1676]), .B(y[1676]), .Z(n13286) );
  NAND U8289 ( .A(n5426), .B(n13286), .Z(n5430) );
  ANDN U8290 ( .B(x[1678]), .A(y[1678]), .Z(n13293) );
  ANDN U8291 ( .B(x[1679]), .A(y[1679]), .Z(n13296) );
  NOR U8292 ( .A(n13293), .B(n13296), .Z(n9182) );
  ANDN U8293 ( .B(x[1677]), .A(y[1677]), .Z(n9178) );
  NANDN U8294 ( .A(n5427), .B(n9178), .Z(n5428) );
  AND U8295 ( .A(n9182), .B(n5428), .Z(n5429) );
  NAND U8296 ( .A(n5430), .B(n5429), .Z(n5431) );
  NANDN U8297 ( .A(x[1679]), .B(y[1679]), .Z(n13295) );
  NAND U8298 ( .A(n5431), .B(n13295), .Z(n5432) );
  NANDN U8299 ( .A(y[1680]), .B(x[1680]), .Z(n13297) );
  NAND U8300 ( .A(n5432), .B(n13297), .Z(n5433) );
  ANDN U8301 ( .B(y[1681]), .A(x[1681]), .Z(n9190) );
  ANDN U8302 ( .B(y[1680]), .A(x[1680]), .Z(n9186) );
  NOR U8303 ( .A(n9190), .B(n9186), .Z(n13301) );
  NAND U8304 ( .A(n5433), .B(n13301), .Z(n5435) );
  IV U8305 ( .A(x[1682]), .Z(n6231) );
  IV U8306 ( .A(y[1682]), .Z(n6230) );
  NANDN U8307 ( .A(n6231), .B(n6230), .Z(n5434) );
  NANDN U8308 ( .A(y[1681]), .B(x[1681]), .Z(n9188) );
  NAND U8309 ( .A(n5434), .B(n9188), .Z(n13303) );
  ANDN U8310 ( .B(n5435), .A(n13303), .Z(n5437) );
  NANDN U8311 ( .A(x[1682]), .B(y[1682]), .Z(n5436) );
  ANDN U8312 ( .B(y[1683]), .A(x[1683]), .Z(n9196) );
  ANDN U8313 ( .B(n5436), .A(n9196), .Z(n13304) );
  NANDN U8314 ( .A(n5437), .B(n13304), .Z(n5438) );
  NANDN U8315 ( .A(n13307), .B(n5438), .Z(n5440) );
  NANDN U8316 ( .A(x[1684]), .B(y[1684]), .Z(n5439) );
  ANDN U8317 ( .B(y[1685]), .A(x[1685]), .Z(n9202) );
  ANDN U8318 ( .B(n5439), .A(n9202), .Z(n13308) );
  NAND U8319 ( .A(n5440), .B(n13308), .Z(n5441) );
  NANDN U8320 ( .A(n13311), .B(n5441), .Z(n5442) );
  NANDN U8321 ( .A(n13312), .B(n5442), .Z(n5443) );
  NANDN U8322 ( .A(n13315), .B(n5443), .Z(n5444) );
  NANDN U8323 ( .A(n13317), .B(n5444), .Z(n5445) );
  AND U8324 ( .A(n13318), .B(n5445), .Z(n5446) );
  NANDN U8325 ( .A(y[1690]), .B(x[1690]), .Z(n6218) );
  NAND U8326 ( .A(n5446), .B(n6218), .Z(n5447) );
  NANDN U8327 ( .A(n13321), .B(n5447), .Z(n5448) );
  IV U8328 ( .A(x[1691]), .Z(n6216) );
  OR U8329 ( .A(n5448), .B(n6216), .Z(n5451) );
  XNOR U8330 ( .A(n5448), .B(x[1691]), .Z(n5449) );
  NANDN U8331 ( .A(y[1691]), .B(n5449), .Z(n5450) );
  NAND U8332 ( .A(n5451), .B(n5450), .Z(n5452) );
  NANDN U8333 ( .A(y[1692]), .B(x[1692]), .Z(n13326) );
  NANDN U8334 ( .A(n5452), .B(n13326), .Z(n5453) );
  AND U8335 ( .A(n5454), .B(n5453), .Z(n5455) );
  ANDN U8336 ( .B(x[1694]), .A(y[1694]), .Z(n9227) );
  ANDN U8337 ( .B(x[1693]), .A(y[1693]), .Z(n9221) );
  NOR U8338 ( .A(n9227), .B(n9221), .Z(n13330) );
  NANDN U8339 ( .A(n5455), .B(n13330), .Z(n5456) );
  NANDN U8340 ( .A(n13333), .B(n5456), .Z(n5458) );
  NANDN U8341 ( .A(y[1695]), .B(x[1695]), .Z(n5457) );
  ANDN U8342 ( .B(x[1696]), .A(y[1696]), .Z(n9236) );
  ANDN U8343 ( .B(n5457), .A(n9236), .Z(n13335) );
  NAND U8344 ( .A(n5458), .B(n13335), .Z(n5459) );
  NAND U8345 ( .A(n5460), .B(n5459), .Z(n5461) );
  ANDN U8346 ( .B(x[1698]), .A(y[1698]), .Z(n13343) );
  NANDN U8347 ( .A(y[1697]), .B(x[1697]), .Z(n9233) );
  NANDN U8348 ( .A(n13343), .B(n9233), .Z(n13339) );
  ANDN U8349 ( .B(n5461), .A(n13339), .Z(n5462) );
  ANDN U8350 ( .B(n13340), .A(n5462), .Z(n5463) );
  NANDN U8351 ( .A(x[1698]), .B(y[1698]), .Z(n9238) );
  NAND U8352 ( .A(n5463), .B(n9238), .Z(n5465) );
  NANDN U8353 ( .A(y[1700]), .B(x[1700]), .Z(n5464) );
  NANDN U8354 ( .A(y[1699]), .B(x[1699]), .Z(n9241) );
  NAND U8355 ( .A(n5464), .B(n9241), .Z(n13346) );
  ANDN U8356 ( .B(n5465), .A(n13346), .Z(n5466) );
  OR U8357 ( .A(n13349), .B(n5466), .Z(n5467) );
  NANDN U8358 ( .A(n13351), .B(n5467), .Z(n5469) );
  NANDN U8359 ( .A(x[1702]), .B(y[1702]), .Z(n5468) );
  ANDN U8360 ( .B(y[1703]), .A(x[1703]), .Z(n9259) );
  ANDN U8361 ( .B(n5468), .A(n9259), .Z(n13352) );
  NAND U8362 ( .A(n5469), .B(n13352), .Z(n5470) );
  NAND U8363 ( .A(n5471), .B(n5470), .Z(n5472) );
  NANDN U8364 ( .A(x[1705]), .B(y[1705]), .Z(n6207) );
  ANDN U8365 ( .B(y[1704]), .A(x[1704]), .Z(n9256) );
  ANDN U8366 ( .B(n6207), .A(n9256), .Z(n13356) );
  NAND U8367 ( .A(n5472), .B(n13356), .Z(n5473) );
  NAND U8368 ( .A(n5474), .B(n5473), .Z(n5476) );
  IV U8369 ( .A(y[1707]), .Z(n9266) );
  OR U8370 ( .A(x[1707]), .B(n9266), .Z(n5475) );
  ANDN U8371 ( .B(y[1706]), .A(x[1706]), .Z(n6208) );
  ANDN U8372 ( .B(n5475), .A(n6208), .Z(n13362) );
  NAND U8373 ( .A(n5476), .B(n13362), .Z(n5477) );
  NANDN U8374 ( .A(n13365), .B(n5477), .Z(n5478) );
  NANDN U8375 ( .A(x[1708]), .B(y[1708]), .Z(n13367) );
  NAND U8376 ( .A(n5478), .B(n13367), .Z(n5480) );
  NANDN U8377 ( .A(y[1709]), .B(x[1709]), .Z(n5479) );
  ANDN U8378 ( .B(x[1710]), .A(y[1710]), .Z(n5481) );
  ANDN U8379 ( .B(n5479), .A(n5481), .Z(n13370) );
  NAND U8380 ( .A(n5480), .B(n13370), .Z(n5483) );
  ANDN U8381 ( .B(y[1710]), .A(x[1710]), .Z(n13373) );
  ANDN U8382 ( .B(y[1709]), .A(x[1709]), .Z(n13369) );
  NANDN U8383 ( .A(n5481), .B(n13369), .Z(n5482) );
  NANDN U8384 ( .A(n13373), .B(n5482), .Z(n9275) );
  ANDN U8385 ( .B(n5483), .A(n9275), .Z(n5484) );
  NANDN U8386 ( .A(y[1711]), .B(x[1711]), .Z(n13375) );
  NANDN U8387 ( .A(n5484), .B(n13375), .Z(n5485) );
  NANDN U8388 ( .A(n13377), .B(n5485), .Z(n5488) );
  NANDN U8389 ( .A(y[1712]), .B(x[1712]), .Z(n5487) );
  NANDN U8390 ( .A(y[1713]), .B(x[1713]), .Z(n5486) );
  AND U8391 ( .A(n5487), .B(n5486), .Z(n13379) );
  NAND U8392 ( .A(n5488), .B(n13379), .Z(n5489) );
  NANDN U8393 ( .A(n13381), .B(n5489), .Z(n5490) );
  NANDN U8394 ( .A(n9282), .B(n5490), .Z(n5491) );
  AND U8395 ( .A(n13384), .B(n5491), .Z(n5492) );
  NANDN U8396 ( .A(y[1716]), .B(x[1716]), .Z(n13388) );
  NANDN U8397 ( .A(n5492), .B(n13388), .Z(n5493) );
  AND U8398 ( .A(n13390), .B(n5493), .Z(n5494) );
  ANDN U8399 ( .B(n13392), .A(n5494), .Z(n5495) );
  NANDN U8400 ( .A(y[1718]), .B(x[1718]), .Z(n6206) );
  NAND U8401 ( .A(n5495), .B(n6206), .Z(n5496) );
  NANDN U8402 ( .A(x[1718]), .B(y[1718]), .Z(n13394) );
  NAND U8403 ( .A(n5496), .B(n13394), .Z(n5497) );
  IV U8404 ( .A(x[1719]), .Z(n6204) );
  OR U8405 ( .A(n5497), .B(n6204), .Z(n5500) );
  XNOR U8406 ( .A(n5497), .B(x[1719]), .Z(n5498) );
  NANDN U8407 ( .A(y[1719]), .B(n5498), .Z(n5499) );
  NAND U8408 ( .A(n5500), .B(n5499), .Z(n5501) );
  NANDN U8409 ( .A(y[1720]), .B(x[1720]), .Z(n13400) );
  NANDN U8410 ( .A(n5501), .B(n13400), .Z(n5503) );
  NANDN U8411 ( .A(x[1721]), .B(y[1721]), .Z(n13402) );
  NANDN U8412 ( .A(x[1720]), .B(y[1720]), .Z(n9289) );
  AND U8413 ( .A(n13402), .B(n9289), .Z(n5502) );
  NAND U8414 ( .A(n5503), .B(n5502), .Z(n5504) );
  NANDN U8415 ( .A(y[1721]), .B(x[1721]), .Z(n9292) );
  XOR U8416 ( .A(x[1722]), .B(y[1722]), .Z(n9296) );
  ANDN U8417 ( .B(n9292), .A(n9296), .Z(n13404) );
  NAND U8418 ( .A(n5504), .B(n13404), .Z(n5505) );
  NANDN U8419 ( .A(n13407), .B(n5505), .Z(n5506) );
  NANDN U8420 ( .A(n13409), .B(n5506), .Z(n5508) );
  IV U8421 ( .A(y[1725]), .Z(n9304) );
  OR U8422 ( .A(x[1725]), .B(n9304), .Z(n5507) );
  NANDN U8423 ( .A(x[1724]), .B(y[1724]), .Z(n9301) );
  NAND U8424 ( .A(n5507), .B(n9301), .Z(n13410) );
  ANDN U8425 ( .B(n5508), .A(n13410), .Z(n5510) );
  NANDN U8426 ( .A(y[1725]), .B(x[1725]), .Z(n5509) );
  ANDN U8427 ( .B(x[1726]), .A(y[1726]), .Z(n9307) );
  ANDN U8428 ( .B(n5509), .A(n9307), .Z(n13413) );
  NANDN U8429 ( .A(n5510), .B(n13413), .Z(n5511) );
  AND U8430 ( .A(n13414), .B(n5511), .Z(n5512) );
  OR U8431 ( .A(n13417), .B(n5512), .Z(n5515) );
  NANDN U8432 ( .A(x[1728]), .B(y[1728]), .Z(n5514) );
  NANDN U8433 ( .A(x[1729]), .B(y[1729]), .Z(n5513) );
  AND U8434 ( .A(n5514), .B(n5513), .Z(n13418) );
  NAND U8435 ( .A(n5515), .B(n13418), .Z(n5516) );
  NANDN U8436 ( .A(y[1730]), .B(x[1730]), .Z(n6201) );
  ANDN U8437 ( .B(x[1729]), .A(y[1729]), .Z(n9313) );
  ANDN U8438 ( .B(n6201), .A(n9313), .Z(n13420) );
  NAND U8439 ( .A(n5516), .B(n13420), .Z(n5518) );
  NANDN U8440 ( .A(x[1730]), .B(y[1730]), .Z(n5517) );
  ANDN U8441 ( .B(y[1731]), .A(x[1731]), .Z(n6203) );
  ANDN U8442 ( .B(n5517), .A(n6203), .Z(n13422) );
  NAND U8443 ( .A(n5518), .B(n13422), .Z(n5519) );
  AND U8444 ( .A(n13423), .B(n5519), .Z(n5520) );
  NANDN U8445 ( .A(y[1732]), .B(x[1732]), .Z(n6200) );
  NAND U8446 ( .A(n5520), .B(n6200), .Z(n5521) );
  NANDN U8447 ( .A(n13424), .B(n5521), .Z(n5522) );
  IV U8448 ( .A(x[1733]), .Z(n6198) );
  OR U8449 ( .A(n5522), .B(n6198), .Z(n5525) );
  XNOR U8450 ( .A(n5522), .B(x[1733]), .Z(n5523) );
  NANDN U8451 ( .A(y[1733]), .B(n5523), .Z(n5524) );
  NAND U8452 ( .A(n5525), .B(n5524), .Z(n5526) );
  NANDN U8453 ( .A(y[1734]), .B(x[1734]), .Z(n13427) );
  NANDN U8454 ( .A(n5526), .B(n13427), .Z(n5527) );
  AND U8455 ( .A(n9319), .B(n5527), .Z(n5528) );
  NANDN U8456 ( .A(x[1735]), .B(y[1735]), .Z(n13428) );
  NAND U8457 ( .A(n5528), .B(n13428), .Z(n5530) );
  NANDN U8458 ( .A(y[1735]), .B(x[1735]), .Z(n9322) );
  NANDN U8459 ( .A(y[1736]), .B(x[1736]), .Z(n5529) );
  NAND U8460 ( .A(n9322), .B(n5529), .Z(n13429) );
  ANDN U8461 ( .B(n5530), .A(n13429), .Z(n5531) );
  OR U8462 ( .A(n13430), .B(n5531), .Z(n5532) );
  NANDN U8463 ( .A(n13431), .B(n5532), .Z(n5533) );
  NANDN U8464 ( .A(x[1739]), .B(y[1739]), .Z(n9340) );
  NAND U8465 ( .A(n5533), .B(n9340), .Z(n5534) );
  NANDN U8466 ( .A(x[1738]), .B(y[1738]), .Z(n13432) );
  NANDN U8467 ( .A(n5534), .B(n13432), .Z(n5535) );
  AND U8468 ( .A(n13433), .B(n5535), .Z(n5537) );
  NANDN U8469 ( .A(x[1740]), .B(y[1740]), .Z(n5536) );
  ANDN U8470 ( .B(y[1741]), .A(x[1741]), .Z(n9345) );
  ANDN U8471 ( .B(n5536), .A(n9345), .Z(n13434) );
  NANDN U8472 ( .A(n5537), .B(n13434), .Z(n5540) );
  XNOR U8473 ( .A(x[1742]), .B(y[1742]), .Z(n5539) );
  NANDN U8474 ( .A(y[1741]), .B(x[1741]), .Z(n5538) );
  AND U8475 ( .A(n5539), .B(n5538), .Z(n13435) );
  NAND U8476 ( .A(n5540), .B(n13435), .Z(n5541) );
  NANDN U8477 ( .A(n13436), .B(n5541), .Z(n5542) );
  NANDN U8478 ( .A(n13437), .B(n5542), .Z(n5545) );
  NANDN U8479 ( .A(x[1745]), .B(y[1745]), .Z(n5544) );
  NANDN U8480 ( .A(x[1744]), .B(y[1744]), .Z(n5543) );
  AND U8481 ( .A(n5544), .B(n5543), .Z(n13439) );
  NAND U8482 ( .A(n5545), .B(n13439), .Z(n5546) );
  NANDN U8483 ( .A(y[1746]), .B(x[1746]), .Z(n9354) );
  NAND U8484 ( .A(n5546), .B(n9354), .Z(n5547) );
  NANDN U8485 ( .A(y[1745]), .B(x[1745]), .Z(n13440) );
  NANDN U8486 ( .A(n5547), .B(n13440), .Z(n5548) );
  AND U8487 ( .A(n6197), .B(n5548), .Z(n5549) );
  NANDN U8488 ( .A(x[1746]), .B(y[1746]), .Z(n13442) );
  NAND U8489 ( .A(n5549), .B(n13442), .Z(n5550) );
  AND U8490 ( .A(n9353), .B(n5550), .Z(n5551) );
  NANDN U8491 ( .A(y[1748]), .B(x[1748]), .Z(n13448) );
  NAND U8492 ( .A(n5551), .B(n13448), .Z(n5552) );
  NAND U8493 ( .A(n5553), .B(n5552), .Z(n5554) );
  NANDN U8494 ( .A(y[1749]), .B(x[1749]), .Z(n6195) );
  ANDN U8495 ( .B(x[1750]), .A(y[1750]), .Z(n9361) );
  ANDN U8496 ( .B(n6195), .A(n9361), .Z(n13452) );
  NAND U8497 ( .A(n5554), .B(n13452), .Z(n5555) );
  NANDN U8498 ( .A(x[1750]), .B(y[1750]), .Z(n13456) );
  NAND U8499 ( .A(n5555), .B(n13456), .Z(n5556) );
  AND U8500 ( .A(n13459), .B(n5556), .Z(n5557) );
  ANDN U8501 ( .B(y[1751]), .A(x[1751]), .Z(n13454) );
  ANDN U8502 ( .B(y[1752]), .A(x[1752]), .Z(n13464) );
  NOR U8503 ( .A(n13454), .B(n13464), .Z(n9364) );
  NANDN U8504 ( .A(n5557), .B(n9364), .Z(n5558) );
  NANDN U8505 ( .A(n9366), .B(n5558), .Z(n5559) );
  NANDN U8506 ( .A(x[1753]), .B(y[1753]), .Z(n6194) );
  NAND U8507 ( .A(n5559), .B(n6194), .Z(n5560) );
  NANDN U8508 ( .A(n13465), .B(n5560), .Z(n5561) );
  IV U8509 ( .A(y[1754]), .Z(n6192) );
  OR U8510 ( .A(n5561), .B(n6192), .Z(n5564) );
  XNOR U8511 ( .A(n5561), .B(y[1754]), .Z(n5562) );
  NANDN U8512 ( .A(x[1754]), .B(n5562), .Z(n5563) );
  NAND U8513 ( .A(n5564), .B(n5563), .Z(n5565) );
  NANDN U8514 ( .A(x[1755]), .B(y[1755]), .Z(n13470) );
  NANDN U8515 ( .A(n5565), .B(n13470), .Z(n5566) );
  ANDN U8516 ( .B(x[1755]), .A(y[1755]), .Z(n9370) );
  ANDN U8517 ( .B(n5566), .A(n9370), .Z(n5567) );
  NANDN U8518 ( .A(y[1756]), .B(x[1756]), .Z(n13472) );
  NAND U8519 ( .A(n5567), .B(n13472), .Z(n5569) );
  IV U8520 ( .A(y[1757]), .Z(n6191) );
  IV U8521 ( .A(x[1757]), .Z(n6190) );
  NANDN U8522 ( .A(n6191), .B(n6190), .Z(n5568) );
  ANDN U8523 ( .B(y[1756]), .A(x[1756]), .Z(n9375) );
  ANDN U8524 ( .B(n5568), .A(n9375), .Z(n13474) );
  NAND U8525 ( .A(n5569), .B(n13474), .Z(n5570) );
  AND U8526 ( .A(n13476), .B(n5570), .Z(n5571) );
  NANDN U8527 ( .A(x[1758]), .B(y[1758]), .Z(n6189) );
  NANDN U8528 ( .A(x[1759]), .B(y[1759]), .Z(n9385) );
  NAND U8529 ( .A(n6189), .B(n9385), .Z(n13478) );
  OR U8530 ( .A(n5571), .B(n13478), .Z(n5572) );
  ANDN U8531 ( .B(x[1760]), .A(y[1760]), .Z(n6186) );
  ANDN U8532 ( .B(n5572), .A(n6186), .Z(n5573) );
  NANDN U8533 ( .A(y[1759]), .B(x[1759]), .Z(n13480) );
  NAND U8534 ( .A(n5573), .B(n13480), .Z(n5574) );
  AND U8535 ( .A(n6185), .B(n5574), .Z(n5575) );
  NANDN U8536 ( .A(x[1760]), .B(y[1760]), .Z(n13482) );
  NAND U8537 ( .A(n5575), .B(n13482), .Z(n5576) );
  NAND U8538 ( .A(n5577), .B(n5576), .Z(n5578) );
  NANDN U8539 ( .A(x[1762]), .B(y[1762]), .Z(n6184) );
  NAND U8540 ( .A(n5578), .B(n6184), .Z(n5579) );
  NANDN U8541 ( .A(x[1763]), .B(y[1763]), .Z(n13490) );
  NANDN U8542 ( .A(n5579), .B(n13490), .Z(n5581) );
  XNOR U8543 ( .A(x[1764]), .B(y[1764]), .Z(n5580) );
  ANDN U8544 ( .B(x[1763]), .A(y[1763]), .Z(n6183) );
  ANDN U8545 ( .B(n5580), .A(n6183), .Z(n13492) );
  NAND U8546 ( .A(n5581), .B(n13492), .Z(n5582) );
  AND U8547 ( .A(n13494), .B(n5582), .Z(n5583) );
  OR U8548 ( .A(n13496), .B(n5583), .Z(n5585) );
  NANDN U8549 ( .A(x[1766]), .B(y[1766]), .Z(n5584) );
  ANDN U8550 ( .B(y[1767]), .A(x[1767]), .Z(n9406) );
  ANDN U8551 ( .B(n5584), .A(n9406), .Z(n13498) );
  NAND U8552 ( .A(n5585), .B(n13498), .Z(n5586) );
  NANDN U8553 ( .A(n13501), .B(n5586), .Z(n5588) );
  NANDN U8554 ( .A(x[1768]), .B(y[1768]), .Z(n5587) );
  ANDN U8555 ( .B(y[1769]), .A(x[1769]), .Z(n9412) );
  ANDN U8556 ( .B(n5587), .A(n9412), .Z(n13502) );
  NAND U8557 ( .A(n5588), .B(n13502), .Z(n5589) );
  NANDN U8558 ( .A(n13505), .B(n5589), .Z(n5590) );
  AND U8559 ( .A(n13506), .B(n5590), .Z(n5591) );
  OR U8560 ( .A(n13508), .B(n5591), .Z(n5593) );
  NANDN U8561 ( .A(x[1772]), .B(y[1772]), .Z(n5592) );
  ANDN U8562 ( .B(y[1773]), .A(x[1773]), .Z(n9428) );
  ANDN U8563 ( .B(n5592), .A(n9428), .Z(n13510) );
  NAND U8564 ( .A(n5593), .B(n13510), .Z(n5594) );
  NANDN U8565 ( .A(y[1774]), .B(x[1774]), .Z(n9431) );
  NAND U8566 ( .A(n5594), .B(n9431), .Z(n5595) );
  NANDN U8567 ( .A(y[1773]), .B(x[1773]), .Z(n13513) );
  NANDN U8568 ( .A(n5595), .B(n13513), .Z(n5597) );
  ANDN U8569 ( .B(y[1775]), .A(x[1775]), .Z(n9433) );
  NANDN U8570 ( .A(x[1774]), .B(y[1774]), .Z(n5596) );
  NANDN U8571 ( .A(n9433), .B(n5596), .Z(n9424) );
  ANDN U8572 ( .B(n5597), .A(n9424), .Z(n5600) );
  ANDN U8573 ( .B(x[1775]), .A(y[1775]), .Z(n9432) );
  NANDN U8574 ( .A(y[1776]), .B(x[1776]), .Z(n5598) );
  NANDN U8575 ( .A(n9432), .B(n5598), .Z(n5599) );
  OR U8576 ( .A(n5600), .B(n5599), .Z(n5601) );
  ANDN U8577 ( .B(y[1777]), .A(x[1777]), .Z(n9429) );
  NANDN U8578 ( .A(x[1776]), .B(y[1776]), .Z(n9430) );
  NANDN U8579 ( .A(n9429), .B(n9430), .Z(n9425) );
  ANDN U8580 ( .B(n5601), .A(n9425), .Z(n5604) );
  NANDN U8581 ( .A(y[1778]), .B(x[1778]), .Z(n5603) );
  NANDN U8582 ( .A(y[1777]), .B(x[1777]), .Z(n5602) );
  AND U8583 ( .A(n5603), .B(n5602), .Z(n9439) );
  NANDN U8584 ( .A(n5604), .B(n9439), .Z(n5605) );
  AND U8585 ( .A(n13518), .B(n5605), .Z(n5606) );
  OR U8586 ( .A(n13521), .B(n5606), .Z(n5608) );
  NANDN U8587 ( .A(x[1780]), .B(y[1780]), .Z(n13522) );
  ANDN U8588 ( .B(y[1781]), .A(x[1781]), .Z(n6171) );
  ANDN U8589 ( .B(n13522), .A(n6171), .Z(n5607) );
  NAND U8590 ( .A(n5608), .B(n5607), .Z(n5609) );
  NANDN U8591 ( .A(n5610), .B(n5609), .Z(n5611) );
  NANDN U8592 ( .A(n5612), .B(n5611), .Z(n5614) );
  NANDN U8593 ( .A(y[1783]), .B(x[1783]), .Z(n9447) );
  IV U8594 ( .A(x[1784]), .Z(n9451) );
  OR U8595 ( .A(y[1784]), .B(n9451), .Z(n5613) );
  NAND U8596 ( .A(n9447), .B(n5613), .Z(n13533) );
  ANDN U8597 ( .B(n5614), .A(n13533), .Z(n5615) );
  OR U8598 ( .A(n13535), .B(n5615), .Z(n5616) );
  NANDN U8599 ( .A(n13537), .B(n5616), .Z(n5617) );
  NANDN U8600 ( .A(n13539), .B(n5617), .Z(n5618) );
  NAND U8601 ( .A(n5619), .B(n5618), .Z(n5620) );
  NANDN U8602 ( .A(n13543), .B(n5620), .Z(n5621) );
  IV U8603 ( .A(x[1789]), .Z(n9465) );
  OR U8604 ( .A(n5621), .B(n9465), .Z(n5624) );
  XNOR U8605 ( .A(n5621), .B(x[1789]), .Z(n5622) );
  NANDN U8606 ( .A(y[1789]), .B(n5622), .Z(n5623) );
  AND U8607 ( .A(n5624), .B(n5623), .Z(n5625) );
  OR U8608 ( .A(n5625), .B(y[1790]), .Z(n5628) );
  XOR U8609 ( .A(y[1790]), .B(n5625), .Z(n5626) );
  NAND U8610 ( .A(n5626), .B(x[1790]), .Z(n5627) );
  NAND U8611 ( .A(n5628), .B(n5627), .Z(n5629) );
  AND U8612 ( .A(n6165), .B(n5629), .Z(n5631) );
  XOR U8613 ( .A(x[1792]), .B(y[1792]), .Z(n6166) );
  NANDN U8614 ( .A(y[1791]), .B(x[1791]), .Z(n5630) );
  NANDN U8615 ( .A(n6166), .B(n5630), .Z(n9470) );
  OR U8616 ( .A(n5631), .B(n9470), .Z(n5632) );
  NANDN U8617 ( .A(n6168), .B(n5632), .Z(n5635) );
  NANDN U8618 ( .A(y[1793]), .B(x[1793]), .Z(n5634) );
  NANDN U8619 ( .A(y[1794]), .B(x[1794]), .Z(n5633) );
  AND U8620 ( .A(n5634), .B(n5633), .Z(n13553) );
  NAND U8621 ( .A(n5635), .B(n13553), .Z(n5636) );
  NANDN U8622 ( .A(n13555), .B(n5636), .Z(n5637) );
  AND U8623 ( .A(n9475), .B(n5637), .Z(n5643) );
  NANDN U8624 ( .A(x[1798]), .B(y[1798]), .Z(n5642) );
  NANDN U8625 ( .A(x[1796]), .B(y[1796]), .Z(n5638) );
  ANDN U8626 ( .B(y[1797]), .A(x[1797]), .Z(n13561) );
  ANDN U8627 ( .B(n5638), .A(n13561), .Z(n5640) );
  NANDN U8628 ( .A(n5640), .B(n5639), .Z(n5641) );
  NAND U8629 ( .A(n5642), .B(n5641), .Z(n9478) );
  OR U8630 ( .A(n5643), .B(n9478), .Z(n5644) );
  AND U8631 ( .A(n9479), .B(n5644), .Z(n5645) );
  NANDN U8632 ( .A(x[1799]), .B(y[1799]), .Z(n13562) );
  NANDN U8633 ( .A(n5645), .B(n13562), .Z(n5646) );
  NANDN U8634 ( .A(y[1800]), .B(x[1800]), .Z(n9991) );
  NAND U8635 ( .A(n5646), .B(n9991), .Z(n5647) );
  NANDN U8636 ( .A(x[1801]), .B(y[1801]), .Z(n9487) );
  ANDN U8637 ( .B(y[1800]), .A(x[1800]), .Z(n9483) );
  ANDN U8638 ( .B(n9487), .A(n9483), .Z(n13563) );
  NAND U8639 ( .A(n5647), .B(n13563), .Z(n5648) );
  NAND U8640 ( .A(n5649), .B(n5648), .Z(n5650) );
  NANDN U8641 ( .A(x[1802]), .B(y[1802]), .Z(n13565) );
  NAND U8642 ( .A(n5650), .B(n13565), .Z(n5651) );
  NANDN U8643 ( .A(x[1803]), .B(y[1803]), .Z(n13567) );
  NANDN U8644 ( .A(n5651), .B(n13567), .Z(n5652) );
  AND U8645 ( .A(n5653), .B(n5652), .Z(n5654) );
  OR U8646 ( .A(n13569), .B(n5654), .Z(n5655) );
  NANDN U8647 ( .A(n13570), .B(n5655), .Z(n5656) );
  NANDN U8648 ( .A(n13571), .B(n5656), .Z(n5657) );
  NANDN U8649 ( .A(n13572), .B(n5657), .Z(n5658) );
  AND U8650 ( .A(n13574), .B(n5658), .Z(n5659) );
  NANDN U8651 ( .A(x[1809]), .B(y[1809]), .Z(n6159) );
  NAND U8652 ( .A(n5659), .B(n6159), .Z(n5660) );
  NAND U8653 ( .A(n5661), .B(n5660), .Z(n5662) );
  NANDN U8654 ( .A(x[1810]), .B(y[1810]), .Z(n6158) );
  NAND U8655 ( .A(n5662), .B(n6158), .Z(n5663) );
  NANDN U8656 ( .A(x[1811]), .B(y[1811]), .Z(n13582) );
  NANDN U8657 ( .A(n5663), .B(n13582), .Z(n5664) );
  NANDN U8658 ( .A(n13584), .B(n5664), .Z(n5665) );
  NANDN U8659 ( .A(n13587), .B(n5665), .Z(n5666) );
  NANDN U8660 ( .A(n13589), .B(n5666), .Z(n5668) );
  NANDN U8661 ( .A(x[1814]), .B(y[1814]), .Z(n5667) );
  ANDN U8662 ( .B(y[1815]), .A(x[1815]), .Z(n9526) );
  ANDN U8663 ( .B(n5667), .A(n9526), .Z(n13590) );
  NAND U8664 ( .A(n5668), .B(n13590), .Z(n5669) );
  AND U8665 ( .A(n13592), .B(n5669), .Z(n5670) );
  NANDN U8666 ( .A(x[1816]), .B(y[1816]), .Z(n13594) );
  NANDN U8667 ( .A(n5670), .B(n13594), .Z(n5673) );
  NANDN U8668 ( .A(y[1816]), .B(x[1816]), .Z(n5672) );
  NANDN U8669 ( .A(y[1817]), .B(x[1817]), .Z(n5671) );
  AND U8670 ( .A(n5672), .B(n5671), .Z(n13597) );
  NAND U8671 ( .A(n5673), .B(n13597), .Z(n5674) );
  NANDN U8672 ( .A(x[1817]), .B(y[1817]), .Z(n9531) );
  NAND U8673 ( .A(n5674), .B(n9531), .Z(n5675) );
  NANDN U8674 ( .A(y[1818]), .B(x[1818]), .Z(n13601) );
  NAND U8675 ( .A(n5675), .B(n13601), .Z(n5676) );
  ANDN U8676 ( .B(y[1818]), .A(x[1818]), .Z(n9530) );
  ANDN U8677 ( .B(n5676), .A(n9530), .Z(n5677) );
  NANDN U8678 ( .A(x[1819]), .B(y[1819]), .Z(n13602) );
  NAND U8679 ( .A(n5677), .B(n13602), .Z(n5678) );
  NANDN U8680 ( .A(n13605), .B(n5678), .Z(n5679) );
  NANDN U8681 ( .A(n13607), .B(n5679), .Z(n5680) );
  NANDN U8682 ( .A(n13609), .B(n5680), .Z(n5681) );
  AND U8683 ( .A(n13610), .B(n5681), .Z(n5682) );
  NANDN U8684 ( .A(x[1823]), .B(y[1823]), .Z(n9552) );
  NAND U8685 ( .A(n5682), .B(n9552), .Z(n5683) );
  NAND U8686 ( .A(n5684), .B(n5683), .Z(n5685) );
  ANDN U8687 ( .B(y[1825]), .A(x[1825]), .Z(n9559) );
  ANDN U8688 ( .B(y[1824]), .A(x[1824]), .Z(n9554) );
  NOR U8689 ( .A(n9559), .B(n9554), .Z(n13618) );
  NAND U8690 ( .A(n5685), .B(n13618), .Z(n5686) );
  AND U8691 ( .A(n13622), .B(n5686), .Z(n5689) );
  NANDN U8692 ( .A(x[1826]), .B(y[1826]), .Z(n5688) );
  ANDN U8693 ( .B(n5688), .A(n5687), .Z(n13624) );
  NANDN U8694 ( .A(n5689), .B(n13624), .Z(n5690) );
  NANDN U8695 ( .A(n9561), .B(n5690), .Z(n5691) );
  NANDN U8696 ( .A(n13629), .B(n5691), .Z(n5692) );
  NAND U8697 ( .A(n5693), .B(n5692), .Z(n5694) );
  NANDN U8698 ( .A(x[1830]), .B(y[1830]), .Z(n13633) );
  NAND U8699 ( .A(n5694), .B(n13633), .Z(n5695) );
  NAND U8700 ( .A(n5696), .B(n5695), .Z(n5697) );
  NANDN U8701 ( .A(x[1831]), .B(y[1831]), .Z(n9569) );
  AND U8702 ( .A(n5697), .B(n9569), .Z(n5698) );
  NANDN U8703 ( .A(y[1832]), .B(x[1832]), .Z(n13638) );
  NANDN U8704 ( .A(n5698), .B(n13638), .Z(n5699) );
  AND U8705 ( .A(n5700), .B(n5699), .Z(n5701) );
  ANDN U8706 ( .B(x[1834]), .A(y[1834]), .Z(n9577) );
  ANDN U8707 ( .B(x[1833]), .A(y[1833]), .Z(n9573) );
  NOR U8708 ( .A(n9577), .B(n9573), .Z(n13642) );
  NANDN U8709 ( .A(n5701), .B(n13642), .Z(n5702) );
  NANDN U8710 ( .A(n13644), .B(n5702), .Z(n5704) );
  NANDN U8711 ( .A(y[1835]), .B(x[1835]), .Z(n5703) );
  ANDN U8712 ( .B(x[1836]), .A(y[1836]), .Z(n9583) );
  ANDN U8713 ( .B(n5703), .A(n9583), .Z(n13646) );
  NAND U8714 ( .A(n5704), .B(n13646), .Z(n5705) );
  NANDN U8715 ( .A(n13649), .B(n5705), .Z(n5707) );
  NANDN U8716 ( .A(y[1837]), .B(x[1837]), .Z(n5706) );
  ANDN U8717 ( .B(x[1838]), .A(y[1838]), .Z(n9589) );
  ANDN U8718 ( .B(n5706), .A(n9589), .Z(n13650) );
  NAND U8719 ( .A(n5707), .B(n13650), .Z(n5708) );
  NANDN U8720 ( .A(n13653), .B(n5708), .Z(n5709) );
  NANDN U8721 ( .A(y[1839]), .B(x[1839]), .Z(n13656) );
  NAND U8722 ( .A(n5709), .B(n13656), .Z(n5710) );
  NANDN U8723 ( .A(x[1840]), .B(y[1840]), .Z(n9989) );
  NAND U8724 ( .A(n5710), .B(n9989), .Z(n5711) );
  ANDN U8725 ( .B(x[1840]), .A(y[1840]), .Z(n13654) );
  ANDN U8726 ( .B(x[1841]), .A(y[1841]), .Z(n13663) );
  NOR U8727 ( .A(n13654), .B(n13663), .Z(n9595) );
  NAND U8728 ( .A(n5711), .B(n9595), .Z(n5712) );
  AND U8729 ( .A(n9988), .B(n5712), .Z(n5713) );
  NANDN U8730 ( .A(y[1842]), .B(x[1842]), .Z(n13661) );
  NANDN U8731 ( .A(n5713), .B(n13661), .Z(n5714) );
  AND U8732 ( .A(n13664), .B(n5714), .Z(n5715) );
  ANDN U8733 ( .B(x[1844]), .A(y[1844]), .Z(n9606) );
  NOR U8734 ( .A(n5715), .B(n9606), .Z(n5716) );
  NANDN U8735 ( .A(y[1843]), .B(x[1843]), .Z(n13667) );
  NAND U8736 ( .A(n5716), .B(n13667), .Z(n5717) );
  NANDN U8737 ( .A(x[1844]), .B(y[1844]), .Z(n13668) );
  NAND U8738 ( .A(n5717), .B(n13668), .Z(n5718) );
  NANDN U8739 ( .A(n9605), .B(n5718), .Z(n5719) );
  NANDN U8740 ( .A(n9609), .B(n5719), .Z(n5720) );
  AND U8741 ( .A(n9610), .B(n5720), .Z(n5721) );
  NANDN U8742 ( .A(x[1847]), .B(y[1847]), .Z(n13678) );
  NANDN U8743 ( .A(n5721), .B(n13678), .Z(n5722) );
  NANDN U8744 ( .A(y[1848]), .B(x[1848]), .Z(n13682) );
  NAND U8745 ( .A(n5722), .B(n13682), .Z(n5723) );
  ANDN U8746 ( .B(y[1848]), .A(x[1848]), .Z(n9612) );
  ANDN U8747 ( .B(y[1849]), .A(x[1849]), .Z(n9620) );
  NOR U8748 ( .A(n9612), .B(n9620), .Z(n13684) );
  NAND U8749 ( .A(n5723), .B(n13684), .Z(n5724) );
  NANDN U8750 ( .A(n13687), .B(n5724), .Z(n5725) );
  AND U8751 ( .A(n13689), .B(n5725), .Z(n5726) );
  NANDN U8752 ( .A(x[1851]), .B(y[1851]), .Z(n9626) );
  NAND U8753 ( .A(n5726), .B(n9626), .Z(n5727) );
  AND U8754 ( .A(n13693), .B(n5727), .Z(n5728) );
  ANDN U8755 ( .B(y[1853]), .A(x[1853]), .Z(n9633) );
  ANDN U8756 ( .B(y[1852]), .A(x[1852]), .Z(n9628) );
  NOR U8757 ( .A(n9633), .B(n9628), .Z(n13694) );
  NANDN U8758 ( .A(n5728), .B(n13694), .Z(n5729) );
  NANDN U8759 ( .A(n13697), .B(n5729), .Z(n5731) );
  NANDN U8760 ( .A(x[1854]), .B(y[1854]), .Z(n5730) );
  ANDN U8761 ( .B(y[1855]), .A(x[1855]), .Z(n9639) );
  ANDN U8762 ( .B(n5730), .A(n9639), .Z(n13699) );
  NAND U8763 ( .A(n5731), .B(n13699), .Z(n5734) );
  NANDN U8764 ( .A(y[1855]), .B(x[1855]), .Z(n5733) );
  NANDN U8765 ( .A(y[1856]), .B(x[1856]), .Z(n5732) );
  AND U8766 ( .A(n5733), .B(n5732), .Z(n13700) );
  NAND U8767 ( .A(n5734), .B(n13700), .Z(n5735) );
  NANDN U8768 ( .A(n13703), .B(n5735), .Z(n5736) );
  NANDN U8769 ( .A(y[1858]), .B(x[1858]), .Z(n6145) );
  NAND U8770 ( .A(n5736), .B(n6145), .Z(n5737) );
  NANDN U8771 ( .A(y[1857]), .B(x[1857]), .Z(n13704) );
  NANDN U8772 ( .A(n5737), .B(n13704), .Z(n5738) );
  NANDN U8773 ( .A(n13707), .B(n5738), .Z(n5739) );
  IV U8774 ( .A(x[1859]), .Z(n6143) );
  OR U8775 ( .A(n5739), .B(n6143), .Z(n5742) );
  XNOR U8776 ( .A(n5739), .B(x[1859]), .Z(n5740) );
  NANDN U8777 ( .A(y[1859]), .B(n5740), .Z(n5741) );
  NAND U8778 ( .A(n5742), .B(n5741), .Z(n5743) );
  NANDN U8779 ( .A(y[1860]), .B(x[1860]), .Z(n13712) );
  NANDN U8780 ( .A(n5743), .B(n13712), .Z(n5745) );
  NANDN U8781 ( .A(x[1861]), .B(y[1861]), .Z(n13714) );
  NANDN U8782 ( .A(x[1860]), .B(y[1860]), .Z(n6141) );
  AND U8783 ( .A(n13714), .B(n6141), .Z(n5744) );
  NAND U8784 ( .A(n5745), .B(n5744), .Z(n5748) );
  NANDN U8785 ( .A(y[1861]), .B(x[1861]), .Z(n5747) );
  NANDN U8786 ( .A(y[1862]), .B(x[1862]), .Z(n5746) );
  AND U8787 ( .A(n5747), .B(n5746), .Z(n13716) );
  NAND U8788 ( .A(n5748), .B(n13716), .Z(n5751) );
  NANDN U8789 ( .A(x[1863]), .B(y[1863]), .Z(n5750) );
  NANDN U8790 ( .A(x[1862]), .B(y[1862]), .Z(n5749) );
  NAND U8791 ( .A(n5750), .B(n5749), .Z(n13719) );
  ANDN U8792 ( .B(n5751), .A(n13719), .Z(n5754) );
  NANDN U8793 ( .A(y[1863]), .B(x[1863]), .Z(n5753) );
  NANDN U8794 ( .A(y[1864]), .B(x[1864]), .Z(n5752) );
  AND U8795 ( .A(n5753), .B(n5752), .Z(n13720) );
  NANDN U8796 ( .A(n5754), .B(n13720), .Z(n5755) );
  NANDN U8797 ( .A(n13722), .B(n5755), .Z(n5758) );
  NANDN U8798 ( .A(y[1865]), .B(x[1865]), .Z(n5757) );
  NANDN U8799 ( .A(y[1866]), .B(x[1866]), .Z(n5756) );
  AND U8800 ( .A(n5757), .B(n5756), .Z(n13724) );
  NAND U8801 ( .A(n5758), .B(n13724), .Z(n5761) );
  NANDN U8802 ( .A(x[1867]), .B(y[1867]), .Z(n5760) );
  NANDN U8803 ( .A(x[1866]), .B(y[1866]), .Z(n5759) );
  NAND U8804 ( .A(n5760), .B(n5759), .Z(n13727) );
  ANDN U8805 ( .B(n5761), .A(n13727), .Z(n5762) );
  ANDN U8806 ( .B(n13730), .A(n5762), .Z(n5763) );
  OR U8807 ( .A(n5763), .B(y[1868]), .Z(n5766) );
  IV U8808 ( .A(x[1868]), .Z(n9656) );
  XOR U8809 ( .A(y[1868]), .B(n5763), .Z(n5764) );
  NANDN U8810 ( .A(n9656), .B(n5764), .Z(n5765) );
  NAND U8811 ( .A(n5766), .B(n5765), .Z(n5767) );
  AND U8812 ( .A(n9985), .B(n5767), .Z(n5770) );
  NANDN U8813 ( .A(y[1870]), .B(x[1870]), .Z(n5768) );
  NAND U8814 ( .A(n5769), .B(n5768), .Z(n9664) );
  NANDN U8815 ( .A(y[1869]), .B(x[1869]), .Z(n9659) );
  NANDN U8816 ( .A(n9664), .B(n9659), .Z(n13735) );
  OR U8817 ( .A(n5770), .B(n13735), .Z(n5771) );
  NANDN U8818 ( .A(n13737), .B(n5771), .Z(n5772) );
  NANDN U8819 ( .A(n13739), .B(n5772), .Z(n5775) );
  NANDN U8820 ( .A(x[1873]), .B(y[1873]), .Z(n5774) );
  NANDN U8821 ( .A(x[1874]), .B(y[1874]), .Z(n5773) );
  NAND U8822 ( .A(n5774), .B(n5773), .Z(n13741) );
  ANDN U8823 ( .B(n5775), .A(n13741), .Z(n5776) );
  NANDN U8824 ( .A(y[1874]), .B(x[1874]), .Z(n13742) );
  NANDN U8825 ( .A(n5776), .B(n13742), .Z(n5777) );
  AND U8826 ( .A(n13745), .B(n5777), .Z(n5778) );
  OR U8827 ( .A(n13747), .B(n5778), .Z(n5779) );
  NANDN U8828 ( .A(n13749), .B(n5779), .Z(n5781) );
  ANDN U8829 ( .B(x[1878]), .A(y[1878]), .Z(n9683) );
  NANDN U8830 ( .A(y[1877]), .B(x[1877]), .Z(n5780) );
  NANDN U8831 ( .A(n9683), .B(n5780), .Z(n13751) );
  ANDN U8832 ( .B(n5781), .A(n13751), .Z(n5782) );
  OR U8833 ( .A(n5783), .B(n5782), .Z(n5784) );
  NANDN U8834 ( .A(n9680), .B(n5784), .Z(n5785) );
  NANDN U8835 ( .A(x[1880]), .B(y[1880]), .Z(n6134) );
  NAND U8836 ( .A(n5785), .B(n6134), .Z(n5786) );
  NANDN U8837 ( .A(x[1881]), .B(y[1881]), .Z(n13761) );
  NANDN U8838 ( .A(n5786), .B(n13761), .Z(n5787) );
  ANDN U8839 ( .B(x[1882]), .A(y[1882]), .Z(n13763) );
  NANDN U8840 ( .A(y[1881]), .B(x[1881]), .Z(n9984) );
  NANDN U8841 ( .A(n13763), .B(n9984), .Z(n9688) );
  ANDN U8842 ( .B(n5787), .A(n9688), .Z(n5790) );
  NANDN U8843 ( .A(x[1882]), .B(y[1882]), .Z(n5789) );
  NANDN U8844 ( .A(x[1883]), .B(y[1883]), .Z(n5788) );
  AND U8845 ( .A(n5789), .B(n5788), .Z(n13765) );
  NANDN U8846 ( .A(n5790), .B(n13765), .Z(n5793) );
  NANDN U8847 ( .A(y[1884]), .B(x[1884]), .Z(n5792) );
  NANDN U8848 ( .A(y[1883]), .B(x[1883]), .Z(n5791) );
  NAND U8849 ( .A(n5792), .B(n5791), .Z(n13767) );
  ANDN U8850 ( .B(n5793), .A(n13767), .Z(n5796) );
  NANDN U8851 ( .A(x[1885]), .B(y[1885]), .Z(n5795) );
  NANDN U8852 ( .A(x[1884]), .B(y[1884]), .Z(n5794) );
  AND U8853 ( .A(n5795), .B(n5794), .Z(n13769) );
  NANDN U8854 ( .A(n5796), .B(n13769), .Z(n5797) );
  ANDN U8855 ( .B(x[1886]), .A(y[1886]), .Z(n9695) );
  ANDN U8856 ( .B(n5797), .A(n9695), .Z(n5798) );
  NANDN U8857 ( .A(y[1885]), .B(x[1885]), .Z(n13770) );
  NAND U8858 ( .A(n5798), .B(n13770), .Z(n5801) );
  NANDN U8859 ( .A(x[1886]), .B(y[1886]), .Z(n5800) );
  NANDN U8860 ( .A(x[1888]), .B(y[1888]), .Z(n5803) );
  NANDN U8861 ( .A(x[1887]), .B(y[1887]), .Z(n5799) );
  NAND U8862 ( .A(n5803), .B(n5799), .Z(n9696) );
  ANDN U8863 ( .B(n5800), .A(n9696), .Z(n13772) );
  NAND U8864 ( .A(n5801), .B(n13772), .Z(n5802) );
  NANDN U8865 ( .A(y[1888]), .B(x[1888]), .Z(n9698) );
  NAND U8866 ( .A(n5802), .B(n9698), .Z(n5805) );
  NANDN U8867 ( .A(y[1887]), .B(x[1887]), .Z(n9694) );
  NANDN U8868 ( .A(n9694), .B(n5803), .Z(n5804) );
  NANDN U8869 ( .A(n5805), .B(n5804), .Z(n5806) );
  NANDN U8870 ( .A(x[1889]), .B(y[1889]), .Z(n13776) );
  NAND U8871 ( .A(n5806), .B(n13776), .Z(n5807) );
  AND U8872 ( .A(n5808), .B(n5807), .Z(n5809) );
  OR U8873 ( .A(n13781), .B(n5809), .Z(n5810) );
  NANDN U8874 ( .A(n13782), .B(n5810), .Z(n5811) );
  NANDN U8875 ( .A(x[1893]), .B(y[1893]), .Z(n6129) );
  NAND U8876 ( .A(n5811), .B(n6129), .Z(n5812) );
  NANDN U8877 ( .A(x[1892]), .B(y[1892]), .Z(n13784) );
  NANDN U8878 ( .A(n5812), .B(n13784), .Z(n5813) );
  NANDN U8879 ( .A(n13786), .B(n5813), .Z(n5816) );
  NANDN U8880 ( .A(x[1895]), .B(y[1895]), .Z(n5815) );
  NANDN U8881 ( .A(x[1894]), .B(y[1894]), .Z(n5814) );
  AND U8882 ( .A(n5815), .B(n5814), .Z(n6130) );
  NAND U8883 ( .A(n5816), .B(n6130), .Z(n5819) );
  NANDN U8884 ( .A(y[1896]), .B(x[1896]), .Z(n5818) );
  NANDN U8885 ( .A(y[1895]), .B(x[1895]), .Z(n5817) );
  NAND U8886 ( .A(n5818), .B(n5817), .Z(n13791) );
  ANDN U8887 ( .B(n5819), .A(n13791), .Z(n5822) );
  NANDN U8888 ( .A(x[1896]), .B(y[1896]), .Z(n5821) );
  NANDN U8889 ( .A(x[1897]), .B(y[1897]), .Z(n5820) );
  AND U8890 ( .A(n5821), .B(n5820), .Z(n13793) );
  NANDN U8891 ( .A(n5822), .B(n13793), .Z(n5823) );
  NANDN U8892 ( .A(n13795), .B(n5823), .Z(n5826) );
  NANDN U8893 ( .A(x[1899]), .B(y[1899]), .Z(n5825) );
  NANDN U8894 ( .A(x[1898]), .B(y[1898]), .Z(n5824) );
  AND U8895 ( .A(n5825), .B(n5824), .Z(n13797) );
  NAND U8896 ( .A(n5826), .B(n13797), .Z(n5827) );
  NAND U8897 ( .A(n5828), .B(n5827), .Z(n5829) );
  NANDN U8898 ( .A(x[1901]), .B(y[1901]), .Z(n6125) );
  NAND U8899 ( .A(n5829), .B(n6125), .Z(n5830) );
  NANDN U8900 ( .A(x[1900]), .B(y[1900]), .Z(n13800) );
  NANDN U8901 ( .A(n5830), .B(n13800), .Z(n5831) );
  AND U8902 ( .A(n6123), .B(n5831), .Z(n5832) );
  NANDN U8903 ( .A(n6127), .B(n5832), .Z(n5833) );
  AND U8904 ( .A(n6120), .B(n5833), .Z(n5834) );
  NANDN U8905 ( .A(x[1902]), .B(y[1902]), .Z(n6124) );
  NAND U8906 ( .A(n5834), .B(n6124), .Z(n5835) );
  NAND U8907 ( .A(n5836), .B(n5835), .Z(n5837) );
  NANDN U8908 ( .A(n6121), .B(n5837), .Z(n5840) );
  NANDN U8909 ( .A(y[1906]), .B(x[1906]), .Z(n5839) );
  NANDN U8910 ( .A(y[1905]), .B(x[1905]), .Z(n5838) );
  NAND U8911 ( .A(n5839), .B(n5838), .Z(n6119) );
  ANDN U8912 ( .B(n5840), .A(n6119), .Z(n5843) );
  NANDN U8913 ( .A(x[1906]), .B(y[1906]), .Z(n5842) );
  NANDN U8914 ( .A(x[1907]), .B(y[1907]), .Z(n5841) );
  AND U8915 ( .A(n5842), .B(n5841), .Z(n13810) );
  NANDN U8916 ( .A(n5843), .B(n13810), .Z(n5846) );
  NANDN U8917 ( .A(y[1908]), .B(x[1908]), .Z(n5845) );
  NANDN U8918 ( .A(y[1907]), .B(x[1907]), .Z(n5844) );
  NAND U8919 ( .A(n5845), .B(n5844), .Z(n13811) );
  ANDN U8920 ( .B(n5846), .A(n13811), .Z(n5849) );
  NANDN U8921 ( .A(x[1908]), .B(y[1908]), .Z(n5848) );
  NANDN U8922 ( .A(x[1909]), .B(y[1909]), .Z(n5847) );
  AND U8923 ( .A(n5848), .B(n5847), .Z(n13812) );
  NANDN U8924 ( .A(n5849), .B(n13812), .Z(n5852) );
  NANDN U8925 ( .A(y[1910]), .B(x[1910]), .Z(n5851) );
  NANDN U8926 ( .A(y[1909]), .B(x[1909]), .Z(n5850) );
  NAND U8927 ( .A(n5851), .B(n5850), .Z(n13813) );
  ANDN U8928 ( .B(n5852), .A(n13813), .Z(n5855) );
  NANDN U8929 ( .A(x[1910]), .B(y[1910]), .Z(n5854) );
  NANDN U8930 ( .A(x[1911]), .B(y[1911]), .Z(n5853) );
  AND U8931 ( .A(n5854), .B(n5853), .Z(n13814) );
  NANDN U8932 ( .A(n5855), .B(n13814), .Z(n5856) );
  NANDN U8933 ( .A(n13815), .B(n5856), .Z(n5857) );
  AND U8934 ( .A(n13816), .B(n5857), .Z(n5858) );
  OR U8935 ( .A(n5859), .B(n5858), .Z(n5860) );
  NANDN U8936 ( .A(n13818), .B(n5860), .Z(n5861) );
  ANDN U8937 ( .B(x[1916]), .A(y[1916]), .Z(n9739) );
  ANDN U8938 ( .B(x[1915]), .A(y[1915]), .Z(n9736) );
  NOR U8939 ( .A(n9739), .B(n9736), .Z(n13820) );
  NAND U8940 ( .A(n5861), .B(n13820), .Z(n5863) );
  IV U8941 ( .A(y[1917]), .Z(n6115) );
  IV U8942 ( .A(x[1917]), .Z(n6114) );
  NANDN U8943 ( .A(n6115), .B(n6114), .Z(n5862) );
  NANDN U8944 ( .A(x[1916]), .B(y[1916]), .Z(n9737) );
  NAND U8945 ( .A(n5862), .B(n9737), .Z(n13821) );
  ANDN U8946 ( .B(n5863), .A(n13821), .Z(n5865) );
  NANDN U8947 ( .A(y[1917]), .B(x[1917]), .Z(n5864) );
  ANDN U8948 ( .B(x[1918]), .A(y[1918]), .Z(n9747) );
  ANDN U8949 ( .B(n5864), .A(n9747), .Z(n13822) );
  NANDN U8950 ( .A(n5865), .B(n13822), .Z(n5866) );
  AND U8951 ( .A(n9982), .B(n5866), .Z(n5867) );
  OR U8952 ( .A(n13823), .B(n5867), .Z(n5871) );
  ANDN U8953 ( .B(y[1920]), .A(x[1920]), .Z(n13825) );
  NANDN U8954 ( .A(x[1919]), .B(y[1919]), .Z(n9981) );
  NANDN U8955 ( .A(n9981), .B(n5868), .Z(n5869) );
  NANDN U8956 ( .A(n13825), .B(n5869), .Z(n9749) );
  ANDN U8957 ( .B(y[1921]), .A(x[1921]), .Z(n9751) );
  NOR U8958 ( .A(n9749), .B(n9751), .Z(n5870) );
  NAND U8959 ( .A(n5871), .B(n5870), .Z(n5872) );
  NAND U8960 ( .A(n6112), .B(n5872), .Z(n5874) );
  NANDN U8961 ( .A(y[1922]), .B(n5874), .Z(n5873) );
  AND U8962 ( .A(n9755), .B(n5873), .Z(n5877) );
  XNOR U8963 ( .A(n5874), .B(y[1922]), .Z(n5875) );
  NAND U8964 ( .A(n5875), .B(x[1922]), .Z(n5876) );
  NAND U8965 ( .A(n5877), .B(n5876), .Z(n5880) );
  NANDN U8966 ( .A(x[1923]), .B(y[1923]), .Z(n5879) );
  NANDN U8967 ( .A(x[1924]), .B(y[1924]), .Z(n5878) );
  AND U8968 ( .A(n5879), .B(n5878), .Z(n13832) );
  NAND U8969 ( .A(n5880), .B(n13832), .Z(n5881) );
  NANDN U8970 ( .A(n13835), .B(n5881), .Z(n5882) );
  NANDN U8971 ( .A(x[1925]), .B(y[1925]), .Z(n13837) );
  NAND U8972 ( .A(n5882), .B(n13837), .Z(n5883) );
  NANDN U8973 ( .A(y[1926]), .B(x[1926]), .Z(n13838) );
  NAND U8974 ( .A(n5883), .B(n13838), .Z(n5886) );
  NANDN U8975 ( .A(x[1926]), .B(y[1926]), .Z(n5885) );
  NANDN U8976 ( .A(x[1927]), .B(y[1927]), .Z(n5884) );
  AND U8977 ( .A(n5885), .B(n5884), .Z(n13840) );
  NAND U8978 ( .A(n5886), .B(n13840), .Z(n5887) );
  AND U8979 ( .A(n13842), .B(n5887), .Z(n5888) );
  NANDN U8980 ( .A(n9764), .B(n5888), .Z(n5889) );
  NANDN U8981 ( .A(n5890), .B(n5889), .Z(n5891) );
  AND U8982 ( .A(n5892), .B(n5891), .Z(n5893) );
  NANDN U8983 ( .A(x[1931]), .B(y[1931]), .Z(n9770) );
  NANDN U8984 ( .A(x[1930]), .B(y[1930]), .Z(n9767) );
  NAND U8985 ( .A(n9770), .B(n9767), .Z(n13852) );
  OR U8986 ( .A(n5893), .B(n13852), .Z(n5896) );
  NANDN U8987 ( .A(y[1932]), .B(x[1932]), .Z(n5895) );
  NANDN U8988 ( .A(y[1931]), .B(x[1931]), .Z(n5894) );
  NAND U8989 ( .A(n5895), .B(n5894), .Z(n13855) );
  ANDN U8990 ( .B(n5896), .A(n13855), .Z(n5899) );
  NANDN U8991 ( .A(x[1932]), .B(y[1932]), .Z(n5898) );
  NANDN U8992 ( .A(x[1933]), .B(y[1933]), .Z(n5897) );
  AND U8993 ( .A(n5898), .B(n5897), .Z(n13857) );
  NANDN U8994 ( .A(n5899), .B(n13857), .Z(n5902) );
  NANDN U8995 ( .A(y[1934]), .B(x[1934]), .Z(n5901) );
  NANDN U8996 ( .A(y[1933]), .B(x[1933]), .Z(n5900) );
  NAND U8997 ( .A(n5901), .B(n5900), .Z(n13859) );
  ANDN U8998 ( .B(n5902), .A(n13859), .Z(n5905) );
  NANDN U8999 ( .A(x[1934]), .B(y[1934]), .Z(n5904) );
  NANDN U9000 ( .A(x[1935]), .B(y[1935]), .Z(n5903) );
  AND U9001 ( .A(n5904), .B(n5903), .Z(n13861) );
  NANDN U9002 ( .A(n5905), .B(n13861), .Z(n5908) );
  NANDN U9003 ( .A(y[1936]), .B(x[1936]), .Z(n5907) );
  NANDN U9004 ( .A(y[1935]), .B(x[1935]), .Z(n5906) );
  NAND U9005 ( .A(n5907), .B(n5906), .Z(n13863) );
  ANDN U9006 ( .B(n5908), .A(n13863), .Z(n5911) );
  NANDN U9007 ( .A(x[1937]), .B(y[1937]), .Z(n5910) );
  NANDN U9008 ( .A(x[1936]), .B(y[1936]), .Z(n5909) );
  NAND U9009 ( .A(n5910), .B(n5909), .Z(n13865) );
  OR U9010 ( .A(n5911), .B(n13865), .Z(n5912) );
  AND U9011 ( .A(n13866), .B(n5912), .Z(n5915) );
  NANDN U9012 ( .A(x[1939]), .B(y[1939]), .Z(n5914) );
  NANDN U9013 ( .A(x[1938]), .B(y[1938]), .Z(n5913) );
  NAND U9014 ( .A(n5914), .B(n5913), .Z(n13868) );
  OR U9015 ( .A(n5915), .B(n13868), .Z(n5916) );
  AND U9016 ( .A(n13870), .B(n5916), .Z(n5918) );
  NANDN U9017 ( .A(x[1940]), .B(y[1940]), .Z(n5917) );
  ANDN U9018 ( .B(y[1941]), .A(x[1941]), .Z(n9784) );
  ANDN U9019 ( .B(n5917), .A(n9784), .Z(n13873) );
  NANDN U9020 ( .A(n5918), .B(n13873), .Z(n5921) );
  NANDN U9021 ( .A(y[1942]), .B(x[1942]), .Z(n5920) );
  NANDN U9022 ( .A(y[1941]), .B(x[1941]), .Z(n5919) );
  NAND U9023 ( .A(n5920), .B(n5919), .Z(n13875) );
  ANDN U9024 ( .B(n5921), .A(n13875), .Z(n5924) );
  NANDN U9025 ( .A(x[1943]), .B(y[1943]), .Z(n5923) );
  NANDN U9026 ( .A(x[1942]), .B(y[1942]), .Z(n5922) );
  NAND U9027 ( .A(n5923), .B(n5922), .Z(n13877) );
  OR U9028 ( .A(n5924), .B(n13877), .Z(n5925) );
  AND U9029 ( .A(n13878), .B(n5925), .Z(n5928) );
  NANDN U9030 ( .A(x[1945]), .B(y[1945]), .Z(n5927) );
  NANDN U9031 ( .A(x[1944]), .B(y[1944]), .Z(n5926) );
  NAND U9032 ( .A(n5927), .B(n5926), .Z(n13880) );
  OR U9033 ( .A(n5928), .B(n13880), .Z(n5931) );
  NANDN U9034 ( .A(y[1945]), .B(x[1945]), .Z(n5930) );
  NANDN U9035 ( .A(y[1946]), .B(x[1946]), .Z(n5929) );
  AND U9036 ( .A(n5930), .B(n5929), .Z(n13882) );
  NAND U9037 ( .A(n5931), .B(n13882), .Z(n5934) );
  NANDN U9038 ( .A(x[1947]), .B(y[1947]), .Z(n5933) );
  NANDN U9039 ( .A(x[1946]), .B(y[1946]), .Z(n5932) );
  NAND U9040 ( .A(n5933), .B(n5932), .Z(n13885) );
  ANDN U9041 ( .B(n5934), .A(n13885), .Z(n5937) );
  NANDN U9042 ( .A(y[1948]), .B(x[1948]), .Z(n5936) );
  NANDN U9043 ( .A(y[1947]), .B(x[1947]), .Z(n5935) );
  AND U9044 ( .A(n5936), .B(n5935), .Z(n13886) );
  NANDN U9045 ( .A(n5937), .B(n13886), .Z(n5938) );
  AND U9046 ( .A(n13894), .B(n5938), .Z(n5939) );
  NANDN U9047 ( .A(x[1948]), .B(y[1948]), .Z(n13888) );
  NAND U9048 ( .A(n5939), .B(n13888), .Z(n5940) );
  NANDN U9049 ( .A(n13891), .B(n5940), .Z(n5941) );
  AND U9050 ( .A(n13893), .B(n5941), .Z(n5943) );
  NANDN U9051 ( .A(x[1950]), .B(y[1950]), .Z(n5942) );
  NAND U9052 ( .A(n5943), .B(n5942), .Z(n5944) );
  AND U9053 ( .A(n13900), .B(n5944), .Z(n5947) );
  NANDN U9054 ( .A(x[1952]), .B(y[1952]), .Z(n5946) );
  NANDN U9055 ( .A(x[1953]), .B(y[1953]), .Z(n5945) );
  NAND U9056 ( .A(n5946), .B(n5945), .Z(n13902) );
  OR U9057 ( .A(n5947), .B(n13902), .Z(n5948) );
  NANDN U9058 ( .A(n13903), .B(n5948), .Z(n5949) );
  NANDN U9059 ( .A(n13904), .B(n5949), .Z(n5954) );
  NANDN U9060 ( .A(y[1956]), .B(x[1956]), .Z(n5951) );
  NANDN U9061 ( .A(y[1955]), .B(x[1955]), .Z(n5950) );
  AND U9062 ( .A(n5951), .B(n5950), .Z(n5953) );
  AND U9063 ( .A(n5953), .B(n5952), .Z(n13905) );
  NAND U9064 ( .A(n5954), .B(n13905), .Z(n5955) );
  NANDN U9065 ( .A(n9812), .B(n5955), .Z(n5956) );
  ANDN U9066 ( .B(x[1958]), .A(y[1958]), .Z(n13907) );
  ANDN U9067 ( .B(x[1959]), .A(y[1959]), .Z(n13911) );
  OR U9068 ( .A(n13907), .B(n13911), .Z(n9813) );
  ANDN U9069 ( .B(n5956), .A(n9813), .Z(n5959) );
  NANDN U9070 ( .A(x[1959]), .B(y[1959]), .Z(n13908) );
  NANDN U9071 ( .A(x[1960]), .B(y[1960]), .Z(n5957) );
  NANDN U9072 ( .A(n5958), .B(n5957), .Z(n13912) );
  ANDN U9073 ( .B(n13908), .A(n13912), .Z(n9815) );
  NANDN U9074 ( .A(n5959), .B(n9815), .Z(n5960) );
  NANDN U9075 ( .A(n9818), .B(n5960), .Z(n5963) );
  NANDN U9076 ( .A(x[1962]), .B(y[1962]), .Z(n5962) );
  NANDN U9077 ( .A(x[1963]), .B(y[1963]), .Z(n5961) );
  AND U9078 ( .A(n5962), .B(n5961), .Z(n13914) );
  NAND U9079 ( .A(n5963), .B(n13914), .Z(n5966) );
  NANDN U9080 ( .A(y[1964]), .B(x[1964]), .Z(n5965) );
  NANDN U9081 ( .A(y[1963]), .B(x[1963]), .Z(n5964) );
  NAND U9082 ( .A(n5965), .B(n5964), .Z(n13915) );
  ANDN U9083 ( .B(n5966), .A(n13915), .Z(n5969) );
  NANDN U9084 ( .A(x[1964]), .B(y[1964]), .Z(n5968) );
  NANDN U9085 ( .A(x[1965]), .B(y[1965]), .Z(n5967) );
  AND U9086 ( .A(n5968), .B(n5967), .Z(n13916) );
  NANDN U9087 ( .A(n5969), .B(n13916), .Z(n5970) );
  NANDN U9088 ( .A(n13917), .B(n5970), .Z(n5973) );
  NANDN U9089 ( .A(x[1966]), .B(y[1966]), .Z(n5972) );
  NANDN U9090 ( .A(x[1967]), .B(y[1967]), .Z(n5971) );
  AND U9091 ( .A(n5972), .B(n5971), .Z(n13918) );
  NAND U9092 ( .A(n5973), .B(n13918), .Z(n5974) );
  NANDN U9093 ( .A(n13919), .B(n5974), .Z(n5977) );
  NANDN U9094 ( .A(x[1969]), .B(y[1969]), .Z(n5976) );
  NANDN U9095 ( .A(x[1968]), .B(y[1968]), .Z(n5975) );
  AND U9096 ( .A(n5976), .B(n5975), .Z(n13920) );
  NAND U9097 ( .A(n5977), .B(n13920), .Z(n5978) );
  NANDN U9098 ( .A(y[1970]), .B(x[1970]), .Z(n9831) );
  NAND U9099 ( .A(n5978), .B(n9831), .Z(n5979) );
  NANDN U9100 ( .A(y[1969]), .B(x[1969]), .Z(n13923) );
  NANDN U9101 ( .A(n5979), .B(n13923), .Z(n5980) );
  AND U9102 ( .A(n13924), .B(n5980), .Z(n5981) );
  NAND U9103 ( .A(n5982), .B(n5981), .Z(n5983) );
  NAND U9104 ( .A(n5984), .B(n5983), .Z(n5985) );
  ANDN U9105 ( .B(y[1972]), .A(x[1972]), .Z(n9833) );
  ANDN U9106 ( .B(n5985), .A(n9833), .Z(n5988) );
  NANDN U9107 ( .A(y[1972]), .B(x[1972]), .Z(n5987) );
  NANDN U9108 ( .A(y[1973]), .B(x[1973]), .Z(n5986) );
  AND U9109 ( .A(n5987), .B(n5986), .Z(n13930) );
  NANDN U9110 ( .A(n5988), .B(n13930), .Z(n5989) );
  NANDN U9111 ( .A(n13933), .B(n5989), .Z(n5990) );
  AND U9112 ( .A(n9838), .B(n5990), .Z(n5991) );
  ANDN U9113 ( .B(y[1976]), .A(x[1976]), .Z(n9979) );
  NANDN U9114 ( .A(x[1975]), .B(y[1975]), .Z(n9980) );
  NANDN U9115 ( .A(n9979), .B(n9980), .Z(n9841) );
  OR U9116 ( .A(n5991), .B(n9841), .Z(n5992) );
  AND U9117 ( .A(n13941), .B(n5992), .Z(n5996) );
  NANDN U9118 ( .A(x[1978]), .B(y[1978]), .Z(n5994) );
  NANDN U9119 ( .A(x[1977]), .B(y[1977]), .Z(n5993) );
  NAND U9120 ( .A(n5994), .B(n5993), .Z(n9844) );
  ANDN U9121 ( .B(n5995), .A(n9844), .Z(n13942) );
  NANDN U9122 ( .A(n5996), .B(n13942), .Z(n5997) );
  NANDN U9123 ( .A(n13944), .B(n5997), .Z(n6000) );
  NANDN U9124 ( .A(x[1980]), .B(y[1980]), .Z(n5999) );
  NANDN U9125 ( .A(x[1981]), .B(y[1981]), .Z(n5998) );
  NAND U9126 ( .A(n5999), .B(n5998), .Z(n13947) );
  ANDN U9127 ( .B(n6000), .A(n13947), .Z(n6001) );
  OR U9128 ( .A(n13949), .B(n6001), .Z(n6002) );
  ANDN U9129 ( .B(y[1982]), .A(x[1982]), .Z(n9857) );
  ANDN U9130 ( .B(y[1983]), .A(x[1983]), .Z(n9862) );
  NOR U9131 ( .A(n9857), .B(n9862), .Z(n13950) );
  NAND U9132 ( .A(n6002), .B(n13950), .Z(n6003) );
  NANDN U9133 ( .A(y[1984]), .B(x[1984]), .Z(n9866) );
  NAND U9134 ( .A(n6003), .B(n9866), .Z(n6004) );
  NANDN U9135 ( .A(y[1983]), .B(x[1983]), .Z(n13952) );
  NANDN U9136 ( .A(n6004), .B(n13952), .Z(n6005) );
  AND U9137 ( .A(n13954), .B(n6005), .Z(n6006) );
  OR U9138 ( .A(n9865), .B(n6006), .Z(n6007) );
  NANDN U9139 ( .A(n13958), .B(n6007), .Z(n6008) );
  NANDN U9140 ( .A(y[1986]), .B(x[1986]), .Z(n13959) );
  NAND U9141 ( .A(n6008), .B(n13959), .Z(n6009) );
  AND U9142 ( .A(n13960), .B(n6009), .Z(n6012) );
  NANDN U9143 ( .A(y[1987]), .B(x[1987]), .Z(n6011) );
  NANDN U9144 ( .A(y[1988]), .B(x[1988]), .Z(n6010) );
  AND U9145 ( .A(n6011), .B(n6010), .Z(n13961) );
  NANDN U9146 ( .A(n6012), .B(n13961), .Z(n6015) );
  NANDN U9147 ( .A(x[1989]), .B(y[1989]), .Z(n6014) );
  NANDN U9148 ( .A(x[1988]), .B(y[1988]), .Z(n6013) );
  NAND U9149 ( .A(n6014), .B(n6013), .Z(n13962) );
  ANDN U9150 ( .B(n6015), .A(n13962), .Z(n6016) );
  NANDN U9151 ( .A(y[1989]), .B(x[1989]), .Z(n9978) );
  NANDN U9152 ( .A(n6016), .B(n9978), .Z(n6017) );
  AND U9153 ( .A(n13963), .B(n6017), .Z(n6018) );
  NANDN U9154 ( .A(y[1990]), .B(x[1990]), .Z(n9977) );
  ANDN U9155 ( .B(x[1991]), .A(y[1991]), .Z(n13964) );
  ANDN U9156 ( .B(n9977), .A(n13964), .Z(n9875) );
  NANDN U9157 ( .A(n6018), .B(n9875), .Z(n6019) );
  AND U9158 ( .A(n6111), .B(n6019), .Z(n6020) );
  NANDN U9159 ( .A(y[1992]), .B(x[1992]), .Z(n13966) );
  NANDN U9160 ( .A(n6020), .B(n13966), .Z(n6021) );
  AND U9161 ( .A(n6022), .B(n6021), .Z(n6024) );
  IV U9162 ( .A(x[1994]), .Z(n6109) );
  IV U9163 ( .A(y[1994]), .Z(n6108) );
  NANDN U9164 ( .A(n6109), .B(n6108), .Z(n6023) );
  ANDN U9165 ( .B(x[1993]), .A(y[1993]), .Z(n9879) );
  ANDN U9166 ( .B(n6023), .A(n9879), .Z(n13968) );
  NANDN U9167 ( .A(n6024), .B(n13968), .Z(n6025) );
  NANDN U9168 ( .A(n13969), .B(n6025), .Z(n6026) );
  NANDN U9169 ( .A(n13970), .B(n6026), .Z(n6027) );
  NANDN U9170 ( .A(n13971), .B(n6027), .Z(n6028) );
  AND U9171 ( .A(n6029), .B(n6028), .Z(n6030) );
  ANDN U9172 ( .B(n13973), .A(n6030), .Z(n6031) );
  NANDN U9173 ( .A(x[1999]), .B(y[1999]), .Z(n6102) );
  NAND U9174 ( .A(n6031), .B(n6102), .Z(n6032) );
  AND U9175 ( .A(n6099), .B(n6032), .Z(n6033) );
  NANDN U9176 ( .A(n6105), .B(n6033), .Z(n6035) );
  NANDN U9177 ( .A(x[2001]), .B(y[2001]), .Z(n6098) );
  NANDN U9178 ( .A(x[2000]), .B(y[2000]), .Z(n6034) );
  NAND U9179 ( .A(n6098), .B(n6034), .Z(n6103) );
  ANDN U9180 ( .B(n6035), .A(n6103), .Z(n6036) );
  OR U9181 ( .A(n6037), .B(n6036), .Z(n6040) );
  NANDN U9182 ( .A(x[2002]), .B(y[2002]), .Z(n6039) );
  NANDN U9183 ( .A(x[2003]), .B(y[2003]), .Z(n6038) );
  AND U9184 ( .A(n6039), .B(n6038), .Z(n13981) );
  NAND U9185 ( .A(n6040), .B(n13981), .Z(n6041) );
  NANDN U9186 ( .A(n13983), .B(n6041), .Z(n6042) );
  NANDN U9187 ( .A(n13984), .B(n6042), .Z(n6043) );
  AND U9188 ( .A(n13986), .B(n6043), .Z(n6046) );
  NANDN U9189 ( .A(x[2007]), .B(y[2007]), .Z(n6045) );
  NANDN U9190 ( .A(x[2006]), .B(y[2006]), .Z(n6044) );
  NAND U9191 ( .A(n6045), .B(n6044), .Z(n13988) );
  OR U9192 ( .A(n6046), .B(n13988), .Z(n6047) );
  AND U9193 ( .A(n13990), .B(n6047), .Z(n6050) );
  NANDN U9194 ( .A(x[2009]), .B(y[2009]), .Z(n6049) );
  NANDN U9195 ( .A(x[2008]), .B(y[2008]), .Z(n6048) );
  NAND U9196 ( .A(n6049), .B(n6048), .Z(n13992) );
  OR U9197 ( .A(n6050), .B(n13992), .Z(n6051) );
  AND U9198 ( .A(n13994), .B(n6051), .Z(n6053) );
  NANDN U9199 ( .A(x[2010]), .B(y[2010]), .Z(n6052) );
  ANDN U9200 ( .B(y[2011]), .A(x[2011]), .Z(n9911) );
  ANDN U9201 ( .B(n6052), .A(n9911), .Z(n13997) );
  NANDN U9202 ( .A(n6053), .B(n13997), .Z(n6054) );
  AND U9203 ( .A(n13998), .B(n6054), .Z(n6057) );
  NANDN U9204 ( .A(x[2013]), .B(y[2013]), .Z(n6056) );
  NANDN U9205 ( .A(x[2012]), .B(y[2012]), .Z(n6055) );
  NAND U9206 ( .A(n6056), .B(n6055), .Z(n14000) );
  OR U9207 ( .A(n6057), .B(n14000), .Z(n6060) );
  NANDN U9208 ( .A(y[2014]), .B(x[2014]), .Z(n6059) );
  NANDN U9209 ( .A(y[2013]), .B(x[2013]), .Z(n6058) );
  NAND U9210 ( .A(n6059), .B(n6058), .Z(n14003) );
  ANDN U9211 ( .B(n6060), .A(n14003), .Z(n6061) );
  OR U9212 ( .A(n14005), .B(n6061), .Z(n6062) );
  NANDN U9213 ( .A(n14007), .B(n6062), .Z(n6065) );
  NANDN U9214 ( .A(x[2017]), .B(y[2017]), .Z(n6064) );
  NANDN U9215 ( .A(x[2018]), .B(y[2018]), .Z(n6063) );
  AND U9216 ( .A(n6064), .B(n6063), .Z(n14009) );
  NAND U9217 ( .A(n6065), .B(n14009), .Z(n6066) );
  NANDN U9218 ( .A(n14011), .B(n6066), .Z(n6067) );
  NANDN U9219 ( .A(x[2019]), .B(y[2019]), .Z(n6095) );
  NAND U9220 ( .A(n6067), .B(n6095), .Z(n6068) );
  NANDN U9221 ( .A(y[2020]), .B(x[2020]), .Z(n14014) );
  NAND U9222 ( .A(n6068), .B(n14014), .Z(n6069) );
  NAND U9223 ( .A(n6070), .B(n6069), .Z(n6071) );
  NANDN U9224 ( .A(y[2021]), .B(x[2021]), .Z(n9921) );
  XOR U9225 ( .A(x[2022]), .B(y[2022]), .Z(n9925) );
  ANDN U9226 ( .B(n9921), .A(n9925), .Z(n14018) );
  NAND U9227 ( .A(n6071), .B(n14018), .Z(n6074) );
  NANDN U9228 ( .A(x[2022]), .B(y[2022]), .Z(n6073) );
  NANDN U9229 ( .A(x[2023]), .B(y[2023]), .Z(n6072) );
  NAND U9230 ( .A(n6073), .B(n6072), .Z(n14021) );
  ANDN U9231 ( .B(n6074), .A(n14021), .Z(n6075) );
  OR U9232 ( .A(n14022), .B(n6075), .Z(n6077) );
  NANDN U9233 ( .A(x[2024]), .B(y[2024]), .Z(n6076) );
  ANDN U9234 ( .B(y[2025]), .A(x[2025]), .Z(n9934) );
  ANDN U9235 ( .B(n6076), .A(n9934), .Z(n14024) );
  NAND U9236 ( .A(n6077), .B(n14024), .Z(n6078) );
  NANDN U9237 ( .A(n6079), .B(n6078), .Z(n6080) );
  NAND U9238 ( .A(n6081), .B(n6080), .Z(n6082) );
  AND U9239 ( .A(n14035), .B(n6082), .Z(n6083) );
  NANDN U9240 ( .A(n6084), .B(n6083), .Z(n6085) );
  AND U9241 ( .A(n14036), .B(n6085), .Z(n6086) );
  XNOR U9242 ( .A(x[2030]), .B(y[2030]), .Z(n9944) );
  ANDN U9243 ( .B(x[2029]), .A(y[2029]), .Z(n9942) );
  ANDN U9244 ( .B(n9944), .A(n9942), .Z(n14040) );
  NANDN U9245 ( .A(n6086), .B(n14040), .Z(n6087) );
  NANDN U9246 ( .A(n14043), .B(n6087), .Z(n6089) );
  NANDN U9247 ( .A(y[2032]), .B(x[2032]), .Z(n6088) );
  ANDN U9248 ( .B(x[2031]), .A(y[2031]), .Z(n9948) );
  ANDN U9249 ( .B(n6088), .A(n9948), .Z(n14044) );
  NAND U9250 ( .A(n6089), .B(n14044), .Z(n6090) );
  NANDN U9251 ( .A(x[2032]), .B(y[2032]), .Z(n9953) );
  ANDN U9252 ( .B(y[2033]), .A(x[2033]), .Z(n9959) );
  ANDN U9253 ( .B(n9953), .A(n9959), .Z(n14046) );
  NAND U9254 ( .A(n6090), .B(n14046), .Z(n6091) );
  NANDN U9255 ( .A(n14048), .B(n6091), .Z(n9967) );
  XNOR U9256 ( .A(y[2032]), .B(x[2032]), .Z(n9951) );
  NANDN U9257 ( .A(y[2030]), .B(x[2030]), .Z(n9947) );
  NAND U9258 ( .A(n6095), .B(n6094), .Z(n14013) );
  NOR U9259 ( .A(n14007), .B(n14003), .Z(n9916) );
  XNOR U9260 ( .A(x[2002]), .B(y[2002]), .Z(n6097) );
  AND U9261 ( .A(n6097), .B(n6096), .Z(n6101) );
  NANDN U9262 ( .A(n6099), .B(n6098), .Z(n6100) );
  NAND U9263 ( .A(n6101), .B(n6100), .Z(n13979) );
  NANDN U9264 ( .A(n6103), .B(n6102), .Z(n13977) );
  NOR U9265 ( .A(n6105), .B(n6104), .Z(n13974) );
  NANDN U9266 ( .A(y[1994]), .B(x[1994]), .Z(n6106) );
  AND U9267 ( .A(n6107), .B(n6106), .Z(n9885) );
  XNOR U9268 ( .A(n6109), .B(n6108), .Z(n9883) );
  NAND U9269 ( .A(n6111), .B(n6110), .Z(n13965) );
  NANDN U9270 ( .A(y[1980]), .B(x[1980]), .Z(n9852) );
  IV U9271 ( .A(n6112), .Z(n13827) );
  NANDN U9272 ( .A(x[1917]), .B(y[1917]), .Z(n6113) );
  AND U9273 ( .A(n9982), .B(n6113), .Z(n9744) );
  XNOR U9274 ( .A(n6115), .B(n6114), .Z(n9742) );
  NANDN U9275 ( .A(n6117), .B(n6116), .Z(n6118) );
  NANDN U9276 ( .A(n6119), .B(n6118), .Z(n13809) );
  NANDN U9277 ( .A(n6121), .B(n6120), .Z(n13808) );
  NAND U9278 ( .A(n6123), .B(n6122), .Z(n13806) );
  NAND U9279 ( .A(n6125), .B(n6124), .Z(n13805) );
  NOR U9280 ( .A(n6127), .B(n6126), .Z(n13802) );
  NANDN U9281 ( .A(n6129), .B(n6128), .Z(n6131) );
  NAND U9282 ( .A(n6131), .B(n6130), .Z(n13788) );
  AND U9283 ( .A(n13784), .B(n6132), .Z(n9707) );
  XNOR U9284 ( .A(y[1891]), .B(x[1891]), .Z(n9705) );
  ANDN U9285 ( .B(n6134), .A(n6133), .Z(n13756) );
  OR U9286 ( .A(n9983), .B(n13756), .Z(n9685) );
  NANDN U9287 ( .A(x[1877]), .B(y[1877]), .Z(n6135) );
  AND U9288 ( .A(n13752), .B(n6135), .Z(n9679) );
  XNOR U9289 ( .A(n6137), .B(n6136), .Z(n9677) );
  XOR U9290 ( .A(x[1876]), .B(n6138), .Z(n9673) );
  AND U9291 ( .A(n13742), .B(n6139), .Z(n9670) );
  ANDN U9292 ( .B(n9985), .A(n6140), .Z(n9662) );
  NANDN U9293 ( .A(x[1859]), .B(y[1859]), .Z(n6142) );
  NAND U9294 ( .A(n6142), .B(n6141), .Z(n13710) );
  OR U9295 ( .A(y[1859]), .B(n6143), .Z(n6144) );
  NAND U9296 ( .A(n6145), .B(n6144), .Z(n13709) );
  XNOR U9297 ( .A(x[1854]), .B(y[1854]), .Z(n9636) );
  NANDN U9298 ( .A(x[1837]), .B(y[1837]), .Z(n6146) );
  AND U9299 ( .A(n6147), .B(n6146), .Z(n9588) );
  XNOR U9300 ( .A(n6149), .B(n6148), .Z(n9586) );
  AND U9301 ( .A(n6151), .B(n6150), .Z(n9582) );
  XNOR U9302 ( .A(y[1835]), .B(x[1835]), .Z(n9580) );
  NANDN U9303 ( .A(y[1814]), .B(x[1814]), .Z(n6152) );
  AND U9304 ( .A(n13592), .B(n6152), .Z(n9525) );
  XNOR U9305 ( .A(n6154), .B(n6153), .Z(n9523) );
  XOR U9306 ( .A(y[1813]), .B(n6155), .Z(n9519) );
  XNOR U9307 ( .A(n6157), .B(n6156), .Z(n9515) );
  NAND U9308 ( .A(n6159), .B(n6158), .Z(n13579) );
  AND U9309 ( .A(n13574), .B(n6160), .Z(n9505) );
  XNOR U9310 ( .A(y[1807]), .B(x[1807]), .Z(n9503) );
  NANDN U9311 ( .A(x[1805]), .B(y[1805]), .Z(n6161) );
  AND U9312 ( .A(n6162), .B(n6161), .Z(n9499) );
  XNOR U9313 ( .A(n6164), .B(n6163), .Z(n9497) );
  OR U9314 ( .A(n6166), .B(n6165), .Z(n6167) );
  NANDN U9315 ( .A(n6168), .B(n6167), .Z(n13551) );
  NANDN U9316 ( .A(x[1789]), .B(y[1789]), .Z(n6170) );
  NANDN U9317 ( .A(x[1790]), .B(y[1790]), .Z(n6169) );
  NAND U9318 ( .A(n6170), .B(n6169), .Z(n13547) );
  NOR U9319 ( .A(n6172), .B(n6171), .Z(n13526) );
  AND U9320 ( .A(n13513), .B(n6173), .Z(n9423) );
  XNOR U9321 ( .A(x[1772]), .B(y[1772]), .Z(n9421) );
  NANDN U9322 ( .A(y[1770]), .B(x[1770]), .Z(n6174) );
  AND U9323 ( .A(n6175), .B(n6174), .Z(n9417) );
  XNOR U9324 ( .A(n6177), .B(n6176), .Z(n9415) );
  NANDN U9325 ( .A(y[1768]), .B(x[1768]), .Z(n6178) );
  AND U9326 ( .A(n6179), .B(n6178), .Z(n9411) );
  XNOR U9327 ( .A(n6181), .B(n6180), .Z(n9409) );
  NANDN U9328 ( .A(y[1764]), .B(x[1764]), .Z(n9394) );
  ANDN U9329 ( .B(n13490), .A(n6182), .Z(n9392) );
  ANDN U9330 ( .B(n13488), .A(n6183), .Z(n9390) );
  NAND U9331 ( .A(n6185), .B(n6184), .Z(n13487) );
  NOR U9332 ( .A(n6187), .B(n6186), .Z(n13484) );
  NANDN U9333 ( .A(x[1757]), .B(y[1757]), .Z(n6188) );
  AND U9334 ( .A(n6189), .B(n6188), .Z(n9380) );
  XNOR U9335 ( .A(n6191), .B(n6190), .Z(n9378) );
  OR U9336 ( .A(x[1754]), .B(n6192), .Z(n6193) );
  NAND U9337 ( .A(n6194), .B(n6193), .Z(n13463) );
  AND U9338 ( .A(n13456), .B(n13451), .Z(n9360) );
  AND U9339 ( .A(n13448), .B(n6195), .Z(n9358) );
  NAND U9340 ( .A(n6197), .B(n6196), .Z(n13447) );
  NANDN U9341 ( .A(y[1740]), .B(x[1740]), .Z(n9344) );
  XNOR U9342 ( .A(x[1740]), .B(y[1740]), .Z(n9342) );
  OR U9343 ( .A(y[1733]), .B(n6198), .Z(n6199) );
  NAND U9344 ( .A(n6200), .B(n6199), .Z(n13425) );
  NAND U9345 ( .A(n6201), .B(n13423), .Z(n6202) );
  NANDN U9346 ( .A(n6203), .B(n6202), .Z(n9316) );
  OR U9347 ( .A(y[1719]), .B(n6204), .Z(n6205) );
  NAND U9348 ( .A(n6206), .B(n6205), .Z(n13397) );
  IV U9349 ( .A(n6207), .Z(n9992) );
  NOR U9350 ( .A(n9992), .B(n6208), .Z(n9264) );
  NANDN U9351 ( .A(y[1702]), .B(x[1702]), .Z(n6209) );
  AND U9352 ( .A(n13354), .B(n6209), .Z(n9255) );
  XNOR U9353 ( .A(n6211), .B(n6210), .Z(n9253) );
  XOR U9354 ( .A(y[1701]), .B(n6212), .Z(n9249) );
  XNOR U9355 ( .A(n6214), .B(n6213), .Z(n9245) );
  AND U9356 ( .A(n13336), .B(n6215), .Z(n9232) );
  XNOR U9357 ( .A(y[1695]), .B(x[1695]), .Z(n9230) );
  OR U9358 ( .A(y[1691]), .B(n6216), .Z(n6217) );
  NAND U9359 ( .A(n6218), .B(n6217), .Z(n13323) );
  NANDN U9360 ( .A(y[1688]), .B(x[1688]), .Z(n6219) );
  AND U9361 ( .A(n13318), .B(n6219), .Z(n9213) );
  XNOR U9362 ( .A(n6221), .B(n6220), .Z(n9211) );
  AND U9363 ( .A(n6223), .B(n6222), .Z(n9207) );
  XNOR U9364 ( .A(x[1686]), .B(y[1686]), .Z(n9205) );
  NANDN U9365 ( .A(y[1684]), .B(x[1684]), .Z(n6224) );
  AND U9366 ( .A(n6225), .B(n6224), .Z(n9201) );
  XNOR U9367 ( .A(n6227), .B(n6226), .Z(n9199) );
  NANDN U9368 ( .A(y[1682]), .B(x[1682]), .Z(n6228) );
  AND U9369 ( .A(n6229), .B(n6228), .Z(n9195) );
  XNOR U9370 ( .A(n6231), .B(n6230), .Z(n9193) );
  ANDN U9371 ( .B(n6233), .A(n6232), .Z(n9171) );
  XOR U9372 ( .A(x[1673]), .B(n6234), .Z(n9169) );
  ANDN U9373 ( .B(y[1671]), .A(x[1671]), .Z(n6240) );
  NANDN U9374 ( .A(n6236), .B(n6235), .Z(n6237) );
  NANDN U9375 ( .A(n6238), .B(n6237), .Z(n6239) );
  NANDN U9376 ( .A(n6240), .B(n6239), .Z(n13275) );
  AND U9377 ( .A(n13270), .B(n6241), .Z(n9160) );
  XNOR U9378 ( .A(y[1667]), .B(x[1667]), .Z(n9158) );
  XOR U9379 ( .A(x[1666]), .B(n6242), .Z(n9154) );
  XNOR U9380 ( .A(y[1653]), .B(x[1653]), .Z(n9129) );
  XNOR U9381 ( .A(x[1652]), .B(y[1652]), .Z(n9125) );
  ANDN U9382 ( .B(n6243), .A(n13231), .Z(n9122) );
  NANDN U9383 ( .A(x[1649]), .B(y[1649]), .Z(n6245) );
  NAND U9384 ( .A(n6245), .B(n6244), .Z(n13229) );
  NANDN U9385 ( .A(y[1649]), .B(x[1649]), .Z(n6247) );
  ANDN U9386 ( .B(n6247), .A(n6246), .Z(n13226) );
  NANDN U9387 ( .A(x[1645]), .B(y[1645]), .Z(n6248) );
  AND U9388 ( .A(n6249), .B(n6248), .Z(n9112) );
  XNOR U9389 ( .A(n6251), .B(n6250), .Z(n9110) );
  NAND U9390 ( .A(n6253), .B(n6252), .Z(n13181) );
  ANDN U9391 ( .B(y[1623]), .A(x[1623]), .Z(n13165) );
  NANDN U9392 ( .A(n13165), .B(n13170), .Z(n9068) );
  NAND U9393 ( .A(n6255), .B(n6254), .Z(n13163) );
  NANDN U9394 ( .A(n6257), .B(n6256), .Z(n6258) );
  NAND U9395 ( .A(n6259), .B(n6258), .Z(n13159) );
  OR U9396 ( .A(y[1619]), .B(n6260), .Z(n6261) );
  NAND U9397 ( .A(n6262), .B(n6261), .Z(n13154) );
  ANDN U9398 ( .B(n13149), .A(n6263), .Z(n9054) );
  NAND U9399 ( .A(n6265), .B(n6264), .Z(n13125) );
  OR U9400 ( .A(n6267), .B(n6266), .Z(n6269) );
  NAND U9401 ( .A(n6269), .B(n6268), .Z(n13112) );
  NANDN U9402 ( .A(n6271), .B(n6270), .Z(n6273) );
  NAND U9403 ( .A(n6273), .B(n6272), .Z(n13089) );
  NAND U9404 ( .A(n6275), .B(n6274), .Z(n13073) );
  ANDN U9405 ( .B(n13066), .A(n6276), .Z(n8993) );
  NANDN U9406 ( .A(n13061), .B(n13065), .Z(n8991) );
  NANDN U9407 ( .A(x[1578]), .B(y[1578]), .Z(n6278) );
  NAND U9408 ( .A(n6278), .B(n6277), .Z(n13055) );
  NANDN U9409 ( .A(n6280), .B(n6279), .Z(n6281) );
  NAND U9410 ( .A(n6282), .B(n6281), .Z(n13045) );
  NANDN U9411 ( .A(x[1571]), .B(y[1571]), .Z(n6284) );
  NAND U9412 ( .A(n6284), .B(n6283), .Z(n13042) );
  NAND U9413 ( .A(n13000), .B(n13005), .Z(n8939) );
  NAND U9414 ( .A(n6286), .B(n6285), .Z(n12985) );
  NANDN U9415 ( .A(n6288), .B(n6287), .Z(n6290) );
  NAND U9416 ( .A(n6290), .B(n6289), .Z(n12977) );
  NANDN U9417 ( .A(n12942), .B(n12945), .Z(n8890) );
  OR U9418 ( .A(x[1530]), .B(n6291), .Z(n6292) );
  NAND U9419 ( .A(n6293), .B(n6292), .Z(n12936) );
  ANDN U9420 ( .B(n12909), .A(n6294), .Z(n8856) );
  NANDN U9421 ( .A(y[1500]), .B(x[1500]), .Z(n6296) );
  NAND U9422 ( .A(n6296), .B(n6295), .Z(n12884) );
  NANDN U9423 ( .A(x[1500]), .B(y[1500]), .Z(n6297) );
  NAND U9424 ( .A(n6298), .B(n6297), .Z(n12882) );
  NANDN U9425 ( .A(n12872), .B(n12876), .Z(n8819) );
  NANDN U9426 ( .A(y[1487]), .B(x[1487]), .Z(n6302) );
  NANDN U9427 ( .A(y[1486]), .B(x[1486]), .Z(n6301) );
  NAND U9428 ( .A(n6302), .B(n6301), .Z(n12856) );
  OR U9429 ( .A(x[1486]), .B(n6303), .Z(n6306) );
  NAND U9430 ( .A(n8797), .B(n6304), .Z(n6305) );
  NAND U9431 ( .A(n6306), .B(n6305), .Z(n12854) );
  NANDN U9432 ( .A(y[1476]), .B(x[1476]), .Z(n6308) );
  NAND U9433 ( .A(n6308), .B(n6307), .Z(n12840) );
  OR U9434 ( .A(x[1476]), .B(n6309), .Z(n6310) );
  NAND U9435 ( .A(n6311), .B(n6310), .Z(n12838) );
  OR U9436 ( .A(n6313), .B(n6312), .Z(n6314) );
  NANDN U9437 ( .A(n6315), .B(n6314), .Z(n12831) );
  NANDN U9438 ( .A(n6317), .B(n6316), .Z(n12790) );
  ANDN U9439 ( .B(n12785), .A(n6318), .Z(n8747) );
  OR U9440 ( .A(n6320), .B(n6319), .Z(n12777) );
  AND U9441 ( .A(n12749), .B(n12745), .Z(n8719) );
  NANDN U9442 ( .A(n6322), .B(n6321), .Z(n6323) );
  NAND U9443 ( .A(n6324), .B(n6323), .Z(n12728) );
  NAND U9444 ( .A(n8692), .B(n6325), .Z(n6326) );
  NANDN U9445 ( .A(n6327), .B(n6326), .Z(n12724) );
  NAND U9446 ( .A(n6329), .B(n6328), .Z(n12705) );
  NANDN U9447 ( .A(y[1404]), .B(x[1404]), .Z(n6330) );
  NAND U9448 ( .A(n6331), .B(n6330), .Z(n12686) );
  NANDN U9449 ( .A(x[1398]), .B(y[1398]), .Z(n6332) );
  NAND U9450 ( .A(n6333), .B(n6332), .Z(n12667) );
  AND U9451 ( .A(n12649), .B(n12645), .Z(n8624) );
  OR U9452 ( .A(y[1381]), .B(n6334), .Z(n6335) );
  NAND U9453 ( .A(n6336), .B(n6335), .Z(n12630) );
  OR U9454 ( .A(y[1378]), .B(n6337), .Z(n6341) );
  NANDN U9455 ( .A(n6339), .B(n6338), .Z(n6340) );
  NAND U9456 ( .A(n6341), .B(n6340), .Z(n12626) );
  OR U9457 ( .A(n6343), .B(n6342), .Z(n6345) );
  NAND U9458 ( .A(n6345), .B(n6344), .Z(n12621) );
  NAND U9459 ( .A(n6347), .B(n6346), .Z(n12582) );
  NAND U9460 ( .A(n12573), .B(n12578), .Z(n8563) );
  ANDN U9461 ( .B(n12545), .A(n12549), .Z(n8536) );
  ANDN U9462 ( .B(n6348), .A(n12520), .Z(n8513) );
  NANDN U9463 ( .A(x[1319]), .B(y[1319]), .Z(n6350) );
  NANDN U9464 ( .A(x[1320]), .B(y[1320]), .Z(n6349) );
  NAND U9465 ( .A(n6350), .B(n6349), .Z(n12504) );
  OR U9466 ( .A(y[1319]), .B(n6351), .Z(n6352) );
  NAND U9467 ( .A(n6353), .B(n6352), .Z(n12502) );
  NOR U9468 ( .A(n12500), .B(n6354), .Z(n8500) );
  NANDN U9469 ( .A(n6356), .B(n6355), .Z(n6357) );
  NAND U9470 ( .A(n6358), .B(n6357), .Z(n12478) );
  ANDN U9471 ( .B(n12471), .A(n6359), .Z(n8476) );
  NANDN U9472 ( .A(x[1297]), .B(y[1297]), .Z(n6361) );
  NAND U9473 ( .A(n6361), .B(n6360), .Z(n12451) );
  NAND U9474 ( .A(n6363), .B(n6362), .Z(n12446) );
  NANDN U9475 ( .A(n12438), .B(n12441), .Z(n8451) );
  NANDN U9476 ( .A(x[1290]), .B(y[1290]), .Z(n6365) );
  NAND U9477 ( .A(n6365), .B(n6364), .Z(n12432) );
  NANDN U9478 ( .A(y[1284]), .B(x[1284]), .Z(n6367) );
  NAND U9479 ( .A(n6367), .B(n6366), .Z(n12422) );
  AND U9480 ( .A(n12413), .B(n6368), .Z(n8428) );
  XNOR U9481 ( .A(x[1280]), .B(y[1280]), .Z(n8426) );
  NANDN U9482 ( .A(y[1275]), .B(x[1275]), .Z(n6369) );
  NAND U9483 ( .A(n6370), .B(n6369), .Z(n12401) );
  NANDN U9484 ( .A(n6372), .B(n6371), .Z(n6373) );
  NAND U9485 ( .A(n6374), .B(n6373), .Z(n12398) );
  NANDN U9486 ( .A(y[1270]), .B(x[1270]), .Z(n6376) );
  NANDN U9487 ( .A(y[1271]), .B(x[1271]), .Z(n6375) );
  NAND U9488 ( .A(n6376), .B(n6375), .Z(n12394) );
  OR U9489 ( .A(x[1270]), .B(n6377), .Z(n6381) );
  NANDN U9490 ( .A(n6379), .B(n6378), .Z(n6380) );
  NAND U9491 ( .A(n6381), .B(n6380), .Z(n12391) );
  NOR U9492 ( .A(n6382), .B(n12384), .Z(n8389) );
  OR U9493 ( .A(n6384), .B(n6383), .Z(n12380) );
  NANDN U9494 ( .A(y[1248]), .B(x[1248]), .Z(n6386) );
  NAND U9495 ( .A(n6386), .B(n6385), .Z(n12371) );
  NANDN U9496 ( .A(n6388), .B(n6387), .Z(n6389) );
  NAND U9497 ( .A(n6390), .B(n6389), .Z(n12370) );
  NAND U9498 ( .A(n12359), .B(n12364), .Z(n8362) );
  NANDN U9499 ( .A(n6392), .B(n6391), .Z(n6393) );
  NAND U9500 ( .A(n6394), .B(n6393), .Z(n12334) );
  ANDN U9501 ( .B(n12330), .A(n6395), .Z(n8340) );
  NANDN U9502 ( .A(y[1223]), .B(x[1223]), .Z(n6396) );
  NAND U9503 ( .A(n6397), .B(n6396), .Z(n12317) );
  ANDN U9504 ( .B(n6398), .A(n12314), .Z(n8318) );
  NAND U9505 ( .A(n6399), .B(n12316), .Z(n12313) );
  ANDN U9506 ( .B(n12311), .A(n6400), .Z(n8315) );
  ANDN U9507 ( .B(n12292), .A(n6401), .Z(n8304) );
  NAND U9508 ( .A(n6403), .B(n6402), .Z(n12281) );
  NANDN U9509 ( .A(x[1187]), .B(y[1187]), .Z(n6405) );
  NAND U9510 ( .A(n6405), .B(n6404), .Z(n12244) );
  NANDN U9511 ( .A(y[1187]), .B(x[1187]), .Z(n6406) );
  NAND U9512 ( .A(n6407), .B(n6406), .Z(n12241) );
  NAND U9513 ( .A(n12233), .B(n12238), .Z(n8258) );
  NANDN U9514 ( .A(x[1181]), .B(y[1181]), .Z(n6408) );
  AND U9515 ( .A(n6409), .B(n6408), .Z(n8250) );
  XNOR U9516 ( .A(n6411), .B(n6410), .Z(n8248) );
  OR U9517 ( .A(x[1175]), .B(n6412), .Z(n6413) );
  NAND U9518 ( .A(n6414), .B(n6413), .Z(n12216) );
  NANDN U9519 ( .A(y[1175]), .B(x[1175]), .Z(n6415) );
  NAND U9520 ( .A(n6416), .B(n6415), .Z(n12213) );
  NANDN U9521 ( .A(y[1164]), .B(x[1164]), .Z(n6418) );
  NANDN U9522 ( .A(y[1165]), .B(x[1165]), .Z(n6417) );
  NAND U9523 ( .A(n6418), .B(n6417), .Z(n12190) );
  OR U9524 ( .A(x[1164]), .B(n6419), .Z(n6420) );
  NAND U9525 ( .A(n6421), .B(n6420), .Z(n12188) );
  NAND U9526 ( .A(n12177), .B(n12182), .Z(n8209) );
  NANDN U9527 ( .A(n6423), .B(n6422), .Z(n6424) );
  NAND U9528 ( .A(n6425), .B(n6424), .Z(n12172) );
  NANDN U9529 ( .A(y[1152]), .B(x[1152]), .Z(n6426) );
  NAND U9530 ( .A(n6427), .B(n6426), .Z(n12160) );
  NAND U9531 ( .A(n6429), .B(n6428), .Z(n12150) );
  ANDN U9532 ( .B(n12148), .A(n12145), .Z(n8173) );
  NANDN U9533 ( .A(x[1139]), .B(y[1139]), .Z(n6431) );
  NANDN U9534 ( .A(x[1140]), .B(y[1140]), .Z(n6430) );
  NAND U9535 ( .A(n6431), .B(n6430), .Z(n12142) );
  NANDN U9536 ( .A(n6433), .B(n6432), .Z(n6434) );
  NAND U9537 ( .A(n6435), .B(n6434), .Z(n12120) );
  NOR U9538 ( .A(n6437), .B(n6436), .Z(n8110) );
  NANDN U9539 ( .A(x[1104]), .B(y[1104]), .Z(n6438) );
  NAND U9540 ( .A(n6439), .B(n6438), .Z(n12072) );
  AND U9541 ( .A(n12061), .B(n12065), .Z(n8092) );
  NANDN U9542 ( .A(y[1098]), .B(x[1098]), .Z(n6442) );
  NAND U9543 ( .A(n6442), .B(n6441), .Z(n12057) );
  NANDN U9544 ( .A(n6445), .B(n6444), .Z(n6446) );
  NAND U9545 ( .A(n6447), .B(n6446), .Z(n12048) );
  ANDN U9546 ( .B(n12043), .A(n6448), .Z(n8077) );
  NANDN U9547 ( .A(x[1067]), .B(y[1067]), .Z(n6450) );
  NANDN U9548 ( .A(x[1068]), .B(y[1068]), .Z(n6449) );
  NAND U9549 ( .A(n6450), .B(n6449), .Z(n11994) );
  OR U9550 ( .A(y[1067]), .B(n6451), .Z(n6452) );
  NAND U9551 ( .A(n6453), .B(n6452), .Z(n11991) );
  NANDN U9552 ( .A(y[1056]), .B(x[1056]), .Z(n6455) );
  ANDN U9553 ( .B(n6455), .A(n6454), .Z(n11967) );
  NANDN U9554 ( .A(x[1056]), .B(y[1056]), .Z(n6456) );
  NAND U9555 ( .A(n6457), .B(n6456), .Z(n11965) );
  OR U9556 ( .A(n11956), .B(n11960), .Z(n8008) );
  NAND U9557 ( .A(n6459), .B(n6458), .Z(n11950) );
  NANDN U9558 ( .A(x[1045]), .B(y[1045]), .Z(n6461) );
  NAND U9559 ( .A(n6461), .B(n6460), .Z(n11941) );
  NAND U9560 ( .A(n6463), .B(n6462), .Z(n11940) );
  NANDN U9561 ( .A(x[1033]), .B(y[1033]), .Z(n6464) );
  NAND U9562 ( .A(n6465), .B(n6464), .Z(n11918) );
  NANDN U9563 ( .A(y[1033]), .B(x[1033]), .Z(n6466) );
  NAND U9564 ( .A(n6467), .B(n6466), .Z(n11916) );
  NAND U9565 ( .A(n6469), .B(n6468), .Z(n11912) );
  AND U9566 ( .A(n11904), .B(n11908), .Z(n7971) );
  NAND U9567 ( .A(n6471), .B(n6470), .Z(n11900) );
  NANDN U9568 ( .A(y[1006]), .B(x[1006]), .Z(n6472) );
  AND U9569 ( .A(n11853), .B(n6472), .Z(n7933) );
  XNOR U9570 ( .A(n6474), .B(n6473), .Z(n7931) );
  NANDN U9571 ( .A(y[946]), .B(x[946]), .Z(n6475) );
  AND U9572 ( .A(n11701), .B(n6475), .Z(n7851) );
  XNOR U9573 ( .A(n6477), .B(n6476), .Z(n7849) );
  ANDN U9574 ( .B(n6479), .A(n6478), .Z(n11690) );
  AND U9575 ( .A(n11643), .B(n6480), .Z(n7817) );
  XOR U9576 ( .A(y[922]), .B(n6481), .Z(n7815) );
  NANDN U9577 ( .A(y[874]), .B(x[874]), .Z(n6482) );
  AND U9578 ( .A(n11517), .B(n6482), .Z(n7754) );
  XNOR U9579 ( .A(n6484), .B(n6483), .Z(n7752) );
  NANDN U9580 ( .A(y[862]), .B(x[862]), .Z(n6485) );
  AND U9581 ( .A(n11487), .B(n6485), .Z(n7734) );
  XNOR U9582 ( .A(n6487), .B(n6486), .Z(n7732) );
  NANDN U9583 ( .A(y[850]), .B(x[850]), .Z(n6488) );
  AND U9584 ( .A(n11457), .B(n6488), .Z(n7714) );
  XNOR U9585 ( .A(n6490), .B(n6489), .Z(n7712) );
  AND U9586 ( .A(n6492), .B(n6491), .Z(n7684) );
  XNOR U9587 ( .A(y[834]), .B(x[834]), .Z(n7682) );
  NANDN U9588 ( .A(x[824]), .B(y[824]), .Z(n6493) );
  AND U9589 ( .A(n6494), .B(n6493), .Z(n6496) );
  NOR U9590 ( .A(n6496), .B(n6495), .Z(n11406) );
  NAND U9591 ( .A(n6498), .B(n6497), .Z(n11387) );
  NANDN U9592 ( .A(y[810]), .B(x[810]), .Z(n6500) );
  NAND U9593 ( .A(n6500), .B(n6499), .Z(n11386) );
  OR U9594 ( .A(n6502), .B(n6501), .Z(n11266) );
  NANDN U9595 ( .A(x[712]), .B(y[712]), .Z(n6503) );
  AND U9596 ( .A(n6504), .B(n6503), .Z(n6505) );
  ANDN U9597 ( .B(n6506), .A(n6505), .Z(n11180) );
  NAND U9598 ( .A(n11171), .B(n11175), .Z(n6507) );
  NANDN U9599 ( .A(n6508), .B(n6507), .Z(n7508) );
  NOR U9600 ( .A(n6510), .B(n6509), .Z(n7443) );
  NANDN U9601 ( .A(x[620]), .B(y[620]), .Z(n6511) );
  AND U9602 ( .A(n6512), .B(n6511), .Z(n6513) );
  OR U9603 ( .A(n6514), .B(n6513), .Z(n6515) );
  NANDN U9604 ( .A(n6516), .B(n6515), .Z(n11069) );
  NANDN U9605 ( .A(x[595]), .B(y[595]), .Z(n6517) );
  AND U9606 ( .A(n6518), .B(n6517), .Z(n7366) );
  XNOR U9607 ( .A(n6520), .B(n6519), .Z(n7364) );
  ANDN U9608 ( .B(n6522), .A(n6521), .Z(n7358) );
  NOR U9609 ( .A(n6524), .B(n6523), .Z(n7289) );
  OR U9610 ( .A(n6526), .B(n6525), .Z(n6528) );
  NAND U9611 ( .A(n6528), .B(n6527), .Z(n10921) );
  ANDN U9612 ( .B(y[522]), .A(x[522]), .Z(n7267) );
  NAND U9613 ( .A(n6530), .B(n6529), .Z(n10893) );
  NOR U9614 ( .A(n6531), .B(n10810), .Z(n7213) );
  NANDN U9615 ( .A(y[434]), .B(x[434]), .Z(n6532) );
  AND U9616 ( .A(n10761), .B(n6532), .Z(n7187) );
  XNOR U9617 ( .A(n6534), .B(n6533), .Z(n7185) );
  ANDN U9618 ( .B(n6536), .A(n6535), .Z(n6537) );
  ANDN U9619 ( .B(n6538), .A(n6537), .Z(n10740) );
  NANDN U9620 ( .A(n6540), .B(n6539), .Z(n6542) );
  NAND U9621 ( .A(n6542), .B(n6541), .Z(n10708) );
  ANDN U9622 ( .B(n6544), .A(n6543), .Z(n6546) );
  NANDN U9623 ( .A(n6546), .B(n6545), .Z(n6547) );
  NANDN U9624 ( .A(n6548), .B(n6547), .Z(n10706) );
  NANDN U9625 ( .A(n6550), .B(n6549), .Z(n10704) );
  ANDN U9626 ( .B(n6552), .A(n6551), .Z(n6553) );
  NOR U9627 ( .A(n6554), .B(n6553), .Z(n10697) );
  ANDN U9628 ( .B(n10602), .A(n6555), .Z(n7070) );
  NAND U9629 ( .A(n10598), .B(n10601), .Z(n7068) );
  ANDN U9630 ( .B(n10035), .A(n6556), .Z(n7066) );
  NAND U9631 ( .A(n6558), .B(n6557), .Z(n6560) );
  NAND U9632 ( .A(n6560), .B(n6559), .Z(n10575) );
  NAND U9633 ( .A(n10465), .B(n10471), .Z(n6984) );
  ANDN U9634 ( .B(n10417), .A(n6561), .Z(n6947) );
  NANDN U9635 ( .A(x[196]), .B(y[196]), .Z(n6562) );
  AND U9636 ( .A(n6563), .B(n6562), .Z(n6564) );
  ANDN U9637 ( .B(n6565), .A(n6564), .Z(n10355) );
  NANDN U9638 ( .A(x[122]), .B(y[122]), .Z(n6811) );
  XNOR U9639 ( .A(n6567), .B(n6566), .Z(n6809) );
  NANDN U9640 ( .A(y[105]), .B(x[105]), .Z(n6568) );
  NAND U9641 ( .A(n6569), .B(n6568), .Z(n10199) );
  ANDN U9642 ( .B(x[40]), .A(y[40]), .Z(n6695) );
  NANDN U9643 ( .A(n6571), .B(n6570), .Z(n6641) );
  AND U9644 ( .A(n6573), .B(n6572), .Z(n6635) );
  AND U9645 ( .A(n6575), .B(n6574), .Z(n6613) );
  AND U9646 ( .A(n6577), .B(n6576), .Z(n6597) );
  NANDN U9647 ( .A(y[0]), .B(x[0]), .Z(n6578) );
  NANDN U9648 ( .A(n6579), .B(n6578), .Z(n6580) );
  AND U9649 ( .A(n6581), .B(n6580), .Z(n6583) );
  NAND U9650 ( .A(n6583), .B(n6582), .Z(n6585) );
  ANDN U9651 ( .B(n6585), .A(n6584), .Z(n6586) );
  NANDN U9652 ( .A(n6587), .B(n6586), .Z(n6589) );
  AND U9653 ( .A(n6589), .B(n6588), .Z(n6591) );
  NAND U9654 ( .A(n6591), .B(n6590), .Z(n6592) );
  NANDN U9655 ( .A(n6593), .B(n6592), .Z(n6594) );
  OR U9656 ( .A(n6595), .B(n6594), .Z(n6596) );
  AND U9657 ( .A(n6597), .B(n6596), .Z(n6598) );
  OR U9658 ( .A(n6599), .B(n6598), .Z(n6601) );
  NAND U9659 ( .A(n6601), .B(n6600), .Z(n6602) );
  NANDN U9660 ( .A(n6603), .B(n6602), .Z(n6604) );
  AND U9661 ( .A(n6605), .B(n6604), .Z(n6607) );
  NAND U9662 ( .A(n6607), .B(n6606), .Z(n6608) );
  NANDN U9663 ( .A(n6609), .B(n6608), .Z(n6610) );
  OR U9664 ( .A(n6611), .B(n6610), .Z(n6612) );
  AND U9665 ( .A(n6613), .B(n6612), .Z(n6617) );
  ANDN U9666 ( .B(n6615), .A(n6614), .Z(n6616) );
  NANDN U9667 ( .A(n6617), .B(n6616), .Z(n6618) );
  AND U9668 ( .A(n6619), .B(n6618), .Z(n6621) );
  NAND U9669 ( .A(n6621), .B(n6620), .Z(n6623) );
  ANDN U9670 ( .B(n6623), .A(n6622), .Z(n6624) );
  NANDN U9671 ( .A(n6625), .B(n6624), .Z(n6627) );
  AND U9672 ( .A(n6627), .B(n6626), .Z(n6629) );
  NAND U9673 ( .A(n6629), .B(n6628), .Z(n6630) );
  NANDN U9674 ( .A(n6631), .B(n6630), .Z(n6632) );
  OR U9675 ( .A(n6633), .B(n6632), .Z(n6634) );
  AND U9676 ( .A(n6635), .B(n6634), .Z(n6639) );
  ANDN U9677 ( .B(n6637), .A(n6636), .Z(n6638) );
  NANDN U9678 ( .A(n6639), .B(n6638), .Z(n6640) );
  AND U9679 ( .A(n6641), .B(n6640), .Z(n6643) );
  NAND U9680 ( .A(n6643), .B(n6642), .Z(n6647) );
  NANDN U9681 ( .A(y[20]), .B(x[20]), .Z(n6645) );
  ANDN U9682 ( .B(n6645), .A(n6644), .Z(n6646) );
  NAND U9683 ( .A(n6647), .B(n6646), .Z(n6648) );
  AND U9684 ( .A(n6649), .B(n6648), .Z(n6650) );
  OR U9685 ( .A(n6651), .B(n6650), .Z(n6652) );
  AND U9686 ( .A(n6653), .B(n6652), .Z(n6655) );
  NANDN U9687 ( .A(x[24]), .B(y[24]), .Z(n6654) );
  NAND U9688 ( .A(n6655), .B(n6654), .Z(n6661) );
  NANDN U9689 ( .A(n6657), .B(n6656), .Z(n6659) );
  ANDN U9690 ( .B(n6659), .A(n6658), .Z(n6660) );
  NAND U9691 ( .A(n6661), .B(n6660), .Z(n6663) );
  ANDN U9692 ( .B(n6663), .A(n6662), .Z(n6665) );
  NAND U9693 ( .A(n6665), .B(n6664), .Z(n6666) );
  NANDN U9694 ( .A(n6667), .B(n6666), .Z(n6668) );
  AND U9695 ( .A(n6669), .B(n6668), .Z(n6670) );
  OR U9696 ( .A(n6671), .B(n6670), .Z(n6673) );
  NAND U9697 ( .A(n6673), .B(n6672), .Z(n6674) );
  NANDN U9698 ( .A(n6675), .B(n6674), .Z(n6676) );
  NANDN U9699 ( .A(n6677), .B(n6676), .Z(n6678) );
  NANDN U9700 ( .A(n6679), .B(n6678), .Z(n6680) );
  AND U9701 ( .A(n6681), .B(n6680), .Z(n6682) );
  OR U9702 ( .A(n6683), .B(n6682), .Z(n6684) );
  NANDN U9703 ( .A(n6685), .B(n6684), .Z(n6686) );
  NANDN U9704 ( .A(n6687), .B(n6686), .Z(n6689) );
  NAND U9705 ( .A(n6689), .B(n6688), .Z(n6690) );
  NANDN U9706 ( .A(n6691), .B(n6690), .Z(n6692) );
  AND U9707 ( .A(n6693), .B(n6692), .Z(n6694) );
  OR U9708 ( .A(n6695), .B(n6694), .Z(n6701) );
  NANDN U9709 ( .A(n6697), .B(n6696), .Z(n6698) );
  AND U9710 ( .A(n6699), .B(n6698), .Z(n6700) );
  NAND U9711 ( .A(n6701), .B(n6700), .Z(n6702) );
  NANDN U9712 ( .A(n6703), .B(n6702), .Z(n6705) );
  NANDN U9713 ( .A(x[42]), .B(y[42]), .Z(n6704) );
  NAND U9714 ( .A(n6705), .B(n6704), .Z(n6711) );
  NANDN U9715 ( .A(n6707), .B(n6706), .Z(n6709) );
  ANDN U9716 ( .B(n6709), .A(n6708), .Z(n6710) );
  NAND U9717 ( .A(n6711), .B(n6710), .Z(n6712) );
  NANDN U9718 ( .A(n6713), .B(n6712), .Z(n10051) );
  NANDN U9719 ( .A(n10051), .B(n10050), .Z(n6715) );
  NAND U9720 ( .A(n6715), .B(n6714), .Z(n6717) );
  ANDN U9721 ( .B(n6717), .A(n6716), .Z(n6718) );
  NAND U9722 ( .A(n6718), .B(n10049), .Z(n6719) );
  NAND U9723 ( .A(n6719), .B(n10057), .Z(n6720) );
  NAND U9724 ( .A(n6720), .B(n10063), .Z(n6722) );
  NANDN U9725 ( .A(n6722), .B(n6721), .Z(n6723) );
  NANDN U9726 ( .A(n6724), .B(n6723), .Z(n6725) );
  NAND U9727 ( .A(n6725), .B(n10067), .Z(n6726) );
  NAND U9728 ( .A(n6726), .B(n10071), .Z(n6727) );
  NAND U9729 ( .A(n6727), .B(n10073), .Z(n6729) );
  ANDN U9730 ( .B(n6729), .A(n6728), .Z(n6730) );
  NANDN U9731 ( .A(n6730), .B(n10079), .Z(n6731) );
  NANDN U9732 ( .A(n6732), .B(n6731), .Z(n6733) );
  NAND U9733 ( .A(n6733), .B(n10083), .Z(n6734) );
  NANDN U9734 ( .A(n10085), .B(n6734), .Z(n6735) );
  NAND U9735 ( .A(n6735), .B(n10087), .Z(n6736) );
  ANDN U9736 ( .B(n6736), .A(n10090), .Z(n6737) );
  NANDN U9737 ( .A(n6737), .B(n10091), .Z(n6738) );
  AND U9738 ( .A(n10095), .B(n6738), .Z(n6739) );
  NANDN U9739 ( .A(n6739), .B(n10097), .Z(n6740) );
  NANDN U9740 ( .A(n6741), .B(n6740), .Z(n6742) );
  NANDN U9741 ( .A(n10104), .B(n6742), .Z(n6743) );
  NANDN U9742 ( .A(n6744), .B(n6743), .Z(n6745) );
  NANDN U9743 ( .A(n6746), .B(n6745), .Z(n6747) );
  NANDN U9744 ( .A(n6748), .B(n6747), .Z(n6749) );
  NANDN U9745 ( .A(n10118), .B(n6749), .Z(n6750) );
  NAND U9746 ( .A(n6750), .B(n10120), .Z(n6751) );
  ANDN U9747 ( .B(n6751), .A(n10122), .Z(n6752) );
  NANDN U9748 ( .A(n6752), .B(n10124), .Z(n6753) );
  NANDN U9749 ( .A(n10128), .B(n6753), .Z(n6754) );
  NANDN U9750 ( .A(n6755), .B(n6754), .Z(n6756) );
  NANDN U9751 ( .A(n10134), .B(n6756), .Z(n6757) );
  NAND U9752 ( .A(n6757), .B(n10136), .Z(n6758) );
  ANDN U9753 ( .B(n6758), .A(n10138), .Z(n6759) );
  NANDN U9754 ( .A(n6759), .B(n10048), .Z(n6760) );
  NAND U9755 ( .A(n6760), .B(n10141), .Z(n6761) );
  NANDN U9756 ( .A(n6762), .B(n6761), .Z(n6763) );
  NANDN U9757 ( .A(n10146), .B(n6763), .Z(n6764) );
  NAND U9758 ( .A(n6764), .B(n10148), .Z(n6765) );
  ANDN U9759 ( .B(n6765), .A(n10152), .Z(n6766) );
  OR U9760 ( .A(n6767), .B(n6766), .Z(n6768) );
  NANDN U9761 ( .A(n10158), .B(n6768), .Z(n6769) );
  NAND U9762 ( .A(n6769), .B(n10161), .Z(n6770) );
  NAND U9763 ( .A(n6770), .B(n10163), .Z(n6771) );
  NANDN U9764 ( .A(n6772), .B(n6771), .Z(n6773) );
  ANDN U9765 ( .B(n6773), .A(n10168), .Z(n6774) );
  NANDN U9766 ( .A(n6774), .B(n10169), .Z(n6775) );
  NANDN U9767 ( .A(n10172), .B(n6775), .Z(n6777) );
  NAND U9768 ( .A(n6777), .B(n6776), .Z(n6778) );
  NANDN U9769 ( .A(n6779), .B(n6778), .Z(n6781) );
  NAND U9770 ( .A(n6781), .B(n6780), .Z(n6783) );
  ANDN U9771 ( .B(n6783), .A(n6782), .Z(n6784) );
  NANDN U9772 ( .A(n6784), .B(n10190), .Z(n6785) );
  NANDN U9773 ( .A(n10193), .B(n6785), .Z(n6788) );
  ANDN U9774 ( .B(n6787), .A(n6786), .Z(n10194) );
  NAND U9775 ( .A(n6788), .B(n10194), .Z(n6789) );
  NANDN U9776 ( .A(n10196), .B(n6789), .Z(n6790) );
  NANDN U9777 ( .A(n10199), .B(n6790), .Z(n6791) );
  ANDN U9778 ( .B(n6791), .A(n10201), .Z(n6792) );
  NANDN U9779 ( .A(n6792), .B(n10204), .Z(n6793) );
  NAND U9780 ( .A(n6793), .B(n10206), .Z(n6794) );
  NANDN U9781 ( .A(n6795), .B(n6794), .Z(n6796) );
  NANDN U9782 ( .A(n10211), .B(n6796), .Z(n6797) );
  NAND U9783 ( .A(n6797), .B(n10212), .Z(n6798) );
  ANDN U9784 ( .B(n6798), .A(n10214), .Z(n6799) );
  NANDN U9785 ( .A(n6799), .B(n10217), .Z(n6800) );
  NAND U9786 ( .A(n6800), .B(n10221), .Z(n6801) );
  NANDN U9787 ( .A(n6802), .B(n6801), .Z(n6803) );
  NANDN U9788 ( .A(n10225), .B(n6803), .Z(n6804) );
  NANDN U9789 ( .A(n10227), .B(n6804), .Z(n6805) );
  NAND U9790 ( .A(n6805), .B(n10228), .Z(n6807) );
  ANDN U9791 ( .B(n6807), .A(n6806), .Z(n6808) );
  NAND U9792 ( .A(n6809), .B(n6808), .Z(n6810) );
  NAND U9793 ( .A(n6811), .B(n6810), .Z(n6812) );
  AND U9794 ( .A(n10235), .B(n6812), .Z(n6813) );
  ANDN U9795 ( .B(n6814), .A(n6813), .Z(n6815) );
  NAND U9796 ( .A(n6815), .B(n10239), .Z(n6817) );
  ANDN U9797 ( .B(n6817), .A(n6816), .Z(n6818) );
  OR U9798 ( .A(n10243), .B(n6818), .Z(n6819) );
  NANDN U9799 ( .A(n10244), .B(n6819), .Z(n6820) );
  NAND U9800 ( .A(n6820), .B(n10246), .Z(n6821) );
  NANDN U9801 ( .A(n10248), .B(n6821), .Z(n6822) );
  NAND U9802 ( .A(n6822), .B(n10252), .Z(n6824) );
  ANDN U9803 ( .B(n6824), .A(n6823), .Z(n6825) );
  NANDN U9804 ( .A(n6825), .B(n10258), .Z(n6826) );
  NANDN U9805 ( .A(n6827), .B(n6826), .Z(n6828) );
  NANDN U9806 ( .A(n10263), .B(n6828), .Z(n6829) );
  NANDN U9807 ( .A(n10265), .B(n6829), .Z(n6830) );
  AND U9808 ( .A(n6831), .B(n6830), .Z(n6832) );
  NAND U9809 ( .A(n6832), .B(n10266), .Z(n6833) );
  AND U9810 ( .A(n10268), .B(n6833), .Z(n6834) );
  NAND U9811 ( .A(n6834), .B(n10274), .Z(n6836) );
  NAND U9812 ( .A(n6836), .B(n6835), .Z(n6837) );
  NANDN U9813 ( .A(n6837), .B(n10276), .Z(n6838) );
  NANDN U9814 ( .A(n6839), .B(n6838), .Z(n6840) );
  NAND U9815 ( .A(n6840), .B(n10282), .Z(n6841) );
  NANDN U9816 ( .A(n6842), .B(n6841), .Z(n6843) );
  NAND U9817 ( .A(n6843), .B(n10285), .Z(n6844) );
  AND U9818 ( .A(n10045), .B(n6844), .Z(n6845) );
  OR U9819 ( .A(n10286), .B(n6845), .Z(n6846) );
  NANDN U9820 ( .A(n6847), .B(n6846), .Z(n6848) );
  NAND U9821 ( .A(n6848), .B(n10288), .Z(n6849) );
  NANDN U9822 ( .A(n10289), .B(n6849), .Z(n6850) );
  NAND U9823 ( .A(n6850), .B(n10290), .Z(n6851) );
  AND U9824 ( .A(n10292), .B(n6851), .Z(n6852) );
  NANDN U9825 ( .A(n6852), .B(n10293), .Z(n6853) );
  NANDN U9826 ( .A(n6854), .B(n6853), .Z(n6855) );
  NAND U9827 ( .A(n6855), .B(n10295), .Z(n6856) );
  NANDN U9828 ( .A(n10296), .B(n6856), .Z(n6857) );
  NAND U9829 ( .A(n6857), .B(n10297), .Z(n6858) );
  ANDN U9830 ( .B(n6858), .A(n10298), .Z(n6861) );
  AND U9831 ( .A(n10299), .B(n6859), .Z(n6860) );
  NANDN U9832 ( .A(n6861), .B(n6860), .Z(n6862) );
  ANDN U9833 ( .B(n6862), .A(n10300), .Z(n6864) );
  NANDN U9834 ( .A(n6864), .B(n6863), .Z(n6865) );
  NANDN U9835 ( .A(n10305), .B(n6865), .Z(n6866) );
  NANDN U9836 ( .A(n10307), .B(n6866), .Z(n6867) );
  NANDN U9837 ( .A(n6868), .B(n6867), .Z(n6869) );
  NANDN U9838 ( .A(n6869), .B(y[176]), .Z(n6872) );
  XNOR U9839 ( .A(n6869), .B(y[176]), .Z(n6870) );
  NANDN U9840 ( .A(x[176]), .B(n6870), .Z(n6871) );
  NAND U9841 ( .A(n6872), .B(n6871), .Z(n6873) );
  NAND U9842 ( .A(n6873), .B(n10314), .Z(n6874) );
  AND U9843 ( .A(n10316), .B(n6874), .Z(n6876) );
  NAND U9844 ( .A(n6876), .B(n6875), .Z(n6877) );
  NANDN U9845 ( .A(n6878), .B(n6877), .Z(n6879) );
  NAND U9846 ( .A(n6879), .B(n10322), .Z(n6881) );
  ANDN U9847 ( .B(n6881), .A(n6880), .Z(n6882) );
  NANDN U9848 ( .A(n6882), .B(n10326), .Z(n6883) );
  NAND U9849 ( .A(n6883), .B(n10328), .Z(n6884) );
  NANDN U9850 ( .A(n10331), .B(n6884), .Z(n6885) );
  NANDN U9851 ( .A(n10332), .B(n6885), .Z(n6886) );
  NAND U9852 ( .A(n6886), .B(n10336), .Z(n6888) );
  ANDN U9853 ( .B(n6888), .A(n6887), .Z(n6889) );
  NANDN U9854 ( .A(n6889), .B(n10340), .Z(n6890) );
  NAND U9855 ( .A(n6890), .B(n10344), .Z(n6891) );
  NAND U9856 ( .A(n6891), .B(n10346), .Z(n6892) );
  NANDN U9857 ( .A(n6893), .B(n6892), .Z(n6894) );
  NAND U9858 ( .A(n6894), .B(n10350), .Z(n6895) );
  AND U9859 ( .A(n10352), .B(n6895), .Z(n6896) );
  OR U9860 ( .A(n10355), .B(n6896), .Z(n6897) );
  NAND U9861 ( .A(n6897), .B(n10356), .Z(n6898) );
  NAND U9862 ( .A(n6898), .B(n10358), .Z(n6899) );
  NAND U9863 ( .A(n6899), .B(n10362), .Z(n6900) );
  NAND U9864 ( .A(n6900), .B(n10364), .Z(n6902) );
  ANDN U9865 ( .B(n6902), .A(n6901), .Z(n6903) );
  NANDN U9866 ( .A(n6903), .B(n10370), .Z(n6904) );
  NANDN U9867 ( .A(n6905), .B(n6904), .Z(n6906) );
  NANDN U9868 ( .A(n10377), .B(n6906), .Z(n6907) );
  NANDN U9869 ( .A(n6908), .B(n6907), .Z(n6909) );
  NAND U9870 ( .A(n6909), .B(n10382), .Z(n6910) );
  NAND U9871 ( .A(n6911), .B(n6910), .Z(n6912) );
  NANDN U9872 ( .A(n6912), .B(y[208]), .Z(n6915) );
  XNOR U9873 ( .A(n6912), .B(y[208]), .Z(n6913) );
  NANDN U9874 ( .A(x[208]), .B(n6913), .Z(n6914) );
  NAND U9875 ( .A(n6915), .B(n6914), .Z(n6916) );
  NAND U9876 ( .A(n6916), .B(n10043), .Z(n6917) );
  ANDN U9877 ( .B(n6917), .A(n10385), .Z(n6919) );
  NAND U9878 ( .A(n6919), .B(n6918), .Z(n6920) );
  NANDN U9879 ( .A(n6921), .B(n6920), .Z(n6922) );
  NAND U9880 ( .A(n6922), .B(n10387), .Z(n6923) );
  ANDN U9881 ( .B(n6923), .A(n10388), .Z(n6924) );
  NANDN U9882 ( .A(n6924), .B(n10389), .Z(n6925) );
  NANDN U9883 ( .A(n10390), .B(n6925), .Z(n6926) );
  NAND U9884 ( .A(n6926), .B(n10391), .Z(n6927) );
  NAND U9885 ( .A(n6927), .B(n10041), .Z(n6928) );
  NANDN U9886 ( .A(n10392), .B(n6928), .Z(n6930) );
  ANDN U9887 ( .B(n6930), .A(n6929), .Z(n6931) );
  OR U9888 ( .A(n10394), .B(n6931), .Z(n6932) );
  NAND U9889 ( .A(n6932), .B(n10395), .Z(n6933) );
  ANDN U9890 ( .B(n6933), .A(n10398), .Z(n6934) );
  OR U9891 ( .A(n10399), .B(n6934), .Z(n6935) );
  NANDN U9892 ( .A(n10402), .B(n6935), .Z(n6936) );
  NANDN U9893 ( .A(n10404), .B(n6936), .Z(n6937) );
  ANDN U9894 ( .B(n6937), .A(n10406), .Z(n6939) );
  NAND U9895 ( .A(n6939), .B(n6938), .Z(n6940) );
  NANDN U9896 ( .A(n10408), .B(n6940), .Z(n6941) );
  NANDN U9897 ( .A(n6942), .B(n6941), .Z(n6943) );
  NANDN U9898 ( .A(n10411), .B(n6943), .Z(n6944) );
  ANDN U9899 ( .B(n6944), .A(n10414), .Z(n6945) );
  NANDN U9900 ( .A(n6945), .B(n10415), .Z(n6946) );
  AND U9901 ( .A(n6947), .B(n6946), .Z(n6948) );
  NANDN U9902 ( .A(n6948), .B(n10419), .Z(n6949) );
  NANDN U9903 ( .A(n6950), .B(n6949), .Z(n6952) );
  NAND U9904 ( .A(n6952), .B(n6951), .Z(n6953) );
  AND U9905 ( .A(n6954), .B(n6953), .Z(n6956) );
  NAND U9906 ( .A(n6956), .B(n6955), .Z(n6957) );
  NANDN U9907 ( .A(n6958), .B(n6957), .Z(n6959) );
  NANDN U9908 ( .A(n6960), .B(n6959), .Z(n6961) );
  NANDN U9909 ( .A(n10428), .B(n6961), .Z(n6962) );
  ANDN U9910 ( .B(n6962), .A(n10430), .Z(n6963) );
  OR U9911 ( .A(n10432), .B(n6963), .Z(n6964) );
  NANDN U9912 ( .A(n6965), .B(n6964), .Z(n6967) );
  NAND U9913 ( .A(n6967), .B(n6966), .Z(n6968) );
  NANDN U9914 ( .A(n6969), .B(n6968), .Z(n6970) );
  NANDN U9915 ( .A(n6971), .B(n6970), .Z(n6972) );
  AND U9916 ( .A(n10449), .B(n6972), .Z(n6974) );
  NANDN U9917 ( .A(n6974), .B(n6973), .Z(n6975) );
  NAND U9918 ( .A(n6975), .B(n10455), .Z(n6976) );
  NANDN U9919 ( .A(n6977), .B(n6976), .Z(n6978) );
  NANDN U9920 ( .A(n10460), .B(n6978), .Z(n6979) );
  NANDN U9921 ( .A(n10462), .B(n6979), .Z(n6981) );
  ANDN U9922 ( .B(n6981), .A(n6980), .Z(n6982) );
  NANDN U9923 ( .A(n10464), .B(n6982), .Z(n6983) );
  NANDN U9924 ( .A(n6984), .B(n6983), .Z(n6986) );
  ANDN U9925 ( .B(n6986), .A(n6985), .Z(n6987) );
  NAND U9926 ( .A(n6987), .B(n10475), .Z(n6989) );
  NAND U9927 ( .A(n6989), .B(n6988), .Z(n6990) );
  AND U9928 ( .A(n6991), .B(n6990), .Z(n6992) );
  NAND U9929 ( .A(n6992), .B(n10474), .Z(n6993) );
  NAND U9930 ( .A(n6993), .B(n10478), .Z(n6994) );
  AND U9931 ( .A(n10485), .B(n6994), .Z(n6996) );
  NAND U9932 ( .A(n6996), .B(n6995), .Z(n6997) );
  AND U9933 ( .A(n6998), .B(n6997), .Z(n7000) );
  NAND U9934 ( .A(n7000), .B(n6999), .Z(n7002) );
  NANDN U9935 ( .A(y[280]), .B(n7002), .Z(n7001) );
  AND U9936 ( .A(n10492), .B(n7001), .Z(n7006) );
  XNOR U9937 ( .A(y[280]), .B(n7002), .Z(n7003) );
  NANDN U9938 ( .A(n7004), .B(n7003), .Z(n7005) );
  NAND U9939 ( .A(n7006), .B(n7005), .Z(n7007) );
  AND U9940 ( .A(n10495), .B(n7007), .Z(n7009) );
  NAND U9941 ( .A(n7009), .B(n7008), .Z(n7010) );
  NANDN U9942 ( .A(n7011), .B(n7010), .Z(n7012) );
  NANDN U9943 ( .A(n10499), .B(n7012), .Z(n7013) );
  NAND U9944 ( .A(n7013), .B(n10502), .Z(n7014) );
  AND U9945 ( .A(n10506), .B(n7014), .Z(n7015) );
  OR U9946 ( .A(n7016), .B(n7015), .Z(n7017) );
  NANDN U9947 ( .A(n10510), .B(n7017), .Z(n7018) );
  NAND U9948 ( .A(n7018), .B(n10511), .Z(n7019) );
  NANDN U9949 ( .A(n10514), .B(n7019), .Z(n7020) );
  NAND U9950 ( .A(n7020), .B(n10515), .Z(n7021) );
  ANDN U9951 ( .B(n7021), .A(n10517), .Z(n7022) );
  NANDN U9952 ( .A(n7022), .B(n10520), .Z(n7023) );
  NAND U9953 ( .A(n7023), .B(n10524), .Z(n7024) );
  NANDN U9954 ( .A(n7025), .B(n7024), .Z(n7026) );
  NANDN U9955 ( .A(n10528), .B(n7026), .Z(n7027) );
  NAND U9956 ( .A(n7027), .B(n10529), .Z(n7028) );
  AND U9957 ( .A(n10533), .B(n7028), .Z(n7030) );
  NANDN U9958 ( .A(n7030), .B(n7029), .Z(n7031) );
  NAND U9959 ( .A(n7031), .B(n10539), .Z(n7032) );
  NANDN U9960 ( .A(n7033), .B(n7032), .Z(n7034) );
  NANDN U9961 ( .A(n10544), .B(n7034), .Z(n7035) );
  NAND U9962 ( .A(n7035), .B(n10039), .Z(n7036) );
  AND U9963 ( .A(n10547), .B(n7036), .Z(n7037) );
  OR U9964 ( .A(n7038), .B(n7037), .Z(n7039) );
  NAND U9965 ( .A(n7039), .B(n10553), .Z(n7041) );
  NAND U9966 ( .A(n7041), .B(n7040), .Z(n7042) );
  NAND U9967 ( .A(n7042), .B(n10559), .Z(n7043) );
  NANDN U9968 ( .A(n7044), .B(n7043), .Z(n7045) );
  NANDN U9969 ( .A(n10564), .B(n7045), .Z(n7046) );
  NANDN U9970 ( .A(n10566), .B(n7046), .Z(n7047) );
  NAND U9971 ( .A(n7047), .B(n10567), .Z(n7048) );
  ANDN U9972 ( .B(n7048), .A(n10570), .Z(n7049) );
  NANDN U9973 ( .A(n7049), .B(n10571), .Z(n7050) );
  NANDN U9974 ( .A(n10573), .B(n7050), .Z(n7051) );
  NANDN U9975 ( .A(n10575), .B(n7051), .Z(n7052) );
  NAND U9976 ( .A(n7052), .B(n10578), .Z(n7053) );
  NAND U9977 ( .A(n7053), .B(n10579), .Z(n7054) );
  AND U9978 ( .A(n10037), .B(n7054), .Z(n7055) );
  NANDN U9979 ( .A(n7055), .B(n10583), .Z(n7056) );
  NANDN U9980 ( .A(n7057), .B(n7056), .Z(n7059) );
  NAND U9981 ( .A(n7059), .B(n7058), .Z(n7060) );
  NAND U9982 ( .A(n7060), .B(n10591), .Z(n7061) );
  AND U9983 ( .A(n10034), .B(n7061), .Z(n7062) );
  NAND U9984 ( .A(n7062), .B(n10594), .Z(n7063) );
  NANDN U9985 ( .A(n7064), .B(n7063), .Z(n7065) );
  AND U9986 ( .A(n7066), .B(n7065), .Z(n7067) );
  OR U9987 ( .A(n7068), .B(n7067), .Z(n7069) );
  AND U9988 ( .A(n7070), .B(n7069), .Z(n7071) );
  OR U9989 ( .A(n7072), .B(n7071), .Z(n7073) );
  NAND U9990 ( .A(n7073), .B(n10605), .Z(n7074) );
  NANDN U9991 ( .A(n7075), .B(n7074), .Z(n7076) );
  NANDN U9992 ( .A(n10607), .B(n7076), .Z(n7077) );
  NAND U9993 ( .A(n7077), .B(n10608), .Z(n7078) );
  AND U9994 ( .A(n10611), .B(n7078), .Z(n7079) );
  OR U9995 ( .A(n7080), .B(n7079), .Z(n7081) );
  NAND U9996 ( .A(n7081), .B(n10616), .Z(n7082) );
  AND U9997 ( .A(n10618), .B(n7082), .Z(n7083) );
  NANDN U9998 ( .A(n7083), .B(n10622), .Z(n7084) );
  NANDN U9999 ( .A(n7085), .B(n7084), .Z(n7086) );
  NANDN U10000 ( .A(n10626), .B(n7086), .Z(n7087) );
  NANDN U10001 ( .A(n10628), .B(n7087), .Z(n7088) );
  NANDN U10002 ( .A(n10632), .B(n7088), .Z(n7090) );
  ANDN U10003 ( .B(n7090), .A(n7089), .Z(n7091) );
  NANDN U10004 ( .A(n7091), .B(n10637), .Z(n7092) );
  NANDN U10005 ( .A(n10639), .B(n7092), .Z(n7093) );
  NAND U10006 ( .A(n7093), .B(n10641), .Z(n7095) );
  NANDN U10007 ( .A(n7095), .B(n7094), .Z(n7096) );
  NANDN U10008 ( .A(n10644), .B(n7096), .Z(n7098) );
  NAND U10009 ( .A(n7098), .B(n7097), .Z(n7099) );
  NANDN U10010 ( .A(n10648), .B(n7099), .Z(n7100) );
  NANDN U10011 ( .A(n10649), .B(n7100), .Z(n7101) );
  NAND U10012 ( .A(n7101), .B(n10651), .Z(n7102) );
  NANDN U10013 ( .A(n10032), .B(n7102), .Z(n7103) );
  NANDN U10014 ( .A(n7104), .B(n7103), .Z(n7105) );
  ANDN U10015 ( .B(n7105), .A(n10653), .Z(n7106) );
  NANDN U10016 ( .A(n7106), .B(n10655), .Z(n7107) );
  NAND U10017 ( .A(n7107), .B(n10656), .Z(n7108) );
  NANDN U10018 ( .A(n7109), .B(n7108), .Z(n7110) );
  NANDN U10019 ( .A(n10658), .B(n7110), .Z(n7111) );
  NANDN U10020 ( .A(n7112), .B(n7111), .Z(n7113) );
  ANDN U10021 ( .B(n7113), .A(n10661), .Z(n7114) );
  NANDN U10022 ( .A(n7114), .B(n10663), .Z(n7115) );
  NAND U10023 ( .A(n7115), .B(n10665), .Z(n7116) );
  NANDN U10024 ( .A(n7117), .B(n7116), .Z(n7118) );
  NANDN U10025 ( .A(n10670), .B(n7118), .Z(n7119) );
  NAND U10026 ( .A(n7119), .B(n10031), .Z(n7120) );
  AND U10027 ( .A(n10673), .B(n7120), .Z(n7121) );
  OR U10028 ( .A(n7122), .B(n7121), .Z(n7123) );
  NANDN U10029 ( .A(n10678), .B(n7123), .Z(n7124) );
  NAND U10030 ( .A(n7124), .B(n10680), .Z(n7125) );
  NAND U10031 ( .A(n7125), .B(n10683), .Z(n7127) );
  NAND U10032 ( .A(n7127), .B(n7126), .Z(n7128) );
  AND U10033 ( .A(n10689), .B(n7128), .Z(n7129) );
  OR U10034 ( .A(n7130), .B(n7129), .Z(n7131) );
  NANDN U10035 ( .A(n10694), .B(n7131), .Z(n7132) );
  NANDN U10036 ( .A(n10696), .B(n7132), .Z(n7133) );
  NANDN U10037 ( .A(n10697), .B(n7133), .Z(n7134) );
  NAND U10038 ( .A(n7134), .B(n10699), .Z(n7135) );
  ANDN U10039 ( .B(n7135), .A(n10702), .Z(n7136) );
  OR U10040 ( .A(n10704), .B(n7136), .Z(n7137) );
  NANDN U10041 ( .A(n10706), .B(n7137), .Z(n7138) );
  NANDN U10042 ( .A(n10708), .B(n7138), .Z(n7139) );
  NANDN U10043 ( .A(n10709), .B(n7139), .Z(n7140) );
  NAND U10044 ( .A(n7140), .B(n10712), .Z(n7141) );
  AND U10045 ( .A(n10716), .B(n7141), .Z(n7142) );
  OR U10046 ( .A(n7143), .B(n7142), .Z(n7144) );
  NANDN U10047 ( .A(n10720), .B(n7144), .Z(n7145) );
  NAND U10048 ( .A(n7145), .B(n10722), .Z(n7146) );
  NAND U10049 ( .A(n7146), .B(n10725), .Z(n7147) );
  NANDN U10050 ( .A(n7148), .B(n7147), .Z(n7149) );
  NAND U10051 ( .A(n7149), .B(n10731), .Z(n7150) );
  NANDN U10052 ( .A(n7151), .B(n7150), .Z(n7152) );
  NAND U10053 ( .A(n7152), .B(n10735), .Z(n7155) );
  NANDN U10054 ( .A(n7154), .B(n7153), .Z(n10738) );
  ANDN U10055 ( .B(n7155), .A(n10738), .Z(n7156) );
  OR U10056 ( .A(n10740), .B(n7156), .Z(n7157) );
  NAND U10057 ( .A(n7157), .B(n10741), .Z(n7158) );
  NAND U10058 ( .A(n7158), .B(n10743), .Z(n7159) );
  NANDN U10059 ( .A(n10744), .B(n7159), .Z(n7160) );
  NAND U10060 ( .A(n7160), .B(n10745), .Z(n7161) );
  ANDN U10061 ( .B(n7161), .A(n10746), .Z(n7162) );
  NANDN U10062 ( .A(n7162), .B(n10747), .Z(n7163) );
  NANDN U10063 ( .A(n10748), .B(n7163), .Z(n7164) );
  NAND U10064 ( .A(n7164), .B(n10749), .Z(n7165) );
  NANDN U10065 ( .A(n7166), .B(n7165), .Z(n7168) );
  NANDN U10066 ( .A(y[426]), .B(n7168), .Z(n7167) );
  AND U10067 ( .A(n10029), .B(n7167), .Z(n7171) );
  XNOR U10068 ( .A(y[426]), .B(n7168), .Z(n7169) );
  NAND U10069 ( .A(n7169), .B(x[426]), .Z(n7170) );
  NAND U10070 ( .A(n7171), .B(n7170), .Z(n7172) );
  AND U10071 ( .A(n10752), .B(n7172), .Z(n7173) );
  NANDN U10072 ( .A(n7174), .B(n7173), .Z(n7176) );
  NAND U10073 ( .A(n7176), .B(n7175), .Z(n7177) );
  AND U10074 ( .A(n7178), .B(n7177), .Z(n7179) );
  NAND U10075 ( .A(n7179), .B(n10025), .Z(n7180) );
  NAND U10076 ( .A(n7180), .B(n10027), .Z(n7182) );
  NANDN U10077 ( .A(n7182), .B(n7181), .Z(n7183) );
  AND U10078 ( .A(n10024), .B(n7183), .Z(n7184) );
  NAND U10079 ( .A(n7185), .B(n7184), .Z(n7186) );
  NAND U10080 ( .A(n7187), .B(n7186), .Z(n7188) );
  AND U10081 ( .A(n10763), .B(n7188), .Z(n7190) );
  NAND U10082 ( .A(n7190), .B(n7189), .Z(n7191) );
  NANDN U10083 ( .A(n7192), .B(n7191), .Z(n7193) );
  NAND U10084 ( .A(n7193), .B(n10769), .Z(n7194) );
  NANDN U10085 ( .A(n7195), .B(n7194), .Z(n7196) );
  ANDN U10086 ( .B(n7196), .A(n10774), .Z(n7197) );
  NANDN U10087 ( .A(n7197), .B(n10775), .Z(n7198) );
  NANDN U10088 ( .A(n10778), .B(n7198), .Z(n7199) );
  NAND U10089 ( .A(n7199), .B(n10780), .Z(n7200) );
  NANDN U10090 ( .A(n10784), .B(n7200), .Z(n7201) );
  NANDN U10091 ( .A(n7202), .B(n7201), .Z(n7203) );
  ANDN U10092 ( .B(n7203), .A(n10790), .Z(n7204) );
  OR U10093 ( .A(n10791), .B(n7204), .Z(n7205) );
  NANDN U10094 ( .A(n10794), .B(n7205), .Z(n7206) );
  NAND U10095 ( .A(n7206), .B(n10796), .Z(n7207) );
  NANDN U10096 ( .A(n10800), .B(n7207), .Z(n7208) );
  NANDN U10097 ( .A(n7209), .B(n7208), .Z(n7210) );
  ANDN U10098 ( .B(n7210), .A(n10806), .Z(n7211) );
  OR U10099 ( .A(n10807), .B(n7211), .Z(n7212) );
  AND U10100 ( .A(n7213), .B(n7212), .Z(n7214) );
  OR U10101 ( .A(n10812), .B(n7214), .Z(n7215) );
  NANDN U10102 ( .A(n7216), .B(n7215), .Z(n7217) );
  NAND U10103 ( .A(n7217), .B(n10815), .Z(n7218) );
  NANDN U10104 ( .A(n10818), .B(n7218), .Z(n7219) );
  NANDN U10105 ( .A(n10819), .B(n7219), .Z(n7220) );
  ANDN U10106 ( .B(n7220), .A(n10822), .Z(n7221) );
  OR U10107 ( .A(n10823), .B(n7221), .Z(n7222) );
  NANDN U10108 ( .A(n10826), .B(n7222), .Z(n7223) );
  NAND U10109 ( .A(n7223), .B(n10827), .Z(n7224) );
  NANDN U10110 ( .A(n7225), .B(n7224), .Z(n7226) );
  NANDN U10111 ( .A(n7227), .B(n7226), .Z(n7228) );
  ANDN U10112 ( .B(n7228), .A(n10840), .Z(n7229) );
  NANDN U10113 ( .A(n7229), .B(n10841), .Z(n7230) );
  NANDN U10114 ( .A(n10844), .B(n7230), .Z(n7231) );
  NAND U10115 ( .A(n7231), .B(n10847), .Z(n7232) );
  NAND U10116 ( .A(n7232), .B(n10849), .Z(n7233) );
  NANDN U10117 ( .A(n7234), .B(n7233), .Z(n7235) );
  ANDN U10118 ( .B(n7235), .A(n10853), .Z(n7236) );
  OR U10119 ( .A(n10856), .B(n7236), .Z(n7237) );
  ANDN U10120 ( .B(n7237), .A(n10858), .Z(n7238) );
  NANDN U10121 ( .A(n7238), .B(n10861), .Z(n7239) );
  NAND U10122 ( .A(n7239), .B(n10864), .Z(n7240) );
  NANDN U10123 ( .A(n7241), .B(n7240), .Z(n7242) );
  NANDN U10124 ( .A(n10869), .B(n7242), .Z(n7243) );
  NAND U10125 ( .A(n7243), .B(n10871), .Z(n7244) );
  ANDN U10126 ( .B(n7244), .A(n10874), .Z(n7245) );
  NANDN U10127 ( .A(n7245), .B(n10875), .Z(n7246) );
  NANDN U10128 ( .A(n10880), .B(n7246), .Z(n7247) );
  NANDN U10129 ( .A(n7248), .B(n7247), .Z(n7249) );
  NANDN U10130 ( .A(n10886), .B(n7249), .Z(n7250) );
  NAND U10131 ( .A(n7250), .B(n10887), .Z(n7251) );
  AND U10132 ( .A(n10889), .B(n7251), .Z(n7252) );
  NANDN U10133 ( .A(n7252), .B(n10891), .Z(n7253) );
  NANDN U10134 ( .A(n10893), .B(n7253), .Z(n7254) );
  NAND U10135 ( .A(n7254), .B(n10896), .Z(n7255) );
  NANDN U10136 ( .A(n10899), .B(n7255), .Z(n7256) );
  NANDN U10137 ( .A(n7257), .B(n7256), .Z(n7258) );
  NAND U10138 ( .A(n7258), .B(n10906), .Z(n7259) );
  NANDN U10139 ( .A(n7260), .B(n7259), .Z(n7261) );
  NAND U10140 ( .A(n7261), .B(n10909), .Z(n7262) );
  ANDN U10141 ( .B(n7262), .A(n10912), .Z(n7263) );
  NANDN U10142 ( .A(n7263), .B(n10913), .Z(n7265) );
  ANDN U10143 ( .B(n7265), .A(n7264), .Z(n7266) );
  OR U10144 ( .A(n7267), .B(n7266), .Z(n7268) );
  NANDN U10145 ( .A(n7269), .B(n7268), .Z(n7271) );
  NAND U10146 ( .A(n7271), .B(n7270), .Z(n7272) );
  NANDN U10147 ( .A(n10920), .B(n7272), .Z(n7273) );
  NANDN U10148 ( .A(n10921), .B(n7273), .Z(n7274) );
  NANDN U10149 ( .A(n10924), .B(n7274), .Z(n7275) );
  NANDN U10150 ( .A(n10926), .B(n7275), .Z(n7276) );
  NAND U10151 ( .A(n7276), .B(n10927), .Z(n7277) );
  ANDN U10152 ( .B(n7277), .A(n10932), .Z(n7278) );
  OR U10153 ( .A(n7279), .B(n7278), .Z(n7280) );
  NANDN U10154 ( .A(n10938), .B(n7280), .Z(n7281) );
  NAND U10155 ( .A(n7281), .B(n10939), .Z(n7282) );
  NANDN U10156 ( .A(n10942), .B(n7282), .Z(n7283) );
  NAND U10157 ( .A(n7283), .B(n10943), .Z(n7285) );
  ANDN U10158 ( .B(n7285), .A(n7284), .Z(n7287) );
  NANDN U10159 ( .A(n7287), .B(n7286), .Z(n7288) );
  AND U10160 ( .A(n7289), .B(n7288), .Z(n7290) );
  OR U10161 ( .A(n7291), .B(n7290), .Z(n7292) );
  NANDN U10162 ( .A(n7293), .B(n7292), .Z(n7295) );
  ANDN U10163 ( .B(n7295), .A(n7294), .Z(n7299) );
  AND U10164 ( .A(n7297), .B(n7296), .Z(n7298) );
  NANDN U10165 ( .A(n7299), .B(n7298), .Z(n7301) );
  ANDN U10166 ( .B(n7301), .A(n7300), .Z(n7303) );
  NANDN U10167 ( .A(n7303), .B(n7302), .Z(n7304) );
  NAND U10168 ( .A(n7304), .B(n10954), .Z(n7305) );
  ANDN U10169 ( .B(n7305), .A(n10955), .Z(n7306) );
  NANDN U10170 ( .A(n7306), .B(n10023), .Z(n7307) );
  NANDN U10171 ( .A(n10020), .B(n7307), .Z(n7308) );
  NANDN U10172 ( .A(n7309), .B(n7308), .Z(n7310) );
  NANDN U10173 ( .A(n10957), .B(n7310), .Z(n7311) );
  NAND U10174 ( .A(n7311), .B(n10959), .Z(n7312) );
  AND U10175 ( .A(n10960), .B(n7312), .Z(n7313) );
  OR U10176 ( .A(n7314), .B(n7313), .Z(n7315) );
  NAND U10177 ( .A(n7315), .B(n10962), .Z(n7316) );
  ANDN U10178 ( .B(n7316), .A(n10963), .Z(n7317) );
  NANDN U10179 ( .A(n7317), .B(n10964), .Z(n7318) );
  NANDN U10180 ( .A(n10965), .B(n7318), .Z(n7319) );
  NAND U10181 ( .A(n7319), .B(n10966), .Z(n7321) );
  NANDN U10182 ( .A(n7321), .B(n7320), .Z(n7322) );
  NAND U10183 ( .A(n7322), .B(n10967), .Z(n7324) );
  NAND U10184 ( .A(n7324), .B(n7323), .Z(n7325) );
  NANDN U10185 ( .A(n7326), .B(n7325), .Z(n7328) );
  NANDN U10186 ( .A(y[570]), .B(n7328), .Z(n7327) );
  AND U10187 ( .A(n10976), .B(n7327), .Z(n7331) );
  XNOR U10188 ( .A(y[570]), .B(n7328), .Z(n7329) );
  NAND U10189 ( .A(n7329), .B(x[570]), .Z(n7330) );
  NAND U10190 ( .A(n7331), .B(n7330), .Z(n7332) );
  AND U10191 ( .A(n10980), .B(n7332), .Z(n7333) );
  NANDN U10192 ( .A(n7334), .B(n7333), .Z(n7335) );
  NANDN U10193 ( .A(n7336), .B(n7335), .Z(n7337) );
  NANDN U10194 ( .A(n10983), .B(n7337), .Z(n7338) );
  NAND U10195 ( .A(n7338), .B(n10985), .Z(n7339) );
  ANDN U10196 ( .B(n7339), .A(n10988), .Z(n7340) );
  NANDN U10197 ( .A(n7340), .B(n10989), .Z(n7341) );
  NAND U10198 ( .A(n7341), .B(n10993), .Z(n7343) );
  ANDN U10199 ( .B(n7343), .A(n7342), .Z(n7344) );
  NANDN U10200 ( .A(n7344), .B(n10999), .Z(n7346) );
  NAND U10201 ( .A(n7346), .B(n7345), .Z(n7347) );
  NANDN U10202 ( .A(n10018), .B(n7347), .Z(n7348) );
  NANDN U10203 ( .A(n7349), .B(n7348), .Z(n7350) );
  NAND U10204 ( .A(n7350), .B(n11010), .Z(n7351) );
  ANDN U10205 ( .B(n7351), .A(n11012), .Z(n7353) );
  NANDN U10206 ( .A(n7353), .B(n7352), .Z(n7354) );
  ANDN U10207 ( .B(n7354), .A(n11016), .Z(n7356) );
  NANDN U10208 ( .A(n7356), .B(n7355), .Z(n7357) );
  NAND U10209 ( .A(n7358), .B(n7357), .Z(n7359) );
  NANDN U10210 ( .A(n7359), .B(y[594]), .Z(n7362) );
  XNOR U10211 ( .A(n7359), .B(y[594]), .Z(n7360) );
  NANDN U10212 ( .A(x[594]), .B(n7360), .Z(n7361) );
  NAND U10213 ( .A(n7362), .B(n7361), .Z(n7363) );
  NAND U10214 ( .A(n7364), .B(n7363), .Z(n7365) );
  NAND U10215 ( .A(n7366), .B(n7365), .Z(n7367) );
  NANDN U10216 ( .A(n7368), .B(n7367), .Z(n7370) );
  NAND U10217 ( .A(n7370), .B(n7369), .Z(n7371) );
  ANDN U10218 ( .B(n7371), .A(n11036), .Z(n7372) );
  NANDN U10219 ( .A(n7372), .B(n11037), .Z(n7373) );
  ANDN U10220 ( .B(n7373), .A(n11040), .Z(n7374) );
  NANDN U10221 ( .A(n7374), .B(n11041), .Z(n7375) );
  NANDN U10222 ( .A(n11044), .B(n7375), .Z(n7377) );
  NAND U10223 ( .A(n7377), .B(n7376), .Z(n7378) );
  NANDN U10224 ( .A(n7378), .B(n11046), .Z(n7379) );
  NANDN U10225 ( .A(n11048), .B(n7379), .Z(n7380) );
  NAND U10226 ( .A(n7380), .B(n11053), .Z(n7382) );
  NANDN U10227 ( .A(n7382), .B(n7381), .Z(n7383) );
  NANDN U10228 ( .A(n7384), .B(n7383), .Z(n7385) );
  NAND U10229 ( .A(n7385), .B(n11058), .Z(n7387) );
  NANDN U10230 ( .A(n7387), .B(n7386), .Z(n7388) );
  NANDN U10231 ( .A(n11060), .B(n7388), .Z(n7390) );
  NAND U10232 ( .A(n7390), .B(n7389), .Z(n7391) );
  NANDN U10233 ( .A(n11064), .B(n7391), .Z(n7392) );
  NAND U10234 ( .A(n7392), .B(n11065), .Z(n7393) );
  ANDN U10235 ( .B(n7393), .A(n11068), .Z(n7394) );
  OR U10236 ( .A(n11069), .B(n7394), .Z(n7395) );
  NAND U10237 ( .A(n7395), .B(n11071), .Z(n7396) );
  ANDN U10238 ( .B(n7396), .A(n11074), .Z(n7397) );
  NANDN U10239 ( .A(n7397), .B(n11075), .Z(n7398) );
  NANDN U10240 ( .A(n11080), .B(n7398), .Z(n7399) );
  NANDN U10241 ( .A(n7400), .B(n7399), .Z(n7401) );
  NANDN U10242 ( .A(n11083), .B(n7401), .Z(n7402) );
  NAND U10243 ( .A(n7402), .B(n11084), .Z(n7403) );
  ANDN U10244 ( .B(n7403), .A(n11085), .Z(n7404) );
  OR U10245 ( .A(n11086), .B(n7404), .Z(n7405) );
  NANDN U10246 ( .A(n11087), .B(n7405), .Z(n7406) );
  NANDN U10247 ( .A(n7407), .B(n7406), .Z(n7408) );
  NANDN U10248 ( .A(n7408), .B(y[642]), .Z(n7411) );
  XNOR U10249 ( .A(n7408), .B(y[642]), .Z(n7409) );
  NANDN U10250 ( .A(x[642]), .B(n7409), .Z(n7410) );
  NAND U10251 ( .A(n7411), .B(n7410), .Z(n7412) );
  NAND U10252 ( .A(n7412), .B(n11091), .Z(n7413) );
  AND U10253 ( .A(n11092), .B(n7413), .Z(n7415) );
  NAND U10254 ( .A(n7415), .B(n7414), .Z(n7416) );
  NANDN U10255 ( .A(n7417), .B(n7416), .Z(n7418) );
  NANDN U10256 ( .A(n11094), .B(n7418), .Z(n7419) );
  NAND U10257 ( .A(n7419), .B(n10017), .Z(n7420) );
  NANDN U10258 ( .A(n11095), .B(n7420), .Z(n7421) );
  NANDN U10259 ( .A(n7422), .B(n7421), .Z(n7423) );
  AND U10260 ( .A(n11099), .B(n7423), .Z(n7424) );
  OR U10261 ( .A(n7425), .B(n7424), .Z(n7426) );
  NANDN U10262 ( .A(n11101), .B(n7426), .Z(n7427) );
  NAND U10263 ( .A(n7427), .B(n11102), .Z(n7428) );
  NANDN U10264 ( .A(n11103), .B(n7428), .Z(n7429) );
  NAND U10265 ( .A(n7429), .B(n11105), .Z(n7430) );
  AND U10266 ( .A(n11106), .B(n7430), .Z(n7431) );
  OR U10267 ( .A(n7432), .B(n7431), .Z(n7433) );
  NAND U10268 ( .A(n7433), .B(n11109), .Z(n7435) );
  ANDN U10269 ( .B(n7435), .A(n7434), .Z(n7436) );
  NANDN U10270 ( .A(n7436), .B(n11111), .Z(n7437) );
  ANDN U10271 ( .B(n7437), .A(n11112), .Z(n7438) );
  NANDN U10272 ( .A(n7438), .B(n11114), .Z(n7440) );
  NAND U10273 ( .A(n7440), .B(n7439), .Z(n7441) );
  NAND U10274 ( .A(n7441), .B(n11116), .Z(n7442) );
  NAND U10275 ( .A(n7443), .B(n7442), .Z(n7444) );
  AND U10276 ( .A(n7445), .B(n7444), .Z(n7448) );
  AND U10277 ( .A(n11120), .B(n7446), .Z(n7447) );
  NANDN U10278 ( .A(n7448), .B(n7447), .Z(n7449) );
  AND U10279 ( .A(n7450), .B(n7449), .Z(n7451) );
  NAND U10280 ( .A(n7451), .B(n11122), .Z(n7452) );
  AND U10281 ( .A(n7453), .B(n7452), .Z(n7454) );
  AND U10282 ( .A(n7455), .B(n7454), .Z(n7456) );
  OR U10283 ( .A(n7456), .B(y[674]), .Z(n7459) );
  XOR U10284 ( .A(y[674]), .B(n7456), .Z(n7457) );
  NAND U10285 ( .A(n7457), .B(x[674]), .Z(n7458) );
  NAND U10286 ( .A(n7459), .B(n7458), .Z(n7460) );
  AND U10287 ( .A(n7461), .B(n7460), .Z(n7462) );
  NANDN U10288 ( .A(n7462), .B(n11125), .Z(n7463) );
  NANDN U10289 ( .A(n11126), .B(n7463), .Z(n7464) );
  NAND U10290 ( .A(n7464), .B(n11128), .Z(n7465) );
  NANDN U10291 ( .A(n11129), .B(n7465), .Z(n7466) );
  NANDN U10292 ( .A(n7467), .B(n7466), .Z(n7469) );
  NAND U10293 ( .A(n7469), .B(n7468), .Z(n7470) );
  NANDN U10294 ( .A(n7471), .B(n7470), .Z(n7472) );
  NAND U10295 ( .A(n7472), .B(n11135), .Z(n7473) );
  AND U10296 ( .A(n11136), .B(n7473), .Z(n7476) );
  ANDN U10297 ( .B(n7475), .A(n7474), .Z(n11138) );
  NOR U10298 ( .A(n7476), .B(n11138), .Z(n7478) );
  NAND U10299 ( .A(n7478), .B(n7477), .Z(n7479) );
  NAND U10300 ( .A(n7479), .B(n11139), .Z(n7481) );
  ANDN U10301 ( .B(n7481), .A(n7480), .Z(n7482) );
  NANDN U10302 ( .A(n7483), .B(n7482), .Z(n7484) );
  NAND U10303 ( .A(n7484), .B(n11141), .Z(n7485) );
  ANDN U10304 ( .B(n7485), .A(n11142), .Z(n7486) );
  NANDN U10305 ( .A(n7486), .B(n11143), .Z(n7487) );
  NANDN U10306 ( .A(n11144), .B(n7487), .Z(n7488) );
  NAND U10307 ( .A(n7488), .B(n11146), .Z(n7489) );
  NAND U10308 ( .A(n7489), .B(n11147), .Z(n7491) );
  NAND U10309 ( .A(n7491), .B(n7490), .Z(n7493) );
  ANDN U10310 ( .B(n7493), .A(n7492), .Z(n7494) );
  OR U10311 ( .A(n7495), .B(n7494), .Z(n7496) );
  NANDN U10312 ( .A(n11152), .B(n7496), .Z(n7497) );
  NAND U10313 ( .A(n7497), .B(n11153), .Z(n7498) );
  NANDN U10314 ( .A(n11156), .B(n7498), .Z(n7499) );
  NAND U10315 ( .A(n7499), .B(n11159), .Z(n7500) );
  AND U10316 ( .A(n11161), .B(n7500), .Z(n7501) );
  OR U10317 ( .A(n7502), .B(n7501), .Z(n7503) );
  NAND U10318 ( .A(n7503), .B(n11167), .Z(n7504) );
  NANDN U10319 ( .A(n7505), .B(n7504), .Z(n7506) );
  NAND U10320 ( .A(n7506), .B(n11173), .Z(n7507) );
  NAND U10321 ( .A(n7508), .B(n7507), .Z(n7509) );
  NANDN U10322 ( .A(n7509), .B(n11177), .Z(n7510) );
  NANDN U10323 ( .A(n11180), .B(n7510), .Z(n7511) );
  NAND U10324 ( .A(n7511), .B(n11182), .Z(n7512) );
  NANDN U10325 ( .A(n11184), .B(n7512), .Z(n7513) );
  NAND U10326 ( .A(n7513), .B(n11185), .Z(n7514) );
  ANDN U10327 ( .B(n7514), .A(n11188), .Z(n7515) );
  NANDN U10328 ( .A(n7515), .B(n11190), .Z(n7516) );
  AND U10329 ( .A(n11193), .B(n7516), .Z(n7518) );
  NANDN U10330 ( .A(n7518), .B(n7517), .Z(n7519) );
  NAND U10331 ( .A(n7519), .B(n11200), .Z(n7520) );
  NANDN U10332 ( .A(n7521), .B(n7520), .Z(n7522) );
  NANDN U10333 ( .A(n11204), .B(n7522), .Z(n7523) );
  NAND U10334 ( .A(n7523), .B(n11205), .Z(n7524) );
  ANDN U10335 ( .B(n7524), .A(n11210), .Z(n7525) );
  OR U10336 ( .A(n7526), .B(n7525), .Z(n7527) );
  ANDN U10337 ( .B(n7527), .A(n11216), .Z(n7528) );
  OR U10338 ( .A(n11218), .B(n7528), .Z(n7529) );
  NAND U10339 ( .A(n7529), .B(n11219), .Z(n7530) );
  AND U10340 ( .A(n11222), .B(n7530), .Z(n7531) );
  NANDN U10341 ( .A(n7531), .B(n11225), .Z(n7532) );
  NANDN U10342 ( .A(n7533), .B(n7532), .Z(n7534) );
  NAND U10343 ( .A(n7534), .B(n11230), .Z(n7535) );
  NANDN U10344 ( .A(n11231), .B(n7535), .Z(n7536) );
  NAND U10345 ( .A(n7536), .B(n11236), .Z(n7537) );
  AND U10346 ( .A(n7538), .B(n7537), .Z(n7539) );
  NANDN U10347 ( .A(n7539), .B(n11238), .Z(n7540) );
  NANDN U10348 ( .A(n11242), .B(n7540), .Z(n7541) );
  NAND U10349 ( .A(n7541), .B(n11243), .Z(n7543) );
  NANDN U10350 ( .A(n7543), .B(n7542), .Z(n7544) );
  NANDN U10351 ( .A(n11245), .B(n7544), .Z(n7546) );
  NAND U10352 ( .A(n7546), .B(n7545), .Z(n7547) );
  NANDN U10353 ( .A(n7548), .B(n7547), .Z(n7550) );
  NAND U10354 ( .A(n7550), .B(n7549), .Z(n7552) );
  ANDN U10355 ( .B(n7552), .A(n7551), .Z(n7555) );
  AND U10356 ( .A(n11259), .B(n7553), .Z(n7554) );
  NANDN U10357 ( .A(n7555), .B(n7554), .Z(n7556) );
  ANDN U10358 ( .B(n7556), .A(n11262), .Z(n7558) );
  NANDN U10359 ( .A(n7558), .B(n7557), .Z(n7559) );
  NANDN U10360 ( .A(n11266), .B(n7559), .Z(n7564) );
  NANDN U10361 ( .A(x[752]), .B(y[752]), .Z(n7560) );
  AND U10362 ( .A(n7561), .B(n7560), .Z(n7562) );
  OR U10363 ( .A(n7563), .B(n7562), .Z(n11268) );
  NAND U10364 ( .A(n7564), .B(n11268), .Z(n7566) );
  NANDN U10365 ( .A(n7566), .B(n7565), .Z(n7567) );
  NANDN U10366 ( .A(n11270), .B(n7567), .Z(n7569) );
  NAND U10367 ( .A(n7569), .B(n7568), .Z(n7570) );
  NANDN U10368 ( .A(n11276), .B(n7570), .Z(n7571) );
  NAND U10369 ( .A(n7571), .B(n11278), .Z(n7573) );
  ANDN U10370 ( .B(n7573), .A(n7572), .Z(n7574) );
  NANDN U10371 ( .A(n7574), .B(n11283), .Z(n7575) );
  NANDN U10372 ( .A(n11286), .B(n7575), .Z(n7576) );
  NAND U10373 ( .A(n7576), .B(n11287), .Z(n7577) );
  NANDN U10374 ( .A(n11290), .B(n7577), .Z(n7578) );
  NAND U10375 ( .A(n7578), .B(n11292), .Z(n7579) );
  ANDN U10376 ( .B(n7579), .A(n11294), .Z(n7580) );
  OR U10377 ( .A(n11296), .B(n7580), .Z(n7581) );
  NAND U10378 ( .A(n7581), .B(n11297), .Z(n7582) );
  AND U10379 ( .A(n11301), .B(n7582), .Z(n7584) );
  NANDN U10380 ( .A(n7584), .B(n7583), .Z(n7585) );
  AND U10381 ( .A(n11307), .B(n7585), .Z(n7586) );
  OR U10382 ( .A(n7587), .B(n7586), .Z(n7588) );
  NANDN U10383 ( .A(n11312), .B(n7588), .Z(n7589) );
  ANDN U10384 ( .B(n7589), .A(n11313), .Z(n7590) );
  NANDN U10385 ( .A(n7590), .B(n11317), .Z(n7592) );
  NAND U10386 ( .A(n7592), .B(n7591), .Z(n7593) );
  NAND U10387 ( .A(n7593), .B(n11323), .Z(n7594) );
  NANDN U10388 ( .A(n7595), .B(n7594), .Z(n7596) );
  NANDN U10389 ( .A(n11328), .B(n7596), .Z(n7597) );
  NAND U10390 ( .A(n7597), .B(n11329), .Z(n7598) );
  NANDN U10391 ( .A(n11331), .B(n7598), .Z(n7599) );
  NAND U10392 ( .A(n7599), .B(n11333), .Z(n7600) );
  ANDN U10393 ( .B(n7600), .A(n11336), .Z(n7601) );
  NANDN U10394 ( .A(n7601), .B(n11337), .Z(n7602) );
  AND U10395 ( .A(n11339), .B(n7602), .Z(n7603) );
  NANDN U10396 ( .A(n7603), .B(n11341), .Z(n7604) );
  NANDN U10397 ( .A(n11343), .B(n7604), .Z(n7605) );
  NAND U10398 ( .A(n7605), .B(n11346), .Z(n7606) );
  NAND U10399 ( .A(n7606), .B(n11350), .Z(n7607) );
  AND U10400 ( .A(n7608), .B(n7607), .Z(n7610) );
  NAND U10401 ( .A(n7610), .B(n7609), .Z(n7612) );
  NANDN U10402 ( .A(y[794]), .B(n7612), .Z(n7611) );
  AND U10403 ( .A(n11357), .B(n7611), .Z(n7616) );
  XNOR U10404 ( .A(y[794]), .B(n7612), .Z(n7613) );
  NANDN U10405 ( .A(n7614), .B(n7613), .Z(n7615) );
  NAND U10406 ( .A(n7616), .B(n7615), .Z(n7617) );
  NANDN U10407 ( .A(n7618), .B(n7617), .Z(n7619) );
  NANDN U10408 ( .A(n7619), .B(n11359), .Z(n7620) );
  NANDN U10409 ( .A(n7621), .B(n7620), .Z(n7622) );
  NANDN U10410 ( .A(n11366), .B(n7622), .Z(n7626) );
  NAND U10411 ( .A(n11363), .B(n11369), .Z(n7624) );
  NAND U10412 ( .A(n7624), .B(n7623), .Z(n7625) );
  AND U10413 ( .A(n7626), .B(n7625), .Z(n7627) );
  NANDN U10414 ( .A(n7627), .B(n11371), .Z(n7628) );
  NANDN U10415 ( .A(n7629), .B(n7628), .Z(n7630) );
  NAND U10416 ( .A(n7630), .B(n11375), .Z(n7631) );
  NANDN U10417 ( .A(n11378), .B(n7631), .Z(n7632) );
  NAND U10418 ( .A(n7632), .B(n11379), .Z(n7633) );
  ANDN U10419 ( .B(n7633), .A(n11382), .Z(n7634) );
  NANDN U10420 ( .A(n7634), .B(n11383), .Z(n7635) );
  NANDN U10421 ( .A(n11384), .B(n7635), .Z(n7636) );
  NAND U10422 ( .A(n7636), .B(n11385), .Z(n7637) );
  NANDN U10423 ( .A(n11386), .B(n7637), .Z(n7638) );
  NANDN U10424 ( .A(n11387), .B(n7638), .Z(n7639) );
  AND U10425 ( .A(n11389), .B(n7639), .Z(n7640) );
  OR U10426 ( .A(n7640), .B(n10009), .Z(n7641) );
  NANDN U10427 ( .A(n7642), .B(n7641), .Z(n7643) );
  NAND U10428 ( .A(n7643), .B(n11391), .Z(n7644) );
  NANDN U10429 ( .A(n11392), .B(n7644), .Z(n7645) );
  AND U10430 ( .A(n7646), .B(n7645), .Z(n7647) );
  NAND U10431 ( .A(n7647), .B(n11393), .Z(n7648) );
  AND U10432 ( .A(n11394), .B(n7648), .Z(n7649) );
  NAND U10433 ( .A(n7649), .B(n11397), .Z(n7651) );
  NAND U10434 ( .A(n7651), .B(n7650), .Z(n7652) );
  NANDN U10435 ( .A(n7652), .B(n11398), .Z(n7653) );
  NANDN U10436 ( .A(n7654), .B(n7653), .Z(n7655) );
  NAND U10437 ( .A(n7655), .B(n11401), .Z(n7656) );
  NAND U10438 ( .A(n7656), .B(n11403), .Z(n7657) );
  NANDN U10439 ( .A(n11406), .B(n7657), .Z(n7658) );
  ANDN U10440 ( .B(n7658), .A(n11408), .Z(n7665) );
  OR U10441 ( .A(n7660), .B(n7659), .Z(n7662) );
  ANDN U10442 ( .B(n7662), .A(n7661), .Z(n7664) );
  ANDN U10443 ( .B(n7664), .A(n7663), .Z(n11410) );
  NANDN U10444 ( .A(n7665), .B(n11410), .Z(n7670) );
  NANDN U10445 ( .A(y[828]), .B(x[828]), .Z(n7666) );
  AND U10446 ( .A(n7667), .B(n7666), .Z(n7668) );
  NOR U10447 ( .A(n7669), .B(n7668), .Z(n11412) );
  ANDN U10448 ( .B(n7670), .A(n11412), .Z(n7672) );
  NAND U10449 ( .A(n7672), .B(n7671), .Z(n7673) );
  NAND U10450 ( .A(n7673), .B(n11413), .Z(n7675) );
  ANDN U10451 ( .B(n7675), .A(n7674), .Z(n7677) );
  NAND U10452 ( .A(n7677), .B(n7676), .Z(n7678) );
  NAND U10453 ( .A(n7678), .B(n11417), .Z(n7679) );
  AND U10454 ( .A(n7680), .B(n7679), .Z(n7681) );
  NAND U10455 ( .A(n7682), .B(n7681), .Z(n7683) );
  NAND U10456 ( .A(n7684), .B(n7683), .Z(n7686) );
  AND U10457 ( .A(n7686), .B(n7685), .Z(n7687) );
  OR U10458 ( .A(n7687), .B(y[836]), .Z(n7690) );
  XOR U10459 ( .A(y[836]), .B(n7687), .Z(n7688) );
  NAND U10460 ( .A(n7688), .B(x[836]), .Z(n7689) );
  NAND U10461 ( .A(n7690), .B(n7689), .Z(n7692) );
  ANDN U10462 ( .B(n7692), .A(n7691), .Z(n7693) );
  NANDN U10463 ( .A(n7693), .B(n11427), .Z(n7694) );
  NANDN U10464 ( .A(n11430), .B(n7694), .Z(n7695) );
  NAND U10465 ( .A(n7695), .B(n11432), .Z(n7696) );
  NAND U10466 ( .A(n7696), .B(n11433), .Z(n7697) );
  NAND U10467 ( .A(n7697), .B(n11438), .Z(n7699) );
  ANDN U10468 ( .B(n7699), .A(n7698), .Z(n7700) );
  NANDN U10469 ( .A(n7700), .B(n11441), .Z(n7701) );
  NANDN U10470 ( .A(n11444), .B(n7701), .Z(n7702) );
  NAND U10471 ( .A(n7702), .B(n11445), .Z(n7703) );
  NANDN U10472 ( .A(n11448), .B(n7703), .Z(n7704) );
  NAND U10473 ( .A(n7704), .B(n11450), .Z(n7706) );
  ANDN U10474 ( .B(n7706), .A(n7705), .Z(n7708) );
  NANDN U10475 ( .A(n7708), .B(n7707), .Z(n7710) );
  ANDN U10476 ( .B(n7710), .A(n7709), .Z(n7711) );
  NAND U10477 ( .A(n7712), .B(n7711), .Z(n7713) );
  NAND U10478 ( .A(n7714), .B(n7713), .Z(n7716) );
  ANDN U10479 ( .B(n7716), .A(n7715), .Z(n7717) );
  NAND U10480 ( .A(n7717), .B(n11459), .Z(n7718) );
  NAND U10481 ( .A(n7718), .B(n11462), .Z(n7719) );
  NANDN U10482 ( .A(n11464), .B(n7719), .Z(n7720) );
  NAND U10483 ( .A(n7720), .B(n11465), .Z(n7721) );
  ANDN U10484 ( .B(n7721), .A(n11468), .Z(n7722) );
  NANDN U10485 ( .A(n7722), .B(n11469), .Z(n7723) );
  NAND U10486 ( .A(n7723), .B(n11472), .Z(n7724) );
  NAND U10487 ( .A(n7724), .B(n11475), .Z(n7725) );
  NANDN U10488 ( .A(n7726), .B(n7725), .Z(n7727) );
  AND U10489 ( .A(n7728), .B(n7727), .Z(n7729) );
  NAND U10490 ( .A(n7729), .B(n11480), .Z(n7730) );
  AND U10491 ( .A(n11481), .B(n7730), .Z(n7731) );
  NAND U10492 ( .A(n7732), .B(n7731), .Z(n7733) );
  NAND U10493 ( .A(n7734), .B(n7733), .Z(n7736) );
  ANDN U10494 ( .B(n7736), .A(n7735), .Z(n7737) );
  NAND U10495 ( .A(n7737), .B(n11489), .Z(n7738) );
  NAND U10496 ( .A(n7738), .B(n11492), .Z(n7739) );
  NANDN U10497 ( .A(n11494), .B(n7739), .Z(n7740) );
  NAND U10498 ( .A(n7740), .B(n11495), .Z(n7741) );
  ANDN U10499 ( .B(n7741), .A(n11498), .Z(n7742) );
  NANDN U10500 ( .A(n7742), .B(n11499), .Z(n7743) );
  NAND U10501 ( .A(n7743), .B(n11502), .Z(n7744) );
  NAND U10502 ( .A(n7744), .B(n11505), .Z(n7745) );
  NANDN U10503 ( .A(n7746), .B(n7745), .Z(n7747) );
  AND U10504 ( .A(n7748), .B(n7747), .Z(n7749) );
  NAND U10505 ( .A(n7749), .B(n11510), .Z(n7750) );
  AND U10506 ( .A(n11511), .B(n7750), .Z(n7751) );
  NAND U10507 ( .A(n7752), .B(n7751), .Z(n7753) );
  NAND U10508 ( .A(n7754), .B(n7753), .Z(n7756) );
  ANDN U10509 ( .B(n7756), .A(n7755), .Z(n7757) );
  NAND U10510 ( .A(n7757), .B(n11519), .Z(n7758) );
  NAND U10511 ( .A(n7758), .B(n11522), .Z(n7759) );
  NANDN U10512 ( .A(n11524), .B(n7759), .Z(n7760) );
  NAND U10513 ( .A(n7760), .B(n11525), .Z(n7761) );
  ANDN U10514 ( .B(n7761), .A(n11528), .Z(n7762) );
  NANDN U10515 ( .A(n7762), .B(n11529), .Z(n7763) );
  NAND U10516 ( .A(n7763), .B(n11532), .Z(n7764) );
  NANDN U10517 ( .A(n11536), .B(n7764), .Z(n7765) );
  NANDN U10518 ( .A(n7766), .B(n7765), .Z(n7767) );
  NAND U10519 ( .A(n7767), .B(n11543), .Z(n7768) );
  ANDN U10520 ( .B(n7768), .A(n11546), .Z(n7769) );
  NANDN U10521 ( .A(n7769), .B(n11547), .Z(n7770) );
  NAND U10522 ( .A(n7770), .B(n11549), .Z(n7771) );
  NAND U10523 ( .A(n7771), .B(n11552), .Z(n7772) );
  NANDN U10524 ( .A(n11554), .B(n7772), .Z(n7773) );
  NAND U10525 ( .A(n7773), .B(n11555), .Z(n7774) );
  ANDN U10526 ( .B(n7774), .A(n11558), .Z(n7775) );
  NANDN U10527 ( .A(n7775), .B(n11559), .Z(n7776) );
  NAND U10528 ( .A(n7776), .B(n11562), .Z(n7777) );
  NAND U10529 ( .A(n7777), .B(n11566), .Z(n7778) );
  NANDN U10530 ( .A(n7779), .B(n7778), .Z(n7781) );
  NAND U10531 ( .A(n7781), .B(n7780), .Z(n7783) );
  ANDN U10532 ( .B(n7783), .A(n7782), .Z(n7784) );
  NANDN U10533 ( .A(n7784), .B(n11578), .Z(n7785) );
  NANDN U10534 ( .A(n11581), .B(n7785), .Z(n7786) );
  NAND U10535 ( .A(n7786), .B(n11582), .Z(n7787) );
  NAND U10536 ( .A(n7787), .B(n11584), .Z(n7788) );
  NANDN U10537 ( .A(n11587), .B(n7788), .Z(n7789) );
  NAND U10538 ( .A(n7789), .B(n11589), .Z(n7790) );
  NANDN U10539 ( .A(n11591), .B(n7790), .Z(n7791) );
  NAND U10540 ( .A(n7791), .B(n11592), .Z(n7792) );
  ANDN U10541 ( .B(n7792), .A(n11595), .Z(n7793) );
  NANDN U10542 ( .A(n7793), .B(n11598), .Z(n7794) );
  NANDN U10543 ( .A(n11601), .B(n7794), .Z(n7796) );
  NAND U10544 ( .A(n7796), .B(n7795), .Z(n7797) );
  NANDN U10545 ( .A(n11609), .B(n7797), .Z(n7798) );
  NANDN U10546 ( .A(n11611), .B(n7798), .Z(n7799) );
  NAND U10547 ( .A(n7799), .B(n11613), .Z(n7800) );
  NAND U10548 ( .A(n7800), .B(n11614), .Z(n7801) );
  NAND U10549 ( .A(n7801), .B(n11616), .Z(n7802) );
  ANDN U10550 ( .B(n7802), .A(n11619), .Z(n7803) );
  NANDN U10551 ( .A(n7803), .B(n11620), .Z(n7804) );
  NANDN U10552 ( .A(n11623), .B(n7804), .Z(n7805) );
  NAND U10553 ( .A(n7805), .B(n11625), .Z(n7806) );
  NAND U10554 ( .A(n7806), .B(n11627), .Z(n7807) );
  NAND U10555 ( .A(n7807), .B(n11631), .Z(n7809) );
  ANDN U10556 ( .B(n7809), .A(n7808), .Z(n7812) );
  AND U10557 ( .A(n11634), .B(n7810), .Z(n7811) );
  NANDN U10558 ( .A(n7812), .B(n7811), .Z(n7813) );
  AND U10559 ( .A(n11636), .B(n7813), .Z(n7814) );
  NAND U10560 ( .A(n7815), .B(n7814), .Z(n7816) );
  AND U10561 ( .A(n7817), .B(n7816), .Z(n7820) );
  ANDN U10562 ( .B(n7818), .A(n11645), .Z(n7819) );
  NANDN U10563 ( .A(n7820), .B(n7819), .Z(n7821) );
  ANDN U10564 ( .B(n7821), .A(n11647), .Z(n7822) );
  NANDN U10565 ( .A(n7822), .B(n11648), .Z(n7823) );
  NANDN U10566 ( .A(n11651), .B(n7823), .Z(n7824) );
  NAND U10567 ( .A(n7824), .B(n11652), .Z(n7825) );
  NANDN U10568 ( .A(n11654), .B(n7825), .Z(n7826) );
  NAND U10569 ( .A(n7826), .B(n11657), .Z(n7827) );
  ANDN U10570 ( .B(n7827), .A(n11660), .Z(n7829) );
  NANDN U10571 ( .A(n7829), .B(n7828), .Z(n7830) );
  NANDN U10572 ( .A(n11667), .B(n7830), .Z(n7831) );
  NAND U10573 ( .A(n7831), .B(n11668), .Z(n7832) );
  NAND U10574 ( .A(n7832), .B(n11671), .Z(n7833) );
  NAND U10575 ( .A(n7833), .B(n11672), .Z(n7834) );
  NAND U10576 ( .A(n7834), .B(n11674), .Z(n7835) );
  NANDN U10577 ( .A(n11677), .B(n7835), .Z(n7836) );
  NAND U10578 ( .A(n7836), .B(n11678), .Z(n7837) );
  ANDN U10579 ( .B(n7837), .A(n11681), .Z(n7838) );
  NANDN U10580 ( .A(n7838), .B(n11683), .Z(n7839) );
  NAND U10581 ( .A(n7839), .B(n11685), .Z(n7840) );
  NAND U10582 ( .A(n7840), .B(n11689), .Z(n7841) );
  AND U10583 ( .A(n11690), .B(n7841), .Z(n7843) );
  NAND U10584 ( .A(n7843), .B(n7842), .Z(n7844) );
  NAND U10585 ( .A(n7844), .B(n11692), .Z(n7846) );
  NANDN U10586 ( .A(n7846), .B(n7845), .Z(n7847) );
  ANDN U10587 ( .B(n7847), .A(n11695), .Z(n7848) );
  NAND U10588 ( .A(n7849), .B(n7848), .Z(n7850) );
  NAND U10589 ( .A(n7851), .B(n7850), .Z(n7853) );
  ANDN U10590 ( .B(n7853), .A(n7852), .Z(n7854) );
  NAND U10591 ( .A(n7854), .B(n11702), .Z(n7855) );
  NAND U10592 ( .A(n7855), .B(n11704), .Z(n7856) );
  NANDN U10593 ( .A(n11707), .B(n7856), .Z(n7857) );
  NAND U10594 ( .A(n7857), .B(n11708), .Z(n7858) );
  ANDN U10595 ( .B(n7858), .A(n11711), .Z(n7859) );
  NANDN U10596 ( .A(n7859), .B(n11713), .Z(n7860) );
  NAND U10597 ( .A(n7860), .B(n11714), .Z(n7861) );
  NAND U10598 ( .A(n7861), .B(n11719), .Z(n7862) );
  NANDN U10599 ( .A(n7863), .B(n7862), .Z(n7865) );
  NAND U10600 ( .A(n7865), .B(n7864), .Z(n7867) );
  ANDN U10601 ( .B(n7867), .A(n7866), .Z(n7868) );
  NANDN U10602 ( .A(n7868), .B(n11731), .Z(n7869) );
  NANDN U10603 ( .A(n7870), .B(n7869), .Z(n7871) );
  NAND U10604 ( .A(n7871), .B(n11736), .Z(n7873) );
  ANDN U10605 ( .B(n7873), .A(n7872), .Z(n7874) );
  NAND U10606 ( .A(n7874), .B(n11737), .Z(n7875) );
  NAND U10607 ( .A(n7875), .B(n11739), .Z(n7876) );
  NANDN U10608 ( .A(n11742), .B(n7876), .Z(n7877) );
  NAND U10609 ( .A(n7877), .B(n11743), .Z(n7878) );
  ANDN U10610 ( .B(n7878), .A(n11746), .Z(n7879) );
  NANDN U10611 ( .A(n7879), .B(n11748), .Z(n7880) );
  NAND U10612 ( .A(n7880), .B(n11749), .Z(n7881) );
  NAND U10613 ( .A(n7881), .B(n11754), .Z(n7882) );
  NANDN U10614 ( .A(n7883), .B(n7882), .Z(n7885) );
  NAND U10615 ( .A(n7885), .B(n7884), .Z(n7887) );
  ANDN U10616 ( .B(n7887), .A(n7886), .Z(n7888) );
  NANDN U10617 ( .A(n7888), .B(n11766), .Z(n7889) );
  NANDN U10618 ( .A(n11769), .B(n7889), .Z(n7890) );
  NAND U10619 ( .A(n7890), .B(n11771), .Z(n7891) );
  NAND U10620 ( .A(n7891), .B(n11772), .Z(n7892) );
  NAND U10621 ( .A(n7892), .B(n11774), .Z(n7893) );
  ANDN U10622 ( .B(n7893), .A(n11777), .Z(n7894) );
  NANDN U10623 ( .A(n7894), .B(n11778), .Z(n7895) );
  NANDN U10624 ( .A(n11781), .B(n7895), .Z(n7896) );
  NAND U10625 ( .A(n7896), .B(n11783), .Z(n7897) );
  NANDN U10626 ( .A(n11785), .B(n7897), .Z(n7898) );
  NAND U10627 ( .A(n7898), .B(n11786), .Z(n7899) );
  ANDN U10628 ( .B(n7899), .A(n11789), .Z(n7900) );
  NANDN U10629 ( .A(n7900), .B(n11790), .Z(n7901) );
  NANDN U10630 ( .A(n11793), .B(n7901), .Z(n7902) );
  NAND U10631 ( .A(n7902), .B(n11795), .Z(n7903) );
  NAND U10632 ( .A(n7903), .B(n11796), .Z(n7904) );
  NAND U10633 ( .A(n7904), .B(n11798), .Z(n7905) );
  ANDN U10634 ( .B(n7905), .A(n11801), .Z(n7906) );
  NANDN U10635 ( .A(n7906), .B(n11802), .Z(n7907) );
  NANDN U10636 ( .A(n11805), .B(n7907), .Z(n7908) );
  NAND U10637 ( .A(n7908), .B(n11807), .Z(n7909) );
  NAND U10638 ( .A(n7909), .B(n11809), .Z(n7910) );
  NANDN U10639 ( .A(n11812), .B(n7910), .Z(n7912) );
  ANDN U10640 ( .B(n7912), .A(n7911), .Z(n7913) );
  NANDN U10641 ( .A(n7913), .B(n11818), .Z(n7914) );
  NANDN U10642 ( .A(n11821), .B(n7914), .Z(n7915) );
  NAND U10643 ( .A(n7915), .B(n11823), .Z(n7916) );
  NAND U10644 ( .A(n7916), .B(n11824), .Z(n7917) );
  NAND U10645 ( .A(n7917), .B(n11827), .Z(n7918) );
  ANDN U10646 ( .B(n7918), .A(n11829), .Z(n7919) );
  NANDN U10647 ( .A(n7919), .B(n11830), .Z(n7920) );
  NANDN U10648 ( .A(n11833), .B(n7920), .Z(n7921) );
  NAND U10649 ( .A(n7921), .B(n11834), .Z(n7922) );
  NAND U10650 ( .A(n7922), .B(n11838), .Z(n7923) );
  NAND U10651 ( .A(n7923), .B(n11841), .Z(n7925) );
  ANDN U10652 ( .B(n7925), .A(n7924), .Z(n7928) );
  ANDN U10653 ( .B(n7926), .A(n11845), .Z(n7927) );
  NANDN U10654 ( .A(n7928), .B(n7927), .Z(n7929) );
  AND U10655 ( .A(n11846), .B(n7929), .Z(n7930) );
  NAND U10656 ( .A(n7931), .B(n7930), .Z(n7932) );
  NAND U10657 ( .A(n7933), .B(n7932), .Z(n7935) );
  ANDN U10658 ( .B(n7935), .A(n7934), .Z(n7936) );
  NAND U10659 ( .A(n7936), .B(n11854), .Z(n7937) );
  NAND U10660 ( .A(n7937), .B(n11857), .Z(n7938) );
  NANDN U10661 ( .A(n11859), .B(n7938), .Z(n7939) );
  NAND U10662 ( .A(n7939), .B(n11860), .Z(n7940) );
  ANDN U10663 ( .B(n7940), .A(n11863), .Z(n7941) );
  NANDN U10664 ( .A(n7941), .B(n11864), .Z(n7942) );
  NAND U10665 ( .A(n7942), .B(n11868), .Z(n7943) );
  NAND U10666 ( .A(n7943), .B(n11870), .Z(n7944) );
  NANDN U10667 ( .A(n7945), .B(n7944), .Z(n7946) );
  NAND U10668 ( .A(n7946), .B(n11874), .Z(n7947) );
  ANDN U10669 ( .B(n7947), .A(n11876), .Z(n7948) );
  NANDN U10670 ( .A(n7948), .B(n11878), .Z(n7949) );
  NANDN U10671 ( .A(n11881), .B(n7949), .Z(n7956) );
  NAND U10672 ( .A(n7951), .B(n7950), .Z(n7952) );
  NANDN U10673 ( .A(n7953), .B(n7952), .Z(n7955) );
  ANDN U10674 ( .B(n7955), .A(n7954), .Z(n11882) );
  NAND U10675 ( .A(n7956), .B(n11882), .Z(n7958) );
  NAND U10676 ( .A(n7958), .B(n7957), .Z(n7960) );
  ANDN U10677 ( .B(n7960), .A(n7959), .Z(n7961) );
  NANDN U10678 ( .A(n7961), .B(n11893), .Z(n7962) );
  NANDN U10679 ( .A(n11896), .B(n7962), .Z(n7965) );
  NANDN U10680 ( .A(x[1026]), .B(y[1026]), .Z(n7964) );
  ANDN U10681 ( .B(n7964), .A(n7963), .Z(n11897) );
  NAND U10682 ( .A(n7965), .B(n11897), .Z(n7966) );
  NANDN U10683 ( .A(n11900), .B(n7966), .Z(n7967) );
  AND U10684 ( .A(n7968), .B(n7967), .Z(n7969) );
  NAND U10685 ( .A(n7969), .B(n11901), .Z(n7970) );
  NAND U10686 ( .A(n7971), .B(n7970), .Z(n7972) );
  AND U10687 ( .A(n11909), .B(n7972), .Z(n7973) );
  NANDN U10688 ( .A(n7974), .B(n7973), .Z(n7975) );
  NANDN U10689 ( .A(n11912), .B(n7975), .Z(n7978) );
  NANDN U10690 ( .A(x[1031]), .B(y[1031]), .Z(n7977) );
  NAND U10691 ( .A(n7977), .B(n7976), .Z(n11913) );
  ANDN U10692 ( .B(n7978), .A(n11913), .Z(n7979) );
  OR U10693 ( .A(n11916), .B(n7979), .Z(n7980) );
  NANDN U10694 ( .A(n11918), .B(n7980), .Z(n7981) );
  NAND U10695 ( .A(n7981), .B(n11919), .Z(n7982) );
  NANDN U10696 ( .A(n11922), .B(n7982), .Z(n7983) );
  NAND U10697 ( .A(n7983), .B(n11923), .Z(n7984) );
  ANDN U10698 ( .B(n7984), .A(n11925), .Z(n7985) );
  NANDN U10699 ( .A(n7985), .B(n11927), .Z(n7986) );
  NANDN U10700 ( .A(n11930), .B(n7986), .Z(n7987) );
  NAND U10701 ( .A(n7987), .B(n11931), .Z(n7988) );
  NAND U10702 ( .A(n7988), .B(n11933), .Z(n7991) );
  ANDN U10703 ( .B(n7990), .A(n7989), .Z(n11935) );
  NAND U10704 ( .A(n7991), .B(n11935), .Z(n7994) );
  NANDN U10705 ( .A(x[1043]), .B(y[1043]), .Z(n7993) );
  NAND U10706 ( .A(n7993), .B(n7992), .Z(n11937) );
  ANDN U10707 ( .B(n7994), .A(n11937), .Z(n7995) );
  OR U10708 ( .A(n11940), .B(n7995), .Z(n7996) );
  NANDN U10709 ( .A(n11941), .B(n7996), .Z(n7997) );
  NAND U10710 ( .A(n7997), .B(n11943), .Z(n7998) );
  ANDN U10711 ( .B(n7998), .A(n11945), .Z(n7999) );
  NANDN U10712 ( .A(n7999), .B(n11947), .Z(n8000) );
  NANDN U10713 ( .A(n11950), .B(n8000), .Z(n8003) );
  NOR U10714 ( .A(n8002), .B(n8001), .Z(n11951) );
  NAND U10715 ( .A(n8003), .B(n11951), .Z(n8005) );
  ANDN U10716 ( .B(n8005), .A(n8004), .Z(n8006) );
  NAND U10717 ( .A(n8006), .B(n11954), .Z(n8007) );
  NANDN U10718 ( .A(n8008), .B(n8007), .Z(n8010) );
  ANDN U10719 ( .B(n8010), .A(n8009), .Z(n8011) );
  NAND U10720 ( .A(n8011), .B(n11961), .Z(n8013) );
  NAND U10721 ( .A(n8013), .B(n11963), .Z(n8014) );
  NANDN U10722 ( .A(n11965), .B(n8014), .Z(n8015) );
  AND U10723 ( .A(n11967), .B(n8015), .Z(n8016) );
  NANDN U10724 ( .A(n8016), .B(n11970), .Z(n8017) );
  NANDN U10725 ( .A(n11972), .B(n8017), .Z(n8018) );
  NAND U10726 ( .A(n8018), .B(n11973), .Z(n8019) );
  ANDN U10727 ( .B(n8019), .A(n11976), .Z(n8022) );
  ANDN U10728 ( .B(n8021), .A(n8020), .Z(n11977) );
  NANDN U10729 ( .A(n8022), .B(n11977), .Z(n8025) );
  NANDN U10730 ( .A(y[1062]), .B(x[1062]), .Z(n8024) );
  NAND U10731 ( .A(n8024), .B(n8023), .Z(n11979) );
  ANDN U10732 ( .B(n8025), .A(n11979), .Z(n8027) );
  XNOR U10733 ( .A(x[1064]), .B(y[1064]), .Z(n8026) );
  NANDN U10734 ( .A(n8027), .B(n8026), .Z(n8028) );
  NANDN U10735 ( .A(n8028), .B(n11981), .Z(n8030) );
  ANDN U10736 ( .B(x[1064]), .A(y[1064]), .Z(n11984) );
  ANDN U10737 ( .B(n11988), .A(n11984), .Z(n8029) );
  NAND U10738 ( .A(n8030), .B(n8029), .Z(n8032) );
  NAND U10739 ( .A(n8032), .B(n8031), .Z(n8033) );
  NANDN U10740 ( .A(n8033), .B(n11989), .Z(n8034) );
  NANDN U10741 ( .A(n11991), .B(n8034), .Z(n8035) );
  NANDN U10742 ( .A(n11994), .B(n8035), .Z(n8039) );
  OR U10743 ( .A(y[1068]), .B(n8036), .Z(n8038) );
  NAND U10744 ( .A(n8038), .B(n8037), .Z(n11996) );
  ANDN U10745 ( .B(n8039), .A(n11996), .Z(n8041) );
  NANDN U10746 ( .A(n8041), .B(n8040), .Z(n8043) );
  ANDN U10747 ( .B(n8043), .A(n8042), .Z(n8044) );
  NANDN U10748 ( .A(n8044), .B(n12003), .Z(n8047) );
  NAND U10749 ( .A(n8046), .B(n8045), .Z(n12009) );
  ANDN U10750 ( .B(n8047), .A(n12009), .Z(n8050) );
  ANDN U10751 ( .B(n8048), .A(n12012), .Z(n8049) );
  NANDN U10752 ( .A(n8050), .B(n8049), .Z(n8051) );
  AND U10753 ( .A(n12017), .B(n8051), .Z(n8052) );
  NAND U10754 ( .A(n8052), .B(n12013), .Z(n8053) );
  ANDN U10755 ( .B(n8053), .A(n12020), .Z(n8054) );
  NANDN U10756 ( .A(n8055), .B(n8054), .Z(n8062) );
  NAND U10757 ( .A(n8057), .B(n8056), .Z(n8058) );
  NANDN U10758 ( .A(n8059), .B(n8058), .Z(n8061) );
  ANDN U10759 ( .B(n8061), .A(n8060), .Z(n12021) );
  NAND U10760 ( .A(n8062), .B(n12021), .Z(n8063) );
  NANDN U10761 ( .A(n12024), .B(n8063), .Z(n8064) );
  NAND U10762 ( .A(n8064), .B(n12025), .Z(n8065) );
  ANDN U10763 ( .B(n8065), .A(n12028), .Z(n8066) );
  NANDN U10764 ( .A(n8066), .B(n12030), .Z(n8067) );
  NAND U10765 ( .A(n8067), .B(n12031), .Z(n8070) );
  NOR U10766 ( .A(n8069), .B(n8068), .Z(n12034) );
  NAND U10767 ( .A(n8070), .B(n12034), .Z(n8071) );
  AND U10768 ( .A(n12035), .B(n8071), .Z(n8072) );
  NANDN U10769 ( .A(n8073), .B(n8072), .Z(n8074) );
  NAND U10770 ( .A(n8074), .B(n12041), .Z(n8075) );
  NANDN U10771 ( .A(n8075), .B(n12037), .Z(n8076) );
  AND U10772 ( .A(n8077), .B(n8076), .Z(n8079) );
  NANDN U10773 ( .A(n8079), .B(n12046), .Z(n8080) );
  NANDN U10774 ( .A(n12048), .B(n8080), .Z(n8083) );
  NANDN U10775 ( .A(y[1092]), .B(x[1092]), .Z(n8081) );
  NANDN U10776 ( .A(n8082), .B(n8081), .Z(n12050) );
  ANDN U10777 ( .B(n8083), .A(n12050), .Z(n8084) );
  NANDN U10778 ( .A(n8084), .B(n12051), .Z(n8085) );
  NANDN U10779 ( .A(n12053), .B(n8085), .Z(n8086) );
  NANDN U10780 ( .A(n12056), .B(n8086), .Z(n8087) );
  NANDN U10781 ( .A(n12057), .B(n8087), .Z(n8088) );
  AND U10782 ( .A(n8089), .B(n8088), .Z(n8090) );
  NAND U10783 ( .A(n8090), .B(n12059), .Z(n8091) );
  NAND U10784 ( .A(n8092), .B(n8091), .Z(n8093) );
  AND U10785 ( .A(n12067), .B(n8093), .Z(n8095) );
  NAND U10786 ( .A(n8095), .B(n8094), .Z(n8096) );
  NANDN U10787 ( .A(n12069), .B(n8096), .Z(n8097) );
  NANDN U10788 ( .A(n12072), .B(n8097), .Z(n8098) );
  NANDN U10789 ( .A(n12074), .B(n8098), .Z(n8101) );
  NANDN U10790 ( .A(x[1105]), .B(y[1105]), .Z(n8100) );
  ANDN U10791 ( .B(n8100), .A(n8099), .Z(n12075) );
  NAND U10792 ( .A(n8101), .B(n12075), .Z(n8102) );
  ANDN U10793 ( .B(n8102), .A(n12078), .Z(n8103) );
  NANDN U10794 ( .A(n8103), .B(n12079), .Z(n8104) );
  NANDN U10795 ( .A(n12081), .B(n8104), .Z(n8105) );
  NANDN U10796 ( .A(n8106), .B(n8105), .Z(n8107) );
  NANDN U10797 ( .A(n8108), .B(n8107), .Z(n8109) );
  AND U10798 ( .A(n8110), .B(n8109), .Z(n8112) );
  NANDN U10799 ( .A(n8112), .B(n8111), .Z(n8113) );
  NANDN U10800 ( .A(n8114), .B(n8113), .Z(n8117) );
  ANDN U10801 ( .B(n8116), .A(n8115), .Z(n12089) );
  NAND U10802 ( .A(n8117), .B(n12089), .Z(n8118) );
  AND U10803 ( .A(n12092), .B(n8118), .Z(n8119) );
  NANDN U10804 ( .A(n8119), .B(n12093), .Z(n8120) );
  ANDN U10805 ( .B(n8120), .A(n12096), .Z(n8121) );
  NANDN U10806 ( .A(n8121), .B(n12097), .Z(n8122) );
  NANDN U10807 ( .A(n12100), .B(n8122), .Z(n8123) );
  NAND U10808 ( .A(n8123), .B(n12101), .Z(n8124) );
  NANDN U10809 ( .A(n12103), .B(n8124), .Z(n8125) );
  NANDN U10810 ( .A(n12106), .B(n8125), .Z(n8127) );
  NAND U10811 ( .A(n8127), .B(n8126), .Z(n8128) );
  NANDN U10812 ( .A(n8128), .B(n12107), .Z(n8130) );
  NOR U10813 ( .A(n12114), .B(n8129), .Z(n12109) );
  NAND U10814 ( .A(n8130), .B(n12109), .Z(n8131) );
  NAND U10815 ( .A(n8131), .B(n12111), .Z(n8133) );
  NANDN U10816 ( .A(n8133), .B(n8132), .Z(n8136) );
  NANDN U10817 ( .A(y[1127]), .B(x[1127]), .Z(n8135) );
  ANDN U10818 ( .B(n8135), .A(n8134), .Z(n12117) );
  NAND U10819 ( .A(n8136), .B(n12117), .Z(n8137) );
  NANDN U10820 ( .A(n12120), .B(n8137), .Z(n8140) );
  NANDN U10821 ( .A(y[1128]), .B(x[1128]), .Z(n8139) );
  ANDN U10822 ( .B(n8139), .A(n8138), .Z(n12121) );
  NAND U10823 ( .A(n8140), .B(n12121), .Z(n8143) );
  ANDN U10824 ( .B(n8143), .A(n12124), .Z(n8144) );
  NANDN U10825 ( .A(n8144), .B(n12125), .Z(n8145) );
  NANDN U10826 ( .A(n12127), .B(n8145), .Z(n8146) );
  NAND U10827 ( .A(n8146), .B(n12129), .Z(n8149) );
  ANDN U10828 ( .B(n8148), .A(n8147), .Z(n12131) );
  NAND U10829 ( .A(n8149), .B(n12131), .Z(n8152) );
  NANDN U10830 ( .A(y[1134]), .B(x[1134]), .Z(n8151) );
  NAND U10831 ( .A(n8151), .B(n8150), .Z(n12134) );
  ANDN U10832 ( .B(n8152), .A(n12134), .Z(n8153) );
  NANDN U10833 ( .A(n8153), .B(n12136), .Z(n8155) );
  NANDN U10834 ( .A(n8155), .B(n8154), .Z(n8157) );
  AND U10835 ( .A(n12137), .B(n12139), .Z(n8156) );
  NAND U10836 ( .A(n8157), .B(n8156), .Z(n8159) );
  NAND U10837 ( .A(n8159), .B(n8158), .Z(n8160) );
  NANDN U10838 ( .A(n8160), .B(n12140), .Z(n8164) );
  OR U10839 ( .A(y[1139]), .B(n8161), .Z(n8162) );
  NAND U10840 ( .A(n8163), .B(n8162), .Z(n12141) );
  ANDN U10841 ( .B(n8164), .A(n12141), .Z(n8165) );
  OR U10842 ( .A(n12142), .B(n8165), .Z(n8168) );
  NANDN U10843 ( .A(y[1140]), .B(x[1140]), .Z(n8167) );
  ANDN U10844 ( .B(n8167), .A(n8166), .Z(n12143) );
  NAND U10845 ( .A(n8168), .B(n12143), .Z(n8169) );
  NAND U10846 ( .A(n8169), .B(n12144), .Z(n8171) );
  NANDN U10847 ( .A(n8171), .B(n8170), .Z(n8172) );
  AND U10848 ( .A(n8173), .B(n8172), .Z(n8176) );
  ANDN U10849 ( .B(n8174), .A(n10002), .Z(n8175) );
  NANDN U10850 ( .A(n8176), .B(n8175), .Z(n8177) );
  AND U10851 ( .A(n8178), .B(n8177), .Z(n8179) );
  NANDN U10852 ( .A(n8179), .B(n12149), .Z(n8180) );
  NANDN U10853 ( .A(n12150), .B(n8180), .Z(n8182) );
  NAND U10854 ( .A(n8182), .B(n8181), .Z(n8183) );
  NANDN U10855 ( .A(n8183), .B(n12151), .Z(n8184) );
  NANDN U10856 ( .A(n12152), .B(n8184), .Z(n8185) );
  NAND U10857 ( .A(n8185), .B(n10001), .Z(n8187) );
  NANDN U10858 ( .A(n8187), .B(n8186), .Z(n8190) );
  NANDN U10859 ( .A(y[1151]), .B(x[1151]), .Z(n8188) );
  NAND U10860 ( .A(n8189), .B(n8188), .Z(n12156) );
  ANDN U10861 ( .B(n8190), .A(n12156), .Z(n8191) );
  OR U10862 ( .A(n12158), .B(n8191), .Z(n8192) );
  NANDN U10863 ( .A(n12160), .B(n8192), .Z(n8193) );
  NAND U10864 ( .A(n8193), .B(n12161), .Z(n8194) );
  NANDN U10865 ( .A(n12164), .B(n8194), .Z(n8195) );
  AND U10866 ( .A(n8195), .B(n12167), .Z(n8196) );
  OR U10867 ( .A(n8196), .B(x[1156]), .Z(n8199) );
  XOR U10868 ( .A(x[1156]), .B(n8196), .Z(n8197) );
  NAND U10869 ( .A(y[1156]), .B(n8197), .Z(n8198) );
  NAND U10870 ( .A(n8199), .B(n8198), .Z(n8200) );
  AND U10871 ( .A(n9999), .B(n8200), .Z(n8201) );
  OR U10872 ( .A(n12172), .B(n8201), .Z(n8204) );
  NANDN U10873 ( .A(y[1158]), .B(x[1158]), .Z(n8203) );
  NAND U10874 ( .A(n8203), .B(n8202), .Z(n12174) );
  ANDN U10875 ( .B(n8204), .A(n12174), .Z(n8207) );
  AND U10876 ( .A(n12175), .B(n8205), .Z(n8206) );
  NANDN U10877 ( .A(n8207), .B(n8206), .Z(n8208) );
  NANDN U10878 ( .A(n8209), .B(n8208), .Z(n8211) );
  ANDN U10879 ( .B(n8211), .A(n8210), .Z(n8212) );
  NAND U10880 ( .A(n8212), .B(n12183), .Z(n8215) );
  NOR U10881 ( .A(n8214), .B(n8213), .Z(n12186) );
  NAND U10882 ( .A(n8215), .B(n12186), .Z(n8216) );
  NANDN U10883 ( .A(n12188), .B(n8216), .Z(n8217) );
  NANDN U10884 ( .A(n12190), .B(n8217), .Z(n8221) );
  OR U10885 ( .A(x[1165]), .B(n8218), .Z(n8220) );
  NAND U10886 ( .A(n8220), .B(n8219), .Z(n12192) );
  ANDN U10887 ( .B(n8221), .A(n12192), .Z(n8222) );
  NANDN U10888 ( .A(n8222), .B(n12193), .Z(n8223) );
  ANDN U10889 ( .B(n8223), .A(n12196), .Z(n8224) );
  OR U10890 ( .A(n12198), .B(n8224), .Z(n8226) );
  NAND U10891 ( .A(n8226), .B(n12199), .Z(n8229) );
  NANDN U10892 ( .A(y[1170]), .B(x[1170]), .Z(n8228) );
  NAND U10893 ( .A(n8228), .B(n8227), .Z(n12201) );
  ANDN U10894 ( .B(n8229), .A(n12201), .Z(n8232) );
  ANDN U10895 ( .B(n8230), .A(n12204), .Z(n8231) );
  NANDN U10896 ( .A(n8232), .B(n8231), .Z(n8233) );
  AND U10897 ( .A(n12209), .B(n8233), .Z(n8234) );
  NAND U10898 ( .A(n8234), .B(n12205), .Z(n8235) );
  AND U10899 ( .A(n8236), .B(n8235), .Z(n8237) );
  NAND U10900 ( .A(n8237), .B(n12211), .Z(n8238) );
  NANDN U10901 ( .A(n12213), .B(n8238), .Z(n8239) );
  NANDN U10902 ( .A(n12216), .B(n8239), .Z(n8240) );
  ANDN U10903 ( .B(n8240), .A(n12217), .Z(n8241) );
  NANDN U10904 ( .A(n8241), .B(n12219), .Z(n8242) );
  ANDN U10905 ( .B(n8242), .A(n12221), .Z(n8245) );
  AND U10906 ( .A(n12223), .B(n8243), .Z(n8244) );
  NANDN U10907 ( .A(n8245), .B(n8244), .Z(n8246) );
  AND U10908 ( .A(n12225), .B(n8246), .Z(n8247) );
  NAND U10909 ( .A(n8248), .B(n8247), .Z(n8249) );
  NAND U10910 ( .A(n8250), .B(n8249), .Z(n8252) );
  ANDN U10911 ( .B(n8252), .A(n8251), .Z(n8256) );
  ANDN U10912 ( .B(n8254), .A(n8253), .Z(n8255) );
  NANDN U10913 ( .A(n8256), .B(n8255), .Z(n8257) );
  NANDN U10914 ( .A(n8258), .B(n8257), .Z(n8260) );
  ANDN U10915 ( .B(n8260), .A(n8259), .Z(n8261) );
  NANDN U10916 ( .A(n12240), .B(n8261), .Z(n8262) );
  NANDN U10917 ( .A(n12241), .B(n8262), .Z(n8263) );
  NANDN U10918 ( .A(n12244), .B(n8263), .Z(n8266) );
  NANDN U10919 ( .A(y[1188]), .B(x[1188]), .Z(n8265) );
  NAND U10920 ( .A(n8265), .B(n8264), .Z(n12245) );
  ANDN U10921 ( .B(n8266), .A(n12245), .Z(n8267) );
  NANDN U10922 ( .A(n8267), .B(n12247), .Z(n8268) );
  NANDN U10923 ( .A(n12250), .B(n8268), .Z(n8269) );
  NAND U10924 ( .A(n8269), .B(n12251), .Z(n8270) );
  ANDN U10925 ( .B(n8270), .A(n12253), .Z(n8273) );
  NANDN U10926 ( .A(x[1194]), .B(y[1194]), .Z(n8271) );
  NAND U10927 ( .A(n8272), .B(n8271), .Z(n12256) );
  OR U10928 ( .A(n8273), .B(n12256), .Z(n8276) );
  NANDN U10929 ( .A(y[1194]), .B(x[1194]), .Z(n8275) );
  NAND U10930 ( .A(n8275), .B(n8274), .Z(n12257) );
  ANDN U10931 ( .B(n8276), .A(n12257), .Z(n8279) );
  AND U10932 ( .A(n12259), .B(n8277), .Z(n8278) );
  NANDN U10933 ( .A(n8279), .B(n8278), .Z(n8280) );
  AND U10934 ( .A(n12265), .B(n8280), .Z(n8281) );
  NAND U10935 ( .A(n8281), .B(n12261), .Z(n8282) );
  ANDN U10936 ( .B(n8282), .A(n12268), .Z(n8283) );
  NANDN U10937 ( .A(n8284), .B(n8283), .Z(n8291) );
  NANDN U10938 ( .A(n8286), .B(n8285), .Z(n8287) );
  NANDN U10939 ( .A(n8288), .B(n8287), .Z(n8290) );
  ANDN U10940 ( .B(n8290), .A(n8289), .Z(n12269) );
  NAND U10941 ( .A(n8291), .B(n12269), .Z(n8292) );
  NANDN U10942 ( .A(n12272), .B(n8292), .Z(n8293) );
  NAND U10943 ( .A(n8293), .B(n12273), .Z(n8294) );
  ANDN U10944 ( .B(n8294), .A(n12276), .Z(n8295) );
  NANDN U10945 ( .A(n8295), .B(n12277), .Z(n8296) );
  NAND U10946 ( .A(n8296), .B(n12279), .Z(n8297) );
  NANDN U10947 ( .A(n12281), .B(n8297), .Z(n8298) );
  ANDN U10948 ( .B(n8298), .A(n12284), .Z(n8299) );
  NANDN U10949 ( .A(n8300), .B(n8299), .Z(n8301) );
  NAND U10950 ( .A(n8301), .B(n12285), .Z(n8302) );
  NANDN U10951 ( .A(n8302), .B(n12289), .Z(n8303) );
  AND U10952 ( .A(n8304), .B(n8303), .Z(n8305) );
  NANDN U10953 ( .A(n8305), .B(n12293), .Z(n8306) );
  ANDN U10954 ( .B(n8306), .A(n12295), .Z(n8307) );
  NANDN U10955 ( .A(n8307), .B(n12297), .Z(n8308) );
  NANDN U10956 ( .A(n12300), .B(n8308), .Z(n8309) );
  NAND U10957 ( .A(n8309), .B(n12301), .Z(n8310) );
  NANDN U10958 ( .A(n12304), .B(n8310), .Z(n8311) );
  NAND U10959 ( .A(n8311), .B(n12305), .Z(n8312) );
  ANDN U10960 ( .B(n8312), .A(n12307), .Z(n8313) );
  NANDN U10961 ( .A(n8313), .B(n12309), .Z(n8314) );
  AND U10962 ( .A(n8315), .B(n8314), .Z(n8316) );
  OR U10963 ( .A(n12313), .B(n8316), .Z(n8317) );
  AND U10964 ( .A(n8318), .B(n8317), .Z(n8319) );
  OR U10965 ( .A(n12317), .B(n8319), .Z(n8320) );
  NANDN U10966 ( .A(n12318), .B(n8320), .Z(n8323) );
  NANDN U10967 ( .A(y[1224]), .B(x[1224]), .Z(n8322) );
  ANDN U10968 ( .B(n8322), .A(n8321), .Z(n12319) );
  NAND U10969 ( .A(n8323), .B(n12319), .Z(n8324) );
  NAND U10970 ( .A(n8324), .B(n12320), .Z(n8325) );
  NAND U10971 ( .A(n8325), .B(n12321), .Z(n8326) );
  ANDN U10972 ( .B(n8326), .A(n12322), .Z(n8327) );
  NANDN U10973 ( .A(n8327), .B(n12323), .Z(n8330) );
  NOR U10974 ( .A(n8329), .B(n8328), .Z(n12324) );
  NAND U10975 ( .A(n8330), .B(n12324), .Z(n8333) );
  ANDN U10976 ( .B(n8332), .A(n8331), .Z(n12325) );
  NAND U10977 ( .A(n8333), .B(n12325), .Z(n8334) );
  ANDN U10978 ( .B(n8334), .A(n12326), .Z(n8335) );
  NANDN U10979 ( .A(n8336), .B(n8335), .Z(n8337) );
  NAND U10980 ( .A(n8337), .B(n12329), .Z(n8338) );
  NANDN U10981 ( .A(n8338), .B(n12327), .Z(n8339) );
  AND U10982 ( .A(n8340), .B(n8339), .Z(n8342) );
  NANDN U10983 ( .A(n8342), .B(n12332), .Z(n8343) );
  NANDN U10984 ( .A(n12334), .B(n8343), .Z(n8346) );
  NANDN U10985 ( .A(y[1236]), .B(x[1236]), .Z(n8345) );
  ANDN U10986 ( .B(n8345), .A(n8344), .Z(n12335) );
  NAND U10987 ( .A(n8346), .B(n12335), .Z(n8348) );
  NAND U10988 ( .A(n8348), .B(n8347), .Z(n8349) );
  NANDN U10989 ( .A(n12339), .B(n8349), .Z(n8351) );
  NAND U10990 ( .A(n8351), .B(n8350), .Z(n8352) );
  NANDN U10991 ( .A(n8353), .B(n8352), .Z(n8354) );
  NAND U10992 ( .A(n8354), .B(n12353), .Z(n8357) );
  NOR U10993 ( .A(n8356), .B(n8355), .Z(n12356) );
  NAND U10994 ( .A(n8357), .B(n12356), .Z(n8359) );
  ANDN U10995 ( .B(n8359), .A(n8358), .Z(n8360) );
  NAND U10996 ( .A(n8360), .B(n12357), .Z(n8361) );
  NANDN U10997 ( .A(n8362), .B(n8361), .Z(n8364) );
  ANDN U10998 ( .B(n8364), .A(n8363), .Z(n8365) );
  NAND U10999 ( .A(n8365), .B(n12365), .Z(n8368) );
  NOR U11000 ( .A(n8367), .B(n8366), .Z(n12367) );
  NAND U11001 ( .A(n8368), .B(n12367), .Z(n8369) );
  NANDN U11002 ( .A(n12370), .B(n8369), .Z(n8370) );
  NANDN U11003 ( .A(n12371), .B(n8370), .Z(n8371) );
  ANDN U11004 ( .B(n8371), .A(n12372), .Z(n8372) );
  NANDN U11005 ( .A(n8372), .B(n12373), .Z(n8373) );
  AND U11006 ( .A(n12374), .B(n8373), .Z(n8374) );
  NANDN U11007 ( .A(n8375), .B(n8374), .Z(n8376) );
  AND U11008 ( .A(n12377), .B(n8376), .Z(n8377) );
  NAND U11009 ( .A(n8377), .B(n12375), .Z(n8379) );
  ANDN U11010 ( .B(n8379), .A(n8378), .Z(n8380) );
  NANDN U11011 ( .A(n8381), .B(n8380), .Z(n8382) );
  NANDN U11012 ( .A(n12380), .B(n8382), .Z(n8383) );
  ANDN U11013 ( .B(n8383), .A(n12381), .Z(n8384) );
  NANDN U11014 ( .A(n8385), .B(n8384), .Z(n8386) );
  NAND U11015 ( .A(n8386), .B(n12383), .Z(n8387) );
  NANDN U11016 ( .A(n8387), .B(n12379), .Z(n8388) );
  NAND U11017 ( .A(n8389), .B(n8388), .Z(n8396) );
  OR U11018 ( .A(n8391), .B(n8390), .Z(n8392) );
  NANDN U11019 ( .A(n8393), .B(n8392), .Z(n8395) );
  ANDN U11020 ( .B(n8395), .A(n8394), .Z(n12385) );
  NAND U11021 ( .A(n8396), .B(n12385), .Z(n8397) );
  ANDN U11022 ( .B(n8397), .A(n12386), .Z(n8398) );
  OR U11023 ( .A(n12387), .B(n8398), .Z(n8399) );
  NANDN U11024 ( .A(n12388), .B(n8399), .Z(n8402) );
  ANDN U11025 ( .B(n8401), .A(n8400), .Z(n12389) );
  NAND U11026 ( .A(n8402), .B(n12389), .Z(n8403) );
  NANDN U11027 ( .A(n12391), .B(n8403), .Z(n8404) );
  NANDN U11028 ( .A(n12394), .B(n8404), .Z(n8408) );
  OR U11029 ( .A(x[1271]), .B(n8405), .Z(n8407) );
  NAND U11030 ( .A(n8407), .B(n8406), .Z(n12396) );
  ANDN U11031 ( .B(n8408), .A(n12396), .Z(n8409) );
  OR U11032 ( .A(n12398), .B(n8409), .Z(n8412) );
  NANDN U11033 ( .A(x[1273]), .B(y[1273]), .Z(n8411) );
  ANDN U11034 ( .B(n8411), .A(n8410), .Z(n12399) );
  NAND U11035 ( .A(n8412), .B(n12399), .Z(n8413) );
  NANDN U11036 ( .A(n12401), .B(n8413), .Z(n8417) );
  OR U11037 ( .A(x[1275]), .B(n8414), .Z(n8415) );
  NAND U11038 ( .A(n8416), .B(n8415), .Z(n12403) );
  ANDN U11039 ( .B(n8417), .A(n12403), .Z(n8418) );
  NANDN U11040 ( .A(n8418), .B(n12405), .Z(n8420) );
  ANDN U11041 ( .B(n8420), .A(n8419), .Z(n8421) );
  OR U11042 ( .A(n8422), .B(n8421), .Z(n8424) );
  ANDN U11043 ( .B(n8424), .A(n8423), .Z(n8425) );
  NAND U11044 ( .A(n8426), .B(n8425), .Z(n8427) );
  NAND U11045 ( .A(n8428), .B(n8427), .Z(n8430) );
  ANDN U11046 ( .B(n8430), .A(n8429), .Z(n8431) );
  NAND U11047 ( .A(n8431), .B(n12415), .Z(n8434) );
  NOR U11048 ( .A(n8433), .B(n8432), .Z(n12417) );
  NAND U11049 ( .A(n8434), .B(n12417), .Z(n8437) );
  NANDN U11050 ( .A(x[1284]), .B(y[1284]), .Z(n8435) );
  NAND U11051 ( .A(n8436), .B(n8435), .Z(n12419) );
  ANDN U11052 ( .B(n8437), .A(n12419), .Z(n8438) );
  OR U11053 ( .A(n12422), .B(n8438), .Z(n8439) );
  NANDN U11054 ( .A(n12424), .B(n8439), .Z(n8440) );
  NAND U11055 ( .A(n8440), .B(n12425), .Z(n8441) );
  ANDN U11056 ( .B(n8441), .A(n12427), .Z(n8442) );
  NANDN U11057 ( .A(n8442), .B(n12429), .Z(n8443) );
  NANDN U11058 ( .A(n12432), .B(n8443), .Z(n8446) );
  ANDN U11059 ( .B(n8445), .A(n8444), .Z(n12433) );
  NAND U11060 ( .A(n8446), .B(n12433), .Z(n8448) );
  AND U11061 ( .A(n8448), .B(n8447), .Z(n8449) );
  NAND U11062 ( .A(n8449), .B(n12436), .Z(n8450) );
  NANDN U11063 ( .A(n8451), .B(n8450), .Z(n8453) );
  AND U11064 ( .A(n8453), .B(n8452), .Z(n8454) );
  NAND U11065 ( .A(n8454), .B(n12443), .Z(n8455) );
  NANDN U11066 ( .A(n12446), .B(n8455), .Z(n8458) );
  NANDN U11067 ( .A(x[1295]), .B(y[1295]), .Z(n8457) );
  ANDN U11068 ( .B(n8457), .A(n8456), .Z(n12448) );
  NAND U11069 ( .A(n8458), .B(n12448), .Z(n8461) );
  NAND U11070 ( .A(n8460), .B(n8459), .Z(n12449) );
  ANDN U11071 ( .B(n8461), .A(n12449), .Z(n8462) );
  OR U11072 ( .A(n12451), .B(n8462), .Z(n8463) );
  NAND U11073 ( .A(n8463), .B(n12453), .Z(n8464) );
  ANDN U11074 ( .B(n8464), .A(n12456), .Z(n8465) );
  NANDN U11075 ( .A(n8465), .B(n12458), .Z(n8466) );
  NAND U11076 ( .A(n8466), .B(n12459), .Z(n8469) );
  ANDN U11077 ( .B(n8468), .A(n8467), .Z(n12462) );
  NAND U11078 ( .A(n8469), .B(n12462), .Z(n8470) );
  AND U11079 ( .A(n12463), .B(n8470), .Z(n8471) );
  NANDN U11080 ( .A(n8472), .B(n8471), .Z(n8473) );
  NAND U11081 ( .A(n8473), .B(n12469), .Z(n8474) );
  NANDN U11082 ( .A(n8474), .B(n12465), .Z(n8475) );
  AND U11083 ( .A(n8476), .B(n8475), .Z(n8479) );
  ANDN U11084 ( .B(n8478), .A(n8477), .Z(n12474) );
  NANDN U11085 ( .A(n8479), .B(n12474), .Z(n8482) );
  NANDN U11086 ( .A(x[1307]), .B(y[1307]), .Z(n8481) );
  ANDN U11087 ( .B(n8481), .A(n8480), .Z(n12475) );
  NAND U11088 ( .A(n8482), .B(n12475), .Z(n8483) );
  NANDN U11089 ( .A(n12478), .B(n8483), .Z(n8486) );
  NANDN U11090 ( .A(x[1309]), .B(y[1309]), .Z(n8485) );
  ANDN U11091 ( .B(n8485), .A(n8484), .Z(n12479) );
  NAND U11092 ( .A(n8486), .B(n12479), .Z(n8487) );
  NAND U11093 ( .A(n8487), .B(n12481), .Z(n8488) );
  ANDN U11094 ( .B(n8488), .A(n12484), .Z(n8489) );
  NANDN U11095 ( .A(n8489), .B(n12486), .Z(n8490) );
  NANDN U11096 ( .A(n12488), .B(n8490), .Z(n8493) );
  NOR U11097 ( .A(n8492), .B(n8491), .Z(n12490) );
  NAND U11098 ( .A(n8493), .B(n12490), .Z(n8494) );
  AND U11099 ( .A(n12491), .B(n8494), .Z(n8495) );
  NANDN U11100 ( .A(n8496), .B(n8495), .Z(n8497) );
  NAND U11101 ( .A(n8497), .B(n12498), .Z(n8498) );
  NANDN U11102 ( .A(n8498), .B(n12493), .Z(n8499) );
  AND U11103 ( .A(n8500), .B(n8499), .Z(n8501) );
  OR U11104 ( .A(n12502), .B(n8501), .Z(n8502) );
  NANDN U11105 ( .A(n12504), .B(n8502), .Z(n8505) );
  NANDN U11106 ( .A(y[1320]), .B(x[1320]), .Z(n8503) );
  AND U11107 ( .A(n8504), .B(n8503), .Z(n12505) );
  NAND U11108 ( .A(n8505), .B(n12505), .Z(n8506) );
  NANDN U11109 ( .A(n12507), .B(n8506), .Z(n8507) );
  NAND U11110 ( .A(n8507), .B(n12509), .Z(n8508) );
  ANDN U11111 ( .B(n8508), .A(n12511), .Z(n8509) );
  NANDN U11112 ( .A(n8509), .B(n12513), .Z(n8510) );
  ANDN U11113 ( .B(n8510), .A(n12515), .Z(n8511) );
  OR U11114 ( .A(n12518), .B(n8511), .Z(n8512) );
  NAND U11115 ( .A(n8513), .B(n8512), .Z(n8514) );
  AND U11116 ( .A(n12525), .B(n8514), .Z(n8515) );
  NAND U11117 ( .A(n8515), .B(n12521), .Z(n8516) );
  AND U11118 ( .A(n12528), .B(n8516), .Z(n8518) );
  NAND U11119 ( .A(n8518), .B(n8517), .Z(n8525) );
  NAND U11120 ( .A(n8520), .B(n8519), .Z(n8521) );
  NANDN U11121 ( .A(n8522), .B(n8521), .Z(n8524) );
  ANDN U11122 ( .B(n8524), .A(n8523), .Z(n12529) );
  NAND U11123 ( .A(n8525), .B(n12529), .Z(n8526) );
  ANDN U11124 ( .B(n8526), .A(n12531), .Z(n8527) );
  NANDN U11125 ( .A(n8527), .B(n12533), .Z(n8528) );
  NANDN U11126 ( .A(n12535), .B(n8528), .Z(n8529) );
  NAND U11127 ( .A(n8529), .B(n12537), .Z(n8530) );
  NANDN U11128 ( .A(n12540), .B(n8530), .Z(n8531) );
  NANDN U11129 ( .A(n12542), .B(n8531), .Z(n8532) );
  NAND U11130 ( .A(n8532), .B(n12544), .Z(n8534) );
  NANDN U11131 ( .A(n8534), .B(n8533), .Z(n8535) );
  AND U11132 ( .A(n8536), .B(n8535), .Z(n8537) );
  ANDN U11133 ( .B(n12551), .A(n8537), .Z(n8538) );
  NANDN U11134 ( .A(n8539), .B(n8538), .Z(n8542) );
  NANDN U11135 ( .A(y[1343]), .B(x[1343]), .Z(n8541) );
  ANDN U11136 ( .B(n8541), .A(n8540), .Z(n12554) );
  NAND U11137 ( .A(n8542), .B(n12554), .Z(n8547) );
  NANDN U11138 ( .A(n8544), .B(n8543), .Z(n8546) );
  NANDN U11139 ( .A(x[1344]), .B(y[1344]), .Z(n8545) );
  NAND U11140 ( .A(n8546), .B(n8545), .Z(n12556) );
  ANDN U11141 ( .B(n8547), .A(n12556), .Z(n8550) );
  NANDN U11142 ( .A(y[1344]), .B(x[1344]), .Z(n8548) );
  AND U11143 ( .A(n8549), .B(n8548), .Z(n12557) );
  NANDN U11144 ( .A(n8550), .B(n12557), .Z(n8551) );
  NANDN U11145 ( .A(n12560), .B(n8551), .Z(n8552) );
  NAND U11146 ( .A(n8552), .B(n12561), .Z(n8553) );
  NANDN U11147 ( .A(n12564), .B(n8553), .Z(n8554) );
  NAND U11148 ( .A(n8554), .B(n12566), .Z(n8555) );
  NAND U11149 ( .A(n8555), .B(n12567), .Z(n8558) );
  NAND U11150 ( .A(n8557), .B(n8556), .Z(n12569) );
  ANDN U11151 ( .B(n8558), .A(n12569), .Z(n8561) );
  ANDN U11152 ( .B(n12571), .A(n8559), .Z(n8560) );
  NANDN U11153 ( .A(n8561), .B(n8560), .Z(n8562) );
  NANDN U11154 ( .A(n8563), .B(n8562), .Z(n8564) );
  AND U11155 ( .A(n12579), .B(n8564), .Z(n8565) );
  NANDN U11156 ( .A(n8566), .B(n8565), .Z(n8567) );
  NANDN U11157 ( .A(n12582), .B(n8567), .Z(n8568) );
  NANDN U11158 ( .A(n12583), .B(n8568), .Z(n8569) );
  NAND U11159 ( .A(n8569), .B(n12585), .Z(n8570) );
  ANDN U11160 ( .B(n8570), .A(n12587), .Z(n8571) );
  NANDN U11161 ( .A(n8571), .B(n12589), .Z(n8572) );
  ANDN U11162 ( .B(n8572), .A(n12591), .Z(n8573) );
  NANDN U11163 ( .A(n8573), .B(n12593), .Z(n8574) );
  NANDN U11164 ( .A(n8575), .B(n8574), .Z(n8577) );
  NAND U11165 ( .A(n8577), .B(n8576), .Z(n8579) );
  ANDN U11166 ( .B(n8579), .A(n8578), .Z(n8581) );
  NAND U11167 ( .A(n8581), .B(n8580), .Z(n8582) );
  NAND U11168 ( .A(n8582), .B(n12601), .Z(n8584) );
  NANDN U11169 ( .A(n8584), .B(n8583), .Z(n8585) );
  AND U11170 ( .A(n8586), .B(n8585), .Z(n8587) );
  NAND U11171 ( .A(n8587), .B(n12603), .Z(n8589) );
  NAND U11172 ( .A(n8589), .B(n12606), .Z(n8594) );
  NANDN U11173 ( .A(n8591), .B(n8590), .Z(n8592) );
  NAND U11174 ( .A(n8593), .B(n8592), .Z(n12608) );
  ANDN U11175 ( .B(n8594), .A(n12608), .Z(n8597) );
  NANDN U11176 ( .A(y[1368]), .B(x[1368]), .Z(n8596) );
  ANDN U11177 ( .B(n8596), .A(n8595), .Z(n12609) );
  NANDN U11178 ( .A(n8597), .B(n12609), .Z(n8598) );
  NANDN U11179 ( .A(n12612), .B(n8598), .Z(n8599) );
  NAND U11180 ( .A(n8599), .B(n12613), .Z(n8600) );
  NAND U11181 ( .A(n8600), .B(n12615), .Z(n8601) );
  ANDN U11182 ( .B(n8601), .A(n12617), .Z(n8602) );
  OR U11183 ( .A(n12620), .B(n8602), .Z(n8603) );
  NANDN U11184 ( .A(n12621), .B(n8603), .Z(n8606) );
  NANDN U11185 ( .A(x[1378]), .B(y[1378]), .Z(n8604) );
  NANDN U11186 ( .A(n8605), .B(n8604), .Z(n12624) );
  ANDN U11187 ( .B(n8606), .A(n12624), .Z(n8607) );
  OR U11188 ( .A(n12626), .B(n8607), .Z(n8610) );
  NANDN U11189 ( .A(x[1379]), .B(y[1379]), .Z(n8609) );
  ANDN U11190 ( .B(n8609), .A(n8608), .Z(n12627) );
  NAND U11191 ( .A(n8610), .B(n12627), .Z(n8611) );
  NANDN U11192 ( .A(n12630), .B(n8611), .Z(n8612) );
  NANDN U11193 ( .A(n12632), .B(n8612), .Z(n8615) );
  NANDN U11194 ( .A(y[1382]), .B(x[1382]), .Z(n8614) );
  NAND U11195 ( .A(n8614), .B(n8613), .Z(n12633) );
  ANDN U11196 ( .B(n8615), .A(n12633), .Z(n8616) );
  NANDN U11197 ( .A(n8616), .B(n12635), .Z(n8617) );
  ANDN U11198 ( .B(n8617), .A(n12637), .Z(n8618) );
  NANDN U11199 ( .A(n8618), .B(n12639), .Z(n8619) );
  NANDN U11200 ( .A(n12641), .B(n8619), .Z(n8620) );
  NAND U11201 ( .A(n8620), .B(n12643), .Z(n8622) );
  NANDN U11202 ( .A(n8622), .B(n8621), .Z(n8623) );
  AND U11203 ( .A(n8624), .B(n8623), .Z(n8627) );
  AND U11204 ( .A(n12651), .B(n8625), .Z(n8626) );
  NANDN U11205 ( .A(n8627), .B(n8626), .Z(n8630) );
  NAND U11206 ( .A(n8629), .B(n8628), .Z(n12653) );
  ANDN U11207 ( .B(n8630), .A(n12653), .Z(n8633) );
  NAND U11208 ( .A(n8632), .B(n8631), .Z(n12656) );
  OR U11209 ( .A(n8633), .B(n12656), .Z(n8636) );
  NANDN U11210 ( .A(y[1392]), .B(x[1392]), .Z(n8635) );
  NAND U11211 ( .A(n8635), .B(n8634), .Z(n12657) );
  ANDN U11212 ( .B(n8636), .A(n12657), .Z(n8637) );
  NANDN U11213 ( .A(n8637), .B(n12659), .Z(n8638) );
  ANDN U11214 ( .B(n8638), .A(n12661), .Z(n8639) );
  NANDN U11215 ( .A(n8639), .B(n12663), .Z(n8640) );
  ANDN U11216 ( .B(n8640), .A(n12665), .Z(n8641) );
  OR U11217 ( .A(n12667), .B(n8641), .Z(n8644) );
  NANDN U11218 ( .A(y[1398]), .B(x[1398]), .Z(n8643) );
  ANDN U11219 ( .B(n8643), .A(n8642), .Z(n12670) );
  NAND U11220 ( .A(n8644), .B(n12670), .Z(n8646) );
  ANDN U11221 ( .B(n8646), .A(n8645), .Z(n8647) );
  NAND U11222 ( .A(n8647), .B(n12671), .Z(n8648) );
  AND U11223 ( .A(n12677), .B(n8648), .Z(n8649) );
  NAND U11224 ( .A(n8649), .B(n12673), .Z(n8651) );
  ANDN U11225 ( .B(n8651), .A(n8650), .Z(n8652) );
  NAND U11226 ( .A(n8652), .B(n12679), .Z(n8655) );
  NOR U11227 ( .A(n8654), .B(n8653), .Z(n12682) );
  NAND U11228 ( .A(n8655), .B(n12682), .Z(n8658) );
  NANDN U11229 ( .A(x[1404]), .B(y[1404]), .Z(n8656) );
  NAND U11230 ( .A(n8657), .B(n8656), .Z(n12684) );
  ANDN U11231 ( .B(n8658), .A(n12684), .Z(n8659) );
  OR U11232 ( .A(n12686), .B(n8659), .Z(n8660) );
  ANDN U11233 ( .B(n8660), .A(n12688), .Z(n8661) );
  OR U11234 ( .A(n12689), .B(n8661), .Z(n8662) );
  NANDN U11235 ( .A(n12692), .B(n8662), .Z(n8663) );
  NAND U11236 ( .A(n8663), .B(n12694), .Z(n8665) );
  ANDN U11237 ( .B(n8665), .A(n8664), .Z(n8666) );
  NAND U11238 ( .A(n8666), .B(n12695), .Z(n8669) );
  AND U11239 ( .A(n8668), .B(n8667), .Z(n12697) );
  NAND U11240 ( .A(n8669), .B(n12697), .Z(n8671) );
  ANDN U11241 ( .B(n8671), .A(n8670), .Z(n8672) );
  NAND U11242 ( .A(n8672), .B(n12699), .Z(n8673) );
  NANDN U11243 ( .A(n12705), .B(n8673), .Z(n8676) );
  NANDN U11244 ( .A(x[1415]), .B(y[1415]), .Z(n8675) );
  ANDN U11245 ( .B(n8675), .A(n8674), .Z(n12707) );
  NAND U11246 ( .A(n8676), .B(n12707), .Z(n8681) );
  NANDN U11247 ( .A(n8678), .B(n8677), .Z(n8679) );
  NAND U11248 ( .A(n8680), .B(n8679), .Z(n12710) );
  ANDN U11249 ( .B(n8681), .A(n12710), .Z(n8684) );
  NANDN U11250 ( .A(x[1417]), .B(y[1417]), .Z(n8683) );
  ANDN U11251 ( .B(n8683), .A(n8682), .Z(n12711) );
  NANDN U11252 ( .A(n8684), .B(n12711), .Z(n8685) );
  NANDN U11253 ( .A(n12714), .B(n8685), .Z(n8686) );
  NAND U11254 ( .A(n8686), .B(n12716), .Z(n8687) );
  NAND U11255 ( .A(n8687), .B(n12717), .Z(n8688) );
  ANDN U11256 ( .B(n8688), .A(n12719), .Z(n8695) );
  OR U11257 ( .A(n8690), .B(n8689), .Z(n8691) );
  AND U11258 ( .A(n8692), .B(n8691), .Z(n8694) );
  AND U11259 ( .A(n8694), .B(n8693), .Z(n12721) );
  NANDN U11260 ( .A(n8695), .B(n12721), .Z(n8696) );
  NANDN U11261 ( .A(n12724), .B(n8696), .Z(n8699) );
  ANDN U11262 ( .B(n8698), .A(n8697), .Z(n12726) );
  NAND U11263 ( .A(n8699), .B(n12726), .Z(n8700) );
  NANDN U11264 ( .A(n12728), .B(n8700), .Z(n8703) );
  NANDN U11265 ( .A(y[1428]), .B(x[1428]), .Z(n8702) );
  NAND U11266 ( .A(n8702), .B(n8701), .Z(n12730) );
  ANDN U11267 ( .B(n8703), .A(n12730), .Z(n8704) );
  NANDN U11268 ( .A(n8704), .B(n12731), .Z(n8705) );
  NANDN U11269 ( .A(n12733), .B(n8705), .Z(n8706) );
  NAND U11270 ( .A(n8706), .B(n12735), .Z(n8708) );
  NANDN U11271 ( .A(n8708), .B(n8707), .Z(n8709) );
  ANDN U11272 ( .B(n8709), .A(n12738), .Z(n8711) );
  NANDN U11273 ( .A(n8711), .B(n8710), .Z(n8714) );
  ANDN U11274 ( .B(n8713), .A(n8712), .Z(n12741) );
  NAND U11275 ( .A(n8714), .B(n12741), .Z(n8715) );
  NAND U11276 ( .A(n8715), .B(n12744), .Z(n8717) );
  NANDN U11277 ( .A(n8717), .B(n8716), .Z(n8718) );
  AND U11278 ( .A(n8719), .B(n8718), .Z(n8722) );
  ANDN U11279 ( .B(n12751), .A(n8720), .Z(n8721) );
  NANDN U11280 ( .A(n8722), .B(n8721), .Z(n8729) );
  NAND U11281 ( .A(n8724), .B(n8723), .Z(n8725) );
  NANDN U11282 ( .A(n8726), .B(n8725), .Z(n8727) );
  NANDN U11283 ( .A(n8728), .B(n8727), .Z(n12754) );
  ANDN U11284 ( .B(n8729), .A(n12754), .Z(n8731) );
  NANDN U11285 ( .A(n8731), .B(n8730), .Z(n8732) );
  NANDN U11286 ( .A(n12758), .B(n8732), .Z(n8734) );
  NAND U11287 ( .A(n8734), .B(n8733), .Z(n8735) );
  ANDN U11288 ( .B(n8735), .A(n12766), .Z(n8738) );
  ANDN U11289 ( .B(n12767), .A(n8736), .Z(n8737) );
  NANDN U11290 ( .A(n8738), .B(n8737), .Z(n8739) );
  NANDN U11291 ( .A(n12777), .B(n8739), .Z(n8741) );
  IV U11292 ( .A(n8740), .Z(n12778) );
  ANDN U11293 ( .B(n8741), .A(n12778), .Z(n8742) );
  NANDN U11294 ( .A(n8743), .B(n8742), .Z(n8744) );
  NAND U11295 ( .A(n8744), .B(n12783), .Z(n8745) );
  NANDN U11296 ( .A(n8745), .B(n12775), .Z(n8746) );
  AND U11297 ( .A(n8747), .B(n8746), .Z(n8750) );
  NOR U11298 ( .A(n8749), .B(n8748), .Z(n12787) );
  NANDN U11299 ( .A(n8750), .B(n12787), .Z(n8751) );
  NANDN U11300 ( .A(n12790), .B(n8751), .Z(n8752) );
  NAND U11301 ( .A(n8752), .B(n12792), .Z(n8753) );
  NAND U11302 ( .A(n8753), .B(n12793), .Z(n8754) );
  NAND U11303 ( .A(n8754), .B(n12795), .Z(n8755) );
  ANDN U11304 ( .B(n8755), .A(n12798), .Z(n8756) );
  NANDN U11305 ( .A(n8756), .B(n12800), .Z(n8759) );
  NOR U11306 ( .A(n8758), .B(n8757), .Z(n12801) );
  NAND U11307 ( .A(n8759), .B(n12801), .Z(n8762) );
  ANDN U11308 ( .B(n8761), .A(n8760), .Z(n12804) );
  NAND U11309 ( .A(n8762), .B(n12804), .Z(n8763) );
  ANDN U11310 ( .B(n8763), .A(n12806), .Z(n8764) );
  NANDN U11311 ( .A(n8765), .B(n8764), .Z(n8766) );
  NAND U11312 ( .A(n8766), .B(n12811), .Z(n8767) );
  NANDN U11313 ( .A(n8767), .B(n12807), .Z(n8768) );
  AND U11314 ( .A(n12813), .B(n8768), .Z(n8769) );
  NANDN U11315 ( .A(n8770), .B(n8769), .Z(n8772) );
  NAND U11316 ( .A(n8772), .B(n12816), .Z(n8777) );
  NANDN U11317 ( .A(n8774), .B(n8773), .Z(n8775) );
  NAND U11318 ( .A(n8776), .B(n8775), .Z(n12818) );
  ANDN U11319 ( .B(n8777), .A(n12818), .Z(n8780) );
  NANDN U11320 ( .A(y[1464]), .B(x[1464]), .Z(n8779) );
  ANDN U11321 ( .B(n8779), .A(n8778), .Z(n12819) );
  NANDN U11322 ( .A(n8780), .B(n12819), .Z(n8781) );
  NANDN U11323 ( .A(n12822), .B(n8781), .Z(n8782) );
  NAND U11324 ( .A(n8782), .B(n12823), .Z(n8783) );
  NANDN U11325 ( .A(n12826), .B(n8783), .Z(n8784) );
  NAND U11326 ( .A(n8784), .B(n12828), .Z(n8785) );
  ANDN U11327 ( .B(n8785), .A(n12830), .Z(n8786) );
  OR U11328 ( .A(n12831), .B(n8786), .Z(n8787) );
  NAND U11329 ( .A(n8787), .B(n12833), .Z(n8788) );
  ANDN U11330 ( .B(n8788), .A(n12836), .Z(n8789) );
  OR U11331 ( .A(n12838), .B(n8789), .Z(n8790) );
  NANDN U11332 ( .A(n12840), .B(n8790), .Z(n8791) );
  NAND U11333 ( .A(n8791), .B(n12841), .Z(n8792) );
  NANDN U11334 ( .A(n12843), .B(n8792), .Z(n8793) );
  NAND U11335 ( .A(n8793), .B(n12845), .Z(n8794) );
  ANDN U11336 ( .B(n8794), .A(n12848), .Z(n8795) );
  NANDN U11337 ( .A(n8795), .B(n12849), .Z(n8802) );
  AND U11338 ( .A(n8797), .B(n8796), .Z(n8801) );
  NANDN U11339 ( .A(n8799), .B(n8798), .Z(n8800) );
  NAND U11340 ( .A(n8801), .B(n8800), .Z(n12852) );
  ANDN U11341 ( .B(n8802), .A(n12852), .Z(n8803) );
  OR U11342 ( .A(n12854), .B(n8803), .Z(n8804) );
  NANDN U11343 ( .A(n12856), .B(n8804), .Z(n8807) );
  NANDN U11344 ( .A(x[1487]), .B(y[1487]), .Z(n8806) );
  NAND U11345 ( .A(n8806), .B(n8805), .Z(n12858) );
  ANDN U11346 ( .B(n8807), .A(n12858), .Z(n8808) );
  NANDN U11347 ( .A(n8808), .B(n12859), .Z(n8809) );
  ANDN U11348 ( .B(n8809), .A(n12861), .Z(n8810) );
  NANDN U11349 ( .A(n8810), .B(n12863), .Z(n8811) );
  NANDN U11350 ( .A(n12866), .B(n8811), .Z(n8814) );
  NOR U11351 ( .A(n8813), .B(n8812), .Z(n12867) );
  NAND U11352 ( .A(n8814), .B(n12867), .Z(n8816) );
  ANDN U11353 ( .B(n8816), .A(n8815), .Z(n8817) );
  NAND U11354 ( .A(n8817), .B(n12869), .Z(n8818) );
  NANDN U11355 ( .A(n8819), .B(n8818), .Z(n8821) );
  ANDN U11356 ( .B(n8821), .A(n8820), .Z(n8822) );
  NAND U11357 ( .A(n8822), .B(n12877), .Z(n8825) );
  NOR U11358 ( .A(n8824), .B(n8823), .Z(n12880) );
  NAND U11359 ( .A(n8825), .B(n12880), .Z(n8826) );
  NANDN U11360 ( .A(n12882), .B(n8826), .Z(n8827) );
  NANDN U11361 ( .A(n12884), .B(n8827), .Z(n8828) );
  ANDN U11362 ( .B(n8828), .A(n12886), .Z(n8829) );
  NANDN U11363 ( .A(n8829), .B(n12887), .Z(n8830) );
  ANDN U11364 ( .B(n8830), .A(n12890), .Z(n8831) );
  NANDN U11365 ( .A(n8831), .B(n12891), .Z(n8832) );
  NANDN U11366 ( .A(n8833), .B(n8832), .Z(n8835) );
  NAND U11367 ( .A(n8835), .B(n8834), .Z(n8837) );
  ANDN U11368 ( .B(n8837), .A(n8836), .Z(n8838) );
  NANDN U11369 ( .A(n8839), .B(n8838), .Z(n8840) );
  NAND U11370 ( .A(n8840), .B(n12899), .Z(n8842) );
  NANDN U11371 ( .A(n8842), .B(n8841), .Z(n8844) );
  ANDN U11372 ( .B(n8844), .A(n8843), .Z(n8845) );
  ANDN U11373 ( .B(n8845), .A(n12902), .Z(n8852) );
  NAND U11374 ( .A(n8847), .B(n8846), .Z(n8848) );
  NANDN U11375 ( .A(n8849), .B(n8848), .Z(n8851) );
  ANDN U11376 ( .B(n8851), .A(n8850), .Z(n12903) );
  NANDN U11377 ( .A(n8852), .B(n12903), .Z(n8853) );
  NANDN U11378 ( .A(n12905), .B(n8853), .Z(n8854) );
  NAND U11379 ( .A(n8854), .B(n12907), .Z(n8855) );
  NAND U11380 ( .A(n8856), .B(n8855), .Z(n8857) );
  AND U11381 ( .A(n12911), .B(n8857), .Z(n8858) );
  OR U11382 ( .A(n8859), .B(n8858), .Z(n8860) );
  NANDN U11383 ( .A(n8861), .B(n8860), .Z(n8863) );
  NAND U11384 ( .A(n8863), .B(n8862), .Z(n8865) );
  NANDN U11385 ( .A(n8865), .B(n8864), .Z(n8867) );
  AND U11386 ( .A(n12917), .B(n12922), .Z(n8866) );
  NAND U11387 ( .A(n8867), .B(n8866), .Z(n8868) );
  NAND U11388 ( .A(n8868), .B(n12923), .Z(n8870) );
  NANDN U11389 ( .A(n8870), .B(n8869), .Z(n8877) );
  NANDN U11390 ( .A(n8872), .B(n8871), .Z(n8873) );
  NANDN U11391 ( .A(n8874), .B(n8873), .Z(n8876) );
  NAND U11392 ( .A(n8876), .B(n8875), .Z(n12926) );
  ANDN U11393 ( .B(n8877), .A(n12926), .Z(n8878) );
  NANDN U11394 ( .A(n8878), .B(n12927), .Z(n8879) );
  NANDN U11395 ( .A(n12930), .B(n8879), .Z(n8880) );
  AND U11396 ( .A(n12931), .B(n8880), .Z(n8881) );
  NANDN U11397 ( .A(n8881), .B(n12933), .Z(n8882) );
  NANDN U11398 ( .A(n12936), .B(n8882), .Z(n8885) );
  NANDN U11399 ( .A(y[1530]), .B(x[1530]), .Z(n8884) );
  ANDN U11400 ( .B(n8884), .A(n8883), .Z(n12937) );
  NAND U11401 ( .A(n8885), .B(n12937), .Z(n8887) );
  ANDN U11402 ( .B(n8887), .A(n8886), .Z(n8888) );
  NAND U11403 ( .A(n8888), .B(n12940), .Z(n8889) );
  NANDN U11404 ( .A(n8890), .B(n8889), .Z(n8891) );
  AND U11405 ( .A(n12948), .B(n8891), .Z(n8892) );
  NANDN U11406 ( .A(n8893), .B(n8892), .Z(n8896) );
  NOR U11407 ( .A(n8895), .B(n8894), .Z(n12949) );
  NAND U11408 ( .A(n8896), .B(n12949), .Z(n8897) );
  NANDN U11409 ( .A(n12951), .B(n8897), .Z(n8898) );
  NAND U11410 ( .A(n8898), .B(n12953), .Z(n8899) );
  ANDN U11411 ( .B(n8899), .A(n12956), .Z(n8900) );
  NANDN U11412 ( .A(n8900), .B(n12957), .Z(n8901) );
  ANDN U11413 ( .B(n8901), .A(n12960), .Z(n8902) );
  NANDN U11414 ( .A(n8902), .B(n12961), .Z(n8903) );
  NANDN U11415 ( .A(n12964), .B(n8903), .Z(n8906) );
  NOR U11416 ( .A(n8905), .B(n8904), .Z(n12965) );
  NAND U11417 ( .A(n8906), .B(n12965), .Z(n8907) );
  AND U11418 ( .A(n12967), .B(n8907), .Z(n8909) );
  NAND U11419 ( .A(n8909), .B(n8908), .Z(n8912) );
  AND U11420 ( .A(n8910), .B(n12970), .Z(n8911) );
  NAND U11421 ( .A(n8912), .B(n8911), .Z(n8913) );
  NANDN U11422 ( .A(n12977), .B(n8913), .Z(n8916) );
  NANDN U11423 ( .A(y[1546]), .B(x[1546]), .Z(n8915) );
  ANDN U11424 ( .B(n8915), .A(n8914), .Z(n12978) );
  NAND U11425 ( .A(n8916), .B(n12978), .Z(n8919) );
  NAND U11426 ( .A(n8918), .B(n8917), .Z(n12980) );
  ANDN U11427 ( .B(n8919), .A(n12980), .Z(n8922) );
  NANDN U11428 ( .A(y[1548]), .B(x[1548]), .Z(n8921) );
  ANDN U11429 ( .B(n8921), .A(n8920), .Z(n12982) );
  NANDN U11430 ( .A(n8922), .B(n12982), .Z(n8923) );
  NANDN U11431 ( .A(n12985), .B(n8923), .Z(n8926) );
  NANDN U11432 ( .A(y[1550]), .B(x[1550]), .Z(n8925) );
  ANDN U11433 ( .B(n8925), .A(n8924), .Z(n12987) );
  NAND U11434 ( .A(n8926), .B(n12987), .Z(n8928) );
  NAND U11435 ( .A(n8928), .B(n8927), .Z(n8930) );
  NAND U11436 ( .A(n8930), .B(n8929), .Z(n8931) );
  NAND U11437 ( .A(n8931), .B(n12994), .Z(n8934) );
  NAND U11438 ( .A(n8933), .B(n8932), .Z(n12997) );
  ANDN U11439 ( .B(n8934), .A(n12997), .Z(n8937) );
  ANDN U11440 ( .B(n12998), .A(n8935), .Z(n8936) );
  NANDN U11441 ( .A(n8937), .B(n8936), .Z(n8938) );
  NANDN U11442 ( .A(n8939), .B(n8938), .Z(n8941) );
  ANDN U11443 ( .B(n8941), .A(n8940), .Z(n8942) );
  NANDN U11444 ( .A(n13007), .B(n8942), .Z(n8945) );
  NANDN U11445 ( .A(y[1559]), .B(x[1559]), .Z(n8944) );
  ANDN U11446 ( .B(n8944), .A(n8943), .Z(n13009) );
  NAND U11447 ( .A(n8945), .B(n13009), .Z(n8946) );
  NANDN U11448 ( .A(n13011), .B(n8946), .Z(n8949) );
  NANDN U11449 ( .A(y[1560]), .B(x[1560]), .Z(n8948) );
  NAND U11450 ( .A(n8948), .B(n8947), .Z(n13012) );
  ANDN U11451 ( .B(n8949), .A(n13012), .Z(n8950) );
  ANDN U11452 ( .B(n8951), .A(n8950), .Z(n8952) );
  NAND U11453 ( .A(n8952), .B(n13014), .Z(n8954) );
  NAND U11454 ( .A(n8954), .B(n8953), .Z(n8956) );
  ANDN U11455 ( .B(n8956), .A(n8955), .Z(n8957) );
  NANDN U11456 ( .A(n13022), .B(n8957), .Z(n8958) );
  NANDN U11457 ( .A(n8959), .B(n8958), .Z(n8960) );
  AND U11458 ( .A(n13026), .B(n8960), .Z(n8963) );
  NOR U11459 ( .A(n8962), .B(n8961), .Z(n13028) );
  NANDN U11460 ( .A(n8963), .B(n13028), .Z(n8964) );
  AND U11461 ( .A(n13030), .B(n8964), .Z(n8965) );
  NANDN U11462 ( .A(n8966), .B(n8965), .Z(n8967) );
  AND U11463 ( .A(n13036), .B(n8967), .Z(n8968) );
  NAND U11464 ( .A(n8968), .B(n13032), .Z(n8970) );
  ANDN U11465 ( .B(n8970), .A(n8969), .Z(n8971) );
  NAND U11466 ( .A(n8971), .B(n13038), .Z(n8974) );
  ANDN U11467 ( .B(n8973), .A(n8972), .Z(n13040) );
  NAND U11468 ( .A(n8974), .B(n13040), .Z(n8975) );
  NANDN U11469 ( .A(n13042), .B(n8975), .Z(n8976) );
  NANDN U11470 ( .A(n13045), .B(n8976), .Z(n8979) );
  NANDN U11471 ( .A(x[1573]), .B(y[1573]), .Z(n8978) );
  NAND U11472 ( .A(n8978), .B(n8977), .Z(n13047) );
  ANDN U11473 ( .B(n8979), .A(n13047), .Z(n8980) );
  NANDN U11474 ( .A(n8980), .B(n13048), .Z(n8981) );
  ANDN U11475 ( .B(n8981), .A(n13050), .Z(n8982) );
  NANDN U11476 ( .A(n8982), .B(n13052), .Z(n8983) );
  NANDN U11477 ( .A(n13055), .B(n8983), .Z(n8986) );
  ANDN U11478 ( .B(n8985), .A(n8984), .Z(n13056) );
  NAND U11479 ( .A(n8986), .B(n13056), .Z(n8988) );
  ANDN U11480 ( .B(n8988), .A(n8987), .Z(n8989) );
  NAND U11481 ( .A(n8989), .B(n13058), .Z(n8990) );
  NANDN U11482 ( .A(n8991), .B(n8990), .Z(n8992) );
  NAND U11483 ( .A(n8993), .B(n8992), .Z(n8998) );
  NANDN U11484 ( .A(n8995), .B(n8994), .Z(n8996) );
  NAND U11485 ( .A(n8997), .B(n8996), .Z(n13069) );
  ANDN U11486 ( .B(n8998), .A(n13069), .Z(n9001) );
  NANDN U11487 ( .A(x[1583]), .B(y[1583]), .Z(n9000) );
  ANDN U11488 ( .B(n9000), .A(n8999), .Z(n13070) );
  NANDN U11489 ( .A(n9001), .B(n13070), .Z(n9002) );
  NANDN U11490 ( .A(n13073), .B(n9002), .Z(n9005) );
  NANDN U11491 ( .A(x[1585]), .B(y[1585]), .Z(n9004) );
  ANDN U11492 ( .B(n9004), .A(n9003), .Z(n13075) );
  NAND U11493 ( .A(n9005), .B(n13075), .Z(n9006) );
  NANDN U11494 ( .A(n13077), .B(n9006), .Z(n9007) );
  NAND U11495 ( .A(n9007), .B(n13078), .Z(n9008) );
  NAND U11496 ( .A(n9008), .B(n13081), .Z(n9009) );
  NANDN U11497 ( .A(n13083), .B(n9009), .Z(n9010) );
  NAND U11498 ( .A(n9010), .B(n13085), .Z(n9011) );
  ANDN U11499 ( .B(n9011), .A(n13087), .Z(n9012) );
  OR U11500 ( .A(n13089), .B(n9012), .Z(n9013) );
  NANDN U11501 ( .A(n13091), .B(n9013), .Z(n9014) );
  NAND U11502 ( .A(n9014), .B(n13092), .Z(n9015) );
  NANDN U11503 ( .A(n13095), .B(n9015), .Z(n9022) );
  NANDN U11504 ( .A(n9017), .B(n9016), .Z(n9018) );
  NANDN U11505 ( .A(n9019), .B(n9018), .Z(n9021) );
  ANDN U11506 ( .B(n9021), .A(n9020), .Z(n13097) );
  NAND U11507 ( .A(n9022), .B(n13097), .Z(n9023) );
  ANDN U11508 ( .B(n9023), .A(n13099), .Z(n9024) );
  NANDN U11509 ( .A(n9024), .B(n13100), .Z(n9026) );
  NAND U11510 ( .A(n9026), .B(n9025), .Z(n9028) );
  NAND U11511 ( .A(n9028), .B(n9027), .Z(n9029) );
  NANDN U11512 ( .A(n13111), .B(n9029), .Z(n9030) );
  NANDN U11513 ( .A(n13112), .B(n9030), .Z(n9031) );
  NAND U11514 ( .A(n9031), .B(n13114), .Z(n9032) );
  NANDN U11515 ( .A(n13117), .B(n9032), .Z(n9033) );
  NANDN U11516 ( .A(n13119), .B(n9033), .Z(n9034) );
  NAND U11517 ( .A(n9034), .B(n13121), .Z(n9035) );
  NANDN U11518 ( .A(n13123), .B(n9035), .Z(n9036) );
  NANDN U11519 ( .A(n13125), .B(n9036), .Z(n9037) );
  AND U11520 ( .A(n13126), .B(n9037), .Z(n9039) );
  NAND U11521 ( .A(n9039), .B(n9038), .Z(n9040) );
  AND U11522 ( .A(n13132), .B(n9040), .Z(n9041) );
  NAND U11523 ( .A(n9041), .B(n13128), .Z(n9042) );
  ANDN U11524 ( .B(n9042), .A(n13135), .Z(n9044) );
  NAND U11525 ( .A(n9044), .B(n9043), .Z(n9047) );
  NOR U11526 ( .A(n9046), .B(n9045), .Z(n13136) );
  NAND U11527 ( .A(n9047), .B(n13136), .Z(n9048) );
  AND U11528 ( .A(n13139), .B(n9048), .Z(n9050) );
  NAND U11529 ( .A(n9050), .B(n9049), .Z(n9051) );
  NAND U11530 ( .A(n9051), .B(n13140), .Z(n9052) );
  NANDN U11531 ( .A(n9052), .B(n13145), .Z(n9053) );
  NAND U11532 ( .A(n9054), .B(n9053), .Z(n9055) );
  NANDN U11533 ( .A(n9056), .B(n9055), .Z(n9057) );
  NANDN U11534 ( .A(n13153), .B(n9057), .Z(n9058) );
  NANDN U11535 ( .A(n13154), .B(n9058), .Z(n9061) );
  NANDN U11536 ( .A(x[1619]), .B(y[1619]), .Z(n9060) );
  NANDN U11537 ( .A(x[1620]), .B(y[1620]), .Z(n9059) );
  NAND U11538 ( .A(n9060), .B(n9059), .Z(n13157) );
  ANDN U11539 ( .B(n9061), .A(n13157), .Z(n9062) );
  OR U11540 ( .A(n13159), .B(n9062), .Z(n9065) );
  NANDN U11541 ( .A(x[1621]), .B(y[1621]), .Z(n9064) );
  ANDN U11542 ( .B(n9064), .A(n9063), .Z(n13160) );
  NAND U11543 ( .A(n9065), .B(n13160), .Z(n9066) );
  NANDN U11544 ( .A(n13163), .B(n9066), .Z(n9067) );
  NANDN U11545 ( .A(n9068), .B(n9067), .Z(n9070) );
  ANDN U11546 ( .B(n9070), .A(n9069), .Z(n9071) );
  OR U11547 ( .A(n9072), .B(n9071), .Z(n9073) );
  NAND U11548 ( .A(n9073), .B(n13176), .Z(n9074) );
  NAND U11549 ( .A(n9074), .B(n13178), .Z(n9075) );
  NANDN U11550 ( .A(n13181), .B(n9075), .Z(n9076) );
  NAND U11551 ( .A(n9076), .B(n13182), .Z(n9077) );
  ANDN U11552 ( .B(n9077), .A(n13185), .Z(n9080) );
  ANDN U11553 ( .B(n9078), .A(n13187), .Z(n9079) );
  NANDN U11554 ( .A(n9080), .B(n9079), .Z(n9081) );
  AND U11555 ( .A(n13188), .B(n9081), .Z(n9084) );
  NOR U11556 ( .A(n9083), .B(n9082), .Z(n13192) );
  NANDN U11557 ( .A(n9084), .B(n13192), .Z(n9087) );
  ANDN U11558 ( .B(n9086), .A(n9085), .Z(n13195) );
  ANDN U11559 ( .B(n9087), .A(n13195), .Z(n9089) );
  NAND U11560 ( .A(n9089), .B(n9088), .Z(n9090) );
  ANDN U11561 ( .B(n9090), .A(n13197), .Z(n9092) );
  NANDN U11562 ( .A(n9092), .B(n9091), .Z(n9093) );
  ANDN U11563 ( .B(n9093), .A(n13201), .Z(n9094) );
  NANDN U11564 ( .A(n9094), .B(n13203), .Z(n9095) );
  NAND U11565 ( .A(n9095), .B(n13204), .Z(n9096) );
  NAND U11566 ( .A(n9096), .B(n13206), .Z(n9101) );
  NANDN U11567 ( .A(n9098), .B(n9097), .Z(n9100) );
  ANDN U11568 ( .B(n9100), .A(n9099), .Z(n13208) );
  NAND U11569 ( .A(n9101), .B(n13208), .Z(n9104) );
  NANDN U11570 ( .A(y[1642]), .B(x[1642]), .Z(n9103) );
  ANDN U11571 ( .B(n9103), .A(n9102), .Z(n13210) );
  NAND U11572 ( .A(n9104), .B(n13210), .Z(n9105) );
  AND U11573 ( .A(n13212), .B(n9105), .Z(n9106) );
  NANDN U11574 ( .A(n9107), .B(n9106), .Z(n9108) );
  ANDN U11575 ( .B(n9108), .A(n13214), .Z(n9109) );
  NAND U11576 ( .A(n9110), .B(n9109), .Z(n9111) );
  NAND U11577 ( .A(n9112), .B(n9111), .Z(n9113) );
  AND U11578 ( .A(n13222), .B(n9113), .Z(n9115) );
  NAND U11579 ( .A(n9115), .B(n9114), .Z(n9116) );
  NAND U11580 ( .A(n9116), .B(n13225), .Z(n9118) );
  NANDN U11581 ( .A(n9118), .B(n9117), .Z(n9119) );
  AND U11582 ( .A(n13226), .B(n9119), .Z(n9120) );
  OR U11583 ( .A(n13229), .B(n9120), .Z(n9121) );
  NAND U11584 ( .A(n9122), .B(n9121), .Z(n9123) );
  NAND U11585 ( .A(n9123), .B(n13232), .Z(n9124) );
  NAND U11586 ( .A(n9125), .B(n9124), .Z(n9126) );
  NAND U11587 ( .A(n9127), .B(n9126), .Z(n9128) );
  NAND U11588 ( .A(n9129), .B(n9128), .Z(n9130) );
  NAND U11589 ( .A(n9131), .B(n9130), .Z(n9133) );
  ANDN U11590 ( .B(n9133), .A(n9132), .Z(n9134) );
  NANDN U11591 ( .A(n9134), .B(n13241), .Z(n9135) );
  ANDN U11592 ( .B(n9135), .A(n13243), .Z(n9136) );
  NANDN U11593 ( .A(n9136), .B(n13244), .Z(n9137) );
  NAND U11594 ( .A(n9137), .B(n13248), .Z(n9138) );
  NAND U11595 ( .A(n9138), .B(n13250), .Z(n9139) );
  NANDN U11596 ( .A(n9140), .B(n9139), .Z(n9141) );
  ANDN U11597 ( .B(n9141), .A(n13255), .Z(n9142) );
  NANDN U11598 ( .A(n9142), .B(n13257), .Z(n9143) );
  NAND U11599 ( .A(n9143), .B(n13258), .Z(n9146) );
  NOR U11600 ( .A(n9145), .B(n9144), .Z(n13260) );
  NAND U11601 ( .A(n9146), .B(n13260), .Z(n9147) );
  NANDN U11602 ( .A(n9148), .B(n9147), .Z(n9150) );
  ANDN U11603 ( .B(n9150), .A(n9149), .Z(n9152) );
  OR U11604 ( .A(n9152), .B(n9151), .Z(n9153) );
  NAND U11605 ( .A(n9154), .B(n9153), .Z(n9155) );
  NAND U11606 ( .A(n9156), .B(n9155), .Z(n9157) );
  NAND U11607 ( .A(n9158), .B(n9157), .Z(n9159) );
  NAND U11608 ( .A(n9160), .B(n9159), .Z(n9161) );
  ANDN U11609 ( .B(n9161), .A(n13273), .Z(n9163) );
  NAND U11610 ( .A(n9163), .B(n9162), .Z(n9164) );
  NANDN U11611 ( .A(n13275), .B(n9164), .Z(n9166) );
  NANDN U11612 ( .A(n9166), .B(n9165), .Z(n9167) );
  AND U11613 ( .A(n13276), .B(n9167), .Z(n9168) );
  NAND U11614 ( .A(n9169), .B(n9168), .Z(n9170) );
  AND U11615 ( .A(n9171), .B(n9170), .Z(n9174) );
  AND U11616 ( .A(n13285), .B(n9172), .Z(n9173) );
  NANDN U11617 ( .A(n9174), .B(n9173), .Z(n9175) );
  AND U11618 ( .A(n13286), .B(n9175), .Z(n9176) );
  NANDN U11619 ( .A(n9177), .B(n9176), .Z(n9180) );
  ANDN U11620 ( .B(n9179), .A(n9178), .Z(n13289) );
  NAND U11621 ( .A(n9180), .B(n13289), .Z(n9181) );
  AND U11622 ( .A(n13290), .B(n9181), .Z(n9183) );
  NANDN U11623 ( .A(n9183), .B(n9182), .Z(n9184) );
  AND U11624 ( .A(n13295), .B(n9184), .Z(n9185) );
  NANDN U11625 ( .A(n9186), .B(n9185), .Z(n9187) );
  AND U11626 ( .A(n9188), .B(n9187), .Z(n9189) );
  NAND U11627 ( .A(n9189), .B(n13297), .Z(n9191) );
  ANDN U11628 ( .B(n9191), .A(n9190), .Z(n9192) );
  NAND U11629 ( .A(n9193), .B(n9192), .Z(n9194) );
  NAND U11630 ( .A(n9195), .B(n9194), .Z(n9197) );
  ANDN U11631 ( .B(n9197), .A(n9196), .Z(n9198) );
  NAND U11632 ( .A(n9199), .B(n9198), .Z(n9200) );
  NAND U11633 ( .A(n9201), .B(n9200), .Z(n9203) );
  ANDN U11634 ( .B(n9203), .A(n9202), .Z(n9204) );
  NAND U11635 ( .A(n9205), .B(n9204), .Z(n9206) );
  NAND U11636 ( .A(n9207), .B(n9206), .Z(n9208) );
  AND U11637 ( .A(n9209), .B(n9208), .Z(n9210) );
  NAND U11638 ( .A(n9211), .B(n9210), .Z(n9212) );
  NAND U11639 ( .A(n9213), .B(n9212), .Z(n9215) );
  AND U11640 ( .A(n9215), .B(n9214), .Z(n9216) );
  NANDN U11641 ( .A(n13321), .B(n9216), .Z(n9217) );
  NANDN U11642 ( .A(n13323), .B(n9217), .Z(n9220) );
  NANDN U11643 ( .A(x[1691]), .B(y[1691]), .Z(n9219) );
  ANDN U11644 ( .B(n9219), .A(n9218), .Z(n13325) );
  NAND U11645 ( .A(n9220), .B(n13325), .Z(n9222) );
  ANDN U11646 ( .B(n9222), .A(n9221), .Z(n9223) );
  NAND U11647 ( .A(n9223), .B(n13326), .Z(n9224) );
  AND U11648 ( .A(n9225), .B(n9224), .Z(n9226) );
  NAND U11649 ( .A(n9226), .B(n13328), .Z(n9228) );
  ANDN U11650 ( .B(n9228), .A(n9227), .Z(n9229) );
  NAND U11651 ( .A(n9230), .B(n9229), .Z(n9231) );
  NAND U11652 ( .A(n9232), .B(n9231), .Z(n9234) );
  AND U11653 ( .A(n9234), .B(n9233), .Z(n9235) );
  NANDN U11654 ( .A(n9236), .B(n9235), .Z(n9239) );
  ANDN U11655 ( .B(n9238), .A(n9237), .Z(n13342) );
  NAND U11656 ( .A(n9239), .B(n13342), .Z(n9240) );
  ANDN U11657 ( .B(n9240), .A(n13343), .Z(n9242) );
  NAND U11658 ( .A(n9242), .B(n9241), .Z(n9243) );
  NAND U11659 ( .A(n9243), .B(n13340), .Z(n9244) );
  NAND U11660 ( .A(n9245), .B(n9244), .Z(n9247) );
  NANDN U11661 ( .A(x[1700]), .B(y[1700]), .Z(n9246) );
  AND U11662 ( .A(n9247), .B(n9246), .Z(n9248) );
  NAND U11663 ( .A(n9249), .B(n9248), .Z(n9250) );
  NAND U11664 ( .A(n9251), .B(n9250), .Z(n9252) );
  NAND U11665 ( .A(n9253), .B(n9252), .Z(n9254) );
  NAND U11666 ( .A(n9255), .B(n9254), .Z(n9257) );
  ANDN U11667 ( .B(n9257), .A(n9256), .Z(n9258) );
  NANDN U11668 ( .A(n9259), .B(n9258), .Z(n9262) );
  NOR U11669 ( .A(n9261), .B(n9260), .Z(n9993) );
  NAND U11670 ( .A(n9262), .B(n9993), .Z(n9263) );
  NAND U11671 ( .A(n9264), .B(n9263), .Z(n9265) );
  NANDN U11672 ( .A(n13358), .B(n9265), .Z(n9267) );
  OR U11673 ( .A(n9267), .B(n9266), .Z(n9270) );
  XNOR U11674 ( .A(n9267), .B(y[1707]), .Z(n9268) );
  NANDN U11675 ( .A(x[1707]), .B(n9268), .Z(n9269) );
  NAND U11676 ( .A(n9270), .B(n9269), .Z(n9271) );
  NANDN U11677 ( .A(n9271), .B(n13367), .Z(n9272) );
  AND U11678 ( .A(n13370), .B(n9272), .Z(n9274) );
  NAND U11679 ( .A(n9274), .B(n9273), .Z(n9276) );
  ANDN U11680 ( .B(n9276), .A(n9275), .Z(n9277) );
  NANDN U11681 ( .A(n9277), .B(n13375), .Z(n9278) );
  ANDN U11682 ( .B(n9278), .A(n13377), .Z(n9279) );
  NANDN U11683 ( .A(n9279), .B(n13379), .Z(n9280) );
  ANDN U11684 ( .B(n9280), .A(n13381), .Z(n9281) );
  OR U11685 ( .A(n9282), .B(n9281), .Z(n9283) );
  NAND U11686 ( .A(n9283), .B(n13384), .Z(n9284) );
  AND U11687 ( .A(n13388), .B(n9284), .Z(n9285) );
  NANDN U11688 ( .A(n9285), .B(n13390), .Z(n9286) );
  AND U11689 ( .A(n13392), .B(n9286), .Z(n9287) );
  NANDN U11690 ( .A(n9287), .B(n13394), .Z(n9288) );
  NANDN U11691 ( .A(n13397), .B(n9288), .Z(n9291) );
  NANDN U11692 ( .A(x[1719]), .B(y[1719]), .Z(n9290) );
  NAND U11693 ( .A(n9290), .B(n9289), .Z(n13398) );
  ANDN U11694 ( .B(n9291), .A(n13398), .Z(n9294) );
  AND U11695 ( .A(n13400), .B(n9292), .Z(n9293) );
  NANDN U11696 ( .A(n9294), .B(n9293), .Z(n9295) );
  AND U11697 ( .A(n13402), .B(n9295), .Z(n9297) );
  OR U11698 ( .A(n9297), .B(n9296), .Z(n9298) );
  ANDN U11699 ( .B(n9298), .A(n13407), .Z(n9299) );
  OR U11700 ( .A(n13409), .B(n9299), .Z(n9300) );
  AND U11701 ( .A(n9301), .B(n9300), .Z(n9302) );
  OR U11702 ( .A(n9302), .B(x[1725]), .Z(n9306) );
  XOR U11703 ( .A(x[1725]), .B(n9302), .Z(n9303) );
  NANDN U11704 ( .A(n9304), .B(n9303), .Z(n9305) );
  NAND U11705 ( .A(n9306), .B(n9305), .Z(n9308) );
  ANDN U11706 ( .B(n9308), .A(n9307), .Z(n9309) );
  NANDN U11707 ( .A(n9309), .B(n13414), .Z(n9310) );
  ANDN U11708 ( .B(n9310), .A(n13417), .Z(n9311) );
  NANDN U11709 ( .A(n9311), .B(n13418), .Z(n9312) );
  NANDN U11710 ( .A(n9313), .B(n9312), .Z(n9314) );
  NAND U11711 ( .A(n9314), .B(n13422), .Z(n9315) );
  NAND U11712 ( .A(n9316), .B(n9315), .Z(n9317) );
  NANDN U11713 ( .A(n13424), .B(n9317), .Z(n9318) );
  NANDN U11714 ( .A(n13425), .B(n9318), .Z(n9321) );
  NANDN U11715 ( .A(x[1733]), .B(y[1733]), .Z(n9320) );
  NAND U11716 ( .A(n9320), .B(n9319), .Z(n13426) );
  ANDN U11717 ( .B(n9321), .A(n13426), .Z(n9324) );
  AND U11718 ( .A(n13427), .B(n9322), .Z(n9323) );
  NANDN U11719 ( .A(n9324), .B(n9323), .Z(n9325) );
  NAND U11720 ( .A(n9325), .B(n13428), .Z(n9326) );
  NANDN U11721 ( .A(n9326), .B(x[1736]), .Z(n9329) );
  XNOR U11722 ( .A(n9326), .B(x[1736]), .Z(n9327) );
  NANDN U11723 ( .A(y[1736]), .B(n9327), .Z(n9328) );
  AND U11724 ( .A(n9329), .B(n9328), .Z(n9330) );
  OR U11725 ( .A(n9330), .B(y[1737]), .Z(n9333) );
  XOR U11726 ( .A(y[1737]), .B(n9330), .Z(n9331) );
  NAND U11727 ( .A(n9331), .B(x[1737]), .Z(n9332) );
  NAND U11728 ( .A(n9333), .B(n9332), .Z(n9334) );
  AND U11729 ( .A(n13432), .B(n9334), .Z(n9338) );
  ANDN U11730 ( .B(n9336), .A(n9335), .Z(n9337) );
  NANDN U11731 ( .A(n9338), .B(n9337), .Z(n9339) );
  AND U11732 ( .A(n9340), .B(n9339), .Z(n9341) );
  NAND U11733 ( .A(n9342), .B(n9341), .Z(n9343) );
  NAND U11734 ( .A(n9344), .B(n9343), .Z(n9346) );
  ANDN U11735 ( .B(n9346), .A(n9345), .Z(n9347) );
  NANDN U11736 ( .A(n9347), .B(n13435), .Z(n9348) );
  ANDN U11737 ( .B(n9348), .A(n13436), .Z(n9349) );
  OR U11738 ( .A(n13437), .B(n9349), .Z(n9350) );
  NAND U11739 ( .A(n9350), .B(n13439), .Z(n9351) );
  AND U11740 ( .A(n13440), .B(n9351), .Z(n9352) );
  NANDN U11741 ( .A(n9352), .B(n13442), .Z(n9355) );
  NAND U11742 ( .A(n9354), .B(n9353), .Z(n13445) );
  ANDN U11743 ( .B(n9355), .A(n13445), .Z(n9356) );
  OR U11744 ( .A(n13447), .B(n9356), .Z(n9357) );
  NAND U11745 ( .A(n9358), .B(n9357), .Z(n9359) );
  NAND U11746 ( .A(n9360), .B(n9359), .Z(n9362) );
  ANDN U11747 ( .B(n9362), .A(n9361), .Z(n9363) );
  NAND U11748 ( .A(n9363), .B(n13459), .Z(n9365) );
  NAND U11749 ( .A(n9365), .B(n9364), .Z(n9368) );
  ANDN U11750 ( .B(n9367), .A(n9366), .Z(n13458) );
  NAND U11751 ( .A(n9368), .B(n13458), .Z(n9369) );
  NANDN U11752 ( .A(n13463), .B(n9369), .Z(n9372) );
  NANDN U11753 ( .A(y[1754]), .B(x[1754]), .Z(n9371) );
  ANDN U11754 ( .B(n9371), .A(n9370), .Z(n13469) );
  NAND U11755 ( .A(n9372), .B(n13469), .Z(n9373) );
  AND U11756 ( .A(n13470), .B(n9373), .Z(n9374) );
  NANDN U11757 ( .A(n9375), .B(n9374), .Z(n9376) );
  AND U11758 ( .A(n13472), .B(n9376), .Z(n9377) );
  NAND U11759 ( .A(n9378), .B(n9377), .Z(n9379) );
  NAND U11760 ( .A(n9380), .B(n9379), .Z(n9381) );
  AND U11761 ( .A(n13480), .B(n9381), .Z(n9382) );
  NANDN U11762 ( .A(n9383), .B(n9382), .Z(n9384) );
  NAND U11763 ( .A(n9384), .B(n13482), .Z(n9386) );
  NANDN U11764 ( .A(n9386), .B(n9385), .Z(n9387) );
  AND U11765 ( .A(n13484), .B(n9387), .Z(n9388) );
  OR U11766 ( .A(n13487), .B(n9388), .Z(n9389) );
  NAND U11767 ( .A(n9390), .B(n9389), .Z(n9391) );
  NAND U11768 ( .A(n9392), .B(n9391), .Z(n9393) );
  NAND U11769 ( .A(n9394), .B(n9393), .Z(n9396) );
  OR U11770 ( .A(n9396), .B(n9395), .Z(n9399) );
  XNOR U11771 ( .A(n9396), .B(y[1765]), .Z(n9397) );
  NANDN U11772 ( .A(x[1765]), .B(n9397), .Z(n9398) );
  AND U11773 ( .A(n9399), .B(n9398), .Z(n9402) );
  NANDN U11774 ( .A(y[1766]), .B(n9402), .Z(n9400) );
  AND U11775 ( .A(n9401), .B(n9400), .Z(n9405) );
  XNOR U11776 ( .A(n9402), .B(y[1766]), .Z(n9403) );
  NAND U11777 ( .A(n9403), .B(x[1766]), .Z(n9404) );
  NAND U11778 ( .A(n9405), .B(n9404), .Z(n9407) );
  ANDN U11779 ( .B(n9407), .A(n9406), .Z(n9408) );
  NAND U11780 ( .A(n9409), .B(n9408), .Z(n9410) );
  NAND U11781 ( .A(n9411), .B(n9410), .Z(n9413) );
  ANDN U11782 ( .B(n9413), .A(n9412), .Z(n9414) );
  NAND U11783 ( .A(n9415), .B(n9414), .Z(n9416) );
  NAND U11784 ( .A(n9417), .B(n9416), .Z(n9419) );
  ANDN U11785 ( .B(n9419), .A(n9418), .Z(n9420) );
  NAND U11786 ( .A(n9421), .B(n9420), .Z(n9422) );
  NAND U11787 ( .A(n9423), .B(n9422), .Z(n9426) );
  OR U11788 ( .A(n9425), .B(n9424), .Z(n13515) );
  ANDN U11789 ( .B(n9426), .A(n13515), .Z(n9427) );
  NANDN U11790 ( .A(n9428), .B(n9427), .Z(n9441) );
  ANDN U11791 ( .B(n9430), .A(n9429), .Z(n9438) );
  NANDN U11792 ( .A(n9432), .B(n9431), .Z(n9434) );
  ANDN U11793 ( .B(n9434), .A(n9433), .Z(n9436) );
  XNOR U11794 ( .A(y[1776]), .B(x[1776]), .Z(n9435) );
  NANDN U11795 ( .A(n9436), .B(n9435), .Z(n9437) );
  NAND U11796 ( .A(n9438), .B(n9437), .Z(n9440) );
  AND U11797 ( .A(n9440), .B(n9439), .Z(n13517) );
  NAND U11798 ( .A(n9441), .B(n13517), .Z(n9442) );
  NAND U11799 ( .A(n9442), .B(n13518), .Z(n9443) );
  ANDN U11800 ( .B(n9443), .A(n13521), .Z(n9444) );
  NANDN U11801 ( .A(n9444), .B(n13522), .Z(n9445) );
  NAND U11802 ( .A(n9445), .B(n13524), .Z(n9446) );
  AND U11803 ( .A(n13526), .B(n9446), .Z(n9449) );
  ANDN U11804 ( .B(n9447), .A(n13528), .Z(n9448) );
  NANDN U11805 ( .A(n9449), .B(n9448), .Z(n9450) );
  NANDN U11806 ( .A(n13531), .B(n9450), .Z(n9452) );
  OR U11807 ( .A(n9452), .B(n9451), .Z(n9455) );
  XNOR U11808 ( .A(n9452), .B(x[1784]), .Z(n9453) );
  NANDN U11809 ( .A(y[1784]), .B(n9453), .Z(n9454) );
  AND U11810 ( .A(n9455), .B(n9454), .Z(n9458) );
  OR U11811 ( .A(n9458), .B(y[1785]), .Z(n9456) );
  AND U11812 ( .A(n9457), .B(n9456), .Z(n9461) );
  XOR U11813 ( .A(n9458), .B(y[1785]), .Z(n9459) );
  NAND U11814 ( .A(n9459), .B(x[1785]), .Z(n9460) );
  NAND U11815 ( .A(n9461), .B(n9460), .Z(n9462) );
  NANDN U11816 ( .A(n13539), .B(n9462), .Z(n9463) );
  NAND U11817 ( .A(n9463), .B(n13541), .Z(n9464) );
  ANDN U11818 ( .B(n9464), .A(n13543), .Z(n9468) );
  OR U11819 ( .A(y[1789]), .B(n9465), .Z(n9467) );
  ANDN U11820 ( .B(n9467), .A(n9466), .Z(n13544) );
  NANDN U11821 ( .A(n9468), .B(n13544), .Z(n9469) );
  NANDN U11822 ( .A(n13547), .B(n9469), .Z(n9471) );
  NAND U11823 ( .A(n9471), .B(n13548), .Z(n9472) );
  NANDN U11824 ( .A(n13551), .B(n9472), .Z(n9473) );
  NAND U11825 ( .A(n9473), .B(n13553), .Z(n9474) );
  ANDN U11826 ( .B(n9474), .A(n13555), .Z(n9476) );
  NANDN U11827 ( .A(n9476), .B(n9475), .Z(n9477) );
  NANDN U11828 ( .A(n9478), .B(n9477), .Z(n9480) );
  NAND U11829 ( .A(n9480), .B(n9479), .Z(n9481) );
  AND U11830 ( .A(n13562), .B(n9481), .Z(n9482) );
  NANDN U11831 ( .A(n9483), .B(n9482), .Z(n9484) );
  NAND U11832 ( .A(n9484), .B(n13564), .Z(n9485) );
  NANDN U11833 ( .A(n9485), .B(n9991), .Z(n9486) );
  AND U11834 ( .A(n13565), .B(n9486), .Z(n9488) );
  NAND U11835 ( .A(n9488), .B(n9487), .Z(n9491) );
  NAND U11836 ( .A(n9490), .B(n9489), .Z(n13566) );
  ANDN U11837 ( .B(n9491), .A(n13566), .Z(n9494) );
  AND U11838 ( .A(n13567), .B(n9492), .Z(n9493) );
  NANDN U11839 ( .A(n9494), .B(n9493), .Z(n9495) );
  AND U11840 ( .A(n13568), .B(n9495), .Z(n9496) );
  NAND U11841 ( .A(n9497), .B(n9496), .Z(n9498) );
  NAND U11842 ( .A(n9499), .B(n9498), .Z(n9500) );
  AND U11843 ( .A(n9501), .B(n9500), .Z(n9502) );
  NAND U11844 ( .A(n9503), .B(n9502), .Z(n9504) );
  NAND U11845 ( .A(n9505), .B(n9504), .Z(n9507) );
  AND U11846 ( .A(n9507), .B(n9506), .Z(n9508) );
  NAND U11847 ( .A(n9508), .B(n13576), .Z(n9509) );
  NANDN U11848 ( .A(n13579), .B(n9509), .Z(n9510) );
  ANDN U11849 ( .B(n9510), .A(n13581), .Z(n9512) );
  NAND U11850 ( .A(n9512), .B(n9511), .Z(n9513) );
  NAND U11851 ( .A(n9513), .B(n13582), .Z(n9514) );
  NAND U11852 ( .A(n9515), .B(n9514), .Z(n9517) );
  NANDN U11853 ( .A(x[1812]), .B(y[1812]), .Z(n9516) );
  AND U11854 ( .A(n9517), .B(n9516), .Z(n9518) );
  NAND U11855 ( .A(n9519), .B(n9518), .Z(n9520) );
  NAND U11856 ( .A(n9521), .B(n9520), .Z(n9522) );
  NAND U11857 ( .A(n9523), .B(n9522), .Z(n9524) );
  NAND U11858 ( .A(n9525), .B(n9524), .Z(n9527) );
  ANDN U11859 ( .B(n9527), .A(n9526), .Z(n9528) );
  NAND U11860 ( .A(n9528), .B(n13594), .Z(n9529) );
  NAND U11861 ( .A(n9529), .B(n13597), .Z(n9532) );
  ANDN U11862 ( .B(n9531), .A(n9530), .Z(n13598) );
  NAND U11863 ( .A(n9532), .B(n13598), .Z(n9533) );
  AND U11864 ( .A(n9534), .B(n9533), .Z(n9535) );
  NAND U11865 ( .A(n9535), .B(n13601), .Z(n9536) );
  NAND U11866 ( .A(n9536), .B(n13602), .Z(n9538) );
  OR U11867 ( .A(n9538), .B(n9537), .Z(n9541) );
  XNOR U11868 ( .A(n9538), .B(x[1820]), .Z(n9539) );
  NANDN U11869 ( .A(y[1820]), .B(n9539), .Z(n9540) );
  AND U11870 ( .A(n9541), .B(n9540), .Z(n9544) );
  OR U11871 ( .A(n9544), .B(y[1821]), .Z(n9542) );
  AND U11872 ( .A(n9543), .B(n9542), .Z(n9547) );
  XOR U11873 ( .A(y[1821]), .B(n9544), .Z(n9545) );
  NAND U11874 ( .A(n9545), .B(x[1821]), .Z(n9546) );
  NAND U11875 ( .A(n9547), .B(n9546), .Z(n9548) );
  NAND U11876 ( .A(n9548), .B(n13610), .Z(n9550) );
  NAND U11877 ( .A(n9550), .B(n9549), .Z(n9551) );
  AND U11878 ( .A(n9552), .B(n9551), .Z(n9553) );
  NANDN U11879 ( .A(n9554), .B(n9553), .Z(n9555) );
  AND U11880 ( .A(n13622), .B(n9555), .Z(n9556) );
  NAND U11881 ( .A(n9556), .B(n13617), .Z(n9557) );
  AND U11882 ( .A(n13624), .B(n9557), .Z(n9558) );
  NANDN U11883 ( .A(n9559), .B(n9558), .Z(n9560) );
  NANDN U11884 ( .A(n9561), .B(n9560), .Z(n9562) );
  NANDN U11885 ( .A(n13629), .B(n9562), .Z(n9563) );
  NANDN U11886 ( .A(n13631), .B(n9563), .Z(n9564) );
  NAND U11887 ( .A(n9564), .B(n13633), .Z(n9567) );
  NANDN U11888 ( .A(y[1831]), .B(x[1831]), .Z(n9566) );
  ANDN U11889 ( .B(n9566), .A(n9565), .Z(n13634) );
  NAND U11890 ( .A(n9567), .B(n13634), .Z(n9570) );
  ANDN U11891 ( .B(n9569), .A(n9568), .Z(n13636) );
  NAND U11892 ( .A(n9570), .B(n13636), .Z(n9571) );
  AND U11893 ( .A(n13638), .B(n9571), .Z(n9572) );
  NANDN U11894 ( .A(n9573), .B(n9572), .Z(n9574) );
  AND U11895 ( .A(n9575), .B(n9574), .Z(n9576) );
  NAND U11896 ( .A(n9576), .B(n13640), .Z(n9578) );
  ANDN U11897 ( .B(n9578), .A(n9577), .Z(n9579) );
  NAND U11898 ( .A(n9580), .B(n9579), .Z(n9581) );
  NAND U11899 ( .A(n9582), .B(n9581), .Z(n9584) );
  ANDN U11900 ( .B(n9584), .A(n9583), .Z(n9585) );
  NAND U11901 ( .A(n9586), .B(n9585), .Z(n9587) );
  NAND U11902 ( .A(n9588), .B(n9587), .Z(n9590) );
  ANDN U11903 ( .B(n9590), .A(n9589), .Z(n9591) );
  NAND U11904 ( .A(n9591), .B(n13656), .Z(n9593) );
  NAND U11905 ( .A(n9593), .B(n9592), .Z(n9594) );
  NANDN U11906 ( .A(n9594), .B(n9989), .Z(n9596) );
  NAND U11907 ( .A(n9596), .B(n9595), .Z(n9597) );
  AND U11908 ( .A(n9988), .B(n9597), .Z(n9598) );
  NANDN U11909 ( .A(n9599), .B(n9598), .Z(n9600) );
  AND U11910 ( .A(n13667), .B(n9600), .Z(n9601) );
  NAND U11911 ( .A(n9601), .B(n13661), .Z(n9602) );
  AND U11912 ( .A(n13668), .B(n9602), .Z(n9603) );
  NANDN U11913 ( .A(n9604), .B(n9603), .Z(n9607) );
  NOR U11914 ( .A(n9606), .B(n9605), .Z(n13671) );
  NAND U11915 ( .A(n9607), .B(n13671), .Z(n9608) );
  NANDN U11916 ( .A(n9609), .B(n9608), .Z(n9611) );
  NAND U11917 ( .A(n9611), .B(n9610), .Z(n9613) );
  ANDN U11918 ( .B(n9613), .A(n9612), .Z(n9614) );
  NAND U11919 ( .A(n9614), .B(n13678), .Z(n9615) );
  AND U11920 ( .A(n9616), .B(n9615), .Z(n9617) );
  NAND U11921 ( .A(n9617), .B(n13682), .Z(n9618) );
  AND U11922 ( .A(n13689), .B(n9618), .Z(n9619) );
  NANDN U11923 ( .A(n9620), .B(n9619), .Z(n9622) );
  NAND U11924 ( .A(n9622), .B(n9621), .Z(n9624) );
  NANDN U11925 ( .A(n9624), .B(n9623), .Z(n9625) );
  AND U11926 ( .A(n9626), .B(n9625), .Z(n9627) );
  NANDN U11927 ( .A(n9628), .B(n9627), .Z(n9629) );
  AND U11928 ( .A(n9630), .B(n9629), .Z(n9632) );
  NAND U11929 ( .A(n9632), .B(n9631), .Z(n9634) );
  ANDN U11930 ( .B(n9634), .A(n9633), .Z(n9635) );
  NAND U11931 ( .A(n9636), .B(n9635), .Z(n9637) );
  NAND U11932 ( .A(n9638), .B(n9637), .Z(n9640) );
  ANDN U11933 ( .B(n9640), .A(n9639), .Z(n9641) );
  NANDN U11934 ( .A(n9641), .B(n13700), .Z(n9642) );
  ANDN U11935 ( .B(n9642), .A(n13703), .Z(n9643) );
  NANDN U11936 ( .A(n9643), .B(n13704), .Z(n9644) );
  NANDN U11937 ( .A(n13707), .B(n9644), .Z(n9645) );
  NANDN U11938 ( .A(n13709), .B(n9645), .Z(n9646) );
  NANDN U11939 ( .A(n13710), .B(n9646), .Z(n9647) );
  NAND U11940 ( .A(n9647), .B(n13712), .Z(n9648) );
  AND U11941 ( .A(n13714), .B(n9648), .Z(n9649) );
  NANDN U11942 ( .A(n9649), .B(n13716), .Z(n9650) );
  NANDN U11943 ( .A(n13719), .B(n9650), .Z(n9651) );
  NAND U11944 ( .A(n9651), .B(n13720), .Z(n9652) );
  NANDN U11945 ( .A(n13722), .B(n9652), .Z(n9653) );
  NAND U11946 ( .A(n9653), .B(n13724), .Z(n9654) );
  ANDN U11947 ( .B(n9654), .A(n13727), .Z(n9655) );
  NANDN U11948 ( .A(n9655), .B(n13730), .Z(n9657) );
  NAND U11949 ( .A(y[1868]), .B(n9656), .Z(n9986) );
  NAND U11950 ( .A(n9657), .B(n9986), .Z(n9658) );
  NANDN U11951 ( .A(n13729), .B(n9658), .Z(n9660) );
  NANDN U11952 ( .A(n9660), .B(n9659), .Z(n9661) );
  NAND U11953 ( .A(n9662), .B(n9661), .Z(n9663) );
  NANDN U11954 ( .A(n9664), .B(n9663), .Z(n9666) );
  NAND U11955 ( .A(n9666), .B(n9665), .Z(n9667) );
  ANDN U11956 ( .B(n9667), .A(n13739), .Z(n9668) );
  OR U11957 ( .A(n13741), .B(n9668), .Z(n9669) );
  NAND U11958 ( .A(n9670), .B(n9669), .Z(n9671) );
  NAND U11959 ( .A(n9671), .B(n13745), .Z(n9672) );
  NAND U11960 ( .A(n9673), .B(n9672), .Z(n9674) );
  NAND U11961 ( .A(n9675), .B(n9674), .Z(n9676) );
  NAND U11962 ( .A(n9677), .B(n9676), .Z(n9678) );
  NAND U11963 ( .A(n9679), .B(n9678), .Z(n9681) );
  ANDN U11964 ( .B(n9681), .A(n9680), .Z(n9682) );
  NANDN U11965 ( .A(n9683), .B(n9682), .Z(n9684) );
  NAND U11966 ( .A(n9685), .B(n9684), .Z(n9686) );
  NANDN U11967 ( .A(n9686), .B(n13761), .Z(n9687) );
  NANDN U11968 ( .A(n9688), .B(n9687), .Z(n9689) );
  NAND U11969 ( .A(n9689), .B(n13765), .Z(n9690) );
  NANDN U11970 ( .A(n13767), .B(n9690), .Z(n9691) );
  NAND U11971 ( .A(n9691), .B(n13769), .Z(n9692) );
  AND U11972 ( .A(n13770), .B(n9692), .Z(n9693) );
  NANDN U11973 ( .A(n9693), .B(n13772), .Z(n9699) );
  ANDN U11974 ( .B(n9699), .A(n13774), .Z(n9702) );
  AND U11975 ( .A(n13776), .B(n9700), .Z(n9701) );
  NANDN U11976 ( .A(n9702), .B(n9701), .Z(n9703) );
  ANDN U11977 ( .B(n9703), .A(n13779), .Z(n9704) );
  NAND U11978 ( .A(n9705), .B(n9704), .Z(n9706) );
  NAND U11979 ( .A(n9707), .B(n9706), .Z(n9708) );
  ANDN U11980 ( .B(n9708), .A(n13786), .Z(n9710) );
  NAND U11981 ( .A(n9710), .B(n9709), .Z(n9711) );
  NANDN U11982 ( .A(n13788), .B(n9711), .Z(n9712) );
  ANDN U11983 ( .B(n9712), .A(n13791), .Z(n9713) );
  NANDN U11984 ( .A(n9713), .B(n13793), .Z(n9714) );
  NANDN U11985 ( .A(n13795), .B(n9714), .Z(n9715) );
  NAND U11986 ( .A(n9715), .B(n13797), .Z(n9716) );
  NAND U11987 ( .A(n9716), .B(n13798), .Z(n9717) );
  NAND U11988 ( .A(n9717), .B(n13800), .Z(n9718) );
  AND U11989 ( .A(n13802), .B(n9718), .Z(n9719) );
  OR U11990 ( .A(n13805), .B(n9719), .Z(n9720) );
  NANDN U11991 ( .A(n13806), .B(n9720), .Z(n9721) );
  NANDN U11992 ( .A(n13808), .B(n9721), .Z(n9722) );
  NANDN U11993 ( .A(n13809), .B(n9722), .Z(n9723) );
  NAND U11994 ( .A(n9723), .B(n13810), .Z(n9724) );
  ANDN U11995 ( .B(n9724), .A(n13811), .Z(n9725) );
  NANDN U11996 ( .A(n9725), .B(n13812), .Z(n9726) );
  ANDN U11997 ( .B(n9726), .A(n13813), .Z(n9727) );
  NANDN U11998 ( .A(n9727), .B(n13814), .Z(n9728) );
  ANDN U11999 ( .B(n9728), .A(n13815), .Z(n9729) );
  NANDN U12000 ( .A(n9729), .B(n13816), .Z(n9730) );
  NANDN U12001 ( .A(n13817), .B(n9730), .Z(n9731) );
  NANDN U12002 ( .A(n13818), .B(n9731), .Z(n9734) );
  NOR U12003 ( .A(n9733), .B(n9732), .Z(n13819) );
  ANDN U12004 ( .B(n9734), .A(n13819), .Z(n9735) );
  NANDN U12005 ( .A(n9736), .B(n9735), .Z(n9738) );
  NAND U12006 ( .A(n9738), .B(n9737), .Z(n9740) );
  ANDN U12007 ( .B(n9740), .A(n9739), .Z(n9741) );
  NAND U12008 ( .A(n9742), .B(n9741), .Z(n9743) );
  NAND U12009 ( .A(n9744), .B(n9743), .Z(n9745) );
  ANDN U12010 ( .B(n9745), .A(n13823), .Z(n9746) );
  NANDN U12011 ( .A(n9747), .B(n9746), .Z(n9748) );
  NANDN U12012 ( .A(n9749), .B(n9748), .Z(n9750) );
  NANDN U12013 ( .A(n13827), .B(n9750), .Z(n9753) );
  NANDN U12014 ( .A(x[1922]), .B(y[1922]), .Z(n9752) );
  ANDN U12015 ( .B(n9752), .A(n9751), .Z(n13829) );
  NAND U12016 ( .A(n9753), .B(n13829), .Z(n9756) );
  NANDN U12017 ( .A(y[1922]), .B(x[1922]), .Z(n9754) );
  NAND U12018 ( .A(n9755), .B(n9754), .Z(n13830) );
  ANDN U12019 ( .B(n9756), .A(n13830), .Z(n9757) );
  NANDN U12020 ( .A(n9757), .B(n13832), .Z(n9758) );
  ANDN U12021 ( .B(n9758), .A(n13835), .Z(n9759) );
  NANDN U12022 ( .A(n9759), .B(n13837), .Z(n9760) );
  NAND U12023 ( .A(n9760), .B(n13838), .Z(n9761) );
  NAND U12024 ( .A(n9761), .B(n13840), .Z(n9762) );
  AND U12025 ( .A(n13842), .B(n9762), .Z(n9763) );
  NANDN U12026 ( .A(n9763), .B(n13844), .Z(n9766) );
  NOR U12027 ( .A(n9765), .B(n9764), .Z(n13846) );
  NAND U12028 ( .A(n9766), .B(n13846), .Z(n9768) );
  NAND U12029 ( .A(n9768), .B(n9767), .Z(n9769) );
  NANDN U12030 ( .A(n13851), .B(n9769), .Z(n9771) );
  NAND U12031 ( .A(n9771), .B(n9770), .Z(n9772) );
  ANDN U12032 ( .B(n9772), .A(n13855), .Z(n9773) );
  NANDN U12033 ( .A(n9773), .B(n13857), .Z(n9774) );
  ANDN U12034 ( .B(n9774), .A(n13859), .Z(n9775) );
  NANDN U12035 ( .A(n9775), .B(n13861), .Z(n9776) );
  ANDN U12036 ( .B(n9776), .A(n13863), .Z(n9777) );
  OR U12037 ( .A(n13865), .B(n9777), .Z(n9778) );
  NAND U12038 ( .A(n9778), .B(n13866), .Z(n9779) );
  ANDN U12039 ( .B(n9779), .A(n13868), .Z(n9781) );
  NANDN U12040 ( .A(n9781), .B(n9780), .Z(n9782) );
  AND U12041 ( .A(n13873), .B(n9782), .Z(n9787) );
  NANDN U12042 ( .A(n9784), .B(n9783), .Z(n9785) );
  ANDN U12043 ( .B(n9785), .A(n13875), .Z(n9786) );
  NANDN U12044 ( .A(n9787), .B(n9786), .Z(n9788) );
  NANDN U12045 ( .A(n13877), .B(n9788), .Z(n9789) );
  NAND U12046 ( .A(n9789), .B(n13878), .Z(n9790) );
  ANDN U12047 ( .B(n9790), .A(n13880), .Z(n9791) );
  NANDN U12048 ( .A(n9791), .B(n13882), .Z(n9792) );
  NANDN U12049 ( .A(n13885), .B(n9792), .Z(n9793) );
  NAND U12050 ( .A(n9793), .B(n13886), .Z(n9794) );
  NAND U12051 ( .A(n9794), .B(n13888), .Z(n9795) );
  ANDN U12052 ( .B(n9795), .A(n13891), .Z(n9797) );
  NAND U12053 ( .A(n9797), .B(n9796), .Z(n9798) );
  AND U12054 ( .A(n13893), .B(n9798), .Z(n9799) );
  OR U12055 ( .A(n9800), .B(n9799), .Z(n9801) );
  NANDN U12056 ( .A(n13902), .B(n9801), .Z(n9803) );
  NAND U12057 ( .A(n9803), .B(n9802), .Z(n9804) );
  NANDN U12058 ( .A(y[1954]), .B(n9804), .Z(n9807) );
  XNOR U12059 ( .A(y[1954]), .B(n9804), .Z(n9805) );
  NAND U12060 ( .A(n9805), .B(x[1954]), .Z(n9806) );
  NAND U12061 ( .A(n9807), .B(n9806), .Z(n9808) );
  AND U12062 ( .A(n9809), .B(n9808), .Z(n9810) );
  NANDN U12063 ( .A(n9810), .B(n13905), .Z(n9811) );
  NANDN U12064 ( .A(n9812), .B(n9811), .Z(n9814) );
  ANDN U12065 ( .B(n9814), .A(n9813), .Z(n9816) );
  NANDN U12066 ( .A(n9816), .B(n9815), .Z(n9817) );
  NANDN U12067 ( .A(n9818), .B(n9817), .Z(n9819) );
  NAND U12068 ( .A(n9819), .B(n13914), .Z(n9820) );
  NANDN U12069 ( .A(n13915), .B(n9820), .Z(n9821) );
  NAND U12070 ( .A(n9821), .B(n13916), .Z(n9822) );
  ANDN U12071 ( .B(n9822), .A(n13917), .Z(n9823) );
  NANDN U12072 ( .A(n9823), .B(n13918), .Z(n9824) );
  ANDN U12073 ( .B(n9824), .A(n13919), .Z(n9825) );
  NANDN U12074 ( .A(n9825), .B(n13920), .Z(n9826) );
  NAND U12075 ( .A(n9826), .B(n13923), .Z(n9827) );
  NAND U12076 ( .A(n9827), .B(n13924), .Z(n9832) );
  NANDN U12077 ( .A(n9829), .B(n9828), .Z(n9830) );
  NAND U12078 ( .A(n9831), .B(n9830), .Z(n13927) );
  ANDN U12079 ( .B(n9832), .A(n13927), .Z(n9835) );
  NANDN U12080 ( .A(x[1971]), .B(y[1971]), .Z(n9834) );
  ANDN U12081 ( .B(n9834), .A(n9833), .Z(n13928) );
  NANDN U12082 ( .A(n9835), .B(n13928), .Z(n9836) );
  NAND U12083 ( .A(n9836), .B(n13930), .Z(n9837) );
  ANDN U12084 ( .B(n9837), .A(n13933), .Z(n9839) );
  NANDN U12085 ( .A(n9839), .B(n9838), .Z(n9840) );
  NANDN U12086 ( .A(n9841), .B(n9840), .Z(n9842) );
  NAND U12087 ( .A(n9842), .B(n13941), .Z(n9843) );
  NANDN U12088 ( .A(n9844), .B(n9843), .Z(n9846) );
  NAND U12089 ( .A(n9846), .B(n9845), .Z(n9848) );
  ANDN U12090 ( .B(n9848), .A(n9847), .Z(n9850) );
  ANDN U12091 ( .B(n9850), .A(n9849), .Z(n9851) );
  ANDN U12092 ( .B(n9852), .A(n9851), .Z(n9853) );
  OR U12093 ( .A(n9853), .B(y[1981]), .Z(n9856) );
  XOR U12094 ( .A(y[1981]), .B(n9853), .Z(n9854) );
  NAND U12095 ( .A(n9854), .B(x[1981]), .Z(n9855) );
  NAND U12096 ( .A(n9856), .B(n9855), .Z(n9858) );
  ANDN U12097 ( .B(n9858), .A(n9857), .Z(n9861) );
  AND U12098 ( .A(n13952), .B(n9859), .Z(n9860) );
  NANDN U12099 ( .A(n9861), .B(n9860), .Z(n9863) );
  ANDN U12100 ( .B(n9863), .A(n9862), .Z(n9864) );
  AND U12101 ( .A(n13954), .B(n9864), .Z(n9867) );
  ANDN U12102 ( .B(n9866), .A(n9865), .Z(n13957) );
  NANDN U12103 ( .A(n9867), .B(n13957), .Z(n9868) );
  NANDN U12104 ( .A(n13958), .B(n9868), .Z(n9869) );
  NAND U12105 ( .A(n9869), .B(n13959), .Z(n9870) );
  AND U12106 ( .A(n13960), .B(n9870), .Z(n9871) );
  NANDN U12107 ( .A(n9871), .B(n13961), .Z(n9872) );
  NANDN U12108 ( .A(n13962), .B(n9872), .Z(n9873) );
  NAND U12109 ( .A(n9873), .B(n9978), .Z(n9874) );
  AND U12110 ( .A(n13963), .B(n9874), .Z(n9876) );
  NANDN U12111 ( .A(n9876), .B(n9875), .Z(n9877) );
  NANDN U12112 ( .A(n13965), .B(n9877), .Z(n9878) );
  AND U12113 ( .A(n13966), .B(n9878), .Z(n9880) );
  ANDN U12114 ( .B(n9880), .A(n9879), .Z(n9881) );
  ANDN U12115 ( .B(n13967), .A(n9881), .Z(n9882) );
  NAND U12116 ( .A(n9883), .B(n9882), .Z(n9884) );
  NAND U12117 ( .A(n9885), .B(n9884), .Z(n9887) );
  AND U12118 ( .A(n9887), .B(n9886), .Z(n9889) );
  NAND U12119 ( .A(n9889), .B(n9888), .Z(n9890) );
  NAND U12120 ( .A(n9890), .B(n13972), .Z(n9892) );
  NANDN U12121 ( .A(n9892), .B(n9891), .Z(n9893) );
  AND U12122 ( .A(n13973), .B(n9893), .Z(n9895) );
  NAND U12123 ( .A(n9895), .B(n9894), .Z(n9896) );
  AND U12124 ( .A(n13974), .B(n9896), .Z(n9897) );
  OR U12125 ( .A(n13977), .B(n9897), .Z(n9898) );
  NANDN U12126 ( .A(n13979), .B(n9898), .Z(n9899) );
  NAND U12127 ( .A(n9899), .B(n13981), .Z(n9900) );
  ANDN U12128 ( .B(n9900), .A(n13983), .Z(n9901) );
  NAND U12129 ( .A(n9901), .B(n13986), .Z(n9902) );
  NANDN U12130 ( .A(n13988), .B(n9902), .Z(n9903) );
  NAND U12131 ( .A(n9903), .B(n13990), .Z(n9904) );
  ANDN U12132 ( .B(n9904), .A(n13992), .Z(n9905) );
  OR U12133 ( .A(n9906), .B(n9905), .Z(n9907) );
  NANDN U12134 ( .A(y[2010]), .B(n9907), .Z(n9910) );
  XNOR U12135 ( .A(y[2010]), .B(n9907), .Z(n9908) );
  NAND U12136 ( .A(n9908), .B(x[2010]), .Z(n9909) );
  NAND U12137 ( .A(n9910), .B(n9909), .Z(n9912) );
  ANDN U12138 ( .B(n9912), .A(n9911), .Z(n9913) );
  NANDN U12139 ( .A(n9913), .B(n13998), .Z(n9914) );
  NANDN U12140 ( .A(n14000), .B(n9914), .Z(n9915) );
  NAND U12141 ( .A(n9916), .B(n9915), .Z(n9917) );
  NAND U12142 ( .A(n9917), .B(n14009), .Z(n9918) );
  NANDN U12143 ( .A(n14011), .B(n9918), .Z(n9919) );
  NANDN U12144 ( .A(n14013), .B(n9919), .Z(n9920) );
  NAND U12145 ( .A(n9920), .B(n14014), .Z(n9922) );
  NANDN U12146 ( .A(n9922), .B(n9921), .Z(n9923) );
  AND U12147 ( .A(n14016), .B(n9923), .Z(n9924) );
  OR U12148 ( .A(n9925), .B(n9924), .Z(n9926) );
  NANDN U12149 ( .A(n14021), .B(n9926), .Z(n9928) );
  NAND U12150 ( .A(n9928), .B(n9927), .Z(n9930) );
  NANDN U12151 ( .A(y[2024]), .B(n9930), .Z(n9929) );
  AND U12152 ( .A(n14027), .B(n9929), .Z(n9933) );
  XNOR U12153 ( .A(y[2024]), .B(n9930), .Z(n9931) );
  NAND U12154 ( .A(n9931), .B(x[2024]), .Z(n9932) );
  NAND U12155 ( .A(n9933), .B(n9932), .Z(n9935) );
  ANDN U12156 ( .B(n9935), .A(n9934), .Z(n9936) );
  NAND U12157 ( .A(n9936), .B(n14028), .Z(n9937) );
  NANDN U12158 ( .A(n14030), .B(n9937), .Z(n9938) );
  NANDN U12159 ( .A(n9939), .B(n9938), .Z(n9940) );
  AND U12160 ( .A(n14035), .B(n9940), .Z(n9941) );
  NANDN U12161 ( .A(n9942), .B(n9941), .Z(n9943) );
  NAND U12162 ( .A(n9943), .B(n14036), .Z(n9945) );
  NANDN U12163 ( .A(n9945), .B(n9944), .Z(n9946) );
  AND U12164 ( .A(n9947), .B(n9946), .Z(n9949) );
  ANDN U12165 ( .B(n9949), .A(n9948), .Z(n9950) );
  NAND U12166 ( .A(n9951), .B(n9950), .Z(n9952) );
  NAND U12167 ( .A(n9953), .B(n9952), .Z(n9954) );
  NANDN U12168 ( .A(n9955), .B(n9954), .Z(n9957) );
  AND U12169 ( .A(n9957), .B(n9956), .Z(n9958) );
  NANDN U12170 ( .A(n9959), .B(n9958), .Z(n9960) );
  NANDN U12171 ( .A(n9961), .B(n9960), .Z(n9963) );
  ANDN U12172 ( .B(n9963), .A(n9962), .Z(n9965) );
  ANDN U12173 ( .B(n9965), .A(n9964), .Z(n9966) );
  ANDN U12174 ( .B(n9967), .A(n9966), .Z(n9968) );
  AND U12175 ( .A(n9969), .B(n9968), .Z(n9970) );
  NANDN U12176 ( .A(ebreg), .B(n9970), .Z(n5) );
  OR U12177 ( .A(n9970), .B(ebreg), .Z(n14077) );
  ANDN U12178 ( .B(y[2041]), .A(x[2041]), .Z(n14061) );
  NANDN U12179 ( .A(y[2040]), .B(x[2040]), .Z(n9972) );
  AND U12180 ( .A(n9972), .B(n9971), .Z(n9976) );
  OR U12181 ( .A(n9974), .B(n9973), .Z(n9975) );
  AND U12182 ( .A(n9976), .B(n9975), .Z(n14059) );
  ANDN U12183 ( .B(n9980), .A(n9979), .Z(n13939) );
  XNOR U12184 ( .A(y[1975]), .B(x[1975]), .Z(n13937) );
  ANDN U12185 ( .B(n9984), .A(n9983), .Z(n13759) );
  AND U12186 ( .A(n9986), .B(n9985), .Z(n13733) );
  XOR U12187 ( .A(n9987), .B(y[1846]), .Z(n13675) );
  NAND U12188 ( .A(n9989), .B(n9988), .Z(n13659) );
  ANDN U12189 ( .B(y[1796]), .A(x[1796]), .Z(n13559) );
  OR U12190 ( .A(n9993), .B(n9992), .Z(n13361) );
  NOR U12191 ( .A(n9995), .B(n9994), .Z(n13021) );
  ANDN U12192 ( .B(n9997), .A(n9996), .Z(n12993) );
  ANDN U12193 ( .B(n9999), .A(n9998), .Z(n12170) );
  ANDN U12194 ( .B(n10001), .A(n10000), .Z(n12154) );
  NAND U12195 ( .A(n10005), .B(n10004), .Z(n11815) );
  NANDN U12196 ( .A(n10007), .B(n10006), .Z(n11663) );
  XOR U12197 ( .A(n10008), .B(x[895]), .Z(n11568) );
  ANDN U12198 ( .B(n10012), .A(n10011), .Z(n11258) );
  ANDN U12199 ( .B(n10031), .A(n10030), .Z(n10672) );
  ANDN U12200 ( .B(n10037), .A(n10036), .Z(n10582) );
  ANDN U12201 ( .B(n10039), .A(n10038), .Z(n10546) );
  XOR U12202 ( .A(n10046), .B(x[97]), .Z(n10176) );
  ANDN U12203 ( .B(n10048), .A(n10047), .Z(n10140) );
  NAND U12204 ( .A(n10050), .B(n10049), .Z(n10054) );
  NANDN U12205 ( .A(n10054), .B(n10053), .Z(n10056) );
  ANDN U12206 ( .B(n10056), .A(n10055), .Z(n10058) );
  NAND U12207 ( .A(n10058), .B(n10057), .Z(n10059) );
  NANDN U12208 ( .A(n10060), .B(n10059), .Z(n10062) );
  ANDN U12209 ( .B(n10062), .A(n10061), .Z(n10064) );
  NANDN U12210 ( .A(n10064), .B(n10063), .Z(n10065) );
  NANDN U12211 ( .A(n10066), .B(n10065), .Z(n10068) );
  NAND U12212 ( .A(n10068), .B(n10067), .Z(n10070) );
  ANDN U12213 ( .B(n10070), .A(n10069), .Z(n10072) );
  NAND U12214 ( .A(n10072), .B(n10071), .Z(n10074) );
  NAND U12215 ( .A(n10074), .B(n10073), .Z(n10076) );
  ANDN U12216 ( .B(n10076), .A(n10075), .Z(n10077) );
  NANDN U12217 ( .A(n10078), .B(n10077), .Z(n10080) );
  NAND U12218 ( .A(n10080), .B(n10079), .Z(n10081) );
  NANDN U12219 ( .A(n10082), .B(n10081), .Z(n10084) );
  NAND U12220 ( .A(n10084), .B(n10083), .Z(n10086) );
  ANDN U12221 ( .B(n10086), .A(n10085), .Z(n10088) );
  NANDN U12222 ( .A(n10088), .B(n10087), .Z(n10089) );
  NANDN U12223 ( .A(n10090), .B(n10089), .Z(n10092) );
  NAND U12224 ( .A(n10092), .B(n10091), .Z(n10094) );
  ANDN U12225 ( .B(n10094), .A(n10093), .Z(n10096) );
  NAND U12226 ( .A(n10096), .B(n10095), .Z(n10098) );
  NAND U12227 ( .A(n10098), .B(n10097), .Z(n10099) );
  AND U12228 ( .A(n10100), .B(n10099), .Z(n10101) );
  NANDN U12229 ( .A(n10102), .B(n10101), .Z(n10103) );
  NANDN U12230 ( .A(n10104), .B(n10103), .Z(n10105) );
  NANDN U12231 ( .A(n10106), .B(n10105), .Z(n10107) );
  NANDN U12232 ( .A(n10108), .B(n10107), .Z(n10110) );
  ANDN U12233 ( .B(n10110), .A(n10109), .Z(n10111) );
  NANDN U12234 ( .A(n10112), .B(n10111), .Z(n10113) );
  NANDN U12235 ( .A(n10114), .B(n10113), .Z(n10116) );
  ANDN U12236 ( .B(n10116), .A(n10115), .Z(n10117) );
  OR U12237 ( .A(n10118), .B(n10117), .Z(n10119) );
  AND U12238 ( .A(n10120), .B(n10119), .Z(n10121) );
  OR U12239 ( .A(n10122), .B(n10121), .Z(n10123) );
  AND U12240 ( .A(n10124), .B(n10123), .Z(n10126) );
  NAND U12241 ( .A(n10126), .B(n10125), .Z(n10127) );
  NANDN U12242 ( .A(n10128), .B(n10127), .Z(n10130) );
  ANDN U12243 ( .B(n10130), .A(n10129), .Z(n10131) );
  NANDN U12244 ( .A(n10132), .B(n10131), .Z(n10133) );
  NANDN U12245 ( .A(n10134), .B(n10133), .Z(n10135) );
  AND U12246 ( .A(n10136), .B(n10135), .Z(n10137) );
  OR U12247 ( .A(n10138), .B(n10137), .Z(n10139) );
  AND U12248 ( .A(n10140), .B(n10139), .Z(n10142) );
  NANDN U12249 ( .A(n10142), .B(n10141), .Z(n10143) );
  NANDN U12250 ( .A(n10144), .B(n10143), .Z(n10145) );
  NANDN U12251 ( .A(n10146), .B(n10145), .Z(n10147) );
  NAND U12252 ( .A(n10148), .B(n10147), .Z(n10150) );
  ANDN U12253 ( .B(x[86]), .A(y[86]), .Z(n10149) );
  OR U12254 ( .A(n10150), .B(n10149), .Z(n10151) );
  NANDN U12255 ( .A(n10152), .B(n10151), .Z(n10153) );
  NANDN U12256 ( .A(n10154), .B(n10153), .Z(n10155) );
  OR U12257 ( .A(n10156), .B(n10155), .Z(n10157) );
  NANDN U12258 ( .A(n10158), .B(n10157), .Z(n10159) );
  NANDN U12259 ( .A(n10160), .B(n10159), .Z(n10162) );
  NANDN U12260 ( .A(n10162), .B(n10161), .Z(n10164) );
  NAND U12261 ( .A(n10164), .B(n10163), .Z(n10166) );
  ANDN U12262 ( .B(n10166), .A(n10165), .Z(n10167) );
  OR U12263 ( .A(n10168), .B(n10167), .Z(n10170) );
  NAND U12264 ( .A(n10170), .B(n10169), .Z(n10171) );
  NANDN U12265 ( .A(n10172), .B(n10171), .Z(n10173) );
  NANDN U12266 ( .A(n10174), .B(n10173), .Z(n10175) );
  NAND U12267 ( .A(n10176), .B(n10175), .Z(n10177) );
  AND U12268 ( .A(n10178), .B(n10177), .Z(n10179) );
  OR U12269 ( .A(n10179), .B(y[98]), .Z(n10183) );
  XNOR U12270 ( .A(n10180), .B(n10179), .Z(n10181) );
  NAND U12271 ( .A(x[98]), .B(n10181), .Z(n10182) );
  NAND U12272 ( .A(n10183), .B(n10182), .Z(n10185) );
  ANDN U12273 ( .B(n10185), .A(n10184), .Z(n10187) );
  OR U12274 ( .A(n10187), .B(n10186), .Z(n10188) );
  NANDN U12275 ( .A(n10189), .B(n10188), .Z(n10191) );
  NAND U12276 ( .A(n10191), .B(n10190), .Z(n10192) );
  NANDN U12277 ( .A(n10193), .B(n10192), .Z(n10195) );
  NAND U12278 ( .A(n10195), .B(n10194), .Z(n10197) );
  ANDN U12279 ( .B(n10197), .A(n10196), .Z(n10198) );
  OR U12280 ( .A(n10199), .B(n10198), .Z(n10200) );
  NANDN U12281 ( .A(n10201), .B(n10200), .Z(n10202) );
  NANDN U12282 ( .A(n10203), .B(n10202), .Z(n10205) );
  NANDN U12283 ( .A(n10205), .B(n10204), .Z(n10207) );
  NAND U12284 ( .A(n10207), .B(n10206), .Z(n10208) );
  NANDN U12285 ( .A(n10209), .B(n10208), .Z(n10210) );
  NANDN U12286 ( .A(n10211), .B(n10210), .Z(n10213) );
  NAND U12287 ( .A(n10213), .B(n10212), .Z(n10215) );
  ANDN U12288 ( .B(n10215), .A(n10214), .Z(n10219) );
  ANDN U12289 ( .B(n10217), .A(n10216), .Z(n10218) );
  NANDN U12290 ( .A(n10219), .B(n10218), .Z(n10220) );
  AND U12291 ( .A(n10221), .B(n10220), .Z(n10222) );
  OR U12292 ( .A(n10223), .B(n10222), .Z(n10224) );
  NANDN U12293 ( .A(n10225), .B(n10224), .Z(n10226) );
  NANDN U12294 ( .A(n10227), .B(n10226), .Z(n10229) );
  NAND U12295 ( .A(n10229), .B(n10228), .Z(n10231) );
  NAND U12296 ( .A(n10231), .B(n10230), .Z(n10233) );
  ANDN U12297 ( .B(n10233), .A(n10232), .Z(n10237) );
  ANDN U12298 ( .B(n10235), .A(n10234), .Z(n10236) );
  NANDN U12299 ( .A(n10237), .B(n10236), .Z(n10238) );
  AND U12300 ( .A(n10239), .B(n10238), .Z(n10241) );
  OR U12301 ( .A(n10241), .B(n10240), .Z(n10242) );
  NANDN U12302 ( .A(n10243), .B(n10242), .Z(n10245) );
  ANDN U12303 ( .B(n10245), .A(n10244), .Z(n10247) );
  NANDN U12304 ( .A(n10247), .B(n10246), .Z(n10249) );
  ANDN U12305 ( .B(n10249), .A(n10248), .Z(n10251) );
  NAND U12306 ( .A(n10251), .B(n10250), .Z(n10253) );
  NAND U12307 ( .A(n10253), .B(n10252), .Z(n10255) );
  ANDN U12308 ( .B(n10255), .A(n10254), .Z(n10256) );
  NANDN U12309 ( .A(n10257), .B(n10256), .Z(n10259) );
  NAND U12310 ( .A(n10259), .B(n10258), .Z(n10261) );
  ANDN U12311 ( .B(n10261), .A(n10260), .Z(n10262) );
  OR U12312 ( .A(n10263), .B(n10262), .Z(n10264) );
  NANDN U12313 ( .A(n10265), .B(n10264), .Z(n10267) );
  NAND U12314 ( .A(n10267), .B(n10266), .Z(n10269) );
  NAND U12315 ( .A(n10269), .B(n10268), .Z(n10270) );
  NANDN U12316 ( .A(n10271), .B(n10270), .Z(n10273) );
  ANDN U12317 ( .B(n10273), .A(n10272), .Z(n10275) );
  NAND U12318 ( .A(n10275), .B(n10274), .Z(n10277) );
  NAND U12319 ( .A(n10277), .B(n10276), .Z(n10279) );
  ANDN U12320 ( .B(n10279), .A(n10278), .Z(n10280) );
  NANDN U12321 ( .A(n10281), .B(n10280), .Z(n10283) );
  ANDN U12322 ( .B(n10301), .A(n10300), .Z(n10303) );
  OR U12323 ( .A(n10303), .B(n10302), .Z(n10304) );
  NANDN U12324 ( .A(n10305), .B(n10304), .Z(n10306) );
  NANDN U12325 ( .A(n10307), .B(n10306), .Z(n10308) );
  NANDN U12326 ( .A(n10309), .B(n10308), .Z(n10310) );
  NANDN U12327 ( .A(n10311), .B(n10310), .Z(n10313) );
  ANDN U12328 ( .B(n10313), .A(n10312), .Z(n10315) );
  NAND U12329 ( .A(n10315), .B(n10314), .Z(n10317) );
  NAND U12330 ( .A(n10317), .B(n10316), .Z(n10319) );
  ANDN U12331 ( .B(n10319), .A(n10318), .Z(n10320) );
  NANDN U12332 ( .A(n10321), .B(n10320), .Z(n10323) );
  NAND U12333 ( .A(n10323), .B(n10322), .Z(n10325) );
  ANDN U12334 ( .B(n10325), .A(n10324), .Z(n10327) );
  NANDN U12335 ( .A(n10327), .B(n10326), .Z(n10329) );
  NAND U12336 ( .A(n10329), .B(n10328), .Z(n10330) );
  NANDN U12337 ( .A(n10331), .B(n10330), .Z(n10333) );
  ANDN U12338 ( .B(n10333), .A(n10332), .Z(n10334) );
  NANDN U12339 ( .A(n10335), .B(n10334), .Z(n10337) );
  NAND U12340 ( .A(n10337), .B(n10336), .Z(n10338) );
  NANDN U12341 ( .A(n10339), .B(n10338), .Z(n10341) );
  NAND U12342 ( .A(n10341), .B(n10340), .Z(n10343) );
  ANDN U12343 ( .B(n10343), .A(n10342), .Z(n10345) );
  NAND U12344 ( .A(n10345), .B(n10344), .Z(n10347) );
  NAND U12345 ( .A(n10347), .B(n10346), .Z(n10349) );
  ANDN U12346 ( .B(n10349), .A(n10348), .Z(n10351) );
  NANDN U12347 ( .A(n10351), .B(n10350), .Z(n10353) );
  NAND U12348 ( .A(n10353), .B(n10352), .Z(n10354) );
  NANDN U12349 ( .A(n10355), .B(n10354), .Z(n10357) );
  NAND U12350 ( .A(n10357), .B(n10356), .Z(n10359) );
  NAND U12351 ( .A(n10359), .B(n10358), .Z(n10361) );
  ANDN U12352 ( .B(n10361), .A(n10360), .Z(n10363) );
  NAND U12353 ( .A(n10363), .B(n10362), .Z(n10365) );
  NAND U12354 ( .A(n10365), .B(n10364), .Z(n10367) );
  ANDN U12355 ( .B(n10367), .A(n10366), .Z(n10368) );
  NANDN U12356 ( .A(n10369), .B(n10368), .Z(n10371) );
  NAND U12357 ( .A(n10371), .B(n10370), .Z(n10373) );
  ANDN U12358 ( .B(n10373), .A(n10372), .Z(n10375) );
  NAND U12359 ( .A(n10375), .B(n10374), .Z(n10376) );
  NANDN U12360 ( .A(n10377), .B(n10376), .Z(n10379) );
  ANDN U12361 ( .B(n10379), .A(n10378), .Z(n10380) );
  NAND U12362 ( .A(n10396), .B(n10395), .Z(n10397) );
  NANDN U12363 ( .A(n10398), .B(n10397), .Z(n10400) );
  ANDN U12364 ( .B(n10400), .A(n10399), .Z(n10401) );
  OR U12365 ( .A(n10402), .B(n10401), .Z(n10403) );
  NANDN U12366 ( .A(n10404), .B(n10403), .Z(n10405) );
  NANDN U12367 ( .A(n10406), .B(n10405), .Z(n10407) );
  NANDN U12368 ( .A(n10408), .B(n10407), .Z(n10409) );
  NANDN U12369 ( .A(n10410), .B(n10409), .Z(n10412) );
  ANDN U12370 ( .B(n10412), .A(n10411), .Z(n10413) );
  OR U12371 ( .A(n10414), .B(n10413), .Z(n10416) );
  NAND U12372 ( .A(n10416), .B(n10415), .Z(n10418) );
  NAND U12373 ( .A(n10418), .B(n10417), .Z(n10420) );
  NAND U12374 ( .A(n10420), .B(n10419), .Z(n10421) );
  NANDN U12375 ( .A(n10422), .B(n10421), .Z(n10424) );
  ANDN U12376 ( .B(n10424), .A(n10423), .Z(n10426) );
  OR U12377 ( .A(n10426), .B(n10425), .Z(n10427) );
  NANDN U12378 ( .A(n10428), .B(n10427), .Z(n10429) );
  NANDN U12379 ( .A(n10430), .B(n10429), .Z(n10431) );
  NANDN U12380 ( .A(n10432), .B(n10431), .Z(n10433) );
  NANDN U12381 ( .A(n10434), .B(n10433), .Z(n10435) );
  AND U12382 ( .A(n10436), .B(n10435), .Z(n10440) );
  ANDN U12383 ( .B(n10438), .A(n10437), .Z(n10439) );
  NANDN U12384 ( .A(n10440), .B(n10439), .Z(n10442) );
  ANDN U12385 ( .B(n10442), .A(n10441), .Z(n10444) );
  OR U12386 ( .A(n10444), .B(n10443), .Z(n10446) );
  ANDN U12387 ( .B(n10446), .A(n10445), .Z(n10448) );
  NAND U12388 ( .A(n10448), .B(n10447), .Z(n10450) );
  NAND U12389 ( .A(n10450), .B(n10449), .Z(n10452) );
  ANDN U12390 ( .B(n10452), .A(n10451), .Z(n10453) );
  NANDN U12391 ( .A(n10454), .B(n10453), .Z(n10456) );
  NAND U12392 ( .A(n10456), .B(n10455), .Z(n10458) );
  ANDN U12393 ( .B(n10458), .A(n10457), .Z(n10459) );
  OR U12394 ( .A(n10460), .B(n10459), .Z(n10461) );
  NANDN U12395 ( .A(n10462), .B(n10461), .Z(n10463) );
  NANDN U12396 ( .A(n10464), .B(n10463), .Z(n10466) );
  NAND U12397 ( .A(n10466), .B(n10465), .Z(n10468) );
  NAND U12398 ( .A(n10468), .B(n10467), .Z(n10470) );
  ANDN U12399 ( .B(n10470), .A(n10469), .Z(n10472) );
  NAND U12400 ( .A(n10472), .B(n10471), .Z(n10473) );
  AND U12401 ( .A(n10474), .B(n10473), .Z(n10476) );
  NAND U12402 ( .A(n10476), .B(n10475), .Z(n10477) );
  AND U12403 ( .A(n10478), .B(n10477), .Z(n10479) );
  NANDN U12404 ( .A(n10480), .B(n10479), .Z(n10481) );
  NANDN U12405 ( .A(n10482), .B(n10481), .Z(n10484) );
  NAND U12406 ( .A(n10484), .B(n10483), .Z(n10486) );
  NAND U12407 ( .A(n10486), .B(n10485), .Z(n10487) );
  NANDN U12408 ( .A(n10488), .B(n10487), .Z(n10489) );
  NANDN U12409 ( .A(n10490), .B(n10489), .Z(n10491) );
  AND U12410 ( .A(n10492), .B(n10491), .Z(n10493) );
  NANDN U12411 ( .A(n10494), .B(n10493), .Z(n10496) );
  NAND U12412 ( .A(n10496), .B(n10495), .Z(n10497) );
  NANDN U12413 ( .A(n10498), .B(n10497), .Z(n10500) );
  ANDN U12414 ( .B(n10500), .A(n10499), .Z(n10504) );
  ANDN U12415 ( .B(n10502), .A(n10501), .Z(n10503) );
  NANDN U12416 ( .A(n10504), .B(n10503), .Z(n10505) );
  AND U12417 ( .A(n10506), .B(n10505), .Z(n10507) );
  OR U12418 ( .A(n10508), .B(n10507), .Z(n10509) );
  NANDN U12419 ( .A(n10510), .B(n10509), .Z(n10512) );
  NAND U12420 ( .A(n10512), .B(n10511), .Z(n10513) );
  NANDN U12421 ( .A(n10514), .B(n10513), .Z(n10516) );
  NAND U12422 ( .A(n10516), .B(n10515), .Z(n10518) );
  ANDN U12423 ( .B(n10518), .A(n10517), .Z(n10522) );
  ANDN U12424 ( .B(n10520), .A(n10519), .Z(n10521) );
  NANDN U12425 ( .A(n10522), .B(n10521), .Z(n10523) );
  AND U12426 ( .A(n10524), .B(n10523), .Z(n10525) );
  OR U12427 ( .A(n10526), .B(n10525), .Z(n10527) );
  NANDN U12428 ( .A(n10528), .B(n10527), .Z(n10530) );
  NAND U12429 ( .A(n10530), .B(n10529), .Z(n10532) );
  ANDN U12430 ( .B(x[298]), .A(y[298]), .Z(n10531) );
  OR U12431 ( .A(n10532), .B(n10531), .Z(n10534) );
  NAND U12432 ( .A(n10534), .B(n10533), .Z(n10535) );
  NANDN U12433 ( .A(n10536), .B(n10535), .Z(n10537) );
  OR U12434 ( .A(n10538), .B(n10537), .Z(n10540) );
  NAND U12435 ( .A(n10540), .B(n10539), .Z(n10542) );
  ANDN U12436 ( .B(n10542), .A(n10541), .Z(n10543) );
  OR U12437 ( .A(n10544), .B(n10543), .Z(n10545) );
  AND U12438 ( .A(n10546), .B(n10545), .Z(n10548) );
  NANDN U12439 ( .A(n10548), .B(n10547), .Z(n10550) );
  ANDN U12440 ( .B(n10550), .A(n10549), .Z(n10552) );
  NAND U12441 ( .A(n10552), .B(n10551), .Z(n10554) );
  NAND U12442 ( .A(n10554), .B(n10553), .Z(n10556) );
  ANDN U12443 ( .B(n10556), .A(n10555), .Z(n10557) );
  NANDN U12444 ( .A(n10558), .B(n10557), .Z(n10560) );
  NAND U12445 ( .A(n10560), .B(n10559), .Z(n10562) );
  ANDN U12446 ( .B(n10562), .A(n10561), .Z(n10563) );
  OR U12447 ( .A(n10564), .B(n10563), .Z(n10565) );
  NANDN U12448 ( .A(n10566), .B(n10565), .Z(n10568) );
  NAND U12449 ( .A(n10568), .B(n10567), .Z(n10569) );
  NANDN U12450 ( .A(n10570), .B(n10569), .Z(n10572) );
  NAND U12451 ( .A(n10572), .B(n10571), .Z(n10574) );
  ANDN U12452 ( .B(n10574), .A(n10573), .Z(n10576) );
  OR U12453 ( .A(n10576), .B(n10575), .Z(n10577) );
  AND U12454 ( .A(n10578), .B(n10577), .Z(n10580) );
  NANDN U12455 ( .A(n10580), .B(n10579), .Z(n10581) );
  AND U12456 ( .A(n10582), .B(n10581), .Z(n10586) );
  OR U12457 ( .A(n10584), .B(n10583), .Z(n10585) );
  NANDN U12458 ( .A(n10586), .B(n10585), .Z(n10588) );
  ANDN U12459 ( .B(n10588), .A(n10587), .Z(n10590) );
  NANDN U12460 ( .A(n10610), .B(n10609), .Z(n10612) );
  NAND U12461 ( .A(n10612), .B(n10611), .Z(n10613) );
  NANDN U12462 ( .A(n10614), .B(n10613), .Z(n10615) );
  AND U12463 ( .A(n10616), .B(n10615), .Z(n10620) );
  ANDN U12464 ( .B(n10618), .A(n10617), .Z(n10619) );
  NANDN U12465 ( .A(n10620), .B(n10619), .Z(n10621) );
  AND U12466 ( .A(n10622), .B(n10621), .Z(n10623) );
  OR U12467 ( .A(n10624), .B(n10623), .Z(n10625) );
  NANDN U12468 ( .A(n10626), .B(n10625), .Z(n10627) );
  NANDN U12469 ( .A(n10628), .B(n10627), .Z(n10630) );
  ANDN U12470 ( .B(x[350]), .A(y[350]), .Z(n10629) );
  OR U12471 ( .A(n10630), .B(n10629), .Z(n10631) );
  NANDN U12472 ( .A(n10632), .B(n10631), .Z(n10633) );
  NANDN U12473 ( .A(n10634), .B(n10633), .Z(n10636) );
  OR U12474 ( .A(n10636), .B(n10635), .Z(n10638) );
  NAND U12475 ( .A(n10638), .B(n10637), .Z(n10640) );
  ANDN U12476 ( .B(n10640), .A(n10639), .Z(n10642) );
  NANDN U12477 ( .A(n10642), .B(n10641), .Z(n10643) );
  NANDN U12478 ( .A(n10644), .B(n10643), .Z(n10645) );
  NANDN U12479 ( .A(n10646), .B(n10645), .Z(n10647) );
  NANDN U12480 ( .A(n10664), .B(n10663), .Z(n10666) );
  NAND U12481 ( .A(n10666), .B(n10665), .Z(n10668) );
  ANDN U12482 ( .B(n10668), .A(n10667), .Z(n10669) );
  OR U12483 ( .A(n10670), .B(n10669), .Z(n10671) );
  AND U12484 ( .A(n10672), .B(n10671), .Z(n10674) );
  NANDN U12485 ( .A(n10674), .B(n10673), .Z(n10675) );
  NANDN U12486 ( .A(n10676), .B(n10675), .Z(n10677) );
  NANDN U12487 ( .A(n10678), .B(n10677), .Z(n10679) );
  AND U12488 ( .A(n10680), .B(n10679), .Z(n10682) );
  NAND U12489 ( .A(n10682), .B(n10681), .Z(n10684) );
  NAND U12490 ( .A(n10684), .B(n10683), .Z(n10686) );
  ANDN U12491 ( .B(n10686), .A(n10685), .Z(n10687) );
  NANDN U12492 ( .A(n10688), .B(n10687), .Z(n10690) );
  NAND U12493 ( .A(n10690), .B(n10689), .Z(n10691) );
  NANDN U12494 ( .A(n10692), .B(n10691), .Z(n10693) );
  NANDN U12495 ( .A(n10694), .B(n10693), .Z(n10695) );
  NANDN U12496 ( .A(n10696), .B(n10695), .Z(n10698) );
  ANDN U12497 ( .B(n10698), .A(n10697), .Z(n10700) );
  NANDN U12498 ( .A(n10700), .B(n10699), .Z(n10701) );
  NANDN U12499 ( .A(n10702), .B(n10701), .Z(n10703) );
  NANDN U12500 ( .A(n10704), .B(n10703), .Z(n10705) );
  NANDN U12501 ( .A(n10706), .B(n10705), .Z(n10707) );
  NANDN U12502 ( .A(n10708), .B(n10707), .Z(n10710) );
  ANDN U12503 ( .B(n10710), .A(n10709), .Z(n10714) );
  ANDN U12504 ( .B(n10712), .A(n10711), .Z(n10713) );
  NANDN U12505 ( .A(n10714), .B(n10713), .Z(n10715) );
  AND U12506 ( .A(n10716), .B(n10715), .Z(n10718) );
  OR U12507 ( .A(n10718), .B(n10717), .Z(n10719) );
  NANDN U12508 ( .A(n10720), .B(n10719), .Z(n10721) );
  AND U12509 ( .A(n10722), .B(n10721), .Z(n10724) );
  NAND U12510 ( .A(n10724), .B(n10723), .Z(n10726) );
  NAND U12511 ( .A(n10726), .B(n10725), .Z(n10728) );
  ANDN U12512 ( .B(n10728), .A(n10727), .Z(n10729) );
  NANDN U12513 ( .A(n10730), .B(n10729), .Z(n10732) );
  NAND U12514 ( .A(n10732), .B(n10731), .Z(n10734) );
  ANDN U12515 ( .B(n10734), .A(n10733), .Z(n10736) );
  NANDN U12516 ( .A(n10736), .B(n10735), .Z(n10737) );
  NANDN U12517 ( .A(n10738), .B(n10737), .Z(n10739) );
  NANDN U12518 ( .A(n10740), .B(n10739), .Z(n10742) );
  OR U12519 ( .A(n10756), .B(n10755), .Z(n10757) );
  NANDN U12520 ( .A(n10758), .B(n10757), .Z(n10759) );
  NANDN U12521 ( .A(n10760), .B(n10759), .Z(n10762) );
  NANDN U12522 ( .A(n10762), .B(n10761), .Z(n10764) );
  NAND U12523 ( .A(n10764), .B(n10763), .Z(n10765) );
  NANDN U12524 ( .A(n10766), .B(n10765), .Z(n10767) );
  OR U12525 ( .A(n10768), .B(n10767), .Z(n10770) );
  NAND U12526 ( .A(n10770), .B(n10769), .Z(n10772) );
  ANDN U12527 ( .B(n10772), .A(n10771), .Z(n10773) );
  OR U12528 ( .A(n10774), .B(n10773), .Z(n10776) );
  NAND U12529 ( .A(n10776), .B(n10775), .Z(n10777) );
  NANDN U12530 ( .A(n10778), .B(n10777), .Z(n10779) );
  AND U12531 ( .A(n10780), .B(n10779), .Z(n10782) );
  NAND U12532 ( .A(n10782), .B(n10781), .Z(n10783) );
  NANDN U12533 ( .A(n10784), .B(n10783), .Z(n10786) );
  ANDN U12534 ( .B(n10786), .A(n10785), .Z(n10787) );
  NANDN U12535 ( .A(n10788), .B(n10787), .Z(n10789) );
  NANDN U12536 ( .A(n10790), .B(n10789), .Z(n10792) );
  ANDN U12537 ( .B(n10792), .A(n10791), .Z(n10793) );
  OR U12538 ( .A(n10794), .B(n10793), .Z(n10795) );
  AND U12539 ( .A(n10796), .B(n10795), .Z(n10798) );
  NAND U12540 ( .A(n10798), .B(n10797), .Z(n10799) );
  NANDN U12541 ( .A(n10800), .B(n10799), .Z(n10802) );
  ANDN U12542 ( .B(n10802), .A(n10801), .Z(n10803) );
  NANDN U12543 ( .A(n10804), .B(n10803), .Z(n10805) );
  NANDN U12544 ( .A(n10806), .B(n10805), .Z(n10808) );
  ANDN U12545 ( .B(n10808), .A(n10807), .Z(n10809) );
  OR U12546 ( .A(n10810), .B(n10809), .Z(n10811) );
  NANDN U12547 ( .A(n10812), .B(n10811), .Z(n10813) );
  NANDN U12548 ( .A(n10814), .B(n10813), .Z(n10816) );
  NAND U12549 ( .A(n10816), .B(n10815), .Z(n10817) );
  NANDN U12550 ( .A(n10818), .B(n10817), .Z(n10820) );
  ANDN U12551 ( .B(n10820), .A(n10819), .Z(n10821) );
  OR U12552 ( .A(n10822), .B(n10821), .Z(n10824) );
  ANDN U12553 ( .B(n10824), .A(n10823), .Z(n10825) );
  OR U12554 ( .A(n10826), .B(n10825), .Z(n10828) );
  NAND U12555 ( .A(n10828), .B(n10827), .Z(n10829) );
  NANDN U12556 ( .A(n10830), .B(n10829), .Z(n10832) );
  NAND U12557 ( .A(n10832), .B(n10831), .Z(n10833) );
  NANDN U12558 ( .A(n10834), .B(n10833), .Z(n10836) );
  ANDN U12559 ( .B(n10836), .A(n10835), .Z(n10837) );
  NANDN U12560 ( .A(n10838), .B(n10837), .Z(n10839) );
  NANDN U12561 ( .A(n10840), .B(n10839), .Z(n10842) );
  NAND U12562 ( .A(n10842), .B(n10841), .Z(n10843) );
  NANDN U12563 ( .A(n10844), .B(n10843), .Z(n10846) );
  ANDN U12564 ( .B(n10846), .A(n10845), .Z(n10848) );
  NAND U12565 ( .A(n10848), .B(n10847), .Z(n10850) );
  NAND U12566 ( .A(n10850), .B(n10849), .Z(n10851) );
  NANDN U12567 ( .A(n10852), .B(n10851), .Z(n10854) );
  ANDN U12568 ( .B(n10854), .A(n10853), .Z(n10855) );
  OR U12569 ( .A(n10856), .B(n10855), .Z(n10857) );
  NANDN U12570 ( .A(n10858), .B(n10857), .Z(n10860) );
  ANDN U12571 ( .B(n10860), .A(n10859), .Z(n10862) );
  NAND U12572 ( .A(n10862), .B(n10861), .Z(n10866) );
  NANDN U12573 ( .A(n10864), .B(n10863), .Z(n10865) );
  NAND U12574 ( .A(n10866), .B(n10865), .Z(n10867) );
  NANDN U12575 ( .A(n10868), .B(n10867), .Z(n10870) );
  ANDN U12576 ( .B(n10870), .A(n10869), .Z(n10872) );
  NANDN U12577 ( .A(n10872), .B(n10871), .Z(n10873) );
  NANDN U12578 ( .A(n10874), .B(n10873), .Z(n10876) );
  NAND U12579 ( .A(n10876), .B(n10875), .Z(n10878) );
  ANDN U12580 ( .B(x[506]), .A(y[506]), .Z(n10877) );
  OR U12581 ( .A(n10878), .B(n10877), .Z(n10879) );
  NANDN U12582 ( .A(n10880), .B(n10879), .Z(n10881) );
  NANDN U12583 ( .A(n10882), .B(n10881), .Z(n10884) );
  OR U12584 ( .A(n10884), .B(n10883), .Z(n10885) );
  NANDN U12585 ( .A(n10886), .B(n10885), .Z(n10888) );
  NAND U12586 ( .A(n10888), .B(n10887), .Z(n10890) );
  NAND U12587 ( .A(n10890), .B(n10889), .Z(n10892) );
  NAND U12588 ( .A(n10892), .B(n10891), .Z(n10894) );
  ANDN U12589 ( .B(n10894), .A(n10893), .Z(n10898) );
  ANDN U12590 ( .B(n10896), .A(n10895), .Z(n10897) );
  NANDN U12591 ( .A(n10898), .B(n10897), .Z(n10900) );
  ANDN U12592 ( .B(n10900), .A(n10899), .Z(n10904) );
  ANDN U12593 ( .B(n10902), .A(n10901), .Z(n10903) );
  NANDN U12594 ( .A(n10904), .B(n10903), .Z(n10905) );
  AND U12595 ( .A(n10906), .B(n10905), .Z(n10907) );
  OR U12596 ( .A(n10908), .B(n10907), .Z(n10910) );
  NAND U12597 ( .A(n10910), .B(n10909), .Z(n10911) );
  NANDN U12598 ( .A(n10912), .B(n10911), .Z(n10914) );
  NAND U12599 ( .A(n10914), .B(n10913), .Z(n10916) );
  NAND U12600 ( .A(n10916), .B(n10915), .Z(n10917) );
  AND U12601 ( .A(n10918), .B(n10917), .Z(n10919) );
  OR U12602 ( .A(n10920), .B(n10919), .Z(n10922) );
  ANDN U12603 ( .B(n10922), .A(n10921), .Z(n10923) );
  OR U12604 ( .A(n10924), .B(n10923), .Z(n10925) );
  NANDN U12605 ( .A(n10926), .B(n10925), .Z(n10928) );
  NAND U12606 ( .A(n10928), .B(n10927), .Z(n10930) );
  ANDN U12607 ( .B(x[532]), .A(y[532]), .Z(n10929) );
  OR U12608 ( .A(n10930), .B(n10929), .Z(n10931) );
  NANDN U12609 ( .A(n10932), .B(n10931), .Z(n10933) );
  NANDN U12610 ( .A(n10934), .B(n10933), .Z(n10935) );
  OR U12611 ( .A(n10936), .B(n10935), .Z(n10937) );
  NANDN U12612 ( .A(n10938), .B(n10937), .Z(n10940) );
  NAND U12613 ( .A(n10940), .B(n10939), .Z(n10941) );
  NANDN U12614 ( .A(n10942), .B(n10941), .Z(n10944) );
  NAND U12615 ( .A(n10944), .B(n10943), .Z(n10946) );
  NAND U12616 ( .A(n10946), .B(n10945), .Z(n10947) );
  NANDN U12617 ( .A(n10948), .B(n10947), .Z(n10950) );
  NAND U12618 ( .A(n10950), .B(n10949), .Z(n10952) );
  NAND U12619 ( .A(n10968), .B(n10967), .Z(n10969) );
  NANDN U12620 ( .A(n10970), .B(n10969), .Z(n10971) );
  NANDN U12621 ( .A(n10972), .B(n10971), .Z(n10973) );
  AND U12622 ( .A(n10974), .B(n10973), .Z(n10978) );
  ANDN U12623 ( .B(n10976), .A(n10975), .Z(n10977) );
  NANDN U12624 ( .A(n10978), .B(n10977), .Z(n10979) );
  AND U12625 ( .A(n10980), .B(n10979), .Z(n10982) );
  OR U12626 ( .A(n10982), .B(n10981), .Z(n10984) );
  ANDN U12627 ( .B(n10984), .A(n10983), .Z(n10986) );
  NANDN U12628 ( .A(n10986), .B(n10985), .Z(n10987) );
  NANDN U12629 ( .A(n10988), .B(n10987), .Z(n10990) );
  NAND U12630 ( .A(n10990), .B(n10989), .Z(n10992) );
  ANDN U12631 ( .B(x[580]), .A(y[580]), .Z(n10991) );
  OR U12632 ( .A(n10992), .B(n10991), .Z(n10994) );
  NAND U12633 ( .A(n10994), .B(n10993), .Z(n10995) );
  NANDN U12634 ( .A(n10996), .B(n10995), .Z(n10997) );
  OR U12635 ( .A(n10998), .B(n10997), .Z(n11000) );
  NAND U12636 ( .A(n11000), .B(n10999), .Z(n11001) );
  NANDN U12637 ( .A(n11002), .B(n11001), .Z(n11003) );
  OR U12638 ( .A(n11004), .B(n11003), .Z(n11005) );
  AND U12639 ( .A(n11006), .B(n11005), .Z(n11008) );
  OR U12640 ( .A(n11008), .B(n11007), .Z(n11009) );
  AND U12641 ( .A(n11010), .B(n11009), .Z(n11011) );
  OR U12642 ( .A(n11012), .B(n11011), .Z(n11013) );
  NANDN U12643 ( .A(n11014), .B(n11013), .Z(n11015) );
  NANDN U12644 ( .A(n11016), .B(n11015), .Z(n11022) );
  NANDN U12645 ( .A(y[591]), .B(n11017), .Z(n11020) );
  XNOR U12646 ( .A(y[591]), .B(n11017), .Z(n11018) );
  NAND U12647 ( .A(n11018), .B(x[591]), .Z(n11019) );
  NAND U12648 ( .A(n11020), .B(n11019), .Z(n11021) );
  AND U12649 ( .A(n11022), .B(n11021), .Z(n11023) );
  OR U12650 ( .A(n11024), .B(n11023), .Z(n11025) );
  NANDN U12651 ( .A(n11026), .B(n11025), .Z(n11028) );
  NAND U12652 ( .A(n11028), .B(n11027), .Z(n11029) );
  NANDN U12653 ( .A(n11030), .B(n11029), .Z(n11031) );
  NANDN U12654 ( .A(n11032), .B(n11031), .Z(n11034) );
  ANDN U12655 ( .B(n11034), .A(n11033), .Z(n11035) );
  OR U12656 ( .A(n11036), .B(n11035), .Z(n11038) );
  NAND U12657 ( .A(n11038), .B(n11037), .Z(n11039) );
  NANDN U12658 ( .A(n11040), .B(n11039), .Z(n11042) );
  NAND U12659 ( .A(n11042), .B(n11041), .Z(n11043) );
  NANDN U12660 ( .A(n11044), .B(n11043), .Z(n11045) );
  AND U12661 ( .A(n11046), .B(n11045), .Z(n11047) );
  OR U12662 ( .A(n11048), .B(n11047), .Z(n11049) );
  NANDN U12663 ( .A(n11050), .B(n11049), .Z(n11051) );
  NANDN U12664 ( .A(n11052), .B(n11051), .Z(n11054) );
  NAND U12665 ( .A(n11054), .B(n11053), .Z(n11055) );
  NANDN U12666 ( .A(n11056), .B(n11055), .Z(n11057) );
  AND U12667 ( .A(n11058), .B(n11057), .Z(n11059) );
  OR U12668 ( .A(n11060), .B(n11059), .Z(n11061) );
  NANDN U12669 ( .A(n11062), .B(n11061), .Z(n11063) );
  NANDN U12670 ( .A(n11064), .B(n11063), .Z(n11066) );
  NAND U12671 ( .A(n11066), .B(n11065), .Z(n11067) );
  NANDN U12672 ( .A(n11068), .B(n11067), .Z(n11070) );
  ANDN U12673 ( .B(n11070), .A(n11069), .Z(n11072) );
  NANDN U12674 ( .A(n11072), .B(n11071), .Z(n11073) );
  NANDN U12675 ( .A(n11074), .B(n11073), .Z(n11076) );
  NAND U12676 ( .A(n11076), .B(n11075), .Z(n11078) );
  ANDN U12677 ( .B(x[628]), .A(y[628]), .Z(n11077) );
  OR U12678 ( .A(n11078), .B(n11077), .Z(n11079) );
  NANDN U12679 ( .A(n11154), .B(n11153), .Z(n11155) );
  NANDN U12680 ( .A(n11156), .B(n11155), .Z(n11157) );
  NANDN U12681 ( .A(n11158), .B(n11157), .Z(n11160) );
  NANDN U12682 ( .A(n11160), .B(n11159), .Z(n11162) );
  NAND U12683 ( .A(n11162), .B(n11161), .Z(n11163) );
  NANDN U12684 ( .A(n11164), .B(n11163), .Z(n11165) );
  OR U12685 ( .A(n11166), .B(n11165), .Z(n11168) );
  NAND U12686 ( .A(n11168), .B(n11167), .Z(n11169) );
  NANDN U12687 ( .A(n11170), .B(n11169), .Z(n11172) );
  NANDN U12688 ( .A(n11172), .B(n11171), .Z(n11174) );
  NAND U12689 ( .A(n11174), .B(n11173), .Z(n11176) );
  NAND U12690 ( .A(n11176), .B(n11175), .Z(n11178) );
  NANDN U12691 ( .A(n11178), .B(n11177), .Z(n11179) );
  NANDN U12692 ( .A(n11180), .B(n11179), .Z(n11181) );
  AND U12693 ( .A(n11182), .B(n11181), .Z(n11183) );
  OR U12694 ( .A(n11184), .B(n11183), .Z(n11186) );
  NAND U12695 ( .A(n11186), .B(n11185), .Z(n11187) );
  NANDN U12696 ( .A(n11188), .B(n11187), .Z(n11189) );
  AND U12697 ( .A(n11190), .B(n11189), .Z(n11192) );
  NAND U12698 ( .A(n11192), .B(n11191), .Z(n11194) );
  NAND U12699 ( .A(n11194), .B(n11193), .Z(n11196) );
  ANDN U12700 ( .B(n11196), .A(n11195), .Z(n11197) );
  NANDN U12701 ( .A(n11198), .B(n11197), .Z(n11199) );
  AND U12702 ( .A(n11200), .B(n11199), .Z(n11201) );
  OR U12703 ( .A(n11202), .B(n11201), .Z(n11203) );
  NANDN U12704 ( .A(n11204), .B(n11203), .Z(n11206) );
  NAND U12705 ( .A(n11206), .B(n11205), .Z(n11208) );
  ANDN U12706 ( .B(x[724]), .A(y[724]), .Z(n11207) );
  OR U12707 ( .A(n11208), .B(n11207), .Z(n11209) );
  NANDN U12708 ( .A(n11210), .B(n11209), .Z(n11211) );
  NANDN U12709 ( .A(n11212), .B(n11211), .Z(n11214) );
  OR U12710 ( .A(n11214), .B(n11213), .Z(n11215) );
  NANDN U12711 ( .A(n11216), .B(n11215), .Z(n11217) );
  NANDN U12712 ( .A(n11218), .B(n11217), .Z(n11220) );
  NAND U12713 ( .A(n11220), .B(n11219), .Z(n11221) );
  AND U12714 ( .A(n11222), .B(n11221), .Z(n11223) );
  NANDN U12715 ( .A(n11224), .B(n11223), .Z(n11226) );
  NAND U12716 ( .A(n11226), .B(n11225), .Z(n11227) );
  NANDN U12717 ( .A(n11228), .B(n11227), .Z(n11229) );
  AND U12718 ( .A(n11230), .B(n11229), .Z(n11232) );
  NOR U12719 ( .A(n11232), .B(n11231), .Z(n11234) );
  NAND U12720 ( .A(n11234), .B(n11233), .Z(n11240) );
  OR U12721 ( .A(n11236), .B(n11235), .Z(n11237) );
  AND U12722 ( .A(n11238), .B(n11237), .Z(n11239) );
  NAND U12723 ( .A(n11240), .B(n11239), .Z(n11241) );
  NANDN U12724 ( .A(n11242), .B(n11241), .Z(n11244) );
  NAND U12725 ( .A(n11244), .B(n11243), .Z(n11246) );
  ANDN U12726 ( .B(n11246), .A(n11245), .Z(n11248) );
  OR U12727 ( .A(n11248), .B(n11247), .Z(n11250) );
  NAND U12728 ( .A(n11250), .B(n11249), .Z(n11251) );
  NANDN U12729 ( .A(n11251), .B(y[745]), .Z(n11254) );
  XNOR U12730 ( .A(n11251), .B(y[745]), .Z(n11252) );
  NANDN U12731 ( .A(x[745]), .B(n11252), .Z(n11253) );
  NAND U12732 ( .A(n11254), .B(n11253), .Z(n11256) );
  XNOR U12733 ( .A(x[746]), .B(y[746]), .Z(n11255) );
  NANDN U12734 ( .A(n11256), .B(n11255), .Z(n11257) );
  NAND U12735 ( .A(n11258), .B(n11257), .Z(n11260) );
  NAND U12736 ( .A(n11260), .B(n11259), .Z(n11261) );
  NANDN U12737 ( .A(n11262), .B(n11261), .Z(n11264) );
  ANDN U12738 ( .B(n11264), .A(n11263), .Z(n11265) );
  OR U12739 ( .A(n11266), .B(n11265), .Z(n11267) );
  AND U12740 ( .A(n11268), .B(n11267), .Z(n11269) );
  OR U12741 ( .A(n11270), .B(n11269), .Z(n11271) );
  NANDN U12742 ( .A(n11272), .B(n11271), .Z(n11274) );
  ANDN U12743 ( .B(n11274), .A(n11273), .Z(n11275) );
  NANDN U12744 ( .A(n11276), .B(n11275), .Z(n11280) );
  NANDN U12745 ( .A(n11278), .B(n11277), .Z(n11279) );
  NAND U12746 ( .A(n11280), .B(n11279), .Z(n11281) );
  NANDN U12747 ( .A(n11282), .B(n11281), .Z(n11284) );
  NAND U12748 ( .A(n11284), .B(n11283), .Z(n11285) );
  NANDN U12749 ( .A(n11286), .B(n11285), .Z(n11288) );
  NAND U12750 ( .A(n11288), .B(n11287), .Z(n11289) );
  NANDN U12751 ( .A(n11290), .B(n11289), .Z(n11291) );
  AND U12752 ( .A(n11292), .B(n11291), .Z(n11293) );
  OR U12753 ( .A(n11294), .B(n11293), .Z(n11295) );
  NANDN U12754 ( .A(n11296), .B(n11295), .Z(n11298) );
  NAND U12755 ( .A(n11298), .B(n11297), .Z(n11300) );
  ANDN U12756 ( .B(x[770]), .A(y[770]), .Z(n11299) );
  OR U12757 ( .A(n11300), .B(n11299), .Z(n11302) );
  NAND U12758 ( .A(n11302), .B(n11301), .Z(n11303) );
  NANDN U12759 ( .A(n11304), .B(n11303), .Z(n11305) );
  OR U12760 ( .A(n11306), .B(n11305), .Z(n11308) );
  NAND U12761 ( .A(n11308), .B(n11307), .Z(n11310) );
  ANDN U12762 ( .B(n11310), .A(n11309), .Z(n11311) );
  OR U12763 ( .A(n11312), .B(n11311), .Z(n11314) );
  ANDN U12764 ( .B(n11314), .A(n11313), .Z(n11316) );
  NAND U12765 ( .A(n11316), .B(n11315), .Z(n11318) );
  NAND U12766 ( .A(n11318), .B(n11317), .Z(n11320) );
  ANDN U12767 ( .B(n11320), .A(n11319), .Z(n11321) );
  NANDN U12768 ( .A(n11322), .B(n11321), .Z(n11324) );
  NAND U12769 ( .A(n11324), .B(n11323), .Z(n11325) );
  NANDN U12770 ( .A(n11326), .B(n11325), .Z(n11327) );
  NANDN U12771 ( .A(n11328), .B(n11327), .Z(n11330) );
  NAND U12772 ( .A(n11330), .B(n11329), .Z(n11332) );
  ANDN U12773 ( .B(n11332), .A(n11331), .Z(n11334) );
  NANDN U12774 ( .A(n11334), .B(n11333), .Z(n11335) );
  NANDN U12775 ( .A(n11336), .B(n11335), .Z(n11338) );
  NAND U12776 ( .A(n11338), .B(n11337), .Z(n11340) );
  NAND U12777 ( .A(n11340), .B(n11339), .Z(n11342) );
  NAND U12778 ( .A(n11342), .B(n11341), .Z(n11344) );
  ANDN U12779 ( .B(n11344), .A(n11343), .Z(n11348) );
  ANDN U12780 ( .B(n11346), .A(n11345), .Z(n11347) );
  NANDN U12781 ( .A(n11348), .B(n11347), .Z(n11349) );
  AND U12782 ( .A(n11350), .B(n11349), .Z(n11351) );
  OR U12783 ( .A(n11352), .B(n11351), .Z(n11354) );
  NAND U12784 ( .A(n11354), .B(n11353), .Z(n11356) );
  ANDN U12785 ( .B(n11356), .A(n11355), .Z(n11358) );
  NAND U12786 ( .A(n11358), .B(n11357), .Z(n11360) );
  NAND U12787 ( .A(n11360), .B(n11359), .Z(n11362) );
  ANDN U12788 ( .B(n11362), .A(n11361), .Z(n11364) );
  NAND U12789 ( .A(n11364), .B(n11363), .Z(n11365) );
  NANDN U12790 ( .A(n11366), .B(n11365), .Z(n11368) );
  ANDN U12791 ( .B(n11368), .A(n11367), .Z(n11370) );
  NAND U12792 ( .A(n11370), .B(n11369), .Z(n11372) );
  NAND U12793 ( .A(n11372), .B(n11371), .Z(n11374) );
  ANDN U12794 ( .B(n11374), .A(n11373), .Z(n11376) );
  NANDN U12795 ( .A(n11376), .B(n11375), .Z(n11377) );
  NANDN U12796 ( .A(n11378), .B(n11377), .Z(n11380) );
  NAND U12797 ( .A(n11380), .B(n11379), .Z(n11381) );
  OR U12798 ( .A(n11400), .B(n11399), .Z(n11402) );
  NAND U12799 ( .A(n11402), .B(n11401), .Z(n11404) );
  NAND U12800 ( .A(n11404), .B(n11403), .Z(n11405) );
  NANDN U12801 ( .A(n11406), .B(n11405), .Z(n11407) );
  NANDN U12802 ( .A(n11408), .B(n11407), .Z(n11409) );
  AND U12803 ( .A(n11410), .B(n11409), .Z(n11411) );
  OR U12804 ( .A(n11412), .B(n11411), .Z(n11414) );
  NAND U12805 ( .A(n11414), .B(n11413), .Z(n11415) );
  NANDN U12806 ( .A(n11416), .B(n11415), .Z(n11418) );
  NAND U12807 ( .A(n11418), .B(n11417), .Z(n11420) );
  ANDN U12808 ( .B(n11420), .A(n11419), .Z(n11422) );
  OR U12809 ( .A(n11422), .B(n11421), .Z(n11423) );
  NANDN U12810 ( .A(n11424), .B(n11423), .Z(n11426) );
  NAND U12811 ( .A(n11426), .B(n11425), .Z(n11428) );
  NAND U12812 ( .A(n11428), .B(n11427), .Z(n11429) );
  NANDN U12813 ( .A(n11430), .B(n11429), .Z(n11431) );
  AND U12814 ( .A(n11432), .B(n11431), .Z(n11436) );
  AND U12815 ( .A(n11434), .B(n11433), .Z(n11435) );
  NANDN U12816 ( .A(n11436), .B(n11435), .Z(n11437) );
  AND U12817 ( .A(n11438), .B(n11437), .Z(n11439) );
  OR U12818 ( .A(n11440), .B(n11439), .Z(n11442) );
  NAND U12819 ( .A(n11442), .B(n11441), .Z(n11443) );
  NANDN U12820 ( .A(n11444), .B(n11443), .Z(n11446) );
  NAND U12821 ( .A(n11446), .B(n11445), .Z(n11447) );
  NANDN U12822 ( .A(n11448), .B(n11447), .Z(n11449) );
  AND U12823 ( .A(n11450), .B(n11449), .Z(n11452) );
  NANDN U12824 ( .A(n11452), .B(n11451), .Z(n11453) );
  NANDN U12825 ( .A(n11454), .B(n11453), .Z(n11456) );
  NAND U12826 ( .A(n11456), .B(n11455), .Z(n11458) );
  NAND U12827 ( .A(n11458), .B(n11457), .Z(n11460) );
  NAND U12828 ( .A(n11460), .B(n11459), .Z(n11461) );
  AND U12829 ( .A(n11462), .B(n11461), .Z(n11463) );
  OR U12830 ( .A(n11464), .B(n11463), .Z(n11466) );
  NAND U12831 ( .A(n11466), .B(n11465), .Z(n11467) );
  NANDN U12832 ( .A(n11468), .B(n11467), .Z(n11470) );
  NAND U12833 ( .A(n11470), .B(n11469), .Z(n11471) );
  AND U12834 ( .A(n11472), .B(n11471), .Z(n11473) );
  NANDN U12835 ( .A(n11474), .B(n11473), .Z(n11476) );
  NAND U12836 ( .A(n11476), .B(n11475), .Z(n11477) );
  NANDN U12837 ( .A(n11478), .B(n11477), .Z(n11479) );
  AND U12838 ( .A(n11480), .B(n11479), .Z(n11482) );
  NANDN U12839 ( .A(n11482), .B(n11481), .Z(n11483) );
  NANDN U12840 ( .A(n11484), .B(n11483), .Z(n11486) );
  NAND U12841 ( .A(n11486), .B(n11485), .Z(n11488) );
  NAND U12842 ( .A(n11488), .B(n11487), .Z(n11490) );
  NAND U12843 ( .A(n11490), .B(n11489), .Z(n11491) );
  AND U12844 ( .A(n11492), .B(n11491), .Z(n11493) );
  OR U12845 ( .A(n11494), .B(n11493), .Z(n11496) );
  NAND U12846 ( .A(n11496), .B(n11495), .Z(n11497) );
  NANDN U12847 ( .A(n11498), .B(n11497), .Z(n11500) );
  NAND U12848 ( .A(n11500), .B(n11499), .Z(n11501) );
  AND U12849 ( .A(n11502), .B(n11501), .Z(n11503) );
  NANDN U12850 ( .A(n11504), .B(n11503), .Z(n11506) );
  NAND U12851 ( .A(n11506), .B(n11505), .Z(n11507) );
  NANDN U12852 ( .A(n11508), .B(n11507), .Z(n11509) );
  AND U12853 ( .A(n11510), .B(n11509), .Z(n11512) );
  NANDN U12854 ( .A(n11512), .B(n11511), .Z(n11513) );
  NANDN U12855 ( .A(n11514), .B(n11513), .Z(n11516) );
  NAND U12856 ( .A(n11516), .B(n11515), .Z(n11518) );
  NAND U12857 ( .A(n11518), .B(n11517), .Z(n11520) );
  NAND U12858 ( .A(n11520), .B(n11519), .Z(n11521) );
  AND U12859 ( .A(n11522), .B(n11521), .Z(n11523) );
  OR U12860 ( .A(n11524), .B(n11523), .Z(n11526) );
  NAND U12861 ( .A(n11526), .B(n11525), .Z(n11527) );
  NANDN U12862 ( .A(n11528), .B(n11527), .Z(n11530) );
  NAND U12863 ( .A(n11530), .B(n11529), .Z(n11531) );
  AND U12864 ( .A(n11532), .B(n11531), .Z(n11533) );
  NANDN U12865 ( .A(n11534), .B(n11533), .Z(n11535) );
  NANDN U12866 ( .A(n11536), .B(n11535), .Z(n11540) );
  NAND U12867 ( .A(n11538), .B(n11537), .Z(n11539) );
  NAND U12868 ( .A(n11540), .B(n11539), .Z(n11542) );
  OR U12869 ( .A(n11542), .B(n11541), .Z(n11544) );
  NAND U12870 ( .A(n11544), .B(n11543), .Z(n11545) );
  NANDN U12871 ( .A(n11546), .B(n11545), .Z(n11548) );
  NAND U12872 ( .A(n11548), .B(n11547), .Z(n11550) );
  NAND U12873 ( .A(n11550), .B(n11549), .Z(n11551) );
  AND U12874 ( .A(n11552), .B(n11551), .Z(n11553) );
  OR U12875 ( .A(n11554), .B(n11553), .Z(n11556) );
  NAND U12876 ( .A(n11556), .B(n11555), .Z(n11557) );
  NANDN U12877 ( .A(n11558), .B(n11557), .Z(n11560) );
  NAND U12878 ( .A(n11560), .B(n11559), .Z(n11561) );
  AND U12879 ( .A(n11562), .B(n11561), .Z(n11563) );
  NANDN U12880 ( .A(n11564), .B(n11563), .Z(n11565) );
  NAND U12881 ( .A(n11566), .B(n11565), .Z(n11567) );
  NAND U12882 ( .A(n11568), .B(n11567), .Z(n11569) );
  AND U12883 ( .A(n11570), .B(n11569), .Z(n11572) );
  OR U12884 ( .A(n11572), .B(y[896]), .Z(n11575) );
  XNOR U12885 ( .A(n11572), .B(n11571), .Z(n11573) );
  NAND U12886 ( .A(x[896]), .B(n11573), .Z(n11574) );
  NAND U12887 ( .A(n11575), .B(n11574), .Z(n11577) );
  ANDN U12888 ( .B(n11577), .A(n11576), .Z(n11579) );
  NANDN U12889 ( .A(n11579), .B(n11578), .Z(n11580) );
  NANDN U12890 ( .A(n11581), .B(n11580), .Z(n11583) );
  NAND U12891 ( .A(n11583), .B(n11582), .Z(n11585) );
  NAND U12892 ( .A(n11585), .B(n11584), .Z(n11586) );
  NANDN U12893 ( .A(n11587), .B(n11586), .Z(n11588) );
  AND U12894 ( .A(n11589), .B(n11588), .Z(n11590) );
  OR U12895 ( .A(n11591), .B(n11590), .Z(n11593) );
  NAND U12896 ( .A(n11593), .B(n11592), .Z(n11594) );
  NANDN U12897 ( .A(n11595), .B(n11594), .Z(n11597) );
  ANDN U12898 ( .B(n11597), .A(n11596), .Z(n11599) );
  NAND U12899 ( .A(n11599), .B(n11598), .Z(n11600) );
  NANDN U12900 ( .A(n11601), .B(n11600), .Z(n11605) );
  NANDN U12901 ( .A(n11603), .B(n11602), .Z(n11604) );
  AND U12902 ( .A(n11605), .B(n11604), .Z(n11606) );
  NANDN U12903 ( .A(n11607), .B(n11606), .Z(n11608) );
  NANDN U12904 ( .A(n11609), .B(n11608), .Z(n11610) );
  NANDN U12905 ( .A(n11611), .B(n11610), .Z(n11612) );
  AND U12906 ( .A(n11613), .B(n11612), .Z(n11615) );
  NANDN U12907 ( .A(n11615), .B(n11614), .Z(n11617) );
  NAND U12908 ( .A(n11617), .B(n11616), .Z(n11618) );
  NANDN U12909 ( .A(n11619), .B(n11618), .Z(n11621) );
  NAND U12910 ( .A(n11621), .B(n11620), .Z(n11622) );
  NANDN U12911 ( .A(n11623), .B(n11622), .Z(n11624) );
  AND U12912 ( .A(n11625), .B(n11624), .Z(n11629) );
  ANDN U12913 ( .B(n11627), .A(n11626), .Z(n11628) );
  NANDN U12914 ( .A(n11629), .B(n11628), .Z(n11630) );
  AND U12915 ( .A(n11631), .B(n11630), .Z(n11632) );
  OR U12916 ( .A(n11633), .B(n11632), .Z(n11635) );
  NAND U12917 ( .A(n11635), .B(n11634), .Z(n11637) );
  NAND U12918 ( .A(n11637), .B(n11636), .Z(n11638) );
  NANDN U12919 ( .A(n11639), .B(n11638), .Z(n11640) );
  NANDN U12920 ( .A(n11641), .B(n11640), .Z(n11642) );
  AND U12921 ( .A(n11643), .B(n11642), .Z(n11644) );
  OR U12922 ( .A(n11645), .B(n11644), .Z(n11646) );
  NANDN U12923 ( .A(n11647), .B(n11646), .Z(n11649) );
  NAND U12924 ( .A(n11649), .B(n11648), .Z(n11650) );
  NANDN U12925 ( .A(n11651), .B(n11650), .Z(n11653) );
  NAND U12926 ( .A(n11653), .B(n11652), .Z(n11655) );
  ANDN U12927 ( .B(n11655), .A(n11654), .Z(n11659) );
  ANDN U12928 ( .B(n11657), .A(n11656), .Z(n11658) );
  NANDN U12929 ( .A(n11659), .B(n11658), .Z(n11661) );
  ANDN U12930 ( .B(n11661), .A(n11660), .Z(n11662) );
  ANDN U12931 ( .B(n11663), .A(n11662), .Z(n11664) );
  NANDN U12932 ( .A(n11665), .B(n11664), .Z(n11666) );
  NANDN U12933 ( .A(n11667), .B(n11666), .Z(n11669) );
  NAND U12934 ( .A(n11669), .B(n11668), .Z(n11670) );
  AND U12935 ( .A(n11671), .B(n11670), .Z(n11673) );
  NANDN U12936 ( .A(n11673), .B(n11672), .Z(n11675) );
  NAND U12937 ( .A(n11675), .B(n11674), .Z(n11676) );
  NANDN U12938 ( .A(n11677), .B(n11676), .Z(n11679) );
  NAND U12939 ( .A(n11679), .B(n11678), .Z(n11680) );
  NANDN U12940 ( .A(n11681), .B(n11680), .Z(n11682) );
  AND U12941 ( .A(n11683), .B(n11682), .Z(n11687) );
  ANDN U12942 ( .B(n11685), .A(n11684), .Z(n11686) );
  NANDN U12943 ( .A(n11687), .B(n11686), .Z(n11688) );
  AND U12944 ( .A(n11689), .B(n11688), .Z(n11691) );
  NANDN U12945 ( .A(n11691), .B(n11690), .Z(n11693) );
  NAND U12946 ( .A(n11693), .B(n11692), .Z(n11694) );
  NANDN U12947 ( .A(n11695), .B(n11694), .Z(n11696) );
  NANDN U12948 ( .A(n11697), .B(n11696), .Z(n11699) );
  NAND U12949 ( .A(n11699), .B(n11698), .Z(n11700) );
  AND U12950 ( .A(n11701), .B(n11700), .Z(n11703) );
  NANDN U12951 ( .A(n11703), .B(n11702), .Z(n11705) );
  NAND U12952 ( .A(n11705), .B(n11704), .Z(n11706) );
  NANDN U12953 ( .A(n11707), .B(n11706), .Z(n11709) );
  NAND U12954 ( .A(n11709), .B(n11708), .Z(n11710) );
  NANDN U12955 ( .A(n11711), .B(n11710), .Z(n11712) );
  AND U12956 ( .A(n11713), .B(n11712), .Z(n11717) );
  AND U12957 ( .A(n11715), .B(n11714), .Z(n11716) );
  NANDN U12958 ( .A(n11717), .B(n11716), .Z(n11718) );
  NAND U12959 ( .A(n11719), .B(n11718), .Z(n11720) );
  NANDN U12960 ( .A(n11720), .B(y[955]), .Z(n11723) );
  XNOR U12961 ( .A(n11720), .B(y[955]), .Z(n11721) );
  NANDN U12962 ( .A(x[955]), .B(n11721), .Z(n11722) );
  AND U12963 ( .A(n11723), .B(n11722), .Z(n11726) );
  OR U12964 ( .A(n11726), .B(x[956]), .Z(n11725) );
  ANDN U12965 ( .B(n11725), .A(n11724), .Z(n11730) );
  XNOR U12966 ( .A(n11727), .B(n11726), .Z(n11728) );
  NAND U12967 ( .A(n11728), .B(y[956]), .Z(n11729) );
  NAND U12968 ( .A(n11730), .B(n11729), .Z(n11732) );
  NAND U12969 ( .A(n11732), .B(n11731), .Z(n11734) );
  NAND U12970 ( .A(n11734), .B(n11733), .Z(n11735) );
  AND U12971 ( .A(n11736), .B(n11735), .Z(n11738) );
  NANDN U12972 ( .A(n11738), .B(n11737), .Z(n11740) );
  NAND U12973 ( .A(n11740), .B(n11739), .Z(n11741) );
  NANDN U12974 ( .A(n11742), .B(n11741), .Z(n11744) );
  NAND U12975 ( .A(n11744), .B(n11743), .Z(n11745) );
  NANDN U12976 ( .A(n11746), .B(n11745), .Z(n11747) );
  AND U12977 ( .A(n11748), .B(n11747), .Z(n11752) );
  AND U12978 ( .A(n11750), .B(n11749), .Z(n11751) );
  NANDN U12979 ( .A(n11752), .B(n11751), .Z(n11753) );
  NAND U12980 ( .A(n11754), .B(n11753), .Z(n11755) );
  NANDN U12981 ( .A(n11755), .B(y[967]), .Z(n11758) );
  XNOR U12982 ( .A(n11755), .B(y[967]), .Z(n11756) );
  NANDN U12983 ( .A(x[967]), .B(n11756), .Z(n11757) );
  AND U12984 ( .A(n11758), .B(n11757), .Z(n11762) );
  OR U12985 ( .A(n11762), .B(x[968]), .Z(n11760) );
  ANDN U12986 ( .B(n11760), .A(n11759), .Z(n11765) );
  XNOR U12987 ( .A(n11762), .B(n11761), .Z(n11763) );
  NAND U12988 ( .A(n11763), .B(y[968]), .Z(n11764) );
  NAND U12989 ( .A(n11765), .B(n11764), .Z(n11767) );
  NAND U12990 ( .A(n11767), .B(n11766), .Z(n11768) );
  NANDN U12991 ( .A(n11769), .B(n11768), .Z(n11770) );
  AND U12992 ( .A(n11771), .B(n11770), .Z(n11773) );
  NANDN U12993 ( .A(n11773), .B(n11772), .Z(n11775) );
  NAND U12994 ( .A(n11775), .B(n11774), .Z(n11776) );
  NANDN U12995 ( .A(n11777), .B(n11776), .Z(n11779) );
  NAND U12996 ( .A(n11779), .B(n11778), .Z(n11780) );
  NANDN U12997 ( .A(n11781), .B(n11780), .Z(n11782) );
  AND U12998 ( .A(n11783), .B(n11782), .Z(n11784) );
  OR U12999 ( .A(n11785), .B(n11784), .Z(n11787) );
  NAND U13000 ( .A(n11787), .B(n11786), .Z(n11788) );
  NANDN U13001 ( .A(n11789), .B(n11788), .Z(n11791) );
  NAND U13002 ( .A(n11791), .B(n11790), .Z(n11792) );
  NANDN U13003 ( .A(n11793), .B(n11792), .Z(n11794) );
  AND U13004 ( .A(n11795), .B(n11794), .Z(n11797) );
  NANDN U13005 ( .A(n11797), .B(n11796), .Z(n11799) );
  NAND U13006 ( .A(n11799), .B(n11798), .Z(n11800) );
  NANDN U13007 ( .A(n11801), .B(n11800), .Z(n11803) );
  NAND U13008 ( .A(n11803), .B(n11802), .Z(n11804) );
  NANDN U13009 ( .A(n11805), .B(n11804), .Z(n11806) );
  AND U13010 ( .A(n11807), .B(n11806), .Z(n11811) );
  ANDN U13011 ( .B(n11809), .A(n11808), .Z(n11810) );
  NANDN U13012 ( .A(n11811), .B(n11810), .Z(n11813) );
  ANDN U13013 ( .B(n11813), .A(n11812), .Z(n11814) );
  ANDN U13014 ( .B(n11815), .A(n11814), .Z(n11816) );
  NANDN U13015 ( .A(n11817), .B(n11816), .Z(n11819) );
  NAND U13016 ( .A(n11819), .B(n11818), .Z(n11820) );
  NANDN U13017 ( .A(n11821), .B(n11820), .Z(n11822) );
  AND U13018 ( .A(n11823), .B(n11822), .Z(n11825) );
  NANDN U13019 ( .A(n11825), .B(n11824), .Z(n11826) );
  AND U13020 ( .A(n11827), .B(n11826), .Z(n11828) );
  OR U13021 ( .A(n11829), .B(n11828), .Z(n11831) );
  NAND U13022 ( .A(n11831), .B(n11830), .Z(n11832) );
  NANDN U13023 ( .A(n11833), .B(n11832), .Z(n11835) );
  NAND U13024 ( .A(n11835), .B(n11834), .Z(n11837) );
  ANDN U13025 ( .B(n11837), .A(n11836), .Z(n11839) );
  NAND U13026 ( .A(n11839), .B(n11838), .Z(n11840) );
  AND U13027 ( .A(n11841), .B(n11840), .Z(n11842) );
  OR U13028 ( .A(n11843), .B(n11842), .Z(n11844) );
  NANDN U13029 ( .A(n11845), .B(n11844), .Z(n11847) );
  NAND U13030 ( .A(n11847), .B(n11846), .Z(n11848) );
  NANDN U13031 ( .A(n11849), .B(n11848), .Z(n11851) );
  NAND U13032 ( .A(n11851), .B(n11850), .Z(n11852) );
  AND U13033 ( .A(n11853), .B(n11852), .Z(n11855) );
  NANDN U13034 ( .A(n11855), .B(n11854), .Z(n11856) );
  AND U13035 ( .A(n11857), .B(n11856), .Z(n11858) );
  OR U13036 ( .A(n11859), .B(n11858), .Z(n11861) );
  NAND U13037 ( .A(n11861), .B(n11860), .Z(n11862) );
  NANDN U13038 ( .A(n11863), .B(n11862), .Z(n11865) );
  NAND U13039 ( .A(n11865), .B(n11864), .Z(n11867) );
  ANDN U13040 ( .B(n11867), .A(n11866), .Z(n11869) );
  NAND U13041 ( .A(n11869), .B(n11868), .Z(n11871) );
  NAND U13042 ( .A(n11871), .B(n11870), .Z(n11873) );
  ANDN U13043 ( .B(n11873), .A(n11872), .Z(n11875) );
  NANDN U13044 ( .A(n11875), .B(n11874), .Z(n11877) );
  ANDN U13045 ( .B(n11877), .A(n11876), .Z(n11879) );
  NANDN U13046 ( .A(n11879), .B(n11878), .Z(n11880) );
  NANDN U13047 ( .A(n11881), .B(n11880), .Z(n11883) );
  NAND U13048 ( .A(n11883), .B(n11882), .Z(n11885) );
  ANDN U13049 ( .B(n11885), .A(n11884), .Z(n11886) );
  OR U13050 ( .A(n11886), .B(x[1022]), .Z(n11890) );
  XNOR U13051 ( .A(n11887), .B(n11886), .Z(n11888) );
  NAND U13052 ( .A(y[1022]), .B(n11888), .Z(n11889) );
  NAND U13053 ( .A(n11890), .B(n11889), .Z(n11892) );
  ANDN U13054 ( .B(n11892), .A(n11891), .Z(n11894) );
  NANDN U13055 ( .A(n11894), .B(n11893), .Z(n11895) );
  NANDN U13056 ( .A(n11896), .B(n11895), .Z(n11898) );
  NAND U13057 ( .A(n11898), .B(n11897), .Z(n11899) );
  NANDN U13058 ( .A(n11900), .B(n11899), .Z(n11902) );
  NAND U13059 ( .A(n11902), .B(n11901), .Z(n11903) );
  AND U13060 ( .A(n11904), .B(n11903), .Z(n11906) );
  NANDN U13061 ( .A(n11906), .B(n11905), .Z(n11907) );
  AND U13062 ( .A(n11908), .B(n11907), .Z(n11910) );
  NANDN U13063 ( .A(n11910), .B(n11909), .Z(n11911) );
  NANDN U13064 ( .A(n11912), .B(n11911), .Z(n11914) );
  ANDN U13065 ( .B(n11914), .A(n11913), .Z(n11915) );
  OR U13066 ( .A(n11916), .B(n11915), .Z(n11917) );
  NANDN U13067 ( .A(n11918), .B(n11917), .Z(n11920) );
  NAND U13068 ( .A(n11920), .B(n11919), .Z(n11921) );
  NANDN U13069 ( .A(n11922), .B(n11921), .Z(n11924) );
  NAND U13070 ( .A(n11924), .B(n11923), .Z(n11926) );
  ANDN U13071 ( .B(n11926), .A(n11925), .Z(n11928) );
  NANDN U13072 ( .A(n11928), .B(n11927), .Z(n11929) );
  NANDN U13073 ( .A(n11930), .B(n11929), .Z(n11932) );
  NAND U13074 ( .A(n11932), .B(n11931), .Z(n11934) );
  NAND U13075 ( .A(n11934), .B(n11933), .Z(n11936) );
  NAND U13076 ( .A(n11936), .B(n11935), .Z(n11938) );
  ANDN U13077 ( .B(n11938), .A(n11937), .Z(n11939) );
  OR U13078 ( .A(n11940), .B(n11939), .Z(n11942) );
  ANDN U13079 ( .B(n11942), .A(n11941), .Z(n11944) );
  NANDN U13080 ( .A(n11944), .B(n11943), .Z(n11946) );
  ANDN U13081 ( .B(n11946), .A(n11945), .Z(n11948) );
  NANDN U13082 ( .A(n11948), .B(n11947), .Z(n11949) );
  NANDN U13083 ( .A(n11950), .B(n11949), .Z(n11952) );
  NAND U13084 ( .A(n11952), .B(n11951), .Z(n11953) );
  AND U13085 ( .A(n11954), .B(n11953), .Z(n11955) );
  OR U13086 ( .A(n11956), .B(n11955), .Z(n11958) );
  NAND U13087 ( .A(n11958), .B(n11957), .Z(n11959) );
  NANDN U13088 ( .A(n11960), .B(n11959), .Z(n11962) );
  NAND U13089 ( .A(n11962), .B(n11961), .Z(n11964) );
  NAND U13090 ( .A(n11964), .B(n11963), .Z(n11966) );
  ANDN U13091 ( .B(n11966), .A(n11965), .Z(n11968) );
  NANDN U13092 ( .A(n11968), .B(n11967), .Z(n11969) );
  AND U13093 ( .A(n11970), .B(n11969), .Z(n11971) );
  OR U13094 ( .A(n11972), .B(n11971), .Z(n11974) );
  NAND U13095 ( .A(n11974), .B(n11973), .Z(n11975) );
  NANDN U13096 ( .A(n11976), .B(n11975), .Z(n11978) );
  NAND U13097 ( .A(n11978), .B(n11977), .Z(n11980) );
  ANDN U13098 ( .B(n11980), .A(n11979), .Z(n11982) );
  NANDN U13099 ( .A(n11982), .B(n11981), .Z(n11983) );
  NANDN U13100 ( .A(n11984), .B(n11983), .Z(n11985) );
  NANDN U13101 ( .A(n11986), .B(n11985), .Z(n11987) );
  AND U13102 ( .A(n11988), .B(n11987), .Z(n11990) );
  NANDN U13103 ( .A(n11990), .B(n11989), .Z(n11992) );
  ANDN U13104 ( .B(n11992), .A(n11991), .Z(n11993) );
  OR U13105 ( .A(n11994), .B(n11993), .Z(n11995) );
  NANDN U13106 ( .A(n11996), .B(n11995), .Z(n11997) );
  NANDN U13107 ( .A(n11998), .B(n11997), .Z(n12000) );
  ANDN U13108 ( .B(n12000), .A(n11999), .Z(n12002) );
  NAND U13109 ( .A(n12002), .B(n12001), .Z(n12004) );
  NAND U13110 ( .A(n12004), .B(n12003), .Z(n12008) );
  NANDN U13111 ( .A(n12006), .B(n12005), .Z(n12007) );
  NANDN U13112 ( .A(n12008), .B(n12007), .Z(n12010) );
  ANDN U13113 ( .B(n12010), .A(n12009), .Z(n12011) );
  OR U13114 ( .A(n12012), .B(n12011), .Z(n12014) );
  NAND U13115 ( .A(n12014), .B(n12013), .Z(n12015) );
  AND U13116 ( .A(n12016), .B(n12015), .Z(n12018) );
  NANDN U13117 ( .A(n12018), .B(n12017), .Z(n12019) );
  NANDN U13118 ( .A(n12020), .B(n12019), .Z(n12022) );
  NAND U13119 ( .A(n12022), .B(n12021), .Z(n12023) );
  NANDN U13120 ( .A(n12024), .B(n12023), .Z(n12026) );
  NAND U13121 ( .A(n12026), .B(n12025), .Z(n12027) );
  NANDN U13122 ( .A(n12028), .B(n12027), .Z(n12029) );
  AND U13123 ( .A(n12030), .B(n12029), .Z(n12032) );
  NANDN U13124 ( .A(n12032), .B(n12031), .Z(n12033) );
  AND U13125 ( .A(n12034), .B(n12033), .Z(n12036) );
  NANDN U13126 ( .A(n12036), .B(n12035), .Z(n12038) );
  NAND U13127 ( .A(n12038), .B(n12037), .Z(n12040) );
  NAND U13128 ( .A(n12040), .B(n12039), .Z(n12042) );
  NAND U13129 ( .A(n12042), .B(n12041), .Z(n12044) );
  NAND U13130 ( .A(n12044), .B(n12043), .Z(n12045) );
  AND U13131 ( .A(n12046), .B(n12045), .Z(n12047) );
  OR U13132 ( .A(n12048), .B(n12047), .Z(n12049) );
  NANDN U13133 ( .A(n12050), .B(n12049), .Z(n12052) );
  NAND U13134 ( .A(n12052), .B(n12051), .Z(n12054) );
  ANDN U13135 ( .B(n12054), .A(n12053), .Z(n12055) );
  OR U13136 ( .A(n12056), .B(n12055), .Z(n12058) );
  ANDN U13137 ( .B(n12058), .A(n12057), .Z(n12060) );
  NANDN U13138 ( .A(n12060), .B(n12059), .Z(n12062) );
  NAND U13139 ( .A(n12062), .B(n12061), .Z(n12063) );
  NANDN U13140 ( .A(n12064), .B(n12063), .Z(n12066) );
  NAND U13141 ( .A(n12066), .B(n12065), .Z(n12068) );
  NAND U13142 ( .A(n12068), .B(n12067), .Z(n12070) );
  ANDN U13143 ( .B(n12070), .A(n12069), .Z(n12071) );
  OR U13144 ( .A(n12072), .B(n12071), .Z(n12073) );
  NANDN U13145 ( .A(n12074), .B(n12073), .Z(n12076) );
  NAND U13146 ( .A(n12076), .B(n12075), .Z(n12077) );
  NANDN U13147 ( .A(n12078), .B(n12077), .Z(n12080) );
  NAND U13148 ( .A(n12080), .B(n12079), .Z(n12082) );
  ANDN U13149 ( .B(n12082), .A(n12081), .Z(n12084) );
  NANDN U13150 ( .A(n12084), .B(n12083), .Z(n12086) );
  ANDN U13151 ( .B(n12086), .A(n12085), .Z(n12088) );
  OR U13152 ( .A(n12088), .B(n12087), .Z(n12090) );
  NAND U13153 ( .A(n12090), .B(n12089), .Z(n12091) );
  AND U13154 ( .A(n12092), .B(n12091), .Z(n12094) );
  NANDN U13155 ( .A(n12094), .B(n12093), .Z(n12095) );
  NANDN U13156 ( .A(n12096), .B(n12095), .Z(n12098) );
  NAND U13157 ( .A(n12098), .B(n12097), .Z(n12099) );
  NANDN U13158 ( .A(n12100), .B(n12099), .Z(n12102) );
  NAND U13159 ( .A(n12102), .B(n12101), .Z(n12104) );
  ANDN U13160 ( .B(n12104), .A(n12103), .Z(n12105) );
  OR U13161 ( .A(n12106), .B(n12105), .Z(n12108) );
  NAND U13162 ( .A(n12108), .B(n12107), .Z(n12110) );
  NAND U13163 ( .A(n12110), .B(n12109), .Z(n12112) );
  AND U13164 ( .A(n12112), .B(n12111), .Z(n12116) );
  OR U13165 ( .A(n12114), .B(n12113), .Z(n12115) );
  AND U13166 ( .A(n12116), .B(n12115), .Z(n12118) );
  NANDN U13167 ( .A(n12118), .B(n12117), .Z(n12119) );
  NANDN U13168 ( .A(n12120), .B(n12119), .Z(n12122) );
  NAND U13169 ( .A(n12122), .B(n12121), .Z(n12123) );
  NANDN U13170 ( .A(n12124), .B(n12123), .Z(n12126) );
  NAND U13171 ( .A(n12126), .B(n12125), .Z(n12128) );
  ANDN U13172 ( .B(n12128), .A(n12127), .Z(n12130) );
  NANDN U13173 ( .A(n12130), .B(n12129), .Z(n12132) );
  NAND U13174 ( .A(n12132), .B(n12131), .Z(n12133) );
  NANDN U13175 ( .A(n12134), .B(n12133), .Z(n12135) );
  AND U13176 ( .A(n12154), .B(n12153), .Z(n12155) );
  OR U13177 ( .A(n12156), .B(n12155), .Z(n12157) );
  NANDN U13178 ( .A(n12158), .B(n12157), .Z(n12159) );
  NANDN U13179 ( .A(n12160), .B(n12159), .Z(n12162) );
  NAND U13180 ( .A(n12162), .B(n12161), .Z(n12163) );
  NANDN U13181 ( .A(n12164), .B(n12163), .Z(n12165) );
  NANDN U13182 ( .A(n12166), .B(n12165), .Z(n12168) );
  NANDN U13183 ( .A(n12168), .B(n12167), .Z(n12169) );
  AND U13184 ( .A(n12170), .B(n12169), .Z(n12171) );
  OR U13185 ( .A(n12172), .B(n12171), .Z(n12173) );
  NANDN U13186 ( .A(n12174), .B(n12173), .Z(n12176) );
  NAND U13187 ( .A(n12176), .B(n12175), .Z(n12178) );
  NAND U13188 ( .A(n12178), .B(n12177), .Z(n12180) );
  NAND U13189 ( .A(n12180), .B(n12179), .Z(n12181) );
  AND U13190 ( .A(n12182), .B(n12181), .Z(n12184) );
  NANDN U13191 ( .A(n12184), .B(n12183), .Z(n12185) );
  AND U13192 ( .A(n12186), .B(n12185), .Z(n12187) );
  NOR U13193 ( .A(n12188), .B(n12187), .Z(n12189) );
  OR U13194 ( .A(n12190), .B(n12189), .Z(n12191) );
  NANDN U13195 ( .A(n12192), .B(n12191), .Z(n12194) );
  NAND U13196 ( .A(n12194), .B(n12193), .Z(n12195) );
  NANDN U13197 ( .A(n12196), .B(n12195), .Z(n12197) );
  NANDN U13198 ( .A(n12198), .B(n12197), .Z(n12200) );
  NAND U13199 ( .A(n12200), .B(n12199), .Z(n12202) );
  ANDN U13200 ( .B(n12202), .A(n12201), .Z(n12203) );
  OR U13201 ( .A(n12204), .B(n12203), .Z(n12206) );
  NAND U13202 ( .A(n12206), .B(n12205), .Z(n12207) );
  NANDN U13203 ( .A(n12208), .B(n12207), .Z(n12210) );
  NAND U13204 ( .A(n12210), .B(n12209), .Z(n12212) );
  NAND U13205 ( .A(n12212), .B(n12211), .Z(n12214) );
  ANDN U13206 ( .B(n12214), .A(n12213), .Z(n12215) );
  OR U13207 ( .A(n12216), .B(n12215), .Z(n12218) );
  ANDN U13208 ( .B(n12218), .A(n12217), .Z(n12220) );
  NANDN U13209 ( .A(n12220), .B(n12219), .Z(n12222) );
  ANDN U13210 ( .B(n12222), .A(n12221), .Z(n12224) );
  NANDN U13211 ( .A(n12224), .B(n12223), .Z(n12226) );
  NAND U13212 ( .A(n12226), .B(n12225), .Z(n12227) );
  NANDN U13213 ( .A(n12228), .B(n12227), .Z(n12229) );
  NANDN U13214 ( .A(n12230), .B(n12229), .Z(n12231) );
  NANDN U13215 ( .A(n12232), .B(n12231), .Z(n12234) );
  NAND U13216 ( .A(n12234), .B(n12233), .Z(n12236) );
  NAND U13217 ( .A(n12236), .B(n12235), .Z(n12237) );
  AND U13218 ( .A(n12238), .B(n12237), .Z(n12239) );
  OR U13219 ( .A(n12240), .B(n12239), .Z(n12242) );
  ANDN U13220 ( .B(n12242), .A(n12241), .Z(n12243) );
  OR U13221 ( .A(n12244), .B(n12243), .Z(n12246) );
  ANDN U13222 ( .B(n12246), .A(n12245), .Z(n12248) );
  NANDN U13223 ( .A(n12248), .B(n12247), .Z(n12249) );
  NANDN U13224 ( .A(n12250), .B(n12249), .Z(n12252) );
  NAND U13225 ( .A(n12252), .B(n12251), .Z(n12254) );
  ANDN U13226 ( .B(n12254), .A(n12253), .Z(n12255) );
  OR U13227 ( .A(n12256), .B(n12255), .Z(n12258) );
  ANDN U13228 ( .B(n12258), .A(n12257), .Z(n12260) );
  NANDN U13229 ( .A(n12260), .B(n12259), .Z(n12262) );
  NAND U13230 ( .A(n12262), .B(n12261), .Z(n12264) );
  NAND U13231 ( .A(n12264), .B(n12263), .Z(n12266) );
  NAND U13232 ( .A(n12266), .B(n12265), .Z(n12267) );
  NANDN U13233 ( .A(n12268), .B(n12267), .Z(n12270) );
  NAND U13234 ( .A(n12270), .B(n12269), .Z(n12271) );
  NANDN U13235 ( .A(n12272), .B(n12271), .Z(n12274) );
  NAND U13236 ( .A(n12274), .B(n12273), .Z(n12275) );
  NANDN U13237 ( .A(n12276), .B(n12275), .Z(n12278) );
  NAND U13238 ( .A(n12278), .B(n12277), .Z(n12280) );
  NAND U13239 ( .A(n12280), .B(n12279), .Z(n12282) );
  ANDN U13240 ( .B(n12282), .A(n12281), .Z(n12283) );
  OR U13241 ( .A(n12284), .B(n12283), .Z(n12286) );
  NAND U13242 ( .A(n12286), .B(n12285), .Z(n12288) );
  NAND U13243 ( .A(n12288), .B(n12287), .Z(n12290) );
  NAND U13244 ( .A(n12290), .B(n12289), .Z(n12291) );
  AND U13245 ( .A(n12292), .B(n12291), .Z(n12294) );
  NANDN U13246 ( .A(n12294), .B(n12293), .Z(n12296) );
  ANDN U13247 ( .B(n12296), .A(n12295), .Z(n12298) );
  NANDN U13248 ( .A(n12298), .B(n12297), .Z(n12299) );
  NANDN U13249 ( .A(n12300), .B(n12299), .Z(n12302) );
  NAND U13250 ( .A(n12302), .B(n12301), .Z(n12303) );
  NANDN U13251 ( .A(n12304), .B(n12303), .Z(n12306) );
  NAND U13252 ( .A(n12306), .B(n12305), .Z(n12308) );
  ANDN U13253 ( .B(n12308), .A(n12307), .Z(n12310) );
  NANDN U13254 ( .A(n12310), .B(n12309), .Z(n12312) );
  AND U13255 ( .A(n12332), .B(n12331), .Z(n12333) );
  OR U13256 ( .A(n12334), .B(n12333), .Z(n12336) );
  NAND U13257 ( .A(n12336), .B(n12335), .Z(n12337) );
  NANDN U13258 ( .A(n12338), .B(n12337), .Z(n12340) );
  ANDN U13259 ( .B(n12340), .A(n12339), .Z(n12341) );
  ANDN U13260 ( .B(n12342), .A(n12341), .Z(n12346) );
  XNOR U13261 ( .A(y[1239]), .B(x[1239]), .Z(n12344) );
  NAND U13262 ( .A(n12344), .B(n12343), .Z(n12345) );
  NAND U13263 ( .A(n12346), .B(n12345), .Z(n12348) );
  NAND U13264 ( .A(n12348), .B(n12347), .Z(n12349) );
  NANDN U13265 ( .A(n12350), .B(n12349), .Z(n12352) );
  ANDN U13266 ( .B(n12352), .A(n12351), .Z(n12354) );
  NANDN U13267 ( .A(n12354), .B(n12353), .Z(n12355) );
  AND U13268 ( .A(n12356), .B(n12355), .Z(n12358) );
  NANDN U13269 ( .A(n12358), .B(n12357), .Z(n12360) );
  NAND U13270 ( .A(n12360), .B(n12359), .Z(n12362) );
  NAND U13271 ( .A(n12362), .B(n12361), .Z(n12363) );
  AND U13272 ( .A(n12364), .B(n12363), .Z(n12366) );
  NANDN U13273 ( .A(n12366), .B(n12365), .Z(n12368) );
  NAND U13274 ( .A(n12368), .B(n12367), .Z(n12369) );
  NAND U13275 ( .A(n12390), .B(n12389), .Z(n12392) );
  ANDN U13276 ( .B(n12392), .A(n12391), .Z(n12393) );
  OR U13277 ( .A(n12394), .B(n12393), .Z(n12395) );
  NANDN U13278 ( .A(n12396), .B(n12395), .Z(n12397) );
  NANDN U13279 ( .A(n12398), .B(n12397), .Z(n12400) );
  NAND U13280 ( .A(n12400), .B(n12399), .Z(n12402) );
  ANDN U13281 ( .B(n12402), .A(n12401), .Z(n12404) );
  OR U13282 ( .A(n12404), .B(n12403), .Z(n12406) );
  NAND U13283 ( .A(n12406), .B(n12405), .Z(n12407) );
  AND U13284 ( .A(n12408), .B(n12407), .Z(n12410) );
  OR U13285 ( .A(n12410), .B(n12409), .Z(n12411) );
  AND U13286 ( .A(n12412), .B(n12411), .Z(n12414) );
  NANDN U13287 ( .A(n12414), .B(n12413), .Z(n12416) );
  NAND U13288 ( .A(n12416), .B(n12415), .Z(n12418) );
  NAND U13289 ( .A(n12418), .B(n12417), .Z(n12420) );
  ANDN U13290 ( .B(n12420), .A(n12419), .Z(n12421) );
  OR U13291 ( .A(n12422), .B(n12421), .Z(n12423) );
  NANDN U13292 ( .A(n12424), .B(n12423), .Z(n12426) );
  NAND U13293 ( .A(n12426), .B(n12425), .Z(n12428) );
  ANDN U13294 ( .B(n12428), .A(n12427), .Z(n12430) );
  NANDN U13295 ( .A(n12430), .B(n12429), .Z(n12431) );
  NANDN U13296 ( .A(n12432), .B(n12431), .Z(n12434) );
  NAND U13297 ( .A(n12434), .B(n12433), .Z(n12435) );
  AND U13298 ( .A(n12436), .B(n12435), .Z(n12437) );
  OR U13299 ( .A(n12438), .B(n12437), .Z(n12439) );
  NANDN U13300 ( .A(n12440), .B(n12439), .Z(n12442) );
  NAND U13301 ( .A(n12442), .B(n12441), .Z(n12444) );
  NAND U13302 ( .A(n12444), .B(n12443), .Z(n12445) );
  NANDN U13303 ( .A(n12446), .B(n12445), .Z(n12447) );
  AND U13304 ( .A(n12448), .B(n12447), .Z(n12450) );
  OR U13305 ( .A(n12450), .B(n12449), .Z(n12452) );
  ANDN U13306 ( .B(n12452), .A(n12451), .Z(n12454) );
  NANDN U13307 ( .A(n12454), .B(n12453), .Z(n12455) );
  NANDN U13308 ( .A(n12456), .B(n12455), .Z(n12457) );
  AND U13309 ( .A(n12458), .B(n12457), .Z(n12460) );
  NANDN U13310 ( .A(n12460), .B(n12459), .Z(n12461) );
  AND U13311 ( .A(n12462), .B(n12461), .Z(n12464) );
  NANDN U13312 ( .A(n12464), .B(n12463), .Z(n12466) );
  NAND U13313 ( .A(n12466), .B(n12465), .Z(n12468) );
  NAND U13314 ( .A(n12468), .B(n12467), .Z(n12470) );
  NAND U13315 ( .A(n12470), .B(n12469), .Z(n12472) );
  NAND U13316 ( .A(n12472), .B(n12471), .Z(n12473) );
  AND U13317 ( .A(n12474), .B(n12473), .Z(n12476) );
  NANDN U13318 ( .A(n12476), .B(n12475), .Z(n12477) );
  NANDN U13319 ( .A(n12478), .B(n12477), .Z(n12480) );
  NAND U13320 ( .A(n12480), .B(n12479), .Z(n12482) );
  NAND U13321 ( .A(n12482), .B(n12481), .Z(n12483) );
  NANDN U13322 ( .A(n12484), .B(n12483), .Z(n12485) );
  AND U13323 ( .A(n12486), .B(n12485), .Z(n12487) );
  OR U13324 ( .A(n12488), .B(n12487), .Z(n12489) );
  AND U13325 ( .A(n12490), .B(n12489), .Z(n12492) );
  NANDN U13326 ( .A(n12492), .B(n12491), .Z(n12494) );
  NAND U13327 ( .A(n12494), .B(n12493), .Z(n12496) );
  NAND U13328 ( .A(n12496), .B(n12495), .Z(n12497) );
  NAND U13329 ( .A(n12498), .B(n12497), .Z(n12499) );
  NANDN U13330 ( .A(n12500), .B(n12499), .Z(n12501) );
  NANDN U13331 ( .A(n12502), .B(n12501), .Z(n12503) );
  NANDN U13332 ( .A(n12504), .B(n12503), .Z(n12506) );
  NAND U13333 ( .A(n12506), .B(n12505), .Z(n12508) );
  ANDN U13334 ( .B(n12508), .A(n12507), .Z(n12510) );
  NANDN U13335 ( .A(n12510), .B(n12509), .Z(n12512) );
  ANDN U13336 ( .B(n12512), .A(n12511), .Z(n12514) );
  NANDN U13337 ( .A(n12514), .B(n12513), .Z(n12516) );
  ANDN U13338 ( .B(n12516), .A(n12515), .Z(n12517) );
  OR U13339 ( .A(n12518), .B(n12517), .Z(n12519) );
  NANDN U13340 ( .A(n12520), .B(n12519), .Z(n12522) );
  NAND U13341 ( .A(n12522), .B(n12521), .Z(n12523) );
  NANDN U13342 ( .A(n12524), .B(n12523), .Z(n12526) );
  NAND U13343 ( .A(n12526), .B(n12525), .Z(n12527) );
  AND U13344 ( .A(n12528), .B(n12527), .Z(n12530) );
  NANDN U13345 ( .A(n12530), .B(n12529), .Z(n12532) );
  ANDN U13346 ( .B(n12532), .A(n12531), .Z(n12534) );
  NANDN U13347 ( .A(n12534), .B(n12533), .Z(n12536) );
  ANDN U13348 ( .B(n12536), .A(n12535), .Z(n12538) );
  NANDN U13349 ( .A(n12538), .B(n12537), .Z(n12539) );
  NANDN U13350 ( .A(n12540), .B(n12539), .Z(n12541) );
  NANDN U13351 ( .A(n12542), .B(n12541), .Z(n12543) );
  NAND U13352 ( .A(n12544), .B(n12543), .Z(n12546) );
  NAND U13353 ( .A(n12546), .B(n12545), .Z(n12548) );
  NAND U13354 ( .A(n12548), .B(n12547), .Z(n12550) );
  ANDN U13355 ( .B(n12550), .A(n12549), .Z(n12552) );
  NANDN U13356 ( .A(n12552), .B(n12551), .Z(n12553) );
  AND U13357 ( .A(n12554), .B(n12553), .Z(n12555) );
  OR U13358 ( .A(n12556), .B(n12555), .Z(n12558) );
  NAND U13359 ( .A(n12558), .B(n12557), .Z(n12559) );
  NANDN U13360 ( .A(n12560), .B(n12559), .Z(n12562) );
  NAND U13361 ( .A(n12562), .B(n12561), .Z(n12563) );
  NANDN U13362 ( .A(n12564), .B(n12563), .Z(n12565) );
  AND U13363 ( .A(n12566), .B(n12565), .Z(n12568) );
  NANDN U13364 ( .A(n12568), .B(n12567), .Z(n12570) );
  ANDN U13365 ( .B(n12570), .A(n12569), .Z(n12572) );
  NANDN U13366 ( .A(n12572), .B(n12571), .Z(n12574) );
  NAND U13367 ( .A(n12574), .B(n12573), .Z(n12576) );
  NAND U13368 ( .A(n12576), .B(n12575), .Z(n12577) );
  AND U13369 ( .A(n12578), .B(n12577), .Z(n12580) );
  NANDN U13370 ( .A(n12580), .B(n12579), .Z(n12581) );
  NANDN U13371 ( .A(n12582), .B(n12581), .Z(n12584) );
  ANDN U13372 ( .B(n12584), .A(n12583), .Z(n12586) );
  NANDN U13373 ( .A(n12586), .B(n12585), .Z(n12588) );
  ANDN U13374 ( .B(n12588), .A(n12587), .Z(n12590) );
  NANDN U13375 ( .A(n12590), .B(n12589), .Z(n12592) );
  ANDN U13376 ( .B(n12592), .A(n12591), .Z(n12594) );
  NANDN U13377 ( .A(n12594), .B(n12593), .Z(n12595) );
  AND U13378 ( .A(n12596), .B(n12595), .Z(n12598) );
  OR U13379 ( .A(n12598), .B(n12597), .Z(n12600) );
  ANDN U13380 ( .B(n12600), .A(n12599), .Z(n12602) );
  NANDN U13381 ( .A(n12602), .B(n12601), .Z(n12604) );
  NAND U13382 ( .A(n12604), .B(n12603), .Z(n12605) );
  AND U13383 ( .A(n12606), .B(n12605), .Z(n12607) );
  OR U13384 ( .A(n12608), .B(n12607), .Z(n12610) );
  NAND U13385 ( .A(n12610), .B(n12609), .Z(n12611) );
  NANDN U13386 ( .A(n12612), .B(n12611), .Z(n12614) );
  NAND U13387 ( .A(n12614), .B(n12613), .Z(n12616) );
  NAND U13388 ( .A(n12616), .B(n12615), .Z(n12618) );
  ANDN U13389 ( .B(n12618), .A(n12617), .Z(n12619) );
  OR U13390 ( .A(n12620), .B(n12619), .Z(n12622) );
  ANDN U13391 ( .B(n12622), .A(n12621), .Z(n12623) );
  OR U13392 ( .A(n12624), .B(n12623), .Z(n12625) );
  NANDN U13393 ( .A(n12626), .B(n12625), .Z(n12628) );
  NAND U13394 ( .A(n12628), .B(n12627), .Z(n12629) );
  NANDN U13395 ( .A(n12630), .B(n12629), .Z(n12631) );
  NANDN U13396 ( .A(n12632), .B(n12631), .Z(n12634) );
  ANDN U13397 ( .B(n12634), .A(n12633), .Z(n12636) );
  NANDN U13398 ( .A(n12636), .B(n12635), .Z(n12638) );
  ANDN U13399 ( .B(n12638), .A(n12637), .Z(n12640) );
  NANDN U13400 ( .A(n12640), .B(n12639), .Z(n12642) );
  ANDN U13401 ( .B(n12642), .A(n12641), .Z(n12644) );
  NANDN U13402 ( .A(n12644), .B(n12643), .Z(n12646) );
  NAND U13403 ( .A(n12646), .B(n12645), .Z(n12647) );
  NANDN U13404 ( .A(n12648), .B(n12647), .Z(n12650) );
  NAND U13405 ( .A(n12650), .B(n12649), .Z(n12652) );
  NAND U13406 ( .A(n12652), .B(n12651), .Z(n12654) );
  ANDN U13407 ( .B(n12654), .A(n12653), .Z(n12655) );
  OR U13408 ( .A(n12656), .B(n12655), .Z(n12658) );
  ANDN U13409 ( .B(n12658), .A(n12657), .Z(n12660) );
  NANDN U13410 ( .A(n12660), .B(n12659), .Z(n12662) );
  ANDN U13411 ( .B(n12662), .A(n12661), .Z(n12664) );
  NANDN U13412 ( .A(n12664), .B(n12663), .Z(n12666) );
  ANDN U13413 ( .B(n12666), .A(n12665), .Z(n12668) );
  OR U13414 ( .A(n12668), .B(n12667), .Z(n12669) );
  AND U13415 ( .A(n12670), .B(n12669), .Z(n12672) );
  NANDN U13416 ( .A(n12672), .B(n12671), .Z(n12674) );
  NAND U13417 ( .A(n12674), .B(n12673), .Z(n12676) );
  NAND U13418 ( .A(n12676), .B(n12675), .Z(n12678) );
  NAND U13419 ( .A(n12678), .B(n12677), .Z(n12680) );
  NAND U13420 ( .A(n12680), .B(n12679), .Z(n12681) );
  AND U13421 ( .A(n12682), .B(n12681), .Z(n12683) );
  OR U13422 ( .A(n12684), .B(n12683), .Z(n12685) );
  NANDN U13423 ( .A(n12686), .B(n12685), .Z(n12687) );
  NANDN U13424 ( .A(n12688), .B(n12687), .Z(n12690) );
  ANDN U13425 ( .B(n12690), .A(n12689), .Z(n12691) );
  OR U13426 ( .A(n12692), .B(n12691), .Z(n12693) );
  AND U13427 ( .A(n12694), .B(n12693), .Z(n12696) );
  NANDN U13428 ( .A(n12696), .B(n12695), .Z(n12698) );
  NAND U13429 ( .A(n12698), .B(n12697), .Z(n12700) );
  NAND U13430 ( .A(n12700), .B(n12699), .Z(n12704) );
  NANDN U13431 ( .A(n12702), .B(n12701), .Z(n12703) );
  NANDN U13432 ( .A(n12704), .B(n12703), .Z(n12706) );
  ANDN U13433 ( .B(n12706), .A(n12705), .Z(n12708) );
  NANDN U13434 ( .A(n12708), .B(n12707), .Z(n12709) );
  NANDN U13435 ( .A(n12710), .B(n12709), .Z(n12712) );
  NAND U13436 ( .A(n12712), .B(n12711), .Z(n12713) );
  NANDN U13437 ( .A(n12714), .B(n12713), .Z(n12715) );
  AND U13438 ( .A(n12716), .B(n12715), .Z(n12718) );
  NANDN U13439 ( .A(n12718), .B(n12717), .Z(n12720) );
  ANDN U13440 ( .B(n12720), .A(n12719), .Z(n12722) );
  NANDN U13441 ( .A(n12722), .B(n12721), .Z(n12723) );
  NANDN U13442 ( .A(n12724), .B(n12723), .Z(n12725) );
  AND U13443 ( .A(n12726), .B(n12725), .Z(n12727) );
  OR U13444 ( .A(n12728), .B(n12727), .Z(n12729) );
  NANDN U13445 ( .A(n12730), .B(n12729), .Z(n12732) );
  NAND U13446 ( .A(n12732), .B(n12731), .Z(n12734) );
  ANDN U13447 ( .B(n12734), .A(n12733), .Z(n12736) );
  NANDN U13448 ( .A(n12736), .B(n12735), .Z(n12737) );
  NANDN U13449 ( .A(n12738), .B(n12737), .Z(n12739) );
  NANDN U13450 ( .A(n12740), .B(n12739), .Z(n12742) );
  NAND U13451 ( .A(n12742), .B(n12741), .Z(n12743) );
  AND U13452 ( .A(n12744), .B(n12743), .Z(n12746) );
  NANDN U13453 ( .A(n12746), .B(n12745), .Z(n12748) );
  ANDN U13454 ( .B(n12748), .A(n12747), .Z(n12750) );
  NANDN U13455 ( .A(n12750), .B(n12749), .Z(n12752) );
  NAND U13456 ( .A(n12752), .B(n12751), .Z(n12753) );
  NANDN U13457 ( .A(n12754), .B(n12753), .Z(n12755) );
  NANDN U13458 ( .A(n12756), .B(n12755), .Z(n12757) );
  NANDN U13459 ( .A(n12758), .B(n12757), .Z(n12764) );
  NANDN U13460 ( .A(y[1443]), .B(n12759), .Z(n12762) );
  XNOR U13461 ( .A(y[1443]), .B(n12759), .Z(n12760) );
  NAND U13462 ( .A(n12760), .B(x[1443]), .Z(n12761) );
  NAND U13463 ( .A(n12762), .B(n12761), .Z(n12763) );
  AND U13464 ( .A(n12764), .B(n12763), .Z(n12765) );
  OR U13465 ( .A(n12766), .B(n12765), .Z(n12774) );
  NANDN U13466 ( .A(n12768), .B(n12767), .Z(n12770) );
  NAND U13467 ( .A(n12770), .B(n12769), .Z(n12771) );
  AND U13468 ( .A(n12772), .B(n12771), .Z(n12773) );
  NAND U13469 ( .A(n12774), .B(n12773), .Z(n12776) );
  NAND U13470 ( .A(n12776), .B(n12775), .Z(n12780) );
  NANDN U13471 ( .A(n12778), .B(n12777), .Z(n12779) );
  NANDN U13472 ( .A(n12780), .B(n12779), .Z(n12781) );
  AND U13473 ( .A(n12782), .B(n12781), .Z(n12784) );
  NANDN U13474 ( .A(n12784), .B(n12783), .Z(n12786) );
  NAND U13475 ( .A(n12786), .B(n12785), .Z(n12788) );
  NAND U13476 ( .A(n12788), .B(n12787), .Z(n12789) );
  NANDN U13477 ( .A(n12790), .B(n12789), .Z(n12791) );
  AND U13478 ( .A(n12792), .B(n12791), .Z(n12794) );
  NANDN U13479 ( .A(n12794), .B(n12793), .Z(n12796) );
  NAND U13480 ( .A(n12796), .B(n12795), .Z(n12797) );
  NANDN U13481 ( .A(n12798), .B(n12797), .Z(n12799) );
  AND U13482 ( .A(n12800), .B(n12799), .Z(n12802) );
  NANDN U13483 ( .A(n12802), .B(n12801), .Z(n12803) );
  AND U13484 ( .A(n12804), .B(n12803), .Z(n12805) );
  OR U13485 ( .A(n12806), .B(n12805), .Z(n12808) );
  NAND U13486 ( .A(n12808), .B(n12807), .Z(n12810) );
  NAND U13487 ( .A(n12810), .B(n12809), .Z(n12812) );
  NAND U13488 ( .A(n12812), .B(n12811), .Z(n12814) );
  NAND U13489 ( .A(n12814), .B(n12813), .Z(n12815) );
  AND U13490 ( .A(n12816), .B(n12815), .Z(n12817) );
  OR U13491 ( .A(n12818), .B(n12817), .Z(n12820) );
  NAND U13492 ( .A(n12820), .B(n12819), .Z(n12821) );
  NANDN U13493 ( .A(n12822), .B(n12821), .Z(n12824) );
  NAND U13494 ( .A(n12824), .B(n12823), .Z(n12825) );
  NANDN U13495 ( .A(n12826), .B(n12825), .Z(n12827) );
  AND U13496 ( .A(n12828), .B(n12827), .Z(n12829) );
  OR U13497 ( .A(n12830), .B(n12829), .Z(n12832) );
  ANDN U13498 ( .B(n12832), .A(n12831), .Z(n12834) );
  NANDN U13499 ( .A(n12834), .B(n12833), .Z(n12835) );
  NANDN U13500 ( .A(n12836), .B(n12835), .Z(n12837) );
  NANDN U13501 ( .A(n12838), .B(n12837), .Z(n12839) );
  NANDN U13502 ( .A(n12840), .B(n12839), .Z(n12842) );
  NAND U13503 ( .A(n12842), .B(n12841), .Z(n12844) );
  ANDN U13504 ( .B(n12844), .A(n12843), .Z(n12846) );
  NANDN U13505 ( .A(n12846), .B(n12845), .Z(n12847) );
  NANDN U13506 ( .A(n12848), .B(n12847), .Z(n12850) );
  NAND U13507 ( .A(n12850), .B(n12849), .Z(n12851) );
  NANDN U13508 ( .A(n12852), .B(n12851), .Z(n12853) );
  NANDN U13509 ( .A(n12854), .B(n12853), .Z(n12855) );
  NANDN U13510 ( .A(n12856), .B(n12855), .Z(n12857) );
  NANDN U13511 ( .A(n12858), .B(n12857), .Z(n12860) );
  NAND U13512 ( .A(n12860), .B(n12859), .Z(n12862) );
  ANDN U13513 ( .B(n12862), .A(n12861), .Z(n12864) );
  NANDN U13514 ( .A(n12864), .B(n12863), .Z(n12865) );
  NANDN U13515 ( .A(n12866), .B(n12865), .Z(n12868) );
  NAND U13516 ( .A(n12868), .B(n12867), .Z(n12870) );
  NAND U13517 ( .A(n12870), .B(n12869), .Z(n12871) );
  NANDN U13518 ( .A(n12872), .B(n12871), .Z(n12874) );
  NAND U13519 ( .A(n12874), .B(n12873), .Z(n12875) );
  AND U13520 ( .A(n12876), .B(n12875), .Z(n12878) );
  NANDN U13521 ( .A(n12878), .B(n12877), .Z(n12879) );
  AND U13522 ( .A(n12880), .B(n12879), .Z(n12881) );
  NOR U13523 ( .A(n12882), .B(n12881), .Z(n12883) );
  OR U13524 ( .A(n12884), .B(n12883), .Z(n12885) );
  NANDN U13525 ( .A(n12886), .B(n12885), .Z(n12888) );
  NAND U13526 ( .A(n12888), .B(n12887), .Z(n12889) );
  NANDN U13527 ( .A(n12890), .B(n12889), .Z(n12892) );
  NAND U13528 ( .A(n12892), .B(n12891), .Z(n12893) );
  AND U13529 ( .A(n12894), .B(n12893), .Z(n12896) );
  OR U13530 ( .A(n12896), .B(n12895), .Z(n12898) );
  NAND U13531 ( .A(n12898), .B(n12897), .Z(n12900) );
  NAND U13532 ( .A(n12900), .B(n12899), .Z(n12901) );
  NANDN U13533 ( .A(n12902), .B(n12901), .Z(n12904) );
  NAND U13534 ( .A(n12904), .B(n12903), .Z(n12906) );
  ANDN U13535 ( .B(n12906), .A(n12905), .Z(n12908) );
  NANDN U13536 ( .A(n12908), .B(n12907), .Z(n12910) );
  NAND U13537 ( .A(n12910), .B(n12909), .Z(n12912) );
  NAND U13538 ( .A(n12912), .B(n12911), .Z(n12914) );
  NAND U13539 ( .A(n12914), .B(n12913), .Z(n12915) );
  AND U13540 ( .A(n12916), .B(n12915), .Z(n12918) );
  NAND U13541 ( .A(n12918), .B(n12917), .Z(n12919) );
  NANDN U13542 ( .A(n12920), .B(n12919), .Z(n12921) );
  AND U13543 ( .A(n12922), .B(n12921), .Z(n12924) );
  NANDN U13544 ( .A(n12924), .B(n12923), .Z(n12925) );
  NANDN U13545 ( .A(n12926), .B(n12925), .Z(n12928) );
  NAND U13546 ( .A(n12928), .B(n12927), .Z(n12929) );
  NANDN U13547 ( .A(n12930), .B(n12929), .Z(n12932) );
  NAND U13548 ( .A(n12932), .B(n12931), .Z(n12934) );
  NAND U13549 ( .A(n12934), .B(n12933), .Z(n12935) );
  NANDN U13550 ( .A(n12936), .B(n12935), .Z(n12938) );
  NAND U13551 ( .A(n12938), .B(n12937), .Z(n12939) );
  AND U13552 ( .A(n12940), .B(n12939), .Z(n12941) );
  OR U13553 ( .A(n12942), .B(n12941), .Z(n12944) );
  NAND U13554 ( .A(n12944), .B(n12943), .Z(n12946) );
  NAND U13555 ( .A(n12946), .B(n12945), .Z(n12947) );
  AND U13556 ( .A(n12948), .B(n12947), .Z(n12950) );
  NANDN U13557 ( .A(n12950), .B(n12949), .Z(n12952) );
  ANDN U13558 ( .B(n12952), .A(n12951), .Z(n12954) );
  NANDN U13559 ( .A(n12954), .B(n12953), .Z(n12955) );
  NANDN U13560 ( .A(n12956), .B(n12955), .Z(n12958) );
  NAND U13561 ( .A(n12958), .B(n12957), .Z(n12959) );
  NANDN U13562 ( .A(n12960), .B(n12959), .Z(n12962) );
  NAND U13563 ( .A(n12962), .B(n12961), .Z(n12963) );
  NANDN U13564 ( .A(n12964), .B(n12963), .Z(n12966) );
  NAND U13565 ( .A(n12966), .B(n12965), .Z(n12968) );
  NAND U13566 ( .A(n12968), .B(n12967), .Z(n12972) );
  OR U13567 ( .A(n12972), .B(y[1544]), .Z(n12969) );
  AND U13568 ( .A(n12970), .B(n12969), .Z(n12975) );
  XNOR U13569 ( .A(n12972), .B(n12971), .Z(n12973) );
  NAND U13570 ( .A(n12973), .B(x[1544]), .Z(n12974) );
  NAND U13571 ( .A(n12975), .B(n12974), .Z(n12976) );
  NANDN U13572 ( .A(n12977), .B(n12976), .Z(n12979) );
  NAND U13573 ( .A(n12979), .B(n12978), .Z(n12981) );
  ANDN U13574 ( .B(n12981), .A(n12980), .Z(n12983) );
  NANDN U13575 ( .A(n12983), .B(n12982), .Z(n12984) );
  NANDN U13576 ( .A(n12985), .B(n12984), .Z(n12986) );
  AND U13577 ( .A(n12987), .B(n12986), .Z(n12988) );
  OR U13578 ( .A(n12989), .B(n12988), .Z(n12990) );
  NANDN U13579 ( .A(n12991), .B(n12990), .Z(n12992) );
  NANDN U13580 ( .A(n12993), .B(n12992), .Z(n12995) );
  NANDN U13581 ( .A(n12995), .B(n12994), .Z(n12996) );
  NANDN U13582 ( .A(n12997), .B(n12996), .Z(n12999) );
  NAND U13583 ( .A(n12999), .B(n12998), .Z(n13001) );
  NAND U13584 ( .A(n13001), .B(n13000), .Z(n13003) );
  NAND U13585 ( .A(n13003), .B(n13002), .Z(n13004) );
  AND U13586 ( .A(n13005), .B(n13004), .Z(n13006) );
  OR U13587 ( .A(n13007), .B(n13006), .Z(n13008) );
  AND U13588 ( .A(n13009), .B(n13008), .Z(n13010) );
  OR U13589 ( .A(n13011), .B(n13010), .Z(n13013) );
  ANDN U13590 ( .B(n13013), .A(n13012), .Z(n13015) );
  NANDN U13591 ( .A(n13015), .B(n13014), .Z(n13016) );
  NANDN U13592 ( .A(n13017), .B(n13016), .Z(n13018) );
  NANDN U13593 ( .A(n13019), .B(n13018), .Z(n13020) );
  NAND U13594 ( .A(n13021), .B(n13020), .Z(n13023) );
  ANDN U13595 ( .B(n13023), .A(n13022), .Z(n13024) );
  OR U13596 ( .A(n13025), .B(n13024), .Z(n13027) );
  NAND U13597 ( .A(n13027), .B(n13026), .Z(n13029) );
  NAND U13598 ( .A(n13029), .B(n13028), .Z(n13031) );
  NAND U13599 ( .A(n13031), .B(n13030), .Z(n13033) );
  NAND U13600 ( .A(n13033), .B(n13032), .Z(n13034) );
  AND U13601 ( .A(n13035), .B(n13034), .Z(n13037) );
  NANDN U13602 ( .A(n13037), .B(n13036), .Z(n13039) );
  NAND U13603 ( .A(n13039), .B(n13038), .Z(n13041) );
  NAND U13604 ( .A(n13041), .B(n13040), .Z(n13043) );
  ANDN U13605 ( .B(n13043), .A(n13042), .Z(n13044) );
  OR U13606 ( .A(n13045), .B(n13044), .Z(n13046) );
  NANDN U13607 ( .A(n13047), .B(n13046), .Z(n13049) );
  NAND U13608 ( .A(n13049), .B(n13048), .Z(n13051) );
  ANDN U13609 ( .B(n13051), .A(n13050), .Z(n13053) );
  NANDN U13610 ( .A(n13053), .B(n13052), .Z(n13054) );
  NANDN U13611 ( .A(n13055), .B(n13054), .Z(n13057) );
  NAND U13612 ( .A(n13057), .B(n13056), .Z(n13059) );
  NAND U13613 ( .A(n13059), .B(n13058), .Z(n13060) );
  NANDN U13614 ( .A(n13061), .B(n13060), .Z(n13063) );
  NAND U13615 ( .A(n13063), .B(n13062), .Z(n13064) );
  AND U13616 ( .A(n13065), .B(n13064), .Z(n13067) );
  NANDN U13617 ( .A(n13067), .B(n13066), .Z(n13068) );
  NANDN U13618 ( .A(n13069), .B(n13068), .Z(n13071) );
  NAND U13619 ( .A(n13071), .B(n13070), .Z(n13072) );
  NANDN U13620 ( .A(n13073), .B(n13072), .Z(n13074) );
  AND U13621 ( .A(n13075), .B(n13074), .Z(n13076) );
  OR U13622 ( .A(n13077), .B(n13076), .Z(n13079) );
  NAND U13623 ( .A(n13079), .B(n13078), .Z(n13080) );
  AND U13624 ( .A(n13081), .B(n13080), .Z(n13082) );
  OR U13625 ( .A(n13083), .B(n13082), .Z(n13084) );
  AND U13626 ( .A(n13085), .B(n13084), .Z(n13086) );
  OR U13627 ( .A(n13087), .B(n13086), .Z(n13088) );
  NANDN U13628 ( .A(n13089), .B(n13088), .Z(n13090) );
  NANDN U13629 ( .A(n13091), .B(n13090), .Z(n13093) );
  NAND U13630 ( .A(n13093), .B(n13092), .Z(n13094) );
  NANDN U13631 ( .A(n13095), .B(n13094), .Z(n13096) );
  AND U13632 ( .A(n13097), .B(n13096), .Z(n13098) );
  OR U13633 ( .A(n13099), .B(n13098), .Z(n13101) );
  NAND U13634 ( .A(n13101), .B(n13100), .Z(n13102) );
  NANDN U13635 ( .A(n13103), .B(n13102), .Z(n13105) );
  NAND U13636 ( .A(n13105), .B(n13104), .Z(n13107) );
  NAND U13637 ( .A(n13107), .B(n13106), .Z(n13109) );
  ANDN U13638 ( .B(n13109), .A(n13108), .Z(n13110) );
  OR U13639 ( .A(n13111), .B(n13110), .Z(n13113) );
  ANDN U13640 ( .B(n13113), .A(n13112), .Z(n13115) );
  NANDN U13641 ( .A(n13115), .B(n13114), .Z(n13116) );
  NANDN U13642 ( .A(n13117), .B(n13116), .Z(n13118) );
  NANDN U13643 ( .A(n13119), .B(n13118), .Z(n13120) );
  AND U13644 ( .A(n13121), .B(n13120), .Z(n13122) );
  OR U13645 ( .A(n13123), .B(n13122), .Z(n13124) );
  NANDN U13646 ( .A(n13125), .B(n13124), .Z(n13127) );
  NAND U13647 ( .A(n13127), .B(n13126), .Z(n13129) );
  NAND U13648 ( .A(n13129), .B(n13128), .Z(n13130) );
  NANDN U13649 ( .A(n13131), .B(n13130), .Z(n13133) );
  NAND U13650 ( .A(n13133), .B(n13132), .Z(n13134) );
  NANDN U13651 ( .A(n13135), .B(n13134), .Z(n13137) );
  NAND U13652 ( .A(n13137), .B(n13136), .Z(n13138) );
  AND U13653 ( .A(n13139), .B(n13138), .Z(n13141) );
  NANDN U13654 ( .A(n13141), .B(n13140), .Z(n13143) );
  ANDN U13655 ( .B(n13143), .A(n13142), .Z(n13147) );
  ANDN U13656 ( .B(n13145), .A(n13144), .Z(n13146) );
  NANDN U13657 ( .A(n13147), .B(n13146), .Z(n13148) );
  AND U13658 ( .A(n13149), .B(n13148), .Z(n13150) );
  OR U13659 ( .A(n13151), .B(n13150), .Z(n13152) );
  NANDN U13660 ( .A(n13153), .B(n13152), .Z(n13155) );
  ANDN U13661 ( .B(n13155), .A(n13154), .Z(n13156) );
  OR U13662 ( .A(n13157), .B(n13156), .Z(n13158) );
  NANDN U13663 ( .A(n13159), .B(n13158), .Z(n13161) );
  NAND U13664 ( .A(n13161), .B(n13160), .Z(n13162) );
  NANDN U13665 ( .A(n13163), .B(n13162), .Z(n13164) );
  NANDN U13666 ( .A(n13165), .B(n13164), .Z(n13166) );
  NANDN U13667 ( .A(n13167), .B(n13166), .Z(n13169) );
  ANDN U13668 ( .B(n13169), .A(n13168), .Z(n13171) );
  NAND U13669 ( .A(n13171), .B(n13170), .Z(n13172) );
  NANDN U13670 ( .A(n13173), .B(n13172), .Z(n13175) );
  ANDN U13671 ( .B(n13175), .A(n13174), .Z(n13177) );
  NANDN U13672 ( .A(n13177), .B(n13176), .Z(n13179) );
  NAND U13673 ( .A(n13179), .B(n13178), .Z(n13180) );
  NANDN U13674 ( .A(n13181), .B(n13180), .Z(n13183) );
  NAND U13675 ( .A(n13183), .B(n13182), .Z(n13184) );
  NANDN U13676 ( .A(n13185), .B(n13184), .Z(n13186) );
  NANDN U13677 ( .A(n13187), .B(n13186), .Z(n13189) );
  NAND U13678 ( .A(n13189), .B(n13188), .Z(n13191) );
  ANDN U13679 ( .B(n13191), .A(n13190), .Z(n13193) );
  NAND U13680 ( .A(n13193), .B(n13192), .Z(n13194) );
  NANDN U13681 ( .A(n13195), .B(n13194), .Z(n13196) );
  NANDN U13682 ( .A(n13197), .B(n13196), .Z(n13199) );
  ANDN U13683 ( .B(n13199), .A(n13198), .Z(n13200) );
  OR U13684 ( .A(n13201), .B(n13200), .Z(n13202) );
  AND U13685 ( .A(n13203), .B(n13202), .Z(n13205) );
  NANDN U13686 ( .A(n13205), .B(n13204), .Z(n13207) );
  NAND U13687 ( .A(n13207), .B(n13206), .Z(n13209) );
  NAND U13688 ( .A(n13209), .B(n13208), .Z(n13211) );
  NAND U13689 ( .A(n13211), .B(n13210), .Z(n13213) );
  NAND U13690 ( .A(n13213), .B(n13212), .Z(n13215) );
  ANDN U13691 ( .B(n13215), .A(n13214), .Z(n13217) );
  NANDN U13692 ( .A(n13217), .B(n13216), .Z(n13218) );
  NANDN U13693 ( .A(n13219), .B(n13218), .Z(n13220) );
  NANDN U13694 ( .A(n13221), .B(n13220), .Z(n13223) );
  NAND U13695 ( .A(n13223), .B(n13222), .Z(n13224) );
  AND U13696 ( .A(n13225), .B(n13224), .Z(n13227) );
  NANDN U13697 ( .A(n13227), .B(n13226), .Z(n13228) );
  NANDN U13698 ( .A(n13229), .B(n13228), .Z(n13230) );
  NANDN U13699 ( .A(n13231), .B(n13230), .Z(n13233) );
  NAND U13700 ( .A(n13233), .B(n13232), .Z(n13234) );
  NANDN U13701 ( .A(n13235), .B(n13234), .Z(n13237) );
  ANDN U13702 ( .B(n13237), .A(n13236), .Z(n13239) );
  NANDN U13703 ( .A(n13239), .B(n13238), .Z(n13240) );
  AND U13704 ( .A(n13241), .B(n13240), .Z(n13242) );
  OR U13705 ( .A(n13243), .B(n13242), .Z(n13245) );
  NAND U13706 ( .A(n13245), .B(n13244), .Z(n13246) );
  NANDN U13707 ( .A(n13247), .B(n13246), .Z(n13249) );
  NANDN U13708 ( .A(n13249), .B(n13248), .Z(n13251) );
  NAND U13709 ( .A(n13251), .B(n13250), .Z(n13253) );
  ANDN U13710 ( .B(n13253), .A(n13252), .Z(n13254) );
  OR U13711 ( .A(n13255), .B(n13254), .Z(n13256) );
  AND U13712 ( .A(n13257), .B(n13256), .Z(n13259) );
  NANDN U13713 ( .A(n13259), .B(n13258), .Z(n13261) );
  NAND U13714 ( .A(n13261), .B(n13260), .Z(n13263) );
  NAND U13715 ( .A(n13263), .B(n13262), .Z(n13265) );
  ANDN U13716 ( .B(n13265), .A(n13264), .Z(n13266) );
  OR U13717 ( .A(n13267), .B(n13266), .Z(n13269) );
  ANDN U13718 ( .B(n13269), .A(n13268), .Z(n13271) );
  NANDN U13719 ( .A(n13271), .B(n13270), .Z(n13272) );
  NANDN U13720 ( .A(n13273), .B(n13272), .Z(n13274) );
  NANDN U13721 ( .A(n13275), .B(n13274), .Z(n13277) );
  NAND U13722 ( .A(n13277), .B(n13276), .Z(n13278) );
  NANDN U13723 ( .A(n13279), .B(n13278), .Z(n13281) );
  ANDN U13724 ( .B(n13281), .A(n13280), .Z(n13283) );
  NANDN U13725 ( .A(n13283), .B(n13282), .Z(n13284) );
  AND U13726 ( .A(n13285), .B(n13284), .Z(n13287) );
  NANDN U13727 ( .A(n13287), .B(n13286), .Z(n13288) );
  AND U13728 ( .A(n13289), .B(n13288), .Z(n13291) );
  NANDN U13729 ( .A(n13291), .B(n13290), .Z(n13292) );
  NANDN U13730 ( .A(n13293), .B(n13292), .Z(n13294) );
  AND U13731 ( .A(n13295), .B(n13294), .Z(n13299) );
  ANDN U13732 ( .B(n13297), .A(n13296), .Z(n13298) );
  NANDN U13733 ( .A(n13299), .B(n13298), .Z(n13300) );
  AND U13734 ( .A(n13301), .B(n13300), .Z(n13302) );
  OR U13735 ( .A(n13303), .B(n13302), .Z(n13305) );
  NAND U13736 ( .A(n13305), .B(n13304), .Z(n13306) );
  NANDN U13737 ( .A(n13307), .B(n13306), .Z(n13309) );
  NAND U13738 ( .A(n13309), .B(n13308), .Z(n13310) );
  NANDN U13739 ( .A(n13311), .B(n13310), .Z(n13313) );
  ANDN U13740 ( .B(n13313), .A(n13312), .Z(n13314) );
  OR U13741 ( .A(n13315), .B(n13314), .Z(n13316) );
  NANDN U13742 ( .A(n13317), .B(n13316), .Z(n13319) );
  NAND U13743 ( .A(n13319), .B(n13318), .Z(n13320) );
  NANDN U13744 ( .A(n13321), .B(n13320), .Z(n13322) );
  NANDN U13745 ( .A(n13323), .B(n13322), .Z(n13324) );
  AND U13746 ( .A(n13325), .B(n13324), .Z(n13327) );
  NANDN U13747 ( .A(n13327), .B(n13326), .Z(n13329) );
  NAND U13748 ( .A(n13329), .B(n13328), .Z(n13331) );
  NAND U13749 ( .A(n13331), .B(n13330), .Z(n13332) );
  NANDN U13750 ( .A(n13333), .B(n13332), .Z(n13334) );
  AND U13751 ( .A(n13335), .B(n13334), .Z(n13337) );
  NANDN U13752 ( .A(n13337), .B(n13336), .Z(n13338) );
  NANDN U13753 ( .A(n13339), .B(n13338), .Z(n13341) );
  NAND U13754 ( .A(n13341), .B(n13340), .Z(n13345) );
  OR U13755 ( .A(n13343), .B(n13342), .Z(n13344) );
  NANDN U13756 ( .A(n13345), .B(n13344), .Z(n13347) );
  ANDN U13757 ( .B(n13347), .A(n13346), .Z(n13348) );
  OR U13758 ( .A(n13349), .B(n13348), .Z(n13350) );
  NANDN U13759 ( .A(n13351), .B(n13350), .Z(n13353) );
  NAND U13760 ( .A(n13353), .B(n13352), .Z(n13355) );
  NAND U13761 ( .A(n13355), .B(n13354), .Z(n13357) );
  NAND U13762 ( .A(n13357), .B(n13356), .Z(n13359) );
  ANDN U13763 ( .B(n13359), .A(n13358), .Z(n13360) );
  NAND U13764 ( .A(n13361), .B(n13360), .Z(n13363) );
  NAND U13765 ( .A(n13363), .B(n13362), .Z(n13364) );
  NANDN U13766 ( .A(n13365), .B(n13364), .Z(n13366) );
  AND U13767 ( .A(n13367), .B(n13366), .Z(n13368) );
  NANDN U13768 ( .A(n13369), .B(n13368), .Z(n13371) );
  NAND U13769 ( .A(n13371), .B(n13370), .Z(n13372) );
  NANDN U13770 ( .A(n13373), .B(n13372), .Z(n13374) );
  AND U13771 ( .A(n13375), .B(n13374), .Z(n13376) );
  OR U13772 ( .A(n13377), .B(n13376), .Z(n13378) );
  AND U13773 ( .A(n13379), .B(n13378), .Z(n13380) );
  OR U13774 ( .A(n13381), .B(n13380), .Z(n13382) );
  NANDN U13775 ( .A(n13383), .B(n13382), .Z(n13385) );
  NAND U13776 ( .A(n13385), .B(n13384), .Z(n13387) );
  ANDN U13777 ( .B(n13387), .A(n13386), .Z(n13389) );
  NAND U13778 ( .A(n13389), .B(n13388), .Z(n13391) );
  NAND U13779 ( .A(n13391), .B(n13390), .Z(n13393) );
  NAND U13780 ( .A(n13393), .B(n13392), .Z(n13395) );
  NAND U13781 ( .A(n13395), .B(n13394), .Z(n13396) );
  NANDN U13782 ( .A(n13397), .B(n13396), .Z(n13399) );
  ANDN U13783 ( .B(n13399), .A(n13398), .Z(n13401) );
  NANDN U13784 ( .A(n13401), .B(n13400), .Z(n13403) );
  NAND U13785 ( .A(n13403), .B(n13402), .Z(n13405) );
  NAND U13786 ( .A(n13405), .B(n13404), .Z(n13406) );
  NANDN U13787 ( .A(n13407), .B(n13406), .Z(n13408) );
  NANDN U13788 ( .A(n13409), .B(n13408), .Z(n13411) );
  ANDN U13789 ( .B(n13411), .A(n13410), .Z(n13412) );
  ANDN U13790 ( .B(n13413), .A(n13412), .Z(n13415) );
  NANDN U13791 ( .A(n13415), .B(n13414), .Z(n13416) );
  NANDN U13792 ( .A(n13417), .B(n13416), .Z(n13419) );
  NAND U13793 ( .A(n13419), .B(n13418), .Z(n13421) );
  AND U13794 ( .A(n13439), .B(n13438), .Z(n13441) );
  NANDN U13795 ( .A(n13441), .B(n13440), .Z(n13443) );
  NAND U13796 ( .A(n13443), .B(n13442), .Z(n13444) );
  NANDN U13797 ( .A(n13445), .B(n13444), .Z(n13446) );
  NANDN U13798 ( .A(n13447), .B(n13446), .Z(n13449) );
  NAND U13799 ( .A(n13449), .B(n13448), .Z(n13450) );
  AND U13800 ( .A(n13451), .B(n13450), .Z(n13453) );
  NANDN U13801 ( .A(n13453), .B(n13452), .Z(n13455) );
  ANDN U13802 ( .B(n13455), .A(n13454), .Z(n13457) );
  NAND U13803 ( .A(n13457), .B(n13456), .Z(n13461) );
  AND U13804 ( .A(n13459), .B(n13458), .Z(n13460) );
  NAND U13805 ( .A(n13461), .B(n13460), .Z(n13462) );
  NANDN U13806 ( .A(n13463), .B(n13462), .Z(n13467) );
  NANDN U13807 ( .A(n13465), .B(n13464), .Z(n13466) );
  NANDN U13808 ( .A(n13467), .B(n13466), .Z(n13468) );
  AND U13809 ( .A(n13469), .B(n13468), .Z(n13471) );
  NANDN U13810 ( .A(n13471), .B(n13470), .Z(n13473) );
  NAND U13811 ( .A(n13473), .B(n13472), .Z(n13475) );
  NAND U13812 ( .A(n13475), .B(n13474), .Z(n13477) );
  NAND U13813 ( .A(n13477), .B(n13476), .Z(n13479) );
  ANDN U13814 ( .B(n13479), .A(n13478), .Z(n13481) );
  NANDN U13815 ( .A(n13481), .B(n13480), .Z(n13483) );
  NAND U13816 ( .A(n13483), .B(n13482), .Z(n13485) );
  NAND U13817 ( .A(n13485), .B(n13484), .Z(n13486) );
  NANDN U13818 ( .A(n13487), .B(n13486), .Z(n13489) );
  NAND U13819 ( .A(n13489), .B(n13488), .Z(n13491) );
  NAND U13820 ( .A(n13491), .B(n13490), .Z(n13493) );
  NAND U13821 ( .A(n13493), .B(n13492), .Z(n13495) );
  NAND U13822 ( .A(n13495), .B(n13494), .Z(n13497) );
  ANDN U13823 ( .B(n13497), .A(n13496), .Z(n13499) );
  NANDN U13824 ( .A(n13499), .B(n13498), .Z(n13500) );
  NANDN U13825 ( .A(n13501), .B(n13500), .Z(n13503) );
  NAND U13826 ( .A(n13503), .B(n13502), .Z(n13504) );
  NANDN U13827 ( .A(n13505), .B(n13504), .Z(n13507) );
  NAND U13828 ( .A(n13507), .B(n13506), .Z(n13509) );
  ANDN U13829 ( .B(n13509), .A(n13508), .Z(n13511) );
  NANDN U13830 ( .A(n13511), .B(n13510), .Z(n13512) );
  AND U13831 ( .A(n13513), .B(n13512), .Z(n13514) );
  OR U13832 ( .A(n13515), .B(n13514), .Z(n13516) );
  AND U13833 ( .A(n13517), .B(n13516), .Z(n13519) );
  NANDN U13834 ( .A(n13519), .B(n13518), .Z(n13520) );
  NANDN U13835 ( .A(n13521), .B(n13520), .Z(n13523) );
  NAND U13836 ( .A(n13523), .B(n13522), .Z(n13525) );
  NAND U13837 ( .A(n13525), .B(n13524), .Z(n13527) );
  NAND U13838 ( .A(n13527), .B(n13526), .Z(n13529) );
  ANDN U13839 ( .B(n13529), .A(n13528), .Z(n13530) );
  OR U13840 ( .A(n13531), .B(n13530), .Z(n13532) );
  NANDN U13841 ( .A(n13533), .B(n13532), .Z(n13534) );
  NANDN U13842 ( .A(n13535), .B(n13534), .Z(n13536) );
  NANDN U13843 ( .A(n13537), .B(n13536), .Z(n13538) );
  NANDN U13844 ( .A(n13539), .B(n13538), .Z(n13540) );
  AND U13845 ( .A(n13541), .B(n13540), .Z(n13542) );
  OR U13846 ( .A(n13543), .B(n13542), .Z(n13545) );
  NAND U13847 ( .A(n13545), .B(n13544), .Z(n13546) );
  NANDN U13848 ( .A(n13547), .B(n13546), .Z(n13549) );
  NAND U13849 ( .A(n13549), .B(n13548), .Z(n13550) );
  NANDN U13850 ( .A(n13551), .B(n13550), .Z(n13552) );
  AND U13851 ( .A(n13553), .B(n13552), .Z(n13554) );
  OR U13852 ( .A(n13555), .B(n13554), .Z(n13557) );
  ANDN U13853 ( .B(n13557), .A(n13556), .Z(n13558) );
  ANDN U13854 ( .B(n13573), .A(n13572), .Z(n13575) );
  NANDN U13855 ( .A(n13575), .B(n13574), .Z(n13577) );
  NAND U13856 ( .A(n13577), .B(n13576), .Z(n13578) );
  NANDN U13857 ( .A(n13579), .B(n13578), .Z(n13580) );
  NANDN U13858 ( .A(n13581), .B(n13580), .Z(n13583) );
  NAND U13859 ( .A(n13583), .B(n13582), .Z(n13585) );
  ANDN U13860 ( .B(n13585), .A(n13584), .Z(n13586) );
  OR U13861 ( .A(n13587), .B(n13586), .Z(n13588) );
  NANDN U13862 ( .A(n13589), .B(n13588), .Z(n13591) );
  NAND U13863 ( .A(n13591), .B(n13590), .Z(n13593) );
  NAND U13864 ( .A(n13593), .B(n13592), .Z(n13595) );
  NAND U13865 ( .A(n13595), .B(n13594), .Z(n13596) );
  AND U13866 ( .A(n13597), .B(n13596), .Z(n13599) );
  NANDN U13867 ( .A(n13599), .B(n13598), .Z(n13600) );
  AND U13868 ( .A(n13601), .B(n13600), .Z(n13603) );
  NANDN U13869 ( .A(n13603), .B(n13602), .Z(n13604) );
  NANDN U13870 ( .A(n13605), .B(n13604), .Z(n13606) );
  NANDN U13871 ( .A(n13607), .B(n13606), .Z(n13608) );
  NANDN U13872 ( .A(n13609), .B(n13608), .Z(n13611) );
  AND U13873 ( .A(n13611), .B(n13610), .Z(n13612) );
  OR U13874 ( .A(n13612), .B(x[1823]), .Z(n13615) );
  XOR U13875 ( .A(x[1823]), .B(n13612), .Z(n13613) );
  NAND U13876 ( .A(y[1823]), .B(n13613), .Z(n13614) );
  NAND U13877 ( .A(n13615), .B(n13614), .Z(n13616) );
  AND U13878 ( .A(n13617), .B(n13616), .Z(n13619) );
  NANDN U13879 ( .A(n13619), .B(n13618), .Z(n13620) );
  NANDN U13880 ( .A(n13621), .B(n13620), .Z(n13623) );
  NANDN U13881 ( .A(n13623), .B(n13622), .Z(n13625) );
  NAND U13882 ( .A(n13625), .B(n13624), .Z(n13626) );
  NANDN U13883 ( .A(n13627), .B(n13626), .Z(n13628) );
  NANDN U13884 ( .A(n13629), .B(n13628), .Z(n13630) );
  NANDN U13885 ( .A(n13631), .B(n13630), .Z(n13632) );
  AND U13886 ( .A(n13633), .B(n13632), .Z(n13635) );
  NANDN U13887 ( .A(n13635), .B(n13634), .Z(n13637) );
  NAND U13888 ( .A(n13637), .B(n13636), .Z(n13639) );
  NAND U13889 ( .A(n13639), .B(n13638), .Z(n13641) );
  NAND U13890 ( .A(n13641), .B(n13640), .Z(n13643) );
  NAND U13891 ( .A(n13643), .B(n13642), .Z(n13645) );
  ANDN U13892 ( .B(n13645), .A(n13644), .Z(n13647) );
  NANDN U13893 ( .A(n13647), .B(n13646), .Z(n13648) );
  NANDN U13894 ( .A(n13649), .B(n13648), .Z(n13651) );
  NAND U13895 ( .A(n13651), .B(n13650), .Z(n13652) );
  NANDN U13896 ( .A(n13653), .B(n13652), .Z(n13655) );
  ANDN U13897 ( .B(n13655), .A(n13654), .Z(n13657) );
  NAND U13898 ( .A(n13657), .B(n13656), .Z(n13658) );
  NANDN U13899 ( .A(n13659), .B(n13658), .Z(n13660) );
  AND U13900 ( .A(n13661), .B(n13660), .Z(n13662) );
  NANDN U13901 ( .A(n13663), .B(n13662), .Z(n13665) );
  NAND U13902 ( .A(n13665), .B(n13664), .Z(n13666) );
  AND U13903 ( .A(n13667), .B(n13666), .Z(n13669) );
  NANDN U13904 ( .A(n13669), .B(n13668), .Z(n13670) );
  AND U13905 ( .A(n13671), .B(n13670), .Z(n13672) );
  OR U13906 ( .A(n13673), .B(n13672), .Z(n13674) );
  NAND U13907 ( .A(n13675), .B(n13674), .Z(n13676) );
  NAND U13908 ( .A(n13677), .B(n13676), .Z(n13679) );
  NANDN U13909 ( .A(n13679), .B(n13678), .Z(n13681) );
  ANDN U13910 ( .B(n13681), .A(n13680), .Z(n13683) );
  NAND U13911 ( .A(n13683), .B(n13682), .Z(n13685) );
  NAND U13912 ( .A(n13685), .B(n13684), .Z(n13686) );
  NANDN U13913 ( .A(n13687), .B(n13686), .Z(n13688) );
  AND U13914 ( .A(n13689), .B(n13688), .Z(n13690) );
  NAND U13915 ( .A(n13691), .B(n13690), .Z(n13692) );
  NAND U13916 ( .A(n13693), .B(n13692), .Z(n13695) );
  NAND U13917 ( .A(n13695), .B(n13694), .Z(n13696) );
  NANDN U13918 ( .A(n13697), .B(n13696), .Z(n13698) );
  AND U13919 ( .A(n13699), .B(n13698), .Z(n13701) );
  NANDN U13920 ( .A(n13701), .B(n13700), .Z(n13702) );
  NANDN U13921 ( .A(n13703), .B(n13702), .Z(n13705) );
  NAND U13922 ( .A(n13705), .B(n13704), .Z(n13706) );
  NANDN U13923 ( .A(n13707), .B(n13706), .Z(n13708) );
  NANDN U13924 ( .A(n13709), .B(n13708), .Z(n13711) );
  ANDN U13925 ( .B(n13711), .A(n13710), .Z(n13713) );
  NANDN U13926 ( .A(n13713), .B(n13712), .Z(n13715) );
  NAND U13927 ( .A(n13715), .B(n13714), .Z(n13717) );
  NAND U13928 ( .A(n13717), .B(n13716), .Z(n13718) );
  NANDN U13929 ( .A(n13719), .B(n13718), .Z(n13721) );
  NAND U13930 ( .A(n13721), .B(n13720), .Z(n13723) );
  ANDN U13931 ( .B(n13723), .A(n13722), .Z(n13725) );
  NANDN U13932 ( .A(n13725), .B(n13724), .Z(n13726) );
  NANDN U13933 ( .A(n13727), .B(n13726), .Z(n13728) );
  NANDN U13934 ( .A(n13729), .B(n13728), .Z(n13731) );
  NANDN U13935 ( .A(n13731), .B(n13730), .Z(n13732) );
  AND U13936 ( .A(n13733), .B(n13732), .Z(n13734) );
  OR U13937 ( .A(n13735), .B(n13734), .Z(n13736) );
  NANDN U13938 ( .A(n13737), .B(n13736), .Z(n13738) );
  NANDN U13939 ( .A(n13739), .B(n13738), .Z(n13740) );
  NANDN U13940 ( .A(n13741), .B(n13740), .Z(n13743) );
  NAND U13941 ( .A(n13743), .B(n13742), .Z(n13744) );
  AND U13942 ( .A(n13745), .B(n13744), .Z(n13746) );
  OR U13943 ( .A(n13747), .B(n13746), .Z(n13748) );
  NANDN U13944 ( .A(n13749), .B(n13748), .Z(n13750) );
  NANDN U13945 ( .A(n13751), .B(n13750), .Z(n13753) );
  NAND U13946 ( .A(n13753), .B(n13752), .Z(n13755) );
  ANDN U13947 ( .B(n13755), .A(n13754), .Z(n13757) );
  NANDN U13948 ( .A(n13757), .B(n13756), .Z(n13758) );
  NAND U13949 ( .A(n13759), .B(n13758), .Z(n13760) );
  NAND U13950 ( .A(n13761), .B(n13760), .Z(n13762) );
  NANDN U13951 ( .A(n13763), .B(n13762), .Z(n13764) );
  AND U13952 ( .A(n13765), .B(n13764), .Z(n13766) );
  OR U13953 ( .A(n13767), .B(n13766), .Z(n13768) );
  AND U13954 ( .A(n13769), .B(n13768), .Z(n13771) );
  NANDN U13955 ( .A(n13771), .B(n13770), .Z(n13773) );
  NAND U13956 ( .A(n13773), .B(n13772), .Z(n13775) );
  ANDN U13957 ( .B(n13775), .A(n13774), .Z(n13777) );
  NANDN U13958 ( .A(n13777), .B(n13776), .Z(n13778) );
  NANDN U13959 ( .A(n13779), .B(n13778), .Z(n13780) );
  NANDN U13960 ( .A(n13781), .B(n13780), .Z(n13783) );
  ANDN U13961 ( .B(n13783), .A(n13782), .Z(n13785) );
  NANDN U13962 ( .A(n13785), .B(n13784), .Z(n13787) );
  ANDN U13963 ( .B(n13787), .A(n13786), .Z(n13789) );
  OR U13964 ( .A(n13789), .B(n13788), .Z(n13790) );
  NANDN U13965 ( .A(n13791), .B(n13790), .Z(n13792) );
  AND U13966 ( .A(n13793), .B(n13792), .Z(n13794) );
  OR U13967 ( .A(n13795), .B(n13794), .Z(n13796) );
  AND U13968 ( .A(n13797), .B(n13796), .Z(n13799) );
  NANDN U13969 ( .A(n13799), .B(n13798), .Z(n13801) );
  NAND U13970 ( .A(n13801), .B(n13800), .Z(n13803) );
  NAND U13971 ( .A(n13803), .B(n13802), .Z(n13804) );
  NANDN U13972 ( .A(n13805), .B(n13804), .Z(n13807) );
  NANDN U13973 ( .A(n13825), .B(n13824), .Z(n13826) );
  NANDN U13974 ( .A(n13827), .B(n13826), .Z(n13828) );
  AND U13975 ( .A(n13829), .B(n13828), .Z(n13831) );
  OR U13976 ( .A(n13831), .B(n13830), .Z(n13833) );
  NAND U13977 ( .A(n13833), .B(n13832), .Z(n13834) );
  NANDN U13978 ( .A(n13835), .B(n13834), .Z(n13836) );
  AND U13979 ( .A(n13837), .B(n13836), .Z(n13839) );
  NANDN U13980 ( .A(n13839), .B(n13838), .Z(n13841) );
  NAND U13981 ( .A(n13841), .B(n13840), .Z(n13843) );
  NAND U13982 ( .A(n13843), .B(n13842), .Z(n13845) );
  NAND U13983 ( .A(n13845), .B(n13844), .Z(n13847) );
  NAND U13984 ( .A(n13847), .B(n13846), .Z(n13849) );
  ANDN U13985 ( .B(n13849), .A(n13848), .Z(n13850) );
  OR U13986 ( .A(n13851), .B(n13850), .Z(n13853) );
  ANDN U13987 ( .B(n13853), .A(n13852), .Z(n13854) );
  OR U13988 ( .A(n13855), .B(n13854), .Z(n13856) );
  AND U13989 ( .A(n13857), .B(n13856), .Z(n13858) );
  OR U13990 ( .A(n13859), .B(n13858), .Z(n13860) );
  AND U13991 ( .A(n13861), .B(n13860), .Z(n13862) );
  OR U13992 ( .A(n13863), .B(n13862), .Z(n13864) );
  NANDN U13993 ( .A(n13865), .B(n13864), .Z(n13867) );
  NAND U13994 ( .A(n13867), .B(n13866), .Z(n13869) );
  ANDN U13995 ( .B(n13869), .A(n13868), .Z(n13871) );
  NANDN U13996 ( .A(n13871), .B(n13870), .Z(n13872) );
  AND U13997 ( .A(n13873), .B(n13872), .Z(n13874) );
  OR U13998 ( .A(n13875), .B(n13874), .Z(n13876) );
  NANDN U13999 ( .A(n13877), .B(n13876), .Z(n13879) );
  NAND U14000 ( .A(n13879), .B(n13878), .Z(n13881) );
  ANDN U14001 ( .B(n13881), .A(n13880), .Z(n13883) );
  NANDN U14002 ( .A(n13883), .B(n13882), .Z(n13884) );
  NANDN U14003 ( .A(n13885), .B(n13884), .Z(n13887) );
  NAND U14004 ( .A(n13887), .B(n13886), .Z(n13889) );
  NAND U14005 ( .A(n13889), .B(n13888), .Z(n13890) );
  NANDN U14006 ( .A(n13891), .B(n13890), .Z(n13892) );
  AND U14007 ( .A(n13893), .B(n13892), .Z(n13899) );
  NANDN U14008 ( .A(y[1950]), .B(n13894), .Z(n13897) );
  XNOR U14009 ( .A(n13894), .B(y[1950]), .Z(n13895) );
  NAND U14010 ( .A(n13895), .B(x[1950]), .Z(n13896) );
  NAND U14011 ( .A(n13897), .B(n13896), .Z(n13898) );
  AND U14012 ( .A(n13899), .B(n13898), .Z(n13901) );
  NAND U14013 ( .A(n13921), .B(n13920), .Z(n13922) );
  AND U14014 ( .A(n13923), .B(n13922), .Z(n13925) );
  NANDN U14015 ( .A(n13925), .B(n13924), .Z(n13926) );
  NANDN U14016 ( .A(n13927), .B(n13926), .Z(n13929) );
  NAND U14017 ( .A(n13929), .B(n13928), .Z(n13931) );
  NAND U14018 ( .A(n13931), .B(n13930), .Z(n13932) );
  NANDN U14019 ( .A(n13933), .B(n13932), .Z(n13935) );
  ANDN U14020 ( .B(n13935), .A(n13934), .Z(n13936) );
  NAND U14021 ( .A(n13937), .B(n13936), .Z(n13938) );
  NAND U14022 ( .A(n13939), .B(n13938), .Z(n13940) );
  AND U14023 ( .A(n13941), .B(n13940), .Z(n13943) );
  NANDN U14024 ( .A(n13943), .B(n13942), .Z(n13945) );
  ANDN U14025 ( .B(n13945), .A(n13944), .Z(n13946) );
  OR U14026 ( .A(n13947), .B(n13946), .Z(n13948) );
  NANDN U14027 ( .A(n13949), .B(n13948), .Z(n13951) );
  NAND U14028 ( .A(n13951), .B(n13950), .Z(n13953) );
  NAND U14029 ( .A(n13953), .B(n13952), .Z(n13955) );
  NAND U14030 ( .A(n13955), .B(n13954), .Z(n13956) );
  NAND U14031 ( .A(n13975), .B(n13974), .Z(n13976) );
  NANDN U14032 ( .A(n13977), .B(n13976), .Z(n13978) );
  NANDN U14033 ( .A(n13979), .B(n13978), .Z(n13980) );
  AND U14034 ( .A(n13981), .B(n13980), .Z(n13982) );
  OR U14035 ( .A(n13983), .B(n13982), .Z(n13985) );
  ANDN U14036 ( .B(n13985), .A(n13984), .Z(n13987) );
  NANDN U14037 ( .A(n13987), .B(n13986), .Z(n13989) );
  ANDN U14038 ( .B(n13989), .A(n13988), .Z(n13991) );
  NANDN U14039 ( .A(n13991), .B(n13990), .Z(n13993) );
  ANDN U14040 ( .B(n13993), .A(n13992), .Z(n13995) );
  NANDN U14041 ( .A(n13995), .B(n13994), .Z(n13996) );
  AND U14042 ( .A(n13997), .B(n13996), .Z(n13999) );
  NANDN U14043 ( .A(n13999), .B(n13998), .Z(n14001) );
  ANDN U14044 ( .B(n14001), .A(n14000), .Z(n14002) );
  OR U14045 ( .A(n14003), .B(n14002), .Z(n14004) );
  NANDN U14046 ( .A(n14005), .B(n14004), .Z(n14006) );
  NANDN U14047 ( .A(n14007), .B(n14006), .Z(n14008) );
  AND U14048 ( .A(n14009), .B(n14008), .Z(n14010) );
  OR U14049 ( .A(n14011), .B(n14010), .Z(n14012) );
  NANDN U14050 ( .A(n14013), .B(n14012), .Z(n14015) );
  NAND U14051 ( .A(n14015), .B(n14014), .Z(n14017) );
  NAND U14052 ( .A(n14017), .B(n14016), .Z(n14019) );
  NAND U14053 ( .A(n14019), .B(n14018), .Z(n14020) );
  NANDN U14054 ( .A(n14021), .B(n14020), .Z(n14023) );
  ANDN U14055 ( .B(n14023), .A(n14022), .Z(n14025) );
  NANDN U14056 ( .A(n14025), .B(n14024), .Z(n14026) );
  AND U14057 ( .A(n14027), .B(n14026), .Z(n14029) );
  NANDN U14058 ( .A(n14029), .B(n14028), .Z(n14031) );
  ANDN U14059 ( .B(n14031), .A(n14030), .Z(n14032) );
  OR U14060 ( .A(n14033), .B(n14032), .Z(n14034) );
  AND U14061 ( .A(n14035), .B(n14034), .Z(n14039) );
  AND U14062 ( .A(n14037), .B(n14036), .Z(n14038) );
  NANDN U14063 ( .A(n14039), .B(n14038), .Z(n14041) );
  NAND U14064 ( .A(n14041), .B(n14040), .Z(n14042) );
  NANDN U14065 ( .A(n14043), .B(n14042), .Z(n14045) );
  NAND U14066 ( .A(n14045), .B(n14044), .Z(n14047) );
  NAND U14067 ( .A(n14047), .B(n14046), .Z(n14049) );
  ANDN U14068 ( .B(n14049), .A(n14048), .Z(n14050) );
  OR U14069 ( .A(n14051), .B(n14050), .Z(n14052) );
  NANDN U14070 ( .A(n14053), .B(n14052), .Z(n14054) );
  NANDN U14071 ( .A(n14055), .B(n14054), .Z(n14056) );
  OR U14072 ( .A(n14057), .B(n14056), .Z(n14058) );
  AND U14073 ( .A(n14059), .B(n14058), .Z(n14060) );
  OR U14074 ( .A(n14061), .B(n14060), .Z(n14063) );
  ANDN U14075 ( .B(n14063), .A(n14062), .Z(n14064) );
  OR U14076 ( .A(n14065), .B(n14064), .Z(n14071) );
  NANDN U14077 ( .A(n14067), .B(n14066), .Z(n14069) );
  ANDN U14078 ( .B(n14069), .A(n14068), .Z(n14070) );
  NAND U14079 ( .A(n14071), .B(n14070), .Z(n14072) );
  NANDN U14080 ( .A(n14073), .B(n14072), .Z(n14075) );
  ANDN U14081 ( .B(n14075), .A(n14074), .Z(n14076) );
  NANDN U14082 ( .A(n14077), .B(n14076), .Z(n14079) );
  NANDN U14083 ( .A(g), .B(n14077), .Z(n14078) );
  AND U14084 ( .A(n14079), .B(n14078), .Z(n4) );
endmodule

