
module mult_N256_CC64 ( clk, rst, a, b, c );
  input [255:0] a;
  input [3:0] b;
  output [511:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008;
  wire   [511:0] sreg;

  DFF \sreg_reg[507]  ( .D(c[511]), .CLK(clk), .RST(rst), .Q(sreg[507]) );
  DFF \sreg_reg[506]  ( .D(c[510]), .CLK(clk), .RST(rst), .Q(sreg[506]) );
  DFF \sreg_reg[505]  ( .D(c[509]), .CLK(clk), .RST(rst), .Q(sreg[505]) );
  DFF \sreg_reg[504]  ( .D(c[508]), .CLK(clk), .RST(rst), .Q(sreg[504]) );
  DFF \sreg_reg[503]  ( .D(c[507]), .CLK(clk), .RST(rst), .Q(sreg[503]) );
  DFF \sreg_reg[502]  ( .D(c[506]), .CLK(clk), .RST(rst), .Q(sreg[502]) );
  DFF \sreg_reg[501]  ( .D(c[505]), .CLK(clk), .RST(rst), .Q(sreg[501]) );
  DFF \sreg_reg[500]  ( .D(c[504]), .CLK(clk), .RST(rst), .Q(sreg[500]) );
  DFF \sreg_reg[499]  ( .D(c[503]), .CLK(clk), .RST(rst), .Q(sreg[499]) );
  DFF \sreg_reg[498]  ( .D(c[502]), .CLK(clk), .RST(rst), .Q(sreg[498]) );
  DFF \sreg_reg[497]  ( .D(c[501]), .CLK(clk), .RST(rst), .Q(sreg[497]) );
  DFF \sreg_reg[496]  ( .D(c[500]), .CLK(clk), .RST(rst), .Q(sreg[496]) );
  DFF \sreg_reg[495]  ( .D(c[499]), .CLK(clk), .RST(rst), .Q(sreg[495]) );
  DFF \sreg_reg[494]  ( .D(c[498]), .CLK(clk), .RST(rst), .Q(sreg[494]) );
  DFF \sreg_reg[493]  ( .D(c[497]), .CLK(clk), .RST(rst), .Q(sreg[493]) );
  DFF \sreg_reg[492]  ( .D(c[496]), .CLK(clk), .RST(rst), .Q(sreg[492]) );
  DFF \sreg_reg[491]  ( .D(c[495]), .CLK(clk), .RST(rst), .Q(sreg[491]) );
  DFF \sreg_reg[490]  ( .D(c[494]), .CLK(clk), .RST(rst), .Q(sreg[490]) );
  DFF \sreg_reg[489]  ( .D(c[493]), .CLK(clk), .RST(rst), .Q(sreg[489]) );
  DFF \sreg_reg[488]  ( .D(c[492]), .CLK(clk), .RST(rst), .Q(sreg[488]) );
  DFF \sreg_reg[487]  ( .D(c[491]), .CLK(clk), .RST(rst), .Q(sreg[487]) );
  DFF \sreg_reg[486]  ( .D(c[490]), .CLK(clk), .RST(rst), .Q(sreg[486]) );
  DFF \sreg_reg[485]  ( .D(c[489]), .CLK(clk), .RST(rst), .Q(sreg[485]) );
  DFF \sreg_reg[484]  ( .D(c[488]), .CLK(clk), .RST(rst), .Q(sreg[484]) );
  DFF \sreg_reg[483]  ( .D(c[487]), .CLK(clk), .RST(rst), .Q(sreg[483]) );
  DFF \sreg_reg[482]  ( .D(c[486]), .CLK(clk), .RST(rst), .Q(sreg[482]) );
  DFF \sreg_reg[481]  ( .D(c[485]), .CLK(clk), .RST(rst), .Q(sreg[481]) );
  DFF \sreg_reg[480]  ( .D(c[484]), .CLK(clk), .RST(rst), .Q(sreg[480]) );
  DFF \sreg_reg[479]  ( .D(c[483]), .CLK(clk), .RST(rst), .Q(sreg[479]) );
  DFF \sreg_reg[478]  ( .D(c[482]), .CLK(clk), .RST(rst), .Q(sreg[478]) );
  DFF \sreg_reg[477]  ( .D(c[481]), .CLK(clk), .RST(rst), .Q(sreg[477]) );
  DFF \sreg_reg[476]  ( .D(c[480]), .CLK(clk), .RST(rst), .Q(sreg[476]) );
  DFF \sreg_reg[475]  ( .D(c[479]), .CLK(clk), .RST(rst), .Q(sreg[475]) );
  DFF \sreg_reg[474]  ( .D(c[478]), .CLK(clk), .RST(rst), .Q(sreg[474]) );
  DFF \sreg_reg[473]  ( .D(c[477]), .CLK(clk), .RST(rst), .Q(sreg[473]) );
  DFF \sreg_reg[472]  ( .D(c[476]), .CLK(clk), .RST(rst), .Q(sreg[472]) );
  DFF \sreg_reg[471]  ( .D(c[475]), .CLK(clk), .RST(rst), .Q(sreg[471]) );
  DFF \sreg_reg[470]  ( .D(c[474]), .CLK(clk), .RST(rst), .Q(sreg[470]) );
  DFF \sreg_reg[469]  ( .D(c[473]), .CLK(clk), .RST(rst), .Q(sreg[469]) );
  DFF \sreg_reg[468]  ( .D(c[472]), .CLK(clk), .RST(rst), .Q(sreg[468]) );
  DFF \sreg_reg[467]  ( .D(c[471]), .CLK(clk), .RST(rst), .Q(sreg[467]) );
  DFF \sreg_reg[466]  ( .D(c[470]), .CLK(clk), .RST(rst), .Q(sreg[466]) );
  DFF \sreg_reg[465]  ( .D(c[469]), .CLK(clk), .RST(rst), .Q(sreg[465]) );
  DFF \sreg_reg[464]  ( .D(c[468]), .CLK(clk), .RST(rst), .Q(sreg[464]) );
  DFF \sreg_reg[463]  ( .D(c[467]), .CLK(clk), .RST(rst), .Q(sreg[463]) );
  DFF \sreg_reg[462]  ( .D(c[466]), .CLK(clk), .RST(rst), .Q(sreg[462]) );
  DFF \sreg_reg[461]  ( .D(c[465]), .CLK(clk), .RST(rst), .Q(sreg[461]) );
  DFF \sreg_reg[460]  ( .D(c[464]), .CLK(clk), .RST(rst), .Q(sreg[460]) );
  DFF \sreg_reg[459]  ( .D(c[463]), .CLK(clk), .RST(rst), .Q(sreg[459]) );
  DFF \sreg_reg[458]  ( .D(c[462]), .CLK(clk), .RST(rst), .Q(sreg[458]) );
  DFF \sreg_reg[457]  ( .D(c[461]), .CLK(clk), .RST(rst), .Q(sreg[457]) );
  DFF \sreg_reg[456]  ( .D(c[460]), .CLK(clk), .RST(rst), .Q(sreg[456]) );
  DFF \sreg_reg[455]  ( .D(c[459]), .CLK(clk), .RST(rst), .Q(sreg[455]) );
  DFF \sreg_reg[454]  ( .D(c[458]), .CLK(clk), .RST(rst), .Q(sreg[454]) );
  DFF \sreg_reg[453]  ( .D(c[457]), .CLK(clk), .RST(rst), .Q(sreg[453]) );
  DFF \sreg_reg[452]  ( .D(c[456]), .CLK(clk), .RST(rst), .Q(sreg[452]) );
  DFF \sreg_reg[451]  ( .D(c[455]), .CLK(clk), .RST(rst), .Q(sreg[451]) );
  DFF \sreg_reg[450]  ( .D(c[454]), .CLK(clk), .RST(rst), .Q(sreg[450]) );
  DFF \sreg_reg[449]  ( .D(c[453]), .CLK(clk), .RST(rst), .Q(sreg[449]) );
  DFF \sreg_reg[448]  ( .D(c[452]), .CLK(clk), .RST(rst), .Q(sreg[448]) );
  DFF \sreg_reg[447]  ( .D(c[451]), .CLK(clk), .RST(rst), .Q(sreg[447]) );
  DFF \sreg_reg[446]  ( .D(c[450]), .CLK(clk), .RST(rst), .Q(sreg[446]) );
  DFF \sreg_reg[445]  ( .D(c[449]), .CLK(clk), .RST(rst), .Q(sreg[445]) );
  DFF \sreg_reg[444]  ( .D(c[448]), .CLK(clk), .RST(rst), .Q(sreg[444]) );
  DFF \sreg_reg[443]  ( .D(c[447]), .CLK(clk), .RST(rst), .Q(sreg[443]) );
  DFF \sreg_reg[442]  ( .D(c[446]), .CLK(clk), .RST(rst), .Q(sreg[442]) );
  DFF \sreg_reg[441]  ( .D(c[445]), .CLK(clk), .RST(rst), .Q(sreg[441]) );
  DFF \sreg_reg[440]  ( .D(c[444]), .CLK(clk), .RST(rst), .Q(sreg[440]) );
  DFF \sreg_reg[439]  ( .D(c[443]), .CLK(clk), .RST(rst), .Q(sreg[439]) );
  DFF \sreg_reg[438]  ( .D(c[442]), .CLK(clk), .RST(rst), .Q(sreg[438]) );
  DFF \sreg_reg[437]  ( .D(c[441]), .CLK(clk), .RST(rst), .Q(sreg[437]) );
  DFF \sreg_reg[436]  ( .D(c[440]), .CLK(clk), .RST(rst), .Q(sreg[436]) );
  DFF \sreg_reg[435]  ( .D(c[439]), .CLK(clk), .RST(rst), .Q(sreg[435]) );
  DFF \sreg_reg[434]  ( .D(c[438]), .CLK(clk), .RST(rst), .Q(sreg[434]) );
  DFF \sreg_reg[433]  ( .D(c[437]), .CLK(clk), .RST(rst), .Q(sreg[433]) );
  DFF \sreg_reg[432]  ( .D(c[436]), .CLK(clk), .RST(rst), .Q(sreg[432]) );
  DFF \sreg_reg[431]  ( .D(c[435]), .CLK(clk), .RST(rst), .Q(sreg[431]) );
  DFF \sreg_reg[430]  ( .D(c[434]), .CLK(clk), .RST(rst), .Q(sreg[430]) );
  DFF \sreg_reg[429]  ( .D(c[433]), .CLK(clk), .RST(rst), .Q(sreg[429]) );
  DFF \sreg_reg[428]  ( .D(c[432]), .CLK(clk), .RST(rst), .Q(sreg[428]) );
  DFF \sreg_reg[427]  ( .D(c[431]), .CLK(clk), .RST(rst), .Q(sreg[427]) );
  DFF \sreg_reg[426]  ( .D(c[430]), .CLK(clk), .RST(rst), .Q(sreg[426]) );
  DFF \sreg_reg[425]  ( .D(c[429]), .CLK(clk), .RST(rst), .Q(sreg[425]) );
  DFF \sreg_reg[424]  ( .D(c[428]), .CLK(clk), .RST(rst), .Q(sreg[424]) );
  DFF \sreg_reg[423]  ( .D(c[427]), .CLK(clk), .RST(rst), .Q(sreg[423]) );
  DFF \sreg_reg[422]  ( .D(c[426]), .CLK(clk), .RST(rst), .Q(sreg[422]) );
  DFF \sreg_reg[421]  ( .D(c[425]), .CLK(clk), .RST(rst), .Q(sreg[421]) );
  DFF \sreg_reg[420]  ( .D(c[424]), .CLK(clk), .RST(rst), .Q(sreg[420]) );
  DFF \sreg_reg[419]  ( .D(c[423]), .CLK(clk), .RST(rst), .Q(sreg[419]) );
  DFF \sreg_reg[418]  ( .D(c[422]), .CLK(clk), .RST(rst), .Q(sreg[418]) );
  DFF \sreg_reg[417]  ( .D(c[421]), .CLK(clk), .RST(rst), .Q(sreg[417]) );
  DFF \sreg_reg[416]  ( .D(c[420]), .CLK(clk), .RST(rst), .Q(sreg[416]) );
  DFF \sreg_reg[415]  ( .D(c[419]), .CLK(clk), .RST(rst), .Q(sreg[415]) );
  DFF \sreg_reg[414]  ( .D(c[418]), .CLK(clk), .RST(rst), .Q(sreg[414]) );
  DFF \sreg_reg[413]  ( .D(c[417]), .CLK(clk), .RST(rst), .Q(sreg[413]) );
  DFF \sreg_reg[412]  ( .D(c[416]), .CLK(clk), .RST(rst), .Q(sreg[412]) );
  DFF \sreg_reg[411]  ( .D(c[415]), .CLK(clk), .RST(rst), .Q(sreg[411]) );
  DFF \sreg_reg[410]  ( .D(c[414]), .CLK(clk), .RST(rst), .Q(sreg[410]) );
  DFF \sreg_reg[409]  ( .D(c[413]), .CLK(clk), .RST(rst), .Q(sreg[409]) );
  DFF \sreg_reg[408]  ( .D(c[412]), .CLK(clk), .RST(rst), .Q(sreg[408]) );
  DFF \sreg_reg[407]  ( .D(c[411]), .CLK(clk), .RST(rst), .Q(sreg[407]) );
  DFF \sreg_reg[406]  ( .D(c[410]), .CLK(clk), .RST(rst), .Q(sreg[406]) );
  DFF \sreg_reg[405]  ( .D(c[409]), .CLK(clk), .RST(rst), .Q(sreg[405]) );
  DFF \sreg_reg[404]  ( .D(c[408]), .CLK(clk), .RST(rst), .Q(sreg[404]) );
  DFF \sreg_reg[403]  ( .D(c[407]), .CLK(clk), .RST(rst), .Q(sreg[403]) );
  DFF \sreg_reg[402]  ( .D(c[406]), .CLK(clk), .RST(rst), .Q(sreg[402]) );
  DFF \sreg_reg[401]  ( .D(c[405]), .CLK(clk), .RST(rst), .Q(sreg[401]) );
  DFF \sreg_reg[400]  ( .D(c[404]), .CLK(clk), .RST(rst), .Q(sreg[400]) );
  DFF \sreg_reg[399]  ( .D(c[403]), .CLK(clk), .RST(rst), .Q(sreg[399]) );
  DFF \sreg_reg[398]  ( .D(c[402]), .CLK(clk), .RST(rst), .Q(sreg[398]) );
  DFF \sreg_reg[397]  ( .D(c[401]), .CLK(clk), .RST(rst), .Q(sreg[397]) );
  DFF \sreg_reg[396]  ( .D(c[400]), .CLK(clk), .RST(rst), .Q(sreg[396]) );
  DFF \sreg_reg[395]  ( .D(c[399]), .CLK(clk), .RST(rst), .Q(sreg[395]) );
  DFF \sreg_reg[394]  ( .D(c[398]), .CLK(clk), .RST(rst), .Q(sreg[394]) );
  DFF \sreg_reg[393]  ( .D(c[397]), .CLK(clk), .RST(rst), .Q(sreg[393]) );
  DFF \sreg_reg[392]  ( .D(c[396]), .CLK(clk), .RST(rst), .Q(sreg[392]) );
  DFF \sreg_reg[391]  ( .D(c[395]), .CLK(clk), .RST(rst), .Q(sreg[391]) );
  DFF \sreg_reg[390]  ( .D(c[394]), .CLK(clk), .RST(rst), .Q(sreg[390]) );
  DFF \sreg_reg[389]  ( .D(c[393]), .CLK(clk), .RST(rst), .Q(sreg[389]) );
  DFF \sreg_reg[388]  ( .D(c[392]), .CLK(clk), .RST(rst), .Q(sreg[388]) );
  DFF \sreg_reg[387]  ( .D(c[391]), .CLK(clk), .RST(rst), .Q(sreg[387]) );
  DFF \sreg_reg[386]  ( .D(c[390]), .CLK(clk), .RST(rst), .Q(sreg[386]) );
  DFF \sreg_reg[385]  ( .D(c[389]), .CLK(clk), .RST(rst), .Q(sreg[385]) );
  DFF \sreg_reg[384]  ( .D(c[388]), .CLK(clk), .RST(rst), .Q(sreg[384]) );
  DFF \sreg_reg[383]  ( .D(c[387]), .CLK(clk), .RST(rst), .Q(sreg[383]) );
  DFF \sreg_reg[382]  ( .D(c[386]), .CLK(clk), .RST(rst), .Q(sreg[382]) );
  DFF \sreg_reg[381]  ( .D(c[385]), .CLK(clk), .RST(rst), .Q(sreg[381]) );
  DFF \sreg_reg[380]  ( .D(c[384]), .CLK(clk), .RST(rst), .Q(sreg[380]) );
  DFF \sreg_reg[379]  ( .D(c[383]), .CLK(clk), .RST(rst), .Q(sreg[379]) );
  DFF \sreg_reg[378]  ( .D(c[382]), .CLK(clk), .RST(rst), .Q(sreg[378]) );
  DFF \sreg_reg[377]  ( .D(c[381]), .CLK(clk), .RST(rst), .Q(sreg[377]) );
  DFF \sreg_reg[376]  ( .D(c[380]), .CLK(clk), .RST(rst), .Q(sreg[376]) );
  DFF \sreg_reg[375]  ( .D(c[379]), .CLK(clk), .RST(rst), .Q(sreg[375]) );
  DFF \sreg_reg[374]  ( .D(c[378]), .CLK(clk), .RST(rst), .Q(sreg[374]) );
  DFF \sreg_reg[373]  ( .D(c[377]), .CLK(clk), .RST(rst), .Q(sreg[373]) );
  DFF \sreg_reg[372]  ( .D(c[376]), .CLK(clk), .RST(rst), .Q(sreg[372]) );
  DFF \sreg_reg[371]  ( .D(c[375]), .CLK(clk), .RST(rst), .Q(sreg[371]) );
  DFF \sreg_reg[370]  ( .D(c[374]), .CLK(clk), .RST(rst), .Q(sreg[370]) );
  DFF \sreg_reg[369]  ( .D(c[373]), .CLK(clk), .RST(rst), .Q(sreg[369]) );
  DFF \sreg_reg[368]  ( .D(c[372]), .CLK(clk), .RST(rst), .Q(sreg[368]) );
  DFF \sreg_reg[367]  ( .D(c[371]), .CLK(clk), .RST(rst), .Q(sreg[367]) );
  DFF \sreg_reg[366]  ( .D(c[370]), .CLK(clk), .RST(rst), .Q(sreg[366]) );
  DFF \sreg_reg[365]  ( .D(c[369]), .CLK(clk), .RST(rst), .Q(sreg[365]) );
  DFF \sreg_reg[364]  ( .D(c[368]), .CLK(clk), .RST(rst), .Q(sreg[364]) );
  DFF \sreg_reg[363]  ( .D(c[367]), .CLK(clk), .RST(rst), .Q(sreg[363]) );
  DFF \sreg_reg[362]  ( .D(c[366]), .CLK(clk), .RST(rst), .Q(sreg[362]) );
  DFF \sreg_reg[361]  ( .D(c[365]), .CLK(clk), .RST(rst), .Q(sreg[361]) );
  DFF \sreg_reg[360]  ( .D(c[364]), .CLK(clk), .RST(rst), .Q(sreg[360]) );
  DFF \sreg_reg[359]  ( .D(c[363]), .CLK(clk), .RST(rst), .Q(sreg[359]) );
  DFF \sreg_reg[358]  ( .D(c[362]), .CLK(clk), .RST(rst), .Q(sreg[358]) );
  DFF \sreg_reg[357]  ( .D(c[361]), .CLK(clk), .RST(rst), .Q(sreg[357]) );
  DFF \sreg_reg[356]  ( .D(c[360]), .CLK(clk), .RST(rst), .Q(sreg[356]) );
  DFF \sreg_reg[355]  ( .D(c[359]), .CLK(clk), .RST(rst), .Q(sreg[355]) );
  DFF \sreg_reg[354]  ( .D(c[358]), .CLK(clk), .RST(rst), .Q(sreg[354]) );
  DFF \sreg_reg[353]  ( .D(c[357]), .CLK(clk), .RST(rst), .Q(sreg[353]) );
  DFF \sreg_reg[352]  ( .D(c[356]), .CLK(clk), .RST(rst), .Q(sreg[352]) );
  DFF \sreg_reg[351]  ( .D(c[355]), .CLK(clk), .RST(rst), .Q(sreg[351]) );
  DFF \sreg_reg[350]  ( .D(c[354]), .CLK(clk), .RST(rst), .Q(sreg[350]) );
  DFF \sreg_reg[349]  ( .D(c[353]), .CLK(clk), .RST(rst), .Q(sreg[349]) );
  DFF \sreg_reg[348]  ( .D(c[352]), .CLK(clk), .RST(rst), .Q(sreg[348]) );
  DFF \sreg_reg[347]  ( .D(c[351]), .CLK(clk), .RST(rst), .Q(sreg[347]) );
  DFF \sreg_reg[346]  ( .D(c[350]), .CLK(clk), .RST(rst), .Q(sreg[346]) );
  DFF \sreg_reg[345]  ( .D(c[349]), .CLK(clk), .RST(rst), .Q(sreg[345]) );
  DFF \sreg_reg[344]  ( .D(c[348]), .CLK(clk), .RST(rst), .Q(sreg[344]) );
  DFF \sreg_reg[343]  ( .D(c[347]), .CLK(clk), .RST(rst), .Q(sreg[343]) );
  DFF \sreg_reg[342]  ( .D(c[346]), .CLK(clk), .RST(rst), .Q(sreg[342]) );
  DFF \sreg_reg[341]  ( .D(c[345]), .CLK(clk), .RST(rst), .Q(sreg[341]) );
  DFF \sreg_reg[340]  ( .D(c[344]), .CLK(clk), .RST(rst), .Q(sreg[340]) );
  DFF \sreg_reg[339]  ( .D(c[343]), .CLK(clk), .RST(rst), .Q(sreg[339]) );
  DFF \sreg_reg[338]  ( .D(c[342]), .CLK(clk), .RST(rst), .Q(sreg[338]) );
  DFF \sreg_reg[337]  ( .D(c[341]), .CLK(clk), .RST(rst), .Q(sreg[337]) );
  DFF \sreg_reg[336]  ( .D(c[340]), .CLK(clk), .RST(rst), .Q(sreg[336]) );
  DFF \sreg_reg[335]  ( .D(c[339]), .CLK(clk), .RST(rst), .Q(sreg[335]) );
  DFF \sreg_reg[334]  ( .D(c[338]), .CLK(clk), .RST(rst), .Q(sreg[334]) );
  DFF \sreg_reg[333]  ( .D(c[337]), .CLK(clk), .RST(rst), .Q(sreg[333]) );
  DFF \sreg_reg[332]  ( .D(c[336]), .CLK(clk), .RST(rst), .Q(sreg[332]) );
  DFF \sreg_reg[331]  ( .D(c[335]), .CLK(clk), .RST(rst), .Q(sreg[331]) );
  DFF \sreg_reg[330]  ( .D(c[334]), .CLK(clk), .RST(rst), .Q(sreg[330]) );
  DFF \sreg_reg[329]  ( .D(c[333]), .CLK(clk), .RST(rst), .Q(sreg[329]) );
  DFF \sreg_reg[328]  ( .D(c[332]), .CLK(clk), .RST(rst), .Q(sreg[328]) );
  DFF \sreg_reg[327]  ( .D(c[331]), .CLK(clk), .RST(rst), .Q(sreg[327]) );
  DFF \sreg_reg[326]  ( .D(c[330]), .CLK(clk), .RST(rst), .Q(sreg[326]) );
  DFF \sreg_reg[325]  ( .D(c[329]), .CLK(clk), .RST(rst), .Q(sreg[325]) );
  DFF \sreg_reg[324]  ( .D(c[328]), .CLK(clk), .RST(rst), .Q(sreg[324]) );
  DFF \sreg_reg[323]  ( .D(c[327]), .CLK(clk), .RST(rst), .Q(sreg[323]) );
  DFF \sreg_reg[322]  ( .D(c[326]), .CLK(clk), .RST(rst), .Q(sreg[322]) );
  DFF \sreg_reg[321]  ( .D(c[325]), .CLK(clk), .RST(rst), .Q(sreg[321]) );
  DFF \sreg_reg[320]  ( .D(c[324]), .CLK(clk), .RST(rst), .Q(sreg[320]) );
  DFF \sreg_reg[319]  ( .D(c[323]), .CLK(clk), .RST(rst), .Q(sreg[319]) );
  DFF \sreg_reg[318]  ( .D(c[322]), .CLK(clk), .RST(rst), .Q(sreg[318]) );
  DFF \sreg_reg[317]  ( .D(c[321]), .CLK(clk), .RST(rst), .Q(sreg[317]) );
  DFF \sreg_reg[316]  ( .D(c[320]), .CLK(clk), .RST(rst), .Q(sreg[316]) );
  DFF \sreg_reg[315]  ( .D(c[319]), .CLK(clk), .RST(rst), .Q(sreg[315]) );
  DFF \sreg_reg[314]  ( .D(c[318]), .CLK(clk), .RST(rst), .Q(sreg[314]) );
  DFF \sreg_reg[313]  ( .D(c[317]), .CLK(clk), .RST(rst), .Q(sreg[313]) );
  DFF \sreg_reg[312]  ( .D(c[316]), .CLK(clk), .RST(rst), .Q(sreg[312]) );
  DFF \sreg_reg[311]  ( .D(c[315]), .CLK(clk), .RST(rst), .Q(sreg[311]) );
  DFF \sreg_reg[310]  ( .D(c[314]), .CLK(clk), .RST(rst), .Q(sreg[310]) );
  DFF \sreg_reg[309]  ( .D(c[313]), .CLK(clk), .RST(rst), .Q(sreg[309]) );
  DFF \sreg_reg[308]  ( .D(c[312]), .CLK(clk), .RST(rst), .Q(sreg[308]) );
  DFF \sreg_reg[307]  ( .D(c[311]), .CLK(clk), .RST(rst), .Q(sreg[307]) );
  DFF \sreg_reg[306]  ( .D(c[310]), .CLK(clk), .RST(rst), .Q(sreg[306]) );
  DFF \sreg_reg[305]  ( .D(c[309]), .CLK(clk), .RST(rst), .Q(sreg[305]) );
  DFF \sreg_reg[304]  ( .D(c[308]), .CLK(clk), .RST(rst), .Q(sreg[304]) );
  DFF \sreg_reg[303]  ( .D(c[307]), .CLK(clk), .RST(rst), .Q(sreg[303]) );
  DFF \sreg_reg[302]  ( .D(c[306]), .CLK(clk), .RST(rst), .Q(sreg[302]) );
  DFF \sreg_reg[301]  ( .D(c[305]), .CLK(clk), .RST(rst), .Q(sreg[301]) );
  DFF \sreg_reg[300]  ( .D(c[304]), .CLK(clk), .RST(rst), .Q(sreg[300]) );
  DFF \sreg_reg[299]  ( .D(c[303]), .CLK(clk), .RST(rst), .Q(sreg[299]) );
  DFF \sreg_reg[298]  ( .D(c[302]), .CLK(clk), .RST(rst), .Q(sreg[298]) );
  DFF \sreg_reg[297]  ( .D(c[301]), .CLK(clk), .RST(rst), .Q(sreg[297]) );
  DFF \sreg_reg[296]  ( .D(c[300]), .CLK(clk), .RST(rst), .Q(sreg[296]) );
  DFF \sreg_reg[295]  ( .D(c[299]), .CLK(clk), .RST(rst), .Q(sreg[295]) );
  DFF \sreg_reg[294]  ( .D(c[298]), .CLK(clk), .RST(rst), .Q(sreg[294]) );
  DFF \sreg_reg[293]  ( .D(c[297]), .CLK(clk), .RST(rst), .Q(sreg[293]) );
  DFF \sreg_reg[292]  ( .D(c[296]), .CLK(clk), .RST(rst), .Q(sreg[292]) );
  DFF \sreg_reg[291]  ( .D(c[295]), .CLK(clk), .RST(rst), .Q(sreg[291]) );
  DFF \sreg_reg[290]  ( .D(c[294]), .CLK(clk), .RST(rst), .Q(sreg[290]) );
  DFF \sreg_reg[289]  ( .D(c[293]), .CLK(clk), .RST(rst), .Q(sreg[289]) );
  DFF \sreg_reg[288]  ( .D(c[292]), .CLK(clk), .RST(rst), .Q(sreg[288]) );
  DFF \sreg_reg[287]  ( .D(c[291]), .CLK(clk), .RST(rst), .Q(sreg[287]) );
  DFF \sreg_reg[286]  ( .D(c[290]), .CLK(clk), .RST(rst), .Q(sreg[286]) );
  DFF \sreg_reg[285]  ( .D(c[289]), .CLK(clk), .RST(rst), .Q(sreg[285]) );
  DFF \sreg_reg[284]  ( .D(c[288]), .CLK(clk), .RST(rst), .Q(sreg[284]) );
  DFF \sreg_reg[283]  ( .D(c[287]), .CLK(clk), .RST(rst), .Q(sreg[283]) );
  DFF \sreg_reg[282]  ( .D(c[286]), .CLK(clk), .RST(rst), .Q(sreg[282]) );
  DFF \sreg_reg[281]  ( .D(c[285]), .CLK(clk), .RST(rst), .Q(sreg[281]) );
  DFF \sreg_reg[280]  ( .D(c[284]), .CLK(clk), .RST(rst), .Q(sreg[280]) );
  DFF \sreg_reg[279]  ( .D(c[283]), .CLK(clk), .RST(rst), .Q(sreg[279]) );
  DFF \sreg_reg[278]  ( .D(c[282]), .CLK(clk), .RST(rst), .Q(sreg[278]) );
  DFF \sreg_reg[277]  ( .D(c[281]), .CLK(clk), .RST(rst), .Q(sreg[277]) );
  DFF \sreg_reg[276]  ( .D(c[280]), .CLK(clk), .RST(rst), .Q(sreg[276]) );
  DFF \sreg_reg[275]  ( .D(c[279]), .CLK(clk), .RST(rst), .Q(sreg[275]) );
  DFF \sreg_reg[274]  ( .D(c[278]), .CLK(clk), .RST(rst), .Q(sreg[274]) );
  DFF \sreg_reg[273]  ( .D(c[277]), .CLK(clk), .RST(rst), .Q(sreg[273]) );
  DFF \sreg_reg[272]  ( .D(c[276]), .CLK(clk), .RST(rst), .Q(sreg[272]) );
  DFF \sreg_reg[271]  ( .D(c[275]), .CLK(clk), .RST(rst), .Q(sreg[271]) );
  DFF \sreg_reg[270]  ( .D(c[274]), .CLK(clk), .RST(rst), .Q(sreg[270]) );
  DFF \sreg_reg[269]  ( .D(c[273]), .CLK(clk), .RST(rst), .Q(sreg[269]) );
  DFF \sreg_reg[268]  ( .D(c[272]), .CLK(clk), .RST(rst), .Q(sreg[268]) );
  DFF \sreg_reg[267]  ( .D(c[271]), .CLK(clk), .RST(rst), .Q(sreg[267]) );
  DFF \sreg_reg[266]  ( .D(c[270]), .CLK(clk), .RST(rst), .Q(sreg[266]) );
  DFF \sreg_reg[265]  ( .D(c[269]), .CLK(clk), .RST(rst), .Q(sreg[265]) );
  DFF \sreg_reg[264]  ( .D(c[268]), .CLK(clk), .RST(rst), .Q(sreg[264]) );
  DFF \sreg_reg[263]  ( .D(c[267]), .CLK(clk), .RST(rst), .Q(sreg[263]) );
  DFF \sreg_reg[262]  ( .D(c[266]), .CLK(clk), .RST(rst), .Q(sreg[262]) );
  DFF \sreg_reg[261]  ( .D(c[265]), .CLK(clk), .RST(rst), .Q(sreg[261]) );
  DFF \sreg_reg[260]  ( .D(c[264]), .CLK(clk), .RST(rst), .Q(sreg[260]) );
  DFF \sreg_reg[259]  ( .D(c[263]), .CLK(clk), .RST(rst), .Q(sreg[259]) );
  DFF \sreg_reg[258]  ( .D(c[262]), .CLK(clk), .RST(rst), .Q(sreg[258]) );
  DFF \sreg_reg[257]  ( .D(c[261]), .CLK(clk), .RST(rst), .Q(sreg[257]) );
  DFF \sreg_reg[256]  ( .D(c[260]), .CLK(clk), .RST(rst), .Q(sreg[256]) );
  DFF \sreg_reg[255]  ( .D(c[259]), .CLK(clk), .RST(rst), .Q(sreg[255]) );
  DFF \sreg_reg[254]  ( .D(c[258]), .CLK(clk), .RST(rst), .Q(sreg[254]) );
  DFF \sreg_reg[253]  ( .D(c[257]), .CLK(clk), .RST(rst), .Q(sreg[253]) );
  DFF \sreg_reg[252]  ( .D(c[256]), .CLK(clk), .RST(rst), .Q(sreg[252]) );
  DFF \sreg_reg[251]  ( .D(c[255]), .CLK(clk), .RST(rst), .Q(c[251]) );
  DFF \sreg_reg[250]  ( .D(c[254]), .CLK(clk), .RST(rst), .Q(c[250]) );
  DFF \sreg_reg[249]  ( .D(c[253]), .CLK(clk), .RST(rst), .Q(c[249]) );
  DFF \sreg_reg[248]  ( .D(c[252]), .CLK(clk), .RST(rst), .Q(c[248]) );
  DFF \sreg_reg[247]  ( .D(c[251]), .CLK(clk), .RST(rst), .Q(c[247]) );
  DFF \sreg_reg[246]  ( .D(c[250]), .CLK(clk), .RST(rst), .Q(c[246]) );
  DFF \sreg_reg[245]  ( .D(c[249]), .CLK(clk), .RST(rst), .Q(c[245]) );
  DFF \sreg_reg[244]  ( .D(c[248]), .CLK(clk), .RST(rst), .Q(c[244]) );
  DFF \sreg_reg[243]  ( .D(c[247]), .CLK(clk), .RST(rst), .Q(c[243]) );
  DFF \sreg_reg[242]  ( .D(c[246]), .CLK(clk), .RST(rst), .Q(c[242]) );
  DFF \sreg_reg[241]  ( .D(c[245]), .CLK(clk), .RST(rst), .Q(c[241]) );
  DFF \sreg_reg[240]  ( .D(c[244]), .CLK(clk), .RST(rst), .Q(c[240]) );
  DFF \sreg_reg[239]  ( .D(c[243]), .CLK(clk), .RST(rst), .Q(c[239]) );
  DFF \sreg_reg[238]  ( .D(c[242]), .CLK(clk), .RST(rst), .Q(c[238]) );
  DFF \sreg_reg[237]  ( .D(c[241]), .CLK(clk), .RST(rst), .Q(c[237]) );
  DFF \sreg_reg[236]  ( .D(c[240]), .CLK(clk), .RST(rst), .Q(c[236]) );
  DFF \sreg_reg[235]  ( .D(c[239]), .CLK(clk), .RST(rst), .Q(c[235]) );
  DFF \sreg_reg[234]  ( .D(c[238]), .CLK(clk), .RST(rst), .Q(c[234]) );
  DFF \sreg_reg[233]  ( .D(c[237]), .CLK(clk), .RST(rst), .Q(c[233]) );
  DFF \sreg_reg[232]  ( .D(c[236]), .CLK(clk), .RST(rst), .Q(c[232]) );
  DFF \sreg_reg[231]  ( .D(c[235]), .CLK(clk), .RST(rst), .Q(c[231]) );
  DFF \sreg_reg[230]  ( .D(c[234]), .CLK(clk), .RST(rst), .Q(c[230]) );
  DFF \sreg_reg[229]  ( .D(c[233]), .CLK(clk), .RST(rst), .Q(c[229]) );
  DFF \sreg_reg[228]  ( .D(c[232]), .CLK(clk), .RST(rst), .Q(c[228]) );
  DFF \sreg_reg[227]  ( .D(c[231]), .CLK(clk), .RST(rst), .Q(c[227]) );
  DFF \sreg_reg[226]  ( .D(c[230]), .CLK(clk), .RST(rst), .Q(c[226]) );
  DFF \sreg_reg[225]  ( .D(c[229]), .CLK(clk), .RST(rst), .Q(c[225]) );
  DFF \sreg_reg[224]  ( .D(c[228]), .CLK(clk), .RST(rst), .Q(c[224]) );
  DFF \sreg_reg[223]  ( .D(c[227]), .CLK(clk), .RST(rst), .Q(c[223]) );
  DFF \sreg_reg[222]  ( .D(c[226]), .CLK(clk), .RST(rst), .Q(c[222]) );
  DFF \sreg_reg[221]  ( .D(c[225]), .CLK(clk), .RST(rst), .Q(c[221]) );
  DFF \sreg_reg[220]  ( .D(c[224]), .CLK(clk), .RST(rst), .Q(c[220]) );
  DFF \sreg_reg[219]  ( .D(c[223]), .CLK(clk), .RST(rst), .Q(c[219]) );
  DFF \sreg_reg[218]  ( .D(c[222]), .CLK(clk), .RST(rst), .Q(c[218]) );
  DFF \sreg_reg[217]  ( .D(c[221]), .CLK(clk), .RST(rst), .Q(c[217]) );
  DFF \sreg_reg[216]  ( .D(c[220]), .CLK(clk), .RST(rst), .Q(c[216]) );
  DFF \sreg_reg[215]  ( .D(c[219]), .CLK(clk), .RST(rst), .Q(c[215]) );
  DFF \sreg_reg[214]  ( .D(c[218]), .CLK(clk), .RST(rst), .Q(c[214]) );
  DFF \sreg_reg[213]  ( .D(c[217]), .CLK(clk), .RST(rst), .Q(c[213]) );
  DFF \sreg_reg[212]  ( .D(c[216]), .CLK(clk), .RST(rst), .Q(c[212]) );
  DFF \sreg_reg[211]  ( .D(c[215]), .CLK(clk), .RST(rst), .Q(c[211]) );
  DFF \sreg_reg[210]  ( .D(c[214]), .CLK(clk), .RST(rst), .Q(c[210]) );
  DFF \sreg_reg[209]  ( .D(c[213]), .CLK(clk), .RST(rst), .Q(c[209]) );
  DFF \sreg_reg[208]  ( .D(c[212]), .CLK(clk), .RST(rst), .Q(c[208]) );
  DFF \sreg_reg[207]  ( .D(c[211]), .CLK(clk), .RST(rst), .Q(c[207]) );
  DFF \sreg_reg[206]  ( .D(c[210]), .CLK(clk), .RST(rst), .Q(c[206]) );
  DFF \sreg_reg[205]  ( .D(c[209]), .CLK(clk), .RST(rst), .Q(c[205]) );
  DFF \sreg_reg[204]  ( .D(c[208]), .CLK(clk), .RST(rst), .Q(c[204]) );
  DFF \sreg_reg[203]  ( .D(c[207]), .CLK(clk), .RST(rst), .Q(c[203]) );
  DFF \sreg_reg[202]  ( .D(c[206]), .CLK(clk), .RST(rst), .Q(c[202]) );
  DFF \sreg_reg[201]  ( .D(c[205]), .CLK(clk), .RST(rst), .Q(c[201]) );
  DFF \sreg_reg[200]  ( .D(c[204]), .CLK(clk), .RST(rst), .Q(c[200]) );
  DFF \sreg_reg[199]  ( .D(c[203]), .CLK(clk), .RST(rst), .Q(c[199]) );
  DFF \sreg_reg[198]  ( .D(c[202]), .CLK(clk), .RST(rst), .Q(c[198]) );
  DFF \sreg_reg[197]  ( .D(c[201]), .CLK(clk), .RST(rst), .Q(c[197]) );
  DFF \sreg_reg[196]  ( .D(c[200]), .CLK(clk), .RST(rst), .Q(c[196]) );
  DFF \sreg_reg[195]  ( .D(c[199]), .CLK(clk), .RST(rst), .Q(c[195]) );
  DFF \sreg_reg[194]  ( .D(c[198]), .CLK(clk), .RST(rst), .Q(c[194]) );
  DFF \sreg_reg[193]  ( .D(c[197]), .CLK(clk), .RST(rst), .Q(c[193]) );
  DFF \sreg_reg[192]  ( .D(c[196]), .CLK(clk), .RST(rst), .Q(c[192]) );
  DFF \sreg_reg[191]  ( .D(c[195]), .CLK(clk), .RST(rst), .Q(c[191]) );
  DFF \sreg_reg[190]  ( .D(c[194]), .CLK(clk), .RST(rst), .Q(c[190]) );
  DFF \sreg_reg[189]  ( .D(c[193]), .CLK(clk), .RST(rst), .Q(c[189]) );
  DFF \sreg_reg[188]  ( .D(c[192]), .CLK(clk), .RST(rst), .Q(c[188]) );
  DFF \sreg_reg[187]  ( .D(c[191]), .CLK(clk), .RST(rst), .Q(c[187]) );
  DFF \sreg_reg[186]  ( .D(c[190]), .CLK(clk), .RST(rst), .Q(c[186]) );
  DFF \sreg_reg[185]  ( .D(c[189]), .CLK(clk), .RST(rst), .Q(c[185]) );
  DFF \sreg_reg[184]  ( .D(c[188]), .CLK(clk), .RST(rst), .Q(c[184]) );
  DFF \sreg_reg[183]  ( .D(c[187]), .CLK(clk), .RST(rst), .Q(c[183]) );
  DFF \sreg_reg[182]  ( .D(c[186]), .CLK(clk), .RST(rst), .Q(c[182]) );
  DFF \sreg_reg[181]  ( .D(c[185]), .CLK(clk), .RST(rst), .Q(c[181]) );
  DFF \sreg_reg[180]  ( .D(c[184]), .CLK(clk), .RST(rst), .Q(c[180]) );
  DFF \sreg_reg[179]  ( .D(c[183]), .CLK(clk), .RST(rst), .Q(c[179]) );
  DFF \sreg_reg[178]  ( .D(c[182]), .CLK(clk), .RST(rst), .Q(c[178]) );
  DFF \sreg_reg[177]  ( .D(c[181]), .CLK(clk), .RST(rst), .Q(c[177]) );
  DFF \sreg_reg[176]  ( .D(c[180]), .CLK(clk), .RST(rst), .Q(c[176]) );
  DFF \sreg_reg[175]  ( .D(c[179]), .CLK(clk), .RST(rst), .Q(c[175]) );
  DFF \sreg_reg[174]  ( .D(c[178]), .CLK(clk), .RST(rst), .Q(c[174]) );
  DFF \sreg_reg[173]  ( .D(c[177]), .CLK(clk), .RST(rst), .Q(c[173]) );
  DFF \sreg_reg[172]  ( .D(c[176]), .CLK(clk), .RST(rst), .Q(c[172]) );
  DFF \sreg_reg[171]  ( .D(c[175]), .CLK(clk), .RST(rst), .Q(c[171]) );
  DFF \sreg_reg[170]  ( .D(c[174]), .CLK(clk), .RST(rst), .Q(c[170]) );
  DFF \sreg_reg[169]  ( .D(c[173]), .CLK(clk), .RST(rst), .Q(c[169]) );
  DFF \sreg_reg[168]  ( .D(c[172]), .CLK(clk), .RST(rst), .Q(c[168]) );
  DFF \sreg_reg[167]  ( .D(c[171]), .CLK(clk), .RST(rst), .Q(c[167]) );
  DFF \sreg_reg[166]  ( .D(c[170]), .CLK(clk), .RST(rst), .Q(c[166]) );
  DFF \sreg_reg[165]  ( .D(c[169]), .CLK(clk), .RST(rst), .Q(c[165]) );
  DFF \sreg_reg[164]  ( .D(c[168]), .CLK(clk), .RST(rst), .Q(c[164]) );
  DFF \sreg_reg[163]  ( .D(c[167]), .CLK(clk), .RST(rst), .Q(c[163]) );
  DFF \sreg_reg[162]  ( .D(c[166]), .CLK(clk), .RST(rst), .Q(c[162]) );
  DFF \sreg_reg[161]  ( .D(c[165]), .CLK(clk), .RST(rst), .Q(c[161]) );
  DFF \sreg_reg[160]  ( .D(c[164]), .CLK(clk), .RST(rst), .Q(c[160]) );
  DFF \sreg_reg[159]  ( .D(c[163]), .CLK(clk), .RST(rst), .Q(c[159]) );
  DFF \sreg_reg[158]  ( .D(c[162]), .CLK(clk), .RST(rst), .Q(c[158]) );
  DFF \sreg_reg[157]  ( .D(c[161]), .CLK(clk), .RST(rst), .Q(c[157]) );
  DFF \sreg_reg[156]  ( .D(c[160]), .CLK(clk), .RST(rst), .Q(c[156]) );
  DFF \sreg_reg[155]  ( .D(c[159]), .CLK(clk), .RST(rst), .Q(c[155]) );
  DFF \sreg_reg[154]  ( .D(c[158]), .CLK(clk), .RST(rst), .Q(c[154]) );
  DFF \sreg_reg[153]  ( .D(c[157]), .CLK(clk), .RST(rst), .Q(c[153]) );
  DFF \sreg_reg[152]  ( .D(c[156]), .CLK(clk), .RST(rst), .Q(c[152]) );
  DFF \sreg_reg[151]  ( .D(c[155]), .CLK(clk), .RST(rst), .Q(c[151]) );
  DFF \sreg_reg[150]  ( .D(c[154]), .CLK(clk), .RST(rst), .Q(c[150]) );
  DFF \sreg_reg[149]  ( .D(c[153]), .CLK(clk), .RST(rst), .Q(c[149]) );
  DFF \sreg_reg[148]  ( .D(c[152]), .CLK(clk), .RST(rst), .Q(c[148]) );
  DFF \sreg_reg[147]  ( .D(c[151]), .CLK(clk), .RST(rst), .Q(c[147]) );
  DFF \sreg_reg[146]  ( .D(c[150]), .CLK(clk), .RST(rst), .Q(c[146]) );
  DFF \sreg_reg[145]  ( .D(c[149]), .CLK(clk), .RST(rst), .Q(c[145]) );
  DFF \sreg_reg[144]  ( .D(c[148]), .CLK(clk), .RST(rst), .Q(c[144]) );
  DFF \sreg_reg[143]  ( .D(c[147]), .CLK(clk), .RST(rst), .Q(c[143]) );
  DFF \sreg_reg[142]  ( .D(c[146]), .CLK(clk), .RST(rst), .Q(c[142]) );
  DFF \sreg_reg[141]  ( .D(c[145]), .CLK(clk), .RST(rst), .Q(c[141]) );
  DFF \sreg_reg[140]  ( .D(c[144]), .CLK(clk), .RST(rst), .Q(c[140]) );
  DFF \sreg_reg[139]  ( .D(c[143]), .CLK(clk), .RST(rst), .Q(c[139]) );
  DFF \sreg_reg[138]  ( .D(c[142]), .CLK(clk), .RST(rst), .Q(c[138]) );
  DFF \sreg_reg[137]  ( .D(c[141]), .CLK(clk), .RST(rst), .Q(c[137]) );
  DFF \sreg_reg[136]  ( .D(c[140]), .CLK(clk), .RST(rst), .Q(c[136]) );
  DFF \sreg_reg[135]  ( .D(c[139]), .CLK(clk), .RST(rst), .Q(c[135]) );
  DFF \sreg_reg[134]  ( .D(c[138]), .CLK(clk), .RST(rst), .Q(c[134]) );
  DFF \sreg_reg[133]  ( .D(c[137]), .CLK(clk), .RST(rst), .Q(c[133]) );
  DFF \sreg_reg[132]  ( .D(c[136]), .CLK(clk), .RST(rst), .Q(c[132]) );
  DFF \sreg_reg[131]  ( .D(c[135]), .CLK(clk), .RST(rst), .Q(c[131]) );
  DFF \sreg_reg[130]  ( .D(c[134]), .CLK(clk), .RST(rst), .Q(c[130]) );
  DFF \sreg_reg[129]  ( .D(c[133]), .CLK(clk), .RST(rst), .Q(c[129]) );
  DFF \sreg_reg[128]  ( .D(c[132]), .CLK(clk), .RST(rst), .Q(c[128]) );
  DFF \sreg_reg[127]  ( .D(c[131]), .CLK(clk), .RST(rst), .Q(c[127]) );
  DFF \sreg_reg[126]  ( .D(c[130]), .CLK(clk), .RST(rst), .Q(c[126]) );
  DFF \sreg_reg[125]  ( .D(c[129]), .CLK(clk), .RST(rst), .Q(c[125]) );
  DFF \sreg_reg[124]  ( .D(c[128]), .CLK(clk), .RST(rst), .Q(c[124]) );
  DFF \sreg_reg[123]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(c[123]) );
  DFF \sreg_reg[122]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(c[122]) );
  DFF \sreg_reg[121]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(c[121]) );
  DFF \sreg_reg[120]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(c[120]) );
  DFF \sreg_reg[119]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(c[119]) );
  DFF \sreg_reg[118]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(c[118]) );
  DFF \sreg_reg[117]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(c[117]) );
  DFF \sreg_reg[116]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(c[116]) );
  DFF \sreg_reg[115]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(c[115]) );
  DFF \sreg_reg[114]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(c[114]) );
  DFF \sreg_reg[113]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(c[113]) );
  DFF \sreg_reg[112]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(c[112]) );
  DFF \sreg_reg[111]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(c[111]) );
  DFF \sreg_reg[110]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(c[110]) );
  DFF \sreg_reg[109]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(c[109]) );
  DFF \sreg_reg[108]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(c[108]) );
  DFF \sreg_reg[107]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(c[107]) );
  DFF \sreg_reg[106]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(c[106]) );
  DFF \sreg_reg[105]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(c[105]) );
  DFF \sreg_reg[104]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(c[104]) );
  DFF \sreg_reg[103]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(c[103]) );
  DFF \sreg_reg[102]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(c[102]) );
  DFF \sreg_reg[101]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(c[101]) );
  DFF \sreg_reg[100]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(c[100]) );
  DFF \sreg_reg[99]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(c[99]) );
  DFF \sreg_reg[98]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(c[98]) );
  DFF \sreg_reg[97]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(c[97]) );
  DFF \sreg_reg[96]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(c[96]) );
  DFF \sreg_reg[95]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(c[95]) );
  DFF \sreg_reg[94]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(c[94]) );
  DFF \sreg_reg[93]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(c[93]) );
  DFF \sreg_reg[92]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(c[92]) );
  DFF \sreg_reg[91]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(c[91]) );
  DFF \sreg_reg[90]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(c[90]) );
  DFF \sreg_reg[89]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(c[89]) );
  DFF \sreg_reg[88]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(c[88]) );
  DFF \sreg_reg[87]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(c[87]) );
  DFF \sreg_reg[86]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(c[86]) );
  DFF \sreg_reg[85]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(c[85]) );
  DFF \sreg_reg[84]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(c[84]) );
  DFF \sreg_reg[83]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(c[83]) );
  DFF \sreg_reg[82]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(c[82]) );
  DFF \sreg_reg[81]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(c[81]) );
  DFF \sreg_reg[80]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(c[80]) );
  DFF \sreg_reg[79]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(c[79]) );
  DFF \sreg_reg[78]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(c[78]) );
  DFF \sreg_reg[77]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(c[77]) );
  DFF \sreg_reg[76]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(c[76]) );
  DFF \sreg_reg[75]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(c[75]) );
  DFF \sreg_reg[74]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(c[74]) );
  DFF \sreg_reg[73]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(c[73]) );
  DFF \sreg_reg[72]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(c[72]) );
  DFF \sreg_reg[71]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(c[71]) );
  DFF \sreg_reg[70]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(c[70]) );
  DFF \sreg_reg[69]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(c[69]) );
  DFF \sreg_reg[68]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(c[68]) );
  DFF \sreg_reg[67]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(c[67]) );
  DFF \sreg_reg[66]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(c[66]) );
  DFF \sreg_reg[65]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(c[65]) );
  DFF \sreg_reg[64]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(c[64]) );
  DFF \sreg_reg[63]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(c[63]) );
  DFF \sreg_reg[62]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(c[62]) );
  DFF \sreg_reg[61]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[60]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[59]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[58]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[57]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[56]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[55]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[54]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[53]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[52]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[51]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[50]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[49]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[48]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[47]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[46]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[45]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[44]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[43]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[42]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[41]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[40]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[39]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[38]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[37]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[36]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[35]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[34]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[33]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[32]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[31]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[30]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[29]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[28]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[27]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[26]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[25]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[24]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[23]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[22]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[21]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[20]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[19]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[18]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[17]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[16]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[15]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[14]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[13]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[12]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[11]  ( .D(c[15]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[10]  ( .D(c[14]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[9]  ( .D(c[13]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[8]  ( .D(c[12]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[7]  ( .D(c[11]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[6]  ( .D(c[10]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[5]  ( .D(c[9]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[4]  ( .D(c[8]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[3]  ( .D(c[7]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[2]  ( .D(c[6]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[1]  ( .D(c[5]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[0]  ( .D(c[4]), .CLK(clk), .RST(rst), .Q(c[0]) );
  OR U7 ( .A(n5903), .B(n5904), .Z(n1) );
  NANDN U8 ( .A(n5906), .B(n5905), .Z(n2) );
  AND U9 ( .A(n1), .B(n2), .Z(n5913) );
  OR U10 ( .A(n5960), .B(n5917), .Z(n3) );
  NANDN U11 ( .A(n5919), .B(n5918), .Z(n4) );
  AND U12 ( .A(n3), .B(n4), .Z(n5948) );
  NANDN U13 ( .A(n2208), .B(n2207), .Z(n5) );
  NANDN U14 ( .A(n2209), .B(n2210), .Z(n6) );
  NAND U15 ( .A(n5), .B(n6), .Z(n2217) );
  NANDN U16 ( .A(n4327), .B(n4326), .Z(n7) );
  NANDN U17 ( .A(n4328), .B(n4329), .Z(n8) );
  NAND U18 ( .A(n7), .B(n8), .Z(n4334) );
  NANDN U19 ( .A(n5729), .B(n5728), .Z(n9) );
  NANDN U20 ( .A(n5730), .B(n5731), .Z(n10) );
  NAND U21 ( .A(n9), .B(n10), .Z(n5753) );
  NANDN U22 ( .A(n5914), .B(n5915), .Z(n11) );
  NANDN U23 ( .A(n5912), .B(n5913), .Z(n12) );
  NAND U24 ( .A(n11), .B(n12), .Z(n5937) );
  XOR U25 ( .A(sreg[260]), .B(n528), .Z(n13) );
  NANDN U26 ( .A(n529), .B(n13), .Z(n14) );
  NAND U27 ( .A(sreg[260]), .B(n528), .Z(n15) );
  AND U28 ( .A(n14), .B(n15), .Z(n568) );
  NAND U29 ( .A(n723), .B(n722), .Z(n16) );
  XOR U30 ( .A(n722), .B(n723), .Z(n17) );
  NANDN U31 ( .A(sreg[268]), .B(n17), .Z(n18) );
  NAND U32 ( .A(n16), .B(n18), .Z(n743) );
  NAND U33 ( .A(n897), .B(sreg[276]), .Z(n19) );
  XOR U34 ( .A(sreg[276]), .B(n897), .Z(n20) );
  NANDN U35 ( .A(n896), .B(n20), .Z(n21) );
  NAND U36 ( .A(n19), .B(n21), .Z(n899) );
  NAND U37 ( .A(n1094), .B(sreg[285]), .Z(n22) );
  XOR U38 ( .A(sreg[285]), .B(n1094), .Z(n23) );
  NAND U39 ( .A(n23), .B(n1093), .Z(n24) );
  NAND U40 ( .A(n22), .B(n24), .Z(n1096) );
  XOR U41 ( .A(n1331), .B(n1330), .Z(n25) );
  NANDN U42 ( .A(sreg[296]), .B(n25), .Z(n26) );
  NAND U43 ( .A(n1331), .B(n1330), .Z(n27) );
  AND U44 ( .A(n26), .B(n27), .Z(n1333) );
  NAND U45 ( .A(n1884), .B(sreg[321]), .Z(n28) );
  XOR U46 ( .A(sreg[321]), .B(n1884), .Z(n29) );
  NAND U47 ( .A(n29), .B(n1883), .Z(n30) );
  NAND U48 ( .A(n28), .B(n30), .Z(n1886) );
  NAND U49 ( .A(sreg[346]), .B(n2434), .Z(n31) );
  XOR U50 ( .A(n2434), .B(sreg[346]), .Z(n32) );
  NANDN U51 ( .A(n2435), .B(n32), .Z(n33) );
  NAND U52 ( .A(n31), .B(n33), .Z(n2437) );
  NAND U53 ( .A(n2542), .B(sreg[351]), .Z(n34) );
  XOR U54 ( .A(sreg[351]), .B(n2542), .Z(n35) );
  NAND U55 ( .A(n35), .B(n2541), .Z(n36) );
  NAND U56 ( .A(n34), .B(n36), .Z(n2563) );
  NAND U57 ( .A(sreg[365]), .B(n2849), .Z(n37) );
  XOR U58 ( .A(n2849), .B(sreg[365]), .Z(n38) );
  NANDN U59 ( .A(n2850), .B(n38), .Z(n39) );
  NAND U60 ( .A(n37), .B(n39), .Z(n2852) );
  XOR U61 ( .A(n3293), .B(sreg[385]), .Z(n40) );
  NANDN U62 ( .A(n3294), .B(n40), .Z(n41) );
  NAND U63 ( .A(n3293), .B(sreg[385]), .Z(n42) );
  AND U64 ( .A(n41), .B(n42), .Z(n3314) );
  NAND U65 ( .A(sreg[390]), .B(n3402), .Z(n43) );
  XOR U66 ( .A(n3402), .B(sreg[390]), .Z(n44) );
  NANDN U67 ( .A(n3403), .B(n44), .Z(n45) );
  NAND U68 ( .A(n43), .B(n45), .Z(n3405) );
  XOR U69 ( .A(n4180), .B(n4179), .Z(n46) );
  NAND U70 ( .A(n46), .B(sreg[425]), .Z(n47) );
  NAND U71 ( .A(n4180), .B(n4179), .Z(n48) );
  AND U72 ( .A(n47), .B(n48), .Z(n4182) );
  NAND U73 ( .A(sreg[441]), .B(n4531), .Z(n49) );
  XOR U74 ( .A(n4531), .B(sreg[441]), .Z(n50) );
  NANDN U75 ( .A(n4532), .B(n50), .Z(n51) );
  NAND U76 ( .A(n49), .B(n51), .Z(n4552) );
  XOR U77 ( .A(n4711), .B(sreg[450]), .Z(n52) );
  NANDN U78 ( .A(n4710), .B(n52), .Z(n53) );
  NAND U79 ( .A(n4711), .B(sreg[450]), .Z(n54) );
  AND U80 ( .A(n53), .B(n54), .Z(n4732) );
  XOR U81 ( .A(sreg[455]), .B(n4837), .Z(n55) );
  NANDN U82 ( .A(n4838), .B(n55), .Z(n56) );
  NAND U83 ( .A(sreg[455]), .B(n4837), .Z(n57) );
  AND U84 ( .A(n56), .B(n57), .Z(n4840) );
  XOR U85 ( .A(n5123), .B(sreg[468]), .Z(n58) );
  NANDN U86 ( .A(n5122), .B(n58), .Z(n59) );
  NAND U87 ( .A(n5123), .B(sreg[468]), .Z(n60) );
  AND U88 ( .A(n59), .B(n60), .Z(n5143) );
  NAND U89 ( .A(n5209), .B(sreg[472]), .Z(n61) );
  XOR U90 ( .A(sreg[472]), .B(n5209), .Z(n62) );
  NANDN U91 ( .A(n5208), .B(n62), .Z(n63) );
  NAND U92 ( .A(n61), .B(n63), .Z(n5230) );
  XOR U93 ( .A(n5364), .B(sreg[479]), .Z(n64) );
  NANDN U94 ( .A(n5363), .B(n64), .Z(n65) );
  NAND U95 ( .A(n5364), .B(sreg[479]), .Z(n66) );
  AND U96 ( .A(n65), .B(n66), .Z(n5366) );
  NAND U97 ( .A(sreg[500]), .B(n5824), .Z(n67) );
  XOR U98 ( .A(n5824), .B(sreg[500]), .Z(n68) );
  NANDN U99 ( .A(n5825), .B(n68), .Z(n69) );
  NAND U100 ( .A(n67), .B(n69), .Z(n5827) );
  AND U101 ( .A(b[0]), .B(a[1]), .Z(n445) );
  NANDN U102 ( .A(n1147), .B(n1146), .Z(n70) );
  NANDN U103 ( .A(n1148), .B(n1149), .Z(n71) );
  NAND U104 ( .A(n70), .B(n71), .Z(n1173) );
  NANDN U105 ( .A(n2578), .B(n2577), .Z(n72) );
  NANDN U106 ( .A(n2579), .B(n2580), .Z(n73) );
  NAND U107 ( .A(n72), .B(n73), .Z(n2582) );
  NAND U108 ( .A(n2199), .B(n2198), .Z(n74) );
  XOR U109 ( .A(n2198), .B(n2199), .Z(n75) );
  NANDN U110 ( .A(n2200), .B(n75), .Z(n76) );
  NAND U111 ( .A(n74), .B(n76), .Z(n2218) );
  NANDN U112 ( .A(n414), .B(n415), .Z(n77) );
  NANDN U113 ( .A(n413), .B(n412), .Z(n78) );
  AND U114 ( .A(n77), .B(n78), .Z(n420) );
  NAND U115 ( .A(n1080), .B(n1078), .Z(n79) );
  XOR U116 ( .A(n1078), .B(n1080), .Z(n80) );
  NANDN U117 ( .A(n1079), .B(n80), .Z(n81) );
  NAND U118 ( .A(n79), .B(n81), .Z(n1101) );
  NAND U119 ( .A(n2504), .B(n2502), .Z(n82) );
  XOR U120 ( .A(n2502), .B(n2504), .Z(n83) );
  NANDN U121 ( .A(n2503), .B(n83), .Z(n84) );
  NAND U122 ( .A(n82), .B(n84), .Z(n2526) );
  NAND U123 ( .A(n4319), .B(n4318), .Z(n85) );
  XOR U124 ( .A(n4318), .B(n4319), .Z(n86) );
  NAND U125 ( .A(n86), .B(n4317), .Z(n87) );
  NAND U126 ( .A(n85), .B(n87), .Z(n4335) );
  NAND U127 ( .A(n5726), .B(n5725), .Z(n88) );
  XOR U128 ( .A(n5725), .B(n5726), .Z(n89) );
  NANDN U129 ( .A(n5727), .B(n89), .Z(n90) );
  NAND U130 ( .A(n88), .B(n90), .Z(n5756) );
  NANDN U131 ( .A(n5936), .B(n5937), .Z(n91) );
  NANDN U132 ( .A(n5934), .B(n5935), .Z(n92) );
  NAND U133 ( .A(n91), .B(n92), .Z(n5956) );
  NAND U134 ( .A(sreg[257]), .B(n481), .Z(n93) );
  XOR U135 ( .A(n481), .B(sreg[257]), .Z(n94) );
  NANDN U136 ( .A(n482), .B(n94), .Z(n95) );
  NAND U137 ( .A(n93), .B(n95), .Z(n484) );
  NAND U138 ( .A(sreg[262]), .B(n590), .Z(n96) );
  XOR U139 ( .A(n590), .B(sreg[262]), .Z(n97) );
  NANDN U140 ( .A(n591), .B(n97), .Z(n98) );
  NAND U141 ( .A(n96), .B(n98), .Z(n593) );
  XOR U142 ( .A(sreg[266]), .B(n660), .Z(n99) );
  NANDN U143 ( .A(n661), .B(n99), .Z(n100) );
  NAND U144 ( .A(sreg[266]), .B(n660), .Z(n101) );
  AND U145 ( .A(n100), .B(n101), .Z(n700) );
  XOR U146 ( .A(sreg[270]), .B(n746), .Z(n102) );
  NANDN U147 ( .A(n747), .B(n102), .Z(n103) );
  NAND U148 ( .A(sreg[270]), .B(n746), .Z(n104) );
  AND U149 ( .A(n103), .B(n104), .Z(n786) );
  NAND U150 ( .A(n835), .B(n834), .Z(n105) );
  XOR U151 ( .A(n834), .B(n835), .Z(n106) );
  NAND U152 ( .A(n106), .B(sreg[274]), .Z(n107) );
  NAND U153 ( .A(n105), .B(n107), .Z(n873) );
  NAND U154 ( .A(n944), .B(sreg[279]), .Z(n108) );
  XOR U155 ( .A(sreg[279]), .B(n944), .Z(n109) );
  NANDN U156 ( .A(n943), .B(n109), .Z(n110) );
  NAND U157 ( .A(n108), .B(n110), .Z(n983) );
  XOR U158 ( .A(sreg[288]), .B(n1141), .Z(n111) );
  NANDN U159 ( .A(n1142), .B(n111), .Z(n112) );
  NAND U160 ( .A(sreg[288]), .B(n1141), .Z(n113) );
  AND U161 ( .A(n112), .B(n113), .Z(n1158) );
  NAND U162 ( .A(n1248), .B(sreg[293]), .Z(n114) );
  XOR U163 ( .A(sreg[293]), .B(n1248), .Z(n115) );
  NANDN U164 ( .A(n1247), .B(n115), .Z(n116) );
  NAND U165 ( .A(n114), .B(n116), .Z(n1286) );
  XOR U166 ( .A(sreg[297]), .B(n1333), .Z(n117) );
  NANDN U167 ( .A(n1334), .B(n117), .Z(n118) );
  NAND U168 ( .A(sreg[297]), .B(n1333), .Z(n119) );
  AND U169 ( .A(n118), .B(n119), .Z(n1373) );
  XOR U170 ( .A(sreg[302]), .B(n1444), .Z(n120) );
  NANDN U171 ( .A(n1445), .B(n120), .Z(n121) );
  NAND U172 ( .A(sreg[302]), .B(n1444), .Z(n122) );
  AND U173 ( .A(n121), .B(n122), .Z(n1484) );
  XOR U174 ( .A(sreg[306]), .B(n1532), .Z(n123) );
  NANDN U175 ( .A(n1533), .B(n123), .Z(n124) );
  NAND U176 ( .A(sreg[306]), .B(n1532), .Z(n125) );
  AND U177 ( .A(n124), .B(n125), .Z(n1572) );
  NAND U178 ( .A(n1644), .B(sreg[311]), .Z(n126) );
  XOR U179 ( .A(sreg[311]), .B(n1644), .Z(n127) );
  NANDN U180 ( .A(n1643), .B(n127), .Z(n128) );
  NAND U181 ( .A(n126), .B(n128), .Z(n1683) );
  XOR U182 ( .A(sreg[316]), .B(n1754), .Z(n129) );
  NANDN U183 ( .A(n1755), .B(n129), .Z(n130) );
  NAND U184 ( .A(sreg[316]), .B(n1754), .Z(n131) );
  AND U185 ( .A(n130), .B(n131), .Z(n1794) );
  XOR U186 ( .A(n1931), .B(n1930), .Z(n132) );
  NANDN U187 ( .A(sreg[324]), .B(n132), .Z(n133) );
  NAND U188 ( .A(n1931), .B(n1930), .Z(n134) );
  AND U189 ( .A(n133), .B(n134), .Z(n1969) );
  NAND U190 ( .A(n2018), .B(sreg[328]), .Z(n135) );
  XOR U191 ( .A(sreg[328]), .B(n2018), .Z(n136) );
  NANDN U192 ( .A(n2019), .B(n136), .Z(n137) );
  NAND U193 ( .A(n135), .B(n137), .Z(n2057) );
  XOR U194 ( .A(sreg[335]), .B(n2177), .Z(n138) );
  NANDN U195 ( .A(n2178), .B(n138), .Z(n139) );
  NAND U196 ( .A(sreg[335]), .B(n2177), .Z(n140) );
  AND U197 ( .A(n139), .B(n140), .Z(n2213) );
  NAND U198 ( .A(n2285), .B(sreg[340]), .Z(n141) );
  XOR U199 ( .A(sreg[340]), .B(n2285), .Z(n142) );
  NANDN U200 ( .A(n2284), .B(n142), .Z(n143) );
  NAND U201 ( .A(n141), .B(n143), .Z(n2323) );
  NAND U202 ( .A(sreg[345]), .B(n2413), .Z(n144) );
  XOR U203 ( .A(n2413), .B(sreg[345]), .Z(n145) );
  NANDN U204 ( .A(n2414), .B(n145), .Z(n146) );
  NAND U205 ( .A(n144), .B(n146), .Z(n2434) );
  NAND U206 ( .A(n2482), .B(n2481), .Z(n147) );
  XOR U207 ( .A(n2481), .B(n2482), .Z(n148) );
  NAND U208 ( .A(n148), .B(sreg[349]), .Z(n149) );
  NAND U209 ( .A(n147), .B(n149), .Z(n2519) );
  NAND U210 ( .A(n2566), .B(sreg[353]), .Z(n150) );
  XOR U211 ( .A(sreg[353]), .B(n2566), .Z(n151) );
  NANDN U212 ( .A(n2567), .B(n151), .Z(n152) );
  NAND U213 ( .A(n150), .B(n152), .Z(n2600) );
  NAND U214 ( .A(sreg[364]), .B(n2828), .Z(n153) );
  XOR U215 ( .A(n2828), .B(sreg[364]), .Z(n154) );
  NANDN U216 ( .A(n2829), .B(n154), .Z(n155) );
  NAND U217 ( .A(n153), .B(n155), .Z(n2849) );
  XOR U218 ( .A(sreg[368]), .B(n2896), .Z(n156) );
  NANDN U219 ( .A(n2897), .B(n156), .Z(n157) );
  NAND U220 ( .A(sreg[368]), .B(n2896), .Z(n158) );
  AND U221 ( .A(n157), .B(n158), .Z(n2918) );
  XOR U222 ( .A(n3008), .B(sreg[373]), .Z(n159) );
  NAND U223 ( .A(n159), .B(n3007), .Z(n160) );
  NAND U224 ( .A(n3008), .B(sreg[373]), .Z(n161) );
  AND U225 ( .A(n160), .B(n161), .Z(n3046) );
  NAND U226 ( .A(n3315), .B(sreg[386]), .Z(n162) );
  XOR U227 ( .A(sreg[386]), .B(n3315), .Z(n163) );
  NANDN U228 ( .A(n3314), .B(n163), .Z(n164) );
  NAND U229 ( .A(n162), .B(n164), .Z(n3317) );
  NAND U230 ( .A(n3406), .B(n3405), .Z(n165) );
  XOR U231 ( .A(n3405), .B(n3406), .Z(n166) );
  NAND U232 ( .A(n166), .B(sreg[391]), .Z(n167) );
  NAND U233 ( .A(n165), .B(n167), .Z(n3427) );
  XOR U234 ( .A(sreg[396]), .B(n3516), .Z(n168) );
  NANDN U235 ( .A(n3517), .B(n168), .Z(n169) );
  NAND U236 ( .A(sreg[396]), .B(n3516), .Z(n170) );
  AND U237 ( .A(n169), .B(n170), .Z(n3538) );
  XOR U238 ( .A(n3651), .B(sreg[402]), .Z(n171) );
  NAND U239 ( .A(n171), .B(n3650), .Z(n172) );
  NAND U240 ( .A(n3651), .B(sreg[402]), .Z(n173) );
  AND U241 ( .A(n172), .B(n173), .Z(n3690) );
  NAND U242 ( .A(sreg[412]), .B(n3892), .Z(n174) );
  XOR U243 ( .A(n3892), .B(sreg[412]), .Z(n175) );
  NANDN U244 ( .A(n3893), .B(n175), .Z(n176) );
  NAND U245 ( .A(n174), .B(n176), .Z(n3895) );
  NAND U246 ( .A(n3963), .B(n3962), .Z(n177) );
  XOR U247 ( .A(n3962), .B(n3963), .Z(n178) );
  NAND U248 ( .A(n178), .B(sreg[416]), .Z(n179) );
  NAND U249 ( .A(n177), .B(n179), .Z(n4001) );
  XOR U250 ( .A(sreg[422]), .B(n4096), .Z(n180) );
  NANDN U251 ( .A(n4097), .B(n180), .Z(n181) );
  NAND U252 ( .A(sreg[422]), .B(n4096), .Z(n182) );
  AND U253 ( .A(n181), .B(n182), .Z(n4136) );
  NAND U254 ( .A(n4183), .B(n4182), .Z(n183) );
  XOR U255 ( .A(n4182), .B(n4183), .Z(n184) );
  NANDN U256 ( .A(sreg[426]), .B(n184), .Z(n185) );
  NAND U257 ( .A(n183), .B(n185), .Z(n4222) );
  XOR U258 ( .A(n4269), .B(sreg[430]), .Z(n186) );
  NAND U259 ( .A(n186), .B(n4268), .Z(n187) );
  NAND U260 ( .A(n4269), .B(sreg[430]), .Z(n188) );
  AND U261 ( .A(n187), .B(n188), .Z(n4309) );
  NAND U262 ( .A(n4553), .B(sreg[442]), .Z(n189) );
  XOR U263 ( .A(sreg[442]), .B(n4553), .Z(n190) );
  NAND U264 ( .A(n190), .B(n4552), .Z(n191) );
  NAND U265 ( .A(n189), .B(n191), .Z(n4555) );
  XOR U266 ( .A(sreg[447]), .B(n4645), .Z(n192) );
  NANDN U267 ( .A(n4646), .B(n192), .Z(n193) );
  NAND U268 ( .A(sreg[447]), .B(n4645), .Z(n194) );
  AND U269 ( .A(n193), .B(n194), .Z(n4684) );
  NAND U270 ( .A(sreg[452]), .B(n4772), .Z(n195) );
  XOR U271 ( .A(n4772), .B(sreg[452]), .Z(n196) );
  NANDN U272 ( .A(n4773), .B(n196), .Z(n197) );
  NAND U273 ( .A(n195), .B(n197), .Z(n4775) );
  XOR U274 ( .A(n4841), .B(sreg[456]), .Z(n198) );
  NANDN U275 ( .A(n4840), .B(n198), .Z(n199) );
  NAND U276 ( .A(n4841), .B(sreg[456]), .Z(n200) );
  AND U277 ( .A(n199), .B(n200), .Z(n4880) );
  XOR U278 ( .A(sreg[460]), .B(n4928), .Z(n201) );
  NANDN U279 ( .A(n4929), .B(n201), .Z(n202) );
  NAND U280 ( .A(sreg[460]), .B(n4928), .Z(n203) );
  AND U281 ( .A(n202), .B(n203), .Z(n4968) );
  XOR U282 ( .A(n5058), .B(sreg[465]), .Z(n204) );
  NANDN U283 ( .A(n5057), .B(n204), .Z(n205) );
  NAND U284 ( .A(n5058), .B(sreg[465]), .Z(n206) );
  AND U285 ( .A(n205), .B(n206), .Z(n5060) );
  XOR U286 ( .A(n5144), .B(n5143), .Z(n207) );
  NANDN U287 ( .A(sreg[469]), .B(n207), .Z(n208) );
  NAND U288 ( .A(n5144), .B(n5143), .Z(n209) );
  AND U289 ( .A(n208), .B(n209), .Z(n5146) );
  NAND U290 ( .A(n5230), .B(sreg[473]), .Z(n210) );
  XOR U291 ( .A(sreg[473]), .B(n5230), .Z(n211) );
  NAND U292 ( .A(n211), .B(n5229), .Z(n212) );
  NAND U293 ( .A(n210), .B(n212), .Z(n5232) );
  NAND U294 ( .A(n5411), .B(sreg[482]), .Z(n213) );
  XOR U295 ( .A(sreg[482]), .B(n5411), .Z(n214) );
  NANDN U296 ( .A(n5410), .B(n214), .Z(n215) );
  NAND U297 ( .A(n213), .B(n215), .Z(n5449) );
  NAND U298 ( .A(n5545), .B(n5544), .Z(n216) );
  XOR U299 ( .A(n5544), .B(n5545), .Z(n217) );
  NAND U300 ( .A(n217), .B(sreg[488]), .Z(n218) );
  NAND U301 ( .A(n216), .B(n218), .Z(n5583) );
  XOR U302 ( .A(sreg[495]), .B(n5699), .Z(n219) );
  NANDN U303 ( .A(n5700), .B(n219), .Z(n220) );
  NAND U304 ( .A(sreg[495]), .B(n5699), .Z(n221) );
  AND U305 ( .A(n220), .B(n221), .Z(n5722) );
  NAND U306 ( .A(n5827), .B(sreg[501]), .Z(n222) );
  XOR U307 ( .A(sreg[501]), .B(n5827), .Z(n223) );
  NANDN U308 ( .A(n5828), .B(n223), .Z(n224) );
  NAND U309 ( .A(n222), .B(n224), .Z(n5866) );
  NAND U310 ( .A(b[2]), .B(a[2]), .Z(n448) );
  XOR U311 ( .A(n469), .B(n470), .Z(n471) );
  NAND U312 ( .A(n1144), .B(n1143), .Z(n225) );
  XOR U313 ( .A(n1143), .B(n1144), .Z(n226) );
  NANDN U314 ( .A(n1145), .B(n226), .Z(n227) );
  NAND U315 ( .A(n225), .B(n227), .Z(n1176) );
  NAND U316 ( .A(n2570), .B(n2569), .Z(n228) );
  XOR U317 ( .A(n2569), .B(n2570), .Z(n229) );
  NAND U318 ( .A(n229), .B(n2568), .Z(n230) );
  NAND U319 ( .A(n228), .B(n230), .Z(n2583) );
  NAND U320 ( .A(n5662), .B(n5660), .Z(n231) );
  XOR U321 ( .A(n5660), .B(n5662), .Z(n232) );
  NANDN U322 ( .A(n5661), .B(n232), .Z(n233) );
  NAND U323 ( .A(n231), .B(n233), .Z(n5678) );
  OR U324 ( .A(n5945), .B(n5946), .Z(n234) );
  NAND U325 ( .A(n5947), .B(n5948), .Z(n235) );
  AND U326 ( .A(n234), .B(n235), .Z(n5954) );
  NANDN U327 ( .A(n5967), .B(n5968), .Z(n236) );
  NANDN U328 ( .A(n5966), .B(n5965), .Z(n237) );
  AND U329 ( .A(n236), .B(n237), .Z(n5971) );
  XOR U330 ( .A(sreg[254]), .B(n416), .Z(n238) );
  NANDN U331 ( .A(n417), .B(n238), .Z(n239) );
  NAND U332 ( .A(sreg[254]), .B(n416), .Z(n240) );
  AND U333 ( .A(n239), .B(n240), .Z(n434) );
  XOR U334 ( .A(n4249), .B(n4248), .Z(n241) );
  NANDN U335 ( .A(n4247), .B(n241), .Z(n242) );
  NAND U336 ( .A(n4249), .B(n4248), .Z(n243) );
  AND U337 ( .A(n242), .B(n243), .Z(n4273) );
  XOR U338 ( .A(n5933), .B(sreg[506]), .Z(n244) );
  NAND U339 ( .A(n244), .B(n5932), .Z(n245) );
  NAND U340 ( .A(n5933), .B(sreg[506]), .Z(n246) );
  AND U341 ( .A(n245), .B(n246), .Z(n5949) );
  NANDN U342 ( .A(n5978), .B(n5977), .Z(n247) );
  NANDN U343 ( .A(n5979), .B(n5980), .Z(n248) );
  NAND U344 ( .A(n247), .B(n248), .Z(n5983) );
  NAND U345 ( .A(n485), .B(n484), .Z(n249) );
  XOR U346 ( .A(n484), .B(n485), .Z(n250) );
  NAND U347 ( .A(n250), .B(sreg[258]), .Z(n251) );
  NAND U348 ( .A(n249), .B(n251), .Z(n523) );
  NAND U349 ( .A(n594), .B(n593), .Z(n252) );
  XOR U350 ( .A(n593), .B(n594), .Z(n253) );
  NAND U351 ( .A(n253), .B(sreg[263]), .Z(n254) );
  NAND U352 ( .A(n252), .B(n254), .Z(n632) );
  NAND U353 ( .A(n744), .B(sreg[269]), .Z(n255) );
  XOR U354 ( .A(sreg[269]), .B(n744), .Z(n256) );
  NANDN U355 ( .A(n743), .B(n256), .Z(n257) );
  NAND U356 ( .A(n255), .B(n257), .Z(n746) );
  NAND U357 ( .A(sreg[273]), .B(n831), .Z(n258) );
  XOR U358 ( .A(n831), .B(sreg[273]), .Z(n259) );
  NANDN U359 ( .A(n832), .B(n259), .Z(n260) );
  NAND U360 ( .A(n258), .B(n260), .Z(n834) );
  NAND U361 ( .A(n900), .B(n899), .Z(n261) );
  XOR U362 ( .A(n899), .B(n900), .Z(n262) );
  NAND U363 ( .A(n262), .B(sreg[277]), .Z(n263) );
  NAND U364 ( .A(n261), .B(n263), .Z(n938) );
  NAND U365 ( .A(n1011), .B(sreg[282]), .Z(n264) );
  XOR U366 ( .A(sreg[282]), .B(n1011), .Z(n265) );
  NANDN U367 ( .A(n1010), .B(n265), .Z(n266) );
  NAND U368 ( .A(n264), .B(n266), .Z(n1049) );
  NAND U369 ( .A(n1096), .B(sreg[286]), .Z(n267) );
  XOR U370 ( .A(sreg[286]), .B(n1096), .Z(n268) );
  NANDN U371 ( .A(n1097), .B(n268), .Z(n269) );
  NAND U372 ( .A(n267), .B(n269), .Z(n1137) );
  XOR U373 ( .A(sreg[291]), .B(n1203), .Z(n270) );
  NANDN U374 ( .A(n1204), .B(n270), .Z(n271) );
  NAND U375 ( .A(sreg[291]), .B(n1203), .Z(n272) );
  AND U376 ( .A(n271), .B(n272), .Z(n1243) );
  XOR U377 ( .A(n1310), .B(sreg[295]), .Z(n273) );
  NANDN U378 ( .A(n1309), .B(n273), .Z(n274) );
  NAND U379 ( .A(n1310), .B(sreg[295]), .Z(n275) );
  AND U380 ( .A(n274), .B(n275), .Z(n1330) );
  XOR U381 ( .A(sreg[299]), .B(n1377), .Z(n276) );
  NANDN U382 ( .A(n1378), .B(n276), .Z(n277) );
  NAND U383 ( .A(sreg[299]), .B(n1377), .Z(n278) );
  AND U384 ( .A(n277), .B(n278), .Z(n1417) );
  XOR U385 ( .A(sreg[304]), .B(n1488), .Z(n279) );
  NANDN U386 ( .A(n1489), .B(n279), .Z(n280) );
  NAND U387 ( .A(sreg[304]), .B(n1488), .Z(n281) );
  AND U388 ( .A(n280), .B(n281), .Z(n1528) );
  XOR U389 ( .A(sreg[309]), .B(n1599), .Z(n282) );
  NANDN U390 ( .A(n1600), .B(n282), .Z(n283) );
  NAND U391 ( .A(sreg[309]), .B(n1599), .Z(n284) );
  AND U392 ( .A(n283), .B(n284), .Z(n1639) );
  XOR U393 ( .A(sreg[313]), .B(n1687), .Z(n285) );
  NANDN U394 ( .A(n1688), .B(n285), .Z(n286) );
  NAND U395 ( .A(sreg[313]), .B(n1687), .Z(n287) );
  AND U396 ( .A(n286), .B(n287), .Z(n1727) );
  XOR U397 ( .A(n1799), .B(sreg[318]), .Z(n288) );
  NAND U398 ( .A(n288), .B(n1798), .Z(n289) );
  NAND U399 ( .A(n1799), .B(sreg[318]), .Z(n290) );
  AND U400 ( .A(n289), .B(n290), .Z(n1838) );
  XOR U401 ( .A(n1887), .B(sreg[322]), .Z(n291) );
  NAND U402 ( .A(n291), .B(n1886), .Z(n292) );
  NAND U403 ( .A(n1887), .B(sreg[322]), .Z(n293) );
  AND U404 ( .A(n292), .B(n293), .Z(n1926) );
  NAND U405 ( .A(sreg[327]), .B(n2015), .Z(n294) );
  XOR U406 ( .A(n2015), .B(sreg[327]), .Z(n295) );
  NANDN U407 ( .A(n2016), .B(n295), .Z(n296) );
  NAND U408 ( .A(n294), .B(n296), .Z(n2018) );
  XOR U409 ( .A(n2086), .B(n2085), .Z(n297) );
  NANDN U410 ( .A(sreg[331]), .B(n297), .Z(n298) );
  NAND U411 ( .A(n2086), .B(n2085), .Z(n299) );
  AND U412 ( .A(n298), .B(n299), .Z(n2106) );
  XOR U413 ( .A(sreg[338]), .B(n2240), .Z(n300) );
  NANDN U414 ( .A(n2241), .B(n300), .Z(n301) );
  NAND U415 ( .A(sreg[338]), .B(n2240), .Z(n302) );
  AND U416 ( .A(n301), .B(n302), .Z(n2280) );
  XOR U417 ( .A(sreg[343]), .B(n2351), .Z(n303) );
  NANDN U418 ( .A(n2352), .B(n303), .Z(n304) );
  NAND U419 ( .A(sreg[343]), .B(n2351), .Z(n305) );
  AND U420 ( .A(n304), .B(n305), .Z(n2391) );
  NAND U421 ( .A(n2438), .B(n2437), .Z(n306) );
  XOR U422 ( .A(n2437), .B(n2438), .Z(n307) );
  NAND U423 ( .A(n307), .B(sreg[347]), .Z(n308) );
  NAND U424 ( .A(n306), .B(n308), .Z(n2459) );
  NAND U425 ( .A(sreg[352]), .B(n2563), .Z(n309) );
  XOR U426 ( .A(n2563), .B(sreg[352]), .Z(n310) );
  NANDN U427 ( .A(n2564), .B(n310), .Z(n311) );
  NAND U428 ( .A(n309), .B(n311), .Z(n2566) );
  XOR U429 ( .A(n2629), .B(n2628), .Z(n312) );
  NANDN U430 ( .A(sreg[356]), .B(n312), .Z(n313) );
  NAND U431 ( .A(n2629), .B(n2628), .Z(n314) );
  AND U432 ( .A(n313), .B(n314), .Z(n2667) );
  XOR U433 ( .A(sreg[366]), .B(n2852), .Z(n315) );
  NANDN U434 ( .A(n2853), .B(n315), .Z(n316) );
  NAND U435 ( .A(sreg[366]), .B(n2852), .Z(n317) );
  AND U436 ( .A(n316), .B(n317), .Z(n2892) );
  XOR U437 ( .A(sreg[371]), .B(n2963), .Z(n318) );
  NANDN U438 ( .A(n2964), .B(n318), .Z(n319) );
  NAND U439 ( .A(sreg[371]), .B(n2963), .Z(n320) );
  AND U440 ( .A(n319), .B(n320), .Z(n3002) );
  XOR U441 ( .A(sreg[375]), .B(n3051), .Z(n321) );
  NANDN U442 ( .A(n3052), .B(n321), .Z(n322) );
  NAND U443 ( .A(sreg[375]), .B(n3051), .Z(n323) );
  AND U444 ( .A(n322), .B(n323), .Z(n3072) );
  XOR U445 ( .A(sreg[379]), .B(n3141), .Z(n324) );
  NANDN U446 ( .A(n3142), .B(n324), .Z(n325) );
  NAND U447 ( .A(sreg[379]), .B(n3141), .Z(n326) );
  AND U448 ( .A(n325), .B(n326), .Z(n3181) );
  XOR U449 ( .A(sreg[383]), .B(n3231), .Z(n327) );
  NANDN U450 ( .A(n3232), .B(n327), .Z(n328) );
  NAND U451 ( .A(sreg[383]), .B(n3231), .Z(n329) );
  AND U452 ( .A(n328), .B(n329), .Z(n3271) );
  XOR U453 ( .A(sreg[387]), .B(n3317), .Z(n330) );
  NANDN U454 ( .A(n3318), .B(n330), .Z(n331) );
  NAND U455 ( .A(sreg[387]), .B(n3317), .Z(n332) );
  AND U456 ( .A(n331), .B(n332), .Z(n3357) );
  NAND U457 ( .A(n3450), .B(n3449), .Z(n333) );
  XOR U458 ( .A(n3449), .B(n3450), .Z(n334) );
  NAND U459 ( .A(n334), .B(sreg[393]), .Z(n335) );
  NAND U460 ( .A(n333), .B(n335), .Z(n3488) );
  NAND U461 ( .A(n3584), .B(n3583), .Z(n336) );
  XOR U462 ( .A(n3583), .B(n3584), .Z(n337) );
  NAND U463 ( .A(n337), .B(sreg[399]), .Z(n338) );
  NAND U464 ( .A(n336), .B(n338), .Z(n3622) );
  XOR U465 ( .A(n3718), .B(sreg[405]), .Z(n339) );
  NAND U466 ( .A(n339), .B(n3717), .Z(n340) );
  NAND U467 ( .A(n3718), .B(sreg[405]), .Z(n341) );
  AND U468 ( .A(n340), .B(n341), .Z(n3757) );
  NAND U469 ( .A(n3808), .B(n3807), .Z(n342) );
  XOR U470 ( .A(n3807), .B(n3808), .Z(n343) );
  NAND U471 ( .A(n343), .B(sreg[409]), .Z(n344) );
  NAND U472 ( .A(n342), .B(n344), .Z(n3846) );
  XOR U473 ( .A(sreg[413]), .B(n3895), .Z(n345) );
  NANDN U474 ( .A(n3896), .B(n345), .Z(n346) );
  NAND U475 ( .A(sreg[413]), .B(n3895), .Z(n347) );
  AND U476 ( .A(n346), .B(n347), .Z(n3935) );
  XOR U477 ( .A(sreg[418]), .B(n4006), .Z(n348) );
  NANDN U478 ( .A(n4007), .B(n348), .Z(n349) );
  NAND U479 ( .A(sreg[418]), .B(n4006), .Z(n350) );
  AND U480 ( .A(n349), .B(n350), .Z(n4046) );
  NAND U481 ( .A(n4159), .B(sreg[424]), .Z(n351) );
  XOR U482 ( .A(sreg[424]), .B(n4159), .Z(n352) );
  NANDN U483 ( .A(n4158), .B(n352), .Z(n353) );
  NAND U484 ( .A(n351), .B(n353), .Z(n4179) );
  XOR U485 ( .A(sreg[428]), .B(n4226), .Z(n354) );
  NANDN U486 ( .A(n4227), .B(n354), .Z(n355) );
  NAND U487 ( .A(sreg[428]), .B(n4226), .Z(n356) );
  AND U488 ( .A(n355), .B(n356), .Z(n4263) );
  NAND U489 ( .A(n4331), .B(sreg[433]), .Z(n357) );
  XOR U490 ( .A(sreg[433]), .B(n4331), .Z(n358) );
  NANDN U491 ( .A(n4332), .B(n358), .Z(n359) );
  NAND U492 ( .A(n357), .B(n359), .Z(n4370) );
  XOR U493 ( .A(n4556), .B(sreg[443]), .Z(n360) );
  NAND U494 ( .A(n360), .B(n4555), .Z(n361) );
  NAND U495 ( .A(n4556), .B(sreg[443]), .Z(n362) );
  AND U496 ( .A(n361), .B(n362), .Z(n4595) );
  XOR U497 ( .A(n4707), .B(sreg[449]), .Z(n363) );
  NANDN U498 ( .A(n4708), .B(n363), .Z(n364) );
  NAND U499 ( .A(n4707), .B(sreg[449]), .Z(n365) );
  AND U500 ( .A(n364), .B(n365), .Z(n4710) );
  XOR U501 ( .A(n4776), .B(sreg[453]), .Z(n366) );
  NAND U502 ( .A(n366), .B(n4775), .Z(n367) );
  NAND U503 ( .A(n4776), .B(sreg[453]), .Z(n368) );
  AND U504 ( .A(n367), .B(n368), .Z(n4797) );
  XOR U505 ( .A(n4885), .B(n4884), .Z(n369) );
  NANDN U506 ( .A(sreg[458]), .B(n369), .Z(n370) );
  NAND U507 ( .A(n4885), .B(n4884), .Z(n371) );
  AND U508 ( .A(n370), .B(n371), .Z(n4923) );
  XOR U509 ( .A(n4973), .B(sreg[462]), .Z(n372) );
  NAND U510 ( .A(n372), .B(n4972), .Z(n373) );
  NAND U511 ( .A(n4973), .B(sreg[462]), .Z(n374) );
  AND U512 ( .A(n373), .B(n374), .Z(n5012) );
  NAND U513 ( .A(n5061), .B(n5060), .Z(n375) );
  XOR U514 ( .A(n5060), .B(n5061), .Z(n376) );
  NANDN U515 ( .A(sreg[466]), .B(n376), .Z(n377) );
  NAND U516 ( .A(n375), .B(n377), .Z(n5100) );
  NAND U517 ( .A(n5147), .B(n5146), .Z(n378) );
  XOR U518 ( .A(n5146), .B(n5147), .Z(n379) );
  NAND U519 ( .A(n379), .B(sreg[470]), .Z(n380) );
  NAND U520 ( .A(n378), .B(n380), .Z(n5185) );
  NAND U521 ( .A(n5233), .B(n5232), .Z(n381) );
  XOR U522 ( .A(n5232), .B(n5233), .Z(n382) );
  NAND U523 ( .A(n382), .B(sreg[474]), .Z(n383) );
  NAND U524 ( .A(n381), .B(n383), .Z(n5271) );
  NAND U525 ( .A(n5367), .B(n5366), .Z(n384) );
  XOR U526 ( .A(n5366), .B(n5367), .Z(n385) );
  NANDN U527 ( .A(sreg[480]), .B(n385), .Z(n386) );
  NAND U528 ( .A(n384), .B(n386), .Z(n5406) );
  XOR U529 ( .A(sreg[484]), .B(n5454), .Z(n387) );
  NANDN U530 ( .A(n5455), .B(n387), .Z(n388) );
  NAND U531 ( .A(sreg[484]), .B(n5454), .Z(n389) );
  AND U532 ( .A(n388), .B(n389), .Z(n5494) );
  NAND U533 ( .A(n5612), .B(n5611), .Z(n390) );
  XOR U534 ( .A(n5611), .B(n5612), .Z(n391) );
  NAND U535 ( .A(n391), .B(sreg[491]), .Z(n392) );
  NAND U536 ( .A(n390), .B(n392), .Z(n5651) );
  XOR U537 ( .A(n5740), .B(sreg[497]), .Z(n393) );
  NAND U538 ( .A(n393), .B(n5739), .Z(n394) );
  NAND U539 ( .A(n5740), .B(sreg[497]), .Z(n395) );
  AND U540 ( .A(n394), .B(n395), .Z(n5779) );
  NAND U541 ( .A(n5872), .B(sreg[503]), .Z(n396) );
  XOR U542 ( .A(sreg[503]), .B(n5872), .Z(n397) );
  NANDN U543 ( .A(n5871), .B(n397), .Z(n398) );
  NAND U544 ( .A(n396), .B(n398), .Z(n5908) );
  IV U545 ( .A(b[1]), .Z(n399) );
  IV U546 ( .A(b[3]), .Z(n400) );
  NAND U547 ( .A(b[0]), .B(a[0]), .Z(n408) );
  XNOR U548 ( .A(n408), .B(sreg[252]), .Z(c[252]) );
  AND U549 ( .A(a[1]), .B(b[0]), .Z(n402) );
  NAND U550 ( .A(b[1]), .B(a[0]), .Z(n401) );
  XNOR U551 ( .A(n402), .B(n401), .Z(n403) );
  XNOR U552 ( .A(sreg[253]), .B(n403), .Z(n405) );
  NANDN U553 ( .A(n408), .B(sreg[252]), .Z(n404) );
  XOR U554 ( .A(n405), .B(n404), .Z(c[253]) );
  NAND U555 ( .A(n403), .B(sreg[253]), .Z(n407) );
  OR U556 ( .A(n405), .B(n404), .Z(n406) );
  AND U557 ( .A(n407), .B(n406), .Z(n417) );
  ANDN U558 ( .B(a[1]), .A(n399), .Z(n428) );
  ANDN U559 ( .B(n428), .A(n408), .Z(n414) );
  AND U560 ( .A(b[2]), .B(a[0]), .Z(n413) );
  NAND U561 ( .A(b[0]), .B(a[2]), .Z(n429) );
  XOR U562 ( .A(n429), .B(n428), .Z(n412) );
  XNOR U563 ( .A(n413), .B(n412), .Z(n415) );
  XOR U564 ( .A(n414), .B(n415), .Z(n416) );
  XNOR U565 ( .A(sreg[254]), .B(n416), .Z(n409) );
  XOR U566 ( .A(n417), .B(n409), .Z(c[254]) );
  ANDN U567 ( .B(a[2]), .A(n445), .Z(n410) );
  NAND U568 ( .A(b[1]), .B(n410), .Z(n431) );
  NAND U569 ( .A(b[3]), .B(a[0]), .Z(n430) );
  XOR U570 ( .A(n431), .B(n430), .Z(n418) );
  AND U571 ( .A(a[3]), .B(b[0]), .Z(n452) );
  NAND U572 ( .A(b[2]), .B(a[1]), .Z(n411) );
  XNOR U573 ( .A(n452), .B(n411), .Z(n419) );
  XNOR U574 ( .A(n418), .B(n419), .Z(n421) );
  XNOR U575 ( .A(n421), .B(n420), .Z(n435) );
  XOR U576 ( .A(n434), .B(sreg[255]), .Z(n436) );
  XNOR U577 ( .A(n435), .B(n436), .Z(c[255]) );
  NAND U578 ( .A(n419), .B(n418), .Z(n423) );
  NANDN U579 ( .A(n421), .B(n420), .Z(n422) );
  NAND U580 ( .A(n423), .B(n422), .Z(n442) );
  AND U581 ( .A(b[2]), .B(a[3]), .Z(n472) );
  NAND U582 ( .A(b[0]), .B(n472), .Z(n424) );
  XNOR U583 ( .A(b[3]), .B(n424), .Z(n425) );
  NAND U584 ( .A(a[1]), .B(n425), .Z(n449) );
  XNOR U585 ( .A(n448), .B(n449), .Z(n454) );
  AND U586 ( .A(a[4]), .B(b[0]), .Z(n427) );
  NAND U587 ( .A(b[1]), .B(a[3]), .Z(n426) );
  XNOR U588 ( .A(n427), .B(n426), .Z(n453) );
  XNOR U589 ( .A(n454), .B(n453), .Z(n439) );
  NANDN U590 ( .A(n429), .B(n428), .Z(n433) );
  OR U591 ( .A(n431), .B(n430), .Z(n432) );
  NAND U592 ( .A(n433), .B(n432), .Z(n440) );
  XOR U593 ( .A(n439), .B(n440), .Z(n441) );
  XOR U594 ( .A(n442), .B(n441), .Z(n457) );
  XNOR U595 ( .A(n457), .B(sreg[256]), .Z(n459) );
  NANDN U596 ( .A(n434), .B(sreg[255]), .Z(n438) );
  NANDN U597 ( .A(n436), .B(n435), .Z(n437) );
  AND U598 ( .A(n438), .B(n437), .Z(n458) );
  XOR U599 ( .A(n459), .B(n458), .Z(c[256]) );
  OR U600 ( .A(n440), .B(n439), .Z(n444) );
  NANDN U601 ( .A(n442), .B(n441), .Z(n443) );
  NAND U602 ( .A(n444), .B(n443), .Z(n466) );
  ANDN U603 ( .B(a[4]), .A(n399), .Z(n469) );
  AND U604 ( .A(b[3]), .B(a[2]), .Z(n470) );
  XNOR U605 ( .A(n472), .B(n471), .Z(n475) );
  NAND U606 ( .A(b[0]), .B(a[5]), .Z(n476) );
  XOR U607 ( .A(n475), .B(n476), .Z(n477) );
  NAND U608 ( .A(n472), .B(n445), .Z(n447) );
  NAND U609 ( .A(b[3]), .B(a[1]), .Z(n446) );
  AND U610 ( .A(n447), .B(n446), .Z(n451) );
  NANDN U611 ( .A(n449), .B(n448), .Z(n450) );
  NANDN U612 ( .A(n451), .B(n450), .Z(n478) );
  XOR U613 ( .A(n477), .B(n478), .Z(n463) );
  NAND U614 ( .A(n469), .B(n452), .Z(n456) );
  NANDN U615 ( .A(n454), .B(n453), .Z(n455) );
  NAND U616 ( .A(n456), .B(n455), .Z(n464) );
  XNOR U617 ( .A(n463), .B(n464), .Z(n465) );
  XOR U618 ( .A(n466), .B(n465), .Z(n482) );
  NAND U619 ( .A(n457), .B(sreg[256]), .Z(n461) );
  OR U620 ( .A(n459), .B(n458), .Z(n460) );
  NAND U621 ( .A(n461), .B(n460), .Z(n481) );
  XNOR U622 ( .A(sreg[257]), .B(n481), .Z(n462) );
  XOR U623 ( .A(n482), .B(n462), .Z(c[257]) );
  NANDN U624 ( .A(n464), .B(n463), .Z(n468) );
  NAND U625 ( .A(n466), .B(n465), .Z(n467) );
  NAND U626 ( .A(n468), .B(n467), .Z(n489) );
  AND U627 ( .A(b[2]), .B(a[4]), .Z(n495) );
  AND U628 ( .A(a[5]), .B(b[1]), .Z(n493) );
  AND U629 ( .A(a[3]), .B(b[3]), .Z(n492) );
  XOR U630 ( .A(n493), .B(n492), .Z(n494) );
  XOR U631 ( .A(n495), .B(n494), .Z(n498) );
  NAND U632 ( .A(b[0]), .B(a[6]), .Z(n499) );
  XOR U633 ( .A(n498), .B(n499), .Z(n501) );
  OR U634 ( .A(n470), .B(n469), .Z(n474) );
  NANDN U635 ( .A(n472), .B(n471), .Z(n473) );
  NAND U636 ( .A(n474), .B(n473), .Z(n500) );
  XNOR U637 ( .A(n501), .B(n500), .Z(n486) );
  OR U638 ( .A(n476), .B(n475), .Z(n480) );
  NANDN U639 ( .A(n478), .B(n477), .Z(n479) );
  NAND U640 ( .A(n480), .B(n479), .Z(n487) );
  XNOR U641 ( .A(n486), .B(n487), .Z(n488) );
  XNOR U642 ( .A(n489), .B(n488), .Z(n485) );
  XOR U643 ( .A(n484), .B(sreg[258]), .Z(n483) );
  XOR U644 ( .A(n485), .B(n483), .Z(c[258]) );
  NANDN U645 ( .A(n487), .B(n486), .Z(n491) );
  NAND U646 ( .A(n489), .B(n488), .Z(n490) );
  NAND U647 ( .A(n491), .B(n490), .Z(n507) );
  AND U648 ( .A(b[2]), .B(a[5]), .Z(n513) );
  AND U649 ( .A(a[6]), .B(b[1]), .Z(n511) );
  AND U650 ( .A(a[4]), .B(b[3]), .Z(n510) );
  XOR U651 ( .A(n511), .B(n510), .Z(n512) );
  XOR U652 ( .A(n513), .B(n512), .Z(n516) );
  NAND U653 ( .A(b[0]), .B(a[7]), .Z(n517) );
  XOR U654 ( .A(n516), .B(n517), .Z(n519) );
  OR U655 ( .A(n493), .B(n492), .Z(n497) );
  NANDN U656 ( .A(n495), .B(n494), .Z(n496) );
  NAND U657 ( .A(n497), .B(n496), .Z(n518) );
  XNOR U658 ( .A(n519), .B(n518), .Z(n504) );
  NANDN U659 ( .A(n499), .B(n498), .Z(n503) );
  OR U660 ( .A(n501), .B(n500), .Z(n502) );
  NAND U661 ( .A(n503), .B(n502), .Z(n505) );
  XNOR U662 ( .A(n504), .B(n505), .Z(n506) );
  XNOR U663 ( .A(n507), .B(n506), .Z(n522) );
  XNOR U664 ( .A(n522), .B(sreg[259]), .Z(n524) );
  XNOR U665 ( .A(n523), .B(n524), .Z(c[259]) );
  NANDN U666 ( .A(n505), .B(n504), .Z(n509) );
  NAND U667 ( .A(n507), .B(n506), .Z(n508) );
  NAND U668 ( .A(n509), .B(n508), .Z(n533) );
  AND U669 ( .A(b[2]), .B(a[6]), .Z(n539) );
  AND U670 ( .A(a[7]), .B(b[1]), .Z(n537) );
  AND U671 ( .A(a[5]), .B(b[3]), .Z(n536) );
  XOR U672 ( .A(n537), .B(n536), .Z(n538) );
  XOR U673 ( .A(n539), .B(n538), .Z(n542) );
  NAND U674 ( .A(b[0]), .B(a[8]), .Z(n543) );
  XOR U675 ( .A(n542), .B(n543), .Z(n545) );
  OR U676 ( .A(n511), .B(n510), .Z(n515) );
  NANDN U677 ( .A(n513), .B(n512), .Z(n514) );
  NAND U678 ( .A(n515), .B(n514), .Z(n544) );
  XNOR U679 ( .A(n545), .B(n544), .Z(n530) );
  NANDN U680 ( .A(n517), .B(n516), .Z(n521) );
  OR U681 ( .A(n519), .B(n518), .Z(n520) );
  NAND U682 ( .A(n521), .B(n520), .Z(n531) );
  XNOR U683 ( .A(n530), .B(n531), .Z(n532) );
  XOR U684 ( .A(n533), .B(n532), .Z(n529) );
  NAND U685 ( .A(n522), .B(sreg[259]), .Z(n526) );
  NANDN U686 ( .A(n524), .B(n523), .Z(n525) );
  NAND U687 ( .A(n526), .B(n525), .Z(n528) );
  XNOR U688 ( .A(sreg[260]), .B(n528), .Z(n527) );
  XOR U689 ( .A(n529), .B(n527), .Z(c[260]) );
  NANDN U690 ( .A(n531), .B(n530), .Z(n535) );
  NAND U691 ( .A(n533), .B(n532), .Z(n534) );
  NAND U692 ( .A(n535), .B(n534), .Z(n551) );
  AND U693 ( .A(b[2]), .B(a[7]), .Z(n557) );
  AND U694 ( .A(a[8]), .B(b[1]), .Z(n555) );
  AND U695 ( .A(a[6]), .B(b[3]), .Z(n554) );
  XOR U696 ( .A(n555), .B(n554), .Z(n556) );
  XOR U697 ( .A(n557), .B(n556), .Z(n560) );
  NAND U698 ( .A(b[0]), .B(a[9]), .Z(n561) );
  XOR U699 ( .A(n560), .B(n561), .Z(n563) );
  OR U700 ( .A(n537), .B(n536), .Z(n541) );
  NANDN U701 ( .A(n539), .B(n538), .Z(n540) );
  NAND U702 ( .A(n541), .B(n540), .Z(n562) );
  XNOR U703 ( .A(n563), .B(n562), .Z(n548) );
  NANDN U704 ( .A(n543), .B(n542), .Z(n547) );
  OR U705 ( .A(n545), .B(n544), .Z(n546) );
  NAND U706 ( .A(n547), .B(n546), .Z(n549) );
  XNOR U707 ( .A(n548), .B(n549), .Z(n550) );
  XNOR U708 ( .A(n551), .B(n550), .Z(n566) );
  XNOR U709 ( .A(n566), .B(sreg[261]), .Z(n567) );
  XOR U710 ( .A(n568), .B(n567), .Z(c[261]) );
  NANDN U711 ( .A(n549), .B(n548), .Z(n553) );
  NAND U712 ( .A(n551), .B(n550), .Z(n552) );
  NAND U713 ( .A(n553), .B(n552), .Z(n575) );
  AND U714 ( .A(b[2]), .B(a[8]), .Z(n581) );
  AND U715 ( .A(a[9]), .B(b[1]), .Z(n579) );
  AND U716 ( .A(a[7]), .B(b[3]), .Z(n578) );
  XOR U717 ( .A(n579), .B(n578), .Z(n580) );
  XOR U718 ( .A(n581), .B(n580), .Z(n584) );
  NAND U719 ( .A(b[0]), .B(a[10]), .Z(n585) );
  XOR U720 ( .A(n584), .B(n585), .Z(n587) );
  OR U721 ( .A(n555), .B(n554), .Z(n559) );
  NANDN U722 ( .A(n557), .B(n556), .Z(n558) );
  NAND U723 ( .A(n559), .B(n558), .Z(n586) );
  XNOR U724 ( .A(n587), .B(n586), .Z(n572) );
  NANDN U725 ( .A(n561), .B(n560), .Z(n565) );
  OR U726 ( .A(n563), .B(n562), .Z(n564) );
  NAND U727 ( .A(n565), .B(n564), .Z(n573) );
  XNOR U728 ( .A(n572), .B(n573), .Z(n574) );
  XOR U729 ( .A(n575), .B(n574), .Z(n591) );
  NAND U730 ( .A(n566), .B(sreg[261]), .Z(n570) );
  OR U731 ( .A(n568), .B(n567), .Z(n569) );
  NAND U732 ( .A(n570), .B(n569), .Z(n590) );
  XNOR U733 ( .A(sreg[262]), .B(n590), .Z(n571) );
  XOR U734 ( .A(n591), .B(n571), .Z(c[262]) );
  NANDN U735 ( .A(n573), .B(n572), .Z(n577) );
  NAND U736 ( .A(n575), .B(n574), .Z(n576) );
  NAND U737 ( .A(n577), .B(n576), .Z(n598) );
  AND U738 ( .A(b[2]), .B(a[9]), .Z(n604) );
  AND U739 ( .A(a[10]), .B(b[1]), .Z(n602) );
  AND U740 ( .A(a[8]), .B(b[3]), .Z(n601) );
  XOR U741 ( .A(n602), .B(n601), .Z(n603) );
  XOR U742 ( .A(n604), .B(n603), .Z(n607) );
  NAND U743 ( .A(b[0]), .B(a[11]), .Z(n608) );
  XOR U744 ( .A(n607), .B(n608), .Z(n610) );
  OR U745 ( .A(n579), .B(n578), .Z(n583) );
  NANDN U746 ( .A(n581), .B(n580), .Z(n582) );
  NAND U747 ( .A(n583), .B(n582), .Z(n609) );
  XNOR U748 ( .A(n610), .B(n609), .Z(n595) );
  NANDN U749 ( .A(n585), .B(n584), .Z(n589) );
  OR U750 ( .A(n587), .B(n586), .Z(n588) );
  NAND U751 ( .A(n589), .B(n588), .Z(n596) );
  XNOR U752 ( .A(n595), .B(n596), .Z(n597) );
  XNOR U753 ( .A(n598), .B(n597), .Z(n594) );
  XOR U754 ( .A(n593), .B(sreg[263]), .Z(n592) );
  XOR U755 ( .A(n594), .B(n592), .Z(c[263]) );
  NANDN U756 ( .A(n596), .B(n595), .Z(n600) );
  NAND U757 ( .A(n598), .B(n597), .Z(n599) );
  NAND U758 ( .A(n600), .B(n599), .Z(n616) );
  AND U759 ( .A(b[2]), .B(a[10]), .Z(n622) );
  AND U760 ( .A(a[11]), .B(b[1]), .Z(n620) );
  AND U761 ( .A(a[9]), .B(b[3]), .Z(n619) );
  XOR U762 ( .A(n620), .B(n619), .Z(n621) );
  XOR U763 ( .A(n622), .B(n621), .Z(n625) );
  NAND U764 ( .A(b[0]), .B(a[12]), .Z(n626) );
  XOR U765 ( .A(n625), .B(n626), .Z(n628) );
  OR U766 ( .A(n602), .B(n601), .Z(n606) );
  NANDN U767 ( .A(n604), .B(n603), .Z(n605) );
  NAND U768 ( .A(n606), .B(n605), .Z(n627) );
  XNOR U769 ( .A(n628), .B(n627), .Z(n613) );
  NANDN U770 ( .A(n608), .B(n607), .Z(n612) );
  OR U771 ( .A(n610), .B(n609), .Z(n611) );
  NAND U772 ( .A(n612), .B(n611), .Z(n614) );
  XNOR U773 ( .A(n613), .B(n614), .Z(n615) );
  XNOR U774 ( .A(n616), .B(n615), .Z(n631) );
  XNOR U775 ( .A(n631), .B(sreg[264]), .Z(n633) );
  XNOR U776 ( .A(n632), .B(n633), .Z(c[264]) );
  NANDN U777 ( .A(n614), .B(n613), .Z(n618) );
  NAND U778 ( .A(n616), .B(n615), .Z(n617) );
  NAND U779 ( .A(n618), .B(n617), .Z(n639) );
  AND U780 ( .A(b[2]), .B(a[11]), .Z(n645) );
  AND U781 ( .A(a[12]), .B(b[1]), .Z(n643) );
  AND U782 ( .A(a[10]), .B(b[3]), .Z(n642) );
  XOR U783 ( .A(n643), .B(n642), .Z(n644) );
  XOR U784 ( .A(n645), .B(n644), .Z(n648) );
  NAND U785 ( .A(b[0]), .B(a[13]), .Z(n649) );
  XOR U786 ( .A(n648), .B(n649), .Z(n651) );
  OR U787 ( .A(n620), .B(n619), .Z(n624) );
  NANDN U788 ( .A(n622), .B(n621), .Z(n623) );
  NAND U789 ( .A(n624), .B(n623), .Z(n650) );
  XNOR U790 ( .A(n651), .B(n650), .Z(n636) );
  NANDN U791 ( .A(n626), .B(n625), .Z(n630) );
  OR U792 ( .A(n628), .B(n627), .Z(n629) );
  NAND U793 ( .A(n630), .B(n629), .Z(n637) );
  XNOR U794 ( .A(n636), .B(n637), .Z(n638) );
  XNOR U795 ( .A(n639), .B(n638), .Z(n654) );
  XOR U796 ( .A(sreg[265]), .B(n654), .Z(n655) );
  NAND U797 ( .A(n631), .B(sreg[264]), .Z(n635) );
  NANDN U798 ( .A(n633), .B(n632), .Z(n634) );
  NAND U799 ( .A(n635), .B(n634), .Z(n656) );
  XOR U800 ( .A(n655), .B(n656), .Z(c[265]) );
  NANDN U801 ( .A(n637), .B(n636), .Z(n641) );
  NAND U802 ( .A(n639), .B(n638), .Z(n640) );
  NAND U803 ( .A(n641), .B(n640), .Z(n665) );
  AND U804 ( .A(b[2]), .B(a[12]), .Z(n671) );
  AND U805 ( .A(a[13]), .B(b[1]), .Z(n669) );
  AND U806 ( .A(a[11]), .B(b[3]), .Z(n668) );
  XOR U807 ( .A(n669), .B(n668), .Z(n670) );
  XOR U808 ( .A(n671), .B(n670), .Z(n674) );
  NAND U809 ( .A(b[0]), .B(a[14]), .Z(n675) );
  XOR U810 ( .A(n674), .B(n675), .Z(n677) );
  OR U811 ( .A(n643), .B(n642), .Z(n647) );
  NANDN U812 ( .A(n645), .B(n644), .Z(n646) );
  NAND U813 ( .A(n647), .B(n646), .Z(n676) );
  XNOR U814 ( .A(n677), .B(n676), .Z(n662) );
  NANDN U815 ( .A(n649), .B(n648), .Z(n653) );
  OR U816 ( .A(n651), .B(n650), .Z(n652) );
  NAND U817 ( .A(n653), .B(n652), .Z(n663) );
  XNOR U818 ( .A(n662), .B(n663), .Z(n664) );
  XOR U819 ( .A(n665), .B(n664), .Z(n661) );
  OR U820 ( .A(n654), .B(sreg[265]), .Z(n658) );
  NANDN U821 ( .A(n656), .B(n655), .Z(n657) );
  AND U822 ( .A(n658), .B(n657), .Z(n660) );
  XNOR U823 ( .A(sreg[266]), .B(n660), .Z(n659) );
  XOR U824 ( .A(n661), .B(n659), .Z(c[266]) );
  NANDN U825 ( .A(n663), .B(n662), .Z(n667) );
  NAND U826 ( .A(n665), .B(n664), .Z(n666) );
  NAND U827 ( .A(n667), .B(n666), .Z(n695) );
  AND U828 ( .A(b[2]), .B(a[13]), .Z(n689) );
  AND U829 ( .A(a[14]), .B(b[1]), .Z(n687) );
  AND U830 ( .A(a[12]), .B(b[3]), .Z(n686) );
  XOR U831 ( .A(n687), .B(n686), .Z(n688) );
  XOR U832 ( .A(n689), .B(n688), .Z(n680) );
  NAND U833 ( .A(b[0]), .B(a[15]), .Z(n681) );
  XOR U834 ( .A(n680), .B(n681), .Z(n683) );
  OR U835 ( .A(n669), .B(n668), .Z(n673) );
  NANDN U836 ( .A(n671), .B(n670), .Z(n672) );
  NAND U837 ( .A(n673), .B(n672), .Z(n682) );
  XNOR U838 ( .A(n683), .B(n682), .Z(n692) );
  NANDN U839 ( .A(n675), .B(n674), .Z(n679) );
  OR U840 ( .A(n677), .B(n676), .Z(n678) );
  NAND U841 ( .A(n679), .B(n678), .Z(n693) );
  XNOR U842 ( .A(n692), .B(n693), .Z(n694) );
  XNOR U843 ( .A(n695), .B(n694), .Z(n698) );
  XNOR U844 ( .A(n698), .B(sreg[267]), .Z(n699) );
  XOR U845 ( .A(n700), .B(n699), .Z(c[267]) );
  NANDN U846 ( .A(n681), .B(n680), .Z(n685) );
  OR U847 ( .A(n683), .B(n682), .Z(n684) );
  NAND U848 ( .A(n685), .B(n684), .Z(n704) );
  AND U849 ( .A(b[2]), .B(a[14]), .Z(n713) );
  AND U850 ( .A(a[15]), .B(b[1]), .Z(n711) );
  AND U851 ( .A(a[13]), .B(b[3]), .Z(n710) );
  XOR U852 ( .A(n711), .B(n710), .Z(n712) );
  XOR U853 ( .A(n713), .B(n712), .Z(n716) );
  NAND U854 ( .A(b[0]), .B(a[16]), .Z(n717) );
  XNOR U855 ( .A(n716), .B(n717), .Z(n718) );
  OR U856 ( .A(n687), .B(n686), .Z(n691) );
  NANDN U857 ( .A(n689), .B(n688), .Z(n690) );
  AND U858 ( .A(n691), .B(n690), .Z(n719) );
  XNOR U859 ( .A(n718), .B(n719), .Z(n705) );
  XNOR U860 ( .A(n704), .B(n705), .Z(n706) );
  NANDN U861 ( .A(n693), .B(n692), .Z(n697) );
  NAND U862 ( .A(n695), .B(n694), .Z(n696) );
  NAND U863 ( .A(n697), .B(n696), .Z(n707) );
  XOR U864 ( .A(n706), .B(n707), .Z(n723) );
  NAND U865 ( .A(n698), .B(sreg[267]), .Z(n702) );
  OR U866 ( .A(n700), .B(n699), .Z(n701) );
  AND U867 ( .A(n702), .B(n701), .Z(n722) );
  XNOR U868 ( .A(n722), .B(sreg[268]), .Z(n703) );
  XNOR U869 ( .A(n723), .B(n703), .Z(c[268]) );
  NANDN U870 ( .A(n705), .B(n704), .Z(n709) );
  NANDN U871 ( .A(n707), .B(n706), .Z(n708) );
  NAND U872 ( .A(n709), .B(n708), .Z(n728) );
  AND U873 ( .A(b[2]), .B(a[15]), .Z(n734) );
  AND U874 ( .A(a[16]), .B(b[1]), .Z(n732) );
  AND U875 ( .A(a[14]), .B(b[3]), .Z(n731) );
  XOR U876 ( .A(n732), .B(n731), .Z(n733) );
  XOR U877 ( .A(n734), .B(n733), .Z(n737) );
  NAND U878 ( .A(b[0]), .B(a[17]), .Z(n738) );
  XOR U879 ( .A(n737), .B(n738), .Z(n740) );
  OR U880 ( .A(n711), .B(n710), .Z(n715) );
  NANDN U881 ( .A(n713), .B(n712), .Z(n714) );
  NAND U882 ( .A(n715), .B(n714), .Z(n739) );
  XNOR U883 ( .A(n740), .B(n739), .Z(n725) );
  NANDN U884 ( .A(n717), .B(n716), .Z(n721) );
  NAND U885 ( .A(n719), .B(n718), .Z(n720) );
  NAND U886 ( .A(n721), .B(n720), .Z(n726) );
  XNOR U887 ( .A(n725), .B(n726), .Z(n727) );
  XOR U888 ( .A(n728), .B(n727), .Z(n744) );
  XOR U889 ( .A(sreg[269]), .B(n743), .Z(n724) );
  XNOR U890 ( .A(n744), .B(n724), .Z(c[269]) );
  NANDN U891 ( .A(n726), .B(n725), .Z(n730) );
  NANDN U892 ( .A(n728), .B(n727), .Z(n729) );
  NAND U893 ( .A(n730), .B(n729), .Z(n751) );
  AND U894 ( .A(b[2]), .B(a[16]), .Z(n757) );
  AND U895 ( .A(a[17]), .B(b[1]), .Z(n755) );
  AND U896 ( .A(a[15]), .B(b[3]), .Z(n754) );
  XOR U897 ( .A(n755), .B(n754), .Z(n756) );
  XOR U898 ( .A(n757), .B(n756), .Z(n760) );
  NAND U899 ( .A(b[0]), .B(a[18]), .Z(n761) );
  XOR U900 ( .A(n760), .B(n761), .Z(n763) );
  OR U901 ( .A(n732), .B(n731), .Z(n736) );
  NANDN U902 ( .A(n734), .B(n733), .Z(n735) );
  NAND U903 ( .A(n736), .B(n735), .Z(n762) );
  XNOR U904 ( .A(n763), .B(n762), .Z(n748) );
  NANDN U905 ( .A(n738), .B(n737), .Z(n742) );
  OR U906 ( .A(n740), .B(n739), .Z(n741) );
  NAND U907 ( .A(n742), .B(n741), .Z(n749) );
  XNOR U908 ( .A(n748), .B(n749), .Z(n750) );
  XOR U909 ( .A(n751), .B(n750), .Z(n747) );
  XNOR U910 ( .A(sreg[270]), .B(n746), .Z(n745) );
  XOR U911 ( .A(n747), .B(n745), .Z(c[270]) );
  NANDN U912 ( .A(n749), .B(n748), .Z(n753) );
  NAND U913 ( .A(n751), .B(n750), .Z(n752) );
  NAND U914 ( .A(n753), .B(n752), .Z(n769) );
  AND U915 ( .A(b[2]), .B(a[17]), .Z(n775) );
  AND U916 ( .A(a[18]), .B(b[1]), .Z(n773) );
  AND U917 ( .A(a[16]), .B(b[3]), .Z(n772) );
  XOR U918 ( .A(n773), .B(n772), .Z(n774) );
  XOR U919 ( .A(n775), .B(n774), .Z(n778) );
  NAND U920 ( .A(b[0]), .B(a[19]), .Z(n779) );
  XOR U921 ( .A(n778), .B(n779), .Z(n781) );
  OR U922 ( .A(n755), .B(n754), .Z(n759) );
  NANDN U923 ( .A(n757), .B(n756), .Z(n758) );
  NAND U924 ( .A(n759), .B(n758), .Z(n780) );
  XNOR U925 ( .A(n781), .B(n780), .Z(n766) );
  NANDN U926 ( .A(n761), .B(n760), .Z(n765) );
  OR U927 ( .A(n763), .B(n762), .Z(n764) );
  NAND U928 ( .A(n765), .B(n764), .Z(n767) );
  XNOR U929 ( .A(n766), .B(n767), .Z(n768) );
  XNOR U930 ( .A(n769), .B(n768), .Z(n784) );
  XNOR U931 ( .A(n784), .B(sreg[271]), .Z(n785) );
  XOR U932 ( .A(n786), .B(n785), .Z(c[271]) );
  NANDN U933 ( .A(n767), .B(n766), .Z(n771) );
  NAND U934 ( .A(n769), .B(n768), .Z(n770) );
  NAND U935 ( .A(n771), .B(n770), .Z(n792) );
  AND U936 ( .A(b[2]), .B(a[18]), .Z(n798) );
  AND U937 ( .A(a[19]), .B(b[1]), .Z(n796) );
  AND U938 ( .A(a[17]), .B(b[3]), .Z(n795) );
  XOR U939 ( .A(n796), .B(n795), .Z(n797) );
  XOR U940 ( .A(n798), .B(n797), .Z(n801) );
  NAND U941 ( .A(b[0]), .B(a[20]), .Z(n802) );
  XOR U942 ( .A(n801), .B(n802), .Z(n804) );
  OR U943 ( .A(n773), .B(n772), .Z(n777) );
  NANDN U944 ( .A(n775), .B(n774), .Z(n776) );
  NAND U945 ( .A(n777), .B(n776), .Z(n803) );
  XNOR U946 ( .A(n804), .B(n803), .Z(n789) );
  NANDN U947 ( .A(n779), .B(n778), .Z(n783) );
  OR U948 ( .A(n781), .B(n780), .Z(n782) );
  NAND U949 ( .A(n783), .B(n782), .Z(n790) );
  XNOR U950 ( .A(n789), .B(n790), .Z(n791) );
  XNOR U951 ( .A(n792), .B(n791), .Z(n807) );
  XOR U952 ( .A(sreg[272]), .B(n807), .Z(n808) );
  NAND U953 ( .A(n784), .B(sreg[271]), .Z(n788) );
  OR U954 ( .A(n786), .B(n785), .Z(n787) );
  NAND U955 ( .A(n788), .B(n787), .Z(n809) );
  XOR U956 ( .A(n808), .B(n809), .Z(c[272]) );
  NANDN U957 ( .A(n790), .B(n789), .Z(n794) );
  NAND U958 ( .A(n792), .B(n791), .Z(n793) );
  NAND U959 ( .A(n794), .B(n793), .Z(n816) );
  AND U960 ( .A(b[2]), .B(a[19]), .Z(n822) );
  AND U961 ( .A(a[20]), .B(b[1]), .Z(n820) );
  AND U962 ( .A(a[18]), .B(b[3]), .Z(n819) );
  XOR U963 ( .A(n820), .B(n819), .Z(n821) );
  XOR U964 ( .A(n822), .B(n821), .Z(n825) );
  NAND U965 ( .A(b[0]), .B(a[21]), .Z(n826) );
  XOR U966 ( .A(n825), .B(n826), .Z(n828) );
  OR U967 ( .A(n796), .B(n795), .Z(n800) );
  NANDN U968 ( .A(n798), .B(n797), .Z(n799) );
  NAND U969 ( .A(n800), .B(n799), .Z(n827) );
  XNOR U970 ( .A(n828), .B(n827), .Z(n813) );
  NANDN U971 ( .A(n802), .B(n801), .Z(n806) );
  OR U972 ( .A(n804), .B(n803), .Z(n805) );
  NAND U973 ( .A(n806), .B(n805), .Z(n814) );
  XNOR U974 ( .A(n813), .B(n814), .Z(n815) );
  XOR U975 ( .A(n816), .B(n815), .Z(n832) );
  OR U976 ( .A(n807), .B(sreg[272]), .Z(n811) );
  NANDN U977 ( .A(n809), .B(n808), .Z(n810) );
  AND U978 ( .A(n811), .B(n810), .Z(n831) );
  XNOR U979 ( .A(sreg[273]), .B(n831), .Z(n812) );
  XOR U980 ( .A(n832), .B(n812), .Z(c[273]) );
  NANDN U981 ( .A(n814), .B(n813), .Z(n818) );
  NAND U982 ( .A(n816), .B(n815), .Z(n817) );
  NAND U983 ( .A(n818), .B(n817), .Z(n839) );
  AND U984 ( .A(b[2]), .B(a[20]), .Z(n845) );
  AND U985 ( .A(a[21]), .B(b[1]), .Z(n843) );
  AND U986 ( .A(a[19]), .B(b[3]), .Z(n842) );
  XOR U987 ( .A(n843), .B(n842), .Z(n844) );
  XOR U988 ( .A(n845), .B(n844), .Z(n848) );
  NAND U989 ( .A(b[0]), .B(a[22]), .Z(n849) );
  XOR U990 ( .A(n848), .B(n849), .Z(n851) );
  OR U991 ( .A(n820), .B(n819), .Z(n824) );
  NANDN U992 ( .A(n822), .B(n821), .Z(n823) );
  NAND U993 ( .A(n824), .B(n823), .Z(n850) );
  XNOR U994 ( .A(n851), .B(n850), .Z(n836) );
  NANDN U995 ( .A(n826), .B(n825), .Z(n830) );
  OR U996 ( .A(n828), .B(n827), .Z(n829) );
  NAND U997 ( .A(n830), .B(n829), .Z(n837) );
  XNOR U998 ( .A(n836), .B(n837), .Z(n838) );
  XNOR U999 ( .A(n839), .B(n838), .Z(n835) );
  XOR U1000 ( .A(n834), .B(sreg[274]), .Z(n833) );
  XOR U1001 ( .A(n835), .B(n833), .Z(c[274]) );
  NANDN U1002 ( .A(n837), .B(n836), .Z(n841) );
  NAND U1003 ( .A(n839), .B(n838), .Z(n840) );
  NAND U1004 ( .A(n841), .B(n840), .Z(n857) );
  AND U1005 ( .A(b[2]), .B(a[21]), .Z(n863) );
  AND U1006 ( .A(a[22]), .B(b[1]), .Z(n861) );
  AND U1007 ( .A(a[20]), .B(b[3]), .Z(n860) );
  XOR U1008 ( .A(n861), .B(n860), .Z(n862) );
  XOR U1009 ( .A(n863), .B(n862), .Z(n866) );
  NAND U1010 ( .A(b[0]), .B(a[23]), .Z(n867) );
  XOR U1011 ( .A(n866), .B(n867), .Z(n869) );
  OR U1012 ( .A(n843), .B(n842), .Z(n847) );
  NANDN U1013 ( .A(n845), .B(n844), .Z(n846) );
  NAND U1014 ( .A(n847), .B(n846), .Z(n868) );
  XNOR U1015 ( .A(n869), .B(n868), .Z(n854) );
  NANDN U1016 ( .A(n849), .B(n848), .Z(n853) );
  OR U1017 ( .A(n851), .B(n850), .Z(n852) );
  NAND U1018 ( .A(n853), .B(n852), .Z(n855) );
  XNOR U1019 ( .A(n854), .B(n855), .Z(n856) );
  XNOR U1020 ( .A(n857), .B(n856), .Z(n872) );
  XNOR U1021 ( .A(n872), .B(sreg[275]), .Z(n874) );
  XNOR U1022 ( .A(n873), .B(n874), .Z(c[275]) );
  NANDN U1023 ( .A(n855), .B(n854), .Z(n859) );
  NAND U1024 ( .A(n857), .B(n856), .Z(n858) );
  NAND U1025 ( .A(n859), .B(n858), .Z(n881) );
  AND U1026 ( .A(b[2]), .B(a[22]), .Z(n887) );
  AND U1027 ( .A(a[23]), .B(b[1]), .Z(n885) );
  AND U1028 ( .A(a[21]), .B(b[3]), .Z(n884) );
  XOR U1029 ( .A(n885), .B(n884), .Z(n886) );
  XOR U1030 ( .A(n887), .B(n886), .Z(n890) );
  NAND U1031 ( .A(b[0]), .B(a[24]), .Z(n891) );
  XOR U1032 ( .A(n890), .B(n891), .Z(n893) );
  OR U1033 ( .A(n861), .B(n860), .Z(n865) );
  NANDN U1034 ( .A(n863), .B(n862), .Z(n864) );
  NAND U1035 ( .A(n865), .B(n864), .Z(n892) );
  XNOR U1036 ( .A(n893), .B(n892), .Z(n878) );
  NANDN U1037 ( .A(n867), .B(n866), .Z(n871) );
  OR U1038 ( .A(n869), .B(n868), .Z(n870) );
  NAND U1039 ( .A(n871), .B(n870), .Z(n879) );
  XNOR U1040 ( .A(n878), .B(n879), .Z(n880) );
  XNOR U1041 ( .A(n881), .B(n880), .Z(n897) );
  NAND U1042 ( .A(n872), .B(sreg[275]), .Z(n876) );
  NANDN U1043 ( .A(n874), .B(n873), .Z(n875) );
  AND U1044 ( .A(n876), .B(n875), .Z(n896) );
  XNOR U1045 ( .A(n896), .B(sreg[276]), .Z(n877) );
  XOR U1046 ( .A(n897), .B(n877), .Z(c[276]) );
  NANDN U1047 ( .A(n879), .B(n878), .Z(n883) );
  NAND U1048 ( .A(n881), .B(n880), .Z(n882) );
  NAND U1049 ( .A(n883), .B(n882), .Z(n904) );
  AND U1050 ( .A(b[2]), .B(a[23]), .Z(n910) );
  AND U1051 ( .A(a[24]), .B(b[1]), .Z(n908) );
  AND U1052 ( .A(a[22]), .B(b[3]), .Z(n907) );
  XOR U1053 ( .A(n908), .B(n907), .Z(n909) );
  XOR U1054 ( .A(n910), .B(n909), .Z(n913) );
  NAND U1055 ( .A(b[0]), .B(a[25]), .Z(n914) );
  XOR U1056 ( .A(n913), .B(n914), .Z(n916) );
  OR U1057 ( .A(n885), .B(n884), .Z(n889) );
  NANDN U1058 ( .A(n887), .B(n886), .Z(n888) );
  NAND U1059 ( .A(n889), .B(n888), .Z(n915) );
  XNOR U1060 ( .A(n916), .B(n915), .Z(n901) );
  NANDN U1061 ( .A(n891), .B(n890), .Z(n895) );
  OR U1062 ( .A(n893), .B(n892), .Z(n894) );
  NAND U1063 ( .A(n895), .B(n894), .Z(n902) );
  XNOR U1064 ( .A(n901), .B(n902), .Z(n903) );
  XNOR U1065 ( .A(n904), .B(n903), .Z(n900) );
  XOR U1066 ( .A(n899), .B(sreg[277]), .Z(n898) );
  XOR U1067 ( .A(n900), .B(n898), .Z(c[277]) );
  NANDN U1068 ( .A(n902), .B(n901), .Z(n906) );
  NAND U1069 ( .A(n904), .B(n903), .Z(n905) );
  NAND U1070 ( .A(n906), .B(n905), .Z(n922) );
  AND U1071 ( .A(b[2]), .B(a[24]), .Z(n928) );
  AND U1072 ( .A(a[25]), .B(b[1]), .Z(n926) );
  AND U1073 ( .A(a[23]), .B(b[3]), .Z(n925) );
  XOR U1074 ( .A(n926), .B(n925), .Z(n927) );
  XOR U1075 ( .A(n928), .B(n927), .Z(n931) );
  NAND U1076 ( .A(b[0]), .B(a[26]), .Z(n932) );
  XOR U1077 ( .A(n931), .B(n932), .Z(n934) );
  OR U1078 ( .A(n908), .B(n907), .Z(n912) );
  NANDN U1079 ( .A(n910), .B(n909), .Z(n911) );
  NAND U1080 ( .A(n912), .B(n911), .Z(n933) );
  XNOR U1081 ( .A(n934), .B(n933), .Z(n919) );
  NANDN U1082 ( .A(n914), .B(n913), .Z(n918) );
  OR U1083 ( .A(n916), .B(n915), .Z(n917) );
  NAND U1084 ( .A(n918), .B(n917), .Z(n920) );
  XNOR U1085 ( .A(n919), .B(n920), .Z(n921) );
  XNOR U1086 ( .A(n922), .B(n921), .Z(n937) );
  XNOR U1087 ( .A(n937), .B(sreg[278]), .Z(n939) );
  XNOR U1088 ( .A(n938), .B(n939), .Z(c[278]) );
  NANDN U1089 ( .A(n920), .B(n919), .Z(n924) );
  NAND U1090 ( .A(n922), .B(n921), .Z(n923) );
  NAND U1091 ( .A(n924), .B(n923), .Z(n948) );
  AND U1092 ( .A(b[2]), .B(a[25]), .Z(n954) );
  AND U1093 ( .A(a[26]), .B(b[1]), .Z(n952) );
  AND U1094 ( .A(a[24]), .B(b[3]), .Z(n951) );
  XOR U1095 ( .A(n952), .B(n951), .Z(n953) );
  XOR U1096 ( .A(n954), .B(n953), .Z(n957) );
  NAND U1097 ( .A(b[0]), .B(a[27]), .Z(n958) );
  XOR U1098 ( .A(n957), .B(n958), .Z(n960) );
  OR U1099 ( .A(n926), .B(n925), .Z(n930) );
  NANDN U1100 ( .A(n928), .B(n927), .Z(n929) );
  NAND U1101 ( .A(n930), .B(n929), .Z(n959) );
  XNOR U1102 ( .A(n960), .B(n959), .Z(n945) );
  NANDN U1103 ( .A(n932), .B(n931), .Z(n936) );
  OR U1104 ( .A(n934), .B(n933), .Z(n935) );
  NAND U1105 ( .A(n936), .B(n935), .Z(n946) );
  XNOR U1106 ( .A(n945), .B(n946), .Z(n947) );
  XNOR U1107 ( .A(n948), .B(n947), .Z(n944) );
  NAND U1108 ( .A(n937), .B(sreg[278]), .Z(n941) );
  NANDN U1109 ( .A(n939), .B(n938), .Z(n940) );
  AND U1110 ( .A(n941), .B(n940), .Z(n943) );
  XNOR U1111 ( .A(n943), .B(sreg[279]), .Z(n942) );
  XOR U1112 ( .A(n944), .B(n942), .Z(c[279]) );
  NANDN U1113 ( .A(n946), .B(n945), .Z(n950) );
  NAND U1114 ( .A(n948), .B(n947), .Z(n949) );
  NAND U1115 ( .A(n950), .B(n949), .Z(n966) );
  AND U1116 ( .A(b[2]), .B(a[26]), .Z(n972) );
  AND U1117 ( .A(a[27]), .B(b[1]), .Z(n970) );
  AND U1118 ( .A(a[25]), .B(b[3]), .Z(n969) );
  XOR U1119 ( .A(n970), .B(n969), .Z(n971) );
  XOR U1120 ( .A(n972), .B(n971), .Z(n975) );
  NAND U1121 ( .A(b[0]), .B(a[28]), .Z(n976) );
  XOR U1122 ( .A(n975), .B(n976), .Z(n978) );
  OR U1123 ( .A(n952), .B(n951), .Z(n956) );
  NANDN U1124 ( .A(n954), .B(n953), .Z(n955) );
  NAND U1125 ( .A(n956), .B(n955), .Z(n977) );
  XNOR U1126 ( .A(n978), .B(n977), .Z(n963) );
  NANDN U1127 ( .A(n958), .B(n957), .Z(n962) );
  OR U1128 ( .A(n960), .B(n959), .Z(n961) );
  NAND U1129 ( .A(n962), .B(n961), .Z(n964) );
  XNOR U1130 ( .A(n963), .B(n964), .Z(n965) );
  XNOR U1131 ( .A(n966), .B(n965), .Z(n981) );
  XOR U1132 ( .A(sreg[280]), .B(n981), .Z(n982) );
  XOR U1133 ( .A(n983), .B(n982), .Z(c[280]) );
  NANDN U1134 ( .A(n964), .B(n963), .Z(n968) );
  NAND U1135 ( .A(n966), .B(n965), .Z(n967) );
  NAND U1136 ( .A(n968), .B(n967), .Z(n989) );
  AND U1137 ( .A(b[2]), .B(a[27]), .Z(n995) );
  AND U1138 ( .A(a[28]), .B(b[1]), .Z(n993) );
  AND U1139 ( .A(a[26]), .B(b[3]), .Z(n992) );
  XOR U1140 ( .A(n993), .B(n992), .Z(n994) );
  XOR U1141 ( .A(n995), .B(n994), .Z(n998) );
  NAND U1142 ( .A(b[0]), .B(a[29]), .Z(n999) );
  XOR U1143 ( .A(n998), .B(n999), .Z(n1001) );
  OR U1144 ( .A(n970), .B(n969), .Z(n974) );
  NANDN U1145 ( .A(n972), .B(n971), .Z(n973) );
  NAND U1146 ( .A(n974), .B(n973), .Z(n1000) );
  XNOR U1147 ( .A(n1001), .B(n1000), .Z(n986) );
  NANDN U1148 ( .A(n976), .B(n975), .Z(n980) );
  OR U1149 ( .A(n978), .B(n977), .Z(n979) );
  NAND U1150 ( .A(n980), .B(n979), .Z(n987) );
  XNOR U1151 ( .A(n986), .B(n987), .Z(n988) );
  XNOR U1152 ( .A(n989), .B(n988), .Z(n1004) );
  XNOR U1153 ( .A(n1004), .B(sreg[281]), .Z(n1006) );
  OR U1154 ( .A(n981), .B(sreg[280]), .Z(n985) );
  NANDN U1155 ( .A(n983), .B(n982), .Z(n984) );
  NAND U1156 ( .A(n985), .B(n984), .Z(n1005) );
  XOR U1157 ( .A(n1006), .B(n1005), .Z(c[281]) );
  NANDN U1158 ( .A(n987), .B(n986), .Z(n991) );
  NAND U1159 ( .A(n989), .B(n988), .Z(n990) );
  NAND U1160 ( .A(n991), .B(n990), .Z(n1015) );
  AND U1161 ( .A(b[2]), .B(a[28]), .Z(n1021) );
  AND U1162 ( .A(a[29]), .B(b[1]), .Z(n1019) );
  AND U1163 ( .A(a[27]), .B(b[3]), .Z(n1018) );
  XOR U1164 ( .A(n1019), .B(n1018), .Z(n1020) );
  XOR U1165 ( .A(n1021), .B(n1020), .Z(n1024) );
  NAND U1166 ( .A(b[0]), .B(a[30]), .Z(n1025) );
  XOR U1167 ( .A(n1024), .B(n1025), .Z(n1027) );
  OR U1168 ( .A(n993), .B(n992), .Z(n997) );
  NANDN U1169 ( .A(n995), .B(n994), .Z(n996) );
  NAND U1170 ( .A(n997), .B(n996), .Z(n1026) );
  XNOR U1171 ( .A(n1027), .B(n1026), .Z(n1012) );
  NANDN U1172 ( .A(n999), .B(n998), .Z(n1003) );
  OR U1173 ( .A(n1001), .B(n1000), .Z(n1002) );
  NAND U1174 ( .A(n1003), .B(n1002), .Z(n1013) );
  XNOR U1175 ( .A(n1012), .B(n1013), .Z(n1014) );
  XNOR U1176 ( .A(n1015), .B(n1014), .Z(n1011) );
  NAND U1177 ( .A(n1004), .B(sreg[281]), .Z(n1008) );
  OR U1178 ( .A(n1006), .B(n1005), .Z(n1007) );
  AND U1179 ( .A(n1008), .B(n1007), .Z(n1010) );
  XNOR U1180 ( .A(n1010), .B(sreg[282]), .Z(n1009) );
  XOR U1181 ( .A(n1011), .B(n1009), .Z(c[282]) );
  NANDN U1182 ( .A(n1013), .B(n1012), .Z(n1017) );
  NAND U1183 ( .A(n1015), .B(n1014), .Z(n1016) );
  NAND U1184 ( .A(n1017), .B(n1016), .Z(n1033) );
  AND U1185 ( .A(b[2]), .B(a[29]), .Z(n1039) );
  AND U1186 ( .A(a[30]), .B(b[1]), .Z(n1037) );
  AND U1187 ( .A(a[28]), .B(b[3]), .Z(n1036) );
  XOR U1188 ( .A(n1037), .B(n1036), .Z(n1038) );
  XOR U1189 ( .A(n1039), .B(n1038), .Z(n1042) );
  NAND U1190 ( .A(b[0]), .B(a[31]), .Z(n1043) );
  XOR U1191 ( .A(n1042), .B(n1043), .Z(n1045) );
  OR U1192 ( .A(n1019), .B(n1018), .Z(n1023) );
  NANDN U1193 ( .A(n1021), .B(n1020), .Z(n1022) );
  NAND U1194 ( .A(n1023), .B(n1022), .Z(n1044) );
  XNOR U1195 ( .A(n1045), .B(n1044), .Z(n1030) );
  NANDN U1196 ( .A(n1025), .B(n1024), .Z(n1029) );
  OR U1197 ( .A(n1027), .B(n1026), .Z(n1028) );
  NAND U1198 ( .A(n1029), .B(n1028), .Z(n1031) );
  XNOR U1199 ( .A(n1030), .B(n1031), .Z(n1032) );
  XNOR U1200 ( .A(n1033), .B(n1032), .Z(n1048) );
  XNOR U1201 ( .A(n1048), .B(sreg[283]), .Z(n1050) );
  XNOR U1202 ( .A(n1049), .B(n1050), .Z(c[283]) );
  NANDN U1203 ( .A(n1031), .B(n1030), .Z(n1035) );
  NAND U1204 ( .A(n1033), .B(n1032), .Z(n1034) );
  NAND U1205 ( .A(n1035), .B(n1034), .Z(n1056) );
  AND U1206 ( .A(b[2]), .B(a[30]), .Z(n1068) );
  AND U1207 ( .A(a[31]), .B(b[1]), .Z(n1066) );
  AND U1208 ( .A(a[29]), .B(b[3]), .Z(n1065) );
  XOR U1209 ( .A(n1066), .B(n1065), .Z(n1067) );
  XOR U1210 ( .A(n1068), .B(n1067), .Z(n1059) );
  NAND U1211 ( .A(b[0]), .B(a[32]), .Z(n1060) );
  XOR U1212 ( .A(n1059), .B(n1060), .Z(n1062) );
  OR U1213 ( .A(n1037), .B(n1036), .Z(n1041) );
  NANDN U1214 ( .A(n1039), .B(n1038), .Z(n1040) );
  NAND U1215 ( .A(n1041), .B(n1040), .Z(n1061) );
  XNOR U1216 ( .A(n1062), .B(n1061), .Z(n1053) );
  NANDN U1217 ( .A(n1043), .B(n1042), .Z(n1047) );
  OR U1218 ( .A(n1045), .B(n1044), .Z(n1046) );
  NAND U1219 ( .A(n1047), .B(n1046), .Z(n1054) );
  XNOR U1220 ( .A(n1053), .B(n1054), .Z(n1055) );
  XNOR U1221 ( .A(n1056), .B(n1055), .Z(n1072) );
  XOR U1222 ( .A(sreg[284]), .B(n1072), .Z(n1073) );
  NAND U1223 ( .A(n1048), .B(sreg[283]), .Z(n1052) );
  NANDN U1224 ( .A(n1050), .B(n1049), .Z(n1051) );
  NAND U1225 ( .A(n1052), .B(n1051), .Z(n1074) );
  XOR U1226 ( .A(n1073), .B(n1074), .Z(c[284]) );
  NANDN U1227 ( .A(n1054), .B(n1053), .Z(n1058) );
  NAND U1228 ( .A(n1056), .B(n1055), .Z(n1057) );
  AND U1229 ( .A(n1058), .B(n1057), .Z(n1080) );
  NANDN U1230 ( .A(n1060), .B(n1059), .Z(n1064) );
  OR U1231 ( .A(n1062), .B(n1061), .Z(n1063) );
  AND U1232 ( .A(n1064), .B(n1063), .Z(n1079) );
  AND U1233 ( .A(b[2]), .B(a[31]), .Z(n1084) );
  AND U1234 ( .A(a[32]), .B(b[1]), .Z(n1082) );
  AND U1235 ( .A(a[30]), .B(b[3]), .Z(n1081) );
  XOR U1236 ( .A(n1082), .B(n1081), .Z(n1083) );
  XOR U1237 ( .A(n1084), .B(n1083), .Z(n1087) );
  NAND U1238 ( .A(b[0]), .B(a[33]), .Z(n1088) );
  XOR U1239 ( .A(n1087), .B(n1088), .Z(n1090) );
  OR U1240 ( .A(n1066), .B(n1065), .Z(n1070) );
  NANDN U1241 ( .A(n1068), .B(n1067), .Z(n1069) );
  NAND U1242 ( .A(n1070), .B(n1069), .Z(n1089) );
  XOR U1243 ( .A(n1090), .B(n1089), .Z(n1078) );
  XNOR U1244 ( .A(n1079), .B(n1078), .Z(n1071) );
  XOR U1245 ( .A(n1080), .B(n1071), .Z(n1094) );
  OR U1246 ( .A(n1072), .B(sreg[284]), .Z(n1076) );
  NANDN U1247 ( .A(n1074), .B(n1073), .Z(n1075) );
  AND U1248 ( .A(n1076), .B(n1075), .Z(n1093) );
  XNOR U1249 ( .A(sreg[285]), .B(n1093), .Z(n1077) );
  XNOR U1250 ( .A(n1094), .B(n1077), .Z(c[285]) );
  AND U1251 ( .A(b[2]), .B(a[32]), .Z(n1107) );
  AND U1252 ( .A(a[33]), .B(b[1]), .Z(n1105) );
  AND U1253 ( .A(a[31]), .B(b[3]), .Z(n1104) );
  XOR U1254 ( .A(n1105), .B(n1104), .Z(n1106) );
  XOR U1255 ( .A(n1107), .B(n1106), .Z(n1110) );
  NAND U1256 ( .A(b[0]), .B(a[34]), .Z(n1111) );
  XOR U1257 ( .A(n1110), .B(n1111), .Z(n1113) );
  OR U1258 ( .A(n1082), .B(n1081), .Z(n1086) );
  NANDN U1259 ( .A(n1084), .B(n1083), .Z(n1085) );
  NAND U1260 ( .A(n1086), .B(n1085), .Z(n1112) );
  XNOR U1261 ( .A(n1113), .B(n1112), .Z(n1098) );
  NANDN U1262 ( .A(n1088), .B(n1087), .Z(n1092) );
  OR U1263 ( .A(n1090), .B(n1089), .Z(n1091) );
  NAND U1264 ( .A(n1092), .B(n1091), .Z(n1099) );
  XNOR U1265 ( .A(n1098), .B(n1099), .Z(n1100) );
  XNOR U1266 ( .A(n1101), .B(n1100), .Z(n1097) );
  XOR U1267 ( .A(n1096), .B(sreg[286]), .Z(n1095) );
  XNOR U1268 ( .A(n1097), .B(n1095), .Z(c[286]) );
  NANDN U1269 ( .A(n1099), .B(n1098), .Z(n1103) );
  NANDN U1270 ( .A(n1101), .B(n1100), .Z(n1102) );
  NAND U1271 ( .A(n1103), .B(n1102), .Z(n1119) );
  AND U1272 ( .A(b[2]), .B(a[33]), .Z(n1125) );
  AND U1273 ( .A(a[34]), .B(b[1]), .Z(n1123) );
  AND U1274 ( .A(a[32]), .B(b[3]), .Z(n1122) );
  XOR U1275 ( .A(n1123), .B(n1122), .Z(n1124) );
  XOR U1276 ( .A(n1125), .B(n1124), .Z(n1128) );
  NAND U1277 ( .A(b[0]), .B(a[35]), .Z(n1129) );
  XOR U1278 ( .A(n1128), .B(n1129), .Z(n1131) );
  OR U1279 ( .A(n1105), .B(n1104), .Z(n1109) );
  NANDN U1280 ( .A(n1107), .B(n1106), .Z(n1108) );
  NAND U1281 ( .A(n1109), .B(n1108), .Z(n1130) );
  XNOR U1282 ( .A(n1131), .B(n1130), .Z(n1116) );
  NANDN U1283 ( .A(n1111), .B(n1110), .Z(n1115) );
  OR U1284 ( .A(n1113), .B(n1112), .Z(n1114) );
  NAND U1285 ( .A(n1115), .B(n1114), .Z(n1117) );
  XNOR U1286 ( .A(n1116), .B(n1117), .Z(n1118) );
  XNOR U1287 ( .A(n1119), .B(n1118), .Z(n1135) );
  XOR U1288 ( .A(sreg[287]), .B(n1135), .Z(n1136) );
  XOR U1289 ( .A(n1137), .B(n1136), .Z(c[287]) );
  NANDN U1290 ( .A(n1117), .B(n1116), .Z(n1121) );
  NAND U1291 ( .A(n1119), .B(n1118), .Z(n1120) );
  AND U1292 ( .A(n1121), .B(n1120), .Z(n1145) );
  AND U1293 ( .A(b[2]), .B(a[34]), .Z(n1153) );
  AND U1294 ( .A(a[35]), .B(b[1]), .Z(n1151) );
  AND U1295 ( .A(a[33]), .B(b[3]), .Z(n1150) );
  XOR U1296 ( .A(n1151), .B(n1150), .Z(n1152) );
  XOR U1297 ( .A(n1153), .B(n1152), .Z(n1146) );
  NAND U1298 ( .A(b[0]), .B(a[36]), .Z(n1147) );
  XOR U1299 ( .A(n1146), .B(n1147), .Z(n1148) );
  OR U1300 ( .A(n1123), .B(n1122), .Z(n1127) );
  NANDN U1301 ( .A(n1125), .B(n1124), .Z(n1126) );
  AND U1302 ( .A(n1127), .B(n1126), .Z(n1149) );
  XOR U1303 ( .A(n1148), .B(n1149), .Z(n1143) );
  NANDN U1304 ( .A(n1129), .B(n1128), .Z(n1133) );
  OR U1305 ( .A(n1131), .B(n1130), .Z(n1132) );
  AND U1306 ( .A(n1133), .B(n1132), .Z(n1144) );
  XOR U1307 ( .A(n1143), .B(n1144), .Z(n1134) );
  XNOR U1308 ( .A(n1145), .B(n1134), .Z(n1142) );
  OR U1309 ( .A(n1135), .B(sreg[287]), .Z(n1139) );
  NANDN U1310 ( .A(n1137), .B(n1136), .Z(n1138) );
  AND U1311 ( .A(n1139), .B(n1138), .Z(n1141) );
  XNOR U1312 ( .A(sreg[288]), .B(n1141), .Z(n1140) );
  XOR U1313 ( .A(n1142), .B(n1140), .Z(c[288]) );
  AND U1314 ( .A(b[2]), .B(a[35]), .Z(n1164) );
  AND U1315 ( .A(a[36]), .B(b[1]), .Z(n1162) );
  AND U1316 ( .A(a[34]), .B(b[3]), .Z(n1161) );
  XOR U1317 ( .A(n1162), .B(n1161), .Z(n1163) );
  XOR U1318 ( .A(n1164), .B(n1163), .Z(n1167) );
  NAND U1319 ( .A(b[0]), .B(a[37]), .Z(n1168) );
  XNOR U1320 ( .A(n1167), .B(n1168), .Z(n1169) );
  OR U1321 ( .A(n1151), .B(n1150), .Z(n1155) );
  NANDN U1322 ( .A(n1153), .B(n1152), .Z(n1154) );
  AND U1323 ( .A(n1155), .B(n1154), .Z(n1170) );
  XNOR U1324 ( .A(n1169), .B(n1170), .Z(n1174) );
  XNOR U1325 ( .A(n1173), .B(n1174), .Z(n1175) );
  XNOR U1326 ( .A(n1176), .B(n1175), .Z(n1156) );
  XNOR U1327 ( .A(sreg[289]), .B(n1156), .Z(n1157) );
  XOR U1328 ( .A(n1158), .B(n1157), .Z(c[289]) );
  NAND U1329 ( .A(sreg[289]), .B(n1156), .Z(n1160) );
  OR U1330 ( .A(n1158), .B(n1157), .Z(n1159) );
  NAND U1331 ( .A(n1160), .B(n1159), .Z(n1199) );
  AND U1332 ( .A(b[2]), .B(a[36]), .Z(n1188) );
  AND U1333 ( .A(a[37]), .B(b[1]), .Z(n1186) );
  AND U1334 ( .A(a[35]), .B(b[3]), .Z(n1185) );
  XOR U1335 ( .A(n1186), .B(n1185), .Z(n1187) );
  XOR U1336 ( .A(n1188), .B(n1187), .Z(n1191) );
  NAND U1337 ( .A(b[0]), .B(a[38]), .Z(n1192) );
  XOR U1338 ( .A(n1191), .B(n1192), .Z(n1194) );
  OR U1339 ( .A(n1162), .B(n1161), .Z(n1166) );
  NANDN U1340 ( .A(n1164), .B(n1163), .Z(n1165) );
  NAND U1341 ( .A(n1166), .B(n1165), .Z(n1193) );
  XNOR U1342 ( .A(n1194), .B(n1193), .Z(n1179) );
  NANDN U1343 ( .A(n1168), .B(n1167), .Z(n1172) );
  NAND U1344 ( .A(n1170), .B(n1169), .Z(n1171) );
  NAND U1345 ( .A(n1172), .B(n1171), .Z(n1180) );
  XNOR U1346 ( .A(n1179), .B(n1180), .Z(n1181) );
  NANDN U1347 ( .A(n1174), .B(n1173), .Z(n1178) );
  NANDN U1348 ( .A(n1176), .B(n1175), .Z(n1177) );
  AND U1349 ( .A(n1178), .B(n1177), .Z(n1182) );
  XNOR U1350 ( .A(n1181), .B(n1182), .Z(n1197) );
  XOR U1351 ( .A(sreg[290]), .B(n1197), .Z(n1198) );
  XOR U1352 ( .A(n1199), .B(n1198), .Z(c[290]) );
  NANDN U1353 ( .A(n1180), .B(n1179), .Z(n1184) );
  NAND U1354 ( .A(n1182), .B(n1181), .Z(n1183) );
  NAND U1355 ( .A(n1184), .B(n1183), .Z(n1220) );
  AND U1356 ( .A(b[2]), .B(a[37]), .Z(n1214) );
  AND U1357 ( .A(a[38]), .B(b[1]), .Z(n1212) );
  AND U1358 ( .A(a[36]), .B(b[3]), .Z(n1211) );
  XOR U1359 ( .A(n1212), .B(n1211), .Z(n1213) );
  XOR U1360 ( .A(n1214), .B(n1213), .Z(n1205) );
  NAND U1361 ( .A(b[0]), .B(a[39]), .Z(n1206) );
  XOR U1362 ( .A(n1205), .B(n1206), .Z(n1208) );
  OR U1363 ( .A(n1186), .B(n1185), .Z(n1190) );
  NANDN U1364 ( .A(n1188), .B(n1187), .Z(n1189) );
  NAND U1365 ( .A(n1190), .B(n1189), .Z(n1207) );
  XNOR U1366 ( .A(n1208), .B(n1207), .Z(n1217) );
  NANDN U1367 ( .A(n1192), .B(n1191), .Z(n1196) );
  OR U1368 ( .A(n1194), .B(n1193), .Z(n1195) );
  NAND U1369 ( .A(n1196), .B(n1195), .Z(n1218) );
  XNOR U1370 ( .A(n1217), .B(n1218), .Z(n1219) );
  XOR U1371 ( .A(n1220), .B(n1219), .Z(n1204) );
  OR U1372 ( .A(n1197), .B(sreg[290]), .Z(n1201) );
  NANDN U1373 ( .A(n1199), .B(n1198), .Z(n1200) );
  AND U1374 ( .A(n1201), .B(n1200), .Z(n1203) );
  XNOR U1375 ( .A(sreg[291]), .B(n1203), .Z(n1202) );
  XOR U1376 ( .A(n1204), .B(n1202), .Z(c[291]) );
  NANDN U1377 ( .A(n1206), .B(n1205), .Z(n1210) );
  OR U1378 ( .A(n1208), .B(n1207), .Z(n1209) );
  NAND U1379 ( .A(n1210), .B(n1209), .Z(n1235) );
  AND U1380 ( .A(b[2]), .B(a[38]), .Z(n1226) );
  AND U1381 ( .A(a[39]), .B(b[1]), .Z(n1224) );
  AND U1382 ( .A(a[37]), .B(b[3]), .Z(n1223) );
  XOR U1383 ( .A(n1224), .B(n1223), .Z(n1225) );
  XOR U1384 ( .A(n1226), .B(n1225), .Z(n1229) );
  NAND U1385 ( .A(b[0]), .B(a[40]), .Z(n1230) );
  XNOR U1386 ( .A(n1229), .B(n1230), .Z(n1231) );
  OR U1387 ( .A(n1212), .B(n1211), .Z(n1216) );
  NANDN U1388 ( .A(n1214), .B(n1213), .Z(n1215) );
  AND U1389 ( .A(n1216), .B(n1215), .Z(n1232) );
  XNOR U1390 ( .A(n1231), .B(n1232), .Z(n1236) );
  XNOR U1391 ( .A(n1235), .B(n1236), .Z(n1237) );
  NANDN U1392 ( .A(n1218), .B(n1217), .Z(n1222) );
  NAND U1393 ( .A(n1220), .B(n1219), .Z(n1221) );
  AND U1394 ( .A(n1222), .B(n1221), .Z(n1238) );
  XOR U1395 ( .A(n1237), .B(n1238), .Z(n1241) );
  XNOR U1396 ( .A(sreg[292]), .B(n1241), .Z(n1242) );
  XOR U1397 ( .A(n1243), .B(n1242), .Z(c[292]) );
  AND U1398 ( .A(b[2]), .B(a[39]), .Z(n1258) );
  AND U1399 ( .A(a[40]), .B(b[1]), .Z(n1256) );
  AND U1400 ( .A(a[38]), .B(b[3]), .Z(n1255) );
  XOR U1401 ( .A(n1256), .B(n1255), .Z(n1257) );
  XOR U1402 ( .A(n1258), .B(n1257), .Z(n1261) );
  NAND U1403 ( .A(b[0]), .B(a[41]), .Z(n1262) );
  XOR U1404 ( .A(n1261), .B(n1262), .Z(n1264) );
  OR U1405 ( .A(n1224), .B(n1223), .Z(n1228) );
  NANDN U1406 ( .A(n1226), .B(n1225), .Z(n1227) );
  NAND U1407 ( .A(n1228), .B(n1227), .Z(n1263) );
  XNOR U1408 ( .A(n1264), .B(n1263), .Z(n1249) );
  NANDN U1409 ( .A(n1230), .B(n1229), .Z(n1234) );
  NAND U1410 ( .A(n1232), .B(n1231), .Z(n1233) );
  NAND U1411 ( .A(n1234), .B(n1233), .Z(n1250) );
  XNOR U1412 ( .A(n1249), .B(n1250), .Z(n1251) );
  NANDN U1413 ( .A(n1236), .B(n1235), .Z(n1240) );
  NAND U1414 ( .A(n1238), .B(n1237), .Z(n1239) );
  AND U1415 ( .A(n1240), .B(n1239), .Z(n1252) );
  XNOR U1416 ( .A(n1251), .B(n1252), .Z(n1248) );
  NAND U1417 ( .A(sreg[292]), .B(n1241), .Z(n1245) );
  OR U1418 ( .A(n1243), .B(n1242), .Z(n1244) );
  AND U1419 ( .A(n1245), .B(n1244), .Z(n1247) );
  XNOR U1420 ( .A(n1247), .B(sreg[293]), .Z(n1246) );
  XOR U1421 ( .A(n1248), .B(n1246), .Z(c[293]) );
  NANDN U1422 ( .A(n1250), .B(n1249), .Z(n1254) );
  NAND U1423 ( .A(n1252), .B(n1251), .Z(n1253) );
  NAND U1424 ( .A(n1254), .B(n1253), .Z(n1270) );
  AND U1425 ( .A(b[2]), .B(a[40]), .Z(n1276) );
  AND U1426 ( .A(a[41]), .B(b[1]), .Z(n1274) );
  AND U1427 ( .A(a[39]), .B(b[3]), .Z(n1273) );
  XOR U1428 ( .A(n1274), .B(n1273), .Z(n1275) );
  XOR U1429 ( .A(n1276), .B(n1275), .Z(n1279) );
  NAND U1430 ( .A(b[0]), .B(a[42]), .Z(n1280) );
  XOR U1431 ( .A(n1279), .B(n1280), .Z(n1282) );
  OR U1432 ( .A(n1256), .B(n1255), .Z(n1260) );
  NANDN U1433 ( .A(n1258), .B(n1257), .Z(n1259) );
  NAND U1434 ( .A(n1260), .B(n1259), .Z(n1281) );
  XNOR U1435 ( .A(n1282), .B(n1281), .Z(n1267) );
  NANDN U1436 ( .A(n1262), .B(n1261), .Z(n1266) );
  OR U1437 ( .A(n1264), .B(n1263), .Z(n1265) );
  NAND U1438 ( .A(n1266), .B(n1265), .Z(n1268) );
  XNOR U1439 ( .A(n1267), .B(n1268), .Z(n1269) );
  XNOR U1440 ( .A(n1270), .B(n1269), .Z(n1285) );
  XNOR U1441 ( .A(n1285), .B(sreg[294]), .Z(n1287) );
  XNOR U1442 ( .A(n1286), .B(n1287), .Z(c[294]) );
  NANDN U1443 ( .A(n1268), .B(n1267), .Z(n1272) );
  NAND U1444 ( .A(n1270), .B(n1269), .Z(n1271) );
  NAND U1445 ( .A(n1272), .B(n1271), .Z(n1294) );
  AND U1446 ( .A(b[2]), .B(a[41]), .Z(n1300) );
  AND U1447 ( .A(a[42]), .B(b[1]), .Z(n1298) );
  AND U1448 ( .A(a[40]), .B(b[3]), .Z(n1297) );
  XOR U1449 ( .A(n1298), .B(n1297), .Z(n1299) );
  XOR U1450 ( .A(n1300), .B(n1299), .Z(n1303) );
  NAND U1451 ( .A(b[0]), .B(a[43]), .Z(n1304) );
  XOR U1452 ( .A(n1303), .B(n1304), .Z(n1306) );
  OR U1453 ( .A(n1274), .B(n1273), .Z(n1278) );
  NANDN U1454 ( .A(n1276), .B(n1275), .Z(n1277) );
  NAND U1455 ( .A(n1278), .B(n1277), .Z(n1305) );
  XNOR U1456 ( .A(n1306), .B(n1305), .Z(n1291) );
  NANDN U1457 ( .A(n1280), .B(n1279), .Z(n1284) );
  OR U1458 ( .A(n1282), .B(n1281), .Z(n1283) );
  NAND U1459 ( .A(n1284), .B(n1283), .Z(n1292) );
  XNOR U1460 ( .A(n1291), .B(n1292), .Z(n1293) );
  XNOR U1461 ( .A(n1294), .B(n1293), .Z(n1310) );
  NAND U1462 ( .A(n1285), .B(sreg[294]), .Z(n1289) );
  NANDN U1463 ( .A(n1287), .B(n1286), .Z(n1288) );
  AND U1464 ( .A(n1289), .B(n1288), .Z(n1309) );
  XNOR U1465 ( .A(n1309), .B(sreg[295]), .Z(n1290) );
  XOR U1466 ( .A(n1310), .B(n1290), .Z(c[295]) );
  NANDN U1467 ( .A(n1292), .B(n1291), .Z(n1296) );
  NAND U1468 ( .A(n1294), .B(n1293), .Z(n1295) );
  NAND U1469 ( .A(n1296), .B(n1295), .Z(n1315) );
  AND U1470 ( .A(b[2]), .B(a[42]), .Z(n1321) );
  AND U1471 ( .A(a[43]), .B(b[1]), .Z(n1319) );
  AND U1472 ( .A(a[41]), .B(b[3]), .Z(n1318) );
  XOR U1473 ( .A(n1319), .B(n1318), .Z(n1320) );
  XOR U1474 ( .A(n1321), .B(n1320), .Z(n1324) );
  NAND U1475 ( .A(b[0]), .B(a[44]), .Z(n1325) );
  XOR U1476 ( .A(n1324), .B(n1325), .Z(n1327) );
  OR U1477 ( .A(n1298), .B(n1297), .Z(n1302) );
  NANDN U1478 ( .A(n1300), .B(n1299), .Z(n1301) );
  NAND U1479 ( .A(n1302), .B(n1301), .Z(n1326) );
  XNOR U1480 ( .A(n1327), .B(n1326), .Z(n1312) );
  NANDN U1481 ( .A(n1304), .B(n1303), .Z(n1308) );
  OR U1482 ( .A(n1306), .B(n1305), .Z(n1307) );
  NAND U1483 ( .A(n1308), .B(n1307), .Z(n1313) );
  XNOR U1484 ( .A(n1312), .B(n1313), .Z(n1314) );
  XOR U1485 ( .A(n1315), .B(n1314), .Z(n1331) );
  XOR U1486 ( .A(sreg[296]), .B(n1330), .Z(n1311) );
  XOR U1487 ( .A(n1331), .B(n1311), .Z(c[296]) );
  NANDN U1488 ( .A(n1313), .B(n1312), .Z(n1317) );
  NAND U1489 ( .A(n1315), .B(n1314), .Z(n1316) );
  NAND U1490 ( .A(n1317), .B(n1316), .Z(n1338) );
  AND U1491 ( .A(b[2]), .B(a[43]), .Z(n1344) );
  AND U1492 ( .A(a[44]), .B(b[1]), .Z(n1342) );
  AND U1493 ( .A(a[42]), .B(b[3]), .Z(n1341) );
  XOR U1494 ( .A(n1342), .B(n1341), .Z(n1343) );
  XOR U1495 ( .A(n1344), .B(n1343), .Z(n1347) );
  NAND U1496 ( .A(b[0]), .B(a[45]), .Z(n1348) );
  XOR U1497 ( .A(n1347), .B(n1348), .Z(n1350) );
  OR U1498 ( .A(n1319), .B(n1318), .Z(n1323) );
  NANDN U1499 ( .A(n1321), .B(n1320), .Z(n1322) );
  NAND U1500 ( .A(n1323), .B(n1322), .Z(n1349) );
  XNOR U1501 ( .A(n1350), .B(n1349), .Z(n1335) );
  NANDN U1502 ( .A(n1325), .B(n1324), .Z(n1329) );
  OR U1503 ( .A(n1327), .B(n1326), .Z(n1328) );
  NAND U1504 ( .A(n1329), .B(n1328), .Z(n1336) );
  XNOR U1505 ( .A(n1335), .B(n1336), .Z(n1337) );
  XOR U1506 ( .A(n1338), .B(n1337), .Z(n1334) );
  XNOR U1507 ( .A(sreg[297]), .B(n1333), .Z(n1332) );
  XOR U1508 ( .A(n1334), .B(n1332), .Z(c[297]) );
  NANDN U1509 ( .A(n1336), .B(n1335), .Z(n1340) );
  NAND U1510 ( .A(n1338), .B(n1337), .Z(n1339) );
  NAND U1511 ( .A(n1340), .B(n1339), .Z(n1356) );
  AND U1512 ( .A(b[2]), .B(a[44]), .Z(n1362) );
  AND U1513 ( .A(a[45]), .B(b[1]), .Z(n1360) );
  AND U1514 ( .A(a[43]), .B(b[3]), .Z(n1359) );
  XOR U1515 ( .A(n1360), .B(n1359), .Z(n1361) );
  XOR U1516 ( .A(n1362), .B(n1361), .Z(n1365) );
  NAND U1517 ( .A(b[0]), .B(a[46]), .Z(n1366) );
  XOR U1518 ( .A(n1365), .B(n1366), .Z(n1368) );
  OR U1519 ( .A(n1342), .B(n1341), .Z(n1346) );
  NANDN U1520 ( .A(n1344), .B(n1343), .Z(n1345) );
  NAND U1521 ( .A(n1346), .B(n1345), .Z(n1367) );
  XNOR U1522 ( .A(n1368), .B(n1367), .Z(n1353) );
  NANDN U1523 ( .A(n1348), .B(n1347), .Z(n1352) );
  OR U1524 ( .A(n1350), .B(n1349), .Z(n1351) );
  NAND U1525 ( .A(n1352), .B(n1351), .Z(n1354) );
  XNOR U1526 ( .A(n1353), .B(n1354), .Z(n1355) );
  XNOR U1527 ( .A(n1356), .B(n1355), .Z(n1371) );
  XNOR U1528 ( .A(n1371), .B(sreg[298]), .Z(n1372) );
  XOR U1529 ( .A(n1373), .B(n1372), .Z(c[298]) );
  NANDN U1530 ( .A(n1354), .B(n1353), .Z(n1358) );
  NAND U1531 ( .A(n1356), .B(n1355), .Z(n1357) );
  NAND U1532 ( .A(n1358), .B(n1357), .Z(n1382) );
  AND U1533 ( .A(b[2]), .B(a[45]), .Z(n1388) );
  AND U1534 ( .A(a[46]), .B(b[1]), .Z(n1386) );
  AND U1535 ( .A(a[44]), .B(b[3]), .Z(n1385) );
  XOR U1536 ( .A(n1386), .B(n1385), .Z(n1387) );
  XOR U1537 ( .A(n1388), .B(n1387), .Z(n1391) );
  NAND U1538 ( .A(b[0]), .B(a[47]), .Z(n1392) );
  XOR U1539 ( .A(n1391), .B(n1392), .Z(n1394) );
  OR U1540 ( .A(n1360), .B(n1359), .Z(n1364) );
  NANDN U1541 ( .A(n1362), .B(n1361), .Z(n1363) );
  NAND U1542 ( .A(n1364), .B(n1363), .Z(n1393) );
  XNOR U1543 ( .A(n1394), .B(n1393), .Z(n1379) );
  NANDN U1544 ( .A(n1366), .B(n1365), .Z(n1370) );
  OR U1545 ( .A(n1368), .B(n1367), .Z(n1369) );
  NAND U1546 ( .A(n1370), .B(n1369), .Z(n1380) );
  XNOR U1547 ( .A(n1379), .B(n1380), .Z(n1381) );
  XOR U1548 ( .A(n1382), .B(n1381), .Z(n1378) );
  NAND U1549 ( .A(n1371), .B(sreg[298]), .Z(n1375) );
  OR U1550 ( .A(n1373), .B(n1372), .Z(n1374) );
  NAND U1551 ( .A(n1375), .B(n1374), .Z(n1377) );
  XNOR U1552 ( .A(sreg[299]), .B(n1377), .Z(n1376) );
  XOR U1553 ( .A(n1378), .B(n1376), .Z(c[299]) );
  NANDN U1554 ( .A(n1380), .B(n1379), .Z(n1384) );
  NAND U1555 ( .A(n1382), .B(n1381), .Z(n1383) );
  NAND U1556 ( .A(n1384), .B(n1383), .Z(n1400) );
  AND U1557 ( .A(b[2]), .B(a[46]), .Z(n1406) );
  AND U1558 ( .A(a[47]), .B(b[1]), .Z(n1404) );
  AND U1559 ( .A(a[45]), .B(b[3]), .Z(n1403) );
  XOR U1560 ( .A(n1404), .B(n1403), .Z(n1405) );
  XOR U1561 ( .A(n1406), .B(n1405), .Z(n1409) );
  NAND U1562 ( .A(b[0]), .B(a[48]), .Z(n1410) );
  XOR U1563 ( .A(n1409), .B(n1410), .Z(n1412) );
  OR U1564 ( .A(n1386), .B(n1385), .Z(n1390) );
  NANDN U1565 ( .A(n1388), .B(n1387), .Z(n1389) );
  NAND U1566 ( .A(n1390), .B(n1389), .Z(n1411) );
  XNOR U1567 ( .A(n1412), .B(n1411), .Z(n1397) );
  NANDN U1568 ( .A(n1392), .B(n1391), .Z(n1396) );
  OR U1569 ( .A(n1394), .B(n1393), .Z(n1395) );
  NAND U1570 ( .A(n1396), .B(n1395), .Z(n1398) );
  XNOR U1571 ( .A(n1397), .B(n1398), .Z(n1399) );
  XNOR U1572 ( .A(n1400), .B(n1399), .Z(n1415) );
  XNOR U1573 ( .A(n1415), .B(sreg[300]), .Z(n1416) );
  XOR U1574 ( .A(n1417), .B(n1416), .Z(c[300]) );
  NANDN U1575 ( .A(n1398), .B(n1397), .Z(n1402) );
  NAND U1576 ( .A(n1400), .B(n1399), .Z(n1401) );
  NAND U1577 ( .A(n1402), .B(n1401), .Z(n1423) );
  AND U1578 ( .A(b[2]), .B(a[47]), .Z(n1429) );
  AND U1579 ( .A(a[48]), .B(b[1]), .Z(n1427) );
  AND U1580 ( .A(a[46]), .B(b[3]), .Z(n1426) );
  XOR U1581 ( .A(n1427), .B(n1426), .Z(n1428) );
  XOR U1582 ( .A(n1429), .B(n1428), .Z(n1432) );
  NAND U1583 ( .A(b[0]), .B(a[49]), .Z(n1433) );
  XOR U1584 ( .A(n1432), .B(n1433), .Z(n1435) );
  OR U1585 ( .A(n1404), .B(n1403), .Z(n1408) );
  NANDN U1586 ( .A(n1406), .B(n1405), .Z(n1407) );
  NAND U1587 ( .A(n1408), .B(n1407), .Z(n1434) );
  XNOR U1588 ( .A(n1435), .B(n1434), .Z(n1420) );
  NANDN U1589 ( .A(n1410), .B(n1409), .Z(n1414) );
  OR U1590 ( .A(n1412), .B(n1411), .Z(n1413) );
  NAND U1591 ( .A(n1414), .B(n1413), .Z(n1421) );
  XNOR U1592 ( .A(n1420), .B(n1421), .Z(n1422) );
  XNOR U1593 ( .A(n1423), .B(n1422), .Z(n1438) );
  XNOR U1594 ( .A(n1438), .B(sreg[301]), .Z(n1440) );
  NAND U1595 ( .A(n1415), .B(sreg[300]), .Z(n1419) );
  OR U1596 ( .A(n1417), .B(n1416), .Z(n1418) );
  AND U1597 ( .A(n1419), .B(n1418), .Z(n1439) );
  XOR U1598 ( .A(n1440), .B(n1439), .Z(c[301]) );
  NANDN U1599 ( .A(n1421), .B(n1420), .Z(n1425) );
  NAND U1600 ( .A(n1423), .B(n1422), .Z(n1424) );
  NAND U1601 ( .A(n1425), .B(n1424), .Z(n1449) );
  AND U1602 ( .A(b[2]), .B(a[48]), .Z(n1455) );
  AND U1603 ( .A(a[49]), .B(b[1]), .Z(n1453) );
  AND U1604 ( .A(a[47]), .B(b[3]), .Z(n1452) );
  XOR U1605 ( .A(n1453), .B(n1452), .Z(n1454) );
  XOR U1606 ( .A(n1455), .B(n1454), .Z(n1458) );
  NAND U1607 ( .A(b[0]), .B(a[50]), .Z(n1459) );
  XOR U1608 ( .A(n1458), .B(n1459), .Z(n1461) );
  OR U1609 ( .A(n1427), .B(n1426), .Z(n1431) );
  NANDN U1610 ( .A(n1429), .B(n1428), .Z(n1430) );
  NAND U1611 ( .A(n1431), .B(n1430), .Z(n1460) );
  XNOR U1612 ( .A(n1461), .B(n1460), .Z(n1446) );
  NANDN U1613 ( .A(n1433), .B(n1432), .Z(n1437) );
  OR U1614 ( .A(n1435), .B(n1434), .Z(n1436) );
  NAND U1615 ( .A(n1437), .B(n1436), .Z(n1447) );
  XNOR U1616 ( .A(n1446), .B(n1447), .Z(n1448) );
  XOR U1617 ( .A(n1449), .B(n1448), .Z(n1445) );
  NAND U1618 ( .A(n1438), .B(sreg[301]), .Z(n1442) );
  OR U1619 ( .A(n1440), .B(n1439), .Z(n1441) );
  NAND U1620 ( .A(n1442), .B(n1441), .Z(n1444) );
  XNOR U1621 ( .A(sreg[302]), .B(n1444), .Z(n1443) );
  XOR U1622 ( .A(n1445), .B(n1443), .Z(c[302]) );
  NANDN U1623 ( .A(n1447), .B(n1446), .Z(n1451) );
  NAND U1624 ( .A(n1449), .B(n1448), .Z(n1450) );
  NAND U1625 ( .A(n1451), .B(n1450), .Z(n1467) );
  AND U1626 ( .A(b[2]), .B(a[49]), .Z(n1473) );
  AND U1627 ( .A(a[50]), .B(b[1]), .Z(n1471) );
  AND U1628 ( .A(a[48]), .B(b[3]), .Z(n1470) );
  XOR U1629 ( .A(n1471), .B(n1470), .Z(n1472) );
  XOR U1630 ( .A(n1473), .B(n1472), .Z(n1476) );
  NAND U1631 ( .A(b[0]), .B(a[51]), .Z(n1477) );
  XOR U1632 ( .A(n1476), .B(n1477), .Z(n1479) );
  OR U1633 ( .A(n1453), .B(n1452), .Z(n1457) );
  NANDN U1634 ( .A(n1455), .B(n1454), .Z(n1456) );
  NAND U1635 ( .A(n1457), .B(n1456), .Z(n1478) );
  XNOR U1636 ( .A(n1479), .B(n1478), .Z(n1464) );
  NANDN U1637 ( .A(n1459), .B(n1458), .Z(n1463) );
  OR U1638 ( .A(n1461), .B(n1460), .Z(n1462) );
  NAND U1639 ( .A(n1463), .B(n1462), .Z(n1465) );
  XNOR U1640 ( .A(n1464), .B(n1465), .Z(n1466) );
  XNOR U1641 ( .A(n1467), .B(n1466), .Z(n1482) );
  XNOR U1642 ( .A(n1482), .B(sreg[303]), .Z(n1483) );
  XOR U1643 ( .A(n1484), .B(n1483), .Z(c[303]) );
  NANDN U1644 ( .A(n1465), .B(n1464), .Z(n1469) );
  NAND U1645 ( .A(n1467), .B(n1466), .Z(n1468) );
  NAND U1646 ( .A(n1469), .B(n1468), .Z(n1493) );
  AND U1647 ( .A(b[2]), .B(a[50]), .Z(n1499) );
  AND U1648 ( .A(a[51]), .B(b[1]), .Z(n1497) );
  AND U1649 ( .A(a[49]), .B(b[3]), .Z(n1496) );
  XOR U1650 ( .A(n1497), .B(n1496), .Z(n1498) );
  XOR U1651 ( .A(n1499), .B(n1498), .Z(n1502) );
  NAND U1652 ( .A(b[0]), .B(a[52]), .Z(n1503) );
  XOR U1653 ( .A(n1502), .B(n1503), .Z(n1505) );
  OR U1654 ( .A(n1471), .B(n1470), .Z(n1475) );
  NANDN U1655 ( .A(n1473), .B(n1472), .Z(n1474) );
  NAND U1656 ( .A(n1475), .B(n1474), .Z(n1504) );
  XNOR U1657 ( .A(n1505), .B(n1504), .Z(n1490) );
  NANDN U1658 ( .A(n1477), .B(n1476), .Z(n1481) );
  OR U1659 ( .A(n1479), .B(n1478), .Z(n1480) );
  NAND U1660 ( .A(n1481), .B(n1480), .Z(n1491) );
  XNOR U1661 ( .A(n1490), .B(n1491), .Z(n1492) );
  XOR U1662 ( .A(n1493), .B(n1492), .Z(n1489) );
  NAND U1663 ( .A(n1482), .B(sreg[303]), .Z(n1486) );
  OR U1664 ( .A(n1484), .B(n1483), .Z(n1485) );
  NAND U1665 ( .A(n1486), .B(n1485), .Z(n1488) );
  XNOR U1666 ( .A(sreg[304]), .B(n1488), .Z(n1487) );
  XOR U1667 ( .A(n1489), .B(n1487), .Z(c[304]) );
  NANDN U1668 ( .A(n1491), .B(n1490), .Z(n1495) );
  NAND U1669 ( .A(n1493), .B(n1492), .Z(n1494) );
  NAND U1670 ( .A(n1495), .B(n1494), .Z(n1511) );
  AND U1671 ( .A(b[2]), .B(a[51]), .Z(n1517) );
  AND U1672 ( .A(a[52]), .B(b[1]), .Z(n1515) );
  AND U1673 ( .A(a[50]), .B(b[3]), .Z(n1514) );
  XOR U1674 ( .A(n1515), .B(n1514), .Z(n1516) );
  XOR U1675 ( .A(n1517), .B(n1516), .Z(n1520) );
  NAND U1676 ( .A(b[0]), .B(a[53]), .Z(n1521) );
  XOR U1677 ( .A(n1520), .B(n1521), .Z(n1523) );
  OR U1678 ( .A(n1497), .B(n1496), .Z(n1501) );
  NANDN U1679 ( .A(n1499), .B(n1498), .Z(n1500) );
  NAND U1680 ( .A(n1501), .B(n1500), .Z(n1522) );
  XNOR U1681 ( .A(n1523), .B(n1522), .Z(n1508) );
  NANDN U1682 ( .A(n1503), .B(n1502), .Z(n1507) );
  OR U1683 ( .A(n1505), .B(n1504), .Z(n1506) );
  NAND U1684 ( .A(n1507), .B(n1506), .Z(n1509) );
  XNOR U1685 ( .A(n1508), .B(n1509), .Z(n1510) );
  XNOR U1686 ( .A(n1511), .B(n1510), .Z(n1526) );
  XNOR U1687 ( .A(n1526), .B(sreg[305]), .Z(n1527) );
  XOR U1688 ( .A(n1528), .B(n1527), .Z(c[305]) );
  NANDN U1689 ( .A(n1509), .B(n1508), .Z(n1513) );
  NAND U1690 ( .A(n1511), .B(n1510), .Z(n1512) );
  NAND U1691 ( .A(n1513), .B(n1512), .Z(n1537) );
  AND U1692 ( .A(b[2]), .B(a[52]), .Z(n1543) );
  AND U1693 ( .A(a[53]), .B(b[1]), .Z(n1541) );
  AND U1694 ( .A(a[51]), .B(b[3]), .Z(n1540) );
  XOR U1695 ( .A(n1541), .B(n1540), .Z(n1542) );
  XOR U1696 ( .A(n1543), .B(n1542), .Z(n1546) );
  NAND U1697 ( .A(b[0]), .B(a[54]), .Z(n1547) );
  XOR U1698 ( .A(n1546), .B(n1547), .Z(n1549) );
  OR U1699 ( .A(n1515), .B(n1514), .Z(n1519) );
  NANDN U1700 ( .A(n1517), .B(n1516), .Z(n1518) );
  NAND U1701 ( .A(n1519), .B(n1518), .Z(n1548) );
  XNOR U1702 ( .A(n1549), .B(n1548), .Z(n1534) );
  NANDN U1703 ( .A(n1521), .B(n1520), .Z(n1525) );
  OR U1704 ( .A(n1523), .B(n1522), .Z(n1524) );
  NAND U1705 ( .A(n1525), .B(n1524), .Z(n1535) );
  XNOR U1706 ( .A(n1534), .B(n1535), .Z(n1536) );
  XOR U1707 ( .A(n1537), .B(n1536), .Z(n1533) );
  NAND U1708 ( .A(n1526), .B(sreg[305]), .Z(n1530) );
  OR U1709 ( .A(n1528), .B(n1527), .Z(n1529) );
  NAND U1710 ( .A(n1530), .B(n1529), .Z(n1532) );
  XNOR U1711 ( .A(sreg[306]), .B(n1532), .Z(n1531) );
  XOR U1712 ( .A(n1533), .B(n1531), .Z(c[306]) );
  NANDN U1713 ( .A(n1535), .B(n1534), .Z(n1539) );
  NAND U1714 ( .A(n1537), .B(n1536), .Z(n1538) );
  NAND U1715 ( .A(n1539), .B(n1538), .Z(n1555) );
  AND U1716 ( .A(b[2]), .B(a[53]), .Z(n1561) );
  AND U1717 ( .A(a[54]), .B(b[1]), .Z(n1559) );
  AND U1718 ( .A(a[52]), .B(b[3]), .Z(n1558) );
  XOR U1719 ( .A(n1559), .B(n1558), .Z(n1560) );
  XOR U1720 ( .A(n1561), .B(n1560), .Z(n1564) );
  NAND U1721 ( .A(b[0]), .B(a[55]), .Z(n1565) );
  XOR U1722 ( .A(n1564), .B(n1565), .Z(n1567) );
  OR U1723 ( .A(n1541), .B(n1540), .Z(n1545) );
  NANDN U1724 ( .A(n1543), .B(n1542), .Z(n1544) );
  NAND U1725 ( .A(n1545), .B(n1544), .Z(n1566) );
  XNOR U1726 ( .A(n1567), .B(n1566), .Z(n1552) );
  NANDN U1727 ( .A(n1547), .B(n1546), .Z(n1551) );
  OR U1728 ( .A(n1549), .B(n1548), .Z(n1550) );
  NAND U1729 ( .A(n1551), .B(n1550), .Z(n1553) );
  XNOR U1730 ( .A(n1552), .B(n1553), .Z(n1554) );
  XNOR U1731 ( .A(n1555), .B(n1554), .Z(n1570) );
  XNOR U1732 ( .A(n1570), .B(sreg[307]), .Z(n1571) );
  XOR U1733 ( .A(n1572), .B(n1571), .Z(c[307]) );
  NANDN U1734 ( .A(n1553), .B(n1552), .Z(n1557) );
  NAND U1735 ( .A(n1555), .B(n1554), .Z(n1556) );
  NAND U1736 ( .A(n1557), .B(n1556), .Z(n1578) );
  AND U1737 ( .A(b[2]), .B(a[54]), .Z(n1584) );
  AND U1738 ( .A(a[55]), .B(b[1]), .Z(n1582) );
  AND U1739 ( .A(a[53]), .B(b[3]), .Z(n1581) );
  XOR U1740 ( .A(n1582), .B(n1581), .Z(n1583) );
  XOR U1741 ( .A(n1584), .B(n1583), .Z(n1587) );
  NAND U1742 ( .A(b[0]), .B(a[56]), .Z(n1588) );
  XOR U1743 ( .A(n1587), .B(n1588), .Z(n1590) );
  OR U1744 ( .A(n1559), .B(n1558), .Z(n1563) );
  NANDN U1745 ( .A(n1561), .B(n1560), .Z(n1562) );
  NAND U1746 ( .A(n1563), .B(n1562), .Z(n1589) );
  XNOR U1747 ( .A(n1590), .B(n1589), .Z(n1575) );
  NANDN U1748 ( .A(n1565), .B(n1564), .Z(n1569) );
  OR U1749 ( .A(n1567), .B(n1566), .Z(n1568) );
  NAND U1750 ( .A(n1569), .B(n1568), .Z(n1576) );
  XNOR U1751 ( .A(n1575), .B(n1576), .Z(n1577) );
  XNOR U1752 ( .A(n1578), .B(n1577), .Z(n1593) );
  XNOR U1753 ( .A(n1593), .B(sreg[308]), .Z(n1595) );
  NAND U1754 ( .A(n1570), .B(sreg[307]), .Z(n1574) );
  OR U1755 ( .A(n1572), .B(n1571), .Z(n1573) );
  AND U1756 ( .A(n1574), .B(n1573), .Z(n1594) );
  XOR U1757 ( .A(n1595), .B(n1594), .Z(c[308]) );
  NANDN U1758 ( .A(n1576), .B(n1575), .Z(n1580) );
  NAND U1759 ( .A(n1578), .B(n1577), .Z(n1579) );
  NAND U1760 ( .A(n1580), .B(n1579), .Z(n1604) );
  AND U1761 ( .A(b[2]), .B(a[55]), .Z(n1610) );
  AND U1762 ( .A(a[56]), .B(b[1]), .Z(n1608) );
  AND U1763 ( .A(a[54]), .B(b[3]), .Z(n1607) );
  XOR U1764 ( .A(n1608), .B(n1607), .Z(n1609) );
  XOR U1765 ( .A(n1610), .B(n1609), .Z(n1613) );
  NAND U1766 ( .A(b[0]), .B(a[57]), .Z(n1614) );
  XOR U1767 ( .A(n1613), .B(n1614), .Z(n1616) );
  OR U1768 ( .A(n1582), .B(n1581), .Z(n1586) );
  NANDN U1769 ( .A(n1584), .B(n1583), .Z(n1585) );
  NAND U1770 ( .A(n1586), .B(n1585), .Z(n1615) );
  XNOR U1771 ( .A(n1616), .B(n1615), .Z(n1601) );
  NANDN U1772 ( .A(n1588), .B(n1587), .Z(n1592) );
  OR U1773 ( .A(n1590), .B(n1589), .Z(n1591) );
  NAND U1774 ( .A(n1592), .B(n1591), .Z(n1602) );
  XNOR U1775 ( .A(n1601), .B(n1602), .Z(n1603) );
  XOR U1776 ( .A(n1604), .B(n1603), .Z(n1600) );
  NAND U1777 ( .A(n1593), .B(sreg[308]), .Z(n1597) );
  OR U1778 ( .A(n1595), .B(n1594), .Z(n1596) );
  NAND U1779 ( .A(n1597), .B(n1596), .Z(n1599) );
  XNOR U1780 ( .A(sreg[309]), .B(n1599), .Z(n1598) );
  XOR U1781 ( .A(n1600), .B(n1598), .Z(c[309]) );
  NANDN U1782 ( .A(n1602), .B(n1601), .Z(n1606) );
  NAND U1783 ( .A(n1604), .B(n1603), .Z(n1605) );
  NAND U1784 ( .A(n1606), .B(n1605), .Z(n1622) );
  AND U1785 ( .A(b[2]), .B(a[56]), .Z(n1628) );
  AND U1786 ( .A(a[57]), .B(b[1]), .Z(n1626) );
  AND U1787 ( .A(a[55]), .B(b[3]), .Z(n1625) );
  XOR U1788 ( .A(n1626), .B(n1625), .Z(n1627) );
  XOR U1789 ( .A(n1628), .B(n1627), .Z(n1631) );
  NAND U1790 ( .A(b[0]), .B(a[58]), .Z(n1632) );
  XOR U1791 ( .A(n1631), .B(n1632), .Z(n1634) );
  OR U1792 ( .A(n1608), .B(n1607), .Z(n1612) );
  NANDN U1793 ( .A(n1610), .B(n1609), .Z(n1611) );
  NAND U1794 ( .A(n1612), .B(n1611), .Z(n1633) );
  XNOR U1795 ( .A(n1634), .B(n1633), .Z(n1619) );
  NANDN U1796 ( .A(n1614), .B(n1613), .Z(n1618) );
  OR U1797 ( .A(n1616), .B(n1615), .Z(n1617) );
  NAND U1798 ( .A(n1618), .B(n1617), .Z(n1620) );
  XNOR U1799 ( .A(n1619), .B(n1620), .Z(n1621) );
  XNOR U1800 ( .A(n1622), .B(n1621), .Z(n1637) );
  XNOR U1801 ( .A(n1637), .B(sreg[310]), .Z(n1638) );
  XOR U1802 ( .A(n1639), .B(n1638), .Z(c[310]) );
  NANDN U1803 ( .A(n1620), .B(n1619), .Z(n1624) );
  NAND U1804 ( .A(n1622), .B(n1621), .Z(n1623) );
  NAND U1805 ( .A(n1624), .B(n1623), .Z(n1648) );
  AND U1806 ( .A(b[2]), .B(a[57]), .Z(n1654) );
  AND U1807 ( .A(a[58]), .B(b[1]), .Z(n1652) );
  AND U1808 ( .A(a[56]), .B(b[3]), .Z(n1651) );
  XOR U1809 ( .A(n1652), .B(n1651), .Z(n1653) );
  XOR U1810 ( .A(n1654), .B(n1653), .Z(n1657) );
  NAND U1811 ( .A(b[0]), .B(a[59]), .Z(n1658) );
  XOR U1812 ( .A(n1657), .B(n1658), .Z(n1660) );
  OR U1813 ( .A(n1626), .B(n1625), .Z(n1630) );
  NANDN U1814 ( .A(n1628), .B(n1627), .Z(n1629) );
  NAND U1815 ( .A(n1630), .B(n1629), .Z(n1659) );
  XNOR U1816 ( .A(n1660), .B(n1659), .Z(n1645) );
  NANDN U1817 ( .A(n1632), .B(n1631), .Z(n1636) );
  OR U1818 ( .A(n1634), .B(n1633), .Z(n1635) );
  NAND U1819 ( .A(n1636), .B(n1635), .Z(n1646) );
  XNOR U1820 ( .A(n1645), .B(n1646), .Z(n1647) );
  XNOR U1821 ( .A(n1648), .B(n1647), .Z(n1644) );
  NAND U1822 ( .A(n1637), .B(sreg[310]), .Z(n1641) );
  OR U1823 ( .A(n1639), .B(n1638), .Z(n1640) );
  AND U1824 ( .A(n1641), .B(n1640), .Z(n1643) );
  XNOR U1825 ( .A(n1643), .B(sreg[311]), .Z(n1642) );
  XOR U1826 ( .A(n1644), .B(n1642), .Z(c[311]) );
  NANDN U1827 ( .A(n1646), .B(n1645), .Z(n1650) );
  NAND U1828 ( .A(n1648), .B(n1647), .Z(n1649) );
  NAND U1829 ( .A(n1650), .B(n1649), .Z(n1666) );
  AND U1830 ( .A(b[2]), .B(a[58]), .Z(n1672) );
  AND U1831 ( .A(a[59]), .B(b[1]), .Z(n1670) );
  AND U1832 ( .A(a[57]), .B(b[3]), .Z(n1669) );
  XOR U1833 ( .A(n1670), .B(n1669), .Z(n1671) );
  XOR U1834 ( .A(n1672), .B(n1671), .Z(n1675) );
  NAND U1835 ( .A(b[0]), .B(a[60]), .Z(n1676) );
  XOR U1836 ( .A(n1675), .B(n1676), .Z(n1678) );
  OR U1837 ( .A(n1652), .B(n1651), .Z(n1656) );
  NANDN U1838 ( .A(n1654), .B(n1653), .Z(n1655) );
  NAND U1839 ( .A(n1656), .B(n1655), .Z(n1677) );
  XNOR U1840 ( .A(n1678), .B(n1677), .Z(n1663) );
  NANDN U1841 ( .A(n1658), .B(n1657), .Z(n1662) );
  OR U1842 ( .A(n1660), .B(n1659), .Z(n1661) );
  NAND U1843 ( .A(n1662), .B(n1661), .Z(n1664) );
  XNOR U1844 ( .A(n1663), .B(n1664), .Z(n1665) );
  XNOR U1845 ( .A(n1666), .B(n1665), .Z(n1681) );
  XOR U1846 ( .A(sreg[312]), .B(n1681), .Z(n1682) );
  XOR U1847 ( .A(n1683), .B(n1682), .Z(c[312]) );
  NANDN U1848 ( .A(n1664), .B(n1663), .Z(n1668) );
  NAND U1849 ( .A(n1666), .B(n1665), .Z(n1667) );
  NAND U1850 ( .A(n1668), .B(n1667), .Z(n1692) );
  AND U1851 ( .A(b[2]), .B(a[59]), .Z(n1698) );
  AND U1852 ( .A(a[60]), .B(b[1]), .Z(n1696) );
  AND U1853 ( .A(a[58]), .B(b[3]), .Z(n1695) );
  XOR U1854 ( .A(n1696), .B(n1695), .Z(n1697) );
  XOR U1855 ( .A(n1698), .B(n1697), .Z(n1701) );
  NAND U1856 ( .A(b[0]), .B(a[61]), .Z(n1702) );
  XOR U1857 ( .A(n1701), .B(n1702), .Z(n1704) );
  OR U1858 ( .A(n1670), .B(n1669), .Z(n1674) );
  NANDN U1859 ( .A(n1672), .B(n1671), .Z(n1673) );
  NAND U1860 ( .A(n1674), .B(n1673), .Z(n1703) );
  XNOR U1861 ( .A(n1704), .B(n1703), .Z(n1689) );
  NANDN U1862 ( .A(n1676), .B(n1675), .Z(n1680) );
  OR U1863 ( .A(n1678), .B(n1677), .Z(n1679) );
  NAND U1864 ( .A(n1680), .B(n1679), .Z(n1690) );
  XNOR U1865 ( .A(n1689), .B(n1690), .Z(n1691) );
  XOR U1866 ( .A(n1692), .B(n1691), .Z(n1688) );
  OR U1867 ( .A(n1681), .B(sreg[312]), .Z(n1685) );
  NANDN U1868 ( .A(n1683), .B(n1682), .Z(n1684) );
  AND U1869 ( .A(n1685), .B(n1684), .Z(n1687) );
  XNOR U1870 ( .A(sreg[313]), .B(n1687), .Z(n1686) );
  XOR U1871 ( .A(n1688), .B(n1686), .Z(c[313]) );
  NANDN U1872 ( .A(n1690), .B(n1689), .Z(n1694) );
  NAND U1873 ( .A(n1692), .B(n1691), .Z(n1693) );
  NAND U1874 ( .A(n1694), .B(n1693), .Z(n1710) );
  AND U1875 ( .A(b[2]), .B(a[60]), .Z(n1716) );
  AND U1876 ( .A(a[61]), .B(b[1]), .Z(n1714) );
  AND U1877 ( .A(a[59]), .B(b[3]), .Z(n1713) );
  XOR U1878 ( .A(n1714), .B(n1713), .Z(n1715) );
  XOR U1879 ( .A(n1716), .B(n1715), .Z(n1719) );
  NAND U1880 ( .A(b[0]), .B(a[62]), .Z(n1720) );
  XOR U1881 ( .A(n1719), .B(n1720), .Z(n1722) );
  OR U1882 ( .A(n1696), .B(n1695), .Z(n1700) );
  NANDN U1883 ( .A(n1698), .B(n1697), .Z(n1699) );
  NAND U1884 ( .A(n1700), .B(n1699), .Z(n1721) );
  XNOR U1885 ( .A(n1722), .B(n1721), .Z(n1707) );
  NANDN U1886 ( .A(n1702), .B(n1701), .Z(n1706) );
  OR U1887 ( .A(n1704), .B(n1703), .Z(n1705) );
  NAND U1888 ( .A(n1706), .B(n1705), .Z(n1708) );
  XNOR U1889 ( .A(n1707), .B(n1708), .Z(n1709) );
  XNOR U1890 ( .A(n1710), .B(n1709), .Z(n1725) );
  XNOR U1891 ( .A(n1725), .B(sreg[314]), .Z(n1726) );
  XOR U1892 ( .A(n1727), .B(n1726), .Z(c[314]) );
  NANDN U1893 ( .A(n1708), .B(n1707), .Z(n1712) );
  NAND U1894 ( .A(n1710), .B(n1709), .Z(n1711) );
  NAND U1895 ( .A(n1712), .B(n1711), .Z(n1733) );
  AND U1896 ( .A(b[2]), .B(a[61]), .Z(n1739) );
  AND U1897 ( .A(a[62]), .B(b[1]), .Z(n1737) );
  AND U1898 ( .A(a[60]), .B(b[3]), .Z(n1736) );
  XOR U1899 ( .A(n1737), .B(n1736), .Z(n1738) );
  XOR U1900 ( .A(n1739), .B(n1738), .Z(n1742) );
  NAND U1901 ( .A(b[0]), .B(a[63]), .Z(n1743) );
  XOR U1902 ( .A(n1742), .B(n1743), .Z(n1745) );
  OR U1903 ( .A(n1714), .B(n1713), .Z(n1718) );
  NANDN U1904 ( .A(n1716), .B(n1715), .Z(n1717) );
  NAND U1905 ( .A(n1718), .B(n1717), .Z(n1744) );
  XNOR U1906 ( .A(n1745), .B(n1744), .Z(n1730) );
  NANDN U1907 ( .A(n1720), .B(n1719), .Z(n1724) );
  OR U1908 ( .A(n1722), .B(n1721), .Z(n1723) );
  NAND U1909 ( .A(n1724), .B(n1723), .Z(n1731) );
  XNOR U1910 ( .A(n1730), .B(n1731), .Z(n1732) );
  XNOR U1911 ( .A(n1733), .B(n1732), .Z(n1748) );
  XOR U1912 ( .A(sreg[315]), .B(n1748), .Z(n1749) );
  NAND U1913 ( .A(n1725), .B(sreg[314]), .Z(n1729) );
  OR U1914 ( .A(n1727), .B(n1726), .Z(n1728) );
  NAND U1915 ( .A(n1729), .B(n1728), .Z(n1750) );
  XOR U1916 ( .A(n1749), .B(n1750), .Z(c[315]) );
  NANDN U1917 ( .A(n1731), .B(n1730), .Z(n1735) );
  NAND U1918 ( .A(n1733), .B(n1732), .Z(n1734) );
  NAND U1919 ( .A(n1735), .B(n1734), .Z(n1771) );
  AND U1920 ( .A(b[2]), .B(a[62]), .Z(n1765) );
  AND U1921 ( .A(a[63]), .B(b[1]), .Z(n1763) );
  AND U1922 ( .A(a[61]), .B(b[3]), .Z(n1762) );
  XOR U1923 ( .A(n1763), .B(n1762), .Z(n1764) );
  XOR U1924 ( .A(n1765), .B(n1764), .Z(n1756) );
  NAND U1925 ( .A(b[0]), .B(a[64]), .Z(n1757) );
  XOR U1926 ( .A(n1756), .B(n1757), .Z(n1759) );
  OR U1927 ( .A(n1737), .B(n1736), .Z(n1741) );
  NANDN U1928 ( .A(n1739), .B(n1738), .Z(n1740) );
  NAND U1929 ( .A(n1741), .B(n1740), .Z(n1758) );
  XNOR U1930 ( .A(n1759), .B(n1758), .Z(n1768) );
  NANDN U1931 ( .A(n1743), .B(n1742), .Z(n1747) );
  OR U1932 ( .A(n1745), .B(n1744), .Z(n1746) );
  NAND U1933 ( .A(n1747), .B(n1746), .Z(n1769) );
  XNOR U1934 ( .A(n1768), .B(n1769), .Z(n1770) );
  XOR U1935 ( .A(n1771), .B(n1770), .Z(n1755) );
  OR U1936 ( .A(n1748), .B(sreg[315]), .Z(n1752) );
  NANDN U1937 ( .A(n1750), .B(n1749), .Z(n1751) );
  AND U1938 ( .A(n1752), .B(n1751), .Z(n1754) );
  XNOR U1939 ( .A(sreg[316]), .B(n1754), .Z(n1753) );
  XOR U1940 ( .A(n1755), .B(n1753), .Z(c[316]) );
  NANDN U1941 ( .A(n1757), .B(n1756), .Z(n1761) );
  OR U1942 ( .A(n1759), .B(n1758), .Z(n1760) );
  NAND U1943 ( .A(n1761), .B(n1760), .Z(n1774) );
  AND U1944 ( .A(b[2]), .B(a[63]), .Z(n1783) );
  AND U1945 ( .A(a[64]), .B(b[1]), .Z(n1781) );
  AND U1946 ( .A(a[62]), .B(b[3]), .Z(n1780) );
  XOR U1947 ( .A(n1781), .B(n1780), .Z(n1782) );
  XOR U1948 ( .A(n1783), .B(n1782), .Z(n1786) );
  NAND U1949 ( .A(b[0]), .B(a[65]), .Z(n1787) );
  XNOR U1950 ( .A(n1786), .B(n1787), .Z(n1788) );
  OR U1951 ( .A(n1763), .B(n1762), .Z(n1767) );
  NANDN U1952 ( .A(n1765), .B(n1764), .Z(n1766) );
  AND U1953 ( .A(n1767), .B(n1766), .Z(n1789) );
  XNOR U1954 ( .A(n1788), .B(n1789), .Z(n1775) );
  XNOR U1955 ( .A(n1774), .B(n1775), .Z(n1776) );
  NANDN U1956 ( .A(n1769), .B(n1768), .Z(n1773) );
  NAND U1957 ( .A(n1771), .B(n1770), .Z(n1772) );
  AND U1958 ( .A(n1773), .B(n1772), .Z(n1777) );
  XOR U1959 ( .A(n1776), .B(n1777), .Z(n1792) );
  XNOR U1960 ( .A(sreg[317]), .B(n1792), .Z(n1793) );
  XOR U1961 ( .A(n1794), .B(n1793), .Z(c[317]) );
  NANDN U1962 ( .A(n1775), .B(n1774), .Z(n1779) );
  NAND U1963 ( .A(n1777), .B(n1776), .Z(n1778) );
  NAND U1964 ( .A(n1779), .B(n1778), .Z(n1803) );
  AND U1965 ( .A(b[2]), .B(a[64]), .Z(n1809) );
  AND U1966 ( .A(a[65]), .B(b[1]), .Z(n1807) );
  AND U1967 ( .A(a[63]), .B(b[3]), .Z(n1806) );
  XOR U1968 ( .A(n1807), .B(n1806), .Z(n1808) );
  XOR U1969 ( .A(n1809), .B(n1808), .Z(n1812) );
  NAND U1970 ( .A(b[0]), .B(a[66]), .Z(n1813) );
  XOR U1971 ( .A(n1812), .B(n1813), .Z(n1815) );
  OR U1972 ( .A(n1781), .B(n1780), .Z(n1785) );
  NANDN U1973 ( .A(n1783), .B(n1782), .Z(n1784) );
  NAND U1974 ( .A(n1785), .B(n1784), .Z(n1814) );
  XNOR U1975 ( .A(n1815), .B(n1814), .Z(n1800) );
  NANDN U1976 ( .A(n1787), .B(n1786), .Z(n1791) );
  NAND U1977 ( .A(n1789), .B(n1788), .Z(n1790) );
  NAND U1978 ( .A(n1791), .B(n1790), .Z(n1801) );
  XNOR U1979 ( .A(n1800), .B(n1801), .Z(n1802) );
  XOR U1980 ( .A(n1803), .B(n1802), .Z(n1799) );
  NAND U1981 ( .A(sreg[317]), .B(n1792), .Z(n1796) );
  OR U1982 ( .A(n1794), .B(n1793), .Z(n1795) );
  NAND U1983 ( .A(n1796), .B(n1795), .Z(n1798) );
  XNOR U1984 ( .A(sreg[318]), .B(n1798), .Z(n1797) );
  XNOR U1985 ( .A(n1799), .B(n1797), .Z(c[318]) );
  NANDN U1986 ( .A(n1801), .B(n1800), .Z(n1805) );
  NANDN U1987 ( .A(n1803), .B(n1802), .Z(n1804) );
  NAND U1988 ( .A(n1805), .B(n1804), .Z(n1821) );
  AND U1989 ( .A(b[2]), .B(a[65]), .Z(n1827) );
  AND U1990 ( .A(a[66]), .B(b[1]), .Z(n1825) );
  AND U1991 ( .A(a[64]), .B(b[3]), .Z(n1824) );
  XOR U1992 ( .A(n1825), .B(n1824), .Z(n1826) );
  XOR U1993 ( .A(n1827), .B(n1826), .Z(n1830) );
  NAND U1994 ( .A(b[0]), .B(a[67]), .Z(n1831) );
  XOR U1995 ( .A(n1830), .B(n1831), .Z(n1833) );
  OR U1996 ( .A(n1807), .B(n1806), .Z(n1811) );
  NANDN U1997 ( .A(n1809), .B(n1808), .Z(n1810) );
  NAND U1998 ( .A(n1811), .B(n1810), .Z(n1832) );
  XNOR U1999 ( .A(n1833), .B(n1832), .Z(n1818) );
  NANDN U2000 ( .A(n1813), .B(n1812), .Z(n1817) );
  OR U2001 ( .A(n1815), .B(n1814), .Z(n1816) );
  NAND U2002 ( .A(n1817), .B(n1816), .Z(n1819) );
  XNOR U2003 ( .A(n1818), .B(n1819), .Z(n1820) );
  XNOR U2004 ( .A(n1821), .B(n1820), .Z(n1836) );
  XNOR U2005 ( .A(n1836), .B(sreg[319]), .Z(n1837) );
  XOR U2006 ( .A(n1838), .B(n1837), .Z(c[319]) );
  NANDN U2007 ( .A(n1819), .B(n1818), .Z(n1823) );
  NAND U2008 ( .A(n1821), .B(n1820), .Z(n1822) );
  NAND U2009 ( .A(n1823), .B(n1822), .Z(n1844) );
  AND U2010 ( .A(b[2]), .B(a[66]), .Z(n1856) );
  AND U2011 ( .A(a[67]), .B(b[1]), .Z(n1854) );
  AND U2012 ( .A(a[65]), .B(b[3]), .Z(n1853) );
  XOR U2013 ( .A(n1854), .B(n1853), .Z(n1855) );
  XOR U2014 ( .A(n1856), .B(n1855), .Z(n1847) );
  NAND U2015 ( .A(b[0]), .B(a[68]), .Z(n1848) );
  XOR U2016 ( .A(n1847), .B(n1848), .Z(n1850) );
  OR U2017 ( .A(n1825), .B(n1824), .Z(n1829) );
  NANDN U2018 ( .A(n1827), .B(n1826), .Z(n1828) );
  NAND U2019 ( .A(n1829), .B(n1828), .Z(n1849) );
  XNOR U2020 ( .A(n1850), .B(n1849), .Z(n1841) );
  NANDN U2021 ( .A(n1831), .B(n1830), .Z(n1835) );
  OR U2022 ( .A(n1833), .B(n1832), .Z(n1834) );
  NAND U2023 ( .A(n1835), .B(n1834), .Z(n1842) );
  XNOR U2024 ( .A(n1841), .B(n1842), .Z(n1843) );
  XNOR U2025 ( .A(n1844), .B(n1843), .Z(n1859) );
  XOR U2026 ( .A(sreg[320]), .B(n1859), .Z(n1860) );
  NAND U2027 ( .A(n1836), .B(sreg[319]), .Z(n1840) );
  OR U2028 ( .A(n1838), .B(n1837), .Z(n1839) );
  NAND U2029 ( .A(n1840), .B(n1839), .Z(n1861) );
  XOR U2030 ( .A(n1860), .B(n1861), .Z(c[320]) );
  NANDN U2031 ( .A(n1842), .B(n1841), .Z(n1846) );
  NAND U2032 ( .A(n1844), .B(n1843), .Z(n1845) );
  NAND U2033 ( .A(n1846), .B(n1845), .Z(n1880) );
  NANDN U2034 ( .A(n1848), .B(n1847), .Z(n1852) );
  OR U2035 ( .A(n1850), .B(n1849), .Z(n1851) );
  NAND U2036 ( .A(n1852), .B(n1851), .Z(n1877) );
  AND U2037 ( .A(b[2]), .B(a[67]), .Z(n1868) );
  AND U2038 ( .A(a[68]), .B(b[1]), .Z(n1866) );
  AND U2039 ( .A(a[66]), .B(b[3]), .Z(n1865) );
  XOR U2040 ( .A(n1866), .B(n1865), .Z(n1867) );
  XOR U2041 ( .A(n1868), .B(n1867), .Z(n1871) );
  NAND U2042 ( .A(b[0]), .B(a[69]), .Z(n1872) );
  XNOR U2043 ( .A(n1871), .B(n1872), .Z(n1873) );
  OR U2044 ( .A(n1854), .B(n1853), .Z(n1858) );
  NANDN U2045 ( .A(n1856), .B(n1855), .Z(n1857) );
  AND U2046 ( .A(n1858), .B(n1857), .Z(n1874) );
  XNOR U2047 ( .A(n1873), .B(n1874), .Z(n1878) );
  XNOR U2048 ( .A(n1877), .B(n1878), .Z(n1879) );
  XNOR U2049 ( .A(n1880), .B(n1879), .Z(n1884) );
  OR U2050 ( .A(n1859), .B(sreg[320]), .Z(n1863) );
  NANDN U2051 ( .A(n1861), .B(n1860), .Z(n1862) );
  AND U2052 ( .A(n1863), .B(n1862), .Z(n1883) );
  XNOR U2053 ( .A(sreg[321]), .B(n1883), .Z(n1864) );
  XNOR U2054 ( .A(n1884), .B(n1864), .Z(c[321]) );
  AND U2055 ( .A(b[2]), .B(a[68]), .Z(n1897) );
  AND U2056 ( .A(a[69]), .B(b[1]), .Z(n1895) );
  AND U2057 ( .A(a[67]), .B(b[3]), .Z(n1894) );
  XOR U2058 ( .A(n1895), .B(n1894), .Z(n1896) );
  XOR U2059 ( .A(n1897), .B(n1896), .Z(n1900) );
  NAND U2060 ( .A(b[0]), .B(a[70]), .Z(n1901) );
  XOR U2061 ( .A(n1900), .B(n1901), .Z(n1903) );
  OR U2062 ( .A(n1866), .B(n1865), .Z(n1870) );
  NANDN U2063 ( .A(n1868), .B(n1867), .Z(n1869) );
  NAND U2064 ( .A(n1870), .B(n1869), .Z(n1902) );
  XNOR U2065 ( .A(n1903), .B(n1902), .Z(n1888) );
  NANDN U2066 ( .A(n1872), .B(n1871), .Z(n1876) );
  NAND U2067 ( .A(n1874), .B(n1873), .Z(n1875) );
  NAND U2068 ( .A(n1876), .B(n1875), .Z(n1889) );
  XNOR U2069 ( .A(n1888), .B(n1889), .Z(n1890) );
  NANDN U2070 ( .A(n1878), .B(n1877), .Z(n1882) );
  NANDN U2071 ( .A(n1880), .B(n1879), .Z(n1881) );
  NAND U2072 ( .A(n1882), .B(n1881), .Z(n1891) );
  XOR U2073 ( .A(n1890), .B(n1891), .Z(n1887) );
  XNOR U2074 ( .A(sreg[322]), .B(n1886), .Z(n1885) );
  XNOR U2075 ( .A(n1887), .B(n1885), .Z(c[322]) );
  NANDN U2076 ( .A(n1889), .B(n1888), .Z(n1893) );
  NANDN U2077 ( .A(n1891), .B(n1890), .Z(n1892) );
  NAND U2078 ( .A(n1893), .B(n1892), .Z(n1921) );
  AND U2079 ( .A(b[2]), .B(a[69]), .Z(n1915) );
  AND U2080 ( .A(a[70]), .B(b[1]), .Z(n1913) );
  AND U2081 ( .A(a[68]), .B(b[3]), .Z(n1912) );
  XOR U2082 ( .A(n1913), .B(n1912), .Z(n1914) );
  XOR U2083 ( .A(n1915), .B(n1914), .Z(n1906) );
  NAND U2084 ( .A(b[0]), .B(a[71]), .Z(n1907) );
  XOR U2085 ( .A(n1906), .B(n1907), .Z(n1909) );
  OR U2086 ( .A(n1895), .B(n1894), .Z(n1899) );
  NANDN U2087 ( .A(n1897), .B(n1896), .Z(n1898) );
  NAND U2088 ( .A(n1899), .B(n1898), .Z(n1908) );
  XNOR U2089 ( .A(n1909), .B(n1908), .Z(n1918) );
  NANDN U2090 ( .A(n1901), .B(n1900), .Z(n1905) );
  OR U2091 ( .A(n1903), .B(n1902), .Z(n1904) );
  NAND U2092 ( .A(n1905), .B(n1904), .Z(n1919) );
  XNOR U2093 ( .A(n1918), .B(n1919), .Z(n1920) );
  XNOR U2094 ( .A(n1921), .B(n1920), .Z(n1924) );
  XNOR U2095 ( .A(n1924), .B(sreg[323]), .Z(n1925) );
  XOR U2096 ( .A(n1926), .B(n1925), .Z(c[323]) );
  NANDN U2097 ( .A(n1907), .B(n1906), .Z(n1911) );
  OR U2098 ( .A(n1909), .B(n1908), .Z(n1910) );
  NAND U2099 ( .A(n1911), .B(n1910), .Z(n1932) );
  AND U2100 ( .A(b[2]), .B(a[70]), .Z(n1941) );
  AND U2101 ( .A(a[71]), .B(b[1]), .Z(n1939) );
  AND U2102 ( .A(a[69]), .B(b[3]), .Z(n1938) );
  XOR U2103 ( .A(n1939), .B(n1938), .Z(n1940) );
  XOR U2104 ( .A(n1941), .B(n1940), .Z(n1944) );
  NAND U2105 ( .A(b[0]), .B(a[72]), .Z(n1945) );
  XNOR U2106 ( .A(n1944), .B(n1945), .Z(n1946) );
  OR U2107 ( .A(n1913), .B(n1912), .Z(n1917) );
  NANDN U2108 ( .A(n1915), .B(n1914), .Z(n1916) );
  AND U2109 ( .A(n1917), .B(n1916), .Z(n1947) );
  XNOR U2110 ( .A(n1946), .B(n1947), .Z(n1933) );
  XNOR U2111 ( .A(n1932), .B(n1933), .Z(n1934) );
  NANDN U2112 ( .A(n1919), .B(n1918), .Z(n1923) );
  NAND U2113 ( .A(n1921), .B(n1920), .Z(n1922) );
  NAND U2114 ( .A(n1923), .B(n1922), .Z(n1935) );
  XOR U2115 ( .A(n1934), .B(n1935), .Z(n1931) );
  NAND U2116 ( .A(n1924), .B(sreg[323]), .Z(n1928) );
  OR U2117 ( .A(n1926), .B(n1925), .Z(n1927) );
  AND U2118 ( .A(n1928), .B(n1927), .Z(n1930) );
  XNOR U2119 ( .A(n1930), .B(sreg[324]), .Z(n1929) );
  XNOR U2120 ( .A(n1931), .B(n1929), .Z(c[324]) );
  NANDN U2121 ( .A(n1933), .B(n1932), .Z(n1937) );
  NANDN U2122 ( .A(n1935), .B(n1934), .Z(n1936) );
  NAND U2123 ( .A(n1937), .B(n1936), .Z(n1953) );
  AND U2124 ( .A(b[2]), .B(a[71]), .Z(n1959) );
  AND U2125 ( .A(a[72]), .B(b[1]), .Z(n1957) );
  AND U2126 ( .A(a[70]), .B(b[3]), .Z(n1956) );
  XOR U2127 ( .A(n1957), .B(n1956), .Z(n1958) );
  XOR U2128 ( .A(n1959), .B(n1958), .Z(n1962) );
  NAND U2129 ( .A(b[0]), .B(a[73]), .Z(n1963) );
  XOR U2130 ( .A(n1962), .B(n1963), .Z(n1965) );
  OR U2131 ( .A(n1939), .B(n1938), .Z(n1943) );
  NANDN U2132 ( .A(n1941), .B(n1940), .Z(n1942) );
  NAND U2133 ( .A(n1943), .B(n1942), .Z(n1964) );
  XNOR U2134 ( .A(n1965), .B(n1964), .Z(n1950) );
  NANDN U2135 ( .A(n1945), .B(n1944), .Z(n1949) );
  NAND U2136 ( .A(n1947), .B(n1946), .Z(n1948) );
  NAND U2137 ( .A(n1949), .B(n1948), .Z(n1951) );
  XNOR U2138 ( .A(n1950), .B(n1951), .Z(n1952) );
  XOR U2139 ( .A(n1953), .B(n1952), .Z(n1968) );
  XNOR U2140 ( .A(n1968), .B(sreg[325]), .Z(n1970) );
  XNOR U2141 ( .A(n1969), .B(n1970), .Z(c[325]) );
  NANDN U2142 ( .A(n1951), .B(n1950), .Z(n1955) );
  NANDN U2143 ( .A(n1953), .B(n1952), .Z(n1954) );
  NAND U2144 ( .A(n1955), .B(n1954), .Z(n1988) );
  AND U2145 ( .A(b[2]), .B(a[72]), .Z(n1982) );
  AND U2146 ( .A(a[73]), .B(b[1]), .Z(n1980) );
  AND U2147 ( .A(a[71]), .B(b[3]), .Z(n1979) );
  XOR U2148 ( .A(n1980), .B(n1979), .Z(n1981) );
  XOR U2149 ( .A(n1982), .B(n1981), .Z(n1973) );
  NAND U2150 ( .A(b[0]), .B(a[74]), .Z(n1974) );
  XOR U2151 ( .A(n1973), .B(n1974), .Z(n1976) );
  OR U2152 ( .A(n1957), .B(n1956), .Z(n1961) );
  NANDN U2153 ( .A(n1959), .B(n1958), .Z(n1960) );
  NAND U2154 ( .A(n1961), .B(n1960), .Z(n1975) );
  XNOR U2155 ( .A(n1976), .B(n1975), .Z(n1985) );
  NANDN U2156 ( .A(n1963), .B(n1962), .Z(n1967) );
  OR U2157 ( .A(n1965), .B(n1964), .Z(n1966) );
  NAND U2158 ( .A(n1967), .B(n1966), .Z(n1986) );
  XNOR U2159 ( .A(n1985), .B(n1986), .Z(n1987) );
  XNOR U2160 ( .A(n1988), .B(n1987), .Z(n1991) );
  XOR U2161 ( .A(sreg[326]), .B(n1991), .Z(n1992) );
  NAND U2162 ( .A(n1968), .B(sreg[325]), .Z(n1972) );
  NANDN U2163 ( .A(n1970), .B(n1969), .Z(n1971) );
  NAND U2164 ( .A(n1972), .B(n1971), .Z(n1993) );
  XOR U2165 ( .A(n1992), .B(n1993), .Z(c[326]) );
  NANDN U2166 ( .A(n1974), .B(n1973), .Z(n1978) );
  OR U2167 ( .A(n1976), .B(n1975), .Z(n1977) );
  NAND U2168 ( .A(n1978), .B(n1977), .Z(n1997) );
  AND U2169 ( .A(b[2]), .B(a[73]), .Z(n2006) );
  AND U2170 ( .A(a[74]), .B(b[1]), .Z(n2004) );
  AND U2171 ( .A(a[72]), .B(b[3]), .Z(n2003) );
  XOR U2172 ( .A(n2004), .B(n2003), .Z(n2005) );
  XOR U2173 ( .A(n2006), .B(n2005), .Z(n2009) );
  NAND U2174 ( .A(b[0]), .B(a[75]), .Z(n2010) );
  XNOR U2175 ( .A(n2009), .B(n2010), .Z(n2011) );
  OR U2176 ( .A(n1980), .B(n1979), .Z(n1984) );
  NANDN U2177 ( .A(n1982), .B(n1981), .Z(n1983) );
  AND U2178 ( .A(n1984), .B(n1983), .Z(n2012) );
  XNOR U2179 ( .A(n2011), .B(n2012), .Z(n1998) );
  XNOR U2180 ( .A(n1997), .B(n1998), .Z(n1999) );
  NANDN U2181 ( .A(n1986), .B(n1985), .Z(n1990) );
  NAND U2182 ( .A(n1988), .B(n1987), .Z(n1989) );
  AND U2183 ( .A(n1990), .B(n1989), .Z(n2000) );
  XNOR U2184 ( .A(n1999), .B(n2000), .Z(n2016) );
  OR U2185 ( .A(n1991), .B(sreg[326]), .Z(n1995) );
  NANDN U2186 ( .A(n1993), .B(n1992), .Z(n1994) );
  AND U2187 ( .A(n1995), .B(n1994), .Z(n2015) );
  XNOR U2188 ( .A(sreg[327]), .B(n2015), .Z(n1996) );
  XOR U2189 ( .A(n2016), .B(n1996), .Z(c[327]) );
  NANDN U2190 ( .A(n1998), .B(n1997), .Z(n2002) );
  NAND U2191 ( .A(n2000), .B(n1999), .Z(n2001) );
  NAND U2192 ( .A(n2002), .B(n2001), .Z(n2023) );
  AND U2193 ( .A(b[2]), .B(a[74]), .Z(n2029) );
  AND U2194 ( .A(a[75]), .B(b[1]), .Z(n2027) );
  AND U2195 ( .A(a[73]), .B(b[3]), .Z(n2026) );
  XOR U2196 ( .A(n2027), .B(n2026), .Z(n2028) );
  XOR U2197 ( .A(n2029), .B(n2028), .Z(n2032) );
  NAND U2198 ( .A(b[0]), .B(a[76]), .Z(n2033) );
  XOR U2199 ( .A(n2032), .B(n2033), .Z(n2035) );
  OR U2200 ( .A(n2004), .B(n2003), .Z(n2008) );
  NANDN U2201 ( .A(n2006), .B(n2005), .Z(n2007) );
  NAND U2202 ( .A(n2008), .B(n2007), .Z(n2034) );
  XNOR U2203 ( .A(n2035), .B(n2034), .Z(n2020) );
  NANDN U2204 ( .A(n2010), .B(n2009), .Z(n2014) );
  NAND U2205 ( .A(n2012), .B(n2011), .Z(n2013) );
  NAND U2206 ( .A(n2014), .B(n2013), .Z(n2021) );
  XNOR U2207 ( .A(n2020), .B(n2021), .Z(n2022) );
  XNOR U2208 ( .A(n2023), .B(n2022), .Z(n2019) );
  XOR U2209 ( .A(n2018), .B(sreg[328]), .Z(n2017) );
  XNOR U2210 ( .A(n2019), .B(n2017), .Z(c[328]) );
  NANDN U2211 ( .A(n2021), .B(n2020), .Z(n2025) );
  NANDN U2212 ( .A(n2023), .B(n2022), .Z(n2024) );
  NAND U2213 ( .A(n2025), .B(n2024), .Z(n2053) );
  AND U2214 ( .A(b[2]), .B(a[75]), .Z(n2047) );
  AND U2215 ( .A(a[76]), .B(b[1]), .Z(n2045) );
  AND U2216 ( .A(a[74]), .B(b[3]), .Z(n2044) );
  XOR U2217 ( .A(n2045), .B(n2044), .Z(n2046) );
  XOR U2218 ( .A(n2047), .B(n2046), .Z(n2038) );
  NAND U2219 ( .A(b[0]), .B(a[77]), .Z(n2039) );
  XOR U2220 ( .A(n2038), .B(n2039), .Z(n2041) );
  OR U2221 ( .A(n2027), .B(n2026), .Z(n2031) );
  NANDN U2222 ( .A(n2029), .B(n2028), .Z(n2030) );
  NAND U2223 ( .A(n2031), .B(n2030), .Z(n2040) );
  XNOR U2224 ( .A(n2041), .B(n2040), .Z(n2050) );
  NANDN U2225 ( .A(n2033), .B(n2032), .Z(n2037) );
  OR U2226 ( .A(n2035), .B(n2034), .Z(n2036) );
  NAND U2227 ( .A(n2037), .B(n2036), .Z(n2051) );
  XNOR U2228 ( .A(n2050), .B(n2051), .Z(n2052) );
  XNOR U2229 ( .A(n2053), .B(n2052), .Z(n2056) );
  XNOR U2230 ( .A(n2056), .B(sreg[329]), .Z(n2058) );
  XNOR U2231 ( .A(n2057), .B(n2058), .Z(c[329]) );
  NANDN U2232 ( .A(n2039), .B(n2038), .Z(n2043) );
  OR U2233 ( .A(n2041), .B(n2040), .Z(n2042) );
  NAND U2234 ( .A(n2043), .B(n2042), .Z(n2061) );
  AND U2235 ( .A(b[2]), .B(a[76]), .Z(n2070) );
  AND U2236 ( .A(a[77]), .B(b[1]), .Z(n2068) );
  AND U2237 ( .A(a[75]), .B(b[3]), .Z(n2067) );
  XOR U2238 ( .A(n2068), .B(n2067), .Z(n2069) );
  XOR U2239 ( .A(n2070), .B(n2069), .Z(n2073) );
  NAND U2240 ( .A(b[0]), .B(a[78]), .Z(n2074) );
  XNOR U2241 ( .A(n2073), .B(n2074), .Z(n2075) );
  OR U2242 ( .A(n2045), .B(n2044), .Z(n2049) );
  NANDN U2243 ( .A(n2047), .B(n2046), .Z(n2048) );
  AND U2244 ( .A(n2049), .B(n2048), .Z(n2076) );
  XNOR U2245 ( .A(n2075), .B(n2076), .Z(n2062) );
  XNOR U2246 ( .A(n2061), .B(n2062), .Z(n2063) );
  NANDN U2247 ( .A(n2051), .B(n2050), .Z(n2055) );
  NAND U2248 ( .A(n2053), .B(n2052), .Z(n2054) );
  AND U2249 ( .A(n2055), .B(n2054), .Z(n2064) );
  XOR U2250 ( .A(n2063), .B(n2064), .Z(n2079) );
  XNOR U2251 ( .A(sreg[330]), .B(n2079), .Z(n2081) );
  NAND U2252 ( .A(n2056), .B(sreg[329]), .Z(n2060) );
  NANDN U2253 ( .A(n2058), .B(n2057), .Z(n2059) );
  AND U2254 ( .A(n2060), .B(n2059), .Z(n2080) );
  XOR U2255 ( .A(n2081), .B(n2080), .Z(c[330]) );
  NANDN U2256 ( .A(n2062), .B(n2061), .Z(n2066) );
  NAND U2257 ( .A(n2064), .B(n2063), .Z(n2065) );
  NAND U2258 ( .A(n2066), .B(n2065), .Z(n2090) );
  AND U2259 ( .A(b[2]), .B(a[77]), .Z(n2096) );
  AND U2260 ( .A(a[78]), .B(b[1]), .Z(n2094) );
  AND U2261 ( .A(a[76]), .B(b[3]), .Z(n2093) );
  XOR U2262 ( .A(n2094), .B(n2093), .Z(n2095) );
  XOR U2263 ( .A(n2096), .B(n2095), .Z(n2099) );
  NAND U2264 ( .A(b[0]), .B(a[79]), .Z(n2100) );
  XOR U2265 ( .A(n2099), .B(n2100), .Z(n2102) );
  OR U2266 ( .A(n2068), .B(n2067), .Z(n2072) );
  NANDN U2267 ( .A(n2070), .B(n2069), .Z(n2071) );
  NAND U2268 ( .A(n2072), .B(n2071), .Z(n2101) );
  XNOR U2269 ( .A(n2102), .B(n2101), .Z(n2087) );
  NANDN U2270 ( .A(n2074), .B(n2073), .Z(n2078) );
  NAND U2271 ( .A(n2076), .B(n2075), .Z(n2077) );
  NAND U2272 ( .A(n2078), .B(n2077), .Z(n2088) );
  XNOR U2273 ( .A(n2087), .B(n2088), .Z(n2089) );
  XNOR U2274 ( .A(n2090), .B(n2089), .Z(n2086) );
  NAND U2275 ( .A(sreg[330]), .B(n2079), .Z(n2083) );
  OR U2276 ( .A(n2081), .B(n2080), .Z(n2082) );
  AND U2277 ( .A(n2083), .B(n2082), .Z(n2085) );
  XNOR U2278 ( .A(n2085), .B(sreg[331]), .Z(n2084) );
  XNOR U2279 ( .A(n2086), .B(n2084), .Z(c[331]) );
  NANDN U2280 ( .A(n2088), .B(n2087), .Z(n2092) );
  NANDN U2281 ( .A(n2090), .B(n2089), .Z(n2091) );
  NAND U2282 ( .A(n2092), .B(n2091), .Z(n2125) );
  AND U2283 ( .A(b[2]), .B(a[78]), .Z(n2119) );
  AND U2284 ( .A(a[79]), .B(b[1]), .Z(n2117) );
  AND U2285 ( .A(a[77]), .B(b[3]), .Z(n2116) );
  XOR U2286 ( .A(n2117), .B(n2116), .Z(n2118) );
  XOR U2287 ( .A(n2119), .B(n2118), .Z(n2110) );
  NAND U2288 ( .A(b[0]), .B(a[80]), .Z(n2111) );
  XOR U2289 ( .A(n2110), .B(n2111), .Z(n2113) );
  OR U2290 ( .A(n2094), .B(n2093), .Z(n2098) );
  NANDN U2291 ( .A(n2096), .B(n2095), .Z(n2097) );
  NAND U2292 ( .A(n2098), .B(n2097), .Z(n2112) );
  XNOR U2293 ( .A(n2113), .B(n2112), .Z(n2122) );
  NANDN U2294 ( .A(n2100), .B(n2099), .Z(n2104) );
  OR U2295 ( .A(n2102), .B(n2101), .Z(n2103) );
  NAND U2296 ( .A(n2104), .B(n2103), .Z(n2123) );
  XNOR U2297 ( .A(n2122), .B(n2123), .Z(n2124) );
  XNOR U2298 ( .A(n2125), .B(n2124), .Z(n2105) );
  XNOR U2299 ( .A(n2105), .B(sreg[332]), .Z(n2107) );
  XNOR U2300 ( .A(n2106), .B(n2107), .Z(c[332]) );
  NAND U2301 ( .A(n2105), .B(sreg[332]), .Z(n2109) );
  NANDN U2302 ( .A(n2107), .B(n2106), .Z(n2108) );
  AND U2303 ( .A(n2109), .B(n2108), .Z(n2130) );
  IV U2304 ( .A(n2130), .Z(n2129) );
  NANDN U2305 ( .A(n2111), .B(n2110), .Z(n2115) );
  OR U2306 ( .A(n2113), .B(n2112), .Z(n2114) );
  NAND U2307 ( .A(n2115), .B(n2114), .Z(n2135) );
  AND U2308 ( .A(b[2]), .B(a[79]), .Z(n2144) );
  AND U2309 ( .A(a[80]), .B(b[1]), .Z(n2142) );
  AND U2310 ( .A(a[78]), .B(b[3]), .Z(n2141) );
  XOR U2311 ( .A(n2142), .B(n2141), .Z(n2143) );
  XOR U2312 ( .A(n2144), .B(n2143), .Z(n2147) );
  NAND U2313 ( .A(b[0]), .B(a[81]), .Z(n2148) );
  XNOR U2314 ( .A(n2147), .B(n2148), .Z(n2149) );
  OR U2315 ( .A(n2117), .B(n2116), .Z(n2121) );
  NANDN U2316 ( .A(n2119), .B(n2118), .Z(n2120) );
  AND U2317 ( .A(n2121), .B(n2120), .Z(n2150) );
  XNOR U2318 ( .A(n2149), .B(n2150), .Z(n2136) );
  XNOR U2319 ( .A(n2135), .B(n2136), .Z(n2137) );
  NANDN U2320 ( .A(n2123), .B(n2122), .Z(n2127) );
  NAND U2321 ( .A(n2125), .B(n2124), .Z(n2126) );
  AND U2322 ( .A(n2127), .B(n2126), .Z(n2138) );
  XNOR U2323 ( .A(n2137), .B(n2138), .Z(n2132) );
  XOR U2324 ( .A(sreg[333]), .B(n2132), .Z(n2128) );
  XNOR U2325 ( .A(n2129), .B(n2128), .Z(c[333]) );
  NAND U2326 ( .A(n2129), .B(sreg[333]), .Z(n2134) );
  NANDN U2327 ( .A(sreg[333]), .B(n2130), .Z(n2131) );
  NANDN U2328 ( .A(n2132), .B(n2131), .Z(n2133) );
  NAND U2329 ( .A(n2134), .B(n2133), .Z(n2173) );
  NANDN U2330 ( .A(n2136), .B(n2135), .Z(n2140) );
  NAND U2331 ( .A(n2138), .B(n2137), .Z(n2139) );
  NAND U2332 ( .A(n2140), .B(n2139), .Z(n2156) );
  AND U2333 ( .A(b[2]), .B(a[80]), .Z(n2162) );
  AND U2334 ( .A(a[81]), .B(b[1]), .Z(n2160) );
  AND U2335 ( .A(a[79]), .B(b[3]), .Z(n2159) );
  XOR U2336 ( .A(n2160), .B(n2159), .Z(n2161) );
  XOR U2337 ( .A(n2162), .B(n2161), .Z(n2165) );
  NAND U2338 ( .A(b[0]), .B(a[82]), .Z(n2166) );
  XOR U2339 ( .A(n2165), .B(n2166), .Z(n2168) );
  OR U2340 ( .A(n2142), .B(n2141), .Z(n2146) );
  NANDN U2341 ( .A(n2144), .B(n2143), .Z(n2145) );
  NAND U2342 ( .A(n2146), .B(n2145), .Z(n2167) );
  XNOR U2343 ( .A(n2168), .B(n2167), .Z(n2153) );
  NANDN U2344 ( .A(n2148), .B(n2147), .Z(n2152) );
  NAND U2345 ( .A(n2150), .B(n2149), .Z(n2151) );
  NAND U2346 ( .A(n2152), .B(n2151), .Z(n2154) );
  XNOR U2347 ( .A(n2153), .B(n2154), .Z(n2155) );
  XNOR U2348 ( .A(n2156), .B(n2155), .Z(n2171) );
  XOR U2349 ( .A(sreg[334]), .B(n2171), .Z(n2172) );
  XNOR U2350 ( .A(n2173), .B(n2172), .Z(c[334]) );
  NANDN U2351 ( .A(n2154), .B(n2153), .Z(n2158) );
  NANDN U2352 ( .A(n2156), .B(n2155), .Z(n2157) );
  NAND U2353 ( .A(n2158), .B(n2157), .Z(n2182) );
  AND U2354 ( .A(b[2]), .B(a[81]), .Z(n2188) );
  AND U2355 ( .A(a[82]), .B(b[1]), .Z(n2186) );
  AND U2356 ( .A(a[80]), .B(b[3]), .Z(n2185) );
  XOR U2357 ( .A(n2186), .B(n2185), .Z(n2187) );
  XOR U2358 ( .A(n2188), .B(n2187), .Z(n2191) );
  NAND U2359 ( .A(b[0]), .B(a[83]), .Z(n2192) );
  XOR U2360 ( .A(n2191), .B(n2192), .Z(n2194) );
  OR U2361 ( .A(n2160), .B(n2159), .Z(n2164) );
  NANDN U2362 ( .A(n2162), .B(n2161), .Z(n2163) );
  NAND U2363 ( .A(n2164), .B(n2163), .Z(n2193) );
  XNOR U2364 ( .A(n2194), .B(n2193), .Z(n2179) );
  NANDN U2365 ( .A(n2166), .B(n2165), .Z(n2170) );
  OR U2366 ( .A(n2168), .B(n2167), .Z(n2169) );
  NAND U2367 ( .A(n2170), .B(n2169), .Z(n2180) );
  XNOR U2368 ( .A(n2179), .B(n2180), .Z(n2181) );
  XOR U2369 ( .A(n2182), .B(n2181), .Z(n2178) );
  NANDN U2370 ( .A(sreg[334]), .B(n2171), .Z(n2175) );
  OR U2371 ( .A(n2173), .B(n2172), .Z(n2174) );
  AND U2372 ( .A(n2175), .B(n2174), .Z(n2177) );
  XNOR U2373 ( .A(sreg[335]), .B(n2177), .Z(n2176) );
  XOR U2374 ( .A(n2178), .B(n2176), .Z(c[335]) );
  NANDN U2375 ( .A(n2180), .B(n2179), .Z(n2184) );
  NAND U2376 ( .A(n2182), .B(n2181), .Z(n2183) );
  AND U2377 ( .A(n2184), .B(n2183), .Z(n2200) );
  AND U2378 ( .A(b[2]), .B(a[82]), .Z(n2204) );
  AND U2379 ( .A(a[83]), .B(b[1]), .Z(n2202) );
  AND U2380 ( .A(a[81]), .B(b[3]), .Z(n2201) );
  XOR U2381 ( .A(n2202), .B(n2201), .Z(n2203) );
  XOR U2382 ( .A(n2204), .B(n2203), .Z(n2207) );
  NAND U2383 ( .A(b[0]), .B(a[84]), .Z(n2208) );
  XOR U2384 ( .A(n2207), .B(n2208), .Z(n2209) );
  OR U2385 ( .A(n2186), .B(n2185), .Z(n2190) );
  NANDN U2386 ( .A(n2188), .B(n2187), .Z(n2189) );
  AND U2387 ( .A(n2190), .B(n2189), .Z(n2210) );
  XOR U2388 ( .A(n2209), .B(n2210), .Z(n2198) );
  NANDN U2389 ( .A(n2192), .B(n2191), .Z(n2196) );
  OR U2390 ( .A(n2194), .B(n2193), .Z(n2195) );
  AND U2391 ( .A(n2196), .B(n2195), .Z(n2199) );
  XOR U2392 ( .A(n2198), .B(n2199), .Z(n2197) );
  XOR U2393 ( .A(n2200), .B(n2197), .Z(n2211) );
  XNOR U2394 ( .A(sreg[336]), .B(n2211), .Z(n2212) );
  XOR U2395 ( .A(n2213), .B(n2212), .Z(c[336]) );
  AND U2396 ( .A(b[2]), .B(a[83]), .Z(n2225) );
  AND U2397 ( .A(a[84]), .B(b[1]), .Z(n2223) );
  AND U2398 ( .A(a[82]), .B(b[3]), .Z(n2222) );
  XOR U2399 ( .A(n2223), .B(n2222), .Z(n2224) );
  XOR U2400 ( .A(n2225), .B(n2224), .Z(n2228) );
  NAND U2401 ( .A(b[0]), .B(a[85]), .Z(n2229) );
  XOR U2402 ( .A(n2228), .B(n2229), .Z(n2231) );
  OR U2403 ( .A(n2202), .B(n2201), .Z(n2206) );
  NANDN U2404 ( .A(n2204), .B(n2203), .Z(n2205) );
  NAND U2405 ( .A(n2206), .B(n2205), .Z(n2230) );
  XNOR U2406 ( .A(n2231), .B(n2230), .Z(n2216) );
  XNOR U2407 ( .A(n2216), .B(n2217), .Z(n2219) );
  XOR U2408 ( .A(n2218), .B(n2219), .Z(n2234) );
  XOR U2409 ( .A(n2234), .B(sreg[337]), .Z(n2236) );
  NAND U2410 ( .A(sreg[336]), .B(n2211), .Z(n2215) );
  OR U2411 ( .A(n2213), .B(n2212), .Z(n2214) );
  AND U2412 ( .A(n2215), .B(n2214), .Z(n2235) );
  XOR U2413 ( .A(n2236), .B(n2235), .Z(c[337]) );
  NANDN U2414 ( .A(n2217), .B(n2216), .Z(n2221) );
  NAND U2415 ( .A(n2219), .B(n2218), .Z(n2220) );
  NAND U2416 ( .A(n2221), .B(n2220), .Z(n2245) );
  AND U2417 ( .A(b[2]), .B(a[84]), .Z(n2251) );
  AND U2418 ( .A(a[85]), .B(b[1]), .Z(n2249) );
  AND U2419 ( .A(a[83]), .B(b[3]), .Z(n2248) );
  XOR U2420 ( .A(n2249), .B(n2248), .Z(n2250) );
  XOR U2421 ( .A(n2251), .B(n2250), .Z(n2254) );
  NAND U2422 ( .A(b[0]), .B(a[86]), .Z(n2255) );
  XOR U2423 ( .A(n2254), .B(n2255), .Z(n2257) );
  OR U2424 ( .A(n2223), .B(n2222), .Z(n2227) );
  NANDN U2425 ( .A(n2225), .B(n2224), .Z(n2226) );
  NAND U2426 ( .A(n2227), .B(n2226), .Z(n2256) );
  XNOR U2427 ( .A(n2257), .B(n2256), .Z(n2242) );
  NANDN U2428 ( .A(n2229), .B(n2228), .Z(n2233) );
  OR U2429 ( .A(n2231), .B(n2230), .Z(n2232) );
  NAND U2430 ( .A(n2233), .B(n2232), .Z(n2243) );
  XNOR U2431 ( .A(n2242), .B(n2243), .Z(n2244) );
  XOR U2432 ( .A(n2245), .B(n2244), .Z(n2241) );
  NANDN U2433 ( .A(n2234), .B(sreg[337]), .Z(n2238) );
  OR U2434 ( .A(n2236), .B(n2235), .Z(n2237) );
  NAND U2435 ( .A(n2238), .B(n2237), .Z(n2240) );
  XNOR U2436 ( .A(sreg[338]), .B(n2240), .Z(n2239) );
  XOR U2437 ( .A(n2241), .B(n2239), .Z(c[338]) );
  NANDN U2438 ( .A(n2243), .B(n2242), .Z(n2247) );
  NAND U2439 ( .A(n2245), .B(n2244), .Z(n2246) );
  NAND U2440 ( .A(n2247), .B(n2246), .Z(n2263) );
  AND U2441 ( .A(b[2]), .B(a[85]), .Z(n2269) );
  AND U2442 ( .A(a[86]), .B(b[1]), .Z(n2267) );
  AND U2443 ( .A(a[84]), .B(b[3]), .Z(n2266) );
  XOR U2444 ( .A(n2267), .B(n2266), .Z(n2268) );
  XOR U2445 ( .A(n2269), .B(n2268), .Z(n2272) );
  NAND U2446 ( .A(b[0]), .B(a[87]), .Z(n2273) );
  XOR U2447 ( .A(n2272), .B(n2273), .Z(n2275) );
  OR U2448 ( .A(n2249), .B(n2248), .Z(n2253) );
  NANDN U2449 ( .A(n2251), .B(n2250), .Z(n2252) );
  NAND U2450 ( .A(n2253), .B(n2252), .Z(n2274) );
  XNOR U2451 ( .A(n2275), .B(n2274), .Z(n2260) );
  NANDN U2452 ( .A(n2255), .B(n2254), .Z(n2259) );
  OR U2453 ( .A(n2257), .B(n2256), .Z(n2258) );
  NAND U2454 ( .A(n2259), .B(n2258), .Z(n2261) );
  XNOR U2455 ( .A(n2260), .B(n2261), .Z(n2262) );
  XNOR U2456 ( .A(n2263), .B(n2262), .Z(n2278) );
  XNOR U2457 ( .A(n2278), .B(sreg[339]), .Z(n2279) );
  XOR U2458 ( .A(n2280), .B(n2279), .Z(c[339]) );
  NANDN U2459 ( .A(n2261), .B(n2260), .Z(n2265) );
  NAND U2460 ( .A(n2263), .B(n2262), .Z(n2264) );
  NAND U2461 ( .A(n2265), .B(n2264), .Z(n2289) );
  AND U2462 ( .A(b[2]), .B(a[86]), .Z(n2295) );
  AND U2463 ( .A(a[87]), .B(b[1]), .Z(n2293) );
  AND U2464 ( .A(a[85]), .B(b[3]), .Z(n2292) );
  XOR U2465 ( .A(n2293), .B(n2292), .Z(n2294) );
  XOR U2466 ( .A(n2295), .B(n2294), .Z(n2298) );
  NAND U2467 ( .A(b[0]), .B(a[88]), .Z(n2299) );
  XOR U2468 ( .A(n2298), .B(n2299), .Z(n2301) );
  OR U2469 ( .A(n2267), .B(n2266), .Z(n2271) );
  NANDN U2470 ( .A(n2269), .B(n2268), .Z(n2270) );
  NAND U2471 ( .A(n2271), .B(n2270), .Z(n2300) );
  XNOR U2472 ( .A(n2301), .B(n2300), .Z(n2286) );
  NANDN U2473 ( .A(n2273), .B(n2272), .Z(n2277) );
  OR U2474 ( .A(n2275), .B(n2274), .Z(n2276) );
  NAND U2475 ( .A(n2277), .B(n2276), .Z(n2287) );
  XNOR U2476 ( .A(n2286), .B(n2287), .Z(n2288) );
  XNOR U2477 ( .A(n2289), .B(n2288), .Z(n2285) );
  NAND U2478 ( .A(n2278), .B(sreg[339]), .Z(n2282) );
  OR U2479 ( .A(n2280), .B(n2279), .Z(n2281) );
  AND U2480 ( .A(n2282), .B(n2281), .Z(n2284) );
  XNOR U2481 ( .A(n2284), .B(sreg[340]), .Z(n2283) );
  XOR U2482 ( .A(n2285), .B(n2283), .Z(c[340]) );
  NANDN U2483 ( .A(n2287), .B(n2286), .Z(n2291) );
  NAND U2484 ( .A(n2289), .B(n2288), .Z(n2290) );
  NAND U2485 ( .A(n2291), .B(n2290), .Z(n2307) );
  AND U2486 ( .A(b[2]), .B(a[87]), .Z(n2313) );
  AND U2487 ( .A(a[88]), .B(b[1]), .Z(n2311) );
  AND U2488 ( .A(a[86]), .B(b[3]), .Z(n2310) );
  XOR U2489 ( .A(n2311), .B(n2310), .Z(n2312) );
  XOR U2490 ( .A(n2313), .B(n2312), .Z(n2316) );
  NAND U2491 ( .A(b[0]), .B(a[89]), .Z(n2317) );
  XOR U2492 ( .A(n2316), .B(n2317), .Z(n2319) );
  OR U2493 ( .A(n2293), .B(n2292), .Z(n2297) );
  NANDN U2494 ( .A(n2295), .B(n2294), .Z(n2296) );
  NAND U2495 ( .A(n2297), .B(n2296), .Z(n2318) );
  XNOR U2496 ( .A(n2319), .B(n2318), .Z(n2304) );
  NANDN U2497 ( .A(n2299), .B(n2298), .Z(n2303) );
  OR U2498 ( .A(n2301), .B(n2300), .Z(n2302) );
  NAND U2499 ( .A(n2303), .B(n2302), .Z(n2305) );
  XNOR U2500 ( .A(n2304), .B(n2305), .Z(n2306) );
  XNOR U2501 ( .A(n2307), .B(n2306), .Z(n2322) );
  XNOR U2502 ( .A(n2322), .B(sreg[341]), .Z(n2324) );
  XNOR U2503 ( .A(n2323), .B(n2324), .Z(c[341]) );
  NANDN U2504 ( .A(n2305), .B(n2304), .Z(n2309) );
  NAND U2505 ( .A(n2307), .B(n2306), .Z(n2308) );
  NAND U2506 ( .A(n2309), .B(n2308), .Z(n2330) );
  AND U2507 ( .A(b[2]), .B(a[88]), .Z(n2336) );
  AND U2508 ( .A(a[89]), .B(b[1]), .Z(n2334) );
  AND U2509 ( .A(a[87]), .B(b[3]), .Z(n2333) );
  XOR U2510 ( .A(n2334), .B(n2333), .Z(n2335) );
  XOR U2511 ( .A(n2336), .B(n2335), .Z(n2339) );
  NAND U2512 ( .A(b[0]), .B(a[90]), .Z(n2340) );
  XOR U2513 ( .A(n2339), .B(n2340), .Z(n2342) );
  OR U2514 ( .A(n2311), .B(n2310), .Z(n2315) );
  NANDN U2515 ( .A(n2313), .B(n2312), .Z(n2314) );
  NAND U2516 ( .A(n2315), .B(n2314), .Z(n2341) );
  XNOR U2517 ( .A(n2342), .B(n2341), .Z(n2327) );
  NANDN U2518 ( .A(n2317), .B(n2316), .Z(n2321) );
  OR U2519 ( .A(n2319), .B(n2318), .Z(n2320) );
  NAND U2520 ( .A(n2321), .B(n2320), .Z(n2328) );
  XNOR U2521 ( .A(n2327), .B(n2328), .Z(n2329) );
  XNOR U2522 ( .A(n2330), .B(n2329), .Z(n2345) );
  XOR U2523 ( .A(sreg[342]), .B(n2345), .Z(n2346) );
  NAND U2524 ( .A(n2322), .B(sreg[341]), .Z(n2326) );
  NANDN U2525 ( .A(n2324), .B(n2323), .Z(n2325) );
  NAND U2526 ( .A(n2326), .B(n2325), .Z(n2347) );
  XOR U2527 ( .A(n2346), .B(n2347), .Z(c[342]) );
  NANDN U2528 ( .A(n2328), .B(n2327), .Z(n2332) );
  NAND U2529 ( .A(n2330), .B(n2329), .Z(n2331) );
  NAND U2530 ( .A(n2332), .B(n2331), .Z(n2356) );
  AND U2531 ( .A(b[2]), .B(a[89]), .Z(n2362) );
  AND U2532 ( .A(a[90]), .B(b[1]), .Z(n2360) );
  AND U2533 ( .A(a[88]), .B(b[3]), .Z(n2359) );
  XOR U2534 ( .A(n2360), .B(n2359), .Z(n2361) );
  XOR U2535 ( .A(n2362), .B(n2361), .Z(n2365) );
  NAND U2536 ( .A(b[0]), .B(a[91]), .Z(n2366) );
  XOR U2537 ( .A(n2365), .B(n2366), .Z(n2368) );
  OR U2538 ( .A(n2334), .B(n2333), .Z(n2338) );
  NANDN U2539 ( .A(n2336), .B(n2335), .Z(n2337) );
  NAND U2540 ( .A(n2338), .B(n2337), .Z(n2367) );
  XNOR U2541 ( .A(n2368), .B(n2367), .Z(n2353) );
  NANDN U2542 ( .A(n2340), .B(n2339), .Z(n2344) );
  OR U2543 ( .A(n2342), .B(n2341), .Z(n2343) );
  NAND U2544 ( .A(n2344), .B(n2343), .Z(n2354) );
  XNOR U2545 ( .A(n2353), .B(n2354), .Z(n2355) );
  XOR U2546 ( .A(n2356), .B(n2355), .Z(n2352) );
  OR U2547 ( .A(n2345), .B(sreg[342]), .Z(n2349) );
  NANDN U2548 ( .A(n2347), .B(n2346), .Z(n2348) );
  AND U2549 ( .A(n2349), .B(n2348), .Z(n2351) );
  XNOR U2550 ( .A(sreg[343]), .B(n2351), .Z(n2350) );
  XOR U2551 ( .A(n2352), .B(n2350), .Z(c[343]) );
  NANDN U2552 ( .A(n2354), .B(n2353), .Z(n2358) );
  NAND U2553 ( .A(n2356), .B(n2355), .Z(n2357) );
  NAND U2554 ( .A(n2358), .B(n2357), .Z(n2374) );
  AND U2555 ( .A(b[2]), .B(a[90]), .Z(n2380) );
  AND U2556 ( .A(a[91]), .B(b[1]), .Z(n2378) );
  AND U2557 ( .A(a[89]), .B(b[3]), .Z(n2377) );
  XOR U2558 ( .A(n2378), .B(n2377), .Z(n2379) );
  XOR U2559 ( .A(n2380), .B(n2379), .Z(n2383) );
  NAND U2560 ( .A(b[0]), .B(a[92]), .Z(n2384) );
  XOR U2561 ( .A(n2383), .B(n2384), .Z(n2386) );
  OR U2562 ( .A(n2360), .B(n2359), .Z(n2364) );
  NANDN U2563 ( .A(n2362), .B(n2361), .Z(n2363) );
  NAND U2564 ( .A(n2364), .B(n2363), .Z(n2385) );
  XNOR U2565 ( .A(n2386), .B(n2385), .Z(n2371) );
  NANDN U2566 ( .A(n2366), .B(n2365), .Z(n2370) );
  OR U2567 ( .A(n2368), .B(n2367), .Z(n2369) );
  NAND U2568 ( .A(n2370), .B(n2369), .Z(n2372) );
  XNOR U2569 ( .A(n2371), .B(n2372), .Z(n2373) );
  XNOR U2570 ( .A(n2374), .B(n2373), .Z(n2389) );
  XNOR U2571 ( .A(n2389), .B(sreg[344]), .Z(n2390) );
  XOR U2572 ( .A(n2391), .B(n2390), .Z(c[344]) );
  NANDN U2573 ( .A(n2372), .B(n2371), .Z(n2376) );
  NAND U2574 ( .A(n2374), .B(n2373), .Z(n2375) );
  NAND U2575 ( .A(n2376), .B(n2375), .Z(n2398) );
  AND U2576 ( .A(b[2]), .B(a[91]), .Z(n2404) );
  AND U2577 ( .A(a[92]), .B(b[1]), .Z(n2402) );
  AND U2578 ( .A(a[90]), .B(b[3]), .Z(n2401) );
  XOR U2579 ( .A(n2402), .B(n2401), .Z(n2403) );
  XOR U2580 ( .A(n2404), .B(n2403), .Z(n2407) );
  NAND U2581 ( .A(b[0]), .B(a[93]), .Z(n2408) );
  XOR U2582 ( .A(n2407), .B(n2408), .Z(n2410) );
  OR U2583 ( .A(n2378), .B(n2377), .Z(n2382) );
  NANDN U2584 ( .A(n2380), .B(n2379), .Z(n2381) );
  NAND U2585 ( .A(n2382), .B(n2381), .Z(n2409) );
  XNOR U2586 ( .A(n2410), .B(n2409), .Z(n2395) );
  NANDN U2587 ( .A(n2384), .B(n2383), .Z(n2388) );
  OR U2588 ( .A(n2386), .B(n2385), .Z(n2387) );
  NAND U2589 ( .A(n2388), .B(n2387), .Z(n2396) );
  XNOR U2590 ( .A(n2395), .B(n2396), .Z(n2397) );
  XOR U2591 ( .A(n2398), .B(n2397), .Z(n2414) );
  NAND U2592 ( .A(n2389), .B(sreg[344]), .Z(n2393) );
  OR U2593 ( .A(n2391), .B(n2390), .Z(n2392) );
  NAND U2594 ( .A(n2393), .B(n2392), .Z(n2413) );
  XNOR U2595 ( .A(sreg[345]), .B(n2413), .Z(n2394) );
  XOR U2596 ( .A(n2414), .B(n2394), .Z(c[345]) );
  NANDN U2597 ( .A(n2396), .B(n2395), .Z(n2400) );
  NAND U2598 ( .A(n2398), .B(n2397), .Z(n2399) );
  NAND U2599 ( .A(n2400), .B(n2399), .Z(n2419) );
  AND U2600 ( .A(b[2]), .B(a[92]), .Z(n2425) );
  AND U2601 ( .A(a[93]), .B(b[1]), .Z(n2423) );
  AND U2602 ( .A(a[91]), .B(b[3]), .Z(n2422) );
  XOR U2603 ( .A(n2423), .B(n2422), .Z(n2424) );
  XOR U2604 ( .A(n2425), .B(n2424), .Z(n2428) );
  NAND U2605 ( .A(b[0]), .B(a[94]), .Z(n2429) );
  XOR U2606 ( .A(n2428), .B(n2429), .Z(n2431) );
  OR U2607 ( .A(n2402), .B(n2401), .Z(n2406) );
  NANDN U2608 ( .A(n2404), .B(n2403), .Z(n2405) );
  NAND U2609 ( .A(n2406), .B(n2405), .Z(n2430) );
  XNOR U2610 ( .A(n2431), .B(n2430), .Z(n2416) );
  NANDN U2611 ( .A(n2408), .B(n2407), .Z(n2412) );
  OR U2612 ( .A(n2410), .B(n2409), .Z(n2411) );
  NAND U2613 ( .A(n2412), .B(n2411), .Z(n2417) );
  XNOR U2614 ( .A(n2416), .B(n2417), .Z(n2418) );
  XOR U2615 ( .A(n2419), .B(n2418), .Z(n2435) );
  XNOR U2616 ( .A(sreg[346]), .B(n2434), .Z(n2415) );
  XOR U2617 ( .A(n2435), .B(n2415), .Z(c[346]) );
  NANDN U2618 ( .A(n2417), .B(n2416), .Z(n2421) );
  NAND U2619 ( .A(n2419), .B(n2418), .Z(n2420) );
  NAND U2620 ( .A(n2421), .B(n2420), .Z(n2442) );
  AND U2621 ( .A(b[2]), .B(a[93]), .Z(n2448) );
  AND U2622 ( .A(a[94]), .B(b[1]), .Z(n2446) );
  AND U2623 ( .A(a[92]), .B(b[3]), .Z(n2445) );
  XOR U2624 ( .A(n2446), .B(n2445), .Z(n2447) );
  XOR U2625 ( .A(n2448), .B(n2447), .Z(n2451) );
  NAND U2626 ( .A(b[0]), .B(a[95]), .Z(n2452) );
  XOR U2627 ( .A(n2451), .B(n2452), .Z(n2454) );
  OR U2628 ( .A(n2423), .B(n2422), .Z(n2427) );
  NANDN U2629 ( .A(n2425), .B(n2424), .Z(n2426) );
  NAND U2630 ( .A(n2427), .B(n2426), .Z(n2453) );
  XNOR U2631 ( .A(n2454), .B(n2453), .Z(n2439) );
  NANDN U2632 ( .A(n2429), .B(n2428), .Z(n2433) );
  OR U2633 ( .A(n2431), .B(n2430), .Z(n2432) );
  NAND U2634 ( .A(n2433), .B(n2432), .Z(n2440) );
  XNOR U2635 ( .A(n2439), .B(n2440), .Z(n2441) );
  XNOR U2636 ( .A(n2442), .B(n2441), .Z(n2438) );
  XOR U2637 ( .A(n2437), .B(sreg[347]), .Z(n2436) );
  XOR U2638 ( .A(n2438), .B(n2436), .Z(c[347]) );
  NANDN U2639 ( .A(n2440), .B(n2439), .Z(n2444) );
  NAND U2640 ( .A(n2442), .B(n2441), .Z(n2443) );
  NAND U2641 ( .A(n2444), .B(n2443), .Z(n2465) );
  AND U2642 ( .A(b[2]), .B(a[94]), .Z(n2471) );
  AND U2643 ( .A(a[95]), .B(b[1]), .Z(n2469) );
  AND U2644 ( .A(a[93]), .B(b[3]), .Z(n2468) );
  XOR U2645 ( .A(n2469), .B(n2468), .Z(n2470) );
  XOR U2646 ( .A(n2471), .B(n2470), .Z(n2474) );
  NAND U2647 ( .A(b[0]), .B(a[96]), .Z(n2475) );
  XOR U2648 ( .A(n2474), .B(n2475), .Z(n2477) );
  OR U2649 ( .A(n2446), .B(n2445), .Z(n2450) );
  NANDN U2650 ( .A(n2448), .B(n2447), .Z(n2449) );
  NAND U2651 ( .A(n2450), .B(n2449), .Z(n2476) );
  XNOR U2652 ( .A(n2477), .B(n2476), .Z(n2462) );
  NANDN U2653 ( .A(n2452), .B(n2451), .Z(n2456) );
  OR U2654 ( .A(n2454), .B(n2453), .Z(n2455) );
  NAND U2655 ( .A(n2456), .B(n2455), .Z(n2463) );
  XNOR U2656 ( .A(n2462), .B(n2463), .Z(n2464) );
  XNOR U2657 ( .A(n2465), .B(n2464), .Z(n2457) );
  XOR U2658 ( .A(sreg[348]), .B(n2457), .Z(n2458) );
  XOR U2659 ( .A(n2459), .B(n2458), .Z(c[348]) );
  OR U2660 ( .A(n2457), .B(sreg[348]), .Z(n2461) );
  NANDN U2661 ( .A(n2459), .B(n2458), .Z(n2460) );
  AND U2662 ( .A(n2461), .B(n2460), .Z(n2481) );
  NANDN U2663 ( .A(n2463), .B(n2462), .Z(n2467) );
  NAND U2664 ( .A(n2465), .B(n2464), .Z(n2466) );
  NAND U2665 ( .A(n2467), .B(n2466), .Z(n2486) );
  AND U2666 ( .A(b[2]), .B(a[95]), .Z(n2498) );
  AND U2667 ( .A(a[96]), .B(b[1]), .Z(n2496) );
  AND U2668 ( .A(a[94]), .B(b[3]), .Z(n2495) );
  XOR U2669 ( .A(n2496), .B(n2495), .Z(n2497) );
  XOR U2670 ( .A(n2498), .B(n2497), .Z(n2489) );
  NAND U2671 ( .A(b[0]), .B(a[97]), .Z(n2490) );
  XOR U2672 ( .A(n2489), .B(n2490), .Z(n2492) );
  OR U2673 ( .A(n2469), .B(n2468), .Z(n2473) );
  NANDN U2674 ( .A(n2471), .B(n2470), .Z(n2472) );
  NAND U2675 ( .A(n2473), .B(n2472), .Z(n2491) );
  XNOR U2676 ( .A(n2492), .B(n2491), .Z(n2483) );
  NANDN U2677 ( .A(n2475), .B(n2474), .Z(n2479) );
  OR U2678 ( .A(n2477), .B(n2476), .Z(n2478) );
  NAND U2679 ( .A(n2479), .B(n2478), .Z(n2484) );
  XNOR U2680 ( .A(n2483), .B(n2484), .Z(n2485) );
  XNOR U2681 ( .A(n2486), .B(n2485), .Z(n2482) );
  XOR U2682 ( .A(sreg[349]), .B(n2482), .Z(n2480) );
  XOR U2683 ( .A(n2481), .B(n2480), .Z(c[349]) );
  NANDN U2684 ( .A(n2484), .B(n2483), .Z(n2488) );
  NAND U2685 ( .A(n2486), .B(n2485), .Z(n2487) );
  AND U2686 ( .A(n2488), .B(n2487), .Z(n2504) );
  NANDN U2687 ( .A(n2490), .B(n2489), .Z(n2494) );
  OR U2688 ( .A(n2492), .B(n2491), .Z(n2493) );
  AND U2689 ( .A(n2494), .B(n2493), .Z(n2503) );
  AND U2690 ( .A(b[2]), .B(a[96]), .Z(n2508) );
  AND U2691 ( .A(a[97]), .B(b[1]), .Z(n2506) );
  AND U2692 ( .A(a[95]), .B(b[3]), .Z(n2505) );
  XOR U2693 ( .A(n2506), .B(n2505), .Z(n2507) );
  XOR U2694 ( .A(n2508), .B(n2507), .Z(n2511) );
  NAND U2695 ( .A(b[0]), .B(a[98]), .Z(n2512) );
  XOR U2696 ( .A(n2511), .B(n2512), .Z(n2514) );
  OR U2697 ( .A(n2496), .B(n2495), .Z(n2500) );
  NANDN U2698 ( .A(n2498), .B(n2497), .Z(n2499) );
  NAND U2699 ( .A(n2500), .B(n2499), .Z(n2513) );
  XOR U2700 ( .A(n2514), .B(n2513), .Z(n2502) );
  XNOR U2701 ( .A(n2503), .B(n2502), .Z(n2501) );
  XOR U2702 ( .A(n2504), .B(n2501), .Z(n2517) );
  XOR U2703 ( .A(n2517), .B(sreg[350]), .Z(n2518) );
  XOR U2704 ( .A(n2519), .B(n2518), .Z(c[350]) );
  AND U2705 ( .A(b[2]), .B(a[97]), .Z(n2532) );
  AND U2706 ( .A(a[98]), .B(b[1]), .Z(n2530) );
  AND U2707 ( .A(a[96]), .B(b[3]), .Z(n2529) );
  XOR U2708 ( .A(n2530), .B(n2529), .Z(n2531) );
  XOR U2709 ( .A(n2532), .B(n2531), .Z(n2535) );
  NAND U2710 ( .A(b[0]), .B(a[99]), .Z(n2536) );
  XOR U2711 ( .A(n2535), .B(n2536), .Z(n2538) );
  OR U2712 ( .A(n2506), .B(n2505), .Z(n2510) );
  NANDN U2713 ( .A(n2508), .B(n2507), .Z(n2509) );
  NAND U2714 ( .A(n2510), .B(n2509), .Z(n2537) );
  XNOR U2715 ( .A(n2538), .B(n2537), .Z(n2523) );
  NANDN U2716 ( .A(n2512), .B(n2511), .Z(n2516) );
  OR U2717 ( .A(n2514), .B(n2513), .Z(n2515) );
  NAND U2718 ( .A(n2516), .B(n2515), .Z(n2524) );
  XNOR U2719 ( .A(n2523), .B(n2524), .Z(n2525) );
  XOR U2720 ( .A(n2526), .B(n2525), .Z(n2542) );
  NAND U2721 ( .A(sreg[350]), .B(n2517), .Z(n2521) );
  NAND U2722 ( .A(n2519), .B(n2518), .Z(n2520) );
  NAND U2723 ( .A(n2521), .B(n2520), .Z(n2541) );
  XNOR U2724 ( .A(sreg[351]), .B(n2541), .Z(n2522) );
  XNOR U2725 ( .A(n2542), .B(n2522), .Z(c[351]) );
  NANDN U2726 ( .A(n2524), .B(n2523), .Z(n2528) );
  NANDN U2727 ( .A(n2526), .B(n2525), .Z(n2527) );
  NAND U2728 ( .A(n2528), .B(n2527), .Z(n2547) );
  AND U2729 ( .A(b[2]), .B(a[98]), .Z(n2553) );
  AND U2730 ( .A(a[99]), .B(b[1]), .Z(n2551) );
  AND U2731 ( .A(a[97]), .B(b[3]), .Z(n2550) );
  XOR U2732 ( .A(n2551), .B(n2550), .Z(n2552) );
  XOR U2733 ( .A(n2553), .B(n2552), .Z(n2556) );
  NAND U2734 ( .A(b[0]), .B(a[100]), .Z(n2557) );
  XOR U2735 ( .A(n2556), .B(n2557), .Z(n2559) );
  OR U2736 ( .A(n2530), .B(n2529), .Z(n2534) );
  NANDN U2737 ( .A(n2532), .B(n2531), .Z(n2533) );
  NAND U2738 ( .A(n2534), .B(n2533), .Z(n2558) );
  XNOR U2739 ( .A(n2559), .B(n2558), .Z(n2544) );
  NANDN U2740 ( .A(n2536), .B(n2535), .Z(n2540) );
  OR U2741 ( .A(n2538), .B(n2537), .Z(n2539) );
  NAND U2742 ( .A(n2540), .B(n2539), .Z(n2545) );
  XNOR U2743 ( .A(n2544), .B(n2545), .Z(n2546) );
  XOR U2744 ( .A(n2547), .B(n2546), .Z(n2564) );
  XNOR U2745 ( .A(sreg[352]), .B(n2563), .Z(n2543) );
  XOR U2746 ( .A(n2564), .B(n2543), .Z(c[352]) );
  NANDN U2747 ( .A(n2545), .B(n2544), .Z(n2549) );
  NAND U2748 ( .A(n2547), .B(n2546), .Z(n2548) );
  NAND U2749 ( .A(n2549), .B(n2548), .Z(n2570) );
  AND U2750 ( .A(b[2]), .B(a[99]), .Z(n2574) );
  AND U2751 ( .A(a[100]), .B(b[1]), .Z(n2572) );
  AND U2752 ( .A(a[98]), .B(b[3]), .Z(n2571) );
  XOR U2753 ( .A(n2572), .B(n2571), .Z(n2573) );
  XOR U2754 ( .A(n2574), .B(n2573), .Z(n2577) );
  NAND U2755 ( .A(b[0]), .B(a[101]), .Z(n2578) );
  XOR U2756 ( .A(n2577), .B(n2578), .Z(n2579) );
  OR U2757 ( .A(n2551), .B(n2550), .Z(n2555) );
  NANDN U2758 ( .A(n2553), .B(n2552), .Z(n2554) );
  AND U2759 ( .A(n2555), .B(n2554), .Z(n2580) );
  XOR U2760 ( .A(n2579), .B(n2580), .Z(n2568) );
  NANDN U2761 ( .A(n2557), .B(n2556), .Z(n2561) );
  OR U2762 ( .A(n2559), .B(n2558), .Z(n2560) );
  AND U2763 ( .A(n2561), .B(n2560), .Z(n2569) );
  XOR U2764 ( .A(n2568), .B(n2569), .Z(n2562) );
  XOR U2765 ( .A(n2570), .B(n2562), .Z(n2567) );
  XOR U2766 ( .A(n2566), .B(sreg[353]), .Z(n2565) );
  XNOR U2767 ( .A(n2567), .B(n2565), .Z(c[353]) );
  AND U2768 ( .A(b[2]), .B(a[100]), .Z(n2590) );
  AND U2769 ( .A(a[101]), .B(b[1]), .Z(n2588) );
  AND U2770 ( .A(a[99]), .B(b[3]), .Z(n2587) );
  XOR U2771 ( .A(n2588), .B(n2587), .Z(n2589) );
  XOR U2772 ( .A(n2590), .B(n2589), .Z(n2593) );
  NAND U2773 ( .A(b[0]), .B(a[102]), .Z(n2594) );
  XOR U2774 ( .A(n2593), .B(n2594), .Z(n2596) );
  OR U2775 ( .A(n2572), .B(n2571), .Z(n2576) );
  NANDN U2776 ( .A(n2574), .B(n2573), .Z(n2575) );
  NAND U2777 ( .A(n2576), .B(n2575), .Z(n2595) );
  XNOR U2778 ( .A(n2596), .B(n2595), .Z(n2581) );
  XNOR U2779 ( .A(n2581), .B(n2582), .Z(n2584) );
  XOR U2780 ( .A(n2583), .B(n2584), .Z(n2599) );
  XOR U2781 ( .A(n2599), .B(sreg[354]), .Z(n2601) );
  XNOR U2782 ( .A(n2600), .B(n2601), .Z(c[354]) );
  NANDN U2783 ( .A(n2582), .B(n2581), .Z(n2586) );
  NAND U2784 ( .A(n2584), .B(n2583), .Z(n2585) );
  NAND U2785 ( .A(n2586), .B(n2585), .Z(n2619) );
  AND U2786 ( .A(b[2]), .B(a[101]), .Z(n2613) );
  AND U2787 ( .A(a[102]), .B(b[1]), .Z(n2611) );
  AND U2788 ( .A(a[100]), .B(b[3]), .Z(n2610) );
  XOR U2789 ( .A(n2611), .B(n2610), .Z(n2612) );
  XOR U2790 ( .A(n2613), .B(n2612), .Z(n2604) );
  NAND U2791 ( .A(b[0]), .B(a[103]), .Z(n2605) );
  XOR U2792 ( .A(n2604), .B(n2605), .Z(n2607) );
  OR U2793 ( .A(n2588), .B(n2587), .Z(n2592) );
  NANDN U2794 ( .A(n2590), .B(n2589), .Z(n2591) );
  NAND U2795 ( .A(n2592), .B(n2591), .Z(n2606) );
  XNOR U2796 ( .A(n2607), .B(n2606), .Z(n2616) );
  NANDN U2797 ( .A(n2594), .B(n2593), .Z(n2598) );
  OR U2798 ( .A(n2596), .B(n2595), .Z(n2597) );
  NAND U2799 ( .A(n2598), .B(n2597), .Z(n2617) );
  XNOR U2800 ( .A(n2616), .B(n2617), .Z(n2618) );
  XNOR U2801 ( .A(n2619), .B(n2618), .Z(n2622) );
  XNOR U2802 ( .A(n2622), .B(sreg[355]), .Z(n2624) );
  NANDN U2803 ( .A(n2599), .B(sreg[354]), .Z(n2603) );
  NANDN U2804 ( .A(n2601), .B(n2600), .Z(n2602) );
  AND U2805 ( .A(n2603), .B(n2602), .Z(n2623) );
  XOR U2806 ( .A(n2624), .B(n2623), .Z(c[355]) );
  NANDN U2807 ( .A(n2605), .B(n2604), .Z(n2609) );
  OR U2808 ( .A(n2607), .B(n2606), .Z(n2608) );
  NAND U2809 ( .A(n2609), .B(n2608), .Z(n2630) );
  AND U2810 ( .A(b[2]), .B(a[102]), .Z(n2639) );
  AND U2811 ( .A(a[103]), .B(b[1]), .Z(n2637) );
  AND U2812 ( .A(a[101]), .B(b[3]), .Z(n2636) );
  XOR U2813 ( .A(n2637), .B(n2636), .Z(n2638) );
  XOR U2814 ( .A(n2639), .B(n2638), .Z(n2642) );
  NAND U2815 ( .A(b[0]), .B(a[104]), .Z(n2643) );
  XNOR U2816 ( .A(n2642), .B(n2643), .Z(n2644) );
  OR U2817 ( .A(n2611), .B(n2610), .Z(n2615) );
  NANDN U2818 ( .A(n2613), .B(n2612), .Z(n2614) );
  AND U2819 ( .A(n2615), .B(n2614), .Z(n2645) );
  XNOR U2820 ( .A(n2644), .B(n2645), .Z(n2631) );
  XNOR U2821 ( .A(n2630), .B(n2631), .Z(n2632) );
  NANDN U2822 ( .A(n2617), .B(n2616), .Z(n2621) );
  NAND U2823 ( .A(n2619), .B(n2618), .Z(n2620) );
  NAND U2824 ( .A(n2621), .B(n2620), .Z(n2633) );
  XOR U2825 ( .A(n2632), .B(n2633), .Z(n2629) );
  NAND U2826 ( .A(n2622), .B(sreg[355]), .Z(n2626) );
  OR U2827 ( .A(n2624), .B(n2623), .Z(n2625) );
  AND U2828 ( .A(n2626), .B(n2625), .Z(n2628) );
  XNOR U2829 ( .A(n2628), .B(sreg[356]), .Z(n2627) );
  XNOR U2830 ( .A(n2629), .B(n2627), .Z(c[356]) );
  NANDN U2831 ( .A(n2631), .B(n2630), .Z(n2635) );
  NANDN U2832 ( .A(n2633), .B(n2632), .Z(n2634) );
  NAND U2833 ( .A(n2635), .B(n2634), .Z(n2651) );
  AND U2834 ( .A(b[2]), .B(a[103]), .Z(n2657) );
  AND U2835 ( .A(a[104]), .B(b[1]), .Z(n2655) );
  AND U2836 ( .A(a[102]), .B(b[3]), .Z(n2654) );
  XOR U2837 ( .A(n2655), .B(n2654), .Z(n2656) );
  XOR U2838 ( .A(n2657), .B(n2656), .Z(n2660) );
  NAND U2839 ( .A(b[0]), .B(a[105]), .Z(n2661) );
  XOR U2840 ( .A(n2660), .B(n2661), .Z(n2663) );
  OR U2841 ( .A(n2637), .B(n2636), .Z(n2641) );
  NANDN U2842 ( .A(n2639), .B(n2638), .Z(n2640) );
  NAND U2843 ( .A(n2641), .B(n2640), .Z(n2662) );
  XNOR U2844 ( .A(n2663), .B(n2662), .Z(n2648) );
  NANDN U2845 ( .A(n2643), .B(n2642), .Z(n2647) );
  NAND U2846 ( .A(n2645), .B(n2644), .Z(n2646) );
  NAND U2847 ( .A(n2647), .B(n2646), .Z(n2649) );
  XNOR U2848 ( .A(n2648), .B(n2649), .Z(n2650) );
  XOR U2849 ( .A(n2651), .B(n2650), .Z(n2666) );
  XNOR U2850 ( .A(n2666), .B(sreg[357]), .Z(n2668) );
  XNOR U2851 ( .A(n2667), .B(n2668), .Z(c[357]) );
  NANDN U2852 ( .A(n2649), .B(n2648), .Z(n2653) );
  NANDN U2853 ( .A(n2651), .B(n2650), .Z(n2652) );
  NAND U2854 ( .A(n2653), .B(n2652), .Z(n2674) );
  AND U2855 ( .A(b[2]), .B(a[104]), .Z(n2680) );
  AND U2856 ( .A(a[105]), .B(b[1]), .Z(n2678) );
  AND U2857 ( .A(a[103]), .B(b[3]), .Z(n2677) );
  XOR U2858 ( .A(n2678), .B(n2677), .Z(n2679) );
  XOR U2859 ( .A(n2680), .B(n2679), .Z(n2683) );
  NAND U2860 ( .A(b[0]), .B(a[106]), .Z(n2684) );
  XOR U2861 ( .A(n2683), .B(n2684), .Z(n2686) );
  OR U2862 ( .A(n2655), .B(n2654), .Z(n2659) );
  NANDN U2863 ( .A(n2657), .B(n2656), .Z(n2658) );
  NAND U2864 ( .A(n2659), .B(n2658), .Z(n2685) );
  XNOR U2865 ( .A(n2686), .B(n2685), .Z(n2671) );
  NANDN U2866 ( .A(n2661), .B(n2660), .Z(n2665) );
  OR U2867 ( .A(n2663), .B(n2662), .Z(n2664) );
  NAND U2868 ( .A(n2665), .B(n2664), .Z(n2672) );
  XNOR U2869 ( .A(n2671), .B(n2672), .Z(n2673) );
  XNOR U2870 ( .A(n2674), .B(n2673), .Z(n2689) );
  XNOR U2871 ( .A(n2689), .B(sreg[358]), .Z(n2691) );
  NAND U2872 ( .A(n2666), .B(sreg[357]), .Z(n2670) );
  NANDN U2873 ( .A(n2668), .B(n2667), .Z(n2669) );
  AND U2874 ( .A(n2670), .B(n2669), .Z(n2690) );
  XOR U2875 ( .A(n2691), .B(n2690), .Z(c[358]) );
  NANDN U2876 ( .A(n2672), .B(n2671), .Z(n2676) );
  NAND U2877 ( .A(n2674), .B(n2673), .Z(n2675) );
  NAND U2878 ( .A(n2676), .B(n2675), .Z(n2697) );
  AND U2879 ( .A(b[2]), .B(a[105]), .Z(n2703) );
  AND U2880 ( .A(a[106]), .B(b[1]), .Z(n2701) );
  AND U2881 ( .A(a[104]), .B(b[3]), .Z(n2700) );
  XOR U2882 ( .A(n2701), .B(n2700), .Z(n2702) );
  XOR U2883 ( .A(n2703), .B(n2702), .Z(n2706) );
  NAND U2884 ( .A(b[0]), .B(a[107]), .Z(n2707) );
  XOR U2885 ( .A(n2706), .B(n2707), .Z(n2709) );
  OR U2886 ( .A(n2678), .B(n2677), .Z(n2682) );
  NANDN U2887 ( .A(n2680), .B(n2679), .Z(n2681) );
  NAND U2888 ( .A(n2682), .B(n2681), .Z(n2708) );
  XNOR U2889 ( .A(n2709), .B(n2708), .Z(n2694) );
  NANDN U2890 ( .A(n2684), .B(n2683), .Z(n2688) );
  OR U2891 ( .A(n2686), .B(n2685), .Z(n2687) );
  NAND U2892 ( .A(n2688), .B(n2687), .Z(n2695) );
  XNOR U2893 ( .A(n2694), .B(n2695), .Z(n2696) );
  XNOR U2894 ( .A(n2697), .B(n2696), .Z(n2712) );
  XNOR U2895 ( .A(n2712), .B(sreg[359]), .Z(n2714) );
  NAND U2896 ( .A(n2689), .B(sreg[358]), .Z(n2693) );
  OR U2897 ( .A(n2691), .B(n2690), .Z(n2692) );
  AND U2898 ( .A(n2693), .B(n2692), .Z(n2713) );
  XOR U2899 ( .A(n2714), .B(n2713), .Z(c[359]) );
  NANDN U2900 ( .A(n2695), .B(n2694), .Z(n2699) );
  NAND U2901 ( .A(n2697), .B(n2696), .Z(n2698) );
  NAND U2902 ( .A(n2699), .B(n2698), .Z(n2720) );
  AND U2903 ( .A(b[2]), .B(a[106]), .Z(n2726) );
  AND U2904 ( .A(a[107]), .B(b[1]), .Z(n2724) );
  AND U2905 ( .A(a[105]), .B(b[3]), .Z(n2723) );
  XOR U2906 ( .A(n2724), .B(n2723), .Z(n2725) );
  XOR U2907 ( .A(n2726), .B(n2725), .Z(n2729) );
  NAND U2908 ( .A(b[0]), .B(a[108]), .Z(n2730) );
  XOR U2909 ( .A(n2729), .B(n2730), .Z(n2732) );
  OR U2910 ( .A(n2701), .B(n2700), .Z(n2705) );
  NANDN U2911 ( .A(n2703), .B(n2702), .Z(n2704) );
  NAND U2912 ( .A(n2705), .B(n2704), .Z(n2731) );
  XNOR U2913 ( .A(n2732), .B(n2731), .Z(n2717) );
  NANDN U2914 ( .A(n2707), .B(n2706), .Z(n2711) );
  OR U2915 ( .A(n2709), .B(n2708), .Z(n2710) );
  NAND U2916 ( .A(n2711), .B(n2710), .Z(n2718) );
  XNOR U2917 ( .A(n2717), .B(n2718), .Z(n2719) );
  XNOR U2918 ( .A(n2720), .B(n2719), .Z(n2735) );
  XNOR U2919 ( .A(n2735), .B(sreg[360]), .Z(n2737) );
  NAND U2920 ( .A(n2712), .B(sreg[359]), .Z(n2716) );
  OR U2921 ( .A(n2714), .B(n2713), .Z(n2715) );
  AND U2922 ( .A(n2716), .B(n2715), .Z(n2736) );
  XOR U2923 ( .A(n2737), .B(n2736), .Z(c[360]) );
  NANDN U2924 ( .A(n2718), .B(n2717), .Z(n2722) );
  NAND U2925 ( .A(n2720), .B(n2719), .Z(n2721) );
  NAND U2926 ( .A(n2722), .B(n2721), .Z(n2743) );
  AND U2927 ( .A(b[2]), .B(a[107]), .Z(n2749) );
  AND U2928 ( .A(a[108]), .B(b[1]), .Z(n2747) );
  AND U2929 ( .A(a[106]), .B(b[3]), .Z(n2746) );
  XOR U2930 ( .A(n2747), .B(n2746), .Z(n2748) );
  XOR U2931 ( .A(n2749), .B(n2748), .Z(n2752) );
  NAND U2932 ( .A(b[0]), .B(a[109]), .Z(n2753) );
  XOR U2933 ( .A(n2752), .B(n2753), .Z(n2755) );
  OR U2934 ( .A(n2724), .B(n2723), .Z(n2728) );
  NANDN U2935 ( .A(n2726), .B(n2725), .Z(n2727) );
  NAND U2936 ( .A(n2728), .B(n2727), .Z(n2754) );
  XNOR U2937 ( .A(n2755), .B(n2754), .Z(n2740) );
  NANDN U2938 ( .A(n2730), .B(n2729), .Z(n2734) );
  OR U2939 ( .A(n2732), .B(n2731), .Z(n2733) );
  NAND U2940 ( .A(n2734), .B(n2733), .Z(n2741) );
  XNOR U2941 ( .A(n2740), .B(n2741), .Z(n2742) );
  XNOR U2942 ( .A(n2743), .B(n2742), .Z(n2758) );
  XNOR U2943 ( .A(n2758), .B(sreg[361]), .Z(n2760) );
  NAND U2944 ( .A(n2735), .B(sreg[360]), .Z(n2739) );
  OR U2945 ( .A(n2737), .B(n2736), .Z(n2738) );
  AND U2946 ( .A(n2739), .B(n2738), .Z(n2759) );
  XOR U2947 ( .A(n2760), .B(n2759), .Z(c[361]) );
  NANDN U2948 ( .A(n2741), .B(n2740), .Z(n2745) );
  NAND U2949 ( .A(n2743), .B(n2742), .Z(n2744) );
  NAND U2950 ( .A(n2745), .B(n2744), .Z(n2766) );
  AND U2951 ( .A(b[2]), .B(a[108]), .Z(n2772) );
  AND U2952 ( .A(a[109]), .B(b[1]), .Z(n2770) );
  AND U2953 ( .A(a[107]), .B(b[3]), .Z(n2769) );
  XOR U2954 ( .A(n2770), .B(n2769), .Z(n2771) );
  XOR U2955 ( .A(n2772), .B(n2771), .Z(n2775) );
  NAND U2956 ( .A(b[0]), .B(a[110]), .Z(n2776) );
  XOR U2957 ( .A(n2775), .B(n2776), .Z(n2778) );
  OR U2958 ( .A(n2747), .B(n2746), .Z(n2751) );
  NANDN U2959 ( .A(n2749), .B(n2748), .Z(n2750) );
  NAND U2960 ( .A(n2751), .B(n2750), .Z(n2777) );
  XNOR U2961 ( .A(n2778), .B(n2777), .Z(n2763) );
  NANDN U2962 ( .A(n2753), .B(n2752), .Z(n2757) );
  OR U2963 ( .A(n2755), .B(n2754), .Z(n2756) );
  NAND U2964 ( .A(n2757), .B(n2756), .Z(n2764) );
  XNOR U2965 ( .A(n2763), .B(n2764), .Z(n2765) );
  XNOR U2966 ( .A(n2766), .B(n2765), .Z(n2781) );
  XNOR U2967 ( .A(n2781), .B(sreg[362]), .Z(n2783) );
  NAND U2968 ( .A(n2758), .B(sreg[361]), .Z(n2762) );
  OR U2969 ( .A(n2760), .B(n2759), .Z(n2761) );
  AND U2970 ( .A(n2762), .B(n2761), .Z(n2782) );
  XOR U2971 ( .A(n2783), .B(n2782), .Z(c[362]) );
  NANDN U2972 ( .A(n2764), .B(n2763), .Z(n2768) );
  NAND U2973 ( .A(n2766), .B(n2765), .Z(n2767) );
  NAND U2974 ( .A(n2768), .B(n2767), .Z(n2789) );
  AND U2975 ( .A(b[2]), .B(a[109]), .Z(n2795) );
  AND U2976 ( .A(a[110]), .B(b[1]), .Z(n2793) );
  AND U2977 ( .A(a[108]), .B(b[3]), .Z(n2792) );
  XOR U2978 ( .A(n2793), .B(n2792), .Z(n2794) );
  XOR U2979 ( .A(n2795), .B(n2794), .Z(n2798) );
  NAND U2980 ( .A(b[0]), .B(a[111]), .Z(n2799) );
  XOR U2981 ( .A(n2798), .B(n2799), .Z(n2801) );
  OR U2982 ( .A(n2770), .B(n2769), .Z(n2774) );
  NANDN U2983 ( .A(n2772), .B(n2771), .Z(n2773) );
  NAND U2984 ( .A(n2774), .B(n2773), .Z(n2800) );
  XNOR U2985 ( .A(n2801), .B(n2800), .Z(n2786) );
  NANDN U2986 ( .A(n2776), .B(n2775), .Z(n2780) );
  OR U2987 ( .A(n2778), .B(n2777), .Z(n2779) );
  NAND U2988 ( .A(n2780), .B(n2779), .Z(n2787) );
  XNOR U2989 ( .A(n2786), .B(n2787), .Z(n2788) );
  XNOR U2990 ( .A(n2789), .B(n2788), .Z(n2804) );
  XNOR U2991 ( .A(n2804), .B(sreg[363]), .Z(n2806) );
  NAND U2992 ( .A(n2781), .B(sreg[362]), .Z(n2785) );
  OR U2993 ( .A(n2783), .B(n2782), .Z(n2784) );
  AND U2994 ( .A(n2785), .B(n2784), .Z(n2805) );
  XOR U2995 ( .A(n2806), .B(n2805), .Z(c[363]) );
  NANDN U2996 ( .A(n2787), .B(n2786), .Z(n2791) );
  NAND U2997 ( .A(n2789), .B(n2788), .Z(n2790) );
  NAND U2998 ( .A(n2791), .B(n2790), .Z(n2813) );
  AND U2999 ( .A(b[2]), .B(a[110]), .Z(n2819) );
  AND U3000 ( .A(a[111]), .B(b[1]), .Z(n2817) );
  AND U3001 ( .A(a[109]), .B(b[3]), .Z(n2816) );
  XOR U3002 ( .A(n2817), .B(n2816), .Z(n2818) );
  XOR U3003 ( .A(n2819), .B(n2818), .Z(n2822) );
  NAND U3004 ( .A(b[0]), .B(a[112]), .Z(n2823) );
  XOR U3005 ( .A(n2822), .B(n2823), .Z(n2825) );
  OR U3006 ( .A(n2793), .B(n2792), .Z(n2797) );
  NANDN U3007 ( .A(n2795), .B(n2794), .Z(n2796) );
  NAND U3008 ( .A(n2797), .B(n2796), .Z(n2824) );
  XNOR U3009 ( .A(n2825), .B(n2824), .Z(n2810) );
  NANDN U3010 ( .A(n2799), .B(n2798), .Z(n2803) );
  OR U3011 ( .A(n2801), .B(n2800), .Z(n2802) );
  NAND U3012 ( .A(n2803), .B(n2802), .Z(n2811) );
  XNOR U3013 ( .A(n2810), .B(n2811), .Z(n2812) );
  XOR U3014 ( .A(n2813), .B(n2812), .Z(n2829) );
  NAND U3015 ( .A(n2804), .B(sreg[363]), .Z(n2808) );
  OR U3016 ( .A(n2806), .B(n2805), .Z(n2807) );
  NAND U3017 ( .A(n2808), .B(n2807), .Z(n2828) );
  XNOR U3018 ( .A(sreg[364]), .B(n2828), .Z(n2809) );
  XOR U3019 ( .A(n2829), .B(n2809), .Z(c[364]) );
  NANDN U3020 ( .A(n2811), .B(n2810), .Z(n2815) );
  NAND U3021 ( .A(n2813), .B(n2812), .Z(n2814) );
  NAND U3022 ( .A(n2815), .B(n2814), .Z(n2834) );
  AND U3023 ( .A(b[2]), .B(a[111]), .Z(n2840) );
  AND U3024 ( .A(a[112]), .B(b[1]), .Z(n2838) );
  AND U3025 ( .A(a[110]), .B(b[3]), .Z(n2837) );
  XOR U3026 ( .A(n2838), .B(n2837), .Z(n2839) );
  XOR U3027 ( .A(n2840), .B(n2839), .Z(n2843) );
  NAND U3028 ( .A(b[0]), .B(a[113]), .Z(n2844) );
  XOR U3029 ( .A(n2843), .B(n2844), .Z(n2846) );
  OR U3030 ( .A(n2817), .B(n2816), .Z(n2821) );
  NANDN U3031 ( .A(n2819), .B(n2818), .Z(n2820) );
  NAND U3032 ( .A(n2821), .B(n2820), .Z(n2845) );
  XNOR U3033 ( .A(n2846), .B(n2845), .Z(n2831) );
  NANDN U3034 ( .A(n2823), .B(n2822), .Z(n2827) );
  OR U3035 ( .A(n2825), .B(n2824), .Z(n2826) );
  NAND U3036 ( .A(n2827), .B(n2826), .Z(n2832) );
  XNOR U3037 ( .A(n2831), .B(n2832), .Z(n2833) );
  XOR U3038 ( .A(n2834), .B(n2833), .Z(n2850) );
  XNOR U3039 ( .A(sreg[365]), .B(n2849), .Z(n2830) );
  XOR U3040 ( .A(n2850), .B(n2830), .Z(c[365]) );
  NANDN U3041 ( .A(n2832), .B(n2831), .Z(n2836) );
  NAND U3042 ( .A(n2834), .B(n2833), .Z(n2835) );
  NAND U3043 ( .A(n2836), .B(n2835), .Z(n2857) );
  AND U3044 ( .A(b[2]), .B(a[112]), .Z(n2863) );
  AND U3045 ( .A(a[113]), .B(b[1]), .Z(n2861) );
  AND U3046 ( .A(a[111]), .B(b[3]), .Z(n2860) );
  XOR U3047 ( .A(n2861), .B(n2860), .Z(n2862) );
  XOR U3048 ( .A(n2863), .B(n2862), .Z(n2866) );
  NAND U3049 ( .A(b[0]), .B(a[114]), .Z(n2867) );
  XOR U3050 ( .A(n2866), .B(n2867), .Z(n2869) );
  OR U3051 ( .A(n2838), .B(n2837), .Z(n2842) );
  NANDN U3052 ( .A(n2840), .B(n2839), .Z(n2841) );
  NAND U3053 ( .A(n2842), .B(n2841), .Z(n2868) );
  XNOR U3054 ( .A(n2869), .B(n2868), .Z(n2854) );
  NANDN U3055 ( .A(n2844), .B(n2843), .Z(n2848) );
  OR U3056 ( .A(n2846), .B(n2845), .Z(n2847) );
  NAND U3057 ( .A(n2848), .B(n2847), .Z(n2855) );
  XNOR U3058 ( .A(n2854), .B(n2855), .Z(n2856) );
  XOR U3059 ( .A(n2857), .B(n2856), .Z(n2853) );
  XNOR U3060 ( .A(sreg[366]), .B(n2852), .Z(n2851) );
  XOR U3061 ( .A(n2853), .B(n2851), .Z(c[366]) );
  NANDN U3062 ( .A(n2855), .B(n2854), .Z(n2859) );
  NAND U3063 ( .A(n2857), .B(n2856), .Z(n2858) );
  NAND U3064 ( .A(n2859), .B(n2858), .Z(n2875) );
  AND U3065 ( .A(b[2]), .B(a[113]), .Z(n2881) );
  AND U3066 ( .A(a[114]), .B(b[1]), .Z(n2879) );
  AND U3067 ( .A(a[112]), .B(b[3]), .Z(n2878) );
  XOR U3068 ( .A(n2879), .B(n2878), .Z(n2880) );
  XOR U3069 ( .A(n2881), .B(n2880), .Z(n2884) );
  NAND U3070 ( .A(b[0]), .B(a[115]), .Z(n2885) );
  XOR U3071 ( .A(n2884), .B(n2885), .Z(n2887) );
  OR U3072 ( .A(n2861), .B(n2860), .Z(n2865) );
  NANDN U3073 ( .A(n2863), .B(n2862), .Z(n2864) );
  NAND U3074 ( .A(n2865), .B(n2864), .Z(n2886) );
  XNOR U3075 ( .A(n2887), .B(n2886), .Z(n2872) );
  NANDN U3076 ( .A(n2867), .B(n2866), .Z(n2871) );
  OR U3077 ( .A(n2869), .B(n2868), .Z(n2870) );
  NAND U3078 ( .A(n2871), .B(n2870), .Z(n2873) );
  XNOR U3079 ( .A(n2872), .B(n2873), .Z(n2874) );
  XNOR U3080 ( .A(n2875), .B(n2874), .Z(n2890) );
  XNOR U3081 ( .A(n2890), .B(sreg[367]), .Z(n2891) );
  XOR U3082 ( .A(n2892), .B(n2891), .Z(c[367]) );
  NANDN U3083 ( .A(n2873), .B(n2872), .Z(n2877) );
  NAND U3084 ( .A(n2875), .B(n2874), .Z(n2876) );
  NAND U3085 ( .A(n2877), .B(n2876), .Z(n2901) );
  AND U3086 ( .A(b[2]), .B(a[114]), .Z(n2913) );
  AND U3087 ( .A(a[115]), .B(b[1]), .Z(n2911) );
  AND U3088 ( .A(a[113]), .B(b[3]), .Z(n2910) );
  XOR U3089 ( .A(n2911), .B(n2910), .Z(n2912) );
  XOR U3090 ( .A(n2913), .B(n2912), .Z(n2904) );
  NAND U3091 ( .A(b[0]), .B(a[116]), .Z(n2905) );
  XOR U3092 ( .A(n2904), .B(n2905), .Z(n2907) );
  OR U3093 ( .A(n2879), .B(n2878), .Z(n2883) );
  NANDN U3094 ( .A(n2881), .B(n2880), .Z(n2882) );
  NAND U3095 ( .A(n2883), .B(n2882), .Z(n2906) );
  XNOR U3096 ( .A(n2907), .B(n2906), .Z(n2898) );
  NANDN U3097 ( .A(n2885), .B(n2884), .Z(n2889) );
  OR U3098 ( .A(n2887), .B(n2886), .Z(n2888) );
  NAND U3099 ( .A(n2889), .B(n2888), .Z(n2899) );
  XNOR U3100 ( .A(n2898), .B(n2899), .Z(n2900) );
  XOR U3101 ( .A(n2901), .B(n2900), .Z(n2897) );
  NAND U3102 ( .A(n2890), .B(sreg[367]), .Z(n2894) );
  OR U3103 ( .A(n2892), .B(n2891), .Z(n2893) );
  NAND U3104 ( .A(n2894), .B(n2893), .Z(n2896) );
  XNOR U3105 ( .A(sreg[368]), .B(n2896), .Z(n2895) );
  XOR U3106 ( .A(n2897), .B(n2895), .Z(c[368]) );
  NANDN U3107 ( .A(n2899), .B(n2898), .Z(n2903) );
  NAND U3108 ( .A(n2901), .B(n2900), .Z(n2902) );
  NAND U3109 ( .A(n2903), .B(n2902), .Z(n2936) );
  NANDN U3110 ( .A(n2905), .B(n2904), .Z(n2909) );
  OR U3111 ( .A(n2907), .B(n2906), .Z(n2908) );
  NAND U3112 ( .A(n2909), .B(n2908), .Z(n2933) );
  AND U3113 ( .A(b[2]), .B(a[115]), .Z(n2924) );
  AND U3114 ( .A(a[116]), .B(b[1]), .Z(n2922) );
  AND U3115 ( .A(a[114]), .B(b[3]), .Z(n2921) );
  XOR U3116 ( .A(n2922), .B(n2921), .Z(n2923) );
  XOR U3117 ( .A(n2924), .B(n2923), .Z(n2927) );
  NAND U3118 ( .A(b[0]), .B(a[117]), .Z(n2928) );
  XNOR U3119 ( .A(n2927), .B(n2928), .Z(n2929) );
  OR U3120 ( .A(n2911), .B(n2910), .Z(n2915) );
  NANDN U3121 ( .A(n2913), .B(n2912), .Z(n2914) );
  AND U3122 ( .A(n2915), .B(n2914), .Z(n2930) );
  XNOR U3123 ( .A(n2929), .B(n2930), .Z(n2934) );
  XNOR U3124 ( .A(n2933), .B(n2934), .Z(n2935) );
  XNOR U3125 ( .A(n2936), .B(n2935), .Z(n2916) );
  XNOR U3126 ( .A(sreg[369]), .B(n2916), .Z(n2917) );
  XOR U3127 ( .A(n2918), .B(n2917), .Z(c[369]) );
  NAND U3128 ( .A(sreg[369]), .B(n2916), .Z(n2920) );
  OR U3129 ( .A(n2918), .B(n2917), .Z(n2919) );
  NAND U3130 ( .A(n2920), .B(n2919), .Z(n2959) );
  AND U3131 ( .A(b[2]), .B(a[116]), .Z(n2948) );
  AND U3132 ( .A(a[117]), .B(b[1]), .Z(n2946) );
  AND U3133 ( .A(a[115]), .B(b[3]), .Z(n2945) );
  XOR U3134 ( .A(n2946), .B(n2945), .Z(n2947) );
  XOR U3135 ( .A(n2948), .B(n2947), .Z(n2951) );
  NAND U3136 ( .A(b[0]), .B(a[118]), .Z(n2952) );
  XOR U3137 ( .A(n2951), .B(n2952), .Z(n2954) );
  OR U3138 ( .A(n2922), .B(n2921), .Z(n2926) );
  NANDN U3139 ( .A(n2924), .B(n2923), .Z(n2925) );
  NAND U3140 ( .A(n2926), .B(n2925), .Z(n2953) );
  XNOR U3141 ( .A(n2954), .B(n2953), .Z(n2939) );
  NANDN U3142 ( .A(n2928), .B(n2927), .Z(n2932) );
  NAND U3143 ( .A(n2930), .B(n2929), .Z(n2931) );
  NAND U3144 ( .A(n2932), .B(n2931), .Z(n2940) );
  XNOR U3145 ( .A(n2939), .B(n2940), .Z(n2941) );
  NANDN U3146 ( .A(n2934), .B(n2933), .Z(n2938) );
  NANDN U3147 ( .A(n2936), .B(n2935), .Z(n2937) );
  AND U3148 ( .A(n2938), .B(n2937), .Z(n2942) );
  XNOR U3149 ( .A(n2941), .B(n2942), .Z(n2957) );
  XOR U3150 ( .A(sreg[370]), .B(n2957), .Z(n2958) );
  XOR U3151 ( .A(n2959), .B(n2958), .Z(c[370]) );
  NANDN U3152 ( .A(n2940), .B(n2939), .Z(n2944) );
  NAND U3153 ( .A(n2942), .B(n2941), .Z(n2943) );
  NAND U3154 ( .A(n2944), .B(n2943), .Z(n2980) );
  AND U3155 ( .A(b[2]), .B(a[117]), .Z(n2974) );
  AND U3156 ( .A(a[118]), .B(b[1]), .Z(n2972) );
  AND U3157 ( .A(a[116]), .B(b[3]), .Z(n2971) );
  XOR U3158 ( .A(n2972), .B(n2971), .Z(n2973) );
  XOR U3159 ( .A(n2974), .B(n2973), .Z(n2965) );
  NAND U3160 ( .A(b[0]), .B(a[119]), .Z(n2966) );
  XOR U3161 ( .A(n2965), .B(n2966), .Z(n2968) );
  OR U3162 ( .A(n2946), .B(n2945), .Z(n2950) );
  NANDN U3163 ( .A(n2948), .B(n2947), .Z(n2949) );
  NAND U3164 ( .A(n2950), .B(n2949), .Z(n2967) );
  XNOR U3165 ( .A(n2968), .B(n2967), .Z(n2977) );
  NANDN U3166 ( .A(n2952), .B(n2951), .Z(n2956) );
  OR U3167 ( .A(n2954), .B(n2953), .Z(n2955) );
  NAND U3168 ( .A(n2956), .B(n2955), .Z(n2978) );
  XNOR U3169 ( .A(n2977), .B(n2978), .Z(n2979) );
  XOR U3170 ( .A(n2980), .B(n2979), .Z(n2964) );
  OR U3171 ( .A(n2957), .B(sreg[370]), .Z(n2961) );
  NANDN U3172 ( .A(n2959), .B(n2958), .Z(n2960) );
  AND U3173 ( .A(n2961), .B(n2960), .Z(n2963) );
  XNOR U3174 ( .A(sreg[371]), .B(n2963), .Z(n2962) );
  XOR U3175 ( .A(n2964), .B(n2962), .Z(c[371]) );
  NANDN U3176 ( .A(n2966), .B(n2965), .Z(n2970) );
  OR U3177 ( .A(n2968), .B(n2967), .Z(n2969) );
  NAND U3178 ( .A(n2970), .B(n2969), .Z(n2995) );
  AND U3179 ( .A(b[2]), .B(a[118]), .Z(n2986) );
  AND U3180 ( .A(a[119]), .B(b[1]), .Z(n2984) );
  AND U3181 ( .A(a[117]), .B(b[3]), .Z(n2983) );
  XOR U3182 ( .A(n2984), .B(n2983), .Z(n2985) );
  XOR U3183 ( .A(n2986), .B(n2985), .Z(n2989) );
  NAND U3184 ( .A(b[0]), .B(a[120]), .Z(n2990) );
  XNOR U3185 ( .A(n2989), .B(n2990), .Z(n2991) );
  OR U3186 ( .A(n2972), .B(n2971), .Z(n2976) );
  NANDN U3187 ( .A(n2974), .B(n2973), .Z(n2975) );
  AND U3188 ( .A(n2976), .B(n2975), .Z(n2992) );
  XNOR U3189 ( .A(n2991), .B(n2992), .Z(n2996) );
  XNOR U3190 ( .A(n2995), .B(n2996), .Z(n2997) );
  NANDN U3191 ( .A(n2978), .B(n2977), .Z(n2982) );
  NAND U3192 ( .A(n2980), .B(n2979), .Z(n2981) );
  NAND U3193 ( .A(n2982), .B(n2981), .Z(n2998) );
  XNOR U3194 ( .A(n2997), .B(n2998), .Z(n3001) );
  XOR U3195 ( .A(sreg[372]), .B(n3001), .Z(n3003) );
  XNOR U3196 ( .A(n3002), .B(n3003), .Z(c[372]) );
  AND U3197 ( .A(b[2]), .B(a[119]), .Z(n3018) );
  AND U3198 ( .A(a[120]), .B(b[1]), .Z(n3016) );
  AND U3199 ( .A(a[118]), .B(b[3]), .Z(n3015) );
  XOR U3200 ( .A(n3016), .B(n3015), .Z(n3017) );
  XOR U3201 ( .A(n3018), .B(n3017), .Z(n3021) );
  NAND U3202 ( .A(b[0]), .B(a[121]), .Z(n3022) );
  XOR U3203 ( .A(n3021), .B(n3022), .Z(n3024) );
  OR U3204 ( .A(n2984), .B(n2983), .Z(n2988) );
  NANDN U3205 ( .A(n2986), .B(n2985), .Z(n2987) );
  NAND U3206 ( .A(n2988), .B(n2987), .Z(n3023) );
  XNOR U3207 ( .A(n3024), .B(n3023), .Z(n3009) );
  NANDN U3208 ( .A(n2990), .B(n2989), .Z(n2994) );
  NAND U3209 ( .A(n2992), .B(n2991), .Z(n2993) );
  NAND U3210 ( .A(n2994), .B(n2993), .Z(n3010) );
  XNOR U3211 ( .A(n3009), .B(n3010), .Z(n3011) );
  NANDN U3212 ( .A(n2996), .B(n2995), .Z(n3000) );
  NANDN U3213 ( .A(n2998), .B(n2997), .Z(n2999) );
  NAND U3214 ( .A(n3000), .B(n2999), .Z(n3012) );
  XOR U3215 ( .A(n3011), .B(n3012), .Z(n3008) );
  OR U3216 ( .A(n3001), .B(sreg[372]), .Z(n3005) );
  NAND U3217 ( .A(n3003), .B(n3002), .Z(n3004) );
  AND U3218 ( .A(n3005), .B(n3004), .Z(n3007) );
  XNOR U3219 ( .A(sreg[373]), .B(n3007), .Z(n3006) );
  XNOR U3220 ( .A(n3008), .B(n3006), .Z(c[373]) );
  NANDN U3221 ( .A(n3010), .B(n3009), .Z(n3014) );
  NANDN U3222 ( .A(n3012), .B(n3011), .Z(n3013) );
  NAND U3223 ( .A(n3014), .B(n3013), .Z(n3030) );
  AND U3224 ( .A(b[2]), .B(a[120]), .Z(n3036) );
  AND U3225 ( .A(a[121]), .B(b[1]), .Z(n3034) );
  AND U3226 ( .A(a[119]), .B(b[3]), .Z(n3033) );
  XOR U3227 ( .A(n3034), .B(n3033), .Z(n3035) );
  XOR U3228 ( .A(n3036), .B(n3035), .Z(n3039) );
  NAND U3229 ( .A(b[0]), .B(a[122]), .Z(n3040) );
  XOR U3230 ( .A(n3039), .B(n3040), .Z(n3042) );
  OR U3231 ( .A(n3016), .B(n3015), .Z(n3020) );
  NANDN U3232 ( .A(n3018), .B(n3017), .Z(n3019) );
  NAND U3233 ( .A(n3020), .B(n3019), .Z(n3041) );
  XNOR U3234 ( .A(n3042), .B(n3041), .Z(n3027) );
  NANDN U3235 ( .A(n3022), .B(n3021), .Z(n3026) );
  OR U3236 ( .A(n3024), .B(n3023), .Z(n3025) );
  NAND U3237 ( .A(n3026), .B(n3025), .Z(n3028) );
  XNOR U3238 ( .A(n3027), .B(n3028), .Z(n3029) );
  XNOR U3239 ( .A(n3030), .B(n3029), .Z(n3045) );
  XOR U3240 ( .A(sreg[374]), .B(n3045), .Z(n3047) );
  XNOR U3241 ( .A(n3046), .B(n3047), .Z(c[374]) );
  NANDN U3242 ( .A(n3028), .B(n3027), .Z(n3032) );
  NAND U3243 ( .A(n3030), .B(n3029), .Z(n3031) );
  NAND U3244 ( .A(n3032), .B(n3031), .Z(n3056) );
  AND U3245 ( .A(b[2]), .B(a[121]), .Z(n3062) );
  AND U3246 ( .A(a[122]), .B(b[1]), .Z(n3060) );
  AND U3247 ( .A(a[120]), .B(b[3]), .Z(n3059) );
  XOR U3248 ( .A(n3060), .B(n3059), .Z(n3061) );
  XOR U3249 ( .A(n3062), .B(n3061), .Z(n3065) );
  NAND U3250 ( .A(b[0]), .B(a[123]), .Z(n3066) );
  XOR U3251 ( .A(n3065), .B(n3066), .Z(n3068) );
  OR U3252 ( .A(n3034), .B(n3033), .Z(n3038) );
  NANDN U3253 ( .A(n3036), .B(n3035), .Z(n3037) );
  NAND U3254 ( .A(n3038), .B(n3037), .Z(n3067) );
  XNOR U3255 ( .A(n3068), .B(n3067), .Z(n3053) );
  NANDN U3256 ( .A(n3040), .B(n3039), .Z(n3044) );
  OR U3257 ( .A(n3042), .B(n3041), .Z(n3043) );
  NAND U3258 ( .A(n3044), .B(n3043), .Z(n3054) );
  XNOR U3259 ( .A(n3053), .B(n3054), .Z(n3055) );
  XOR U3260 ( .A(n3056), .B(n3055), .Z(n3052) );
  OR U3261 ( .A(n3045), .B(sreg[374]), .Z(n3049) );
  NAND U3262 ( .A(n3047), .B(n3046), .Z(n3048) );
  AND U3263 ( .A(n3049), .B(n3048), .Z(n3051) );
  XNOR U3264 ( .A(sreg[375]), .B(n3051), .Z(n3050) );
  XOR U3265 ( .A(n3052), .B(n3050), .Z(c[375]) );
  NANDN U3266 ( .A(n3054), .B(n3053), .Z(n3058) );
  NAND U3267 ( .A(n3056), .B(n3055), .Z(n3057) );
  NAND U3268 ( .A(n3058), .B(n3057), .Z(n3079) );
  AND U3269 ( .A(b[2]), .B(a[122]), .Z(n3085) );
  AND U3270 ( .A(a[123]), .B(b[1]), .Z(n3083) );
  AND U3271 ( .A(a[121]), .B(b[3]), .Z(n3082) );
  XOR U3272 ( .A(n3083), .B(n3082), .Z(n3084) );
  XOR U3273 ( .A(n3085), .B(n3084), .Z(n3088) );
  NAND U3274 ( .A(b[0]), .B(a[124]), .Z(n3089) );
  XOR U3275 ( .A(n3088), .B(n3089), .Z(n3091) );
  OR U3276 ( .A(n3060), .B(n3059), .Z(n3064) );
  NANDN U3277 ( .A(n3062), .B(n3061), .Z(n3063) );
  NAND U3278 ( .A(n3064), .B(n3063), .Z(n3090) );
  XNOR U3279 ( .A(n3091), .B(n3090), .Z(n3076) );
  NANDN U3280 ( .A(n3066), .B(n3065), .Z(n3070) );
  OR U3281 ( .A(n3068), .B(n3067), .Z(n3069) );
  NAND U3282 ( .A(n3070), .B(n3069), .Z(n3077) );
  XNOR U3283 ( .A(n3076), .B(n3077), .Z(n3078) );
  XNOR U3284 ( .A(n3079), .B(n3078), .Z(n3071) );
  XOR U3285 ( .A(sreg[376]), .B(n3071), .Z(n3073) );
  XNOR U3286 ( .A(n3072), .B(n3073), .Z(c[376]) );
  OR U3287 ( .A(n3071), .B(sreg[376]), .Z(n3075) );
  NAND U3288 ( .A(n3073), .B(n3072), .Z(n3074) );
  NAND U3289 ( .A(n3075), .B(n3074), .Z(n3114) );
  NANDN U3290 ( .A(n3077), .B(n3076), .Z(n3081) );
  NAND U3291 ( .A(n3079), .B(n3078), .Z(n3080) );
  NAND U3292 ( .A(n3081), .B(n3080), .Z(n3097) );
  AND U3293 ( .A(b[2]), .B(a[123]), .Z(n3103) );
  AND U3294 ( .A(a[124]), .B(b[1]), .Z(n3101) );
  AND U3295 ( .A(a[122]), .B(b[3]), .Z(n3100) );
  XOR U3296 ( .A(n3101), .B(n3100), .Z(n3102) );
  XOR U3297 ( .A(n3103), .B(n3102), .Z(n3106) );
  NAND U3298 ( .A(b[0]), .B(a[125]), .Z(n3107) );
  XOR U3299 ( .A(n3106), .B(n3107), .Z(n3109) );
  OR U3300 ( .A(n3083), .B(n3082), .Z(n3087) );
  NANDN U3301 ( .A(n3085), .B(n3084), .Z(n3086) );
  NAND U3302 ( .A(n3087), .B(n3086), .Z(n3108) );
  XNOR U3303 ( .A(n3109), .B(n3108), .Z(n3094) );
  NANDN U3304 ( .A(n3089), .B(n3088), .Z(n3093) );
  OR U3305 ( .A(n3091), .B(n3090), .Z(n3092) );
  NAND U3306 ( .A(n3093), .B(n3092), .Z(n3095) );
  XNOR U3307 ( .A(n3094), .B(n3095), .Z(n3096) );
  XNOR U3308 ( .A(n3097), .B(n3096), .Z(n3112) );
  XNOR U3309 ( .A(n3112), .B(sreg[377]), .Z(n3113) );
  XOR U3310 ( .A(n3114), .B(n3113), .Z(c[377]) );
  NANDN U3311 ( .A(n3095), .B(n3094), .Z(n3099) );
  NAND U3312 ( .A(n3097), .B(n3096), .Z(n3098) );
  NAND U3313 ( .A(n3099), .B(n3098), .Z(n3120) );
  AND U3314 ( .A(b[2]), .B(a[124]), .Z(n3126) );
  AND U3315 ( .A(a[125]), .B(b[1]), .Z(n3124) );
  AND U3316 ( .A(a[123]), .B(b[3]), .Z(n3123) );
  XOR U3317 ( .A(n3124), .B(n3123), .Z(n3125) );
  XOR U3318 ( .A(n3126), .B(n3125), .Z(n3129) );
  NAND U3319 ( .A(b[0]), .B(a[126]), .Z(n3130) );
  XOR U3320 ( .A(n3129), .B(n3130), .Z(n3132) );
  OR U3321 ( .A(n3101), .B(n3100), .Z(n3105) );
  NANDN U3322 ( .A(n3103), .B(n3102), .Z(n3104) );
  NAND U3323 ( .A(n3105), .B(n3104), .Z(n3131) );
  XNOR U3324 ( .A(n3132), .B(n3131), .Z(n3117) );
  NANDN U3325 ( .A(n3107), .B(n3106), .Z(n3111) );
  OR U3326 ( .A(n3109), .B(n3108), .Z(n3110) );
  NAND U3327 ( .A(n3111), .B(n3110), .Z(n3118) );
  XNOR U3328 ( .A(n3117), .B(n3118), .Z(n3119) );
  XNOR U3329 ( .A(n3120), .B(n3119), .Z(n3135) );
  XOR U3330 ( .A(sreg[378]), .B(n3135), .Z(n3136) );
  NAND U3331 ( .A(n3112), .B(sreg[377]), .Z(n3116) );
  OR U3332 ( .A(n3114), .B(n3113), .Z(n3115) );
  NAND U3333 ( .A(n3116), .B(n3115), .Z(n3137) );
  XOR U3334 ( .A(n3136), .B(n3137), .Z(c[378]) );
  NANDN U3335 ( .A(n3118), .B(n3117), .Z(n3122) );
  NAND U3336 ( .A(n3120), .B(n3119), .Z(n3121) );
  NAND U3337 ( .A(n3122), .B(n3121), .Z(n3146) );
  AND U3338 ( .A(b[2]), .B(a[125]), .Z(n3152) );
  AND U3339 ( .A(a[126]), .B(b[1]), .Z(n3150) );
  AND U3340 ( .A(a[124]), .B(b[3]), .Z(n3149) );
  XOR U3341 ( .A(n3150), .B(n3149), .Z(n3151) );
  XOR U3342 ( .A(n3152), .B(n3151), .Z(n3155) );
  NAND U3343 ( .A(b[0]), .B(a[127]), .Z(n3156) );
  XOR U3344 ( .A(n3155), .B(n3156), .Z(n3158) );
  OR U3345 ( .A(n3124), .B(n3123), .Z(n3128) );
  NANDN U3346 ( .A(n3126), .B(n3125), .Z(n3127) );
  NAND U3347 ( .A(n3128), .B(n3127), .Z(n3157) );
  XNOR U3348 ( .A(n3158), .B(n3157), .Z(n3143) );
  NANDN U3349 ( .A(n3130), .B(n3129), .Z(n3134) );
  OR U3350 ( .A(n3132), .B(n3131), .Z(n3133) );
  NAND U3351 ( .A(n3134), .B(n3133), .Z(n3144) );
  XNOR U3352 ( .A(n3143), .B(n3144), .Z(n3145) );
  XOR U3353 ( .A(n3146), .B(n3145), .Z(n3142) );
  OR U3354 ( .A(n3135), .B(sreg[378]), .Z(n3139) );
  NANDN U3355 ( .A(n3137), .B(n3136), .Z(n3138) );
  AND U3356 ( .A(n3139), .B(n3138), .Z(n3141) );
  XNOR U3357 ( .A(sreg[379]), .B(n3141), .Z(n3140) );
  XOR U3358 ( .A(n3142), .B(n3140), .Z(c[379]) );
  NANDN U3359 ( .A(n3144), .B(n3143), .Z(n3148) );
  NAND U3360 ( .A(n3146), .B(n3145), .Z(n3147) );
  NAND U3361 ( .A(n3148), .B(n3147), .Z(n3164) );
  AND U3362 ( .A(b[2]), .B(a[126]), .Z(n3170) );
  AND U3363 ( .A(a[127]), .B(b[1]), .Z(n3168) );
  AND U3364 ( .A(a[125]), .B(b[3]), .Z(n3167) );
  XOR U3365 ( .A(n3168), .B(n3167), .Z(n3169) );
  XOR U3366 ( .A(n3170), .B(n3169), .Z(n3173) );
  NAND U3367 ( .A(b[0]), .B(a[128]), .Z(n3174) );
  XOR U3368 ( .A(n3173), .B(n3174), .Z(n3176) );
  OR U3369 ( .A(n3150), .B(n3149), .Z(n3154) );
  NANDN U3370 ( .A(n3152), .B(n3151), .Z(n3153) );
  NAND U3371 ( .A(n3154), .B(n3153), .Z(n3175) );
  XNOR U3372 ( .A(n3176), .B(n3175), .Z(n3161) );
  NANDN U3373 ( .A(n3156), .B(n3155), .Z(n3160) );
  OR U3374 ( .A(n3158), .B(n3157), .Z(n3159) );
  NAND U3375 ( .A(n3160), .B(n3159), .Z(n3162) );
  XNOR U3376 ( .A(n3161), .B(n3162), .Z(n3163) );
  XNOR U3377 ( .A(n3164), .B(n3163), .Z(n3179) );
  XNOR U3378 ( .A(n3179), .B(sreg[380]), .Z(n3180) );
  XOR U3379 ( .A(n3181), .B(n3180), .Z(c[380]) );
  NANDN U3380 ( .A(n3162), .B(n3161), .Z(n3166) );
  NAND U3381 ( .A(n3164), .B(n3163), .Z(n3165) );
  NAND U3382 ( .A(n3166), .B(n3165), .Z(n3187) );
  AND U3383 ( .A(b[2]), .B(a[127]), .Z(n3193) );
  AND U3384 ( .A(a[128]), .B(b[1]), .Z(n3191) );
  AND U3385 ( .A(a[126]), .B(b[3]), .Z(n3190) );
  XOR U3386 ( .A(n3191), .B(n3190), .Z(n3192) );
  XOR U3387 ( .A(n3193), .B(n3192), .Z(n3196) );
  NAND U3388 ( .A(b[0]), .B(a[129]), .Z(n3197) );
  XOR U3389 ( .A(n3196), .B(n3197), .Z(n3199) );
  OR U3390 ( .A(n3168), .B(n3167), .Z(n3172) );
  NANDN U3391 ( .A(n3170), .B(n3169), .Z(n3171) );
  NAND U3392 ( .A(n3172), .B(n3171), .Z(n3198) );
  XNOR U3393 ( .A(n3199), .B(n3198), .Z(n3184) );
  NANDN U3394 ( .A(n3174), .B(n3173), .Z(n3178) );
  OR U3395 ( .A(n3176), .B(n3175), .Z(n3177) );
  NAND U3396 ( .A(n3178), .B(n3177), .Z(n3185) );
  XNOR U3397 ( .A(n3184), .B(n3185), .Z(n3186) );
  XNOR U3398 ( .A(n3187), .B(n3186), .Z(n3202) );
  XOR U3399 ( .A(sreg[381]), .B(n3202), .Z(n3203) );
  NAND U3400 ( .A(n3179), .B(sreg[380]), .Z(n3183) );
  OR U3401 ( .A(n3181), .B(n3180), .Z(n3182) );
  NAND U3402 ( .A(n3183), .B(n3182), .Z(n3204) );
  XOR U3403 ( .A(n3203), .B(n3204), .Z(c[381]) );
  NANDN U3404 ( .A(n3185), .B(n3184), .Z(n3189) );
  NAND U3405 ( .A(n3187), .B(n3186), .Z(n3188) );
  NAND U3406 ( .A(n3189), .B(n3188), .Z(n3210) );
  AND U3407 ( .A(b[2]), .B(a[128]), .Z(n3216) );
  AND U3408 ( .A(a[129]), .B(b[1]), .Z(n3214) );
  AND U3409 ( .A(a[127]), .B(b[3]), .Z(n3213) );
  XOR U3410 ( .A(n3214), .B(n3213), .Z(n3215) );
  XOR U3411 ( .A(n3216), .B(n3215), .Z(n3219) );
  NAND U3412 ( .A(b[0]), .B(a[130]), .Z(n3220) );
  XOR U3413 ( .A(n3219), .B(n3220), .Z(n3222) );
  OR U3414 ( .A(n3191), .B(n3190), .Z(n3195) );
  NANDN U3415 ( .A(n3193), .B(n3192), .Z(n3194) );
  NAND U3416 ( .A(n3195), .B(n3194), .Z(n3221) );
  XNOR U3417 ( .A(n3222), .B(n3221), .Z(n3207) );
  NANDN U3418 ( .A(n3197), .B(n3196), .Z(n3201) );
  OR U3419 ( .A(n3199), .B(n3198), .Z(n3200) );
  NAND U3420 ( .A(n3201), .B(n3200), .Z(n3208) );
  XNOR U3421 ( .A(n3207), .B(n3208), .Z(n3209) );
  XNOR U3422 ( .A(n3210), .B(n3209), .Z(n3225) );
  XOR U3423 ( .A(sreg[382]), .B(n3225), .Z(n3226) );
  OR U3424 ( .A(n3202), .B(sreg[381]), .Z(n3206) );
  NANDN U3425 ( .A(n3204), .B(n3203), .Z(n3205) );
  AND U3426 ( .A(n3206), .B(n3205), .Z(n3227) );
  XOR U3427 ( .A(n3226), .B(n3227), .Z(c[382]) );
  NANDN U3428 ( .A(n3208), .B(n3207), .Z(n3212) );
  NAND U3429 ( .A(n3210), .B(n3209), .Z(n3211) );
  NAND U3430 ( .A(n3212), .B(n3211), .Z(n3236) );
  AND U3431 ( .A(b[2]), .B(a[129]), .Z(n3242) );
  AND U3432 ( .A(a[130]), .B(b[1]), .Z(n3240) );
  AND U3433 ( .A(a[128]), .B(b[3]), .Z(n3239) );
  XOR U3434 ( .A(n3240), .B(n3239), .Z(n3241) );
  XOR U3435 ( .A(n3242), .B(n3241), .Z(n3245) );
  NAND U3436 ( .A(b[0]), .B(a[131]), .Z(n3246) );
  XOR U3437 ( .A(n3245), .B(n3246), .Z(n3248) );
  OR U3438 ( .A(n3214), .B(n3213), .Z(n3218) );
  NANDN U3439 ( .A(n3216), .B(n3215), .Z(n3217) );
  NAND U3440 ( .A(n3218), .B(n3217), .Z(n3247) );
  XNOR U3441 ( .A(n3248), .B(n3247), .Z(n3233) );
  NANDN U3442 ( .A(n3220), .B(n3219), .Z(n3224) );
  OR U3443 ( .A(n3222), .B(n3221), .Z(n3223) );
  NAND U3444 ( .A(n3224), .B(n3223), .Z(n3234) );
  XNOR U3445 ( .A(n3233), .B(n3234), .Z(n3235) );
  XOR U3446 ( .A(n3236), .B(n3235), .Z(n3232) );
  OR U3447 ( .A(n3225), .B(sreg[382]), .Z(n3229) );
  NANDN U3448 ( .A(n3227), .B(n3226), .Z(n3228) );
  AND U3449 ( .A(n3229), .B(n3228), .Z(n3231) );
  XNOR U3450 ( .A(sreg[383]), .B(n3231), .Z(n3230) );
  XOR U3451 ( .A(n3232), .B(n3230), .Z(c[383]) );
  NANDN U3452 ( .A(n3234), .B(n3233), .Z(n3238) );
  NAND U3453 ( .A(n3236), .B(n3235), .Z(n3237) );
  NAND U3454 ( .A(n3238), .B(n3237), .Z(n3254) );
  AND U3455 ( .A(b[2]), .B(a[130]), .Z(n3266) );
  AND U3456 ( .A(a[131]), .B(b[1]), .Z(n3264) );
  AND U3457 ( .A(a[129]), .B(b[3]), .Z(n3263) );
  XOR U3458 ( .A(n3264), .B(n3263), .Z(n3265) );
  XOR U3459 ( .A(n3266), .B(n3265), .Z(n3257) );
  NAND U3460 ( .A(b[0]), .B(a[132]), .Z(n3258) );
  XOR U3461 ( .A(n3257), .B(n3258), .Z(n3260) );
  OR U3462 ( .A(n3240), .B(n3239), .Z(n3244) );
  NANDN U3463 ( .A(n3242), .B(n3241), .Z(n3243) );
  NAND U3464 ( .A(n3244), .B(n3243), .Z(n3259) );
  XNOR U3465 ( .A(n3260), .B(n3259), .Z(n3251) );
  NANDN U3466 ( .A(n3246), .B(n3245), .Z(n3250) );
  OR U3467 ( .A(n3248), .B(n3247), .Z(n3249) );
  NAND U3468 ( .A(n3250), .B(n3249), .Z(n3252) );
  XNOR U3469 ( .A(n3251), .B(n3252), .Z(n3253) );
  XOR U3470 ( .A(n3254), .B(n3253), .Z(n3269) );
  XNOR U3471 ( .A(sreg[384]), .B(n3269), .Z(n3270) );
  XNOR U3472 ( .A(n3271), .B(n3270), .Z(c[384]) );
  NANDN U3473 ( .A(n3252), .B(n3251), .Z(n3256) );
  NAND U3474 ( .A(n3254), .B(n3253), .Z(n3255) );
  NAND U3475 ( .A(n3256), .B(n3255), .Z(n3290) );
  NANDN U3476 ( .A(n3258), .B(n3257), .Z(n3262) );
  OR U3477 ( .A(n3260), .B(n3259), .Z(n3261) );
  NAND U3478 ( .A(n3262), .B(n3261), .Z(n3287) );
  AND U3479 ( .A(b[2]), .B(a[131]), .Z(n3278) );
  AND U3480 ( .A(a[132]), .B(b[1]), .Z(n3276) );
  AND U3481 ( .A(a[130]), .B(b[3]), .Z(n3275) );
  XOR U3482 ( .A(n3276), .B(n3275), .Z(n3277) );
  XOR U3483 ( .A(n3278), .B(n3277), .Z(n3281) );
  NAND U3484 ( .A(b[0]), .B(a[133]), .Z(n3282) );
  XNOR U3485 ( .A(n3281), .B(n3282), .Z(n3283) );
  OR U3486 ( .A(n3264), .B(n3263), .Z(n3268) );
  NANDN U3487 ( .A(n3266), .B(n3265), .Z(n3267) );
  AND U3488 ( .A(n3268), .B(n3267), .Z(n3284) );
  XNOR U3489 ( .A(n3283), .B(n3284), .Z(n3288) );
  XNOR U3490 ( .A(n3287), .B(n3288), .Z(n3289) );
  XOR U3491 ( .A(n3290), .B(n3289), .Z(n3294) );
  NANDN U3492 ( .A(sreg[384]), .B(n3269), .Z(n3273) );
  NAND U3493 ( .A(n3271), .B(n3270), .Z(n3272) );
  AND U3494 ( .A(n3273), .B(n3272), .Z(n3293) );
  XOR U3495 ( .A(sreg[385]), .B(n3293), .Z(n3274) );
  XNOR U3496 ( .A(n3294), .B(n3274), .Z(c[385]) );
  AND U3497 ( .A(b[2]), .B(a[132]), .Z(n3305) );
  AND U3498 ( .A(a[133]), .B(b[1]), .Z(n3303) );
  AND U3499 ( .A(a[131]), .B(b[3]), .Z(n3302) );
  XOR U3500 ( .A(n3303), .B(n3302), .Z(n3304) );
  XOR U3501 ( .A(n3305), .B(n3304), .Z(n3308) );
  NAND U3502 ( .A(b[0]), .B(a[134]), .Z(n3309) );
  XOR U3503 ( .A(n3308), .B(n3309), .Z(n3311) );
  OR U3504 ( .A(n3276), .B(n3275), .Z(n3280) );
  NANDN U3505 ( .A(n3278), .B(n3277), .Z(n3279) );
  NAND U3506 ( .A(n3280), .B(n3279), .Z(n3310) );
  XNOR U3507 ( .A(n3311), .B(n3310), .Z(n3296) );
  NANDN U3508 ( .A(n3282), .B(n3281), .Z(n3286) );
  NAND U3509 ( .A(n3284), .B(n3283), .Z(n3285) );
  NAND U3510 ( .A(n3286), .B(n3285), .Z(n3297) );
  XNOR U3511 ( .A(n3296), .B(n3297), .Z(n3298) );
  NANDN U3512 ( .A(n3288), .B(n3287), .Z(n3292) );
  NANDN U3513 ( .A(n3290), .B(n3289), .Z(n3291) );
  NAND U3514 ( .A(n3292), .B(n3291), .Z(n3299) );
  XOR U3515 ( .A(n3298), .B(n3299), .Z(n3315) );
  XOR U3516 ( .A(sreg[386]), .B(n3314), .Z(n3295) );
  XNOR U3517 ( .A(n3315), .B(n3295), .Z(c[386]) );
  NANDN U3518 ( .A(n3297), .B(n3296), .Z(n3301) );
  NANDN U3519 ( .A(n3299), .B(n3298), .Z(n3300) );
  NAND U3520 ( .A(n3301), .B(n3300), .Z(n3334) );
  AND U3521 ( .A(b[2]), .B(a[133]), .Z(n3328) );
  AND U3522 ( .A(a[134]), .B(b[1]), .Z(n3326) );
  AND U3523 ( .A(a[132]), .B(b[3]), .Z(n3325) );
  XOR U3524 ( .A(n3326), .B(n3325), .Z(n3327) );
  XOR U3525 ( .A(n3328), .B(n3327), .Z(n3319) );
  NAND U3526 ( .A(b[0]), .B(a[135]), .Z(n3320) );
  XOR U3527 ( .A(n3319), .B(n3320), .Z(n3322) );
  OR U3528 ( .A(n3303), .B(n3302), .Z(n3307) );
  NANDN U3529 ( .A(n3305), .B(n3304), .Z(n3306) );
  NAND U3530 ( .A(n3307), .B(n3306), .Z(n3321) );
  XNOR U3531 ( .A(n3322), .B(n3321), .Z(n3331) );
  NANDN U3532 ( .A(n3309), .B(n3308), .Z(n3313) );
  OR U3533 ( .A(n3311), .B(n3310), .Z(n3312) );
  NAND U3534 ( .A(n3313), .B(n3312), .Z(n3332) );
  XNOR U3535 ( .A(n3331), .B(n3332), .Z(n3333) );
  XOR U3536 ( .A(n3334), .B(n3333), .Z(n3318) );
  XNOR U3537 ( .A(sreg[387]), .B(n3317), .Z(n3316) );
  XOR U3538 ( .A(n3318), .B(n3316), .Z(c[387]) );
  NANDN U3539 ( .A(n3320), .B(n3319), .Z(n3324) );
  OR U3540 ( .A(n3322), .B(n3321), .Z(n3323) );
  NAND U3541 ( .A(n3324), .B(n3323), .Z(n3349) );
  AND U3542 ( .A(b[2]), .B(a[134]), .Z(n3340) );
  AND U3543 ( .A(a[135]), .B(b[1]), .Z(n3338) );
  AND U3544 ( .A(a[133]), .B(b[3]), .Z(n3337) );
  XOR U3545 ( .A(n3338), .B(n3337), .Z(n3339) );
  XOR U3546 ( .A(n3340), .B(n3339), .Z(n3343) );
  NAND U3547 ( .A(b[0]), .B(a[136]), .Z(n3344) );
  XNOR U3548 ( .A(n3343), .B(n3344), .Z(n3345) );
  OR U3549 ( .A(n3326), .B(n3325), .Z(n3330) );
  NANDN U3550 ( .A(n3328), .B(n3327), .Z(n3329) );
  AND U3551 ( .A(n3330), .B(n3329), .Z(n3346) );
  XNOR U3552 ( .A(n3345), .B(n3346), .Z(n3350) );
  XNOR U3553 ( .A(n3349), .B(n3350), .Z(n3351) );
  NANDN U3554 ( .A(n3332), .B(n3331), .Z(n3336) );
  NAND U3555 ( .A(n3334), .B(n3333), .Z(n3335) );
  AND U3556 ( .A(n3336), .B(n3335), .Z(n3352) );
  XOR U3557 ( .A(n3351), .B(n3352), .Z(n3355) );
  XNOR U3558 ( .A(sreg[388]), .B(n3355), .Z(n3356) );
  XOR U3559 ( .A(n3357), .B(n3356), .Z(c[388]) );
  AND U3560 ( .A(b[2]), .B(a[135]), .Z(n3369) );
  AND U3561 ( .A(a[136]), .B(b[1]), .Z(n3367) );
  AND U3562 ( .A(a[134]), .B(b[3]), .Z(n3366) );
  XOR U3563 ( .A(n3367), .B(n3366), .Z(n3368) );
  XOR U3564 ( .A(n3369), .B(n3368), .Z(n3372) );
  NAND U3565 ( .A(b[0]), .B(a[137]), .Z(n3373) );
  XOR U3566 ( .A(n3372), .B(n3373), .Z(n3375) );
  OR U3567 ( .A(n3338), .B(n3337), .Z(n3342) );
  NANDN U3568 ( .A(n3340), .B(n3339), .Z(n3341) );
  NAND U3569 ( .A(n3342), .B(n3341), .Z(n3374) );
  XNOR U3570 ( .A(n3375), .B(n3374), .Z(n3360) );
  NANDN U3571 ( .A(n3344), .B(n3343), .Z(n3348) );
  NAND U3572 ( .A(n3346), .B(n3345), .Z(n3347) );
  NAND U3573 ( .A(n3348), .B(n3347), .Z(n3361) );
  XNOR U3574 ( .A(n3360), .B(n3361), .Z(n3362) );
  NANDN U3575 ( .A(n3350), .B(n3349), .Z(n3354) );
  NAND U3576 ( .A(n3352), .B(n3351), .Z(n3353) );
  NAND U3577 ( .A(n3354), .B(n3353), .Z(n3363) );
  XOR U3578 ( .A(n3362), .B(n3363), .Z(n3378) );
  XNOR U3579 ( .A(n3378), .B(sreg[389]), .Z(n3380) );
  NAND U3580 ( .A(sreg[388]), .B(n3355), .Z(n3359) );
  OR U3581 ( .A(n3357), .B(n3356), .Z(n3358) );
  AND U3582 ( .A(n3359), .B(n3358), .Z(n3379) );
  XOR U3583 ( .A(n3380), .B(n3379), .Z(c[389]) );
  NANDN U3584 ( .A(n3361), .B(n3360), .Z(n3365) );
  NANDN U3585 ( .A(n3363), .B(n3362), .Z(n3364) );
  NAND U3586 ( .A(n3365), .B(n3364), .Z(n3387) );
  AND U3587 ( .A(b[2]), .B(a[136]), .Z(n3393) );
  AND U3588 ( .A(a[137]), .B(b[1]), .Z(n3391) );
  AND U3589 ( .A(a[135]), .B(b[3]), .Z(n3390) );
  XOR U3590 ( .A(n3391), .B(n3390), .Z(n3392) );
  XOR U3591 ( .A(n3393), .B(n3392), .Z(n3396) );
  NAND U3592 ( .A(b[0]), .B(a[138]), .Z(n3397) );
  XOR U3593 ( .A(n3396), .B(n3397), .Z(n3399) );
  OR U3594 ( .A(n3367), .B(n3366), .Z(n3371) );
  NANDN U3595 ( .A(n3369), .B(n3368), .Z(n3370) );
  NAND U3596 ( .A(n3371), .B(n3370), .Z(n3398) );
  XNOR U3597 ( .A(n3399), .B(n3398), .Z(n3384) );
  NANDN U3598 ( .A(n3373), .B(n3372), .Z(n3377) );
  OR U3599 ( .A(n3375), .B(n3374), .Z(n3376) );
  NAND U3600 ( .A(n3377), .B(n3376), .Z(n3385) );
  XNOR U3601 ( .A(n3384), .B(n3385), .Z(n3386) );
  XOR U3602 ( .A(n3387), .B(n3386), .Z(n3403) );
  NAND U3603 ( .A(n3378), .B(sreg[389]), .Z(n3382) );
  OR U3604 ( .A(n3380), .B(n3379), .Z(n3381) );
  NAND U3605 ( .A(n3382), .B(n3381), .Z(n3402) );
  XNOR U3606 ( .A(sreg[390]), .B(n3402), .Z(n3383) );
  XOR U3607 ( .A(n3403), .B(n3383), .Z(c[390]) );
  NANDN U3608 ( .A(n3385), .B(n3384), .Z(n3389) );
  NAND U3609 ( .A(n3387), .B(n3386), .Z(n3388) );
  NAND U3610 ( .A(n3389), .B(n3388), .Z(n3410) );
  AND U3611 ( .A(b[2]), .B(a[137]), .Z(n3416) );
  AND U3612 ( .A(a[138]), .B(b[1]), .Z(n3414) );
  AND U3613 ( .A(a[136]), .B(b[3]), .Z(n3413) );
  XOR U3614 ( .A(n3414), .B(n3413), .Z(n3415) );
  XOR U3615 ( .A(n3416), .B(n3415), .Z(n3419) );
  NAND U3616 ( .A(b[0]), .B(a[139]), .Z(n3420) );
  XOR U3617 ( .A(n3419), .B(n3420), .Z(n3422) );
  OR U3618 ( .A(n3391), .B(n3390), .Z(n3395) );
  NANDN U3619 ( .A(n3393), .B(n3392), .Z(n3394) );
  NAND U3620 ( .A(n3395), .B(n3394), .Z(n3421) );
  XNOR U3621 ( .A(n3422), .B(n3421), .Z(n3407) );
  NANDN U3622 ( .A(n3397), .B(n3396), .Z(n3401) );
  OR U3623 ( .A(n3399), .B(n3398), .Z(n3400) );
  NAND U3624 ( .A(n3401), .B(n3400), .Z(n3408) );
  XNOR U3625 ( .A(n3407), .B(n3408), .Z(n3409) );
  XNOR U3626 ( .A(n3410), .B(n3409), .Z(n3406) );
  XOR U3627 ( .A(n3405), .B(sreg[391]), .Z(n3404) );
  XOR U3628 ( .A(n3406), .B(n3404), .Z(c[391]) );
  NANDN U3629 ( .A(n3408), .B(n3407), .Z(n3412) );
  NAND U3630 ( .A(n3410), .B(n3409), .Z(n3411) );
  NAND U3631 ( .A(n3412), .B(n3411), .Z(n3433) );
  AND U3632 ( .A(b[2]), .B(a[138]), .Z(n3439) );
  AND U3633 ( .A(a[139]), .B(b[1]), .Z(n3437) );
  AND U3634 ( .A(a[137]), .B(b[3]), .Z(n3436) );
  XOR U3635 ( .A(n3437), .B(n3436), .Z(n3438) );
  XOR U3636 ( .A(n3439), .B(n3438), .Z(n3442) );
  NAND U3637 ( .A(b[0]), .B(a[140]), .Z(n3443) );
  XOR U3638 ( .A(n3442), .B(n3443), .Z(n3445) );
  OR U3639 ( .A(n3414), .B(n3413), .Z(n3418) );
  NANDN U3640 ( .A(n3416), .B(n3415), .Z(n3417) );
  NAND U3641 ( .A(n3418), .B(n3417), .Z(n3444) );
  XNOR U3642 ( .A(n3445), .B(n3444), .Z(n3430) );
  NANDN U3643 ( .A(n3420), .B(n3419), .Z(n3424) );
  OR U3644 ( .A(n3422), .B(n3421), .Z(n3423) );
  NAND U3645 ( .A(n3424), .B(n3423), .Z(n3431) );
  XNOR U3646 ( .A(n3430), .B(n3431), .Z(n3432) );
  XNOR U3647 ( .A(n3433), .B(n3432), .Z(n3425) );
  XOR U3648 ( .A(sreg[392]), .B(n3425), .Z(n3426) );
  XOR U3649 ( .A(n3427), .B(n3426), .Z(c[392]) );
  OR U3650 ( .A(n3425), .B(sreg[392]), .Z(n3429) );
  NANDN U3651 ( .A(n3427), .B(n3426), .Z(n3428) );
  AND U3652 ( .A(n3429), .B(n3428), .Z(n3449) );
  NANDN U3653 ( .A(n3431), .B(n3430), .Z(n3435) );
  NAND U3654 ( .A(n3433), .B(n3432), .Z(n3434) );
  NAND U3655 ( .A(n3435), .B(n3434), .Z(n3454) );
  AND U3656 ( .A(b[2]), .B(a[139]), .Z(n3460) );
  AND U3657 ( .A(a[140]), .B(b[1]), .Z(n3458) );
  AND U3658 ( .A(a[138]), .B(b[3]), .Z(n3457) );
  XOR U3659 ( .A(n3458), .B(n3457), .Z(n3459) );
  XOR U3660 ( .A(n3460), .B(n3459), .Z(n3463) );
  NAND U3661 ( .A(b[0]), .B(a[141]), .Z(n3464) );
  XOR U3662 ( .A(n3463), .B(n3464), .Z(n3466) );
  OR U3663 ( .A(n3437), .B(n3436), .Z(n3441) );
  NANDN U3664 ( .A(n3439), .B(n3438), .Z(n3440) );
  NAND U3665 ( .A(n3441), .B(n3440), .Z(n3465) );
  XNOR U3666 ( .A(n3466), .B(n3465), .Z(n3451) );
  NANDN U3667 ( .A(n3443), .B(n3442), .Z(n3447) );
  OR U3668 ( .A(n3445), .B(n3444), .Z(n3446) );
  NAND U3669 ( .A(n3447), .B(n3446), .Z(n3452) );
  XNOR U3670 ( .A(n3451), .B(n3452), .Z(n3453) );
  XNOR U3671 ( .A(n3454), .B(n3453), .Z(n3450) );
  XOR U3672 ( .A(sreg[393]), .B(n3450), .Z(n3448) );
  XOR U3673 ( .A(n3449), .B(n3448), .Z(c[393]) );
  NANDN U3674 ( .A(n3452), .B(n3451), .Z(n3456) );
  NAND U3675 ( .A(n3454), .B(n3453), .Z(n3455) );
  NAND U3676 ( .A(n3456), .B(n3455), .Z(n3472) );
  AND U3677 ( .A(b[2]), .B(a[140]), .Z(n3478) );
  AND U3678 ( .A(a[141]), .B(b[1]), .Z(n3476) );
  AND U3679 ( .A(a[139]), .B(b[3]), .Z(n3475) );
  XOR U3680 ( .A(n3476), .B(n3475), .Z(n3477) );
  XOR U3681 ( .A(n3478), .B(n3477), .Z(n3481) );
  NAND U3682 ( .A(b[0]), .B(a[142]), .Z(n3482) );
  XOR U3683 ( .A(n3481), .B(n3482), .Z(n3484) );
  OR U3684 ( .A(n3458), .B(n3457), .Z(n3462) );
  NANDN U3685 ( .A(n3460), .B(n3459), .Z(n3461) );
  NAND U3686 ( .A(n3462), .B(n3461), .Z(n3483) );
  XNOR U3687 ( .A(n3484), .B(n3483), .Z(n3469) );
  NANDN U3688 ( .A(n3464), .B(n3463), .Z(n3468) );
  OR U3689 ( .A(n3466), .B(n3465), .Z(n3467) );
  NAND U3690 ( .A(n3468), .B(n3467), .Z(n3470) );
  XNOR U3691 ( .A(n3469), .B(n3470), .Z(n3471) );
  XOR U3692 ( .A(n3472), .B(n3471), .Z(n3487) );
  XOR U3693 ( .A(sreg[394]), .B(n3487), .Z(n3489) );
  XNOR U3694 ( .A(n3488), .B(n3489), .Z(c[394]) );
  NANDN U3695 ( .A(n3470), .B(n3469), .Z(n3474) );
  NAND U3696 ( .A(n3472), .B(n3471), .Z(n3473) );
  NAND U3697 ( .A(n3474), .B(n3473), .Z(n3495) );
  AND U3698 ( .A(b[2]), .B(a[141]), .Z(n3501) );
  AND U3699 ( .A(a[142]), .B(b[1]), .Z(n3499) );
  AND U3700 ( .A(a[140]), .B(b[3]), .Z(n3498) );
  XOR U3701 ( .A(n3499), .B(n3498), .Z(n3500) );
  XOR U3702 ( .A(n3501), .B(n3500), .Z(n3504) );
  NAND U3703 ( .A(b[0]), .B(a[143]), .Z(n3505) );
  XOR U3704 ( .A(n3504), .B(n3505), .Z(n3507) );
  OR U3705 ( .A(n3476), .B(n3475), .Z(n3480) );
  NANDN U3706 ( .A(n3478), .B(n3477), .Z(n3479) );
  NAND U3707 ( .A(n3480), .B(n3479), .Z(n3506) );
  XNOR U3708 ( .A(n3507), .B(n3506), .Z(n3492) );
  NANDN U3709 ( .A(n3482), .B(n3481), .Z(n3486) );
  OR U3710 ( .A(n3484), .B(n3483), .Z(n3485) );
  NAND U3711 ( .A(n3486), .B(n3485), .Z(n3493) );
  XNOR U3712 ( .A(n3492), .B(n3493), .Z(n3494) );
  XNOR U3713 ( .A(n3495), .B(n3494), .Z(n3510) );
  XOR U3714 ( .A(sreg[395]), .B(n3510), .Z(n3511) );
  NANDN U3715 ( .A(n3487), .B(sreg[394]), .Z(n3491) );
  NANDN U3716 ( .A(n3489), .B(n3488), .Z(n3490) );
  NAND U3717 ( .A(n3491), .B(n3490), .Z(n3512) );
  XOR U3718 ( .A(n3511), .B(n3512), .Z(c[395]) );
  NANDN U3719 ( .A(n3493), .B(n3492), .Z(n3497) );
  NAND U3720 ( .A(n3495), .B(n3494), .Z(n3496) );
  NAND U3721 ( .A(n3497), .B(n3496), .Z(n3521) );
  AND U3722 ( .A(b[2]), .B(a[142]), .Z(n3527) );
  AND U3723 ( .A(a[143]), .B(b[1]), .Z(n3525) );
  AND U3724 ( .A(a[141]), .B(b[3]), .Z(n3524) );
  XOR U3725 ( .A(n3525), .B(n3524), .Z(n3526) );
  XOR U3726 ( .A(n3527), .B(n3526), .Z(n3530) );
  NAND U3727 ( .A(b[0]), .B(a[144]), .Z(n3531) );
  XOR U3728 ( .A(n3530), .B(n3531), .Z(n3533) );
  OR U3729 ( .A(n3499), .B(n3498), .Z(n3503) );
  NANDN U3730 ( .A(n3501), .B(n3500), .Z(n3502) );
  NAND U3731 ( .A(n3503), .B(n3502), .Z(n3532) );
  XNOR U3732 ( .A(n3533), .B(n3532), .Z(n3518) );
  NANDN U3733 ( .A(n3505), .B(n3504), .Z(n3509) );
  OR U3734 ( .A(n3507), .B(n3506), .Z(n3508) );
  NAND U3735 ( .A(n3509), .B(n3508), .Z(n3519) );
  XNOR U3736 ( .A(n3518), .B(n3519), .Z(n3520) );
  XOR U3737 ( .A(n3521), .B(n3520), .Z(n3517) );
  OR U3738 ( .A(n3510), .B(sreg[395]), .Z(n3514) );
  NANDN U3739 ( .A(n3512), .B(n3511), .Z(n3513) );
  AND U3740 ( .A(n3514), .B(n3513), .Z(n3516) );
  XNOR U3741 ( .A(sreg[396]), .B(n3516), .Z(n3515) );
  XOR U3742 ( .A(n3517), .B(n3515), .Z(c[396]) );
  NANDN U3743 ( .A(n3519), .B(n3518), .Z(n3523) );
  NAND U3744 ( .A(n3521), .B(n3520), .Z(n3522) );
  NAND U3745 ( .A(n3523), .B(n3522), .Z(n3544) );
  AND U3746 ( .A(b[2]), .B(a[143]), .Z(n3550) );
  AND U3747 ( .A(a[144]), .B(b[1]), .Z(n3548) );
  AND U3748 ( .A(a[142]), .B(b[3]), .Z(n3547) );
  XOR U3749 ( .A(n3548), .B(n3547), .Z(n3549) );
  XOR U3750 ( .A(n3550), .B(n3549), .Z(n3553) );
  NAND U3751 ( .A(b[0]), .B(a[145]), .Z(n3554) );
  XOR U3752 ( .A(n3553), .B(n3554), .Z(n3556) );
  OR U3753 ( .A(n3525), .B(n3524), .Z(n3529) );
  NANDN U3754 ( .A(n3527), .B(n3526), .Z(n3528) );
  NAND U3755 ( .A(n3529), .B(n3528), .Z(n3555) );
  XNOR U3756 ( .A(n3556), .B(n3555), .Z(n3541) );
  NANDN U3757 ( .A(n3531), .B(n3530), .Z(n3535) );
  OR U3758 ( .A(n3533), .B(n3532), .Z(n3534) );
  NAND U3759 ( .A(n3535), .B(n3534), .Z(n3542) );
  XNOR U3760 ( .A(n3541), .B(n3542), .Z(n3543) );
  XNOR U3761 ( .A(n3544), .B(n3543), .Z(n3536) );
  XNOR U3762 ( .A(n3536), .B(sreg[397]), .Z(n3537) );
  XOR U3763 ( .A(n3538), .B(n3537), .Z(c[397]) );
  NAND U3764 ( .A(n3536), .B(sreg[397]), .Z(n3540) );
  OR U3765 ( .A(n3538), .B(n3537), .Z(n3539) );
  NAND U3766 ( .A(n3540), .B(n3539), .Z(n3561) );
  NANDN U3767 ( .A(n3542), .B(n3541), .Z(n3546) );
  NAND U3768 ( .A(n3544), .B(n3543), .Z(n3545) );
  NAND U3769 ( .A(n3546), .B(n3545), .Z(n3567) );
  AND U3770 ( .A(b[2]), .B(a[144]), .Z(n3573) );
  AND U3771 ( .A(a[145]), .B(b[1]), .Z(n3571) );
  AND U3772 ( .A(a[143]), .B(b[3]), .Z(n3570) );
  XOR U3773 ( .A(n3571), .B(n3570), .Z(n3572) );
  XOR U3774 ( .A(n3573), .B(n3572), .Z(n3576) );
  NAND U3775 ( .A(b[0]), .B(a[146]), .Z(n3577) );
  XOR U3776 ( .A(n3576), .B(n3577), .Z(n3579) );
  OR U3777 ( .A(n3548), .B(n3547), .Z(n3552) );
  NANDN U3778 ( .A(n3550), .B(n3549), .Z(n3551) );
  NAND U3779 ( .A(n3552), .B(n3551), .Z(n3578) );
  XNOR U3780 ( .A(n3579), .B(n3578), .Z(n3564) );
  NANDN U3781 ( .A(n3554), .B(n3553), .Z(n3558) );
  OR U3782 ( .A(n3556), .B(n3555), .Z(n3557) );
  NAND U3783 ( .A(n3558), .B(n3557), .Z(n3565) );
  XNOR U3784 ( .A(n3564), .B(n3565), .Z(n3566) );
  XNOR U3785 ( .A(n3567), .B(n3566), .Z(n3559) );
  XOR U3786 ( .A(sreg[398]), .B(n3559), .Z(n3560) );
  XOR U3787 ( .A(n3561), .B(n3560), .Z(c[398]) );
  OR U3788 ( .A(n3559), .B(sreg[398]), .Z(n3563) );
  NANDN U3789 ( .A(n3561), .B(n3560), .Z(n3562) );
  AND U3790 ( .A(n3563), .B(n3562), .Z(n3583) );
  NANDN U3791 ( .A(n3565), .B(n3564), .Z(n3569) );
  NAND U3792 ( .A(n3567), .B(n3566), .Z(n3568) );
  NAND U3793 ( .A(n3569), .B(n3568), .Z(n3588) );
  AND U3794 ( .A(b[2]), .B(a[145]), .Z(n3594) );
  AND U3795 ( .A(a[146]), .B(b[1]), .Z(n3592) );
  AND U3796 ( .A(a[144]), .B(b[3]), .Z(n3591) );
  XOR U3797 ( .A(n3592), .B(n3591), .Z(n3593) );
  XOR U3798 ( .A(n3594), .B(n3593), .Z(n3597) );
  NAND U3799 ( .A(b[0]), .B(a[147]), .Z(n3598) );
  XOR U3800 ( .A(n3597), .B(n3598), .Z(n3600) );
  OR U3801 ( .A(n3571), .B(n3570), .Z(n3575) );
  NANDN U3802 ( .A(n3573), .B(n3572), .Z(n3574) );
  NAND U3803 ( .A(n3575), .B(n3574), .Z(n3599) );
  XNOR U3804 ( .A(n3600), .B(n3599), .Z(n3585) );
  NANDN U3805 ( .A(n3577), .B(n3576), .Z(n3581) );
  OR U3806 ( .A(n3579), .B(n3578), .Z(n3580) );
  NAND U3807 ( .A(n3581), .B(n3580), .Z(n3586) );
  XNOR U3808 ( .A(n3585), .B(n3586), .Z(n3587) );
  XNOR U3809 ( .A(n3588), .B(n3587), .Z(n3584) );
  XOR U3810 ( .A(sreg[399]), .B(n3584), .Z(n3582) );
  XOR U3811 ( .A(n3583), .B(n3582), .Z(c[399]) );
  NANDN U3812 ( .A(n3586), .B(n3585), .Z(n3590) );
  NAND U3813 ( .A(n3588), .B(n3587), .Z(n3589) );
  NAND U3814 ( .A(n3590), .B(n3589), .Z(n3606) );
  AND U3815 ( .A(b[2]), .B(a[146]), .Z(n3618) );
  AND U3816 ( .A(a[147]), .B(b[1]), .Z(n3616) );
  AND U3817 ( .A(a[145]), .B(b[3]), .Z(n3615) );
  XOR U3818 ( .A(n3616), .B(n3615), .Z(n3617) );
  XOR U3819 ( .A(n3618), .B(n3617), .Z(n3609) );
  NAND U3820 ( .A(b[0]), .B(a[148]), .Z(n3610) );
  XOR U3821 ( .A(n3609), .B(n3610), .Z(n3612) );
  OR U3822 ( .A(n3592), .B(n3591), .Z(n3596) );
  NANDN U3823 ( .A(n3594), .B(n3593), .Z(n3595) );
  NAND U3824 ( .A(n3596), .B(n3595), .Z(n3611) );
  XNOR U3825 ( .A(n3612), .B(n3611), .Z(n3603) );
  NANDN U3826 ( .A(n3598), .B(n3597), .Z(n3602) );
  OR U3827 ( .A(n3600), .B(n3599), .Z(n3601) );
  NAND U3828 ( .A(n3602), .B(n3601), .Z(n3604) );
  XNOR U3829 ( .A(n3603), .B(n3604), .Z(n3605) );
  XNOR U3830 ( .A(n3606), .B(n3605), .Z(n3621) );
  XNOR U3831 ( .A(n3621), .B(sreg[400]), .Z(n3623) );
  XNOR U3832 ( .A(n3622), .B(n3623), .Z(c[400]) );
  NANDN U3833 ( .A(n3604), .B(n3603), .Z(n3608) );
  NAND U3834 ( .A(n3606), .B(n3605), .Z(n3607) );
  NAND U3835 ( .A(n3608), .B(n3607), .Z(n3641) );
  NANDN U3836 ( .A(n3610), .B(n3609), .Z(n3614) );
  OR U3837 ( .A(n3612), .B(n3611), .Z(n3613) );
  NAND U3838 ( .A(n3614), .B(n3613), .Z(n3638) );
  AND U3839 ( .A(b[2]), .B(a[147]), .Z(n3629) );
  AND U3840 ( .A(a[148]), .B(b[1]), .Z(n3627) );
  AND U3841 ( .A(a[146]), .B(b[3]), .Z(n3626) );
  XOR U3842 ( .A(n3627), .B(n3626), .Z(n3628) );
  XOR U3843 ( .A(n3629), .B(n3628), .Z(n3632) );
  NAND U3844 ( .A(b[0]), .B(a[149]), .Z(n3633) );
  XNOR U3845 ( .A(n3632), .B(n3633), .Z(n3634) );
  OR U3846 ( .A(n3616), .B(n3615), .Z(n3620) );
  NANDN U3847 ( .A(n3618), .B(n3617), .Z(n3619) );
  AND U3848 ( .A(n3620), .B(n3619), .Z(n3635) );
  XNOR U3849 ( .A(n3634), .B(n3635), .Z(n3639) );
  XNOR U3850 ( .A(n3638), .B(n3639), .Z(n3640) );
  XNOR U3851 ( .A(n3641), .B(n3640), .Z(n3644) );
  XOR U3852 ( .A(sreg[401]), .B(n3644), .Z(n3645) );
  NAND U3853 ( .A(n3621), .B(sreg[400]), .Z(n3625) );
  NANDN U3854 ( .A(n3623), .B(n3622), .Z(n3624) );
  NAND U3855 ( .A(n3625), .B(n3624), .Z(n3646) );
  XOR U3856 ( .A(n3645), .B(n3646), .Z(c[401]) );
  AND U3857 ( .A(b[2]), .B(a[148]), .Z(n3661) );
  AND U3858 ( .A(a[149]), .B(b[1]), .Z(n3659) );
  AND U3859 ( .A(a[147]), .B(b[3]), .Z(n3658) );
  XOR U3860 ( .A(n3659), .B(n3658), .Z(n3660) );
  XOR U3861 ( .A(n3661), .B(n3660), .Z(n3664) );
  NAND U3862 ( .A(b[0]), .B(a[150]), .Z(n3665) );
  XOR U3863 ( .A(n3664), .B(n3665), .Z(n3667) );
  OR U3864 ( .A(n3627), .B(n3626), .Z(n3631) );
  NANDN U3865 ( .A(n3629), .B(n3628), .Z(n3630) );
  NAND U3866 ( .A(n3631), .B(n3630), .Z(n3666) );
  XNOR U3867 ( .A(n3667), .B(n3666), .Z(n3652) );
  NANDN U3868 ( .A(n3633), .B(n3632), .Z(n3637) );
  NAND U3869 ( .A(n3635), .B(n3634), .Z(n3636) );
  NAND U3870 ( .A(n3637), .B(n3636), .Z(n3653) );
  XNOR U3871 ( .A(n3652), .B(n3653), .Z(n3654) );
  NANDN U3872 ( .A(n3639), .B(n3638), .Z(n3643) );
  NANDN U3873 ( .A(n3641), .B(n3640), .Z(n3642) );
  NAND U3874 ( .A(n3643), .B(n3642), .Z(n3655) );
  XOR U3875 ( .A(n3654), .B(n3655), .Z(n3651) );
  OR U3876 ( .A(n3644), .B(sreg[401]), .Z(n3648) );
  NANDN U3877 ( .A(n3646), .B(n3645), .Z(n3647) );
  AND U3878 ( .A(n3648), .B(n3647), .Z(n3650) );
  XNOR U3879 ( .A(sreg[402]), .B(n3650), .Z(n3649) );
  XNOR U3880 ( .A(n3651), .B(n3649), .Z(c[402]) );
  NANDN U3881 ( .A(n3653), .B(n3652), .Z(n3657) );
  NANDN U3882 ( .A(n3655), .B(n3654), .Z(n3656) );
  NAND U3883 ( .A(n3657), .B(n3656), .Z(n3685) );
  AND U3884 ( .A(b[2]), .B(a[149]), .Z(n3679) );
  AND U3885 ( .A(a[150]), .B(b[1]), .Z(n3677) );
  AND U3886 ( .A(a[148]), .B(b[3]), .Z(n3676) );
  XOR U3887 ( .A(n3677), .B(n3676), .Z(n3678) );
  XOR U3888 ( .A(n3679), .B(n3678), .Z(n3670) );
  NAND U3889 ( .A(b[0]), .B(a[151]), .Z(n3671) );
  XOR U3890 ( .A(n3670), .B(n3671), .Z(n3673) );
  OR U3891 ( .A(n3659), .B(n3658), .Z(n3663) );
  NANDN U3892 ( .A(n3661), .B(n3660), .Z(n3662) );
  NAND U3893 ( .A(n3663), .B(n3662), .Z(n3672) );
  XNOR U3894 ( .A(n3673), .B(n3672), .Z(n3682) );
  NANDN U3895 ( .A(n3665), .B(n3664), .Z(n3669) );
  OR U3896 ( .A(n3667), .B(n3666), .Z(n3668) );
  NAND U3897 ( .A(n3669), .B(n3668), .Z(n3683) );
  XNOR U3898 ( .A(n3682), .B(n3683), .Z(n3684) );
  XNOR U3899 ( .A(n3685), .B(n3684), .Z(n3688) );
  XNOR U3900 ( .A(n3688), .B(sreg[403]), .Z(n3689) );
  XOR U3901 ( .A(n3690), .B(n3689), .Z(c[403]) );
  NANDN U3902 ( .A(n3671), .B(n3670), .Z(n3675) );
  OR U3903 ( .A(n3673), .B(n3672), .Z(n3674) );
  NAND U3904 ( .A(n3675), .B(n3674), .Z(n3705) );
  AND U3905 ( .A(b[2]), .B(a[150]), .Z(n3696) );
  AND U3906 ( .A(a[151]), .B(b[1]), .Z(n3694) );
  AND U3907 ( .A(a[149]), .B(b[3]), .Z(n3693) );
  XOR U3908 ( .A(n3694), .B(n3693), .Z(n3695) );
  XOR U3909 ( .A(n3696), .B(n3695), .Z(n3699) );
  NAND U3910 ( .A(b[0]), .B(a[152]), .Z(n3700) );
  XNOR U3911 ( .A(n3699), .B(n3700), .Z(n3701) );
  OR U3912 ( .A(n3677), .B(n3676), .Z(n3681) );
  NANDN U3913 ( .A(n3679), .B(n3678), .Z(n3680) );
  AND U3914 ( .A(n3681), .B(n3680), .Z(n3702) );
  XNOR U3915 ( .A(n3701), .B(n3702), .Z(n3706) );
  XNOR U3916 ( .A(n3705), .B(n3706), .Z(n3707) );
  NANDN U3917 ( .A(n3683), .B(n3682), .Z(n3687) );
  NAND U3918 ( .A(n3685), .B(n3684), .Z(n3686) );
  NAND U3919 ( .A(n3687), .B(n3686), .Z(n3708) );
  XNOR U3920 ( .A(n3707), .B(n3708), .Z(n3711) );
  XOR U3921 ( .A(sreg[404]), .B(n3711), .Z(n3712) );
  NAND U3922 ( .A(n3688), .B(sreg[403]), .Z(n3692) );
  OR U3923 ( .A(n3690), .B(n3689), .Z(n3691) );
  NAND U3924 ( .A(n3692), .B(n3691), .Z(n3713) );
  XOR U3925 ( .A(n3712), .B(n3713), .Z(c[404]) );
  AND U3926 ( .A(b[2]), .B(a[151]), .Z(n3728) );
  AND U3927 ( .A(a[152]), .B(b[1]), .Z(n3726) );
  AND U3928 ( .A(a[150]), .B(b[3]), .Z(n3725) );
  XOR U3929 ( .A(n3726), .B(n3725), .Z(n3727) );
  XOR U3930 ( .A(n3728), .B(n3727), .Z(n3731) );
  NAND U3931 ( .A(b[0]), .B(a[153]), .Z(n3732) );
  XOR U3932 ( .A(n3731), .B(n3732), .Z(n3734) );
  OR U3933 ( .A(n3694), .B(n3693), .Z(n3698) );
  NANDN U3934 ( .A(n3696), .B(n3695), .Z(n3697) );
  NAND U3935 ( .A(n3698), .B(n3697), .Z(n3733) );
  XNOR U3936 ( .A(n3734), .B(n3733), .Z(n3719) );
  NANDN U3937 ( .A(n3700), .B(n3699), .Z(n3704) );
  NAND U3938 ( .A(n3702), .B(n3701), .Z(n3703) );
  NAND U3939 ( .A(n3704), .B(n3703), .Z(n3720) );
  XNOR U3940 ( .A(n3719), .B(n3720), .Z(n3721) );
  NANDN U3941 ( .A(n3706), .B(n3705), .Z(n3710) );
  NANDN U3942 ( .A(n3708), .B(n3707), .Z(n3709) );
  NAND U3943 ( .A(n3710), .B(n3709), .Z(n3722) );
  XOR U3944 ( .A(n3721), .B(n3722), .Z(n3718) );
  OR U3945 ( .A(n3711), .B(sreg[404]), .Z(n3715) );
  NANDN U3946 ( .A(n3713), .B(n3712), .Z(n3714) );
  AND U3947 ( .A(n3715), .B(n3714), .Z(n3717) );
  XNOR U3948 ( .A(sreg[405]), .B(n3717), .Z(n3716) );
  XNOR U3949 ( .A(n3718), .B(n3716), .Z(c[405]) );
  NANDN U3950 ( .A(n3720), .B(n3719), .Z(n3724) );
  NANDN U3951 ( .A(n3722), .B(n3721), .Z(n3723) );
  NAND U3952 ( .A(n3724), .B(n3723), .Z(n3740) );
  AND U3953 ( .A(b[2]), .B(a[152]), .Z(n3746) );
  AND U3954 ( .A(a[153]), .B(b[1]), .Z(n3744) );
  AND U3955 ( .A(a[151]), .B(b[3]), .Z(n3743) );
  XOR U3956 ( .A(n3744), .B(n3743), .Z(n3745) );
  XOR U3957 ( .A(n3746), .B(n3745), .Z(n3749) );
  NAND U3958 ( .A(b[0]), .B(a[154]), .Z(n3750) );
  XOR U3959 ( .A(n3749), .B(n3750), .Z(n3752) );
  OR U3960 ( .A(n3726), .B(n3725), .Z(n3730) );
  NANDN U3961 ( .A(n3728), .B(n3727), .Z(n3729) );
  NAND U3962 ( .A(n3730), .B(n3729), .Z(n3751) );
  XNOR U3963 ( .A(n3752), .B(n3751), .Z(n3737) );
  NANDN U3964 ( .A(n3732), .B(n3731), .Z(n3736) );
  OR U3965 ( .A(n3734), .B(n3733), .Z(n3735) );
  NAND U3966 ( .A(n3736), .B(n3735), .Z(n3738) );
  XNOR U3967 ( .A(n3737), .B(n3738), .Z(n3739) );
  XNOR U3968 ( .A(n3740), .B(n3739), .Z(n3755) );
  XNOR U3969 ( .A(n3755), .B(sreg[406]), .Z(n3756) );
  XOR U3970 ( .A(n3757), .B(n3756), .Z(c[406]) );
  NANDN U3971 ( .A(n3738), .B(n3737), .Z(n3742) );
  NAND U3972 ( .A(n3740), .B(n3739), .Z(n3741) );
  NAND U3973 ( .A(n3742), .B(n3741), .Z(n3763) );
  AND U3974 ( .A(b[2]), .B(a[153]), .Z(n3769) );
  AND U3975 ( .A(a[154]), .B(b[1]), .Z(n3767) );
  AND U3976 ( .A(a[152]), .B(b[3]), .Z(n3766) );
  XOR U3977 ( .A(n3767), .B(n3766), .Z(n3768) );
  XOR U3978 ( .A(n3769), .B(n3768), .Z(n3772) );
  NAND U3979 ( .A(b[0]), .B(a[155]), .Z(n3773) );
  XOR U3980 ( .A(n3772), .B(n3773), .Z(n3775) );
  OR U3981 ( .A(n3744), .B(n3743), .Z(n3748) );
  NANDN U3982 ( .A(n3746), .B(n3745), .Z(n3747) );
  NAND U3983 ( .A(n3748), .B(n3747), .Z(n3774) );
  XNOR U3984 ( .A(n3775), .B(n3774), .Z(n3760) );
  NANDN U3985 ( .A(n3750), .B(n3749), .Z(n3754) );
  OR U3986 ( .A(n3752), .B(n3751), .Z(n3753) );
  NAND U3987 ( .A(n3754), .B(n3753), .Z(n3761) );
  XNOR U3988 ( .A(n3760), .B(n3761), .Z(n3762) );
  XNOR U3989 ( .A(n3763), .B(n3762), .Z(n3778) );
  XNOR U3990 ( .A(n3778), .B(sreg[407]), .Z(n3780) );
  NAND U3991 ( .A(n3755), .B(sreg[406]), .Z(n3759) );
  OR U3992 ( .A(n3757), .B(n3756), .Z(n3758) );
  AND U3993 ( .A(n3759), .B(n3758), .Z(n3779) );
  XOR U3994 ( .A(n3780), .B(n3779), .Z(c[407]) );
  NANDN U3995 ( .A(n3761), .B(n3760), .Z(n3765) );
  NAND U3996 ( .A(n3763), .B(n3762), .Z(n3764) );
  NAND U3997 ( .A(n3765), .B(n3764), .Z(n3791) );
  AND U3998 ( .A(b[2]), .B(a[154]), .Z(n3797) );
  AND U3999 ( .A(a[155]), .B(b[1]), .Z(n3795) );
  AND U4000 ( .A(a[153]), .B(b[3]), .Z(n3794) );
  XOR U4001 ( .A(n3795), .B(n3794), .Z(n3796) );
  XOR U4002 ( .A(n3797), .B(n3796), .Z(n3800) );
  NAND U4003 ( .A(b[0]), .B(a[156]), .Z(n3801) );
  XOR U4004 ( .A(n3800), .B(n3801), .Z(n3803) );
  OR U4005 ( .A(n3767), .B(n3766), .Z(n3771) );
  NANDN U4006 ( .A(n3769), .B(n3768), .Z(n3770) );
  NAND U4007 ( .A(n3771), .B(n3770), .Z(n3802) );
  XNOR U4008 ( .A(n3803), .B(n3802), .Z(n3788) );
  NANDN U4009 ( .A(n3773), .B(n3772), .Z(n3777) );
  OR U4010 ( .A(n3775), .B(n3774), .Z(n3776) );
  NAND U4011 ( .A(n3777), .B(n3776), .Z(n3789) );
  XNOR U4012 ( .A(n3788), .B(n3789), .Z(n3790) );
  XNOR U4013 ( .A(n3791), .B(n3790), .Z(n3783) );
  XOR U4014 ( .A(sreg[408]), .B(n3783), .Z(n3784) );
  NAND U4015 ( .A(n3778), .B(sreg[407]), .Z(n3782) );
  OR U4016 ( .A(n3780), .B(n3779), .Z(n3781) );
  NAND U4017 ( .A(n3782), .B(n3781), .Z(n3785) );
  XOR U4018 ( .A(n3784), .B(n3785), .Z(c[408]) );
  OR U4019 ( .A(n3783), .B(sreg[408]), .Z(n3787) );
  NANDN U4020 ( .A(n3785), .B(n3784), .Z(n3786) );
  AND U4021 ( .A(n3787), .B(n3786), .Z(n3807) );
  NANDN U4022 ( .A(n3789), .B(n3788), .Z(n3793) );
  NAND U4023 ( .A(n3791), .B(n3790), .Z(n3792) );
  NAND U4024 ( .A(n3793), .B(n3792), .Z(n3812) );
  AND U4025 ( .A(b[2]), .B(a[155]), .Z(n3818) );
  AND U4026 ( .A(a[156]), .B(b[1]), .Z(n3816) );
  AND U4027 ( .A(a[154]), .B(b[3]), .Z(n3815) );
  XOR U4028 ( .A(n3816), .B(n3815), .Z(n3817) );
  XOR U4029 ( .A(n3818), .B(n3817), .Z(n3821) );
  NAND U4030 ( .A(b[0]), .B(a[157]), .Z(n3822) );
  XOR U4031 ( .A(n3821), .B(n3822), .Z(n3824) );
  OR U4032 ( .A(n3795), .B(n3794), .Z(n3799) );
  NANDN U4033 ( .A(n3797), .B(n3796), .Z(n3798) );
  NAND U4034 ( .A(n3799), .B(n3798), .Z(n3823) );
  XNOR U4035 ( .A(n3824), .B(n3823), .Z(n3809) );
  NANDN U4036 ( .A(n3801), .B(n3800), .Z(n3805) );
  OR U4037 ( .A(n3803), .B(n3802), .Z(n3804) );
  NAND U4038 ( .A(n3805), .B(n3804), .Z(n3810) );
  XNOR U4039 ( .A(n3809), .B(n3810), .Z(n3811) );
  XNOR U4040 ( .A(n3812), .B(n3811), .Z(n3808) );
  XOR U4041 ( .A(sreg[409]), .B(n3808), .Z(n3806) );
  XOR U4042 ( .A(n3807), .B(n3806), .Z(c[409]) );
  NANDN U4043 ( .A(n3810), .B(n3809), .Z(n3814) );
  NAND U4044 ( .A(n3812), .B(n3811), .Z(n3813) );
  NAND U4045 ( .A(n3814), .B(n3813), .Z(n3830) );
  AND U4046 ( .A(b[2]), .B(a[156]), .Z(n3836) );
  AND U4047 ( .A(a[157]), .B(b[1]), .Z(n3834) );
  AND U4048 ( .A(a[155]), .B(b[3]), .Z(n3833) );
  XOR U4049 ( .A(n3834), .B(n3833), .Z(n3835) );
  XOR U4050 ( .A(n3836), .B(n3835), .Z(n3839) );
  NAND U4051 ( .A(b[0]), .B(a[158]), .Z(n3840) );
  XOR U4052 ( .A(n3839), .B(n3840), .Z(n3842) );
  OR U4053 ( .A(n3816), .B(n3815), .Z(n3820) );
  NANDN U4054 ( .A(n3818), .B(n3817), .Z(n3819) );
  NAND U4055 ( .A(n3820), .B(n3819), .Z(n3841) );
  XNOR U4056 ( .A(n3842), .B(n3841), .Z(n3827) );
  NANDN U4057 ( .A(n3822), .B(n3821), .Z(n3826) );
  OR U4058 ( .A(n3824), .B(n3823), .Z(n3825) );
  NAND U4059 ( .A(n3826), .B(n3825), .Z(n3828) );
  XNOR U4060 ( .A(n3827), .B(n3828), .Z(n3829) );
  XOR U4061 ( .A(n3830), .B(n3829), .Z(n3845) );
  XOR U4062 ( .A(sreg[410]), .B(n3845), .Z(n3847) );
  XNOR U4063 ( .A(n3846), .B(n3847), .Z(c[410]) );
  NANDN U4064 ( .A(n3828), .B(n3827), .Z(n3832) );
  NAND U4065 ( .A(n3830), .B(n3829), .Z(n3831) );
  NAND U4066 ( .A(n3832), .B(n3831), .Z(n3853) );
  AND U4067 ( .A(b[2]), .B(a[157]), .Z(n3859) );
  AND U4068 ( .A(a[158]), .B(b[1]), .Z(n3857) );
  AND U4069 ( .A(a[156]), .B(b[3]), .Z(n3856) );
  XOR U4070 ( .A(n3857), .B(n3856), .Z(n3858) );
  XOR U4071 ( .A(n3859), .B(n3858), .Z(n3862) );
  NAND U4072 ( .A(b[0]), .B(a[159]), .Z(n3863) );
  XOR U4073 ( .A(n3862), .B(n3863), .Z(n3865) );
  OR U4074 ( .A(n3834), .B(n3833), .Z(n3838) );
  NANDN U4075 ( .A(n3836), .B(n3835), .Z(n3837) );
  NAND U4076 ( .A(n3838), .B(n3837), .Z(n3864) );
  XNOR U4077 ( .A(n3865), .B(n3864), .Z(n3850) );
  NANDN U4078 ( .A(n3840), .B(n3839), .Z(n3844) );
  OR U4079 ( .A(n3842), .B(n3841), .Z(n3843) );
  NAND U4080 ( .A(n3844), .B(n3843), .Z(n3851) );
  XNOR U4081 ( .A(n3850), .B(n3851), .Z(n3852) );
  XNOR U4082 ( .A(n3853), .B(n3852), .Z(n3868) );
  XOR U4083 ( .A(sreg[411]), .B(n3868), .Z(n3869) );
  NANDN U4084 ( .A(n3845), .B(sreg[410]), .Z(n3849) );
  NANDN U4085 ( .A(n3847), .B(n3846), .Z(n3848) );
  NAND U4086 ( .A(n3849), .B(n3848), .Z(n3870) );
  XOR U4087 ( .A(n3869), .B(n3870), .Z(c[411]) );
  NANDN U4088 ( .A(n3851), .B(n3850), .Z(n3855) );
  NAND U4089 ( .A(n3853), .B(n3852), .Z(n3854) );
  NAND U4090 ( .A(n3855), .B(n3854), .Z(n3877) );
  AND U4091 ( .A(b[2]), .B(a[158]), .Z(n3883) );
  AND U4092 ( .A(a[159]), .B(b[1]), .Z(n3881) );
  AND U4093 ( .A(a[157]), .B(b[3]), .Z(n3880) );
  XOR U4094 ( .A(n3881), .B(n3880), .Z(n3882) );
  XOR U4095 ( .A(n3883), .B(n3882), .Z(n3886) );
  NAND U4096 ( .A(b[0]), .B(a[160]), .Z(n3887) );
  XOR U4097 ( .A(n3886), .B(n3887), .Z(n3889) );
  OR U4098 ( .A(n3857), .B(n3856), .Z(n3861) );
  NANDN U4099 ( .A(n3859), .B(n3858), .Z(n3860) );
  NAND U4100 ( .A(n3861), .B(n3860), .Z(n3888) );
  XNOR U4101 ( .A(n3889), .B(n3888), .Z(n3874) );
  NANDN U4102 ( .A(n3863), .B(n3862), .Z(n3867) );
  OR U4103 ( .A(n3865), .B(n3864), .Z(n3866) );
  NAND U4104 ( .A(n3867), .B(n3866), .Z(n3875) );
  XNOR U4105 ( .A(n3874), .B(n3875), .Z(n3876) );
  XOR U4106 ( .A(n3877), .B(n3876), .Z(n3893) );
  OR U4107 ( .A(n3868), .B(sreg[411]), .Z(n3872) );
  NANDN U4108 ( .A(n3870), .B(n3869), .Z(n3871) );
  AND U4109 ( .A(n3872), .B(n3871), .Z(n3892) );
  XNOR U4110 ( .A(sreg[412]), .B(n3892), .Z(n3873) );
  XOR U4111 ( .A(n3893), .B(n3873), .Z(c[412]) );
  NANDN U4112 ( .A(n3875), .B(n3874), .Z(n3879) );
  NAND U4113 ( .A(n3877), .B(n3876), .Z(n3878) );
  NAND U4114 ( .A(n3879), .B(n3878), .Z(n3900) );
  AND U4115 ( .A(b[2]), .B(a[159]), .Z(n3906) );
  AND U4116 ( .A(a[160]), .B(b[1]), .Z(n3904) );
  AND U4117 ( .A(a[158]), .B(b[3]), .Z(n3903) );
  XOR U4118 ( .A(n3904), .B(n3903), .Z(n3905) );
  XOR U4119 ( .A(n3906), .B(n3905), .Z(n3909) );
  NAND U4120 ( .A(b[0]), .B(a[161]), .Z(n3910) );
  XOR U4121 ( .A(n3909), .B(n3910), .Z(n3912) );
  OR U4122 ( .A(n3881), .B(n3880), .Z(n3885) );
  NANDN U4123 ( .A(n3883), .B(n3882), .Z(n3884) );
  NAND U4124 ( .A(n3885), .B(n3884), .Z(n3911) );
  XNOR U4125 ( .A(n3912), .B(n3911), .Z(n3897) );
  NANDN U4126 ( .A(n3887), .B(n3886), .Z(n3891) );
  OR U4127 ( .A(n3889), .B(n3888), .Z(n3890) );
  NAND U4128 ( .A(n3891), .B(n3890), .Z(n3898) );
  XNOR U4129 ( .A(n3897), .B(n3898), .Z(n3899) );
  XOR U4130 ( .A(n3900), .B(n3899), .Z(n3896) );
  XNOR U4131 ( .A(sreg[413]), .B(n3895), .Z(n3894) );
  XOR U4132 ( .A(n3896), .B(n3894), .Z(c[413]) );
  NANDN U4133 ( .A(n3898), .B(n3897), .Z(n3902) );
  NAND U4134 ( .A(n3900), .B(n3899), .Z(n3901) );
  NAND U4135 ( .A(n3902), .B(n3901), .Z(n3918) );
  AND U4136 ( .A(b[2]), .B(a[160]), .Z(n3924) );
  AND U4137 ( .A(a[161]), .B(b[1]), .Z(n3922) );
  AND U4138 ( .A(a[159]), .B(b[3]), .Z(n3921) );
  XOR U4139 ( .A(n3922), .B(n3921), .Z(n3923) );
  XOR U4140 ( .A(n3924), .B(n3923), .Z(n3927) );
  NAND U4141 ( .A(b[0]), .B(a[162]), .Z(n3928) );
  XOR U4142 ( .A(n3927), .B(n3928), .Z(n3930) );
  OR U4143 ( .A(n3904), .B(n3903), .Z(n3908) );
  NANDN U4144 ( .A(n3906), .B(n3905), .Z(n3907) );
  NAND U4145 ( .A(n3908), .B(n3907), .Z(n3929) );
  XNOR U4146 ( .A(n3930), .B(n3929), .Z(n3915) );
  NANDN U4147 ( .A(n3910), .B(n3909), .Z(n3914) );
  OR U4148 ( .A(n3912), .B(n3911), .Z(n3913) );
  NAND U4149 ( .A(n3914), .B(n3913), .Z(n3916) );
  XNOR U4150 ( .A(n3915), .B(n3916), .Z(n3917) );
  XNOR U4151 ( .A(n3918), .B(n3917), .Z(n3933) );
  XNOR U4152 ( .A(n3933), .B(sreg[414]), .Z(n3934) );
  XOR U4153 ( .A(n3935), .B(n3934), .Z(c[414]) );
  NANDN U4154 ( .A(n3916), .B(n3915), .Z(n3920) );
  NAND U4155 ( .A(n3918), .B(n3917), .Z(n3919) );
  NAND U4156 ( .A(n3920), .B(n3919), .Z(n3946) );
  AND U4157 ( .A(b[2]), .B(a[161]), .Z(n3952) );
  AND U4158 ( .A(a[162]), .B(b[1]), .Z(n3950) );
  AND U4159 ( .A(a[160]), .B(b[3]), .Z(n3949) );
  XOR U4160 ( .A(n3950), .B(n3949), .Z(n3951) );
  XOR U4161 ( .A(n3952), .B(n3951), .Z(n3955) );
  NAND U4162 ( .A(b[0]), .B(a[163]), .Z(n3956) );
  XOR U4163 ( .A(n3955), .B(n3956), .Z(n3958) );
  OR U4164 ( .A(n3922), .B(n3921), .Z(n3926) );
  NANDN U4165 ( .A(n3924), .B(n3923), .Z(n3925) );
  NAND U4166 ( .A(n3926), .B(n3925), .Z(n3957) );
  XNOR U4167 ( .A(n3958), .B(n3957), .Z(n3943) );
  NANDN U4168 ( .A(n3928), .B(n3927), .Z(n3932) );
  OR U4169 ( .A(n3930), .B(n3929), .Z(n3931) );
  NAND U4170 ( .A(n3932), .B(n3931), .Z(n3944) );
  XNOR U4171 ( .A(n3943), .B(n3944), .Z(n3945) );
  XNOR U4172 ( .A(n3946), .B(n3945), .Z(n3938) );
  XOR U4173 ( .A(sreg[415]), .B(n3938), .Z(n3939) );
  NAND U4174 ( .A(n3933), .B(sreg[414]), .Z(n3937) );
  OR U4175 ( .A(n3935), .B(n3934), .Z(n3936) );
  NAND U4176 ( .A(n3937), .B(n3936), .Z(n3940) );
  XOR U4177 ( .A(n3939), .B(n3940), .Z(c[415]) );
  OR U4178 ( .A(n3938), .B(sreg[415]), .Z(n3942) );
  NANDN U4179 ( .A(n3940), .B(n3939), .Z(n3941) );
  AND U4180 ( .A(n3942), .B(n3941), .Z(n3962) );
  NANDN U4181 ( .A(n3944), .B(n3943), .Z(n3948) );
  NAND U4182 ( .A(n3946), .B(n3945), .Z(n3947) );
  NAND U4183 ( .A(n3948), .B(n3947), .Z(n3967) );
  AND U4184 ( .A(b[2]), .B(a[162]), .Z(n3973) );
  AND U4185 ( .A(a[163]), .B(b[1]), .Z(n3971) );
  AND U4186 ( .A(a[161]), .B(b[3]), .Z(n3970) );
  XOR U4187 ( .A(n3971), .B(n3970), .Z(n3972) );
  XOR U4188 ( .A(n3973), .B(n3972), .Z(n3976) );
  NAND U4189 ( .A(b[0]), .B(a[164]), .Z(n3977) );
  XOR U4190 ( .A(n3976), .B(n3977), .Z(n3979) );
  OR U4191 ( .A(n3950), .B(n3949), .Z(n3954) );
  NANDN U4192 ( .A(n3952), .B(n3951), .Z(n3953) );
  NAND U4193 ( .A(n3954), .B(n3953), .Z(n3978) );
  XNOR U4194 ( .A(n3979), .B(n3978), .Z(n3964) );
  NANDN U4195 ( .A(n3956), .B(n3955), .Z(n3960) );
  OR U4196 ( .A(n3958), .B(n3957), .Z(n3959) );
  NAND U4197 ( .A(n3960), .B(n3959), .Z(n3965) );
  XNOR U4198 ( .A(n3964), .B(n3965), .Z(n3966) );
  XNOR U4199 ( .A(n3967), .B(n3966), .Z(n3963) );
  XOR U4200 ( .A(sreg[416]), .B(n3963), .Z(n3961) );
  XOR U4201 ( .A(n3962), .B(n3961), .Z(c[416]) );
  NANDN U4202 ( .A(n3965), .B(n3964), .Z(n3969) );
  NAND U4203 ( .A(n3967), .B(n3966), .Z(n3968) );
  NAND U4204 ( .A(n3969), .B(n3968), .Z(n3985) );
  AND U4205 ( .A(b[2]), .B(a[163]), .Z(n3991) );
  AND U4206 ( .A(a[164]), .B(b[1]), .Z(n3989) );
  AND U4207 ( .A(a[162]), .B(b[3]), .Z(n3988) );
  XOR U4208 ( .A(n3989), .B(n3988), .Z(n3990) );
  XOR U4209 ( .A(n3991), .B(n3990), .Z(n3994) );
  NAND U4210 ( .A(b[0]), .B(a[165]), .Z(n3995) );
  XOR U4211 ( .A(n3994), .B(n3995), .Z(n3997) );
  OR U4212 ( .A(n3971), .B(n3970), .Z(n3975) );
  NANDN U4213 ( .A(n3973), .B(n3972), .Z(n3974) );
  NAND U4214 ( .A(n3975), .B(n3974), .Z(n3996) );
  XNOR U4215 ( .A(n3997), .B(n3996), .Z(n3982) );
  NANDN U4216 ( .A(n3977), .B(n3976), .Z(n3981) );
  OR U4217 ( .A(n3979), .B(n3978), .Z(n3980) );
  NAND U4218 ( .A(n3981), .B(n3980), .Z(n3983) );
  XNOR U4219 ( .A(n3982), .B(n3983), .Z(n3984) );
  XNOR U4220 ( .A(n3985), .B(n3984), .Z(n4000) );
  XNOR U4221 ( .A(n4000), .B(sreg[417]), .Z(n4002) );
  XNOR U4222 ( .A(n4001), .B(n4002), .Z(c[417]) );
  NANDN U4223 ( .A(n3983), .B(n3982), .Z(n3987) );
  NAND U4224 ( .A(n3985), .B(n3984), .Z(n3986) );
  NAND U4225 ( .A(n3987), .B(n3986), .Z(n4011) );
  AND U4226 ( .A(b[2]), .B(a[164]), .Z(n4017) );
  AND U4227 ( .A(a[165]), .B(b[1]), .Z(n4015) );
  AND U4228 ( .A(a[163]), .B(b[3]), .Z(n4014) );
  XOR U4229 ( .A(n4015), .B(n4014), .Z(n4016) );
  XOR U4230 ( .A(n4017), .B(n4016), .Z(n4020) );
  NAND U4231 ( .A(b[0]), .B(a[166]), .Z(n4021) );
  XOR U4232 ( .A(n4020), .B(n4021), .Z(n4023) );
  OR U4233 ( .A(n3989), .B(n3988), .Z(n3993) );
  NANDN U4234 ( .A(n3991), .B(n3990), .Z(n3992) );
  NAND U4235 ( .A(n3993), .B(n3992), .Z(n4022) );
  XNOR U4236 ( .A(n4023), .B(n4022), .Z(n4008) );
  NANDN U4237 ( .A(n3995), .B(n3994), .Z(n3999) );
  OR U4238 ( .A(n3997), .B(n3996), .Z(n3998) );
  NAND U4239 ( .A(n3999), .B(n3998), .Z(n4009) );
  XNOR U4240 ( .A(n4008), .B(n4009), .Z(n4010) );
  XOR U4241 ( .A(n4011), .B(n4010), .Z(n4007) );
  NAND U4242 ( .A(n4000), .B(sreg[417]), .Z(n4004) );
  NANDN U4243 ( .A(n4002), .B(n4001), .Z(n4003) );
  NAND U4244 ( .A(n4004), .B(n4003), .Z(n4006) );
  XNOR U4245 ( .A(sreg[418]), .B(n4006), .Z(n4005) );
  XOR U4246 ( .A(n4007), .B(n4005), .Z(c[418]) );
  NANDN U4247 ( .A(n4009), .B(n4008), .Z(n4013) );
  NAND U4248 ( .A(n4011), .B(n4010), .Z(n4012) );
  NAND U4249 ( .A(n4013), .B(n4012), .Z(n4029) );
  AND U4250 ( .A(b[2]), .B(a[165]), .Z(n4035) );
  AND U4251 ( .A(a[166]), .B(b[1]), .Z(n4033) );
  AND U4252 ( .A(a[164]), .B(b[3]), .Z(n4032) );
  XOR U4253 ( .A(n4033), .B(n4032), .Z(n4034) );
  XOR U4254 ( .A(n4035), .B(n4034), .Z(n4038) );
  NAND U4255 ( .A(b[0]), .B(a[167]), .Z(n4039) );
  XOR U4256 ( .A(n4038), .B(n4039), .Z(n4041) );
  OR U4257 ( .A(n4015), .B(n4014), .Z(n4019) );
  NANDN U4258 ( .A(n4017), .B(n4016), .Z(n4018) );
  NAND U4259 ( .A(n4019), .B(n4018), .Z(n4040) );
  XNOR U4260 ( .A(n4041), .B(n4040), .Z(n4026) );
  NANDN U4261 ( .A(n4021), .B(n4020), .Z(n4025) );
  OR U4262 ( .A(n4023), .B(n4022), .Z(n4024) );
  NAND U4263 ( .A(n4025), .B(n4024), .Z(n4027) );
  XNOR U4264 ( .A(n4026), .B(n4027), .Z(n4028) );
  XNOR U4265 ( .A(n4029), .B(n4028), .Z(n4044) );
  XNOR U4266 ( .A(n4044), .B(sreg[419]), .Z(n4045) );
  XOR U4267 ( .A(n4046), .B(n4045), .Z(c[419]) );
  NANDN U4268 ( .A(n4027), .B(n4026), .Z(n4031) );
  NAND U4269 ( .A(n4029), .B(n4028), .Z(n4030) );
  NAND U4270 ( .A(n4031), .B(n4030), .Z(n4052) );
  AND U4271 ( .A(b[2]), .B(a[166]), .Z(n4058) );
  AND U4272 ( .A(a[167]), .B(b[1]), .Z(n4056) );
  AND U4273 ( .A(a[165]), .B(b[3]), .Z(n4055) );
  XOR U4274 ( .A(n4056), .B(n4055), .Z(n4057) );
  XOR U4275 ( .A(n4058), .B(n4057), .Z(n4061) );
  NAND U4276 ( .A(b[0]), .B(a[168]), .Z(n4062) );
  XOR U4277 ( .A(n4061), .B(n4062), .Z(n4064) );
  OR U4278 ( .A(n4033), .B(n4032), .Z(n4037) );
  NANDN U4279 ( .A(n4035), .B(n4034), .Z(n4036) );
  NAND U4280 ( .A(n4037), .B(n4036), .Z(n4063) );
  XNOR U4281 ( .A(n4064), .B(n4063), .Z(n4049) );
  NANDN U4282 ( .A(n4039), .B(n4038), .Z(n4043) );
  OR U4283 ( .A(n4041), .B(n4040), .Z(n4042) );
  NAND U4284 ( .A(n4043), .B(n4042), .Z(n4050) );
  XNOR U4285 ( .A(n4049), .B(n4050), .Z(n4051) );
  XNOR U4286 ( .A(n4052), .B(n4051), .Z(n4067) );
  XNOR U4287 ( .A(n4067), .B(sreg[420]), .Z(n4069) );
  NAND U4288 ( .A(n4044), .B(sreg[419]), .Z(n4048) );
  OR U4289 ( .A(n4046), .B(n4045), .Z(n4047) );
  AND U4290 ( .A(n4048), .B(n4047), .Z(n4068) );
  XOR U4291 ( .A(n4069), .B(n4068), .Z(c[420]) );
  NANDN U4292 ( .A(n4050), .B(n4049), .Z(n4054) );
  NAND U4293 ( .A(n4052), .B(n4051), .Z(n4053) );
  NAND U4294 ( .A(n4054), .B(n4053), .Z(n4075) );
  AND U4295 ( .A(b[2]), .B(a[167]), .Z(n4081) );
  AND U4296 ( .A(a[168]), .B(b[1]), .Z(n4079) );
  AND U4297 ( .A(a[166]), .B(b[3]), .Z(n4078) );
  XOR U4298 ( .A(n4079), .B(n4078), .Z(n4080) );
  XOR U4299 ( .A(n4081), .B(n4080), .Z(n4084) );
  NAND U4300 ( .A(b[0]), .B(a[169]), .Z(n4085) );
  XOR U4301 ( .A(n4084), .B(n4085), .Z(n4087) );
  OR U4302 ( .A(n4056), .B(n4055), .Z(n4060) );
  NANDN U4303 ( .A(n4058), .B(n4057), .Z(n4059) );
  NAND U4304 ( .A(n4060), .B(n4059), .Z(n4086) );
  XNOR U4305 ( .A(n4087), .B(n4086), .Z(n4072) );
  NANDN U4306 ( .A(n4062), .B(n4061), .Z(n4066) );
  OR U4307 ( .A(n4064), .B(n4063), .Z(n4065) );
  NAND U4308 ( .A(n4066), .B(n4065), .Z(n4073) );
  XNOR U4309 ( .A(n4072), .B(n4073), .Z(n4074) );
  XNOR U4310 ( .A(n4075), .B(n4074), .Z(n4090) );
  XNOR U4311 ( .A(n4090), .B(sreg[421]), .Z(n4092) );
  NAND U4312 ( .A(n4067), .B(sreg[420]), .Z(n4071) );
  OR U4313 ( .A(n4069), .B(n4068), .Z(n4070) );
  AND U4314 ( .A(n4071), .B(n4070), .Z(n4091) );
  XOR U4315 ( .A(n4092), .B(n4091), .Z(c[421]) );
  NANDN U4316 ( .A(n4073), .B(n4072), .Z(n4077) );
  NAND U4317 ( .A(n4075), .B(n4074), .Z(n4076) );
  NAND U4318 ( .A(n4077), .B(n4076), .Z(n4101) );
  AND U4319 ( .A(b[2]), .B(a[168]), .Z(n4107) );
  AND U4320 ( .A(a[169]), .B(b[1]), .Z(n4105) );
  AND U4321 ( .A(a[167]), .B(b[3]), .Z(n4104) );
  XOR U4322 ( .A(n4105), .B(n4104), .Z(n4106) );
  XOR U4323 ( .A(n4107), .B(n4106), .Z(n4110) );
  NAND U4324 ( .A(b[0]), .B(a[170]), .Z(n4111) );
  XOR U4325 ( .A(n4110), .B(n4111), .Z(n4113) );
  OR U4326 ( .A(n4079), .B(n4078), .Z(n4083) );
  NANDN U4327 ( .A(n4081), .B(n4080), .Z(n4082) );
  NAND U4328 ( .A(n4083), .B(n4082), .Z(n4112) );
  XNOR U4329 ( .A(n4113), .B(n4112), .Z(n4098) );
  NANDN U4330 ( .A(n4085), .B(n4084), .Z(n4089) );
  OR U4331 ( .A(n4087), .B(n4086), .Z(n4088) );
  NAND U4332 ( .A(n4089), .B(n4088), .Z(n4099) );
  XNOR U4333 ( .A(n4098), .B(n4099), .Z(n4100) );
  XOR U4334 ( .A(n4101), .B(n4100), .Z(n4097) );
  NAND U4335 ( .A(n4090), .B(sreg[421]), .Z(n4094) );
  OR U4336 ( .A(n4092), .B(n4091), .Z(n4093) );
  NAND U4337 ( .A(n4094), .B(n4093), .Z(n4096) );
  XNOR U4338 ( .A(sreg[422]), .B(n4096), .Z(n4095) );
  XOR U4339 ( .A(n4097), .B(n4095), .Z(c[422]) );
  NANDN U4340 ( .A(n4099), .B(n4098), .Z(n4103) );
  NAND U4341 ( .A(n4101), .B(n4100), .Z(n4102) );
  NAND U4342 ( .A(n4103), .B(n4102), .Z(n4119) );
  AND U4343 ( .A(b[2]), .B(a[169]), .Z(n4125) );
  AND U4344 ( .A(a[170]), .B(b[1]), .Z(n4123) );
  AND U4345 ( .A(a[168]), .B(b[3]), .Z(n4122) );
  XOR U4346 ( .A(n4123), .B(n4122), .Z(n4124) );
  XOR U4347 ( .A(n4125), .B(n4124), .Z(n4128) );
  NAND U4348 ( .A(b[0]), .B(a[171]), .Z(n4129) );
  XOR U4349 ( .A(n4128), .B(n4129), .Z(n4131) );
  OR U4350 ( .A(n4105), .B(n4104), .Z(n4109) );
  NANDN U4351 ( .A(n4107), .B(n4106), .Z(n4108) );
  NAND U4352 ( .A(n4109), .B(n4108), .Z(n4130) );
  XNOR U4353 ( .A(n4131), .B(n4130), .Z(n4116) );
  NANDN U4354 ( .A(n4111), .B(n4110), .Z(n4115) );
  OR U4355 ( .A(n4113), .B(n4112), .Z(n4114) );
  NAND U4356 ( .A(n4115), .B(n4114), .Z(n4117) );
  XNOR U4357 ( .A(n4116), .B(n4117), .Z(n4118) );
  XNOR U4358 ( .A(n4119), .B(n4118), .Z(n4134) );
  XNOR U4359 ( .A(n4134), .B(sreg[423]), .Z(n4135) );
  XOR U4360 ( .A(n4136), .B(n4135), .Z(c[423]) );
  NANDN U4361 ( .A(n4117), .B(n4116), .Z(n4121) );
  NAND U4362 ( .A(n4119), .B(n4118), .Z(n4120) );
  NAND U4363 ( .A(n4121), .B(n4120), .Z(n4143) );
  AND U4364 ( .A(b[2]), .B(a[170]), .Z(n4149) );
  AND U4365 ( .A(a[171]), .B(b[1]), .Z(n4147) );
  AND U4366 ( .A(a[169]), .B(b[3]), .Z(n4146) );
  XOR U4367 ( .A(n4147), .B(n4146), .Z(n4148) );
  XOR U4368 ( .A(n4149), .B(n4148), .Z(n4152) );
  NAND U4369 ( .A(b[0]), .B(a[172]), .Z(n4153) );
  XOR U4370 ( .A(n4152), .B(n4153), .Z(n4155) );
  OR U4371 ( .A(n4123), .B(n4122), .Z(n4127) );
  NANDN U4372 ( .A(n4125), .B(n4124), .Z(n4126) );
  NAND U4373 ( .A(n4127), .B(n4126), .Z(n4154) );
  XNOR U4374 ( .A(n4155), .B(n4154), .Z(n4140) );
  NANDN U4375 ( .A(n4129), .B(n4128), .Z(n4133) );
  OR U4376 ( .A(n4131), .B(n4130), .Z(n4132) );
  NAND U4377 ( .A(n4133), .B(n4132), .Z(n4141) );
  XNOR U4378 ( .A(n4140), .B(n4141), .Z(n4142) );
  XNOR U4379 ( .A(n4143), .B(n4142), .Z(n4159) );
  NAND U4380 ( .A(n4134), .B(sreg[423]), .Z(n4138) );
  OR U4381 ( .A(n4136), .B(n4135), .Z(n4137) );
  AND U4382 ( .A(n4138), .B(n4137), .Z(n4158) );
  XNOR U4383 ( .A(n4158), .B(sreg[424]), .Z(n4139) );
  XOR U4384 ( .A(n4159), .B(n4139), .Z(c[424]) );
  NANDN U4385 ( .A(n4141), .B(n4140), .Z(n4145) );
  NAND U4386 ( .A(n4143), .B(n4142), .Z(n4144) );
  NAND U4387 ( .A(n4145), .B(n4144), .Z(n4164) );
  AND U4388 ( .A(b[2]), .B(a[171]), .Z(n4170) );
  AND U4389 ( .A(a[172]), .B(b[1]), .Z(n4168) );
  AND U4390 ( .A(a[170]), .B(b[3]), .Z(n4167) );
  XOR U4391 ( .A(n4168), .B(n4167), .Z(n4169) );
  XOR U4392 ( .A(n4170), .B(n4169), .Z(n4173) );
  NAND U4393 ( .A(b[0]), .B(a[173]), .Z(n4174) );
  XOR U4394 ( .A(n4173), .B(n4174), .Z(n4176) );
  OR U4395 ( .A(n4147), .B(n4146), .Z(n4151) );
  NANDN U4396 ( .A(n4149), .B(n4148), .Z(n4150) );
  NAND U4397 ( .A(n4151), .B(n4150), .Z(n4175) );
  XNOR U4398 ( .A(n4176), .B(n4175), .Z(n4161) );
  NANDN U4399 ( .A(n4153), .B(n4152), .Z(n4157) );
  OR U4400 ( .A(n4155), .B(n4154), .Z(n4156) );
  NAND U4401 ( .A(n4157), .B(n4156), .Z(n4162) );
  XNOR U4402 ( .A(n4161), .B(n4162), .Z(n4163) );
  XNOR U4403 ( .A(n4164), .B(n4163), .Z(n4180) );
  XOR U4404 ( .A(n4179), .B(sreg[425]), .Z(n4160) );
  XOR U4405 ( .A(n4180), .B(n4160), .Z(c[425]) );
  NANDN U4406 ( .A(n4162), .B(n4161), .Z(n4166) );
  NAND U4407 ( .A(n4164), .B(n4163), .Z(n4165) );
  NAND U4408 ( .A(n4166), .B(n4165), .Z(n4187) );
  AND U4409 ( .A(b[2]), .B(a[172]), .Z(n4193) );
  AND U4410 ( .A(a[173]), .B(b[1]), .Z(n4191) );
  AND U4411 ( .A(a[171]), .B(b[3]), .Z(n4190) );
  XOR U4412 ( .A(n4191), .B(n4190), .Z(n4192) );
  XOR U4413 ( .A(n4193), .B(n4192), .Z(n4196) );
  NAND U4414 ( .A(b[0]), .B(a[174]), .Z(n4197) );
  XOR U4415 ( .A(n4196), .B(n4197), .Z(n4199) );
  OR U4416 ( .A(n4168), .B(n4167), .Z(n4172) );
  NANDN U4417 ( .A(n4170), .B(n4169), .Z(n4171) );
  NAND U4418 ( .A(n4172), .B(n4171), .Z(n4198) );
  XNOR U4419 ( .A(n4199), .B(n4198), .Z(n4184) );
  NANDN U4420 ( .A(n4174), .B(n4173), .Z(n4178) );
  OR U4421 ( .A(n4176), .B(n4175), .Z(n4177) );
  NAND U4422 ( .A(n4178), .B(n4177), .Z(n4185) );
  XNOR U4423 ( .A(n4184), .B(n4185), .Z(n4186) );
  XOR U4424 ( .A(n4187), .B(n4186), .Z(n4183) );
  XOR U4425 ( .A(sreg[426]), .B(n4182), .Z(n4181) );
  XOR U4426 ( .A(n4183), .B(n4181), .Z(c[426]) );
  NANDN U4427 ( .A(n4185), .B(n4184), .Z(n4189) );
  NAND U4428 ( .A(n4187), .B(n4186), .Z(n4188) );
  NAND U4429 ( .A(n4189), .B(n4188), .Z(n4205) );
  AND U4430 ( .A(b[2]), .B(a[173]), .Z(n4211) );
  AND U4431 ( .A(a[174]), .B(b[1]), .Z(n4209) );
  AND U4432 ( .A(a[172]), .B(b[3]), .Z(n4208) );
  XOR U4433 ( .A(n4209), .B(n4208), .Z(n4210) );
  XOR U4434 ( .A(n4211), .B(n4210), .Z(n4214) );
  NAND U4435 ( .A(b[0]), .B(a[175]), .Z(n4215) );
  XOR U4436 ( .A(n4214), .B(n4215), .Z(n4217) );
  OR U4437 ( .A(n4191), .B(n4190), .Z(n4195) );
  NANDN U4438 ( .A(n4193), .B(n4192), .Z(n4194) );
  NAND U4439 ( .A(n4195), .B(n4194), .Z(n4216) );
  XNOR U4440 ( .A(n4217), .B(n4216), .Z(n4202) );
  NANDN U4441 ( .A(n4197), .B(n4196), .Z(n4201) );
  OR U4442 ( .A(n4199), .B(n4198), .Z(n4200) );
  NAND U4443 ( .A(n4201), .B(n4200), .Z(n4203) );
  XNOR U4444 ( .A(n4202), .B(n4203), .Z(n4204) );
  XNOR U4445 ( .A(n4205), .B(n4204), .Z(n4220) );
  XNOR U4446 ( .A(n4220), .B(sreg[427]), .Z(n4221) );
  XOR U4447 ( .A(n4222), .B(n4221), .Z(c[427]) );
  NANDN U4448 ( .A(n4203), .B(n4202), .Z(n4207) );
  NAND U4449 ( .A(n4205), .B(n4204), .Z(n4206) );
  NAND U4450 ( .A(n4207), .B(n4206), .Z(n4231) );
  AND U4451 ( .A(b[2]), .B(a[174]), .Z(n4243) );
  AND U4452 ( .A(a[175]), .B(b[1]), .Z(n4241) );
  AND U4453 ( .A(a[173]), .B(b[3]), .Z(n4240) );
  XOR U4454 ( .A(n4241), .B(n4240), .Z(n4242) );
  XOR U4455 ( .A(n4243), .B(n4242), .Z(n4234) );
  NAND U4456 ( .A(b[0]), .B(a[176]), .Z(n4235) );
  XOR U4457 ( .A(n4234), .B(n4235), .Z(n4237) );
  OR U4458 ( .A(n4209), .B(n4208), .Z(n4213) );
  NANDN U4459 ( .A(n4211), .B(n4210), .Z(n4212) );
  NAND U4460 ( .A(n4213), .B(n4212), .Z(n4236) );
  XNOR U4461 ( .A(n4237), .B(n4236), .Z(n4228) );
  NANDN U4462 ( .A(n4215), .B(n4214), .Z(n4219) );
  OR U4463 ( .A(n4217), .B(n4216), .Z(n4218) );
  NAND U4464 ( .A(n4219), .B(n4218), .Z(n4229) );
  XNOR U4465 ( .A(n4228), .B(n4229), .Z(n4230) );
  XOR U4466 ( .A(n4231), .B(n4230), .Z(n4227) );
  NAND U4467 ( .A(n4220), .B(sreg[427]), .Z(n4224) );
  OR U4468 ( .A(n4222), .B(n4221), .Z(n4223) );
  NAND U4469 ( .A(n4224), .B(n4223), .Z(n4226) );
  XNOR U4470 ( .A(sreg[428]), .B(n4226), .Z(n4225) );
  XOR U4471 ( .A(n4227), .B(n4225), .Z(c[428]) );
  NANDN U4472 ( .A(n4229), .B(n4228), .Z(n4233) );
  NAND U4473 ( .A(n4231), .B(n4230), .Z(n4232) );
  NAND U4474 ( .A(n4233), .B(n4232), .Z(n4249) );
  NANDN U4475 ( .A(n4235), .B(n4234), .Z(n4239) );
  OR U4476 ( .A(n4237), .B(n4236), .Z(n4238) );
  AND U4477 ( .A(n4239), .B(n4238), .Z(n4248) );
  AND U4478 ( .A(b[2]), .B(a[175]), .Z(n4253) );
  AND U4479 ( .A(a[176]), .B(b[1]), .Z(n4251) );
  AND U4480 ( .A(a[174]), .B(b[3]), .Z(n4250) );
  XOR U4481 ( .A(n4251), .B(n4250), .Z(n4252) );
  XOR U4482 ( .A(n4253), .B(n4252), .Z(n4256) );
  NAND U4483 ( .A(b[0]), .B(a[177]), .Z(n4257) );
  XOR U4484 ( .A(n4256), .B(n4257), .Z(n4259) );
  OR U4485 ( .A(n4241), .B(n4240), .Z(n4245) );
  NANDN U4486 ( .A(n4243), .B(n4242), .Z(n4244) );
  NAND U4487 ( .A(n4245), .B(n4244), .Z(n4258) );
  XOR U4488 ( .A(n4259), .B(n4258), .Z(n4247) );
  XNOR U4489 ( .A(n4248), .B(n4247), .Z(n4246) );
  XNOR U4490 ( .A(n4249), .B(n4246), .Z(n4262) );
  XOR U4491 ( .A(sreg[429]), .B(n4262), .Z(n4264) );
  XNOR U4492 ( .A(n4263), .B(n4264), .Z(c[429]) );
  AND U4493 ( .A(b[2]), .B(a[176]), .Z(n4279) );
  AND U4494 ( .A(a[177]), .B(b[1]), .Z(n4277) );
  AND U4495 ( .A(a[175]), .B(b[3]), .Z(n4276) );
  XOR U4496 ( .A(n4277), .B(n4276), .Z(n4278) );
  XOR U4497 ( .A(n4279), .B(n4278), .Z(n4282) );
  NAND U4498 ( .A(b[0]), .B(a[178]), .Z(n4283) );
  XOR U4499 ( .A(n4282), .B(n4283), .Z(n4285) );
  OR U4500 ( .A(n4251), .B(n4250), .Z(n4255) );
  NANDN U4501 ( .A(n4253), .B(n4252), .Z(n4254) );
  NAND U4502 ( .A(n4255), .B(n4254), .Z(n4284) );
  XNOR U4503 ( .A(n4285), .B(n4284), .Z(n4270) );
  NANDN U4504 ( .A(n4257), .B(n4256), .Z(n4261) );
  OR U4505 ( .A(n4259), .B(n4258), .Z(n4260) );
  NAND U4506 ( .A(n4261), .B(n4260), .Z(n4271) );
  XNOR U4507 ( .A(n4270), .B(n4271), .Z(n4272) );
  XOR U4508 ( .A(n4273), .B(n4272), .Z(n4269) );
  OR U4509 ( .A(n4262), .B(sreg[429]), .Z(n4266) );
  NAND U4510 ( .A(n4264), .B(n4263), .Z(n4265) );
  AND U4511 ( .A(n4266), .B(n4265), .Z(n4268) );
  XNOR U4512 ( .A(sreg[430]), .B(n4268), .Z(n4267) );
  XNOR U4513 ( .A(n4269), .B(n4267), .Z(c[430]) );
  NANDN U4514 ( .A(n4271), .B(n4270), .Z(n4275) );
  NANDN U4515 ( .A(n4273), .B(n4272), .Z(n4274) );
  NAND U4516 ( .A(n4275), .B(n4274), .Z(n4291) );
  AND U4517 ( .A(b[2]), .B(a[177]), .Z(n4297) );
  AND U4518 ( .A(a[178]), .B(b[1]), .Z(n4295) );
  AND U4519 ( .A(a[176]), .B(b[3]), .Z(n4294) );
  XOR U4520 ( .A(n4295), .B(n4294), .Z(n4296) );
  XOR U4521 ( .A(n4297), .B(n4296), .Z(n4300) );
  NAND U4522 ( .A(b[0]), .B(a[179]), .Z(n4301) );
  XOR U4523 ( .A(n4300), .B(n4301), .Z(n4303) );
  OR U4524 ( .A(n4277), .B(n4276), .Z(n4281) );
  NANDN U4525 ( .A(n4279), .B(n4278), .Z(n4280) );
  NAND U4526 ( .A(n4281), .B(n4280), .Z(n4302) );
  XNOR U4527 ( .A(n4303), .B(n4302), .Z(n4288) );
  NANDN U4528 ( .A(n4283), .B(n4282), .Z(n4287) );
  OR U4529 ( .A(n4285), .B(n4284), .Z(n4286) );
  NAND U4530 ( .A(n4287), .B(n4286), .Z(n4289) );
  XNOR U4531 ( .A(n4288), .B(n4289), .Z(n4290) );
  XNOR U4532 ( .A(n4291), .B(n4290), .Z(n4307) );
  XNOR U4533 ( .A(n4307), .B(sreg[431]), .Z(n4308) );
  XOR U4534 ( .A(n4309), .B(n4308), .Z(c[431]) );
  NANDN U4535 ( .A(n4289), .B(n4288), .Z(n4293) );
  NAND U4536 ( .A(n4291), .B(n4290), .Z(n4292) );
  NAND U4537 ( .A(n4293), .B(n4292), .Z(n4319) );
  AND U4538 ( .A(b[2]), .B(a[178]), .Z(n4323) );
  AND U4539 ( .A(a[179]), .B(b[1]), .Z(n4321) );
  AND U4540 ( .A(a[177]), .B(b[3]), .Z(n4320) );
  XOR U4541 ( .A(n4321), .B(n4320), .Z(n4322) );
  XOR U4542 ( .A(n4323), .B(n4322), .Z(n4326) );
  NAND U4543 ( .A(b[0]), .B(a[180]), .Z(n4327) );
  XOR U4544 ( .A(n4326), .B(n4327), .Z(n4328) );
  OR U4545 ( .A(n4295), .B(n4294), .Z(n4299) );
  NANDN U4546 ( .A(n4297), .B(n4296), .Z(n4298) );
  AND U4547 ( .A(n4299), .B(n4298), .Z(n4329) );
  XOR U4548 ( .A(n4328), .B(n4329), .Z(n4317) );
  NANDN U4549 ( .A(n4301), .B(n4300), .Z(n4305) );
  OR U4550 ( .A(n4303), .B(n4302), .Z(n4304) );
  AND U4551 ( .A(n4305), .B(n4304), .Z(n4318) );
  XOR U4552 ( .A(n4317), .B(n4318), .Z(n4306) );
  XOR U4553 ( .A(n4319), .B(n4306), .Z(n4312) );
  XOR U4554 ( .A(sreg[432]), .B(n4312), .Z(n4314) );
  NAND U4555 ( .A(n4307), .B(sreg[431]), .Z(n4311) );
  OR U4556 ( .A(n4309), .B(n4308), .Z(n4310) );
  NAND U4557 ( .A(n4311), .B(n4310), .Z(n4313) );
  XNOR U4558 ( .A(n4314), .B(n4313), .Z(c[432]) );
  NANDN U4559 ( .A(sreg[432]), .B(n4312), .Z(n4316) );
  OR U4560 ( .A(n4314), .B(n4313), .Z(n4315) );
  AND U4561 ( .A(n4316), .B(n4315), .Z(n4331) );
  AND U4562 ( .A(b[2]), .B(a[179]), .Z(n4342) );
  AND U4563 ( .A(a[180]), .B(b[1]), .Z(n4340) );
  AND U4564 ( .A(a[178]), .B(b[3]), .Z(n4339) );
  XOR U4565 ( .A(n4340), .B(n4339), .Z(n4341) );
  XOR U4566 ( .A(n4342), .B(n4341), .Z(n4345) );
  NAND U4567 ( .A(b[0]), .B(a[181]), .Z(n4346) );
  XOR U4568 ( .A(n4345), .B(n4346), .Z(n4348) );
  OR U4569 ( .A(n4321), .B(n4320), .Z(n4325) );
  NANDN U4570 ( .A(n4323), .B(n4322), .Z(n4324) );
  NAND U4571 ( .A(n4325), .B(n4324), .Z(n4347) );
  XNOR U4572 ( .A(n4348), .B(n4347), .Z(n4333) );
  XNOR U4573 ( .A(n4333), .B(n4334), .Z(n4336) );
  XOR U4574 ( .A(n4335), .B(n4336), .Z(n4332) );
  XNOR U4575 ( .A(sreg[433]), .B(n4332), .Z(n4330) );
  XOR U4576 ( .A(n4331), .B(n4330), .Z(c[433]) );
  NANDN U4577 ( .A(n4334), .B(n4333), .Z(n4338) );
  NAND U4578 ( .A(n4336), .B(n4335), .Z(n4337) );
  NAND U4579 ( .A(n4338), .B(n4337), .Z(n4354) );
  AND U4580 ( .A(b[2]), .B(a[180]), .Z(n4360) );
  AND U4581 ( .A(a[181]), .B(b[1]), .Z(n4358) );
  AND U4582 ( .A(a[179]), .B(b[3]), .Z(n4357) );
  XOR U4583 ( .A(n4358), .B(n4357), .Z(n4359) );
  XOR U4584 ( .A(n4360), .B(n4359), .Z(n4363) );
  NAND U4585 ( .A(b[0]), .B(a[182]), .Z(n4364) );
  XOR U4586 ( .A(n4363), .B(n4364), .Z(n4366) );
  OR U4587 ( .A(n4340), .B(n4339), .Z(n4344) );
  NANDN U4588 ( .A(n4342), .B(n4341), .Z(n4343) );
  NAND U4589 ( .A(n4344), .B(n4343), .Z(n4365) );
  XNOR U4590 ( .A(n4366), .B(n4365), .Z(n4351) );
  NANDN U4591 ( .A(n4346), .B(n4345), .Z(n4350) );
  OR U4592 ( .A(n4348), .B(n4347), .Z(n4349) );
  NAND U4593 ( .A(n4350), .B(n4349), .Z(n4352) );
  XNOR U4594 ( .A(n4351), .B(n4352), .Z(n4353) );
  XNOR U4595 ( .A(n4354), .B(n4353), .Z(n4369) );
  XNOR U4596 ( .A(n4369), .B(sreg[434]), .Z(n4371) );
  XNOR U4597 ( .A(n4370), .B(n4371), .Z(c[434]) );
  NANDN U4598 ( .A(n4352), .B(n4351), .Z(n4356) );
  NAND U4599 ( .A(n4354), .B(n4353), .Z(n4355) );
  NAND U4600 ( .A(n4356), .B(n4355), .Z(n4377) );
  AND U4601 ( .A(b[2]), .B(a[181]), .Z(n4383) );
  AND U4602 ( .A(a[182]), .B(b[1]), .Z(n4381) );
  AND U4603 ( .A(a[180]), .B(b[3]), .Z(n4380) );
  XOR U4604 ( .A(n4381), .B(n4380), .Z(n4382) );
  XOR U4605 ( .A(n4383), .B(n4382), .Z(n4386) );
  NAND U4606 ( .A(b[0]), .B(a[183]), .Z(n4387) );
  XOR U4607 ( .A(n4386), .B(n4387), .Z(n4389) );
  OR U4608 ( .A(n4358), .B(n4357), .Z(n4362) );
  NANDN U4609 ( .A(n4360), .B(n4359), .Z(n4361) );
  NAND U4610 ( .A(n4362), .B(n4361), .Z(n4388) );
  XNOR U4611 ( .A(n4389), .B(n4388), .Z(n4374) );
  NANDN U4612 ( .A(n4364), .B(n4363), .Z(n4368) );
  OR U4613 ( .A(n4366), .B(n4365), .Z(n4367) );
  NAND U4614 ( .A(n4368), .B(n4367), .Z(n4375) );
  XNOR U4615 ( .A(n4374), .B(n4375), .Z(n4376) );
  XNOR U4616 ( .A(n4377), .B(n4376), .Z(n4392) );
  XOR U4617 ( .A(sreg[435]), .B(n4392), .Z(n4393) );
  NAND U4618 ( .A(n4369), .B(sreg[434]), .Z(n4373) );
  NANDN U4619 ( .A(n4371), .B(n4370), .Z(n4372) );
  NAND U4620 ( .A(n4373), .B(n4372), .Z(n4394) );
  XOR U4621 ( .A(n4393), .B(n4394), .Z(c[435]) );
  NANDN U4622 ( .A(n4375), .B(n4374), .Z(n4379) );
  NAND U4623 ( .A(n4377), .B(n4376), .Z(n4378) );
  NAND U4624 ( .A(n4379), .B(n4378), .Z(n4400) );
  AND U4625 ( .A(b[2]), .B(a[182]), .Z(n4406) );
  AND U4626 ( .A(a[183]), .B(b[1]), .Z(n4404) );
  AND U4627 ( .A(a[181]), .B(b[3]), .Z(n4403) );
  XOR U4628 ( .A(n4404), .B(n4403), .Z(n4405) );
  XOR U4629 ( .A(n4406), .B(n4405), .Z(n4409) );
  NAND U4630 ( .A(b[0]), .B(a[184]), .Z(n4410) );
  XOR U4631 ( .A(n4409), .B(n4410), .Z(n4412) );
  OR U4632 ( .A(n4381), .B(n4380), .Z(n4385) );
  NANDN U4633 ( .A(n4383), .B(n4382), .Z(n4384) );
  NAND U4634 ( .A(n4385), .B(n4384), .Z(n4411) );
  XNOR U4635 ( .A(n4412), .B(n4411), .Z(n4397) );
  NANDN U4636 ( .A(n4387), .B(n4386), .Z(n4391) );
  OR U4637 ( .A(n4389), .B(n4388), .Z(n4390) );
  NAND U4638 ( .A(n4391), .B(n4390), .Z(n4398) );
  XNOR U4639 ( .A(n4397), .B(n4398), .Z(n4399) );
  XNOR U4640 ( .A(n4400), .B(n4399), .Z(n4415) );
  XNOR U4641 ( .A(n4415), .B(sreg[436]), .Z(n4417) );
  OR U4642 ( .A(n4392), .B(sreg[435]), .Z(n4396) );
  NANDN U4643 ( .A(n4394), .B(n4393), .Z(n4395) );
  NAND U4644 ( .A(n4396), .B(n4395), .Z(n4416) );
  XOR U4645 ( .A(n4417), .B(n4416), .Z(c[436]) );
  NANDN U4646 ( .A(n4398), .B(n4397), .Z(n4402) );
  NAND U4647 ( .A(n4400), .B(n4399), .Z(n4401) );
  NAND U4648 ( .A(n4402), .B(n4401), .Z(n4428) );
  AND U4649 ( .A(b[2]), .B(a[183]), .Z(n4434) );
  AND U4650 ( .A(a[184]), .B(b[1]), .Z(n4432) );
  AND U4651 ( .A(a[182]), .B(b[3]), .Z(n4431) );
  XOR U4652 ( .A(n4432), .B(n4431), .Z(n4433) );
  XOR U4653 ( .A(n4434), .B(n4433), .Z(n4437) );
  NAND U4654 ( .A(b[0]), .B(a[185]), .Z(n4438) );
  XOR U4655 ( .A(n4437), .B(n4438), .Z(n4440) );
  OR U4656 ( .A(n4404), .B(n4403), .Z(n4408) );
  NANDN U4657 ( .A(n4406), .B(n4405), .Z(n4407) );
  NAND U4658 ( .A(n4408), .B(n4407), .Z(n4439) );
  XNOR U4659 ( .A(n4440), .B(n4439), .Z(n4425) );
  NANDN U4660 ( .A(n4410), .B(n4409), .Z(n4414) );
  OR U4661 ( .A(n4412), .B(n4411), .Z(n4413) );
  NAND U4662 ( .A(n4414), .B(n4413), .Z(n4426) );
  XNOR U4663 ( .A(n4425), .B(n4426), .Z(n4427) );
  XNOR U4664 ( .A(n4428), .B(n4427), .Z(n4420) );
  XNOR U4665 ( .A(n4420), .B(sreg[437]), .Z(n4422) );
  NAND U4666 ( .A(n4415), .B(sreg[436]), .Z(n4419) );
  OR U4667 ( .A(n4417), .B(n4416), .Z(n4418) );
  AND U4668 ( .A(n4419), .B(n4418), .Z(n4421) );
  XOR U4669 ( .A(n4422), .B(n4421), .Z(c[437]) );
  NAND U4670 ( .A(n4420), .B(sreg[437]), .Z(n4424) );
  OR U4671 ( .A(n4422), .B(n4421), .Z(n4423) );
  NAND U4672 ( .A(n4424), .B(n4423), .Z(n4463) );
  NANDN U4673 ( .A(n4426), .B(n4425), .Z(n4430) );
  NAND U4674 ( .A(n4428), .B(n4427), .Z(n4429) );
  NAND U4675 ( .A(n4430), .B(n4429), .Z(n4446) );
  AND U4676 ( .A(b[2]), .B(a[184]), .Z(n4452) );
  AND U4677 ( .A(a[185]), .B(b[1]), .Z(n4450) );
  AND U4678 ( .A(a[183]), .B(b[3]), .Z(n4449) );
  XOR U4679 ( .A(n4450), .B(n4449), .Z(n4451) );
  XOR U4680 ( .A(n4452), .B(n4451), .Z(n4455) );
  NAND U4681 ( .A(b[0]), .B(a[186]), .Z(n4456) );
  XOR U4682 ( .A(n4455), .B(n4456), .Z(n4458) );
  OR U4683 ( .A(n4432), .B(n4431), .Z(n4436) );
  NANDN U4684 ( .A(n4434), .B(n4433), .Z(n4435) );
  NAND U4685 ( .A(n4436), .B(n4435), .Z(n4457) );
  XNOR U4686 ( .A(n4458), .B(n4457), .Z(n4443) );
  NANDN U4687 ( .A(n4438), .B(n4437), .Z(n4442) );
  OR U4688 ( .A(n4440), .B(n4439), .Z(n4441) );
  NAND U4689 ( .A(n4442), .B(n4441), .Z(n4444) );
  XNOR U4690 ( .A(n4443), .B(n4444), .Z(n4445) );
  XNOR U4691 ( .A(n4446), .B(n4445), .Z(n4461) );
  XOR U4692 ( .A(sreg[438]), .B(n4461), .Z(n4462) );
  XOR U4693 ( .A(n4463), .B(n4462), .Z(c[438]) );
  NANDN U4694 ( .A(n4444), .B(n4443), .Z(n4448) );
  NAND U4695 ( .A(n4446), .B(n4445), .Z(n4447) );
  NAND U4696 ( .A(n4448), .B(n4447), .Z(n4469) );
  AND U4697 ( .A(b[2]), .B(a[185]), .Z(n4475) );
  AND U4698 ( .A(a[186]), .B(b[1]), .Z(n4473) );
  AND U4699 ( .A(a[184]), .B(b[3]), .Z(n4472) );
  XOR U4700 ( .A(n4473), .B(n4472), .Z(n4474) );
  XOR U4701 ( .A(n4475), .B(n4474), .Z(n4478) );
  NAND U4702 ( .A(b[0]), .B(a[187]), .Z(n4479) );
  XOR U4703 ( .A(n4478), .B(n4479), .Z(n4481) );
  OR U4704 ( .A(n4450), .B(n4449), .Z(n4454) );
  NANDN U4705 ( .A(n4452), .B(n4451), .Z(n4453) );
  NAND U4706 ( .A(n4454), .B(n4453), .Z(n4480) );
  XNOR U4707 ( .A(n4481), .B(n4480), .Z(n4466) );
  NANDN U4708 ( .A(n4456), .B(n4455), .Z(n4460) );
  OR U4709 ( .A(n4458), .B(n4457), .Z(n4459) );
  NAND U4710 ( .A(n4460), .B(n4459), .Z(n4467) );
  XNOR U4711 ( .A(n4466), .B(n4467), .Z(n4468) );
  XNOR U4712 ( .A(n4469), .B(n4468), .Z(n4484) );
  XNOR U4713 ( .A(n4484), .B(sreg[439]), .Z(n4486) );
  OR U4714 ( .A(n4461), .B(sreg[438]), .Z(n4465) );
  NANDN U4715 ( .A(n4463), .B(n4462), .Z(n4464) );
  NAND U4716 ( .A(n4465), .B(n4464), .Z(n4485) );
  XOR U4717 ( .A(n4486), .B(n4485), .Z(c[439]) );
  NANDN U4718 ( .A(n4467), .B(n4466), .Z(n4471) );
  NAND U4719 ( .A(n4469), .B(n4468), .Z(n4470) );
  NAND U4720 ( .A(n4471), .B(n4470), .Z(n4492) );
  AND U4721 ( .A(b[2]), .B(a[186]), .Z(n4498) );
  AND U4722 ( .A(a[187]), .B(b[1]), .Z(n4496) );
  AND U4723 ( .A(a[185]), .B(b[3]), .Z(n4495) );
  XOR U4724 ( .A(n4496), .B(n4495), .Z(n4497) );
  XOR U4725 ( .A(n4498), .B(n4497), .Z(n4501) );
  NAND U4726 ( .A(b[0]), .B(a[188]), .Z(n4502) );
  XOR U4727 ( .A(n4501), .B(n4502), .Z(n4504) );
  OR U4728 ( .A(n4473), .B(n4472), .Z(n4477) );
  NANDN U4729 ( .A(n4475), .B(n4474), .Z(n4476) );
  NAND U4730 ( .A(n4477), .B(n4476), .Z(n4503) );
  XNOR U4731 ( .A(n4504), .B(n4503), .Z(n4489) );
  NANDN U4732 ( .A(n4479), .B(n4478), .Z(n4483) );
  OR U4733 ( .A(n4481), .B(n4480), .Z(n4482) );
  NAND U4734 ( .A(n4483), .B(n4482), .Z(n4490) );
  XNOR U4735 ( .A(n4489), .B(n4490), .Z(n4491) );
  XNOR U4736 ( .A(n4492), .B(n4491), .Z(n4507) );
  XNOR U4737 ( .A(n4507), .B(sreg[440]), .Z(n4509) );
  NAND U4738 ( .A(n4484), .B(sreg[439]), .Z(n4488) );
  OR U4739 ( .A(n4486), .B(n4485), .Z(n4487) );
  AND U4740 ( .A(n4488), .B(n4487), .Z(n4508) );
  XOR U4741 ( .A(n4509), .B(n4508), .Z(c[440]) );
  NANDN U4742 ( .A(n4490), .B(n4489), .Z(n4494) );
  NAND U4743 ( .A(n4492), .B(n4491), .Z(n4493) );
  NAND U4744 ( .A(n4494), .B(n4493), .Z(n4516) );
  AND U4745 ( .A(b[2]), .B(a[187]), .Z(n4528) );
  AND U4746 ( .A(a[188]), .B(b[1]), .Z(n4526) );
  AND U4747 ( .A(a[186]), .B(b[3]), .Z(n4525) );
  XOR U4748 ( .A(n4526), .B(n4525), .Z(n4527) );
  XOR U4749 ( .A(n4528), .B(n4527), .Z(n4519) );
  NAND U4750 ( .A(b[0]), .B(a[189]), .Z(n4520) );
  XOR U4751 ( .A(n4519), .B(n4520), .Z(n4522) );
  OR U4752 ( .A(n4496), .B(n4495), .Z(n4500) );
  NANDN U4753 ( .A(n4498), .B(n4497), .Z(n4499) );
  NAND U4754 ( .A(n4500), .B(n4499), .Z(n4521) );
  XNOR U4755 ( .A(n4522), .B(n4521), .Z(n4513) );
  NANDN U4756 ( .A(n4502), .B(n4501), .Z(n4506) );
  OR U4757 ( .A(n4504), .B(n4503), .Z(n4505) );
  NAND U4758 ( .A(n4506), .B(n4505), .Z(n4514) );
  XNOR U4759 ( .A(n4513), .B(n4514), .Z(n4515) );
  XOR U4760 ( .A(n4516), .B(n4515), .Z(n4532) );
  NAND U4761 ( .A(n4507), .B(sreg[440]), .Z(n4511) );
  OR U4762 ( .A(n4509), .B(n4508), .Z(n4510) );
  NAND U4763 ( .A(n4511), .B(n4510), .Z(n4531) );
  XNOR U4764 ( .A(sreg[441]), .B(n4531), .Z(n4512) );
  XOR U4765 ( .A(n4532), .B(n4512), .Z(c[441]) );
  NANDN U4766 ( .A(n4514), .B(n4513), .Z(n4518) );
  NAND U4767 ( .A(n4516), .B(n4515), .Z(n4517) );
  NAND U4768 ( .A(n4518), .B(n4517), .Z(n4549) );
  NANDN U4769 ( .A(n4520), .B(n4519), .Z(n4524) );
  OR U4770 ( .A(n4522), .B(n4521), .Z(n4523) );
  NAND U4771 ( .A(n4524), .B(n4523), .Z(n4546) );
  AND U4772 ( .A(b[2]), .B(a[188]), .Z(n4537) );
  AND U4773 ( .A(a[189]), .B(b[1]), .Z(n4535) );
  AND U4774 ( .A(a[187]), .B(b[3]), .Z(n4534) );
  XOR U4775 ( .A(n4535), .B(n4534), .Z(n4536) );
  XOR U4776 ( .A(n4537), .B(n4536), .Z(n4540) );
  NAND U4777 ( .A(b[0]), .B(a[190]), .Z(n4541) );
  XNOR U4778 ( .A(n4540), .B(n4541), .Z(n4542) );
  OR U4779 ( .A(n4526), .B(n4525), .Z(n4530) );
  NANDN U4780 ( .A(n4528), .B(n4527), .Z(n4529) );
  AND U4781 ( .A(n4530), .B(n4529), .Z(n4543) );
  XNOR U4782 ( .A(n4542), .B(n4543), .Z(n4547) );
  XNOR U4783 ( .A(n4546), .B(n4547), .Z(n4548) );
  XNOR U4784 ( .A(n4549), .B(n4548), .Z(n4553) );
  XNOR U4785 ( .A(sreg[442]), .B(n4552), .Z(n4533) );
  XNOR U4786 ( .A(n4553), .B(n4533), .Z(c[442]) );
  AND U4787 ( .A(b[2]), .B(a[189]), .Z(n4566) );
  AND U4788 ( .A(a[190]), .B(b[1]), .Z(n4564) );
  AND U4789 ( .A(a[188]), .B(b[3]), .Z(n4563) );
  XOR U4790 ( .A(n4564), .B(n4563), .Z(n4565) );
  XOR U4791 ( .A(n4566), .B(n4565), .Z(n4569) );
  NAND U4792 ( .A(b[0]), .B(a[191]), .Z(n4570) );
  XOR U4793 ( .A(n4569), .B(n4570), .Z(n4572) );
  OR U4794 ( .A(n4535), .B(n4534), .Z(n4539) );
  NANDN U4795 ( .A(n4537), .B(n4536), .Z(n4538) );
  NAND U4796 ( .A(n4539), .B(n4538), .Z(n4571) );
  XNOR U4797 ( .A(n4572), .B(n4571), .Z(n4557) );
  NANDN U4798 ( .A(n4541), .B(n4540), .Z(n4545) );
  NAND U4799 ( .A(n4543), .B(n4542), .Z(n4544) );
  NAND U4800 ( .A(n4545), .B(n4544), .Z(n4558) );
  XNOR U4801 ( .A(n4557), .B(n4558), .Z(n4559) );
  NANDN U4802 ( .A(n4547), .B(n4546), .Z(n4551) );
  NANDN U4803 ( .A(n4549), .B(n4548), .Z(n4550) );
  NAND U4804 ( .A(n4551), .B(n4550), .Z(n4560) );
  XOR U4805 ( .A(n4559), .B(n4560), .Z(n4556) );
  XNOR U4806 ( .A(sreg[443]), .B(n4555), .Z(n4554) );
  XNOR U4807 ( .A(n4556), .B(n4554), .Z(c[443]) );
  NANDN U4808 ( .A(n4558), .B(n4557), .Z(n4562) );
  NANDN U4809 ( .A(n4560), .B(n4559), .Z(n4561) );
  NAND U4810 ( .A(n4562), .B(n4561), .Z(n4590) );
  AND U4811 ( .A(b[2]), .B(a[190]), .Z(n4584) );
  AND U4812 ( .A(a[191]), .B(b[1]), .Z(n4582) );
  AND U4813 ( .A(a[189]), .B(b[3]), .Z(n4581) );
  XOR U4814 ( .A(n4582), .B(n4581), .Z(n4583) );
  XOR U4815 ( .A(n4584), .B(n4583), .Z(n4575) );
  NAND U4816 ( .A(b[0]), .B(a[192]), .Z(n4576) );
  XOR U4817 ( .A(n4575), .B(n4576), .Z(n4578) );
  OR U4818 ( .A(n4564), .B(n4563), .Z(n4568) );
  NANDN U4819 ( .A(n4566), .B(n4565), .Z(n4567) );
  NAND U4820 ( .A(n4568), .B(n4567), .Z(n4577) );
  XNOR U4821 ( .A(n4578), .B(n4577), .Z(n4587) );
  NANDN U4822 ( .A(n4570), .B(n4569), .Z(n4574) );
  OR U4823 ( .A(n4572), .B(n4571), .Z(n4573) );
  NAND U4824 ( .A(n4574), .B(n4573), .Z(n4588) );
  XNOR U4825 ( .A(n4587), .B(n4588), .Z(n4589) );
  XNOR U4826 ( .A(n4590), .B(n4589), .Z(n4593) );
  XNOR U4827 ( .A(n4593), .B(sreg[444]), .Z(n4594) );
  XOR U4828 ( .A(n4595), .B(n4594), .Z(c[444]) );
  NANDN U4829 ( .A(n4576), .B(n4575), .Z(n4580) );
  OR U4830 ( .A(n4578), .B(n4577), .Z(n4579) );
  NAND U4831 ( .A(n4580), .B(n4579), .Z(n4610) );
  AND U4832 ( .A(b[2]), .B(a[191]), .Z(n4601) );
  AND U4833 ( .A(a[192]), .B(b[1]), .Z(n4599) );
  AND U4834 ( .A(a[190]), .B(b[3]), .Z(n4598) );
  XOR U4835 ( .A(n4599), .B(n4598), .Z(n4600) );
  XOR U4836 ( .A(n4601), .B(n4600), .Z(n4604) );
  NAND U4837 ( .A(b[0]), .B(a[193]), .Z(n4605) );
  XNOR U4838 ( .A(n4604), .B(n4605), .Z(n4606) );
  OR U4839 ( .A(n4582), .B(n4581), .Z(n4586) );
  NANDN U4840 ( .A(n4584), .B(n4583), .Z(n4585) );
  AND U4841 ( .A(n4586), .B(n4585), .Z(n4607) );
  XNOR U4842 ( .A(n4606), .B(n4607), .Z(n4611) );
  XNOR U4843 ( .A(n4610), .B(n4611), .Z(n4612) );
  NANDN U4844 ( .A(n4588), .B(n4587), .Z(n4592) );
  NAND U4845 ( .A(n4590), .B(n4589), .Z(n4591) );
  NAND U4846 ( .A(n4592), .B(n4591), .Z(n4613) );
  XNOR U4847 ( .A(n4612), .B(n4613), .Z(n4616) );
  XOR U4848 ( .A(sreg[445]), .B(n4616), .Z(n4617) );
  NAND U4849 ( .A(n4593), .B(sreg[444]), .Z(n4597) );
  OR U4850 ( .A(n4595), .B(n4594), .Z(n4596) );
  NAND U4851 ( .A(n4597), .B(n4596), .Z(n4618) );
  XOR U4852 ( .A(n4617), .B(n4618), .Z(c[445]) );
  AND U4853 ( .A(b[2]), .B(a[192]), .Z(n4630) );
  AND U4854 ( .A(a[193]), .B(b[1]), .Z(n4628) );
  AND U4855 ( .A(a[191]), .B(b[3]), .Z(n4627) );
  XOR U4856 ( .A(n4628), .B(n4627), .Z(n4629) );
  XOR U4857 ( .A(n4630), .B(n4629), .Z(n4633) );
  NAND U4858 ( .A(b[0]), .B(a[194]), .Z(n4634) );
  XOR U4859 ( .A(n4633), .B(n4634), .Z(n4636) );
  OR U4860 ( .A(n4599), .B(n4598), .Z(n4603) );
  NANDN U4861 ( .A(n4601), .B(n4600), .Z(n4602) );
  NAND U4862 ( .A(n4603), .B(n4602), .Z(n4635) );
  XNOR U4863 ( .A(n4636), .B(n4635), .Z(n4621) );
  NANDN U4864 ( .A(n4605), .B(n4604), .Z(n4609) );
  NAND U4865 ( .A(n4607), .B(n4606), .Z(n4608) );
  NAND U4866 ( .A(n4609), .B(n4608), .Z(n4622) );
  XNOR U4867 ( .A(n4621), .B(n4622), .Z(n4623) );
  NANDN U4868 ( .A(n4611), .B(n4610), .Z(n4615) );
  NANDN U4869 ( .A(n4613), .B(n4612), .Z(n4614) );
  AND U4870 ( .A(n4615), .B(n4614), .Z(n4624) );
  XNOR U4871 ( .A(n4623), .B(n4624), .Z(n4639) );
  XOR U4872 ( .A(sreg[446]), .B(n4639), .Z(n4640) );
  OR U4873 ( .A(n4616), .B(sreg[445]), .Z(n4620) );
  NANDN U4874 ( .A(n4618), .B(n4617), .Z(n4619) );
  AND U4875 ( .A(n4620), .B(n4619), .Z(n4641) );
  XOR U4876 ( .A(n4640), .B(n4641), .Z(c[446]) );
  NANDN U4877 ( .A(n4622), .B(n4621), .Z(n4626) );
  NAND U4878 ( .A(n4624), .B(n4623), .Z(n4625) );
  NAND U4879 ( .A(n4626), .B(n4625), .Z(n4650) );
  AND U4880 ( .A(b[2]), .B(a[193]), .Z(n4656) );
  AND U4881 ( .A(a[194]), .B(b[1]), .Z(n4654) );
  AND U4882 ( .A(a[192]), .B(b[3]), .Z(n4653) );
  XOR U4883 ( .A(n4654), .B(n4653), .Z(n4655) );
  XOR U4884 ( .A(n4656), .B(n4655), .Z(n4659) );
  NAND U4885 ( .A(b[0]), .B(a[195]), .Z(n4660) );
  XOR U4886 ( .A(n4659), .B(n4660), .Z(n4662) );
  OR U4887 ( .A(n4628), .B(n4627), .Z(n4632) );
  NANDN U4888 ( .A(n4630), .B(n4629), .Z(n4631) );
  NAND U4889 ( .A(n4632), .B(n4631), .Z(n4661) );
  XNOR U4890 ( .A(n4662), .B(n4661), .Z(n4647) );
  NANDN U4891 ( .A(n4634), .B(n4633), .Z(n4638) );
  OR U4892 ( .A(n4636), .B(n4635), .Z(n4637) );
  NAND U4893 ( .A(n4638), .B(n4637), .Z(n4648) );
  XNOR U4894 ( .A(n4647), .B(n4648), .Z(n4649) );
  XOR U4895 ( .A(n4650), .B(n4649), .Z(n4646) );
  OR U4896 ( .A(n4639), .B(sreg[446]), .Z(n4643) );
  NANDN U4897 ( .A(n4641), .B(n4640), .Z(n4642) );
  AND U4898 ( .A(n4643), .B(n4642), .Z(n4645) );
  XNOR U4899 ( .A(sreg[447]), .B(n4645), .Z(n4644) );
  XOR U4900 ( .A(n4646), .B(n4644), .Z(c[447]) );
  NANDN U4901 ( .A(n4648), .B(n4647), .Z(n4652) );
  NAND U4902 ( .A(n4650), .B(n4649), .Z(n4651) );
  NAND U4903 ( .A(n4652), .B(n4651), .Z(n4668) );
  AND U4904 ( .A(b[2]), .B(a[194]), .Z(n4680) );
  AND U4905 ( .A(a[195]), .B(b[1]), .Z(n4678) );
  AND U4906 ( .A(a[193]), .B(b[3]), .Z(n4677) );
  XOR U4907 ( .A(n4678), .B(n4677), .Z(n4679) );
  XOR U4908 ( .A(n4680), .B(n4679), .Z(n4671) );
  NAND U4909 ( .A(b[0]), .B(a[196]), .Z(n4672) );
  XOR U4910 ( .A(n4671), .B(n4672), .Z(n4674) );
  OR U4911 ( .A(n4654), .B(n4653), .Z(n4658) );
  NANDN U4912 ( .A(n4656), .B(n4655), .Z(n4657) );
  NAND U4913 ( .A(n4658), .B(n4657), .Z(n4673) );
  XNOR U4914 ( .A(n4674), .B(n4673), .Z(n4665) );
  NANDN U4915 ( .A(n4660), .B(n4659), .Z(n4664) );
  OR U4916 ( .A(n4662), .B(n4661), .Z(n4663) );
  NAND U4917 ( .A(n4664), .B(n4663), .Z(n4666) );
  XNOR U4918 ( .A(n4665), .B(n4666), .Z(n4667) );
  XNOR U4919 ( .A(n4668), .B(n4667), .Z(n4683) );
  XOR U4920 ( .A(sreg[448]), .B(n4683), .Z(n4685) );
  XNOR U4921 ( .A(n4684), .B(n4685), .Z(c[448]) );
  NANDN U4922 ( .A(n4666), .B(n4665), .Z(n4670) );
  NAND U4923 ( .A(n4668), .B(n4667), .Z(n4669) );
  NAND U4924 ( .A(n4670), .B(n4669), .Z(n4704) );
  NANDN U4925 ( .A(n4672), .B(n4671), .Z(n4676) );
  OR U4926 ( .A(n4674), .B(n4673), .Z(n4675) );
  NAND U4927 ( .A(n4676), .B(n4675), .Z(n4701) );
  AND U4928 ( .A(b[2]), .B(a[195]), .Z(n4692) );
  AND U4929 ( .A(a[196]), .B(b[1]), .Z(n4690) );
  AND U4930 ( .A(a[194]), .B(b[3]), .Z(n4689) );
  XOR U4931 ( .A(n4690), .B(n4689), .Z(n4691) );
  XOR U4932 ( .A(n4692), .B(n4691), .Z(n4695) );
  NAND U4933 ( .A(b[0]), .B(a[197]), .Z(n4696) );
  XNOR U4934 ( .A(n4695), .B(n4696), .Z(n4697) );
  OR U4935 ( .A(n4678), .B(n4677), .Z(n4682) );
  NANDN U4936 ( .A(n4680), .B(n4679), .Z(n4681) );
  AND U4937 ( .A(n4682), .B(n4681), .Z(n4698) );
  XNOR U4938 ( .A(n4697), .B(n4698), .Z(n4702) );
  XNOR U4939 ( .A(n4701), .B(n4702), .Z(n4703) );
  XOR U4940 ( .A(n4704), .B(n4703), .Z(n4708) );
  OR U4941 ( .A(n4683), .B(sreg[448]), .Z(n4687) );
  NAND U4942 ( .A(n4685), .B(n4684), .Z(n4686) );
  AND U4943 ( .A(n4687), .B(n4686), .Z(n4707) );
  XOR U4944 ( .A(sreg[449]), .B(n4707), .Z(n4688) );
  XNOR U4945 ( .A(n4708), .B(n4688), .Z(c[449]) );
  AND U4946 ( .A(b[2]), .B(a[196]), .Z(n4721) );
  AND U4947 ( .A(a[197]), .B(b[1]), .Z(n4719) );
  AND U4948 ( .A(a[195]), .B(b[3]), .Z(n4718) );
  XOR U4949 ( .A(n4719), .B(n4718), .Z(n4720) );
  XOR U4950 ( .A(n4721), .B(n4720), .Z(n4724) );
  NAND U4951 ( .A(b[0]), .B(a[198]), .Z(n4725) );
  XOR U4952 ( .A(n4724), .B(n4725), .Z(n4727) );
  OR U4953 ( .A(n4690), .B(n4689), .Z(n4694) );
  NANDN U4954 ( .A(n4692), .B(n4691), .Z(n4693) );
  NAND U4955 ( .A(n4694), .B(n4693), .Z(n4726) );
  XNOR U4956 ( .A(n4727), .B(n4726), .Z(n4712) );
  NANDN U4957 ( .A(n4696), .B(n4695), .Z(n4700) );
  NAND U4958 ( .A(n4698), .B(n4697), .Z(n4699) );
  NAND U4959 ( .A(n4700), .B(n4699), .Z(n4713) );
  XNOR U4960 ( .A(n4712), .B(n4713), .Z(n4714) );
  NANDN U4961 ( .A(n4702), .B(n4701), .Z(n4706) );
  NANDN U4962 ( .A(n4704), .B(n4703), .Z(n4705) );
  NAND U4963 ( .A(n4706), .B(n4705), .Z(n4715) );
  XOR U4964 ( .A(n4714), .B(n4715), .Z(n4711) );
  XOR U4965 ( .A(sreg[450]), .B(n4710), .Z(n4709) );
  XNOR U4966 ( .A(n4711), .B(n4709), .Z(c[450]) );
  NANDN U4967 ( .A(n4713), .B(n4712), .Z(n4717) );
  NANDN U4968 ( .A(n4715), .B(n4714), .Z(n4716) );
  NAND U4969 ( .A(n4717), .B(n4716), .Z(n4750) );
  AND U4970 ( .A(b[2]), .B(a[197]), .Z(n4744) );
  AND U4971 ( .A(a[198]), .B(b[1]), .Z(n4742) );
  AND U4972 ( .A(a[196]), .B(b[3]), .Z(n4741) );
  XOR U4973 ( .A(n4742), .B(n4741), .Z(n4743) );
  XOR U4974 ( .A(n4744), .B(n4743), .Z(n4735) );
  NAND U4975 ( .A(b[0]), .B(a[199]), .Z(n4736) );
  XOR U4976 ( .A(n4735), .B(n4736), .Z(n4738) );
  OR U4977 ( .A(n4719), .B(n4718), .Z(n4723) );
  NANDN U4978 ( .A(n4721), .B(n4720), .Z(n4722) );
  NAND U4979 ( .A(n4723), .B(n4722), .Z(n4737) );
  XNOR U4980 ( .A(n4738), .B(n4737), .Z(n4747) );
  NANDN U4981 ( .A(n4725), .B(n4724), .Z(n4729) );
  OR U4982 ( .A(n4727), .B(n4726), .Z(n4728) );
  NAND U4983 ( .A(n4729), .B(n4728), .Z(n4748) );
  XNOR U4984 ( .A(n4747), .B(n4748), .Z(n4749) );
  XNOR U4985 ( .A(n4750), .B(n4749), .Z(n4730) );
  XNOR U4986 ( .A(n4730), .B(sreg[451]), .Z(n4731) );
  XOR U4987 ( .A(n4732), .B(n4731), .Z(c[451]) );
  NAND U4988 ( .A(n4730), .B(sreg[451]), .Z(n4734) );
  OR U4989 ( .A(n4732), .B(n4731), .Z(n4733) );
  AND U4990 ( .A(n4734), .B(n4733), .Z(n4773) );
  NANDN U4991 ( .A(n4736), .B(n4735), .Z(n4740) );
  OR U4992 ( .A(n4738), .B(n4737), .Z(n4739) );
  NAND U4993 ( .A(n4740), .B(n4739), .Z(n4766) );
  AND U4994 ( .A(b[2]), .B(a[198]), .Z(n4757) );
  AND U4995 ( .A(a[199]), .B(b[1]), .Z(n4755) );
  AND U4996 ( .A(a[197]), .B(b[3]), .Z(n4754) );
  XOR U4997 ( .A(n4755), .B(n4754), .Z(n4756) );
  XOR U4998 ( .A(n4757), .B(n4756), .Z(n4760) );
  NAND U4999 ( .A(b[0]), .B(a[200]), .Z(n4761) );
  XNOR U5000 ( .A(n4760), .B(n4761), .Z(n4762) );
  OR U5001 ( .A(n4742), .B(n4741), .Z(n4746) );
  NANDN U5002 ( .A(n4744), .B(n4743), .Z(n4745) );
  AND U5003 ( .A(n4746), .B(n4745), .Z(n4763) );
  XNOR U5004 ( .A(n4762), .B(n4763), .Z(n4767) );
  XNOR U5005 ( .A(n4766), .B(n4767), .Z(n4768) );
  NANDN U5006 ( .A(n4748), .B(n4747), .Z(n4752) );
  NAND U5007 ( .A(n4750), .B(n4749), .Z(n4751) );
  AND U5008 ( .A(n4752), .B(n4751), .Z(n4769) );
  XOR U5009 ( .A(n4768), .B(n4769), .Z(n4772) );
  XNOR U5010 ( .A(sreg[452]), .B(n4772), .Z(n4753) );
  XOR U5011 ( .A(n4773), .B(n4753), .Z(c[452]) );
  AND U5012 ( .A(b[2]), .B(a[199]), .Z(n4786) );
  AND U5013 ( .A(a[200]), .B(b[1]), .Z(n4784) );
  AND U5014 ( .A(a[198]), .B(b[3]), .Z(n4783) );
  XOR U5015 ( .A(n4784), .B(n4783), .Z(n4785) );
  XOR U5016 ( .A(n4786), .B(n4785), .Z(n4789) );
  NAND U5017 ( .A(b[0]), .B(a[201]), .Z(n4790) );
  XOR U5018 ( .A(n4789), .B(n4790), .Z(n4792) );
  OR U5019 ( .A(n4755), .B(n4754), .Z(n4759) );
  NANDN U5020 ( .A(n4757), .B(n4756), .Z(n4758) );
  NAND U5021 ( .A(n4759), .B(n4758), .Z(n4791) );
  XNOR U5022 ( .A(n4792), .B(n4791), .Z(n4777) );
  NANDN U5023 ( .A(n4761), .B(n4760), .Z(n4765) );
  NAND U5024 ( .A(n4763), .B(n4762), .Z(n4764) );
  NAND U5025 ( .A(n4765), .B(n4764), .Z(n4778) );
  XNOR U5026 ( .A(n4777), .B(n4778), .Z(n4779) );
  NANDN U5027 ( .A(n4767), .B(n4766), .Z(n4771) );
  NAND U5028 ( .A(n4769), .B(n4768), .Z(n4770) );
  NAND U5029 ( .A(n4771), .B(n4770), .Z(n4780) );
  XOR U5030 ( .A(n4779), .B(n4780), .Z(n4776) );
  XNOR U5031 ( .A(sreg[453]), .B(n4775), .Z(n4774) );
  XNOR U5032 ( .A(n4776), .B(n4774), .Z(c[453]) );
  NANDN U5033 ( .A(n4778), .B(n4777), .Z(n4782) );
  NANDN U5034 ( .A(n4780), .B(n4779), .Z(n4781) );
  NAND U5035 ( .A(n4782), .B(n4781), .Z(n4815) );
  AND U5036 ( .A(b[2]), .B(a[200]), .Z(n4809) );
  AND U5037 ( .A(a[201]), .B(b[1]), .Z(n4807) );
  AND U5038 ( .A(a[199]), .B(b[3]), .Z(n4806) );
  XOR U5039 ( .A(n4807), .B(n4806), .Z(n4808) );
  XOR U5040 ( .A(n4809), .B(n4808), .Z(n4800) );
  NAND U5041 ( .A(b[0]), .B(a[202]), .Z(n4801) );
  XOR U5042 ( .A(n4800), .B(n4801), .Z(n4803) );
  OR U5043 ( .A(n4784), .B(n4783), .Z(n4788) );
  NANDN U5044 ( .A(n4786), .B(n4785), .Z(n4787) );
  NAND U5045 ( .A(n4788), .B(n4787), .Z(n4802) );
  XNOR U5046 ( .A(n4803), .B(n4802), .Z(n4812) );
  NANDN U5047 ( .A(n4790), .B(n4789), .Z(n4794) );
  OR U5048 ( .A(n4792), .B(n4791), .Z(n4793) );
  NAND U5049 ( .A(n4794), .B(n4793), .Z(n4813) );
  XNOR U5050 ( .A(n4812), .B(n4813), .Z(n4814) );
  XNOR U5051 ( .A(n4815), .B(n4814), .Z(n4795) );
  XNOR U5052 ( .A(n4795), .B(sreg[454]), .Z(n4796) );
  XOR U5053 ( .A(n4797), .B(n4796), .Z(c[454]) );
  NAND U5054 ( .A(n4795), .B(sreg[454]), .Z(n4799) );
  OR U5055 ( .A(n4797), .B(n4796), .Z(n4798) );
  NAND U5056 ( .A(n4799), .B(n4798), .Z(n4837) );
  NANDN U5057 ( .A(n4801), .B(n4800), .Z(n4805) );
  OR U5058 ( .A(n4803), .B(n4802), .Z(n4804) );
  NAND U5059 ( .A(n4805), .B(n4804), .Z(n4831) );
  AND U5060 ( .A(b[2]), .B(a[201]), .Z(n4822) );
  AND U5061 ( .A(a[202]), .B(b[1]), .Z(n4820) );
  AND U5062 ( .A(a[200]), .B(b[3]), .Z(n4819) );
  XOR U5063 ( .A(n4820), .B(n4819), .Z(n4821) );
  XOR U5064 ( .A(n4822), .B(n4821), .Z(n4825) );
  NAND U5065 ( .A(b[0]), .B(a[203]), .Z(n4826) );
  XNOR U5066 ( .A(n4825), .B(n4826), .Z(n4827) );
  OR U5067 ( .A(n4807), .B(n4806), .Z(n4811) );
  NANDN U5068 ( .A(n4809), .B(n4808), .Z(n4810) );
  AND U5069 ( .A(n4811), .B(n4810), .Z(n4828) );
  XNOR U5070 ( .A(n4827), .B(n4828), .Z(n4832) );
  XNOR U5071 ( .A(n4831), .B(n4832), .Z(n4833) );
  NANDN U5072 ( .A(n4813), .B(n4812), .Z(n4817) );
  NAND U5073 ( .A(n4815), .B(n4814), .Z(n4816) );
  AND U5074 ( .A(n4817), .B(n4816), .Z(n4834) );
  XNOR U5075 ( .A(n4833), .B(n4834), .Z(n4838) );
  XOR U5076 ( .A(sreg[455]), .B(n4838), .Z(n4818) );
  XNOR U5077 ( .A(n4837), .B(n4818), .Z(c[455]) );
  AND U5078 ( .A(b[2]), .B(a[202]), .Z(n4851) );
  AND U5079 ( .A(a[203]), .B(b[1]), .Z(n4849) );
  AND U5080 ( .A(a[201]), .B(b[3]), .Z(n4848) );
  XOR U5081 ( .A(n4849), .B(n4848), .Z(n4850) );
  XOR U5082 ( .A(n4851), .B(n4850), .Z(n4854) );
  NAND U5083 ( .A(b[0]), .B(a[204]), .Z(n4855) );
  XOR U5084 ( .A(n4854), .B(n4855), .Z(n4857) );
  OR U5085 ( .A(n4820), .B(n4819), .Z(n4824) );
  NANDN U5086 ( .A(n4822), .B(n4821), .Z(n4823) );
  NAND U5087 ( .A(n4824), .B(n4823), .Z(n4856) );
  XNOR U5088 ( .A(n4857), .B(n4856), .Z(n4842) );
  NANDN U5089 ( .A(n4826), .B(n4825), .Z(n4830) );
  NAND U5090 ( .A(n4828), .B(n4827), .Z(n4829) );
  NAND U5091 ( .A(n4830), .B(n4829), .Z(n4843) );
  XNOR U5092 ( .A(n4842), .B(n4843), .Z(n4844) );
  NANDN U5093 ( .A(n4832), .B(n4831), .Z(n4836) );
  NAND U5094 ( .A(n4834), .B(n4833), .Z(n4835) );
  AND U5095 ( .A(n4836), .B(n4835), .Z(n4845) );
  XNOR U5096 ( .A(n4844), .B(n4845), .Z(n4841) );
  XNOR U5097 ( .A(sreg[456]), .B(n4840), .Z(n4839) );
  XOR U5098 ( .A(n4841), .B(n4839), .Z(c[456]) );
  NANDN U5099 ( .A(n4843), .B(n4842), .Z(n4847) );
  NAND U5100 ( .A(n4845), .B(n4844), .Z(n4846) );
  NAND U5101 ( .A(n4847), .B(n4846), .Z(n4875) );
  AND U5102 ( .A(b[2]), .B(a[203]), .Z(n4869) );
  AND U5103 ( .A(a[204]), .B(b[1]), .Z(n4867) );
  AND U5104 ( .A(a[202]), .B(b[3]), .Z(n4866) );
  XOR U5105 ( .A(n4867), .B(n4866), .Z(n4868) );
  XOR U5106 ( .A(n4869), .B(n4868), .Z(n4860) );
  NAND U5107 ( .A(b[0]), .B(a[205]), .Z(n4861) );
  XOR U5108 ( .A(n4860), .B(n4861), .Z(n4863) );
  OR U5109 ( .A(n4849), .B(n4848), .Z(n4853) );
  NANDN U5110 ( .A(n4851), .B(n4850), .Z(n4852) );
  NAND U5111 ( .A(n4853), .B(n4852), .Z(n4862) );
  XNOR U5112 ( .A(n4863), .B(n4862), .Z(n4872) );
  NANDN U5113 ( .A(n4855), .B(n4854), .Z(n4859) );
  OR U5114 ( .A(n4857), .B(n4856), .Z(n4858) );
  NAND U5115 ( .A(n4859), .B(n4858), .Z(n4873) );
  XNOR U5116 ( .A(n4872), .B(n4873), .Z(n4874) );
  XNOR U5117 ( .A(n4875), .B(n4874), .Z(n4878) );
  XNOR U5118 ( .A(n4878), .B(sreg[457]), .Z(n4879) );
  XOR U5119 ( .A(n4880), .B(n4879), .Z(c[457]) );
  NANDN U5120 ( .A(n4861), .B(n4860), .Z(n4865) );
  OR U5121 ( .A(n4863), .B(n4862), .Z(n4864) );
  NAND U5122 ( .A(n4865), .B(n4864), .Z(n4898) );
  AND U5123 ( .A(b[2]), .B(a[204]), .Z(n4889) );
  AND U5124 ( .A(a[205]), .B(b[1]), .Z(n4887) );
  AND U5125 ( .A(a[203]), .B(b[3]), .Z(n4886) );
  XOR U5126 ( .A(n4887), .B(n4886), .Z(n4888) );
  XOR U5127 ( .A(n4889), .B(n4888), .Z(n4892) );
  NAND U5128 ( .A(b[0]), .B(a[206]), .Z(n4893) );
  XNOR U5129 ( .A(n4892), .B(n4893), .Z(n4894) );
  OR U5130 ( .A(n4867), .B(n4866), .Z(n4871) );
  NANDN U5131 ( .A(n4869), .B(n4868), .Z(n4870) );
  AND U5132 ( .A(n4871), .B(n4870), .Z(n4895) );
  XNOR U5133 ( .A(n4894), .B(n4895), .Z(n4899) );
  XNOR U5134 ( .A(n4898), .B(n4899), .Z(n4900) );
  NANDN U5135 ( .A(n4873), .B(n4872), .Z(n4877) );
  NAND U5136 ( .A(n4875), .B(n4874), .Z(n4876) );
  NAND U5137 ( .A(n4877), .B(n4876), .Z(n4901) );
  XOR U5138 ( .A(n4900), .B(n4901), .Z(n4885) );
  NAND U5139 ( .A(n4878), .B(sreg[457]), .Z(n4882) );
  OR U5140 ( .A(n4880), .B(n4879), .Z(n4881) );
  AND U5141 ( .A(n4882), .B(n4881), .Z(n4884) );
  XNOR U5142 ( .A(n4884), .B(sreg[458]), .Z(n4883) );
  XNOR U5143 ( .A(n4885), .B(n4883), .Z(c[458]) );
  AND U5144 ( .A(b[2]), .B(a[205]), .Z(n4913) );
  AND U5145 ( .A(a[206]), .B(b[1]), .Z(n4911) );
  AND U5146 ( .A(a[204]), .B(b[3]), .Z(n4910) );
  XOR U5147 ( .A(n4911), .B(n4910), .Z(n4912) );
  XOR U5148 ( .A(n4913), .B(n4912), .Z(n4916) );
  NAND U5149 ( .A(b[0]), .B(a[207]), .Z(n4917) );
  XOR U5150 ( .A(n4916), .B(n4917), .Z(n4919) );
  OR U5151 ( .A(n4887), .B(n4886), .Z(n4891) );
  NANDN U5152 ( .A(n4889), .B(n4888), .Z(n4890) );
  NAND U5153 ( .A(n4891), .B(n4890), .Z(n4918) );
  XNOR U5154 ( .A(n4919), .B(n4918), .Z(n4904) );
  NANDN U5155 ( .A(n4893), .B(n4892), .Z(n4897) );
  NAND U5156 ( .A(n4895), .B(n4894), .Z(n4896) );
  NAND U5157 ( .A(n4897), .B(n4896), .Z(n4905) );
  XNOR U5158 ( .A(n4904), .B(n4905), .Z(n4906) );
  NANDN U5159 ( .A(n4899), .B(n4898), .Z(n4903) );
  NANDN U5160 ( .A(n4901), .B(n4900), .Z(n4902) );
  NAND U5161 ( .A(n4903), .B(n4902), .Z(n4907) );
  XOR U5162 ( .A(n4906), .B(n4907), .Z(n4922) );
  XNOR U5163 ( .A(n4922), .B(sreg[459]), .Z(n4924) );
  XNOR U5164 ( .A(n4923), .B(n4924), .Z(c[459]) );
  NANDN U5165 ( .A(n4905), .B(n4904), .Z(n4909) );
  NANDN U5166 ( .A(n4907), .B(n4906), .Z(n4908) );
  NAND U5167 ( .A(n4909), .B(n4908), .Z(n4945) );
  AND U5168 ( .A(b[2]), .B(a[206]), .Z(n4939) );
  AND U5169 ( .A(a[207]), .B(b[1]), .Z(n4937) );
  AND U5170 ( .A(a[205]), .B(b[3]), .Z(n4936) );
  XOR U5171 ( .A(n4937), .B(n4936), .Z(n4938) );
  XOR U5172 ( .A(n4939), .B(n4938), .Z(n4930) );
  NAND U5173 ( .A(b[0]), .B(a[208]), .Z(n4931) );
  XOR U5174 ( .A(n4930), .B(n4931), .Z(n4933) );
  OR U5175 ( .A(n4911), .B(n4910), .Z(n4915) );
  NANDN U5176 ( .A(n4913), .B(n4912), .Z(n4914) );
  NAND U5177 ( .A(n4915), .B(n4914), .Z(n4932) );
  XNOR U5178 ( .A(n4933), .B(n4932), .Z(n4942) );
  NANDN U5179 ( .A(n4917), .B(n4916), .Z(n4921) );
  OR U5180 ( .A(n4919), .B(n4918), .Z(n4920) );
  NAND U5181 ( .A(n4921), .B(n4920), .Z(n4943) );
  XNOR U5182 ( .A(n4942), .B(n4943), .Z(n4944) );
  XOR U5183 ( .A(n4945), .B(n4944), .Z(n4929) );
  NAND U5184 ( .A(n4922), .B(sreg[459]), .Z(n4926) );
  NANDN U5185 ( .A(n4924), .B(n4923), .Z(n4925) );
  NAND U5186 ( .A(n4926), .B(n4925), .Z(n4928) );
  XNOR U5187 ( .A(sreg[460]), .B(n4928), .Z(n4927) );
  XOR U5188 ( .A(n4929), .B(n4927), .Z(c[460]) );
  NANDN U5189 ( .A(n4931), .B(n4930), .Z(n4935) );
  OR U5190 ( .A(n4933), .B(n4932), .Z(n4934) );
  NAND U5191 ( .A(n4935), .B(n4934), .Z(n4948) );
  AND U5192 ( .A(b[2]), .B(a[207]), .Z(n4957) );
  AND U5193 ( .A(a[208]), .B(b[1]), .Z(n4955) );
  AND U5194 ( .A(a[206]), .B(b[3]), .Z(n4954) );
  XOR U5195 ( .A(n4955), .B(n4954), .Z(n4956) );
  XOR U5196 ( .A(n4957), .B(n4956), .Z(n4960) );
  NAND U5197 ( .A(b[0]), .B(a[209]), .Z(n4961) );
  XNOR U5198 ( .A(n4960), .B(n4961), .Z(n4962) );
  OR U5199 ( .A(n4937), .B(n4936), .Z(n4941) );
  NANDN U5200 ( .A(n4939), .B(n4938), .Z(n4940) );
  AND U5201 ( .A(n4941), .B(n4940), .Z(n4963) );
  XNOR U5202 ( .A(n4962), .B(n4963), .Z(n4949) );
  XNOR U5203 ( .A(n4948), .B(n4949), .Z(n4950) );
  NANDN U5204 ( .A(n4943), .B(n4942), .Z(n4947) );
  NAND U5205 ( .A(n4945), .B(n4944), .Z(n4946) );
  AND U5206 ( .A(n4947), .B(n4946), .Z(n4951) );
  XOR U5207 ( .A(n4950), .B(n4951), .Z(n4966) );
  XNOR U5208 ( .A(sreg[461]), .B(n4966), .Z(n4967) );
  XOR U5209 ( .A(n4968), .B(n4967), .Z(c[461]) );
  NANDN U5210 ( .A(n4949), .B(n4948), .Z(n4953) );
  NAND U5211 ( .A(n4951), .B(n4950), .Z(n4952) );
  NAND U5212 ( .A(n4953), .B(n4952), .Z(n4977) );
  AND U5213 ( .A(b[2]), .B(a[208]), .Z(n4983) );
  AND U5214 ( .A(a[209]), .B(b[1]), .Z(n4981) );
  AND U5215 ( .A(a[207]), .B(b[3]), .Z(n4980) );
  XOR U5216 ( .A(n4981), .B(n4980), .Z(n4982) );
  XOR U5217 ( .A(n4983), .B(n4982), .Z(n4986) );
  NAND U5218 ( .A(b[0]), .B(a[210]), .Z(n4987) );
  XOR U5219 ( .A(n4986), .B(n4987), .Z(n4989) );
  OR U5220 ( .A(n4955), .B(n4954), .Z(n4959) );
  NANDN U5221 ( .A(n4957), .B(n4956), .Z(n4958) );
  NAND U5222 ( .A(n4959), .B(n4958), .Z(n4988) );
  XNOR U5223 ( .A(n4989), .B(n4988), .Z(n4974) );
  NANDN U5224 ( .A(n4961), .B(n4960), .Z(n4965) );
  NAND U5225 ( .A(n4963), .B(n4962), .Z(n4964) );
  NAND U5226 ( .A(n4965), .B(n4964), .Z(n4975) );
  XNOR U5227 ( .A(n4974), .B(n4975), .Z(n4976) );
  XOR U5228 ( .A(n4977), .B(n4976), .Z(n4973) );
  NAND U5229 ( .A(sreg[461]), .B(n4966), .Z(n4970) );
  OR U5230 ( .A(n4968), .B(n4967), .Z(n4969) );
  NAND U5231 ( .A(n4970), .B(n4969), .Z(n4972) );
  XNOR U5232 ( .A(sreg[462]), .B(n4972), .Z(n4971) );
  XNOR U5233 ( .A(n4973), .B(n4971), .Z(c[462]) );
  NANDN U5234 ( .A(n4975), .B(n4974), .Z(n4979) );
  NANDN U5235 ( .A(n4977), .B(n4976), .Z(n4978) );
  NAND U5236 ( .A(n4979), .B(n4978), .Z(n4995) );
  AND U5237 ( .A(b[2]), .B(a[209]), .Z(n5001) );
  AND U5238 ( .A(a[210]), .B(b[1]), .Z(n4999) );
  AND U5239 ( .A(a[208]), .B(b[3]), .Z(n4998) );
  XOR U5240 ( .A(n4999), .B(n4998), .Z(n5000) );
  XOR U5241 ( .A(n5001), .B(n5000), .Z(n5004) );
  NAND U5242 ( .A(b[0]), .B(a[211]), .Z(n5005) );
  XOR U5243 ( .A(n5004), .B(n5005), .Z(n5007) );
  OR U5244 ( .A(n4981), .B(n4980), .Z(n4985) );
  NANDN U5245 ( .A(n4983), .B(n4982), .Z(n4984) );
  NAND U5246 ( .A(n4985), .B(n4984), .Z(n5006) );
  XNOR U5247 ( .A(n5007), .B(n5006), .Z(n4992) );
  NANDN U5248 ( .A(n4987), .B(n4986), .Z(n4991) );
  OR U5249 ( .A(n4989), .B(n4988), .Z(n4990) );
  NAND U5250 ( .A(n4991), .B(n4990), .Z(n4993) );
  XNOR U5251 ( .A(n4992), .B(n4993), .Z(n4994) );
  XNOR U5252 ( .A(n4995), .B(n4994), .Z(n5010) );
  XNOR U5253 ( .A(n5010), .B(sreg[463]), .Z(n5011) );
  XOR U5254 ( .A(n5012), .B(n5011), .Z(c[463]) );
  NANDN U5255 ( .A(n4993), .B(n4992), .Z(n4997) );
  NAND U5256 ( .A(n4995), .B(n4994), .Z(n4996) );
  NAND U5257 ( .A(n4997), .B(n4996), .Z(n5018) );
  AND U5258 ( .A(b[2]), .B(a[210]), .Z(n5024) );
  AND U5259 ( .A(a[211]), .B(b[1]), .Z(n5022) );
  AND U5260 ( .A(a[209]), .B(b[3]), .Z(n5021) );
  XOR U5261 ( .A(n5022), .B(n5021), .Z(n5023) );
  XOR U5262 ( .A(n5024), .B(n5023), .Z(n5027) );
  NAND U5263 ( .A(b[0]), .B(a[212]), .Z(n5028) );
  XOR U5264 ( .A(n5027), .B(n5028), .Z(n5030) );
  OR U5265 ( .A(n4999), .B(n4998), .Z(n5003) );
  NANDN U5266 ( .A(n5001), .B(n5000), .Z(n5002) );
  NAND U5267 ( .A(n5003), .B(n5002), .Z(n5029) );
  XNOR U5268 ( .A(n5030), .B(n5029), .Z(n5015) );
  NANDN U5269 ( .A(n5005), .B(n5004), .Z(n5009) );
  OR U5270 ( .A(n5007), .B(n5006), .Z(n5008) );
  NAND U5271 ( .A(n5009), .B(n5008), .Z(n5016) );
  XNOR U5272 ( .A(n5015), .B(n5016), .Z(n5017) );
  XNOR U5273 ( .A(n5018), .B(n5017), .Z(n5033) );
  XNOR U5274 ( .A(n5033), .B(sreg[464]), .Z(n5035) );
  NAND U5275 ( .A(n5010), .B(sreg[463]), .Z(n5014) );
  OR U5276 ( .A(n5012), .B(n5011), .Z(n5013) );
  AND U5277 ( .A(n5014), .B(n5013), .Z(n5034) );
  XOR U5278 ( .A(n5035), .B(n5034), .Z(c[464]) );
  NANDN U5279 ( .A(n5016), .B(n5015), .Z(n5020) );
  NAND U5280 ( .A(n5018), .B(n5017), .Z(n5019) );
  NAND U5281 ( .A(n5020), .B(n5019), .Z(n5042) );
  AND U5282 ( .A(b[2]), .B(a[211]), .Z(n5048) );
  AND U5283 ( .A(a[212]), .B(b[1]), .Z(n5046) );
  AND U5284 ( .A(a[210]), .B(b[3]), .Z(n5045) );
  XOR U5285 ( .A(n5046), .B(n5045), .Z(n5047) );
  XOR U5286 ( .A(n5048), .B(n5047), .Z(n5051) );
  NAND U5287 ( .A(b[0]), .B(a[213]), .Z(n5052) );
  XOR U5288 ( .A(n5051), .B(n5052), .Z(n5054) );
  OR U5289 ( .A(n5022), .B(n5021), .Z(n5026) );
  NANDN U5290 ( .A(n5024), .B(n5023), .Z(n5025) );
  NAND U5291 ( .A(n5026), .B(n5025), .Z(n5053) );
  XNOR U5292 ( .A(n5054), .B(n5053), .Z(n5039) );
  NANDN U5293 ( .A(n5028), .B(n5027), .Z(n5032) );
  OR U5294 ( .A(n5030), .B(n5029), .Z(n5031) );
  NAND U5295 ( .A(n5032), .B(n5031), .Z(n5040) );
  XNOR U5296 ( .A(n5039), .B(n5040), .Z(n5041) );
  XNOR U5297 ( .A(n5042), .B(n5041), .Z(n5058) );
  NAND U5298 ( .A(n5033), .B(sreg[464]), .Z(n5037) );
  OR U5299 ( .A(n5035), .B(n5034), .Z(n5036) );
  AND U5300 ( .A(n5037), .B(n5036), .Z(n5057) );
  XNOR U5301 ( .A(n5057), .B(sreg[465]), .Z(n5038) );
  XOR U5302 ( .A(n5058), .B(n5038), .Z(c[465]) );
  NANDN U5303 ( .A(n5040), .B(n5039), .Z(n5044) );
  NAND U5304 ( .A(n5042), .B(n5041), .Z(n5043) );
  NAND U5305 ( .A(n5044), .B(n5043), .Z(n5065) );
  AND U5306 ( .A(b[2]), .B(a[212]), .Z(n5071) );
  AND U5307 ( .A(a[213]), .B(b[1]), .Z(n5069) );
  AND U5308 ( .A(a[211]), .B(b[3]), .Z(n5068) );
  XOR U5309 ( .A(n5069), .B(n5068), .Z(n5070) );
  XOR U5310 ( .A(n5071), .B(n5070), .Z(n5074) );
  NAND U5311 ( .A(b[0]), .B(a[214]), .Z(n5075) );
  XOR U5312 ( .A(n5074), .B(n5075), .Z(n5077) );
  OR U5313 ( .A(n5046), .B(n5045), .Z(n5050) );
  NANDN U5314 ( .A(n5048), .B(n5047), .Z(n5049) );
  NAND U5315 ( .A(n5050), .B(n5049), .Z(n5076) );
  XNOR U5316 ( .A(n5077), .B(n5076), .Z(n5062) );
  NANDN U5317 ( .A(n5052), .B(n5051), .Z(n5056) );
  OR U5318 ( .A(n5054), .B(n5053), .Z(n5055) );
  NAND U5319 ( .A(n5056), .B(n5055), .Z(n5063) );
  XNOR U5320 ( .A(n5062), .B(n5063), .Z(n5064) );
  XOR U5321 ( .A(n5065), .B(n5064), .Z(n5061) );
  XOR U5322 ( .A(sreg[466]), .B(n5060), .Z(n5059) );
  XOR U5323 ( .A(n5061), .B(n5059), .Z(c[466]) );
  NANDN U5324 ( .A(n5063), .B(n5062), .Z(n5067) );
  NAND U5325 ( .A(n5065), .B(n5064), .Z(n5066) );
  NAND U5326 ( .A(n5067), .B(n5066), .Z(n5083) );
  AND U5327 ( .A(b[2]), .B(a[213]), .Z(n5089) );
  AND U5328 ( .A(a[214]), .B(b[1]), .Z(n5087) );
  AND U5329 ( .A(a[212]), .B(b[3]), .Z(n5086) );
  XOR U5330 ( .A(n5087), .B(n5086), .Z(n5088) );
  XOR U5331 ( .A(n5089), .B(n5088), .Z(n5092) );
  NAND U5332 ( .A(b[0]), .B(a[215]), .Z(n5093) );
  XOR U5333 ( .A(n5092), .B(n5093), .Z(n5095) );
  OR U5334 ( .A(n5069), .B(n5068), .Z(n5073) );
  NANDN U5335 ( .A(n5071), .B(n5070), .Z(n5072) );
  NAND U5336 ( .A(n5073), .B(n5072), .Z(n5094) );
  XNOR U5337 ( .A(n5095), .B(n5094), .Z(n5080) );
  NANDN U5338 ( .A(n5075), .B(n5074), .Z(n5079) );
  OR U5339 ( .A(n5077), .B(n5076), .Z(n5078) );
  NAND U5340 ( .A(n5079), .B(n5078), .Z(n5081) );
  XNOR U5341 ( .A(n5080), .B(n5081), .Z(n5082) );
  XNOR U5342 ( .A(n5083), .B(n5082), .Z(n5098) );
  XNOR U5343 ( .A(n5098), .B(sreg[467]), .Z(n5099) );
  XOR U5344 ( .A(n5100), .B(n5099), .Z(c[467]) );
  NANDN U5345 ( .A(n5081), .B(n5080), .Z(n5085) );
  NAND U5346 ( .A(n5083), .B(n5082), .Z(n5084) );
  NAND U5347 ( .A(n5085), .B(n5084), .Z(n5107) );
  AND U5348 ( .A(b[2]), .B(a[214]), .Z(n5113) );
  AND U5349 ( .A(a[215]), .B(b[1]), .Z(n5111) );
  AND U5350 ( .A(a[213]), .B(b[3]), .Z(n5110) );
  XOR U5351 ( .A(n5111), .B(n5110), .Z(n5112) );
  XOR U5352 ( .A(n5113), .B(n5112), .Z(n5116) );
  NAND U5353 ( .A(b[0]), .B(a[216]), .Z(n5117) );
  XOR U5354 ( .A(n5116), .B(n5117), .Z(n5119) );
  OR U5355 ( .A(n5087), .B(n5086), .Z(n5091) );
  NANDN U5356 ( .A(n5089), .B(n5088), .Z(n5090) );
  NAND U5357 ( .A(n5091), .B(n5090), .Z(n5118) );
  XNOR U5358 ( .A(n5119), .B(n5118), .Z(n5104) );
  NANDN U5359 ( .A(n5093), .B(n5092), .Z(n5097) );
  OR U5360 ( .A(n5095), .B(n5094), .Z(n5096) );
  NAND U5361 ( .A(n5097), .B(n5096), .Z(n5105) );
  XNOR U5362 ( .A(n5104), .B(n5105), .Z(n5106) );
  XNOR U5363 ( .A(n5107), .B(n5106), .Z(n5123) );
  NAND U5364 ( .A(n5098), .B(sreg[467]), .Z(n5102) );
  OR U5365 ( .A(n5100), .B(n5099), .Z(n5101) );
  AND U5366 ( .A(n5102), .B(n5101), .Z(n5122) );
  XNOR U5367 ( .A(n5122), .B(sreg[468]), .Z(n5103) );
  XOR U5368 ( .A(n5123), .B(n5103), .Z(c[468]) );
  NANDN U5369 ( .A(n5105), .B(n5104), .Z(n5109) );
  NAND U5370 ( .A(n5107), .B(n5106), .Z(n5108) );
  NAND U5371 ( .A(n5109), .B(n5108), .Z(n5128) );
  AND U5372 ( .A(b[2]), .B(a[215]), .Z(n5134) );
  AND U5373 ( .A(a[216]), .B(b[1]), .Z(n5132) );
  AND U5374 ( .A(a[214]), .B(b[3]), .Z(n5131) );
  XOR U5375 ( .A(n5132), .B(n5131), .Z(n5133) );
  XOR U5376 ( .A(n5134), .B(n5133), .Z(n5137) );
  NAND U5377 ( .A(b[0]), .B(a[217]), .Z(n5138) );
  XOR U5378 ( .A(n5137), .B(n5138), .Z(n5140) );
  OR U5379 ( .A(n5111), .B(n5110), .Z(n5115) );
  NANDN U5380 ( .A(n5113), .B(n5112), .Z(n5114) );
  NAND U5381 ( .A(n5115), .B(n5114), .Z(n5139) );
  XNOR U5382 ( .A(n5140), .B(n5139), .Z(n5125) );
  NANDN U5383 ( .A(n5117), .B(n5116), .Z(n5121) );
  OR U5384 ( .A(n5119), .B(n5118), .Z(n5120) );
  NAND U5385 ( .A(n5121), .B(n5120), .Z(n5126) );
  XNOR U5386 ( .A(n5125), .B(n5126), .Z(n5127) );
  XOR U5387 ( .A(n5128), .B(n5127), .Z(n5144) );
  XOR U5388 ( .A(sreg[469]), .B(n5143), .Z(n5124) );
  XOR U5389 ( .A(n5144), .B(n5124), .Z(c[469]) );
  NANDN U5390 ( .A(n5126), .B(n5125), .Z(n5130) );
  NAND U5391 ( .A(n5128), .B(n5127), .Z(n5129) );
  NAND U5392 ( .A(n5130), .B(n5129), .Z(n5151) );
  AND U5393 ( .A(b[2]), .B(a[216]), .Z(n5157) );
  AND U5394 ( .A(a[217]), .B(b[1]), .Z(n5155) );
  AND U5395 ( .A(a[215]), .B(b[3]), .Z(n5154) );
  XOR U5396 ( .A(n5155), .B(n5154), .Z(n5156) );
  XOR U5397 ( .A(n5157), .B(n5156), .Z(n5160) );
  NAND U5398 ( .A(b[0]), .B(a[218]), .Z(n5161) );
  XOR U5399 ( .A(n5160), .B(n5161), .Z(n5163) );
  OR U5400 ( .A(n5132), .B(n5131), .Z(n5136) );
  NANDN U5401 ( .A(n5134), .B(n5133), .Z(n5135) );
  NAND U5402 ( .A(n5136), .B(n5135), .Z(n5162) );
  XNOR U5403 ( .A(n5163), .B(n5162), .Z(n5148) );
  NANDN U5404 ( .A(n5138), .B(n5137), .Z(n5142) );
  OR U5405 ( .A(n5140), .B(n5139), .Z(n5141) );
  NAND U5406 ( .A(n5142), .B(n5141), .Z(n5149) );
  XNOR U5407 ( .A(n5148), .B(n5149), .Z(n5150) );
  XNOR U5408 ( .A(n5151), .B(n5150), .Z(n5147) );
  XOR U5409 ( .A(n5146), .B(sreg[470]), .Z(n5145) );
  XOR U5410 ( .A(n5147), .B(n5145), .Z(c[470]) );
  NANDN U5411 ( .A(n5149), .B(n5148), .Z(n5153) );
  NAND U5412 ( .A(n5151), .B(n5150), .Z(n5152) );
  NAND U5413 ( .A(n5153), .B(n5152), .Z(n5169) );
  AND U5414 ( .A(b[2]), .B(a[217]), .Z(n5175) );
  AND U5415 ( .A(a[218]), .B(b[1]), .Z(n5173) );
  AND U5416 ( .A(a[216]), .B(b[3]), .Z(n5172) );
  XOR U5417 ( .A(n5173), .B(n5172), .Z(n5174) );
  XOR U5418 ( .A(n5175), .B(n5174), .Z(n5178) );
  NAND U5419 ( .A(b[0]), .B(a[219]), .Z(n5179) );
  XOR U5420 ( .A(n5178), .B(n5179), .Z(n5181) );
  OR U5421 ( .A(n5155), .B(n5154), .Z(n5159) );
  NANDN U5422 ( .A(n5157), .B(n5156), .Z(n5158) );
  NAND U5423 ( .A(n5159), .B(n5158), .Z(n5180) );
  XNOR U5424 ( .A(n5181), .B(n5180), .Z(n5166) );
  NANDN U5425 ( .A(n5161), .B(n5160), .Z(n5165) );
  OR U5426 ( .A(n5163), .B(n5162), .Z(n5164) );
  NAND U5427 ( .A(n5165), .B(n5164), .Z(n5167) );
  XNOR U5428 ( .A(n5166), .B(n5167), .Z(n5168) );
  XNOR U5429 ( .A(n5169), .B(n5168), .Z(n5184) );
  XNOR U5430 ( .A(n5184), .B(sreg[471]), .Z(n5186) );
  XNOR U5431 ( .A(n5185), .B(n5186), .Z(c[471]) );
  NANDN U5432 ( .A(n5167), .B(n5166), .Z(n5171) );
  NAND U5433 ( .A(n5169), .B(n5168), .Z(n5170) );
  NAND U5434 ( .A(n5171), .B(n5170), .Z(n5193) );
  AND U5435 ( .A(b[2]), .B(a[218]), .Z(n5199) );
  AND U5436 ( .A(a[219]), .B(b[1]), .Z(n5197) );
  AND U5437 ( .A(a[217]), .B(b[3]), .Z(n5196) );
  XOR U5438 ( .A(n5197), .B(n5196), .Z(n5198) );
  XOR U5439 ( .A(n5199), .B(n5198), .Z(n5202) );
  NAND U5440 ( .A(b[0]), .B(a[220]), .Z(n5203) );
  XOR U5441 ( .A(n5202), .B(n5203), .Z(n5205) );
  OR U5442 ( .A(n5173), .B(n5172), .Z(n5177) );
  NANDN U5443 ( .A(n5175), .B(n5174), .Z(n5176) );
  NAND U5444 ( .A(n5177), .B(n5176), .Z(n5204) );
  XNOR U5445 ( .A(n5205), .B(n5204), .Z(n5190) );
  NANDN U5446 ( .A(n5179), .B(n5178), .Z(n5183) );
  OR U5447 ( .A(n5181), .B(n5180), .Z(n5182) );
  NAND U5448 ( .A(n5183), .B(n5182), .Z(n5191) );
  XNOR U5449 ( .A(n5190), .B(n5191), .Z(n5192) );
  XNOR U5450 ( .A(n5193), .B(n5192), .Z(n5209) );
  NAND U5451 ( .A(n5184), .B(sreg[471]), .Z(n5188) );
  NANDN U5452 ( .A(n5186), .B(n5185), .Z(n5187) );
  AND U5453 ( .A(n5188), .B(n5187), .Z(n5208) );
  XNOR U5454 ( .A(n5208), .B(sreg[472]), .Z(n5189) );
  XOR U5455 ( .A(n5209), .B(n5189), .Z(c[472]) );
  NANDN U5456 ( .A(n5191), .B(n5190), .Z(n5195) );
  NAND U5457 ( .A(n5193), .B(n5192), .Z(n5194) );
  NAND U5458 ( .A(n5195), .B(n5194), .Z(n5214) );
  AND U5459 ( .A(b[2]), .B(a[219]), .Z(n5220) );
  AND U5460 ( .A(a[220]), .B(b[1]), .Z(n5218) );
  AND U5461 ( .A(a[218]), .B(b[3]), .Z(n5217) );
  XOR U5462 ( .A(n5218), .B(n5217), .Z(n5219) );
  XOR U5463 ( .A(n5220), .B(n5219), .Z(n5223) );
  NAND U5464 ( .A(b[0]), .B(a[221]), .Z(n5224) );
  XOR U5465 ( .A(n5223), .B(n5224), .Z(n5226) );
  OR U5466 ( .A(n5197), .B(n5196), .Z(n5201) );
  NANDN U5467 ( .A(n5199), .B(n5198), .Z(n5200) );
  NAND U5468 ( .A(n5201), .B(n5200), .Z(n5225) );
  XNOR U5469 ( .A(n5226), .B(n5225), .Z(n5211) );
  NANDN U5470 ( .A(n5203), .B(n5202), .Z(n5207) );
  OR U5471 ( .A(n5205), .B(n5204), .Z(n5206) );
  NAND U5472 ( .A(n5207), .B(n5206), .Z(n5212) );
  XNOR U5473 ( .A(n5211), .B(n5212), .Z(n5213) );
  XNOR U5474 ( .A(n5214), .B(n5213), .Z(n5229) );
  XNOR U5475 ( .A(sreg[473]), .B(n5230), .Z(n5210) );
  XNOR U5476 ( .A(n5229), .B(n5210), .Z(c[473]) );
  NANDN U5477 ( .A(n5212), .B(n5211), .Z(n5216) );
  NAND U5478 ( .A(n5214), .B(n5213), .Z(n5215) );
  NAND U5479 ( .A(n5216), .B(n5215), .Z(n5237) );
  AND U5480 ( .A(b[2]), .B(a[220]), .Z(n5243) );
  AND U5481 ( .A(a[221]), .B(b[1]), .Z(n5241) );
  AND U5482 ( .A(a[219]), .B(b[3]), .Z(n5240) );
  XOR U5483 ( .A(n5241), .B(n5240), .Z(n5242) );
  XOR U5484 ( .A(n5243), .B(n5242), .Z(n5246) );
  NAND U5485 ( .A(b[0]), .B(a[222]), .Z(n5247) );
  XOR U5486 ( .A(n5246), .B(n5247), .Z(n5249) );
  OR U5487 ( .A(n5218), .B(n5217), .Z(n5222) );
  NANDN U5488 ( .A(n5220), .B(n5219), .Z(n5221) );
  NAND U5489 ( .A(n5222), .B(n5221), .Z(n5248) );
  XNOR U5490 ( .A(n5249), .B(n5248), .Z(n5234) );
  NANDN U5491 ( .A(n5224), .B(n5223), .Z(n5228) );
  OR U5492 ( .A(n5226), .B(n5225), .Z(n5227) );
  NAND U5493 ( .A(n5228), .B(n5227), .Z(n5235) );
  XNOR U5494 ( .A(n5234), .B(n5235), .Z(n5236) );
  XNOR U5495 ( .A(n5237), .B(n5236), .Z(n5233) );
  XOR U5496 ( .A(n5232), .B(sreg[474]), .Z(n5231) );
  XOR U5497 ( .A(n5233), .B(n5231), .Z(c[474]) );
  NANDN U5498 ( .A(n5235), .B(n5234), .Z(n5239) );
  NAND U5499 ( .A(n5237), .B(n5236), .Z(n5238) );
  NAND U5500 ( .A(n5239), .B(n5238), .Z(n5255) );
  AND U5501 ( .A(b[2]), .B(a[221]), .Z(n5261) );
  AND U5502 ( .A(a[222]), .B(b[1]), .Z(n5259) );
  AND U5503 ( .A(a[220]), .B(b[3]), .Z(n5258) );
  XOR U5504 ( .A(n5259), .B(n5258), .Z(n5260) );
  XOR U5505 ( .A(n5261), .B(n5260), .Z(n5264) );
  NAND U5506 ( .A(b[0]), .B(a[223]), .Z(n5265) );
  XOR U5507 ( .A(n5264), .B(n5265), .Z(n5267) );
  OR U5508 ( .A(n5241), .B(n5240), .Z(n5245) );
  NANDN U5509 ( .A(n5243), .B(n5242), .Z(n5244) );
  NAND U5510 ( .A(n5245), .B(n5244), .Z(n5266) );
  XNOR U5511 ( .A(n5267), .B(n5266), .Z(n5252) );
  NANDN U5512 ( .A(n5247), .B(n5246), .Z(n5251) );
  OR U5513 ( .A(n5249), .B(n5248), .Z(n5250) );
  NAND U5514 ( .A(n5251), .B(n5250), .Z(n5253) );
  XNOR U5515 ( .A(n5252), .B(n5253), .Z(n5254) );
  XNOR U5516 ( .A(n5255), .B(n5254), .Z(n5270) );
  XNOR U5517 ( .A(n5270), .B(sreg[475]), .Z(n5272) );
  XNOR U5518 ( .A(n5271), .B(n5272), .Z(c[475]) );
  NANDN U5519 ( .A(n5253), .B(n5252), .Z(n5257) );
  NAND U5520 ( .A(n5255), .B(n5254), .Z(n5256) );
  NAND U5521 ( .A(n5257), .B(n5256), .Z(n5283) );
  AND U5522 ( .A(b[2]), .B(a[222]), .Z(n5289) );
  AND U5523 ( .A(a[223]), .B(b[1]), .Z(n5287) );
  AND U5524 ( .A(a[221]), .B(b[3]), .Z(n5286) );
  XOR U5525 ( .A(n5287), .B(n5286), .Z(n5288) );
  XOR U5526 ( .A(n5289), .B(n5288), .Z(n5292) );
  NAND U5527 ( .A(b[0]), .B(a[224]), .Z(n5293) );
  XOR U5528 ( .A(n5292), .B(n5293), .Z(n5295) );
  OR U5529 ( .A(n5259), .B(n5258), .Z(n5263) );
  NANDN U5530 ( .A(n5261), .B(n5260), .Z(n5262) );
  NAND U5531 ( .A(n5263), .B(n5262), .Z(n5294) );
  XNOR U5532 ( .A(n5295), .B(n5294), .Z(n5280) );
  NANDN U5533 ( .A(n5265), .B(n5264), .Z(n5269) );
  OR U5534 ( .A(n5267), .B(n5266), .Z(n5268) );
  NAND U5535 ( .A(n5269), .B(n5268), .Z(n5281) );
  XNOR U5536 ( .A(n5280), .B(n5281), .Z(n5282) );
  XNOR U5537 ( .A(n5283), .B(n5282), .Z(n5275) );
  XOR U5538 ( .A(sreg[476]), .B(n5275), .Z(n5276) );
  NAND U5539 ( .A(n5270), .B(sreg[475]), .Z(n5274) );
  NANDN U5540 ( .A(n5272), .B(n5271), .Z(n5273) );
  NAND U5541 ( .A(n5274), .B(n5273), .Z(n5277) );
  XOR U5542 ( .A(n5276), .B(n5277), .Z(c[476]) );
  OR U5543 ( .A(n5275), .B(sreg[476]), .Z(n5279) );
  NANDN U5544 ( .A(n5277), .B(n5276), .Z(n5278) );
  NAND U5545 ( .A(n5279), .B(n5278), .Z(n5318) );
  NANDN U5546 ( .A(n5281), .B(n5280), .Z(n5285) );
  NAND U5547 ( .A(n5283), .B(n5282), .Z(n5284) );
  NAND U5548 ( .A(n5285), .B(n5284), .Z(n5301) );
  AND U5549 ( .A(b[2]), .B(a[223]), .Z(n5307) );
  AND U5550 ( .A(a[224]), .B(b[1]), .Z(n5305) );
  AND U5551 ( .A(a[222]), .B(b[3]), .Z(n5304) );
  XOR U5552 ( .A(n5305), .B(n5304), .Z(n5306) );
  XOR U5553 ( .A(n5307), .B(n5306), .Z(n5310) );
  NAND U5554 ( .A(b[0]), .B(a[225]), .Z(n5311) );
  XOR U5555 ( .A(n5310), .B(n5311), .Z(n5313) );
  OR U5556 ( .A(n5287), .B(n5286), .Z(n5291) );
  NANDN U5557 ( .A(n5289), .B(n5288), .Z(n5290) );
  NAND U5558 ( .A(n5291), .B(n5290), .Z(n5312) );
  XNOR U5559 ( .A(n5313), .B(n5312), .Z(n5298) );
  NANDN U5560 ( .A(n5293), .B(n5292), .Z(n5297) );
  OR U5561 ( .A(n5295), .B(n5294), .Z(n5296) );
  NAND U5562 ( .A(n5297), .B(n5296), .Z(n5299) );
  XNOR U5563 ( .A(n5298), .B(n5299), .Z(n5300) );
  XNOR U5564 ( .A(n5301), .B(n5300), .Z(n5316) );
  XNOR U5565 ( .A(n5316), .B(sreg[477]), .Z(n5317) );
  XOR U5566 ( .A(n5318), .B(n5317), .Z(c[477]) );
  NANDN U5567 ( .A(n5299), .B(n5298), .Z(n5303) );
  NAND U5568 ( .A(n5301), .B(n5300), .Z(n5302) );
  NAND U5569 ( .A(n5303), .B(n5302), .Z(n5324) );
  AND U5570 ( .A(b[2]), .B(a[224]), .Z(n5330) );
  AND U5571 ( .A(a[225]), .B(b[1]), .Z(n5328) );
  AND U5572 ( .A(a[223]), .B(b[3]), .Z(n5327) );
  XOR U5573 ( .A(n5328), .B(n5327), .Z(n5329) );
  XOR U5574 ( .A(n5330), .B(n5329), .Z(n5333) );
  NAND U5575 ( .A(b[0]), .B(a[226]), .Z(n5334) );
  XOR U5576 ( .A(n5333), .B(n5334), .Z(n5336) );
  OR U5577 ( .A(n5305), .B(n5304), .Z(n5309) );
  NANDN U5578 ( .A(n5307), .B(n5306), .Z(n5308) );
  NAND U5579 ( .A(n5309), .B(n5308), .Z(n5335) );
  XNOR U5580 ( .A(n5336), .B(n5335), .Z(n5321) );
  NANDN U5581 ( .A(n5311), .B(n5310), .Z(n5315) );
  OR U5582 ( .A(n5313), .B(n5312), .Z(n5314) );
  NAND U5583 ( .A(n5315), .B(n5314), .Z(n5322) );
  XNOR U5584 ( .A(n5321), .B(n5322), .Z(n5323) );
  XNOR U5585 ( .A(n5324), .B(n5323), .Z(n5339) );
  XNOR U5586 ( .A(n5339), .B(sreg[478]), .Z(n5341) );
  NAND U5587 ( .A(n5316), .B(sreg[477]), .Z(n5320) );
  OR U5588 ( .A(n5318), .B(n5317), .Z(n5319) );
  AND U5589 ( .A(n5320), .B(n5319), .Z(n5340) );
  XOR U5590 ( .A(n5341), .B(n5340), .Z(c[478]) );
  NANDN U5591 ( .A(n5322), .B(n5321), .Z(n5326) );
  NAND U5592 ( .A(n5324), .B(n5323), .Z(n5325) );
  NAND U5593 ( .A(n5326), .B(n5325), .Z(n5348) );
  AND U5594 ( .A(b[2]), .B(a[225]), .Z(n5354) );
  AND U5595 ( .A(a[226]), .B(b[1]), .Z(n5352) );
  AND U5596 ( .A(a[224]), .B(b[3]), .Z(n5351) );
  XOR U5597 ( .A(n5352), .B(n5351), .Z(n5353) );
  XOR U5598 ( .A(n5354), .B(n5353), .Z(n5357) );
  NAND U5599 ( .A(b[0]), .B(a[227]), .Z(n5358) );
  XOR U5600 ( .A(n5357), .B(n5358), .Z(n5360) );
  OR U5601 ( .A(n5328), .B(n5327), .Z(n5332) );
  NANDN U5602 ( .A(n5330), .B(n5329), .Z(n5331) );
  NAND U5603 ( .A(n5332), .B(n5331), .Z(n5359) );
  XNOR U5604 ( .A(n5360), .B(n5359), .Z(n5345) );
  NANDN U5605 ( .A(n5334), .B(n5333), .Z(n5338) );
  OR U5606 ( .A(n5336), .B(n5335), .Z(n5337) );
  NAND U5607 ( .A(n5338), .B(n5337), .Z(n5346) );
  XNOR U5608 ( .A(n5345), .B(n5346), .Z(n5347) );
  XNOR U5609 ( .A(n5348), .B(n5347), .Z(n5364) );
  NAND U5610 ( .A(n5339), .B(sreg[478]), .Z(n5343) );
  OR U5611 ( .A(n5341), .B(n5340), .Z(n5342) );
  AND U5612 ( .A(n5343), .B(n5342), .Z(n5363) );
  XNOR U5613 ( .A(n5363), .B(sreg[479]), .Z(n5344) );
  XOR U5614 ( .A(n5364), .B(n5344), .Z(c[479]) );
  NANDN U5615 ( .A(n5346), .B(n5345), .Z(n5350) );
  NAND U5616 ( .A(n5348), .B(n5347), .Z(n5349) );
  NAND U5617 ( .A(n5350), .B(n5349), .Z(n5371) );
  AND U5618 ( .A(b[2]), .B(a[226]), .Z(n5377) );
  AND U5619 ( .A(a[227]), .B(b[1]), .Z(n5375) );
  AND U5620 ( .A(a[225]), .B(b[3]), .Z(n5374) );
  XOR U5621 ( .A(n5375), .B(n5374), .Z(n5376) );
  XOR U5622 ( .A(n5377), .B(n5376), .Z(n5380) );
  NAND U5623 ( .A(b[0]), .B(a[228]), .Z(n5381) );
  XOR U5624 ( .A(n5380), .B(n5381), .Z(n5383) );
  OR U5625 ( .A(n5352), .B(n5351), .Z(n5356) );
  NANDN U5626 ( .A(n5354), .B(n5353), .Z(n5355) );
  NAND U5627 ( .A(n5356), .B(n5355), .Z(n5382) );
  XNOR U5628 ( .A(n5383), .B(n5382), .Z(n5368) );
  NANDN U5629 ( .A(n5358), .B(n5357), .Z(n5362) );
  OR U5630 ( .A(n5360), .B(n5359), .Z(n5361) );
  NAND U5631 ( .A(n5362), .B(n5361), .Z(n5369) );
  XNOR U5632 ( .A(n5368), .B(n5369), .Z(n5370) );
  XOR U5633 ( .A(n5371), .B(n5370), .Z(n5367) );
  XOR U5634 ( .A(sreg[480]), .B(n5366), .Z(n5365) );
  XOR U5635 ( .A(n5367), .B(n5365), .Z(c[480]) );
  NANDN U5636 ( .A(n5369), .B(n5368), .Z(n5373) );
  NAND U5637 ( .A(n5371), .B(n5370), .Z(n5372) );
  NAND U5638 ( .A(n5373), .B(n5372), .Z(n5389) );
  AND U5639 ( .A(b[2]), .B(a[227]), .Z(n5395) );
  AND U5640 ( .A(a[228]), .B(b[1]), .Z(n5393) );
  AND U5641 ( .A(a[226]), .B(b[3]), .Z(n5392) );
  XOR U5642 ( .A(n5393), .B(n5392), .Z(n5394) );
  XOR U5643 ( .A(n5395), .B(n5394), .Z(n5398) );
  NAND U5644 ( .A(b[0]), .B(a[229]), .Z(n5399) );
  XOR U5645 ( .A(n5398), .B(n5399), .Z(n5401) );
  OR U5646 ( .A(n5375), .B(n5374), .Z(n5379) );
  NANDN U5647 ( .A(n5377), .B(n5376), .Z(n5378) );
  NAND U5648 ( .A(n5379), .B(n5378), .Z(n5400) );
  XNOR U5649 ( .A(n5401), .B(n5400), .Z(n5386) );
  NANDN U5650 ( .A(n5381), .B(n5380), .Z(n5385) );
  OR U5651 ( .A(n5383), .B(n5382), .Z(n5384) );
  NAND U5652 ( .A(n5385), .B(n5384), .Z(n5387) );
  XNOR U5653 ( .A(n5386), .B(n5387), .Z(n5388) );
  XNOR U5654 ( .A(n5389), .B(n5388), .Z(n5404) );
  XNOR U5655 ( .A(n5404), .B(sreg[481]), .Z(n5405) );
  XOR U5656 ( .A(n5406), .B(n5405), .Z(c[481]) );
  NANDN U5657 ( .A(n5387), .B(n5386), .Z(n5391) );
  NAND U5658 ( .A(n5389), .B(n5388), .Z(n5390) );
  NAND U5659 ( .A(n5391), .B(n5390), .Z(n5415) );
  AND U5660 ( .A(b[2]), .B(a[228]), .Z(n5421) );
  AND U5661 ( .A(a[229]), .B(b[1]), .Z(n5419) );
  AND U5662 ( .A(a[227]), .B(b[3]), .Z(n5418) );
  XOR U5663 ( .A(n5419), .B(n5418), .Z(n5420) );
  XOR U5664 ( .A(n5421), .B(n5420), .Z(n5424) );
  NAND U5665 ( .A(b[0]), .B(a[230]), .Z(n5425) );
  XOR U5666 ( .A(n5424), .B(n5425), .Z(n5427) );
  OR U5667 ( .A(n5393), .B(n5392), .Z(n5397) );
  NANDN U5668 ( .A(n5395), .B(n5394), .Z(n5396) );
  NAND U5669 ( .A(n5397), .B(n5396), .Z(n5426) );
  XNOR U5670 ( .A(n5427), .B(n5426), .Z(n5412) );
  NANDN U5671 ( .A(n5399), .B(n5398), .Z(n5403) );
  OR U5672 ( .A(n5401), .B(n5400), .Z(n5402) );
  NAND U5673 ( .A(n5403), .B(n5402), .Z(n5413) );
  XNOR U5674 ( .A(n5412), .B(n5413), .Z(n5414) );
  XNOR U5675 ( .A(n5415), .B(n5414), .Z(n5411) );
  NAND U5676 ( .A(n5404), .B(sreg[481]), .Z(n5408) );
  OR U5677 ( .A(n5406), .B(n5405), .Z(n5407) );
  AND U5678 ( .A(n5408), .B(n5407), .Z(n5410) );
  XNOR U5679 ( .A(n5410), .B(sreg[482]), .Z(n5409) );
  XOR U5680 ( .A(n5411), .B(n5409), .Z(c[482]) );
  NANDN U5681 ( .A(n5413), .B(n5412), .Z(n5417) );
  NAND U5682 ( .A(n5415), .B(n5414), .Z(n5416) );
  NAND U5683 ( .A(n5417), .B(n5416), .Z(n5433) );
  AND U5684 ( .A(b[2]), .B(a[229]), .Z(n5439) );
  AND U5685 ( .A(a[230]), .B(b[1]), .Z(n5437) );
  AND U5686 ( .A(a[228]), .B(b[3]), .Z(n5436) );
  XOR U5687 ( .A(n5437), .B(n5436), .Z(n5438) );
  XOR U5688 ( .A(n5439), .B(n5438), .Z(n5442) );
  NAND U5689 ( .A(b[0]), .B(a[231]), .Z(n5443) );
  XOR U5690 ( .A(n5442), .B(n5443), .Z(n5445) );
  OR U5691 ( .A(n5419), .B(n5418), .Z(n5423) );
  NANDN U5692 ( .A(n5421), .B(n5420), .Z(n5422) );
  NAND U5693 ( .A(n5423), .B(n5422), .Z(n5444) );
  XNOR U5694 ( .A(n5445), .B(n5444), .Z(n5430) );
  NANDN U5695 ( .A(n5425), .B(n5424), .Z(n5429) );
  OR U5696 ( .A(n5427), .B(n5426), .Z(n5428) );
  NAND U5697 ( .A(n5429), .B(n5428), .Z(n5431) );
  XNOR U5698 ( .A(n5430), .B(n5431), .Z(n5432) );
  XNOR U5699 ( .A(n5433), .B(n5432), .Z(n5448) );
  XNOR U5700 ( .A(n5448), .B(sreg[483]), .Z(n5450) );
  XNOR U5701 ( .A(n5449), .B(n5450), .Z(c[483]) );
  NANDN U5702 ( .A(n5431), .B(n5430), .Z(n5435) );
  NAND U5703 ( .A(n5433), .B(n5432), .Z(n5434) );
  NAND U5704 ( .A(n5435), .B(n5434), .Z(n5459) );
  AND U5705 ( .A(b[2]), .B(a[230]), .Z(n5465) );
  AND U5706 ( .A(a[231]), .B(b[1]), .Z(n5463) );
  AND U5707 ( .A(a[229]), .B(b[3]), .Z(n5462) );
  XOR U5708 ( .A(n5463), .B(n5462), .Z(n5464) );
  XOR U5709 ( .A(n5465), .B(n5464), .Z(n5468) );
  NAND U5710 ( .A(b[0]), .B(a[232]), .Z(n5469) );
  XOR U5711 ( .A(n5468), .B(n5469), .Z(n5471) );
  OR U5712 ( .A(n5437), .B(n5436), .Z(n5441) );
  NANDN U5713 ( .A(n5439), .B(n5438), .Z(n5440) );
  NAND U5714 ( .A(n5441), .B(n5440), .Z(n5470) );
  XNOR U5715 ( .A(n5471), .B(n5470), .Z(n5456) );
  NANDN U5716 ( .A(n5443), .B(n5442), .Z(n5447) );
  OR U5717 ( .A(n5445), .B(n5444), .Z(n5446) );
  NAND U5718 ( .A(n5447), .B(n5446), .Z(n5457) );
  XNOR U5719 ( .A(n5456), .B(n5457), .Z(n5458) );
  XOR U5720 ( .A(n5459), .B(n5458), .Z(n5455) );
  NAND U5721 ( .A(n5448), .B(sreg[483]), .Z(n5452) );
  NANDN U5722 ( .A(n5450), .B(n5449), .Z(n5451) );
  NAND U5723 ( .A(n5452), .B(n5451), .Z(n5454) );
  XNOR U5724 ( .A(sreg[484]), .B(n5454), .Z(n5453) );
  XOR U5725 ( .A(n5455), .B(n5453), .Z(c[484]) );
  NANDN U5726 ( .A(n5457), .B(n5456), .Z(n5461) );
  NAND U5727 ( .A(n5459), .B(n5458), .Z(n5460) );
  NAND U5728 ( .A(n5461), .B(n5460), .Z(n5477) );
  AND U5729 ( .A(b[2]), .B(a[231]), .Z(n5483) );
  AND U5730 ( .A(a[232]), .B(b[1]), .Z(n5481) );
  AND U5731 ( .A(a[230]), .B(b[3]), .Z(n5480) );
  XOR U5732 ( .A(n5481), .B(n5480), .Z(n5482) );
  XOR U5733 ( .A(n5483), .B(n5482), .Z(n5486) );
  NAND U5734 ( .A(b[0]), .B(a[233]), .Z(n5487) );
  XOR U5735 ( .A(n5486), .B(n5487), .Z(n5489) );
  OR U5736 ( .A(n5463), .B(n5462), .Z(n5467) );
  NANDN U5737 ( .A(n5465), .B(n5464), .Z(n5466) );
  NAND U5738 ( .A(n5467), .B(n5466), .Z(n5488) );
  XNOR U5739 ( .A(n5489), .B(n5488), .Z(n5474) );
  NANDN U5740 ( .A(n5469), .B(n5468), .Z(n5473) );
  OR U5741 ( .A(n5471), .B(n5470), .Z(n5472) );
  NAND U5742 ( .A(n5473), .B(n5472), .Z(n5475) );
  XNOR U5743 ( .A(n5474), .B(n5475), .Z(n5476) );
  XNOR U5744 ( .A(n5477), .B(n5476), .Z(n5492) );
  XNOR U5745 ( .A(n5492), .B(sreg[485]), .Z(n5493) );
  XOR U5746 ( .A(n5494), .B(n5493), .Z(c[485]) );
  NANDN U5747 ( .A(n5475), .B(n5474), .Z(n5479) );
  NAND U5748 ( .A(n5477), .B(n5476), .Z(n5478) );
  NAND U5749 ( .A(n5479), .B(n5478), .Z(n5500) );
  AND U5750 ( .A(b[2]), .B(a[232]), .Z(n5506) );
  AND U5751 ( .A(a[233]), .B(b[1]), .Z(n5504) );
  AND U5752 ( .A(a[231]), .B(b[3]), .Z(n5503) );
  XOR U5753 ( .A(n5504), .B(n5503), .Z(n5505) );
  XOR U5754 ( .A(n5506), .B(n5505), .Z(n5509) );
  NAND U5755 ( .A(b[0]), .B(a[234]), .Z(n5510) );
  XOR U5756 ( .A(n5509), .B(n5510), .Z(n5512) );
  OR U5757 ( .A(n5481), .B(n5480), .Z(n5485) );
  NANDN U5758 ( .A(n5483), .B(n5482), .Z(n5484) );
  NAND U5759 ( .A(n5485), .B(n5484), .Z(n5511) );
  XNOR U5760 ( .A(n5512), .B(n5511), .Z(n5497) );
  NANDN U5761 ( .A(n5487), .B(n5486), .Z(n5491) );
  OR U5762 ( .A(n5489), .B(n5488), .Z(n5490) );
  NAND U5763 ( .A(n5491), .B(n5490), .Z(n5498) );
  XNOR U5764 ( .A(n5497), .B(n5498), .Z(n5499) );
  XNOR U5765 ( .A(n5500), .B(n5499), .Z(n5515) );
  XOR U5766 ( .A(sreg[486]), .B(n5515), .Z(n5516) );
  NAND U5767 ( .A(n5492), .B(sreg[485]), .Z(n5496) );
  OR U5768 ( .A(n5494), .B(n5493), .Z(n5495) );
  NAND U5769 ( .A(n5496), .B(n5495), .Z(n5517) );
  XOR U5770 ( .A(n5516), .B(n5517), .Z(c[486]) );
  NANDN U5771 ( .A(n5498), .B(n5497), .Z(n5502) );
  NAND U5772 ( .A(n5500), .B(n5499), .Z(n5501) );
  NAND U5773 ( .A(n5502), .B(n5501), .Z(n5528) );
  AND U5774 ( .A(b[2]), .B(a[233]), .Z(n5534) );
  AND U5775 ( .A(a[234]), .B(b[1]), .Z(n5532) );
  AND U5776 ( .A(a[232]), .B(b[3]), .Z(n5531) );
  XOR U5777 ( .A(n5532), .B(n5531), .Z(n5533) );
  XOR U5778 ( .A(n5534), .B(n5533), .Z(n5537) );
  NAND U5779 ( .A(b[0]), .B(a[235]), .Z(n5538) );
  XOR U5780 ( .A(n5537), .B(n5538), .Z(n5540) );
  OR U5781 ( .A(n5504), .B(n5503), .Z(n5508) );
  NANDN U5782 ( .A(n5506), .B(n5505), .Z(n5507) );
  NAND U5783 ( .A(n5508), .B(n5507), .Z(n5539) );
  XNOR U5784 ( .A(n5540), .B(n5539), .Z(n5525) );
  NANDN U5785 ( .A(n5510), .B(n5509), .Z(n5514) );
  OR U5786 ( .A(n5512), .B(n5511), .Z(n5513) );
  NAND U5787 ( .A(n5514), .B(n5513), .Z(n5526) );
  XNOR U5788 ( .A(n5525), .B(n5526), .Z(n5527) );
  XNOR U5789 ( .A(n5528), .B(n5527), .Z(n5520) );
  XOR U5790 ( .A(sreg[487]), .B(n5520), .Z(n5521) );
  OR U5791 ( .A(n5515), .B(sreg[486]), .Z(n5519) );
  NANDN U5792 ( .A(n5517), .B(n5516), .Z(n5518) );
  AND U5793 ( .A(n5519), .B(n5518), .Z(n5522) );
  XOR U5794 ( .A(n5521), .B(n5522), .Z(c[487]) );
  OR U5795 ( .A(n5520), .B(sreg[487]), .Z(n5524) );
  NANDN U5796 ( .A(n5522), .B(n5521), .Z(n5523) );
  AND U5797 ( .A(n5524), .B(n5523), .Z(n5544) );
  NANDN U5798 ( .A(n5526), .B(n5525), .Z(n5530) );
  NAND U5799 ( .A(n5528), .B(n5527), .Z(n5529) );
  NAND U5800 ( .A(n5530), .B(n5529), .Z(n5549) );
  AND U5801 ( .A(b[2]), .B(a[234]), .Z(n5555) );
  AND U5802 ( .A(a[235]), .B(b[1]), .Z(n5553) );
  AND U5803 ( .A(a[233]), .B(b[3]), .Z(n5552) );
  XOR U5804 ( .A(n5553), .B(n5552), .Z(n5554) );
  XOR U5805 ( .A(n5555), .B(n5554), .Z(n5558) );
  NAND U5806 ( .A(b[0]), .B(a[236]), .Z(n5559) );
  XOR U5807 ( .A(n5558), .B(n5559), .Z(n5561) );
  OR U5808 ( .A(n5532), .B(n5531), .Z(n5536) );
  NANDN U5809 ( .A(n5534), .B(n5533), .Z(n5535) );
  NAND U5810 ( .A(n5536), .B(n5535), .Z(n5560) );
  XNOR U5811 ( .A(n5561), .B(n5560), .Z(n5546) );
  NANDN U5812 ( .A(n5538), .B(n5537), .Z(n5542) );
  OR U5813 ( .A(n5540), .B(n5539), .Z(n5541) );
  NAND U5814 ( .A(n5542), .B(n5541), .Z(n5547) );
  XNOR U5815 ( .A(n5546), .B(n5547), .Z(n5548) );
  XNOR U5816 ( .A(n5549), .B(n5548), .Z(n5545) );
  XOR U5817 ( .A(sreg[488]), .B(n5545), .Z(n5543) );
  XOR U5818 ( .A(n5544), .B(n5543), .Z(c[488]) );
  NANDN U5819 ( .A(n5547), .B(n5546), .Z(n5551) );
  NAND U5820 ( .A(n5549), .B(n5548), .Z(n5550) );
  NAND U5821 ( .A(n5551), .B(n5550), .Z(n5567) );
  AND U5822 ( .A(b[2]), .B(a[235]), .Z(n5573) );
  AND U5823 ( .A(a[236]), .B(b[1]), .Z(n5571) );
  AND U5824 ( .A(a[234]), .B(b[3]), .Z(n5570) );
  XOR U5825 ( .A(n5571), .B(n5570), .Z(n5572) );
  XOR U5826 ( .A(n5573), .B(n5572), .Z(n5576) );
  NAND U5827 ( .A(b[0]), .B(a[237]), .Z(n5577) );
  XOR U5828 ( .A(n5576), .B(n5577), .Z(n5579) );
  OR U5829 ( .A(n5553), .B(n5552), .Z(n5557) );
  NANDN U5830 ( .A(n5555), .B(n5554), .Z(n5556) );
  NAND U5831 ( .A(n5557), .B(n5556), .Z(n5578) );
  XNOR U5832 ( .A(n5579), .B(n5578), .Z(n5564) );
  NANDN U5833 ( .A(n5559), .B(n5558), .Z(n5563) );
  OR U5834 ( .A(n5561), .B(n5560), .Z(n5562) );
  NAND U5835 ( .A(n5563), .B(n5562), .Z(n5565) );
  XNOR U5836 ( .A(n5564), .B(n5565), .Z(n5566) );
  XNOR U5837 ( .A(n5567), .B(n5566), .Z(n5582) );
  XNOR U5838 ( .A(n5582), .B(sreg[489]), .Z(n5584) );
  XNOR U5839 ( .A(n5583), .B(n5584), .Z(c[489]) );
  NANDN U5840 ( .A(n5565), .B(n5564), .Z(n5569) );
  NAND U5841 ( .A(n5567), .B(n5566), .Z(n5568) );
  NAND U5842 ( .A(n5569), .B(n5568), .Z(n5595) );
  AND U5843 ( .A(b[2]), .B(a[236]), .Z(n5601) );
  AND U5844 ( .A(a[237]), .B(b[1]), .Z(n5599) );
  AND U5845 ( .A(a[235]), .B(b[3]), .Z(n5598) );
  XOR U5846 ( .A(n5599), .B(n5598), .Z(n5600) );
  XOR U5847 ( .A(n5601), .B(n5600), .Z(n5604) );
  NAND U5848 ( .A(b[0]), .B(a[238]), .Z(n5605) );
  XOR U5849 ( .A(n5604), .B(n5605), .Z(n5607) );
  OR U5850 ( .A(n5571), .B(n5570), .Z(n5575) );
  NANDN U5851 ( .A(n5573), .B(n5572), .Z(n5574) );
  NAND U5852 ( .A(n5575), .B(n5574), .Z(n5606) );
  XNOR U5853 ( .A(n5607), .B(n5606), .Z(n5592) );
  NANDN U5854 ( .A(n5577), .B(n5576), .Z(n5581) );
  OR U5855 ( .A(n5579), .B(n5578), .Z(n5580) );
  NAND U5856 ( .A(n5581), .B(n5580), .Z(n5593) );
  XNOR U5857 ( .A(n5592), .B(n5593), .Z(n5594) );
  XNOR U5858 ( .A(n5595), .B(n5594), .Z(n5587) );
  XOR U5859 ( .A(sreg[490]), .B(n5587), .Z(n5588) );
  NAND U5860 ( .A(n5582), .B(sreg[489]), .Z(n5586) );
  NANDN U5861 ( .A(n5584), .B(n5583), .Z(n5585) );
  NAND U5862 ( .A(n5586), .B(n5585), .Z(n5589) );
  XOR U5863 ( .A(n5588), .B(n5589), .Z(c[490]) );
  OR U5864 ( .A(n5587), .B(sreg[490]), .Z(n5591) );
  NANDN U5865 ( .A(n5589), .B(n5588), .Z(n5590) );
  AND U5866 ( .A(n5591), .B(n5590), .Z(n5611) );
  NANDN U5867 ( .A(n5593), .B(n5592), .Z(n5597) );
  NAND U5868 ( .A(n5595), .B(n5594), .Z(n5596) );
  NAND U5869 ( .A(n5597), .B(n5596), .Z(n5616) );
  AND U5870 ( .A(b[2]), .B(a[237]), .Z(n5622) );
  AND U5871 ( .A(a[238]), .B(b[1]), .Z(n5620) );
  AND U5872 ( .A(a[236]), .B(b[3]), .Z(n5619) );
  XOR U5873 ( .A(n5620), .B(n5619), .Z(n5621) );
  XOR U5874 ( .A(n5622), .B(n5621), .Z(n5625) );
  NAND U5875 ( .A(b[0]), .B(a[239]), .Z(n5626) );
  XOR U5876 ( .A(n5625), .B(n5626), .Z(n5628) );
  OR U5877 ( .A(n5599), .B(n5598), .Z(n5603) );
  NANDN U5878 ( .A(n5601), .B(n5600), .Z(n5602) );
  NAND U5879 ( .A(n5603), .B(n5602), .Z(n5627) );
  XNOR U5880 ( .A(n5628), .B(n5627), .Z(n5613) );
  NANDN U5881 ( .A(n5605), .B(n5604), .Z(n5609) );
  OR U5882 ( .A(n5607), .B(n5606), .Z(n5608) );
  NAND U5883 ( .A(n5609), .B(n5608), .Z(n5614) );
  XNOR U5884 ( .A(n5613), .B(n5614), .Z(n5615) );
  XNOR U5885 ( .A(n5616), .B(n5615), .Z(n5612) );
  XOR U5886 ( .A(sreg[491]), .B(n5612), .Z(n5610) );
  XOR U5887 ( .A(n5611), .B(n5610), .Z(c[491]) );
  NANDN U5888 ( .A(n5614), .B(n5613), .Z(n5618) );
  NAND U5889 ( .A(n5616), .B(n5615), .Z(n5617) );
  NAND U5890 ( .A(n5618), .B(n5617), .Z(n5634) );
  AND U5891 ( .A(b[2]), .B(a[238]), .Z(n5646) );
  AND U5892 ( .A(a[239]), .B(b[1]), .Z(n5644) );
  AND U5893 ( .A(a[237]), .B(b[3]), .Z(n5643) );
  XOR U5894 ( .A(n5644), .B(n5643), .Z(n5645) );
  XOR U5895 ( .A(n5646), .B(n5645), .Z(n5637) );
  NAND U5896 ( .A(b[0]), .B(a[240]), .Z(n5638) );
  XOR U5897 ( .A(n5637), .B(n5638), .Z(n5640) );
  OR U5898 ( .A(n5620), .B(n5619), .Z(n5624) );
  NANDN U5899 ( .A(n5622), .B(n5621), .Z(n5623) );
  NAND U5900 ( .A(n5624), .B(n5623), .Z(n5639) );
  XNOR U5901 ( .A(n5640), .B(n5639), .Z(n5631) );
  NANDN U5902 ( .A(n5626), .B(n5625), .Z(n5630) );
  OR U5903 ( .A(n5628), .B(n5627), .Z(n5629) );
  NAND U5904 ( .A(n5630), .B(n5629), .Z(n5632) );
  XNOR U5905 ( .A(n5631), .B(n5632), .Z(n5633) );
  XOR U5906 ( .A(n5634), .B(n5633), .Z(n5650) );
  XOR U5907 ( .A(sreg[492]), .B(n5650), .Z(n5652) );
  XNOR U5908 ( .A(n5651), .B(n5652), .Z(c[492]) );
  NANDN U5909 ( .A(n5632), .B(n5631), .Z(n5636) );
  NAND U5910 ( .A(n5634), .B(n5633), .Z(n5635) );
  AND U5911 ( .A(n5636), .B(n5635), .Z(n5662) );
  NANDN U5912 ( .A(n5638), .B(n5637), .Z(n5642) );
  OR U5913 ( .A(n5640), .B(n5639), .Z(n5641) );
  AND U5914 ( .A(n5642), .B(n5641), .Z(n5661) );
  AND U5915 ( .A(b[2]), .B(a[239]), .Z(n5666) );
  AND U5916 ( .A(a[240]), .B(b[1]), .Z(n5664) );
  AND U5917 ( .A(a[238]), .B(b[3]), .Z(n5663) );
  XOR U5918 ( .A(n5664), .B(n5663), .Z(n5665) );
  XOR U5919 ( .A(n5666), .B(n5665), .Z(n5669) );
  NAND U5920 ( .A(b[0]), .B(a[241]), .Z(n5670) );
  XOR U5921 ( .A(n5669), .B(n5670), .Z(n5672) );
  OR U5922 ( .A(n5644), .B(n5643), .Z(n5648) );
  NANDN U5923 ( .A(n5646), .B(n5645), .Z(n5647) );
  NAND U5924 ( .A(n5648), .B(n5647), .Z(n5671) );
  XOR U5925 ( .A(n5672), .B(n5671), .Z(n5660) );
  XNOR U5926 ( .A(n5661), .B(n5660), .Z(n5649) );
  XOR U5927 ( .A(n5662), .B(n5649), .Z(n5655) );
  XNOR U5928 ( .A(sreg[493]), .B(n5655), .Z(n5657) );
  NANDN U5929 ( .A(n5650), .B(sreg[492]), .Z(n5654) );
  NANDN U5930 ( .A(n5652), .B(n5651), .Z(n5653) );
  AND U5931 ( .A(n5654), .B(n5653), .Z(n5656) );
  XOR U5932 ( .A(n5657), .B(n5656), .Z(c[493]) );
  NAND U5933 ( .A(sreg[493]), .B(n5655), .Z(n5659) );
  OR U5934 ( .A(n5657), .B(n5656), .Z(n5658) );
  NAND U5935 ( .A(n5659), .B(n5658), .Z(n5695) );
  AND U5936 ( .A(b[2]), .B(a[240]), .Z(n5684) );
  AND U5937 ( .A(a[241]), .B(b[1]), .Z(n5682) );
  AND U5938 ( .A(a[239]), .B(b[3]), .Z(n5681) );
  XOR U5939 ( .A(n5682), .B(n5681), .Z(n5683) );
  XOR U5940 ( .A(n5684), .B(n5683), .Z(n5687) );
  NAND U5941 ( .A(b[0]), .B(a[242]), .Z(n5688) );
  XOR U5942 ( .A(n5687), .B(n5688), .Z(n5690) );
  OR U5943 ( .A(n5664), .B(n5663), .Z(n5668) );
  NANDN U5944 ( .A(n5666), .B(n5665), .Z(n5667) );
  NAND U5945 ( .A(n5668), .B(n5667), .Z(n5689) );
  XNOR U5946 ( .A(n5690), .B(n5689), .Z(n5675) );
  NANDN U5947 ( .A(n5670), .B(n5669), .Z(n5674) );
  OR U5948 ( .A(n5672), .B(n5671), .Z(n5673) );
  NAND U5949 ( .A(n5674), .B(n5673), .Z(n5676) );
  XNOR U5950 ( .A(n5675), .B(n5676), .Z(n5677) );
  XNOR U5951 ( .A(n5678), .B(n5677), .Z(n5693) );
  XOR U5952 ( .A(sreg[494]), .B(n5693), .Z(n5694) );
  XNOR U5953 ( .A(n5695), .B(n5694), .Z(c[494]) );
  NANDN U5954 ( .A(n5676), .B(n5675), .Z(n5680) );
  NANDN U5955 ( .A(n5678), .B(n5677), .Z(n5679) );
  NAND U5956 ( .A(n5680), .B(n5679), .Z(n5704) );
  AND U5957 ( .A(b[2]), .B(a[241]), .Z(n5710) );
  AND U5958 ( .A(a[242]), .B(b[1]), .Z(n5708) );
  AND U5959 ( .A(a[240]), .B(b[3]), .Z(n5707) );
  XOR U5960 ( .A(n5708), .B(n5707), .Z(n5709) );
  XOR U5961 ( .A(n5710), .B(n5709), .Z(n5713) );
  NAND U5962 ( .A(b[0]), .B(a[243]), .Z(n5714) );
  XOR U5963 ( .A(n5713), .B(n5714), .Z(n5716) );
  OR U5964 ( .A(n5682), .B(n5681), .Z(n5686) );
  NANDN U5965 ( .A(n5684), .B(n5683), .Z(n5685) );
  NAND U5966 ( .A(n5686), .B(n5685), .Z(n5715) );
  XNOR U5967 ( .A(n5716), .B(n5715), .Z(n5701) );
  NANDN U5968 ( .A(n5688), .B(n5687), .Z(n5692) );
  OR U5969 ( .A(n5690), .B(n5689), .Z(n5691) );
  NAND U5970 ( .A(n5692), .B(n5691), .Z(n5702) );
  XNOR U5971 ( .A(n5701), .B(n5702), .Z(n5703) );
  XOR U5972 ( .A(n5704), .B(n5703), .Z(n5700) );
  NANDN U5973 ( .A(sreg[494]), .B(n5693), .Z(n5697) );
  OR U5974 ( .A(n5695), .B(n5694), .Z(n5696) );
  AND U5975 ( .A(n5697), .B(n5696), .Z(n5699) );
  XNOR U5976 ( .A(sreg[495]), .B(n5699), .Z(n5698) );
  XOR U5977 ( .A(n5700), .B(n5698), .Z(c[495]) );
  NANDN U5978 ( .A(n5702), .B(n5701), .Z(n5706) );
  NAND U5979 ( .A(n5704), .B(n5703), .Z(n5705) );
  AND U5980 ( .A(n5706), .B(n5705), .Z(n5727) );
  AND U5981 ( .A(b[2]), .B(a[242]), .Z(n5735) );
  AND U5982 ( .A(a[243]), .B(b[1]), .Z(n5733) );
  AND U5983 ( .A(a[241]), .B(b[3]), .Z(n5732) );
  XOR U5984 ( .A(n5733), .B(n5732), .Z(n5734) );
  XOR U5985 ( .A(n5735), .B(n5734), .Z(n5728) );
  NAND U5986 ( .A(b[0]), .B(a[244]), .Z(n5729) );
  XOR U5987 ( .A(n5728), .B(n5729), .Z(n5730) );
  OR U5988 ( .A(n5708), .B(n5707), .Z(n5712) );
  NANDN U5989 ( .A(n5710), .B(n5709), .Z(n5711) );
  AND U5990 ( .A(n5712), .B(n5711), .Z(n5731) );
  XOR U5991 ( .A(n5730), .B(n5731), .Z(n5725) );
  NANDN U5992 ( .A(n5714), .B(n5713), .Z(n5718) );
  OR U5993 ( .A(n5716), .B(n5715), .Z(n5717) );
  AND U5994 ( .A(n5718), .B(n5717), .Z(n5726) );
  XOR U5995 ( .A(n5725), .B(n5726), .Z(n5719) );
  XOR U5996 ( .A(n5727), .B(n5719), .Z(n5720) );
  XNOR U5997 ( .A(sreg[496]), .B(n5720), .Z(n5721) );
  XOR U5998 ( .A(n5722), .B(n5721), .Z(c[496]) );
  NAND U5999 ( .A(sreg[496]), .B(n5720), .Z(n5724) );
  OR U6000 ( .A(n5722), .B(n5721), .Z(n5723) );
  NAND U6001 ( .A(n5724), .B(n5723), .Z(n5739) );
  AND U6002 ( .A(b[2]), .B(a[243]), .Z(n5744) );
  AND U6003 ( .A(a[244]), .B(b[1]), .Z(n5742) );
  AND U6004 ( .A(a[242]), .B(b[3]), .Z(n5741) );
  XOR U6005 ( .A(n5742), .B(n5741), .Z(n5743) );
  XOR U6006 ( .A(n5744), .B(n5743), .Z(n5747) );
  NAND U6007 ( .A(b[0]), .B(a[245]), .Z(n5748) );
  XNOR U6008 ( .A(n5747), .B(n5748), .Z(n5749) );
  OR U6009 ( .A(n5733), .B(n5732), .Z(n5737) );
  NANDN U6010 ( .A(n5735), .B(n5734), .Z(n5736) );
  AND U6011 ( .A(n5737), .B(n5736), .Z(n5750) );
  XNOR U6012 ( .A(n5749), .B(n5750), .Z(n5754) );
  XNOR U6013 ( .A(n5753), .B(n5754), .Z(n5755) );
  XNOR U6014 ( .A(n5756), .B(n5755), .Z(n5740) );
  XNOR U6015 ( .A(sreg[497]), .B(n5740), .Z(n5738) );
  XNOR U6016 ( .A(n5739), .B(n5738), .Z(c[497]) );
  AND U6017 ( .A(b[2]), .B(a[244]), .Z(n5768) );
  AND U6018 ( .A(a[245]), .B(b[1]), .Z(n5766) );
  AND U6019 ( .A(a[243]), .B(b[3]), .Z(n5765) );
  XOR U6020 ( .A(n5766), .B(n5765), .Z(n5767) );
  XOR U6021 ( .A(n5768), .B(n5767), .Z(n5771) );
  NAND U6022 ( .A(b[0]), .B(a[246]), .Z(n5772) );
  XOR U6023 ( .A(n5771), .B(n5772), .Z(n5774) );
  OR U6024 ( .A(n5742), .B(n5741), .Z(n5746) );
  NANDN U6025 ( .A(n5744), .B(n5743), .Z(n5745) );
  NAND U6026 ( .A(n5746), .B(n5745), .Z(n5773) );
  XNOR U6027 ( .A(n5774), .B(n5773), .Z(n5759) );
  NANDN U6028 ( .A(n5748), .B(n5747), .Z(n5752) );
  NAND U6029 ( .A(n5750), .B(n5749), .Z(n5751) );
  NAND U6030 ( .A(n5752), .B(n5751), .Z(n5760) );
  XNOR U6031 ( .A(n5759), .B(n5760), .Z(n5761) );
  NANDN U6032 ( .A(n5754), .B(n5753), .Z(n5758) );
  NANDN U6033 ( .A(n5756), .B(n5755), .Z(n5757) );
  NAND U6034 ( .A(n5758), .B(n5757), .Z(n5762) );
  XOR U6035 ( .A(n5761), .B(n5762), .Z(n5777) );
  XNOR U6036 ( .A(n5777), .B(sreg[498]), .Z(n5778) );
  XOR U6037 ( .A(n5779), .B(n5778), .Z(c[498]) );
  NANDN U6038 ( .A(n5760), .B(n5759), .Z(n5764) );
  NANDN U6039 ( .A(n5762), .B(n5761), .Z(n5763) );
  NAND U6040 ( .A(n5764), .B(n5763), .Z(n5802) );
  AND U6041 ( .A(b[2]), .B(a[245]), .Z(n5796) );
  AND U6042 ( .A(a[246]), .B(b[1]), .Z(n5794) );
  AND U6043 ( .A(a[244]), .B(b[3]), .Z(n5793) );
  XOR U6044 ( .A(n5794), .B(n5793), .Z(n5795) );
  XOR U6045 ( .A(n5796), .B(n5795), .Z(n5787) );
  NAND U6046 ( .A(b[0]), .B(a[247]), .Z(n5788) );
  XOR U6047 ( .A(n5787), .B(n5788), .Z(n5790) );
  OR U6048 ( .A(n5766), .B(n5765), .Z(n5770) );
  NANDN U6049 ( .A(n5768), .B(n5767), .Z(n5769) );
  NAND U6050 ( .A(n5770), .B(n5769), .Z(n5789) );
  XNOR U6051 ( .A(n5790), .B(n5789), .Z(n5799) );
  NANDN U6052 ( .A(n5772), .B(n5771), .Z(n5776) );
  OR U6053 ( .A(n5774), .B(n5773), .Z(n5775) );
  NAND U6054 ( .A(n5776), .B(n5775), .Z(n5800) );
  XNOR U6055 ( .A(n5799), .B(n5800), .Z(n5801) );
  XNOR U6056 ( .A(n5802), .B(n5801), .Z(n5782) );
  XNOR U6057 ( .A(n5782), .B(sreg[499]), .Z(n5784) );
  NAND U6058 ( .A(n5777), .B(sreg[498]), .Z(n5781) );
  OR U6059 ( .A(n5779), .B(n5778), .Z(n5780) );
  AND U6060 ( .A(n5781), .B(n5780), .Z(n5783) );
  XOR U6061 ( .A(n5784), .B(n5783), .Z(c[499]) );
  NAND U6062 ( .A(n5782), .B(sreg[499]), .Z(n5786) );
  OR U6063 ( .A(n5784), .B(n5783), .Z(n5785) );
  NAND U6064 ( .A(n5786), .B(n5785), .Z(n5824) );
  NANDN U6065 ( .A(n5788), .B(n5787), .Z(n5792) );
  OR U6066 ( .A(n5790), .B(n5789), .Z(n5791) );
  NAND U6067 ( .A(n5792), .B(n5791), .Z(n5806) );
  AND U6068 ( .A(b[2]), .B(a[246]), .Z(n5815) );
  AND U6069 ( .A(a[247]), .B(b[1]), .Z(n5813) );
  AND U6070 ( .A(a[245]), .B(b[3]), .Z(n5812) );
  XOR U6071 ( .A(n5813), .B(n5812), .Z(n5814) );
  XOR U6072 ( .A(n5815), .B(n5814), .Z(n5818) );
  NAND U6073 ( .A(b[0]), .B(a[248]), .Z(n5819) );
  XNOR U6074 ( .A(n5818), .B(n5819), .Z(n5820) );
  OR U6075 ( .A(n5794), .B(n5793), .Z(n5798) );
  NANDN U6076 ( .A(n5796), .B(n5795), .Z(n5797) );
  AND U6077 ( .A(n5798), .B(n5797), .Z(n5821) );
  XNOR U6078 ( .A(n5820), .B(n5821), .Z(n5807) );
  XNOR U6079 ( .A(n5806), .B(n5807), .Z(n5808) );
  NANDN U6080 ( .A(n5800), .B(n5799), .Z(n5804) );
  NAND U6081 ( .A(n5802), .B(n5801), .Z(n5803) );
  AND U6082 ( .A(n5804), .B(n5803), .Z(n5809) );
  XNOR U6083 ( .A(n5808), .B(n5809), .Z(n5825) );
  XOR U6084 ( .A(sreg[500]), .B(n5825), .Z(n5805) );
  XNOR U6085 ( .A(n5824), .B(n5805), .Z(c[500]) );
  NANDN U6086 ( .A(n5807), .B(n5806), .Z(n5811) );
  NAND U6087 ( .A(n5809), .B(n5808), .Z(n5810) );
  NAND U6088 ( .A(n5811), .B(n5810), .Z(n5832) );
  AND U6089 ( .A(b[2]), .B(a[247]), .Z(n5838) );
  AND U6090 ( .A(a[248]), .B(b[1]), .Z(n5836) );
  AND U6091 ( .A(a[246]), .B(b[3]), .Z(n5835) );
  XOR U6092 ( .A(n5836), .B(n5835), .Z(n5837) );
  XOR U6093 ( .A(n5838), .B(n5837), .Z(n5841) );
  NAND U6094 ( .A(b[0]), .B(a[249]), .Z(n5842) );
  XOR U6095 ( .A(n5841), .B(n5842), .Z(n5844) );
  OR U6096 ( .A(n5813), .B(n5812), .Z(n5817) );
  NANDN U6097 ( .A(n5815), .B(n5814), .Z(n5816) );
  NAND U6098 ( .A(n5817), .B(n5816), .Z(n5843) );
  XNOR U6099 ( .A(n5844), .B(n5843), .Z(n5829) );
  NANDN U6100 ( .A(n5819), .B(n5818), .Z(n5823) );
  NAND U6101 ( .A(n5821), .B(n5820), .Z(n5822) );
  NAND U6102 ( .A(n5823), .B(n5822), .Z(n5830) );
  XNOR U6103 ( .A(n5829), .B(n5830), .Z(n5831) );
  XNOR U6104 ( .A(n5832), .B(n5831), .Z(n5828) );
  XOR U6105 ( .A(n5827), .B(sreg[501]), .Z(n5826) );
  XNOR U6106 ( .A(n5828), .B(n5826), .Z(c[501]) );
  NANDN U6107 ( .A(n5830), .B(n5829), .Z(n5834) );
  NANDN U6108 ( .A(n5832), .B(n5831), .Z(n5833) );
  NAND U6109 ( .A(n5834), .B(n5833), .Z(n5850) );
  AND U6110 ( .A(b[2]), .B(a[248]), .Z(n5856) );
  AND U6111 ( .A(a[249]), .B(b[1]), .Z(n5854) );
  AND U6112 ( .A(a[247]), .B(b[3]), .Z(n5853) );
  XOR U6113 ( .A(n5854), .B(n5853), .Z(n5855) );
  XOR U6114 ( .A(n5856), .B(n5855), .Z(n5859) );
  NAND U6115 ( .A(b[0]), .B(a[250]), .Z(n5860) );
  XOR U6116 ( .A(n5859), .B(n5860), .Z(n5862) );
  OR U6117 ( .A(n5836), .B(n5835), .Z(n5840) );
  NANDN U6118 ( .A(n5838), .B(n5837), .Z(n5839) );
  NAND U6119 ( .A(n5840), .B(n5839), .Z(n5861) );
  XNOR U6120 ( .A(n5862), .B(n5861), .Z(n5847) );
  NANDN U6121 ( .A(n5842), .B(n5841), .Z(n5846) );
  OR U6122 ( .A(n5844), .B(n5843), .Z(n5845) );
  NAND U6123 ( .A(n5846), .B(n5845), .Z(n5848) );
  XNOR U6124 ( .A(n5847), .B(n5848), .Z(n5849) );
  XNOR U6125 ( .A(n5850), .B(n5849), .Z(n5865) );
  XNOR U6126 ( .A(n5865), .B(sreg[502]), .Z(n5867) );
  XNOR U6127 ( .A(n5866), .B(n5867), .Z(c[502]) );
  NANDN U6128 ( .A(n5848), .B(n5847), .Z(n5852) );
  NAND U6129 ( .A(n5850), .B(n5849), .Z(n5851) );
  NAND U6130 ( .A(n5852), .B(n5851), .Z(n5876) );
  AND U6131 ( .A(b[2]), .B(a[249]), .Z(n5882) );
  AND U6132 ( .A(a[250]), .B(b[1]), .Z(n5880) );
  AND U6133 ( .A(a[248]), .B(b[3]), .Z(n5879) );
  XOR U6134 ( .A(n5880), .B(n5879), .Z(n5881) );
  XOR U6135 ( .A(n5882), .B(n5881), .Z(n5885) );
  NAND U6136 ( .A(a[251]), .B(b[0]), .Z(n5886) );
  XOR U6137 ( .A(n5885), .B(n5886), .Z(n5888) );
  OR U6138 ( .A(n5854), .B(n5853), .Z(n5858) );
  NANDN U6139 ( .A(n5856), .B(n5855), .Z(n5857) );
  NAND U6140 ( .A(n5858), .B(n5857), .Z(n5887) );
  XNOR U6141 ( .A(n5888), .B(n5887), .Z(n5873) );
  NANDN U6142 ( .A(n5860), .B(n5859), .Z(n5864) );
  OR U6143 ( .A(n5862), .B(n5861), .Z(n5863) );
  NAND U6144 ( .A(n5864), .B(n5863), .Z(n5874) );
  XNOR U6145 ( .A(n5873), .B(n5874), .Z(n5875) );
  XNOR U6146 ( .A(n5876), .B(n5875), .Z(n5872) );
  NAND U6147 ( .A(n5865), .B(sreg[502]), .Z(n5869) );
  NANDN U6148 ( .A(n5867), .B(n5866), .Z(n5868) );
  AND U6149 ( .A(n5869), .B(n5868), .Z(n5871) );
  XNOR U6150 ( .A(n5871), .B(sreg[503]), .Z(n5870) );
  XOR U6151 ( .A(n5872), .B(n5870), .Z(c[503]) );
  NANDN U6152 ( .A(n5874), .B(n5873), .Z(n5878) );
  NAND U6153 ( .A(n5876), .B(n5875), .Z(n5877) );
  NAND U6154 ( .A(n5878), .B(n5877), .Z(n5894) );
  AND U6155 ( .A(b[2]), .B(a[250]), .Z(n5899) );
  IV U6156 ( .A(a[251]), .Z(n5916) );
  NANDN U6157 ( .A(n5916), .B(b[1]), .Z(n5898) );
  NANDN U6158 ( .A(n400), .B(a[249]), .Z(n5897) );
  XNOR U6159 ( .A(n5898), .B(n5897), .Z(n5900) );
  XOR U6160 ( .A(n5899), .B(n5900), .Z(n5903) );
  NAND U6161 ( .A(b[0]), .B(a[252]), .Z(n5904) );
  XOR U6162 ( .A(n5903), .B(n5904), .Z(n5905) );
  OR U6163 ( .A(n5880), .B(n5879), .Z(n5884) );
  NANDN U6164 ( .A(n5882), .B(n5881), .Z(n5883) );
  NAND U6165 ( .A(n5884), .B(n5883), .Z(n5906) );
  XOR U6166 ( .A(n5905), .B(n5906), .Z(n5891) );
  NANDN U6167 ( .A(n5886), .B(n5885), .Z(n5890) );
  OR U6168 ( .A(n5888), .B(n5887), .Z(n5889) );
  NAND U6169 ( .A(n5890), .B(n5889), .Z(n5892) );
  XNOR U6170 ( .A(n5891), .B(n5892), .Z(n5893) );
  XOR U6171 ( .A(n5894), .B(n5893), .Z(n5907) );
  XOR U6172 ( .A(sreg[504]), .B(n5907), .Z(n5909) );
  XNOR U6173 ( .A(n5908), .B(n5909), .Z(c[504]) );
  NANDN U6174 ( .A(n5892), .B(n5891), .Z(n5896) );
  NAND U6175 ( .A(n5894), .B(n5893), .Z(n5895) );
  NAND U6176 ( .A(n5896), .B(n5895), .Z(n5915) );
  AND U6177 ( .A(b[2]), .B(a[251]), .Z(n5919) );
  AND U6178 ( .A(a[252]), .B(b[1]), .Z(n5960) );
  ANDN U6179 ( .B(a[250]), .A(n400), .Z(n5917) );
  XOR U6180 ( .A(n5960), .B(n5917), .Z(n5918) );
  XOR U6181 ( .A(n5919), .B(n5918), .Z(n5920) );
  NAND U6182 ( .A(b[0]), .B(a[253]), .Z(n5921) );
  XNOR U6183 ( .A(n5920), .B(n5921), .Z(n5922) );
  NAND U6184 ( .A(n5898), .B(n5897), .Z(n5902) );
  OR U6185 ( .A(n5900), .B(n5899), .Z(n5901) );
  AND U6186 ( .A(n5902), .B(n5901), .Z(n5923) );
  XOR U6187 ( .A(n5922), .B(n5923), .Z(n5912) );
  XOR U6188 ( .A(n5912), .B(n5913), .Z(n5914) );
  XOR U6189 ( .A(n5915), .B(n5914), .Z(n5926) );
  XNOR U6190 ( .A(n5926), .B(sreg[505]), .Z(n5928) );
  NANDN U6191 ( .A(n5907), .B(sreg[504]), .Z(n5911) );
  NANDN U6192 ( .A(n5909), .B(n5908), .Z(n5910) );
  AND U6193 ( .A(n5911), .B(n5910), .Z(n5927) );
  XOR U6194 ( .A(n5928), .B(n5927), .Z(c[505]) );
  AND U6195 ( .A(b[2]), .B(a[252]), .Z(n5941) );
  NANDN U6196 ( .A(n399), .B(a[253]), .Z(n5940) );
  NANDN U6197 ( .A(n5916), .B(b[3]), .Z(n5939) );
  XNOR U6198 ( .A(n5940), .B(n5939), .Z(n5942) );
  XOR U6199 ( .A(n5941), .B(n5942), .Z(n5945) );
  NAND U6200 ( .A(b[0]), .B(a[254]), .Z(n5946) );
  XOR U6201 ( .A(n5945), .B(n5946), .Z(n5947) );
  XOR U6202 ( .A(n5947), .B(n5948), .Z(n5934) );
  NANDN U6203 ( .A(n5921), .B(n5920), .Z(n5925) );
  NAND U6204 ( .A(n5923), .B(n5922), .Z(n5924) );
  AND U6205 ( .A(n5925), .B(n5924), .Z(n5935) );
  XOR U6206 ( .A(n5934), .B(n5935), .Z(n5936) );
  XOR U6207 ( .A(n5937), .B(n5936), .Z(n5933) );
  NAND U6208 ( .A(n5926), .B(sreg[505]), .Z(n5930) );
  OR U6209 ( .A(n5928), .B(n5927), .Z(n5929) );
  NAND U6210 ( .A(n5930), .B(n5929), .Z(n5932) );
  XNOR U6211 ( .A(sreg[506]), .B(n5932), .Z(n5931) );
  XNOR U6212 ( .A(n5933), .B(n5931), .Z(c[506]) );
  XOR U6213 ( .A(n5949), .B(sreg[507]), .Z(n5951) );
  AND U6214 ( .A(a[252]), .B(b[3]), .Z(n5938) );
  NAND U6215 ( .A(b[1]), .B(a[254]), .Z(n5981) );
  XOR U6216 ( .A(n5938), .B(n5981), .Z(n5962) );
  NAND U6217 ( .A(a[253]), .B(b[2]), .Z(n5961) );
  XOR U6218 ( .A(n5962), .B(n5961), .Z(n5965) );
  NAND U6219 ( .A(b[0]), .B(a[255]), .Z(n5966) );
  XOR U6220 ( .A(n5965), .B(n5966), .Z(n5967) );
  NAND U6221 ( .A(n5940), .B(n5939), .Z(n5944) );
  OR U6222 ( .A(n5942), .B(n5941), .Z(n5943) );
  AND U6223 ( .A(n5944), .B(n5943), .Z(n5968) );
  XNOR U6224 ( .A(n5967), .B(n5968), .Z(n5955) );
  XNOR U6225 ( .A(n5955), .B(n5954), .Z(n5957) );
  XOR U6226 ( .A(n5956), .B(n5957), .Z(n5950) );
  XOR U6227 ( .A(n5951), .B(n5950), .Z(c[507]) );
  NANDN U6228 ( .A(n5949), .B(sreg[507]), .Z(n5953) );
  OR U6229 ( .A(n5951), .B(n5950), .Z(n5952) );
  AND U6230 ( .A(n5953), .B(n5952), .Z(n5970) );
  NANDN U6231 ( .A(n5955), .B(n5954), .Z(n5959) );
  NAND U6232 ( .A(n5957), .B(n5956), .Z(n5958) );
  NAND U6233 ( .A(n5959), .B(n5958), .Z(n5973) );
  AND U6234 ( .A(a[254]), .B(b[3]), .Z(n5991) );
  NAND U6235 ( .A(n5960), .B(n5991), .Z(n5964) );
  OR U6236 ( .A(n5962), .B(n5961), .Z(n5963) );
  NAND U6237 ( .A(n5964), .B(n5963), .Z(n5980) );
  NAND U6238 ( .A(b[2]), .B(a[254]), .Z(n5990) );
  AND U6239 ( .A(a[255]), .B(b[1]), .Z(n5989) );
  XNOR U6240 ( .A(n5990), .B(n5989), .Z(n5977) );
  NAND U6241 ( .A(b[3]), .B(a[253]), .Z(n5978) );
  XOR U6242 ( .A(n5977), .B(n5978), .Z(n5979) );
  XNOR U6243 ( .A(n5980), .B(n5979), .Z(n5972) );
  XNOR U6244 ( .A(n5972), .B(n5971), .Z(n5974) );
  XOR U6245 ( .A(n5973), .B(n5974), .Z(n5969) );
  XOR U6246 ( .A(n5970), .B(n5969), .Z(c[508]) );
  OR U6247 ( .A(n5970), .B(n5969), .Z(n5995) );
  NANDN U6248 ( .A(n5972), .B(n5971), .Z(n5976) );
  NAND U6249 ( .A(n5974), .B(n5973), .Z(n5975) );
  NAND U6250 ( .A(n5976), .B(n5975), .Z(n5986) );
  AND U6251 ( .A(n5981), .B(a[255]), .Z(n5982) );
  NAND U6252 ( .A(b[2]), .B(n5982), .Z(n5992) );
  XNOR U6253 ( .A(n5991), .B(n5992), .Z(n5984) );
  XOR U6254 ( .A(n5983), .B(n5984), .Z(n5985) );
  XOR U6255 ( .A(n5986), .B(n5985), .Z(n5996) );
  XOR U6256 ( .A(n5995), .B(n5996), .Z(c[509]) );
  NAND U6257 ( .A(n5984), .B(n5983), .Z(n5988) );
  NANDN U6258 ( .A(n5986), .B(n5985), .Z(n5987) );
  NAND U6259 ( .A(n5988), .B(n5987), .Z(n6003) );
  NAND U6260 ( .A(b[3]), .B(a[255]), .Z(n6000) );
  XOR U6261 ( .A(n6003), .B(n6000), .Z(n5998) );
  NANDN U6262 ( .A(n5990), .B(n5989), .Z(n5994) );
  NANDN U6263 ( .A(n5992), .B(n5991), .Z(n5993) );
  NAND U6264 ( .A(n5994), .B(n5993), .Z(n6001) );
  NOR U6265 ( .A(n5996), .B(n5995), .Z(n6002) );
  XOR U6266 ( .A(n6001), .B(n6002), .Z(n5997) );
  XNOR U6267 ( .A(n5998), .B(n5997), .Z(c[510]) );
  XNOR U6268 ( .A(n6002), .B(n6001), .Z(n6004) );
  XNOR U6269 ( .A(n6003), .B(n6004), .Z(n5999) );
  NANDN U6270 ( .A(n6000), .B(n5999), .Z(n6008) );
  OR U6271 ( .A(n6002), .B(n6001), .Z(n6006) );
  OR U6272 ( .A(n6004), .B(n6003), .Z(n6005) );
  NAND U6273 ( .A(n6006), .B(n6005), .Z(n6007) );
  NAND U6274 ( .A(n6008), .B(n6007), .Z(c[511]) );
endmodule

