
module compare_N16384_CC128 ( clk, rst, x, y, g, e );
  input [127:0] x;
  input [127:0] y;
  input clk, rst;
  output g, e;
  wire   ebreg, n4, n5, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651;

  DFF ebreg_reg ( .D(n5), .CLK(clk), .RST(rst), .Q(ebreg) );
  DFF greg_reg ( .D(n4), .CLK(clk), .RST(rst), .Q(g) );
  XNOR U10 ( .A(x[1]), .B(n519), .Z(n8) );
  ANDN U11 ( .B(n8), .A(y[1]), .Z(n9) );
  ANDN U12 ( .B(n520), .A(n9), .Z(n10) );
  NANDN U13 ( .A(n519), .B(x[1]), .Z(n11) );
  NAND U14 ( .A(n10), .B(n11), .Z(n521) );
  NANDN U15 ( .A(n541), .B(n540), .Z(n12) );
  AND U16 ( .A(n542), .B(n12), .Z(n13) );
  ANDN U17 ( .B(n543), .A(n13), .Z(n14) );
  NANDN U18 ( .A(y[21]), .B(x[21]), .Z(n15) );
  AND U19 ( .A(n14), .B(n15), .Z(n16) );
  NANDN U20 ( .A(y[23]), .B(x[23]), .Z(n17) );
  NANDN U21 ( .A(n16), .B(n544), .Z(n18) );
  NAND U22 ( .A(n17), .B(n18), .Z(n19) );
  NANDN U23 ( .A(n19), .B(n545), .Z(n20) );
  AND U24 ( .A(n546), .B(n20), .Z(n21) );
  ANDN U25 ( .B(n547), .A(n21), .Z(n22) );
  NANDN U26 ( .A(y[25]), .B(x[25]), .Z(n23) );
  AND U27 ( .A(n22), .B(n23), .Z(n24) );
  NANDN U28 ( .A(n24), .B(n548), .Z(n25) );
  NANDN U29 ( .A(y[27]), .B(x[27]), .Z(n26) );
  AND U30 ( .A(n25), .B(n26), .Z(n27) );
  NAND U31 ( .A(n549), .B(n27), .Z(n28) );
  NAND U32 ( .A(n550), .B(n28), .Z(n551) );
  AND U33 ( .A(n571), .B(n572), .Z(n29) );
  NANDN U34 ( .A(y[47]), .B(x[47]), .Z(n30) );
  AND U35 ( .A(n29), .B(n30), .Z(n31) );
  NANDN U36 ( .A(y[49]), .B(x[49]), .Z(n32) );
  NANDN U37 ( .A(n31), .B(n573), .Z(n33) );
  NAND U38 ( .A(n32), .B(n33), .Z(n34) );
  NANDN U39 ( .A(n34), .B(n574), .Z(n35) );
  AND U40 ( .A(n575), .B(n35), .Z(n36) );
  ANDN U41 ( .B(n576), .A(n36), .Z(n37) );
  NANDN U42 ( .A(y[51]), .B(x[51]), .Z(n38) );
  AND U43 ( .A(n37), .B(n38), .Z(n39) );
  NANDN U44 ( .A(y[53]), .B(x[53]), .Z(n40) );
  NANDN U45 ( .A(n39), .B(n577), .Z(n41) );
  NAND U46 ( .A(n40), .B(n41), .Z(n42) );
  ANDN U47 ( .B(x[55]), .A(y[55]), .Z(n43) );
  NANDN U48 ( .A(n42), .B(n578), .Z(n44) );
  NAND U49 ( .A(n579), .B(n44), .Z(n45) );
  NANDN U50 ( .A(n43), .B(n45), .Z(n582) );
  OR U51 ( .A(n599), .B(n600), .Z(n46) );
  NAND U52 ( .A(n601), .B(n46), .Z(n47) );
  AND U53 ( .A(n602), .B(n47), .Z(n48) );
  NANDN U54 ( .A(y[75]), .B(x[75]), .Z(n49) );
  NAND U55 ( .A(n48), .B(n49), .Z(n50) );
  NAND U56 ( .A(n603), .B(n50), .Z(n51) );
  AND U57 ( .A(n51), .B(n604), .Z(n52) );
  NANDN U58 ( .A(y[77]), .B(x[77]), .Z(n53) );
  AND U59 ( .A(n52), .B(n53), .Z(n54) );
  NANDN U60 ( .A(n54), .B(n605), .Z(n55) );
  AND U61 ( .A(n515), .B(n55), .Z(n56) );
  NANDN U62 ( .A(y[79]), .B(x[79]), .Z(n57) );
  NAND U63 ( .A(n56), .B(n57), .Z(n58) );
  AND U64 ( .A(n606), .B(n58), .Z(n59) );
  ANDN U65 ( .B(n514), .A(n59), .Z(n60) );
  NANDN U66 ( .A(y[81]), .B(x[81]), .Z(n61) );
  NAND U67 ( .A(n60), .B(n61), .Z(n62) );
  NAND U68 ( .A(n607), .B(n62), .Z(n608) );
  OR U69 ( .A(n626), .B(n627), .Z(n63) );
  NAND U70 ( .A(n628), .B(n63), .Z(n64) );
  AND U71 ( .A(n509), .B(n64), .Z(n65) );
  NANDN U72 ( .A(y[103]), .B(x[103]), .Z(n66) );
  NAND U73 ( .A(n65), .B(n66), .Z(n67) );
  NAND U74 ( .A(n629), .B(n67), .Z(n68) );
  AND U75 ( .A(n68), .B(n508), .Z(n69) );
  NANDN U76 ( .A(y[105]), .B(x[105]), .Z(n70) );
  AND U77 ( .A(n69), .B(n70), .Z(n71) );
  NANDN U78 ( .A(n71), .B(n630), .Z(n72) );
  AND U79 ( .A(n631), .B(n72), .Z(n73) );
  NANDN U80 ( .A(y[107]), .B(x[107]), .Z(n74) );
  NAND U81 ( .A(n73), .B(n74), .Z(n75) );
  AND U82 ( .A(n632), .B(n75), .Z(n76) );
  ANDN U83 ( .B(n633), .A(n76), .Z(n77) );
  NANDN U84 ( .A(y[109]), .B(x[109]), .Z(n78) );
  NAND U85 ( .A(n77), .B(n78), .Z(n79) );
  NAND U86 ( .A(n634), .B(n79), .Z(n635) );
  NAND U87 ( .A(n522), .B(n521), .Z(n80) );
  NANDN U88 ( .A(y[3]), .B(x[3]), .Z(n81) );
  NAND U89 ( .A(n80), .B(n81), .Z(n82) );
  NANDN U90 ( .A(n82), .B(n523), .Z(n83) );
  AND U91 ( .A(n524), .B(n83), .Z(n84) );
  ANDN U92 ( .B(n525), .A(n84), .Z(n85) );
  NANDN U93 ( .A(y[5]), .B(x[5]), .Z(n86) );
  AND U94 ( .A(n85), .B(n86), .Z(n87) );
  NANDN U95 ( .A(y[7]), .B(x[7]), .Z(n88) );
  NANDN U96 ( .A(n87), .B(n526), .Z(n89) );
  NAND U97 ( .A(n88), .B(n89), .Z(n90) );
  NANDN U98 ( .A(n90), .B(n527), .Z(n91) );
  AND U99 ( .A(n528), .B(n91), .Z(n92) );
  ANDN U100 ( .B(n529), .A(n92), .Z(n93) );
  NANDN U101 ( .A(y[9]), .B(x[9]), .Z(n94) );
  NAND U102 ( .A(n93), .B(n94), .Z(n95) );
  NAND U103 ( .A(n530), .B(n95), .Z(n531) );
  AND U104 ( .A(n552), .B(n551), .Z(n96) );
  NANDN U105 ( .A(y[29]), .B(x[29]), .Z(n97) );
  AND U106 ( .A(n96), .B(n97), .Z(n98) );
  NANDN U107 ( .A(y[31]), .B(x[31]), .Z(n99) );
  NANDN U108 ( .A(n98), .B(n553), .Z(n100) );
  NAND U109 ( .A(n99), .B(n100), .Z(n101) );
  NANDN U110 ( .A(n101), .B(n554), .Z(n102) );
  AND U111 ( .A(n555), .B(n102), .Z(n103) );
  ANDN U112 ( .B(n556), .A(n103), .Z(n104) );
  NANDN U113 ( .A(y[33]), .B(x[33]), .Z(n105) );
  AND U114 ( .A(n104), .B(n105), .Z(n106) );
  NANDN U115 ( .A(y[35]), .B(x[35]), .Z(n107) );
  NANDN U116 ( .A(n106), .B(n557), .Z(n108) );
  NAND U117 ( .A(n107), .B(n108), .Z(n109) );
  ANDN U118 ( .B(x[37]), .A(y[37]), .Z(n110) );
  NANDN U119 ( .A(n109), .B(n558), .Z(n111) );
  NAND U120 ( .A(n559), .B(n111), .Z(n112) );
  NANDN U121 ( .A(n110), .B(n112), .Z(n561) );
  OR U122 ( .A(n581), .B(n582), .Z(n113) );
  AND U123 ( .A(n583), .B(n113), .Z(n114) );
  ANDN U124 ( .B(n584), .A(n114), .Z(n115) );
  NANDN U125 ( .A(y[57]), .B(x[57]), .Z(n116) );
  AND U126 ( .A(n115), .B(n116), .Z(n117) );
  NANDN U127 ( .A(y[59]), .B(x[59]), .Z(n118) );
  NANDN U128 ( .A(n117), .B(n585), .Z(n119) );
  NAND U129 ( .A(n118), .B(n119), .Z(n120) );
  NANDN U130 ( .A(n120), .B(n586), .Z(n121) );
  AND U131 ( .A(n587), .B(n121), .Z(n122) );
  ANDN U132 ( .B(n588), .A(n122), .Z(n123) );
  NANDN U133 ( .A(y[61]), .B(x[61]), .Z(n124) );
  AND U134 ( .A(n123), .B(n124), .Z(n125) );
  NANDN U135 ( .A(n125), .B(n589), .Z(n126) );
  NANDN U136 ( .A(y[63]), .B(x[63]), .Z(n127) );
  AND U137 ( .A(n126), .B(n127), .Z(n128) );
  NAND U138 ( .A(n128), .B(n590), .Z(n129) );
  NAND U139 ( .A(n591), .B(n129), .Z(n592) );
  ANDN U140 ( .B(n608), .A(n610), .Z(n130) );
  NAND U141 ( .A(n609), .B(n130), .Z(n131) );
  NAND U142 ( .A(n611), .B(n131), .Z(n132) );
  AND U143 ( .A(n132), .B(n612), .Z(n133) );
  NANDN U144 ( .A(y[85]), .B(x[85]), .Z(n134) );
  AND U145 ( .A(n133), .B(n134), .Z(n135) );
  NANDN U146 ( .A(n135), .B(n613), .Z(n136) );
  AND U147 ( .A(n513), .B(n136), .Z(n137) );
  NANDN U148 ( .A(y[87]), .B(x[87]), .Z(n138) );
  NAND U149 ( .A(n137), .B(n138), .Z(n139) );
  AND U150 ( .A(n614), .B(n139), .Z(n140) );
  ANDN U151 ( .B(n512), .A(n140), .Z(n141) );
  NANDN U152 ( .A(y[89]), .B(x[89]), .Z(n142) );
  NAND U153 ( .A(n141), .B(n142), .Z(n143) );
  AND U154 ( .A(n615), .B(n143), .Z(n144) );
  ANDN U155 ( .B(n616), .A(n144), .Z(n145) );
  NANDN U156 ( .A(y[91]), .B(x[91]), .Z(n146) );
  NAND U157 ( .A(n145), .B(n146), .Z(n617) );
  NOR U158 ( .A(n637), .B(n636), .Z(n147) );
  NAND U159 ( .A(n635), .B(n147), .Z(n148) );
  NAND U160 ( .A(n638), .B(n148), .Z(n149) );
  AND U161 ( .A(n149), .B(n506), .Z(n150) );
  NANDN U162 ( .A(y[113]), .B(x[113]), .Z(n151) );
  AND U163 ( .A(n150), .B(n151), .Z(n152) );
  NANDN U164 ( .A(n152), .B(n639), .Z(n153) );
  AND U165 ( .A(n640), .B(n153), .Z(n154) );
  NANDN U166 ( .A(y[115]), .B(x[115]), .Z(n155) );
  NAND U167 ( .A(n154), .B(n155), .Z(n156) );
  AND U168 ( .A(n641), .B(n156), .Z(n157) );
  ANDN U169 ( .B(n642), .A(n157), .Z(n158) );
  NANDN U170 ( .A(y[117]), .B(x[117]), .Z(n159) );
  NAND U171 ( .A(n158), .B(n159), .Z(n160) );
  AND U172 ( .A(n643), .B(n160), .Z(n161) );
  ANDN U173 ( .B(n505), .A(n161), .Z(n162) );
  NANDN U174 ( .A(y[119]), .B(x[119]), .Z(n163) );
  NAND U175 ( .A(n162), .B(n163), .Z(n644) );
  AND U176 ( .A(n532), .B(n531), .Z(n164) );
  NANDN U177 ( .A(y[11]), .B(x[11]), .Z(n165) );
  AND U178 ( .A(n164), .B(n165), .Z(n166) );
  NANDN U179 ( .A(y[13]), .B(x[13]), .Z(n167) );
  NANDN U180 ( .A(n166), .B(n533), .Z(n168) );
  NAND U181 ( .A(n167), .B(n168), .Z(n169) );
  NANDN U182 ( .A(n169), .B(n534), .Z(n170) );
  AND U183 ( .A(n535), .B(n170), .Z(n171) );
  ANDN U184 ( .B(n536), .A(n171), .Z(n172) );
  NANDN U185 ( .A(y[15]), .B(x[15]), .Z(n173) );
  AND U186 ( .A(n172), .B(n173), .Z(n174) );
  NANDN U187 ( .A(n174), .B(n537), .Z(n175) );
  NANDN U188 ( .A(y[17]), .B(x[17]), .Z(n176) );
  AND U189 ( .A(n175), .B(n176), .Z(n177) );
  ANDN U190 ( .B(x[19]), .A(y[19]), .Z(n178) );
  NAND U191 ( .A(n538), .B(n177), .Z(n179) );
  NAND U192 ( .A(n539), .B(n179), .Z(n180) );
  NANDN U193 ( .A(n178), .B(n180), .Z(n541) );
  NANDN U194 ( .A(n561), .B(n560), .Z(n181) );
  AND U195 ( .A(n562), .B(n181), .Z(n182) );
  ANDN U196 ( .B(n563), .A(n182), .Z(n183) );
  NANDN U197 ( .A(y[39]), .B(x[39]), .Z(n184) );
  AND U198 ( .A(n183), .B(n184), .Z(n185) );
  NANDN U199 ( .A(y[41]), .B(x[41]), .Z(n186) );
  NANDN U200 ( .A(n185), .B(n564), .Z(n187) );
  NAND U201 ( .A(n186), .B(n187), .Z(n188) );
  NANDN U202 ( .A(n188), .B(n565), .Z(n189) );
  AND U203 ( .A(n566), .B(n189), .Z(n190) );
  ANDN U204 ( .B(n567), .A(n190), .Z(n191) );
  NANDN U205 ( .A(y[43]), .B(x[43]), .Z(n192) );
  AND U206 ( .A(n191), .B(n192), .Z(n193) );
  NANDN U207 ( .A(n193), .B(n568), .Z(n194) );
  NANDN U208 ( .A(y[45]), .B(x[45]), .Z(n195) );
  AND U209 ( .A(n194), .B(n195), .Z(n196) );
  NAND U210 ( .A(n569), .B(n196), .Z(n197) );
  NAND U211 ( .A(n570), .B(n197), .Z(n571) );
  AND U212 ( .A(n518), .B(n592), .Z(n198) );
  NANDN U213 ( .A(y[65]), .B(x[65]), .Z(n199) );
  AND U214 ( .A(n198), .B(n199), .Z(n200) );
  NANDN U215 ( .A(n200), .B(n593), .Z(n201) );
  AND U216 ( .A(n594), .B(n201), .Z(n202) );
  NANDN U217 ( .A(y[67]), .B(x[67]), .Z(n203) );
  NAND U218 ( .A(n202), .B(n203), .Z(n204) );
  NAND U219 ( .A(n595), .B(n204), .Z(n205) );
  AND U220 ( .A(n205), .B(n596), .Z(n206) );
  NANDN U221 ( .A(y[69]), .B(x[69]), .Z(n207) );
  AND U222 ( .A(n206), .B(n207), .Z(n208) );
  NANDN U223 ( .A(n208), .B(n597), .Z(n209) );
  AND U224 ( .A(n517), .B(n209), .Z(n210) );
  NANDN U225 ( .A(y[71]), .B(x[71]), .Z(n211) );
  NAND U226 ( .A(n210), .B(n211), .Z(n212) );
  NAND U227 ( .A(n598), .B(n212), .Z(n213) );
  NAND U228 ( .A(n516), .B(n213), .Z(n600) );
  NAND U229 ( .A(n617), .B(n618), .Z(n214) );
  AND U230 ( .A(n619), .B(n214), .Z(n215) );
  NANDN U231 ( .A(y[93]), .B(x[93]), .Z(n216) );
  NAND U232 ( .A(n215), .B(n216), .Z(n217) );
  NAND U233 ( .A(n620), .B(n217), .Z(n218) );
  AND U234 ( .A(n218), .B(n511), .Z(n219) );
  NANDN U235 ( .A(y[95]), .B(x[95]), .Z(n220) );
  AND U236 ( .A(n219), .B(n220), .Z(n221) );
  NANDN U237 ( .A(n221), .B(n621), .Z(n222) );
  AND U238 ( .A(n510), .B(n222), .Z(n223) );
  NANDN U239 ( .A(y[97]), .B(x[97]), .Z(n224) );
  NAND U240 ( .A(n223), .B(n224), .Z(n225) );
  AND U241 ( .A(n622), .B(n225), .Z(n226) );
  ANDN U242 ( .B(n623), .A(n226), .Z(n227) );
  NANDN U243 ( .A(y[99]), .B(x[99]), .Z(n228) );
  NAND U244 ( .A(n227), .B(n228), .Z(n229) );
  NAND U245 ( .A(n624), .B(n229), .Z(n230) );
  NAND U246 ( .A(n625), .B(n230), .Z(n627) );
  AND U247 ( .A(e), .B(n651), .Z(n231) );
  NAND U248 ( .A(n645), .B(n644), .Z(n232) );
  AND U249 ( .A(n504), .B(n232), .Z(n233) );
  NANDN U250 ( .A(y[121]), .B(x[121]), .Z(n234) );
  NAND U251 ( .A(n233), .B(n234), .Z(n235) );
  NAND U252 ( .A(n646), .B(n235), .Z(n236) );
  AND U253 ( .A(n236), .B(n647), .Z(n237) );
  NANDN U254 ( .A(y[123]), .B(x[123]), .Z(n238) );
  AND U255 ( .A(n237), .B(n238), .Z(n239) );
  NANDN U256 ( .A(n239), .B(n648), .Z(n240) );
  AND U257 ( .A(n649), .B(n240), .Z(n241) );
  NANDN U258 ( .A(y[125]), .B(x[125]), .Z(n242) );
  AND U259 ( .A(n241), .B(n242), .Z(n243) );
  NANDN U260 ( .A(y[127]), .B(x[127]), .Z(n244) );
  NANDN U261 ( .A(n243), .B(n650), .Z(n245) );
  NAND U262 ( .A(n244), .B(n245), .Z(n246) );
  NAND U263 ( .A(n246), .B(n231), .Z(n247) );
  NANDN U264 ( .A(n231), .B(g), .Z(n248) );
  NAND U265 ( .A(n247), .B(n248), .Z(n4) );
  IV U266 ( .A(ebreg), .Z(e) );
  XNOR U267 ( .A(x[95]), .B(y[95]), .Z(n250) );
  NANDN U268 ( .A(x[94]), .B(y[94]), .Z(n249) );
  AND U269 ( .A(n250), .B(n249), .Z(n620) );
  XNOR U270 ( .A(x[89]), .B(y[89]), .Z(n252) );
  NANDN U271 ( .A(x[88]), .B(y[88]), .Z(n251) );
  AND U272 ( .A(n252), .B(n251), .Z(n614) );
  AND U273 ( .A(n620), .B(n614), .Z(n258) );
  XNOR U274 ( .A(x[93]), .B(y[93]), .Z(n254) );
  NANDN U275 ( .A(x[92]), .B(y[92]), .Z(n253) );
  AND U276 ( .A(n254), .B(n253), .Z(n618) );
  XNOR U277 ( .A(x[91]), .B(y[91]), .Z(n256) );
  NANDN U278 ( .A(x[90]), .B(y[90]), .Z(n255) );
  AND U279 ( .A(n256), .B(n255), .Z(n615) );
  AND U280 ( .A(n618), .B(n615), .Z(n257) );
  AND U281 ( .A(n258), .B(n257), .Z(n270) );
  XNOR U282 ( .A(x[71]), .B(y[71]), .Z(n260) );
  NANDN U283 ( .A(x[70]), .B(y[70]), .Z(n259) );
  AND U284 ( .A(n260), .B(n259), .Z(n597) );
  XNOR U285 ( .A(x[65]), .B(y[65]), .Z(n262) );
  NANDN U286 ( .A(x[64]), .B(y[64]), .Z(n261) );
  AND U287 ( .A(n262), .B(n261), .Z(n591) );
  AND U288 ( .A(n597), .B(n591), .Z(n268) );
  XNOR U289 ( .A(x[69]), .B(y[69]), .Z(n264) );
  NANDN U290 ( .A(x[68]), .B(y[68]), .Z(n263) );
  AND U291 ( .A(n264), .B(n263), .Z(n595) );
  XNOR U292 ( .A(x[67]), .B(y[67]), .Z(n266) );
  NANDN U293 ( .A(x[66]), .B(y[66]), .Z(n265) );
  AND U294 ( .A(n266), .B(n265), .Z(n593) );
  AND U295 ( .A(n595), .B(n593), .Z(n267) );
  AND U296 ( .A(n268), .B(n267), .Z(n269) );
  AND U297 ( .A(n270), .B(n269), .Z(n294) );
  XNOR U298 ( .A(x[87]), .B(y[87]), .Z(n272) );
  NANDN U299 ( .A(x[86]), .B(y[86]), .Z(n271) );
  AND U300 ( .A(n272), .B(n271), .Z(n613) );
  XNOR U301 ( .A(x[81]), .B(y[81]), .Z(n274) );
  NANDN U302 ( .A(x[80]), .B(y[80]), .Z(n273) );
  AND U303 ( .A(n274), .B(n273), .Z(n606) );
  AND U304 ( .A(n613), .B(n606), .Z(n280) );
  XNOR U305 ( .A(x[85]), .B(y[85]), .Z(n276) );
  NANDN U306 ( .A(x[84]), .B(y[84]), .Z(n275) );
  AND U307 ( .A(n276), .B(n275), .Z(n611) );
  XNOR U308 ( .A(x[83]), .B(y[83]), .Z(n278) );
  NANDN U309 ( .A(x[82]), .B(y[82]), .Z(n277) );
  AND U310 ( .A(n278), .B(n277), .Z(n607) );
  AND U311 ( .A(n611), .B(n607), .Z(n279) );
  AND U312 ( .A(n280), .B(n279), .Z(n292) );
  XNOR U313 ( .A(x[79]), .B(y[79]), .Z(n282) );
  NANDN U314 ( .A(x[78]), .B(y[78]), .Z(n281) );
  AND U315 ( .A(n282), .B(n281), .Z(n605) );
  XNOR U316 ( .A(x[73]), .B(y[73]), .Z(n284) );
  NANDN U317 ( .A(x[72]), .B(y[72]), .Z(n283) );
  AND U318 ( .A(n284), .B(n283), .Z(n598) );
  AND U319 ( .A(n605), .B(n598), .Z(n290) );
  XNOR U320 ( .A(x[77]), .B(y[77]), .Z(n286) );
  NANDN U321 ( .A(x[76]), .B(y[76]), .Z(n285) );
  AND U322 ( .A(n286), .B(n285), .Z(n603) );
  XNOR U323 ( .A(x[75]), .B(y[75]), .Z(n288) );
  NANDN U324 ( .A(x[74]), .B(y[74]), .Z(n287) );
  AND U325 ( .A(n288), .B(n287), .Z(n601) );
  AND U326 ( .A(n603), .B(n601), .Z(n289) );
  AND U327 ( .A(n290), .B(n289), .Z(n291) );
  AND U328 ( .A(n292), .B(n291), .Z(n293) );
  AND U329 ( .A(n294), .B(n293), .Z(n503) );
  XNOR U330 ( .A(y[23]), .B(x[23]), .Z(n296) );
  NANDN U331 ( .A(x[22]), .B(y[22]), .Z(n295) );
  AND U332 ( .A(n296), .B(n295), .Z(n544) );
  XNOR U333 ( .A(y[17]), .B(x[17]), .Z(n298) );
  NANDN U334 ( .A(x[16]), .B(y[16]), .Z(n297) );
  AND U335 ( .A(n298), .B(n297), .Z(n537) );
  AND U336 ( .A(n544), .B(n537), .Z(n304) );
  XNOR U337 ( .A(y[21]), .B(x[21]), .Z(n300) );
  NANDN U338 ( .A(x[20]), .B(y[20]), .Z(n299) );
  AND U339 ( .A(n300), .B(n299), .Z(n542) );
  XNOR U340 ( .A(y[19]), .B(x[19]), .Z(n302) );
  NANDN U341 ( .A(x[18]), .B(y[18]), .Z(n301) );
  AND U342 ( .A(n302), .B(n301), .Z(n539) );
  AND U343 ( .A(n542), .B(n539), .Z(n303) );
  AND U344 ( .A(n304), .B(n303), .Z(n317) );
  XNOR U345 ( .A(y[1]), .B(x[1]), .Z(n306) );
  NANDN U346 ( .A(x[0]), .B(y[0]), .Z(n305) );
  AND U347 ( .A(n306), .B(n305), .Z(n309) );
  XNOR U348 ( .A(y[13]), .B(x[13]), .Z(n308) );
  NANDN U349 ( .A(x[12]), .B(y[12]), .Z(n307) );
  AND U350 ( .A(n308), .B(n307), .Z(n533) );
  AND U351 ( .A(n309), .B(n533), .Z(n315) );
  XNOR U352 ( .A(y[3]), .B(x[3]), .Z(n311) );
  NANDN U353 ( .A(x[2]), .B(y[2]), .Z(n310) );
  AND U354 ( .A(n311), .B(n310), .Z(n522) );
  XNOR U355 ( .A(y[15]), .B(x[15]), .Z(n313) );
  NANDN U356 ( .A(x[14]), .B(y[14]), .Z(n312) );
  AND U357 ( .A(n313), .B(n312), .Z(n535) );
  AND U358 ( .A(n522), .B(n535), .Z(n314) );
  AND U359 ( .A(n315), .B(n314), .Z(n316) );
  AND U360 ( .A(n317), .B(n316), .Z(n341) );
  XNOR U361 ( .A(y[31]), .B(x[31]), .Z(n319) );
  NANDN U362 ( .A(x[30]), .B(y[30]), .Z(n318) );
  AND U363 ( .A(n319), .B(n318), .Z(n553) );
  XNOR U364 ( .A(y[25]), .B(x[25]), .Z(n321) );
  NANDN U365 ( .A(x[24]), .B(y[24]), .Z(n320) );
  AND U366 ( .A(n321), .B(n320), .Z(n546) );
  AND U367 ( .A(n553), .B(n546), .Z(n327) );
  XNOR U368 ( .A(y[29]), .B(x[29]), .Z(n323) );
  NANDN U369 ( .A(x[28]), .B(y[28]), .Z(n322) );
  AND U370 ( .A(n323), .B(n322), .Z(n550) );
  XNOR U371 ( .A(y[27]), .B(x[27]), .Z(n325) );
  NANDN U372 ( .A(x[26]), .B(y[26]), .Z(n324) );
  AND U373 ( .A(n325), .B(n324), .Z(n548) );
  AND U374 ( .A(n550), .B(n548), .Z(n326) );
  AND U375 ( .A(n327), .B(n326), .Z(n339) );
  XNOR U376 ( .A(y[11]), .B(x[11]), .Z(n329) );
  NANDN U377 ( .A(x[10]), .B(y[10]), .Z(n328) );
  AND U378 ( .A(n329), .B(n328), .Z(n530) );
  XNOR U379 ( .A(y[5]), .B(x[5]), .Z(n331) );
  NANDN U380 ( .A(x[4]), .B(y[4]), .Z(n330) );
  AND U381 ( .A(n331), .B(n330), .Z(n524) );
  AND U382 ( .A(n530), .B(n524), .Z(n337) );
  XNOR U383 ( .A(y[9]), .B(x[9]), .Z(n333) );
  NANDN U384 ( .A(x[8]), .B(y[8]), .Z(n332) );
  AND U385 ( .A(n333), .B(n332), .Z(n528) );
  XNOR U386 ( .A(y[7]), .B(x[7]), .Z(n335) );
  NANDN U387 ( .A(x[6]), .B(y[6]), .Z(n334) );
  AND U388 ( .A(n335), .B(n334), .Z(n526) );
  AND U389 ( .A(n528), .B(n526), .Z(n336) );
  AND U390 ( .A(n337), .B(n336), .Z(n338) );
  AND U391 ( .A(n339), .B(n338), .Z(n340) );
  AND U392 ( .A(n341), .B(n340), .Z(n389) );
  XNOR U393 ( .A(x[127]), .B(y[127]), .Z(n343) );
  NANDN U394 ( .A(x[126]), .B(y[126]), .Z(n342) );
  AND U395 ( .A(n343), .B(n342), .Z(n650) );
  XNOR U396 ( .A(x[121]), .B(y[121]), .Z(n345) );
  NANDN U397 ( .A(x[120]), .B(y[120]), .Z(n344) );
  AND U398 ( .A(n345), .B(n344), .Z(n645) );
  AND U399 ( .A(n650), .B(n645), .Z(n351) );
  XNOR U400 ( .A(x[125]), .B(y[125]), .Z(n347) );
  NANDN U401 ( .A(x[124]), .B(y[124]), .Z(n346) );
  AND U402 ( .A(n347), .B(n346), .Z(n648) );
  XNOR U403 ( .A(x[123]), .B(y[123]), .Z(n349) );
  NANDN U404 ( .A(x[122]), .B(y[122]), .Z(n348) );
  AND U405 ( .A(n349), .B(n348), .Z(n646) );
  AND U406 ( .A(n648), .B(n646), .Z(n350) );
  AND U407 ( .A(n351), .B(n350), .Z(n363) );
  XNOR U408 ( .A(x[103]), .B(y[103]), .Z(n353) );
  NANDN U409 ( .A(x[102]), .B(y[102]), .Z(n352) );
  AND U410 ( .A(n353), .B(n352), .Z(n628) );
  XNOR U411 ( .A(x[97]), .B(y[97]), .Z(n355) );
  NANDN U412 ( .A(x[96]), .B(y[96]), .Z(n354) );
  AND U413 ( .A(n355), .B(n354), .Z(n621) );
  AND U414 ( .A(n628), .B(n621), .Z(n361) );
  XNOR U415 ( .A(x[101]), .B(y[101]), .Z(n357) );
  NANDN U416 ( .A(x[100]), .B(y[100]), .Z(n356) );
  AND U417 ( .A(n357), .B(n356), .Z(n624) );
  XNOR U418 ( .A(x[99]), .B(y[99]), .Z(n359) );
  NANDN U419 ( .A(x[98]), .B(y[98]), .Z(n358) );
  AND U420 ( .A(n359), .B(n358), .Z(n622) );
  AND U421 ( .A(n624), .B(n622), .Z(n360) );
  AND U422 ( .A(n361), .B(n360), .Z(n362) );
  AND U423 ( .A(n363), .B(n362), .Z(n387) );
  XNOR U424 ( .A(x[119]), .B(y[119]), .Z(n365) );
  NANDN U425 ( .A(x[118]), .B(y[118]), .Z(n364) );
  AND U426 ( .A(n365), .B(n364), .Z(n643) );
  XNOR U427 ( .A(x[113]), .B(y[113]), .Z(n367) );
  NANDN U428 ( .A(x[112]), .B(y[112]), .Z(n366) );
  AND U429 ( .A(n367), .B(n366), .Z(n638) );
  AND U430 ( .A(n643), .B(n638), .Z(n373) );
  XNOR U431 ( .A(x[117]), .B(y[117]), .Z(n369) );
  NANDN U432 ( .A(x[116]), .B(y[116]), .Z(n368) );
  AND U433 ( .A(n369), .B(n368), .Z(n641) );
  XNOR U434 ( .A(x[115]), .B(y[115]), .Z(n371) );
  NANDN U435 ( .A(x[114]), .B(y[114]), .Z(n370) );
  AND U436 ( .A(n371), .B(n370), .Z(n639) );
  AND U437 ( .A(n641), .B(n639), .Z(n372) );
  AND U438 ( .A(n373), .B(n372), .Z(n385) );
  XNOR U439 ( .A(x[111]), .B(y[111]), .Z(n375) );
  NANDN U440 ( .A(x[110]), .B(y[110]), .Z(n374) );
  AND U441 ( .A(n375), .B(n374), .Z(n634) );
  XNOR U442 ( .A(x[105]), .B(y[105]), .Z(n377) );
  NANDN U443 ( .A(x[104]), .B(y[104]), .Z(n376) );
  AND U444 ( .A(n377), .B(n376), .Z(n629) );
  AND U445 ( .A(n634), .B(n629), .Z(n383) );
  XNOR U446 ( .A(x[109]), .B(y[109]), .Z(n379) );
  NANDN U447 ( .A(x[108]), .B(y[108]), .Z(n378) );
  AND U448 ( .A(n379), .B(n378), .Z(n632) );
  XNOR U449 ( .A(x[107]), .B(y[107]), .Z(n381) );
  NANDN U450 ( .A(x[106]), .B(y[106]), .Z(n380) );
  AND U451 ( .A(n381), .B(n380), .Z(n630) );
  AND U452 ( .A(n632), .B(n630), .Z(n382) );
  AND U453 ( .A(n383), .B(n382), .Z(n384) );
  AND U454 ( .A(n385), .B(n384), .Z(n386) );
  AND U455 ( .A(n387), .B(n386), .Z(n388) );
  AND U456 ( .A(n389), .B(n388), .Z(n501) );
  XNOR U457 ( .A(y[55]), .B(x[55]), .Z(n391) );
  NANDN U458 ( .A(x[54]), .B(y[54]), .Z(n390) );
  AND U459 ( .A(n391), .B(n390), .Z(n579) );
  XNOR U460 ( .A(y[49]), .B(x[49]), .Z(n393) );
  NANDN U461 ( .A(x[48]), .B(y[48]), .Z(n392) );
  AND U462 ( .A(n393), .B(n392), .Z(n573) );
  AND U463 ( .A(n579), .B(n573), .Z(n399) );
  XNOR U464 ( .A(y[53]), .B(x[53]), .Z(n395) );
  NANDN U465 ( .A(x[52]), .B(y[52]), .Z(n394) );
  AND U466 ( .A(n395), .B(n394), .Z(n577) );
  XNOR U467 ( .A(y[51]), .B(x[51]), .Z(n397) );
  NANDN U468 ( .A(x[50]), .B(y[50]), .Z(n396) );
  AND U469 ( .A(n397), .B(n396), .Z(n575) );
  AND U470 ( .A(n577), .B(n575), .Z(n398) );
  AND U471 ( .A(n399), .B(n398), .Z(n411) );
  XNOR U472 ( .A(y[47]), .B(x[47]), .Z(n401) );
  NANDN U473 ( .A(x[46]), .B(y[46]), .Z(n400) );
  AND U474 ( .A(n401), .B(n400), .Z(n570) );
  XNOR U475 ( .A(y[41]), .B(x[41]), .Z(n403) );
  NANDN U476 ( .A(x[40]), .B(y[40]), .Z(n402) );
  AND U477 ( .A(n403), .B(n402), .Z(n564) );
  AND U478 ( .A(n570), .B(n564), .Z(n409) );
  XNOR U479 ( .A(y[45]), .B(x[45]), .Z(n405) );
  NANDN U480 ( .A(x[44]), .B(y[44]), .Z(n404) );
  AND U481 ( .A(n405), .B(n404), .Z(n568) );
  XNOR U482 ( .A(y[43]), .B(x[43]), .Z(n407) );
  NANDN U483 ( .A(x[42]), .B(y[42]), .Z(n406) );
  AND U484 ( .A(n407), .B(n406), .Z(n566) );
  AND U485 ( .A(n568), .B(n566), .Z(n408) );
  AND U486 ( .A(n409), .B(n408), .Z(n410) );
  AND U487 ( .A(n411), .B(n410), .Z(n435) );
  XNOR U488 ( .A(y[63]), .B(x[63]), .Z(n413) );
  NANDN U489 ( .A(x[62]), .B(y[62]), .Z(n412) );
  AND U490 ( .A(n413), .B(n412), .Z(n589) );
  XNOR U491 ( .A(y[57]), .B(x[57]), .Z(n415) );
  NANDN U492 ( .A(x[56]), .B(y[56]), .Z(n414) );
  AND U493 ( .A(n415), .B(n414), .Z(n583) );
  AND U494 ( .A(n589), .B(n583), .Z(n421) );
  XNOR U495 ( .A(y[61]), .B(x[61]), .Z(n417) );
  NANDN U496 ( .A(x[60]), .B(y[60]), .Z(n416) );
  AND U497 ( .A(n417), .B(n416), .Z(n587) );
  XNOR U498 ( .A(y[59]), .B(x[59]), .Z(n419) );
  NANDN U499 ( .A(x[58]), .B(y[58]), .Z(n418) );
  AND U500 ( .A(n419), .B(n418), .Z(n585) );
  AND U501 ( .A(n587), .B(n585), .Z(n420) );
  AND U502 ( .A(n421), .B(n420), .Z(n433) );
  XNOR U503 ( .A(y[39]), .B(x[39]), .Z(n423) );
  NANDN U504 ( .A(x[38]), .B(y[38]), .Z(n422) );
  AND U505 ( .A(n423), .B(n422), .Z(n562) );
  XNOR U506 ( .A(y[33]), .B(x[33]), .Z(n425) );
  NANDN U507 ( .A(x[32]), .B(y[32]), .Z(n424) );
  AND U508 ( .A(n425), .B(n424), .Z(n555) );
  AND U509 ( .A(n562), .B(n555), .Z(n431) );
  XNOR U510 ( .A(y[37]), .B(x[37]), .Z(n427) );
  NANDN U511 ( .A(x[36]), .B(y[36]), .Z(n426) );
  AND U512 ( .A(n427), .B(n426), .Z(n559) );
  XNOR U513 ( .A(y[35]), .B(x[35]), .Z(n429) );
  NANDN U514 ( .A(x[34]), .B(y[34]), .Z(n428) );
  AND U515 ( .A(n429), .B(n428), .Z(n557) );
  AND U516 ( .A(n559), .B(n557), .Z(n430) );
  AND U517 ( .A(n431), .B(n430), .Z(n432) );
  AND U518 ( .A(n433), .B(n432), .Z(n434) );
  AND U519 ( .A(n435), .B(n434), .Z(n499) );
  NANDN U520 ( .A(y[126]), .B(x[126]), .Z(n649) );
  NANDN U521 ( .A(y[120]), .B(x[120]), .Z(n505) );
  AND U522 ( .A(n649), .B(n505), .Z(n437) );
  NANDN U523 ( .A(y[124]), .B(x[124]), .Z(n647) );
  NANDN U524 ( .A(y[122]), .B(x[122]), .Z(n504) );
  AND U525 ( .A(n647), .B(n504), .Z(n436) );
  AND U526 ( .A(n437), .B(n436), .Z(n441) );
  NANDN U527 ( .A(y[102]), .B(x[102]), .Z(n625) );
  NANDN U528 ( .A(y[96]), .B(x[96]), .Z(n511) );
  AND U529 ( .A(n625), .B(n511), .Z(n439) );
  NANDN U530 ( .A(y[100]), .B(x[100]), .Z(n623) );
  NANDN U531 ( .A(y[98]), .B(x[98]), .Z(n510) );
  AND U532 ( .A(n623), .B(n510), .Z(n438) );
  AND U533 ( .A(n439), .B(n438), .Z(n440) );
  AND U534 ( .A(n441), .B(n440), .Z(n449) );
  NANDN U535 ( .A(y[118]), .B(x[118]), .Z(n642) );
  NANDN U536 ( .A(y[112]), .B(x[112]), .Z(n507) );
  AND U537 ( .A(n642), .B(n507), .Z(n443) );
  NANDN U538 ( .A(y[116]), .B(x[116]), .Z(n640) );
  NANDN U539 ( .A(y[114]), .B(x[114]), .Z(n506) );
  AND U540 ( .A(n640), .B(n506), .Z(n442) );
  AND U541 ( .A(n443), .B(n442), .Z(n447) );
  NANDN U542 ( .A(y[110]), .B(x[110]), .Z(n633) );
  NANDN U543 ( .A(y[104]), .B(x[104]), .Z(n509) );
  AND U544 ( .A(n633), .B(n509), .Z(n445) );
  NANDN U545 ( .A(y[108]), .B(x[108]), .Z(n631) );
  NANDN U546 ( .A(y[106]), .B(x[106]), .Z(n508) );
  AND U547 ( .A(n631), .B(n508), .Z(n444) );
  AND U548 ( .A(n445), .B(n444), .Z(n446) );
  AND U549 ( .A(n447), .B(n446), .Z(n448) );
  AND U550 ( .A(n449), .B(n448), .Z(n465) );
  NANDN U551 ( .A(y[30]), .B(x[30]), .Z(n552) );
  NANDN U552 ( .A(y[24]), .B(x[24]), .Z(n545) );
  AND U553 ( .A(n552), .B(n545), .Z(n451) );
  NANDN U554 ( .A(y[28]), .B(x[28]), .Z(n549) );
  NANDN U555 ( .A(y[26]), .B(x[26]), .Z(n547) );
  AND U556 ( .A(n549), .B(n547), .Z(n450) );
  AND U557 ( .A(n451), .B(n450), .Z(n455) );
  NANDN U558 ( .A(y[6]), .B(x[6]), .Z(n525) );
  NANDN U559 ( .A(y[4]), .B(x[4]), .Z(n523) );
  AND U560 ( .A(n525), .B(n523), .Z(n453) );
  NANDN U561 ( .A(y[2]), .B(x[2]), .Z(n520) );
  NANDN U562 ( .A(y[0]), .B(x[0]), .Z(n519) );
  AND U563 ( .A(n520), .B(n519), .Z(n452) );
  AND U564 ( .A(n453), .B(n452), .Z(n454) );
  AND U565 ( .A(n455), .B(n454), .Z(n463) );
  NANDN U566 ( .A(y[22]), .B(x[22]), .Z(n543) );
  NANDN U567 ( .A(y[16]), .B(x[16]), .Z(n536) );
  AND U568 ( .A(n543), .B(n536), .Z(n457) );
  NANDN U569 ( .A(y[20]), .B(x[20]), .Z(n540) );
  NANDN U570 ( .A(y[18]), .B(x[18]), .Z(n538) );
  AND U571 ( .A(n540), .B(n538), .Z(n456) );
  AND U572 ( .A(n457), .B(n456), .Z(n461) );
  NANDN U573 ( .A(y[14]), .B(x[14]), .Z(n534) );
  NANDN U574 ( .A(y[8]), .B(x[8]), .Z(n527) );
  AND U575 ( .A(n534), .B(n527), .Z(n459) );
  NANDN U576 ( .A(y[12]), .B(x[12]), .Z(n532) );
  NANDN U577 ( .A(y[10]), .B(x[10]), .Z(n529) );
  AND U578 ( .A(n532), .B(n529), .Z(n458) );
  AND U579 ( .A(n459), .B(n458), .Z(n460) );
  AND U580 ( .A(n461), .B(n460), .Z(n462) );
  AND U581 ( .A(n463), .B(n462), .Z(n464) );
  AND U582 ( .A(n465), .B(n464), .Z(n497) );
  NANDN U583 ( .A(y[94]), .B(x[94]), .Z(n619) );
  NANDN U584 ( .A(y[88]), .B(x[88]), .Z(n513) );
  AND U585 ( .A(n619), .B(n513), .Z(n467) );
  NANDN U586 ( .A(y[92]), .B(x[92]), .Z(n616) );
  NANDN U587 ( .A(y[90]), .B(x[90]), .Z(n512) );
  AND U588 ( .A(n616), .B(n512), .Z(n466) );
  AND U589 ( .A(n467), .B(n466), .Z(n471) );
  NANDN U590 ( .A(y[70]), .B(x[70]), .Z(n596) );
  NANDN U591 ( .A(y[64]), .B(x[64]), .Z(n590) );
  AND U592 ( .A(n596), .B(n590), .Z(n469) );
  NANDN U593 ( .A(y[68]), .B(x[68]), .Z(n594) );
  NANDN U594 ( .A(y[66]), .B(x[66]), .Z(n518) );
  AND U595 ( .A(n594), .B(n518), .Z(n468) );
  AND U596 ( .A(n469), .B(n468), .Z(n470) );
  AND U597 ( .A(n471), .B(n470), .Z(n479) );
  NANDN U598 ( .A(y[86]), .B(x[86]), .Z(n612) );
  NANDN U599 ( .A(y[80]), .B(x[80]), .Z(n515) );
  AND U600 ( .A(n612), .B(n515), .Z(n473) );
  NANDN U601 ( .A(y[84]), .B(x[84]), .Z(n609) );
  NANDN U602 ( .A(y[82]), .B(x[82]), .Z(n514) );
  AND U603 ( .A(n609), .B(n514), .Z(n472) );
  AND U604 ( .A(n473), .B(n472), .Z(n477) );
  NANDN U605 ( .A(y[78]), .B(x[78]), .Z(n604) );
  NANDN U606 ( .A(y[72]), .B(x[72]), .Z(n517) );
  AND U607 ( .A(n604), .B(n517), .Z(n475) );
  NANDN U608 ( .A(y[76]), .B(x[76]), .Z(n602) );
  NANDN U609 ( .A(y[74]), .B(x[74]), .Z(n516) );
  AND U610 ( .A(n602), .B(n516), .Z(n474) );
  AND U611 ( .A(n475), .B(n474), .Z(n476) );
  AND U612 ( .A(n477), .B(n476), .Z(n478) );
  AND U613 ( .A(n479), .B(n478), .Z(n495) );
  NANDN U614 ( .A(y[62]), .B(x[62]), .Z(n588) );
  NANDN U615 ( .A(y[56]), .B(x[56]), .Z(n580) );
  AND U616 ( .A(n588), .B(n580), .Z(n481) );
  NANDN U617 ( .A(y[60]), .B(x[60]), .Z(n586) );
  NANDN U618 ( .A(y[58]), .B(x[58]), .Z(n584) );
  AND U619 ( .A(n586), .B(n584), .Z(n480) );
  AND U620 ( .A(n481), .B(n480), .Z(n485) );
  NANDN U621 ( .A(y[38]), .B(x[38]), .Z(n560) );
  NANDN U622 ( .A(y[32]), .B(x[32]), .Z(n554) );
  AND U623 ( .A(n560), .B(n554), .Z(n483) );
  NANDN U624 ( .A(y[36]), .B(x[36]), .Z(n558) );
  NANDN U625 ( .A(y[34]), .B(x[34]), .Z(n556) );
  AND U626 ( .A(n558), .B(n556), .Z(n482) );
  AND U627 ( .A(n483), .B(n482), .Z(n484) );
  AND U628 ( .A(n485), .B(n484), .Z(n493) );
  NANDN U629 ( .A(y[54]), .B(x[54]), .Z(n578) );
  NANDN U630 ( .A(y[48]), .B(x[48]), .Z(n572) );
  AND U631 ( .A(n578), .B(n572), .Z(n487) );
  NANDN U632 ( .A(y[52]), .B(x[52]), .Z(n576) );
  NANDN U633 ( .A(y[50]), .B(x[50]), .Z(n574) );
  AND U634 ( .A(n576), .B(n574), .Z(n486) );
  AND U635 ( .A(n487), .B(n486), .Z(n491) );
  NANDN U636 ( .A(y[46]), .B(x[46]), .Z(n569) );
  NANDN U637 ( .A(y[40]), .B(x[40]), .Z(n563) );
  AND U638 ( .A(n569), .B(n563), .Z(n489) );
  NANDN U639 ( .A(y[44]), .B(x[44]), .Z(n567) );
  NANDN U640 ( .A(y[42]), .B(x[42]), .Z(n565) );
  AND U641 ( .A(n567), .B(n565), .Z(n488) );
  AND U642 ( .A(n489), .B(n488), .Z(n490) );
  AND U643 ( .A(n491), .B(n490), .Z(n492) );
  AND U644 ( .A(n493), .B(n492), .Z(n494) );
  AND U645 ( .A(n495), .B(n494), .Z(n496) );
  AND U646 ( .A(n497), .B(n496), .Z(n498) );
  AND U647 ( .A(n499), .B(n498), .Z(n500) );
  AND U648 ( .A(n501), .B(n500), .Z(n502) );
  NAND U649 ( .A(n503), .B(n502), .Z(n651) );
  NANDN U650 ( .A(n651), .B(e), .Z(n5) );
  IV U651 ( .A(n507), .Z(n636) );
  IV U652 ( .A(n580), .Z(n581) );
  ANDN U653 ( .B(x[73]), .A(y[73]), .Z(n599) );
  ANDN U654 ( .B(x[83]), .A(y[83]), .Z(n610) );
  ANDN U655 ( .B(x[101]), .A(y[101]), .Z(n626) );
  ANDN U656 ( .B(x[111]), .A(y[111]), .Z(n637) );
endmodule

