
module sum_N262144_CC512 ( clk, rst, a, b, c );
  input [511:0] a;
  input [511:0] b;
  output [511:0] c;
  input clk, rst;
  wire   carry_on, carry_on_d, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048;

  DFF carry_on_reg ( .D(carry_on_d), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        carry_on) );
  XOR U4 ( .A(a[1]), .B(n2044), .Z(n1342) );
  XOR U5 ( .A(a[4]), .B(n2035), .Z(n109) );
  XOR U6 ( .A(a[7]), .B(n2026), .Z(n28) );
  XOR U7 ( .A(a[10]), .B(n2017), .Z(n1712) );
  XOR U8 ( .A(a[13]), .B(n2008), .Z(n1589) );
  XOR U9 ( .A(a[16]), .B(n1999), .Z(n1466) );
  XOR U10 ( .A(a[19]), .B(n1990), .Z(n1343) );
  XOR U11 ( .A(a[22]), .B(n1981), .Z(n1219) );
  XOR U12 ( .A(a[25]), .B(n1972), .Z(n1096) );
  XOR U13 ( .A(a[28]), .B(n1963), .Z(n973) );
  XOR U14 ( .A(a[31]), .B(n1954), .Z(n849) );
  XOR U15 ( .A(a[34]), .B(n1945), .Z(n726) );
  XOR U16 ( .A(a[37]), .B(n1936), .Z(n603) );
  XOR U17 ( .A(a[40]), .B(n1927), .Z(n479) );
  XOR U18 ( .A(a[43]), .B(n1918), .Z(n356) );
  XOR U19 ( .A(a[46]), .B(n1909), .Z(n233) );
  XOR U20 ( .A(a[49]), .B(n1900), .Z(n110) );
  XOR U21 ( .A(a[52]), .B(n1891), .Z(n58) );
  XOR U22 ( .A(a[55]), .B(n1882), .Z(n55) );
  XOR U23 ( .A(a[58]), .B(n1873), .Z(n52) );
  XOR U24 ( .A(a[61]), .B(n1864), .Z(n48) );
  XOR U25 ( .A(a[64]), .B(n1855), .Z(n45) );
  XOR U26 ( .A(a[67]), .B(n1846), .Z(n42) );
  XOR U27 ( .A(a[70]), .B(n1837), .Z(n38) );
  XOR U28 ( .A(a[73]), .B(n1828), .Z(n35) );
  XOR U29 ( .A(a[76]), .B(n1819), .Z(n32) );
  XOR U30 ( .A(a[79]), .B(n1810), .Z(n29) );
  XOR U31 ( .A(a[82]), .B(n1801), .Z(n25) );
  XOR U32 ( .A(a[85]), .B(n1792), .Z(n22) );
  XOR U33 ( .A(a[88]), .B(n1783), .Z(n19) );
  XOR U34 ( .A(a[91]), .B(n1774), .Z(n15) );
  XOR U35 ( .A(a[94]), .B(n1765), .Z(n12) );
  XOR U36 ( .A(a[97]), .B(n1756), .Z(n9) );
  XOR U37 ( .A(a[100]), .B(n1746), .Z(n1748) );
  XOR U38 ( .A(a[103]), .B(n1734), .Z(n1736) );
  XOR U39 ( .A(a[106]), .B(n1722), .Z(n1724) );
  XOR U40 ( .A(a[109]), .B(n1709), .Z(n1711) );
  XOR U41 ( .A(a[112]), .B(n1697), .Z(n1699) );
  XOR U42 ( .A(a[115]), .B(n1685), .Z(n1687) );
  XOR U43 ( .A(a[118]), .B(n1673), .Z(n1675) );
  XOR U44 ( .A(a[121]), .B(n1660), .Z(n1662) );
  XOR U45 ( .A(a[124]), .B(n1648), .Z(n1650) );
  XOR U46 ( .A(a[127]), .B(n1636), .Z(n1638) );
  XOR U47 ( .A(a[130]), .B(n1623), .Z(n1625) );
  XOR U48 ( .A(a[133]), .B(n1611), .Z(n1613) );
  XOR U49 ( .A(a[136]), .B(n1599), .Z(n1601) );
  XOR U50 ( .A(a[139]), .B(n1586), .Z(n1588) );
  XOR U51 ( .A(a[142]), .B(n1574), .Z(n1576) );
  XOR U52 ( .A(a[145]), .B(n1562), .Z(n1564) );
  XOR U53 ( .A(a[148]), .B(n1550), .Z(n1552) );
  XOR U54 ( .A(a[151]), .B(n1537), .Z(n1539) );
  XOR U55 ( .A(a[154]), .B(n1525), .Z(n1527) );
  XOR U56 ( .A(a[157]), .B(n1513), .Z(n1515) );
  XOR U57 ( .A(a[160]), .B(n1500), .Z(n1502) );
  XOR U58 ( .A(a[163]), .B(n1488), .Z(n1490) );
  XOR U59 ( .A(a[166]), .B(n1476), .Z(n1478) );
  XOR U60 ( .A(a[169]), .B(n1463), .Z(n1465) );
  XOR U61 ( .A(a[172]), .B(n1451), .Z(n1453) );
  XOR U62 ( .A(a[175]), .B(n1439), .Z(n1441) );
  XOR U63 ( .A(a[178]), .B(n1427), .Z(n1429) );
  XOR U64 ( .A(a[181]), .B(n1414), .Z(n1416) );
  XOR U65 ( .A(a[184]), .B(n1402), .Z(n1404) );
  XOR U66 ( .A(a[187]), .B(n1390), .Z(n1392) );
  XOR U67 ( .A(a[190]), .B(n1377), .Z(n1379) );
  XOR U68 ( .A(a[193]), .B(n1365), .Z(n1367) );
  XOR U69 ( .A(a[196]), .B(n1353), .Z(n1355) );
  XOR U70 ( .A(a[199]), .B(n1339), .Z(n1341) );
  XOR U71 ( .A(a[202]), .B(n1327), .Z(n1329) );
  XOR U72 ( .A(a[205]), .B(n1315), .Z(n1317) );
  XOR U73 ( .A(a[208]), .B(n1303), .Z(n1305) );
  XOR U74 ( .A(a[211]), .B(n1290), .Z(n1292) );
  XOR U75 ( .A(a[214]), .B(n1278), .Z(n1280) );
  XOR U76 ( .A(a[217]), .B(n1266), .Z(n1268) );
  XOR U77 ( .A(a[220]), .B(n1253), .Z(n1255) );
  XOR U78 ( .A(a[223]), .B(n1241), .Z(n1243) );
  XOR U79 ( .A(a[226]), .B(n1229), .Z(n1231) );
  XOR U80 ( .A(a[229]), .B(n1216), .Z(n1218) );
  XOR U81 ( .A(a[232]), .B(n1204), .Z(n1206) );
  XOR U82 ( .A(a[235]), .B(n1192), .Z(n1194) );
  XOR U83 ( .A(a[238]), .B(n1180), .Z(n1182) );
  XOR U84 ( .A(a[241]), .B(n1167), .Z(n1169) );
  XOR U85 ( .A(a[244]), .B(n1155), .Z(n1157) );
  XOR U86 ( .A(a[247]), .B(n1143), .Z(n1145) );
  XOR U87 ( .A(a[250]), .B(n1130), .Z(n1132) );
  XOR U88 ( .A(a[253]), .B(n1118), .Z(n1120) );
  XOR U89 ( .A(a[256]), .B(n1106), .Z(n1108) );
  XOR U90 ( .A(a[259]), .B(n1093), .Z(n1095) );
  XOR U91 ( .A(a[262]), .B(n1081), .Z(n1083) );
  XOR U92 ( .A(a[265]), .B(n1069), .Z(n1071) );
  XOR U93 ( .A(a[268]), .B(n1057), .Z(n1059) );
  XOR U94 ( .A(a[271]), .B(n1044), .Z(n1046) );
  XOR U95 ( .A(a[274]), .B(n1032), .Z(n1034) );
  XOR U96 ( .A(a[277]), .B(n1020), .Z(n1022) );
  XOR U97 ( .A(a[280]), .B(n1007), .Z(n1009) );
  XOR U98 ( .A(a[283]), .B(n995), .Z(n997) );
  XOR U99 ( .A(a[286]), .B(n983), .Z(n985) );
  XOR U100 ( .A(a[289]), .B(n970), .Z(n972) );
  XOR U101 ( .A(a[292]), .B(n958), .Z(n960) );
  XOR U102 ( .A(a[295]), .B(n946), .Z(n948) );
  XOR U103 ( .A(a[298]), .B(n934), .Z(n936) );
  XOR U104 ( .A(a[301]), .B(n920), .Z(n922) );
  XOR U105 ( .A(a[304]), .B(n908), .Z(n910) );
  XOR U106 ( .A(a[307]), .B(n896), .Z(n898) );
  XOR U107 ( .A(a[310]), .B(n883), .Z(n885) );
  XOR U108 ( .A(a[313]), .B(n871), .Z(n873) );
  XOR U109 ( .A(a[316]), .B(n859), .Z(n861) );
  XOR U110 ( .A(a[319]), .B(n846), .Z(n848) );
  XOR U111 ( .A(a[322]), .B(n834), .Z(n836) );
  XOR U112 ( .A(a[325]), .B(n822), .Z(n824) );
  XOR U113 ( .A(a[328]), .B(n810), .Z(n812) );
  XOR U114 ( .A(a[331]), .B(n797), .Z(n799) );
  XOR U115 ( .A(a[334]), .B(n785), .Z(n787) );
  XOR U116 ( .A(a[337]), .B(n773), .Z(n775) );
  XOR U117 ( .A(a[340]), .B(n760), .Z(n762) );
  XOR U118 ( .A(a[343]), .B(n748), .Z(n750) );
  XOR U119 ( .A(a[346]), .B(n736), .Z(n738) );
  XOR U120 ( .A(a[349]), .B(n723), .Z(n725) );
  XOR U121 ( .A(a[352]), .B(n711), .Z(n713) );
  XOR U122 ( .A(a[355]), .B(n699), .Z(n701) );
  XOR U123 ( .A(a[358]), .B(n687), .Z(n689) );
  XOR U124 ( .A(a[361]), .B(n674), .Z(n676) );
  XOR U125 ( .A(a[364]), .B(n662), .Z(n664) );
  XOR U126 ( .A(a[367]), .B(n650), .Z(n652) );
  XOR U127 ( .A(a[370]), .B(n637), .Z(n639) );
  XOR U128 ( .A(a[373]), .B(n625), .Z(n627) );
  XOR U129 ( .A(a[376]), .B(n613), .Z(n615) );
  XOR U130 ( .A(a[379]), .B(n600), .Z(n602) );
  XOR U131 ( .A(a[382]), .B(n588), .Z(n590) );
  XOR U132 ( .A(a[385]), .B(n576), .Z(n578) );
  XOR U133 ( .A(a[388]), .B(n564), .Z(n566) );
  XOR U134 ( .A(a[391]), .B(n551), .Z(n553) );
  XOR U135 ( .A(a[394]), .B(n539), .Z(n541) );
  XOR U136 ( .A(a[397]), .B(n527), .Z(n529) );
  XOR U137 ( .A(a[400]), .B(n513), .Z(n515) );
  XOR U138 ( .A(a[403]), .B(n501), .Z(n503) );
  XOR U139 ( .A(a[406]), .B(n489), .Z(n491) );
  XOR U140 ( .A(a[409]), .B(n476), .Z(n478) );
  XOR U141 ( .A(a[412]), .B(n464), .Z(n466) );
  XOR U142 ( .A(a[415]), .B(n452), .Z(n454) );
  XOR U143 ( .A(a[418]), .B(n440), .Z(n442) );
  XOR U144 ( .A(a[421]), .B(n427), .Z(n429) );
  XOR U145 ( .A(a[424]), .B(n415), .Z(n417) );
  XOR U146 ( .A(a[427]), .B(n403), .Z(n405) );
  XOR U147 ( .A(a[430]), .B(n390), .Z(n392) );
  XOR U148 ( .A(a[433]), .B(n378), .Z(n380) );
  XOR U149 ( .A(a[436]), .B(n366), .Z(n368) );
  XOR U150 ( .A(a[439]), .B(n353), .Z(n355) );
  XOR U151 ( .A(a[442]), .B(n341), .Z(n343) );
  XOR U152 ( .A(a[445]), .B(n329), .Z(n331) );
  XOR U153 ( .A(a[448]), .B(n317), .Z(n319) );
  XOR U154 ( .A(a[451]), .B(n304), .Z(n306) );
  XOR U155 ( .A(a[454]), .B(n292), .Z(n294) );
  XOR U156 ( .A(a[457]), .B(n280), .Z(n282) );
  XOR U157 ( .A(a[460]), .B(n267), .Z(n269) );
  XOR U158 ( .A(a[463]), .B(n255), .Z(n257) );
  XOR U159 ( .A(a[466]), .B(n243), .Z(n245) );
  XOR U160 ( .A(a[469]), .B(n230), .Z(n232) );
  XOR U161 ( .A(a[472]), .B(n218), .Z(n220) );
  XOR U162 ( .A(a[475]), .B(n206), .Z(n208) );
  XOR U163 ( .A(a[478]), .B(n194), .Z(n196) );
  XOR U164 ( .A(a[481]), .B(n181), .Z(n183) );
  XOR U165 ( .A(a[484]), .B(n169), .Z(n171) );
  XOR U166 ( .A(a[487]), .B(n157), .Z(n159) );
  XOR U167 ( .A(a[490]), .B(n144), .Z(n146) );
  XOR U168 ( .A(a[493]), .B(n132), .Z(n134) );
  XOR U169 ( .A(a[496]), .B(n120), .Z(n122) );
  XOR U170 ( .A(a[499]), .B(n106), .Z(n108) );
  XOR U171 ( .A(a[502]), .B(n94), .Z(n96) );
  XOR U172 ( .A(a[505]), .B(n82), .Z(n84) );
  XOR U173 ( .A(a[508]), .B(n70), .Z(n72) );
  XOR U174 ( .A(a[2]), .B(n2041), .Z(n931) );
  XOR U175 ( .A(a[5]), .B(n2032), .Z(n50) );
  XOR U176 ( .A(a[8]), .B(n2023), .Z(n17) );
  XOR U177 ( .A(a[11]), .B(n2014), .Z(n1671) );
  XOR U178 ( .A(a[14]), .B(n2005), .Z(n1548) );
  XOR U179 ( .A(a[17]), .B(n1996), .Z(n1425) );
  XOR U180 ( .A(a[20]), .B(n1987), .Z(n1301) );
  XOR U181 ( .A(a[23]), .B(n1978), .Z(n1178) );
  XOR U182 ( .A(a[26]), .B(n1969), .Z(n1055) );
  XOR U183 ( .A(a[29]), .B(n1960), .Z(n932) );
  XOR U184 ( .A(a[32]), .B(n1951), .Z(n808) );
  XOR U185 ( .A(a[35]), .B(n1942), .Z(n685) );
  XOR U186 ( .A(a[38]), .B(n1933), .Z(n562) );
  XOR U187 ( .A(a[41]), .B(n1924), .Z(n438) );
  XOR U188 ( .A(a[44]), .B(n1915), .Z(n315) );
  XOR U189 ( .A(a[47]), .B(n1906), .Z(n192) );
  XOR U190 ( .A(a[50]), .B(n1897), .Z(n68) );
  XOR U191 ( .A(a[53]), .B(n1888), .Z(n57) );
  XOR U192 ( .A(a[56]), .B(n1879), .Z(n54) );
  XOR U193 ( .A(a[59]), .B(n1870), .Z(n51) );
  XOR U194 ( .A(a[62]), .B(n1861), .Z(n47) );
  XOR U195 ( .A(a[65]), .B(n1852), .Z(n44) );
  XOR U196 ( .A(a[68]), .B(n1843), .Z(n41) );
  XOR U197 ( .A(a[71]), .B(n1834), .Z(n37) );
  XOR U198 ( .A(a[74]), .B(n1825), .Z(n34) );
  XOR U199 ( .A(a[77]), .B(n1816), .Z(n31) );
  XOR U200 ( .A(a[80]), .B(n1807), .Z(n27) );
  XOR U201 ( .A(a[83]), .B(n1798), .Z(n24) );
  XOR U202 ( .A(a[86]), .B(n1789), .Z(n21) );
  XOR U203 ( .A(a[89]), .B(n1780), .Z(n18) );
  XOR U204 ( .A(a[92]), .B(n1771), .Z(n14) );
  XOR U205 ( .A(a[95]), .B(n1762), .Z(n11) );
  XOR U206 ( .A(a[98]), .B(n1753), .Z(n8) );
  XOR U207 ( .A(a[101]), .B(n1742), .Z(n1744) );
  XOR U208 ( .A(a[104]), .B(n1730), .Z(n1732) );
  XOR U209 ( .A(a[107]), .B(n1718), .Z(n1720) );
  XOR U210 ( .A(a[110]), .B(n1705), .Z(n1707) );
  XOR U211 ( .A(a[113]), .B(n1693), .Z(n1695) );
  XOR U212 ( .A(a[116]), .B(n1681), .Z(n1683) );
  XOR U213 ( .A(a[119]), .B(n1668), .Z(n1670) );
  XOR U214 ( .A(a[122]), .B(n1656), .Z(n1658) );
  XOR U215 ( .A(a[125]), .B(n1644), .Z(n1646) );
  XOR U216 ( .A(a[128]), .B(n1632), .Z(n1634) );
  XOR U217 ( .A(a[131]), .B(n1619), .Z(n1621) );
  XOR U218 ( .A(a[134]), .B(n1607), .Z(n1609) );
  XOR U219 ( .A(a[137]), .B(n1595), .Z(n1597) );
  XOR U220 ( .A(a[140]), .B(n1582), .Z(n1584) );
  XOR U221 ( .A(a[143]), .B(n1570), .Z(n1572) );
  XOR U222 ( .A(a[146]), .B(n1558), .Z(n1560) );
  XOR U223 ( .A(a[149]), .B(n1545), .Z(n1547) );
  XOR U224 ( .A(a[152]), .B(n1533), .Z(n1535) );
  XOR U225 ( .A(a[155]), .B(n1521), .Z(n1523) );
  XOR U226 ( .A(a[158]), .B(n1509), .Z(n1511) );
  XOR U227 ( .A(a[161]), .B(n1496), .Z(n1498) );
  XOR U228 ( .A(a[164]), .B(n1484), .Z(n1486) );
  XOR U229 ( .A(a[167]), .B(n1472), .Z(n1474) );
  XOR U230 ( .A(a[170]), .B(n1459), .Z(n1461) );
  XOR U231 ( .A(a[173]), .B(n1447), .Z(n1449) );
  XOR U232 ( .A(a[176]), .B(n1435), .Z(n1437) );
  XOR U233 ( .A(a[179]), .B(n1422), .Z(n1424) );
  XOR U234 ( .A(a[182]), .B(n1410), .Z(n1412) );
  XOR U235 ( .A(a[185]), .B(n1398), .Z(n1400) );
  XOR U236 ( .A(a[188]), .B(n1386), .Z(n1388) );
  XOR U237 ( .A(a[191]), .B(n1373), .Z(n1375) );
  XOR U238 ( .A(a[194]), .B(n1361), .Z(n1363) );
  XOR U239 ( .A(a[197]), .B(n1349), .Z(n1351) );
  XOR U240 ( .A(a[200]), .B(n1335), .Z(n1337) );
  XOR U241 ( .A(a[203]), .B(n1323), .Z(n1325) );
  XOR U242 ( .A(a[206]), .B(n1311), .Z(n1313) );
  XOR U243 ( .A(a[209]), .B(n1298), .Z(n1300) );
  XOR U244 ( .A(a[212]), .B(n1286), .Z(n1288) );
  XOR U245 ( .A(a[215]), .B(n1274), .Z(n1276) );
  XOR U246 ( .A(a[218]), .B(n1262), .Z(n1264) );
  XOR U247 ( .A(a[221]), .B(n1249), .Z(n1251) );
  XOR U248 ( .A(a[224]), .B(n1237), .Z(n1239) );
  XOR U249 ( .A(a[227]), .B(n1225), .Z(n1227) );
  XOR U250 ( .A(a[230]), .B(n1212), .Z(n1214) );
  XOR U251 ( .A(a[233]), .B(n1200), .Z(n1202) );
  XOR U252 ( .A(a[236]), .B(n1188), .Z(n1190) );
  XOR U253 ( .A(a[239]), .B(n1175), .Z(n1177) );
  XOR U254 ( .A(a[242]), .B(n1163), .Z(n1165) );
  XOR U255 ( .A(a[245]), .B(n1151), .Z(n1153) );
  XOR U256 ( .A(a[248]), .B(n1139), .Z(n1141) );
  XOR U257 ( .A(a[251]), .B(n1126), .Z(n1128) );
  XOR U258 ( .A(a[254]), .B(n1114), .Z(n1116) );
  XOR U259 ( .A(a[257]), .B(n1102), .Z(n1104) );
  XOR U260 ( .A(a[260]), .B(n1089), .Z(n1091) );
  XOR U261 ( .A(a[263]), .B(n1077), .Z(n1079) );
  XOR U262 ( .A(a[266]), .B(n1065), .Z(n1067) );
  XOR U263 ( .A(a[269]), .B(n1052), .Z(n1054) );
  XOR U264 ( .A(a[272]), .B(n1040), .Z(n1042) );
  XOR U265 ( .A(a[275]), .B(n1028), .Z(n1030) );
  XOR U266 ( .A(a[278]), .B(n1016), .Z(n1018) );
  XOR U267 ( .A(a[281]), .B(n1003), .Z(n1005) );
  XOR U268 ( .A(a[284]), .B(n991), .Z(n993) );
  XOR U269 ( .A(a[287]), .B(n979), .Z(n981) );
  XOR U270 ( .A(a[290]), .B(n966), .Z(n968) );
  XOR U271 ( .A(a[293]), .B(n954), .Z(n956) );
  XOR U272 ( .A(a[296]), .B(n942), .Z(n944) );
  XOR U273 ( .A(a[299]), .B(n928), .Z(n930) );
  XOR U274 ( .A(a[302]), .B(n916), .Z(n918) );
  XOR U275 ( .A(a[305]), .B(n904), .Z(n906) );
  XOR U276 ( .A(a[308]), .B(n892), .Z(n894) );
  XOR U277 ( .A(a[311]), .B(n879), .Z(n881) );
  XOR U278 ( .A(a[314]), .B(n867), .Z(n869) );
  XOR U279 ( .A(a[317]), .B(n855), .Z(n857) );
  XOR U280 ( .A(a[320]), .B(n842), .Z(n844) );
  XOR U281 ( .A(a[323]), .B(n830), .Z(n832) );
  XOR U282 ( .A(a[326]), .B(n818), .Z(n820) );
  XOR U283 ( .A(a[329]), .B(n805), .Z(n807) );
  XOR U284 ( .A(a[332]), .B(n793), .Z(n795) );
  XOR U285 ( .A(a[335]), .B(n781), .Z(n783) );
  XOR U286 ( .A(a[338]), .B(n769), .Z(n771) );
  XOR U287 ( .A(a[341]), .B(n756), .Z(n758) );
  XOR U288 ( .A(a[344]), .B(n744), .Z(n746) );
  XOR U289 ( .A(a[347]), .B(n732), .Z(n734) );
  XOR U290 ( .A(a[350]), .B(n719), .Z(n721) );
  XOR U291 ( .A(a[353]), .B(n707), .Z(n709) );
  XOR U292 ( .A(a[356]), .B(n695), .Z(n697) );
  XOR U293 ( .A(a[359]), .B(n682), .Z(n684) );
  XOR U294 ( .A(a[362]), .B(n670), .Z(n672) );
  XOR U295 ( .A(a[365]), .B(n658), .Z(n660) );
  XOR U296 ( .A(a[368]), .B(n646), .Z(n648) );
  XOR U297 ( .A(a[371]), .B(n633), .Z(n635) );
  XOR U298 ( .A(a[374]), .B(n621), .Z(n623) );
  XOR U299 ( .A(a[377]), .B(n609), .Z(n611) );
  XOR U300 ( .A(a[380]), .B(n596), .Z(n598) );
  XOR U301 ( .A(a[383]), .B(n584), .Z(n586) );
  XOR U302 ( .A(a[386]), .B(n572), .Z(n574) );
  XOR U303 ( .A(a[389]), .B(n559), .Z(n561) );
  XOR U304 ( .A(a[392]), .B(n547), .Z(n549) );
  XOR U305 ( .A(a[395]), .B(n535), .Z(n537) );
  XOR U306 ( .A(a[398]), .B(n523), .Z(n525) );
  XOR U307 ( .A(a[401]), .B(n509), .Z(n511) );
  XOR U308 ( .A(a[404]), .B(n497), .Z(n499) );
  XOR U309 ( .A(a[407]), .B(n485), .Z(n487) );
  XOR U310 ( .A(a[410]), .B(n472), .Z(n474) );
  XOR U311 ( .A(a[413]), .B(n460), .Z(n462) );
  XOR U312 ( .A(a[416]), .B(n448), .Z(n450) );
  XOR U313 ( .A(a[419]), .B(n435), .Z(n437) );
  XOR U314 ( .A(a[422]), .B(n423), .Z(n425) );
  XOR U315 ( .A(a[425]), .B(n411), .Z(n413) );
  XOR U316 ( .A(a[428]), .B(n399), .Z(n401) );
  XOR U317 ( .A(a[431]), .B(n386), .Z(n388) );
  XOR U318 ( .A(a[434]), .B(n374), .Z(n376) );
  XOR U319 ( .A(a[437]), .B(n362), .Z(n364) );
  XOR U320 ( .A(a[440]), .B(n349), .Z(n351) );
  XOR U321 ( .A(a[443]), .B(n337), .Z(n339) );
  XOR U322 ( .A(a[446]), .B(n325), .Z(n327) );
  XOR U323 ( .A(a[449]), .B(n312), .Z(n314) );
  XOR U324 ( .A(a[452]), .B(n300), .Z(n302) );
  XOR U325 ( .A(a[455]), .B(n288), .Z(n290) );
  XOR U326 ( .A(a[458]), .B(n276), .Z(n278) );
  XOR U327 ( .A(a[461]), .B(n263), .Z(n265) );
  XOR U328 ( .A(a[464]), .B(n251), .Z(n253) );
  XOR U329 ( .A(a[467]), .B(n239), .Z(n241) );
  XOR U330 ( .A(a[470]), .B(n226), .Z(n228) );
  XOR U331 ( .A(a[473]), .B(n214), .Z(n216) );
  XOR U332 ( .A(a[476]), .B(n202), .Z(n204) );
  XOR U333 ( .A(a[479]), .B(n189), .Z(n191) );
  XOR U334 ( .A(a[482]), .B(n177), .Z(n179) );
  XOR U335 ( .A(a[485]), .B(n165), .Z(n167) );
  XOR U336 ( .A(a[488]), .B(n153), .Z(n155) );
  XOR U337 ( .A(a[491]), .B(n140), .Z(n142) );
  XOR U338 ( .A(a[494]), .B(n128), .Z(n130) );
  XOR U339 ( .A(a[497]), .B(n116), .Z(n118) );
  XOR U340 ( .A(a[500]), .B(n102), .Z(n104) );
  XOR U341 ( .A(a[503]), .B(n90), .Z(n92) );
  XOR U342 ( .A(a[506]), .B(n78), .Z(n80) );
  XOR U343 ( .A(a[509]), .B(n65), .Z(n67) );
  XOR U344 ( .A(a[3]), .B(n2038), .Z(n520) );
  XOR U345 ( .A(a[6]), .B(n2029), .Z(n39) );
  XOR U346 ( .A(a[9]), .B(n2020), .Z(n6) );
  XOR U347 ( .A(a[12]), .B(n2011), .Z(n1630) );
  XOR U348 ( .A(a[15]), .B(n2002), .Z(n1507) );
  XOR U349 ( .A(a[18]), .B(n1993), .Z(n1384) );
  XOR U350 ( .A(a[21]), .B(n1984), .Z(n1260) );
  XOR U351 ( .A(a[24]), .B(n1975), .Z(n1137) );
  XOR U352 ( .A(a[27]), .B(n1966), .Z(n1014) );
  XOR U353 ( .A(a[30]), .B(n1957), .Z(n890) );
  XOR U354 ( .A(a[33]), .B(n1948), .Z(n767) );
  XOR U355 ( .A(a[36]), .B(n1939), .Z(n644) );
  XOR U356 ( .A(a[39]), .B(n1930), .Z(n521) );
  XOR U357 ( .A(a[42]), .B(n1921), .Z(n397) );
  XOR U358 ( .A(a[45]), .B(n1912), .Z(n274) );
  XOR U359 ( .A(a[48]), .B(n1903), .Z(n151) );
  XOR U360 ( .A(a[51]), .B(n1894), .Z(n59) );
  XOR U361 ( .A(a[54]), .B(n1885), .Z(n56) );
  XOR U362 ( .A(a[57]), .B(n1876), .Z(n53) );
  XOR U363 ( .A(a[60]), .B(n1867), .Z(n49) );
  XOR U364 ( .A(a[63]), .B(n1858), .Z(n46) );
  XOR U365 ( .A(a[66]), .B(n1849), .Z(n43) );
  XOR U366 ( .A(a[69]), .B(n1840), .Z(n40) );
  XOR U367 ( .A(a[72]), .B(n1831), .Z(n36) );
  XOR U368 ( .A(a[75]), .B(n1822), .Z(n33) );
  XOR U369 ( .A(a[78]), .B(n1813), .Z(n30) );
  XOR U370 ( .A(a[81]), .B(n1804), .Z(n26) );
  XOR U371 ( .A(a[84]), .B(n1795), .Z(n23) );
  XOR U372 ( .A(a[87]), .B(n1786), .Z(n20) );
  XOR U373 ( .A(a[90]), .B(n1777), .Z(n16) );
  XOR U374 ( .A(a[93]), .B(n1768), .Z(n13) );
  XOR U375 ( .A(a[96]), .B(n1759), .Z(n10) );
  XOR U376 ( .A(a[99]), .B(n1750), .Z(n7) );
  XOR U377 ( .A(a[102]), .B(n1738), .Z(n1740) );
  XOR U378 ( .A(a[105]), .B(n1726), .Z(n1728) );
  XOR U379 ( .A(a[108]), .B(n1714), .Z(n1716) );
  XOR U380 ( .A(a[111]), .B(n1701), .Z(n1703) );
  XOR U381 ( .A(a[114]), .B(n1689), .Z(n1691) );
  XOR U382 ( .A(a[117]), .B(n1677), .Z(n1679) );
  XOR U383 ( .A(a[120]), .B(n1664), .Z(n1666) );
  XOR U384 ( .A(a[123]), .B(n1652), .Z(n1654) );
  XOR U385 ( .A(a[126]), .B(n1640), .Z(n1642) );
  XOR U386 ( .A(a[129]), .B(n1627), .Z(n1629) );
  XOR U387 ( .A(a[132]), .B(n1615), .Z(n1617) );
  XOR U388 ( .A(a[135]), .B(n1603), .Z(n1605) );
  XOR U389 ( .A(a[138]), .B(n1591), .Z(n1593) );
  XOR U390 ( .A(a[141]), .B(n1578), .Z(n1580) );
  XOR U391 ( .A(a[144]), .B(n1566), .Z(n1568) );
  XOR U392 ( .A(a[147]), .B(n1554), .Z(n1556) );
  XOR U393 ( .A(a[150]), .B(n1541), .Z(n1543) );
  XOR U394 ( .A(a[153]), .B(n1529), .Z(n1531) );
  XOR U395 ( .A(a[156]), .B(n1517), .Z(n1519) );
  XOR U396 ( .A(a[159]), .B(n1504), .Z(n1506) );
  XOR U397 ( .A(a[162]), .B(n1492), .Z(n1494) );
  XOR U398 ( .A(a[165]), .B(n1480), .Z(n1482) );
  XOR U399 ( .A(a[168]), .B(n1468), .Z(n1470) );
  XOR U400 ( .A(a[171]), .B(n1455), .Z(n1457) );
  XOR U401 ( .A(a[174]), .B(n1443), .Z(n1445) );
  XOR U402 ( .A(a[177]), .B(n1431), .Z(n1433) );
  XOR U403 ( .A(a[180]), .B(n1418), .Z(n1420) );
  XOR U404 ( .A(a[183]), .B(n1406), .Z(n1408) );
  XOR U405 ( .A(a[186]), .B(n1394), .Z(n1396) );
  XOR U406 ( .A(a[189]), .B(n1381), .Z(n1383) );
  XOR U407 ( .A(a[192]), .B(n1369), .Z(n1371) );
  XOR U408 ( .A(a[195]), .B(n1357), .Z(n1359) );
  XOR U409 ( .A(a[198]), .B(n1345), .Z(n1347) );
  XOR U410 ( .A(a[201]), .B(n1331), .Z(n1333) );
  XOR U411 ( .A(a[204]), .B(n1319), .Z(n1321) );
  XOR U412 ( .A(a[207]), .B(n1307), .Z(n1309) );
  XOR U413 ( .A(a[210]), .B(n1294), .Z(n1296) );
  XOR U414 ( .A(a[213]), .B(n1282), .Z(n1284) );
  XOR U415 ( .A(a[216]), .B(n1270), .Z(n1272) );
  XOR U416 ( .A(a[219]), .B(n1257), .Z(n1259) );
  XOR U417 ( .A(a[222]), .B(n1245), .Z(n1247) );
  XOR U418 ( .A(a[225]), .B(n1233), .Z(n1235) );
  XOR U419 ( .A(a[228]), .B(n1221), .Z(n1223) );
  XOR U420 ( .A(a[231]), .B(n1208), .Z(n1210) );
  XOR U421 ( .A(a[234]), .B(n1196), .Z(n1198) );
  XOR U422 ( .A(a[237]), .B(n1184), .Z(n1186) );
  XOR U423 ( .A(a[240]), .B(n1171), .Z(n1173) );
  XOR U424 ( .A(a[243]), .B(n1159), .Z(n1161) );
  XOR U425 ( .A(a[246]), .B(n1147), .Z(n1149) );
  XOR U426 ( .A(a[249]), .B(n1134), .Z(n1136) );
  XOR U427 ( .A(a[252]), .B(n1122), .Z(n1124) );
  XOR U428 ( .A(a[255]), .B(n1110), .Z(n1112) );
  XOR U429 ( .A(a[258]), .B(n1098), .Z(n1100) );
  XOR U430 ( .A(a[261]), .B(n1085), .Z(n1087) );
  XOR U431 ( .A(a[264]), .B(n1073), .Z(n1075) );
  XOR U432 ( .A(a[267]), .B(n1061), .Z(n1063) );
  XOR U433 ( .A(a[270]), .B(n1048), .Z(n1050) );
  XOR U434 ( .A(a[273]), .B(n1036), .Z(n1038) );
  XOR U435 ( .A(a[276]), .B(n1024), .Z(n1026) );
  XOR U436 ( .A(a[279]), .B(n1011), .Z(n1013) );
  XOR U437 ( .A(a[282]), .B(n999), .Z(n1001) );
  XOR U438 ( .A(a[285]), .B(n987), .Z(n989) );
  XOR U439 ( .A(a[288]), .B(n975), .Z(n977) );
  XOR U440 ( .A(a[291]), .B(n962), .Z(n964) );
  XOR U441 ( .A(a[294]), .B(n950), .Z(n952) );
  XOR U442 ( .A(a[297]), .B(n938), .Z(n940) );
  XOR U443 ( .A(a[300]), .B(n924), .Z(n926) );
  XOR U444 ( .A(a[303]), .B(n912), .Z(n914) );
  XOR U445 ( .A(a[306]), .B(n900), .Z(n902) );
  XOR U446 ( .A(a[309]), .B(n887), .Z(n889) );
  XOR U447 ( .A(a[312]), .B(n875), .Z(n877) );
  XOR U448 ( .A(a[315]), .B(n863), .Z(n865) );
  XOR U449 ( .A(a[318]), .B(n851), .Z(n853) );
  XOR U450 ( .A(a[321]), .B(n838), .Z(n840) );
  XOR U451 ( .A(a[324]), .B(n826), .Z(n828) );
  XOR U452 ( .A(a[327]), .B(n814), .Z(n816) );
  XOR U453 ( .A(a[330]), .B(n801), .Z(n803) );
  XOR U454 ( .A(a[333]), .B(n789), .Z(n791) );
  XOR U455 ( .A(a[336]), .B(n777), .Z(n779) );
  XOR U456 ( .A(a[339]), .B(n764), .Z(n766) );
  XOR U457 ( .A(a[342]), .B(n752), .Z(n754) );
  XOR U458 ( .A(a[345]), .B(n740), .Z(n742) );
  XOR U459 ( .A(a[348]), .B(n728), .Z(n730) );
  XOR U460 ( .A(a[351]), .B(n715), .Z(n717) );
  XOR U461 ( .A(a[354]), .B(n703), .Z(n705) );
  XOR U462 ( .A(a[357]), .B(n691), .Z(n693) );
  XOR U463 ( .A(a[360]), .B(n678), .Z(n680) );
  XOR U464 ( .A(a[363]), .B(n666), .Z(n668) );
  XOR U465 ( .A(a[366]), .B(n654), .Z(n656) );
  XOR U466 ( .A(a[369]), .B(n641), .Z(n643) );
  XOR U467 ( .A(a[372]), .B(n629), .Z(n631) );
  XOR U468 ( .A(a[375]), .B(n617), .Z(n619) );
  XOR U469 ( .A(a[378]), .B(n605), .Z(n607) );
  XOR U470 ( .A(a[381]), .B(n592), .Z(n594) );
  XOR U471 ( .A(a[384]), .B(n580), .Z(n582) );
  XOR U472 ( .A(a[387]), .B(n568), .Z(n570) );
  XOR U473 ( .A(a[390]), .B(n555), .Z(n557) );
  XOR U474 ( .A(a[393]), .B(n543), .Z(n545) );
  XOR U475 ( .A(a[396]), .B(n531), .Z(n533) );
  XOR U476 ( .A(a[399]), .B(n517), .Z(n519) );
  XOR U477 ( .A(a[402]), .B(n505), .Z(n507) );
  XOR U478 ( .A(a[405]), .B(n493), .Z(n495) );
  XOR U479 ( .A(a[408]), .B(n481), .Z(n483) );
  XOR U480 ( .A(a[411]), .B(n468), .Z(n470) );
  XOR U481 ( .A(a[414]), .B(n456), .Z(n458) );
  XOR U482 ( .A(a[417]), .B(n444), .Z(n446) );
  XOR U483 ( .A(a[420]), .B(n431), .Z(n433) );
  XOR U484 ( .A(a[423]), .B(n419), .Z(n421) );
  XOR U485 ( .A(a[426]), .B(n407), .Z(n409) );
  XOR U486 ( .A(a[429]), .B(n394), .Z(n396) );
  XOR U487 ( .A(a[432]), .B(n382), .Z(n384) );
  XOR U488 ( .A(a[435]), .B(n370), .Z(n372) );
  XOR U489 ( .A(a[438]), .B(n358), .Z(n360) );
  XOR U490 ( .A(a[441]), .B(n345), .Z(n347) );
  XOR U491 ( .A(a[444]), .B(n333), .Z(n335) );
  XOR U492 ( .A(a[447]), .B(n321), .Z(n323) );
  XOR U493 ( .A(a[450]), .B(n308), .Z(n310) );
  XOR U494 ( .A(a[453]), .B(n296), .Z(n298) );
  XOR U495 ( .A(a[456]), .B(n284), .Z(n286) );
  XOR U496 ( .A(a[459]), .B(n271), .Z(n273) );
  XOR U497 ( .A(a[462]), .B(n259), .Z(n261) );
  XOR U498 ( .A(a[465]), .B(n247), .Z(n249) );
  XOR U499 ( .A(a[468]), .B(n235), .Z(n237) );
  XOR U500 ( .A(a[471]), .B(n222), .Z(n224) );
  XOR U501 ( .A(a[474]), .B(n210), .Z(n212) );
  XOR U502 ( .A(a[477]), .B(n198), .Z(n200) );
  XOR U503 ( .A(a[480]), .B(n185), .Z(n187) );
  XOR U504 ( .A(a[483]), .B(n173), .Z(n175) );
  XOR U505 ( .A(a[486]), .B(n161), .Z(n163) );
  XOR U506 ( .A(a[489]), .B(n148), .Z(n150) );
  XOR U507 ( .A(a[492]), .B(n136), .Z(n138) );
  XOR U508 ( .A(a[495]), .B(n124), .Z(n126) );
  XOR U509 ( .A(a[498]), .B(n112), .Z(n114) );
  XOR U510 ( .A(a[501]), .B(n98), .Z(n100) );
  XOR U511 ( .A(a[504]), .B(n86), .Z(n88) );
  XOR U512 ( .A(a[507]), .B(n74), .Z(n76) );
  XOR U513 ( .A(a[510]), .B(n61), .Z(n63) );
  XOR U514 ( .A(n2), .B(n3), .Z(carry_on_d) );
  ANDN U515 ( .B(n4), .A(n5), .Z(n2) );
  XOR U516 ( .A(b[511]), .B(n3), .Z(n4) );
  XNOR U517 ( .A(b[9]), .B(n6), .Z(c[9]) );
  XNOR U518 ( .A(b[99]), .B(n7), .Z(c[99]) );
  XNOR U519 ( .A(b[98]), .B(n8), .Z(c[98]) );
  XNOR U520 ( .A(b[97]), .B(n9), .Z(c[97]) );
  XNOR U521 ( .A(b[96]), .B(n10), .Z(c[96]) );
  XNOR U522 ( .A(b[95]), .B(n11), .Z(c[95]) );
  XNOR U523 ( .A(b[94]), .B(n12), .Z(c[94]) );
  XNOR U524 ( .A(b[93]), .B(n13), .Z(c[93]) );
  XNOR U525 ( .A(b[92]), .B(n14), .Z(c[92]) );
  XNOR U526 ( .A(b[91]), .B(n15), .Z(c[91]) );
  XNOR U527 ( .A(b[90]), .B(n16), .Z(c[90]) );
  XNOR U528 ( .A(b[8]), .B(n17), .Z(c[8]) );
  XNOR U529 ( .A(b[89]), .B(n18), .Z(c[89]) );
  XNOR U530 ( .A(b[88]), .B(n19), .Z(c[88]) );
  XNOR U531 ( .A(b[87]), .B(n20), .Z(c[87]) );
  XNOR U532 ( .A(b[86]), .B(n21), .Z(c[86]) );
  XNOR U533 ( .A(b[85]), .B(n22), .Z(c[85]) );
  XNOR U534 ( .A(b[84]), .B(n23), .Z(c[84]) );
  XNOR U535 ( .A(b[83]), .B(n24), .Z(c[83]) );
  XNOR U536 ( .A(b[82]), .B(n25), .Z(c[82]) );
  XNOR U537 ( .A(b[81]), .B(n26), .Z(c[81]) );
  XNOR U538 ( .A(b[80]), .B(n27), .Z(c[80]) );
  XNOR U539 ( .A(b[7]), .B(n28), .Z(c[7]) );
  XNOR U540 ( .A(b[79]), .B(n29), .Z(c[79]) );
  XNOR U541 ( .A(b[78]), .B(n30), .Z(c[78]) );
  XNOR U542 ( .A(b[77]), .B(n31), .Z(c[77]) );
  XNOR U543 ( .A(b[76]), .B(n32), .Z(c[76]) );
  XNOR U544 ( .A(b[75]), .B(n33), .Z(c[75]) );
  XNOR U545 ( .A(b[74]), .B(n34), .Z(c[74]) );
  XNOR U546 ( .A(b[73]), .B(n35), .Z(c[73]) );
  XNOR U547 ( .A(b[72]), .B(n36), .Z(c[72]) );
  XNOR U548 ( .A(b[71]), .B(n37), .Z(c[71]) );
  XNOR U549 ( .A(b[70]), .B(n38), .Z(c[70]) );
  XNOR U550 ( .A(b[6]), .B(n39), .Z(c[6]) );
  XNOR U551 ( .A(b[69]), .B(n40), .Z(c[69]) );
  XNOR U552 ( .A(b[68]), .B(n41), .Z(c[68]) );
  XNOR U553 ( .A(b[67]), .B(n42), .Z(c[67]) );
  XNOR U554 ( .A(b[66]), .B(n43), .Z(c[66]) );
  XNOR U555 ( .A(b[65]), .B(n44), .Z(c[65]) );
  XNOR U556 ( .A(b[64]), .B(n45), .Z(c[64]) );
  XNOR U557 ( .A(b[63]), .B(n46), .Z(c[63]) );
  XNOR U558 ( .A(b[62]), .B(n47), .Z(c[62]) );
  XNOR U559 ( .A(b[61]), .B(n48), .Z(c[61]) );
  XNOR U560 ( .A(b[60]), .B(n49), .Z(c[60]) );
  XNOR U561 ( .A(b[5]), .B(n50), .Z(c[5]) );
  XNOR U562 ( .A(b[59]), .B(n51), .Z(c[59]) );
  XNOR U563 ( .A(b[58]), .B(n52), .Z(c[58]) );
  XNOR U564 ( .A(b[57]), .B(n53), .Z(c[57]) );
  XNOR U565 ( .A(b[56]), .B(n54), .Z(c[56]) );
  XNOR U566 ( .A(b[55]), .B(n55), .Z(c[55]) );
  XNOR U567 ( .A(b[54]), .B(n56), .Z(c[54]) );
  XNOR U568 ( .A(b[53]), .B(n57), .Z(c[53]) );
  XNOR U569 ( .A(b[52]), .B(n58), .Z(c[52]) );
  XNOR U570 ( .A(b[51]), .B(n59), .Z(c[51]) );
  XNOR U571 ( .A(b[511]), .B(n5), .Z(c[511]) );
  XNOR U572 ( .A(a[511]), .B(n3), .Z(n5) );
  XNOR U573 ( .A(n60), .B(n61), .Z(n3) );
  ANDN U574 ( .B(n62), .A(n63), .Z(n60) );
  XNOR U575 ( .A(b[510]), .B(n61), .Z(n62) );
  XNOR U576 ( .A(b[510]), .B(n63), .Z(c[510]) );
  XOR U577 ( .A(n64), .B(n65), .Z(n61) );
  ANDN U578 ( .B(n66), .A(n67), .Z(n64) );
  XNOR U579 ( .A(b[509]), .B(n65), .Z(n66) );
  XNOR U580 ( .A(b[50]), .B(n68), .Z(c[50]) );
  XNOR U581 ( .A(b[509]), .B(n67), .Z(c[509]) );
  XOR U582 ( .A(n69), .B(n70), .Z(n65) );
  ANDN U583 ( .B(n71), .A(n72), .Z(n69) );
  XNOR U584 ( .A(b[508]), .B(n70), .Z(n71) );
  XNOR U585 ( .A(b[508]), .B(n72), .Z(c[508]) );
  XOR U586 ( .A(n73), .B(n74), .Z(n70) );
  ANDN U587 ( .B(n75), .A(n76), .Z(n73) );
  XNOR U588 ( .A(b[507]), .B(n74), .Z(n75) );
  XNOR U589 ( .A(b[507]), .B(n76), .Z(c[507]) );
  XOR U590 ( .A(n77), .B(n78), .Z(n74) );
  ANDN U591 ( .B(n79), .A(n80), .Z(n77) );
  XNOR U592 ( .A(b[506]), .B(n78), .Z(n79) );
  XNOR U593 ( .A(b[506]), .B(n80), .Z(c[506]) );
  XOR U594 ( .A(n81), .B(n82), .Z(n78) );
  ANDN U595 ( .B(n83), .A(n84), .Z(n81) );
  XNOR U596 ( .A(b[505]), .B(n82), .Z(n83) );
  XNOR U597 ( .A(b[505]), .B(n84), .Z(c[505]) );
  XOR U598 ( .A(n85), .B(n86), .Z(n82) );
  ANDN U599 ( .B(n87), .A(n88), .Z(n85) );
  XNOR U600 ( .A(b[504]), .B(n86), .Z(n87) );
  XNOR U601 ( .A(b[504]), .B(n88), .Z(c[504]) );
  XOR U602 ( .A(n89), .B(n90), .Z(n86) );
  ANDN U603 ( .B(n91), .A(n92), .Z(n89) );
  XNOR U604 ( .A(b[503]), .B(n90), .Z(n91) );
  XNOR U605 ( .A(b[503]), .B(n92), .Z(c[503]) );
  XOR U606 ( .A(n93), .B(n94), .Z(n90) );
  ANDN U607 ( .B(n95), .A(n96), .Z(n93) );
  XNOR U608 ( .A(b[502]), .B(n94), .Z(n95) );
  XNOR U609 ( .A(b[502]), .B(n96), .Z(c[502]) );
  XOR U610 ( .A(n97), .B(n98), .Z(n94) );
  ANDN U611 ( .B(n99), .A(n100), .Z(n97) );
  XNOR U612 ( .A(b[501]), .B(n98), .Z(n99) );
  XNOR U613 ( .A(b[501]), .B(n100), .Z(c[501]) );
  XOR U614 ( .A(n101), .B(n102), .Z(n98) );
  ANDN U615 ( .B(n103), .A(n104), .Z(n101) );
  XNOR U616 ( .A(b[500]), .B(n102), .Z(n103) );
  XNOR U617 ( .A(b[500]), .B(n104), .Z(c[500]) );
  XOR U618 ( .A(n105), .B(n106), .Z(n102) );
  ANDN U619 ( .B(n107), .A(n108), .Z(n105) );
  XNOR U620 ( .A(b[499]), .B(n106), .Z(n107) );
  XNOR U621 ( .A(b[4]), .B(n109), .Z(c[4]) );
  XNOR U622 ( .A(b[49]), .B(n110), .Z(c[49]) );
  XNOR U623 ( .A(b[499]), .B(n108), .Z(c[499]) );
  XOR U624 ( .A(n111), .B(n112), .Z(n106) );
  ANDN U625 ( .B(n113), .A(n114), .Z(n111) );
  XNOR U626 ( .A(b[498]), .B(n112), .Z(n113) );
  XNOR U627 ( .A(b[498]), .B(n114), .Z(c[498]) );
  XOR U628 ( .A(n115), .B(n116), .Z(n112) );
  ANDN U629 ( .B(n117), .A(n118), .Z(n115) );
  XNOR U630 ( .A(b[497]), .B(n116), .Z(n117) );
  XNOR U631 ( .A(b[497]), .B(n118), .Z(c[497]) );
  XOR U632 ( .A(n119), .B(n120), .Z(n116) );
  ANDN U633 ( .B(n121), .A(n122), .Z(n119) );
  XNOR U634 ( .A(b[496]), .B(n120), .Z(n121) );
  XNOR U635 ( .A(b[496]), .B(n122), .Z(c[496]) );
  XOR U636 ( .A(n123), .B(n124), .Z(n120) );
  ANDN U637 ( .B(n125), .A(n126), .Z(n123) );
  XNOR U638 ( .A(b[495]), .B(n124), .Z(n125) );
  XNOR U639 ( .A(b[495]), .B(n126), .Z(c[495]) );
  XOR U640 ( .A(n127), .B(n128), .Z(n124) );
  ANDN U641 ( .B(n129), .A(n130), .Z(n127) );
  XNOR U642 ( .A(b[494]), .B(n128), .Z(n129) );
  XNOR U643 ( .A(b[494]), .B(n130), .Z(c[494]) );
  XOR U644 ( .A(n131), .B(n132), .Z(n128) );
  ANDN U645 ( .B(n133), .A(n134), .Z(n131) );
  XNOR U646 ( .A(b[493]), .B(n132), .Z(n133) );
  XNOR U647 ( .A(b[493]), .B(n134), .Z(c[493]) );
  XOR U648 ( .A(n135), .B(n136), .Z(n132) );
  ANDN U649 ( .B(n137), .A(n138), .Z(n135) );
  XNOR U650 ( .A(b[492]), .B(n136), .Z(n137) );
  XNOR U651 ( .A(b[492]), .B(n138), .Z(c[492]) );
  XOR U652 ( .A(n139), .B(n140), .Z(n136) );
  ANDN U653 ( .B(n141), .A(n142), .Z(n139) );
  XNOR U654 ( .A(b[491]), .B(n140), .Z(n141) );
  XNOR U655 ( .A(b[491]), .B(n142), .Z(c[491]) );
  XOR U656 ( .A(n143), .B(n144), .Z(n140) );
  ANDN U657 ( .B(n145), .A(n146), .Z(n143) );
  XNOR U658 ( .A(b[490]), .B(n144), .Z(n145) );
  XNOR U659 ( .A(b[490]), .B(n146), .Z(c[490]) );
  XOR U660 ( .A(n147), .B(n148), .Z(n144) );
  ANDN U661 ( .B(n149), .A(n150), .Z(n147) );
  XNOR U662 ( .A(b[489]), .B(n148), .Z(n149) );
  XNOR U663 ( .A(b[48]), .B(n151), .Z(c[48]) );
  XNOR U664 ( .A(b[489]), .B(n150), .Z(c[489]) );
  XOR U665 ( .A(n152), .B(n153), .Z(n148) );
  ANDN U666 ( .B(n154), .A(n155), .Z(n152) );
  XNOR U667 ( .A(b[488]), .B(n153), .Z(n154) );
  XNOR U668 ( .A(b[488]), .B(n155), .Z(c[488]) );
  XOR U669 ( .A(n156), .B(n157), .Z(n153) );
  ANDN U670 ( .B(n158), .A(n159), .Z(n156) );
  XNOR U671 ( .A(b[487]), .B(n157), .Z(n158) );
  XNOR U672 ( .A(b[487]), .B(n159), .Z(c[487]) );
  XOR U673 ( .A(n160), .B(n161), .Z(n157) );
  ANDN U674 ( .B(n162), .A(n163), .Z(n160) );
  XNOR U675 ( .A(b[486]), .B(n161), .Z(n162) );
  XNOR U676 ( .A(b[486]), .B(n163), .Z(c[486]) );
  XOR U677 ( .A(n164), .B(n165), .Z(n161) );
  ANDN U678 ( .B(n166), .A(n167), .Z(n164) );
  XNOR U679 ( .A(b[485]), .B(n165), .Z(n166) );
  XNOR U680 ( .A(b[485]), .B(n167), .Z(c[485]) );
  XOR U681 ( .A(n168), .B(n169), .Z(n165) );
  ANDN U682 ( .B(n170), .A(n171), .Z(n168) );
  XNOR U683 ( .A(b[484]), .B(n169), .Z(n170) );
  XNOR U684 ( .A(b[484]), .B(n171), .Z(c[484]) );
  XOR U685 ( .A(n172), .B(n173), .Z(n169) );
  ANDN U686 ( .B(n174), .A(n175), .Z(n172) );
  XNOR U687 ( .A(b[483]), .B(n173), .Z(n174) );
  XNOR U688 ( .A(b[483]), .B(n175), .Z(c[483]) );
  XOR U689 ( .A(n176), .B(n177), .Z(n173) );
  ANDN U690 ( .B(n178), .A(n179), .Z(n176) );
  XNOR U691 ( .A(b[482]), .B(n177), .Z(n178) );
  XNOR U692 ( .A(b[482]), .B(n179), .Z(c[482]) );
  XOR U693 ( .A(n180), .B(n181), .Z(n177) );
  ANDN U694 ( .B(n182), .A(n183), .Z(n180) );
  XNOR U695 ( .A(b[481]), .B(n181), .Z(n182) );
  XNOR U696 ( .A(b[481]), .B(n183), .Z(c[481]) );
  XOR U697 ( .A(n184), .B(n185), .Z(n181) );
  ANDN U698 ( .B(n186), .A(n187), .Z(n184) );
  XNOR U699 ( .A(b[480]), .B(n185), .Z(n186) );
  XNOR U700 ( .A(b[480]), .B(n187), .Z(c[480]) );
  XOR U701 ( .A(n188), .B(n189), .Z(n185) );
  ANDN U702 ( .B(n190), .A(n191), .Z(n188) );
  XNOR U703 ( .A(b[479]), .B(n189), .Z(n190) );
  XNOR U704 ( .A(b[47]), .B(n192), .Z(c[47]) );
  XNOR U705 ( .A(b[479]), .B(n191), .Z(c[479]) );
  XOR U706 ( .A(n193), .B(n194), .Z(n189) );
  ANDN U707 ( .B(n195), .A(n196), .Z(n193) );
  XNOR U708 ( .A(b[478]), .B(n194), .Z(n195) );
  XNOR U709 ( .A(b[478]), .B(n196), .Z(c[478]) );
  XOR U710 ( .A(n197), .B(n198), .Z(n194) );
  ANDN U711 ( .B(n199), .A(n200), .Z(n197) );
  XNOR U712 ( .A(b[477]), .B(n198), .Z(n199) );
  XNOR U713 ( .A(b[477]), .B(n200), .Z(c[477]) );
  XOR U714 ( .A(n201), .B(n202), .Z(n198) );
  ANDN U715 ( .B(n203), .A(n204), .Z(n201) );
  XNOR U716 ( .A(b[476]), .B(n202), .Z(n203) );
  XNOR U717 ( .A(b[476]), .B(n204), .Z(c[476]) );
  XOR U718 ( .A(n205), .B(n206), .Z(n202) );
  ANDN U719 ( .B(n207), .A(n208), .Z(n205) );
  XNOR U720 ( .A(b[475]), .B(n206), .Z(n207) );
  XNOR U721 ( .A(b[475]), .B(n208), .Z(c[475]) );
  XOR U722 ( .A(n209), .B(n210), .Z(n206) );
  ANDN U723 ( .B(n211), .A(n212), .Z(n209) );
  XNOR U724 ( .A(b[474]), .B(n210), .Z(n211) );
  XNOR U725 ( .A(b[474]), .B(n212), .Z(c[474]) );
  XOR U726 ( .A(n213), .B(n214), .Z(n210) );
  ANDN U727 ( .B(n215), .A(n216), .Z(n213) );
  XNOR U728 ( .A(b[473]), .B(n214), .Z(n215) );
  XNOR U729 ( .A(b[473]), .B(n216), .Z(c[473]) );
  XOR U730 ( .A(n217), .B(n218), .Z(n214) );
  ANDN U731 ( .B(n219), .A(n220), .Z(n217) );
  XNOR U732 ( .A(b[472]), .B(n218), .Z(n219) );
  XNOR U733 ( .A(b[472]), .B(n220), .Z(c[472]) );
  XOR U734 ( .A(n221), .B(n222), .Z(n218) );
  ANDN U735 ( .B(n223), .A(n224), .Z(n221) );
  XNOR U736 ( .A(b[471]), .B(n222), .Z(n223) );
  XNOR U737 ( .A(b[471]), .B(n224), .Z(c[471]) );
  XOR U738 ( .A(n225), .B(n226), .Z(n222) );
  ANDN U739 ( .B(n227), .A(n228), .Z(n225) );
  XNOR U740 ( .A(b[470]), .B(n226), .Z(n227) );
  XNOR U741 ( .A(b[470]), .B(n228), .Z(c[470]) );
  XOR U742 ( .A(n229), .B(n230), .Z(n226) );
  ANDN U743 ( .B(n231), .A(n232), .Z(n229) );
  XNOR U744 ( .A(b[469]), .B(n230), .Z(n231) );
  XNOR U745 ( .A(b[46]), .B(n233), .Z(c[46]) );
  XNOR U746 ( .A(b[469]), .B(n232), .Z(c[469]) );
  XOR U747 ( .A(n234), .B(n235), .Z(n230) );
  ANDN U748 ( .B(n236), .A(n237), .Z(n234) );
  XNOR U749 ( .A(b[468]), .B(n235), .Z(n236) );
  XNOR U750 ( .A(b[468]), .B(n237), .Z(c[468]) );
  XOR U751 ( .A(n238), .B(n239), .Z(n235) );
  ANDN U752 ( .B(n240), .A(n241), .Z(n238) );
  XNOR U753 ( .A(b[467]), .B(n239), .Z(n240) );
  XNOR U754 ( .A(b[467]), .B(n241), .Z(c[467]) );
  XOR U755 ( .A(n242), .B(n243), .Z(n239) );
  ANDN U756 ( .B(n244), .A(n245), .Z(n242) );
  XNOR U757 ( .A(b[466]), .B(n243), .Z(n244) );
  XNOR U758 ( .A(b[466]), .B(n245), .Z(c[466]) );
  XOR U759 ( .A(n246), .B(n247), .Z(n243) );
  ANDN U760 ( .B(n248), .A(n249), .Z(n246) );
  XNOR U761 ( .A(b[465]), .B(n247), .Z(n248) );
  XNOR U762 ( .A(b[465]), .B(n249), .Z(c[465]) );
  XOR U763 ( .A(n250), .B(n251), .Z(n247) );
  ANDN U764 ( .B(n252), .A(n253), .Z(n250) );
  XNOR U765 ( .A(b[464]), .B(n251), .Z(n252) );
  XNOR U766 ( .A(b[464]), .B(n253), .Z(c[464]) );
  XOR U767 ( .A(n254), .B(n255), .Z(n251) );
  ANDN U768 ( .B(n256), .A(n257), .Z(n254) );
  XNOR U769 ( .A(b[463]), .B(n255), .Z(n256) );
  XNOR U770 ( .A(b[463]), .B(n257), .Z(c[463]) );
  XOR U771 ( .A(n258), .B(n259), .Z(n255) );
  ANDN U772 ( .B(n260), .A(n261), .Z(n258) );
  XNOR U773 ( .A(b[462]), .B(n259), .Z(n260) );
  XNOR U774 ( .A(b[462]), .B(n261), .Z(c[462]) );
  XOR U775 ( .A(n262), .B(n263), .Z(n259) );
  ANDN U776 ( .B(n264), .A(n265), .Z(n262) );
  XNOR U777 ( .A(b[461]), .B(n263), .Z(n264) );
  XNOR U778 ( .A(b[461]), .B(n265), .Z(c[461]) );
  XOR U779 ( .A(n266), .B(n267), .Z(n263) );
  ANDN U780 ( .B(n268), .A(n269), .Z(n266) );
  XNOR U781 ( .A(b[460]), .B(n267), .Z(n268) );
  XNOR U782 ( .A(b[460]), .B(n269), .Z(c[460]) );
  XOR U783 ( .A(n270), .B(n271), .Z(n267) );
  ANDN U784 ( .B(n272), .A(n273), .Z(n270) );
  XNOR U785 ( .A(b[459]), .B(n271), .Z(n272) );
  XNOR U786 ( .A(b[45]), .B(n274), .Z(c[45]) );
  XNOR U787 ( .A(b[459]), .B(n273), .Z(c[459]) );
  XOR U788 ( .A(n275), .B(n276), .Z(n271) );
  ANDN U789 ( .B(n277), .A(n278), .Z(n275) );
  XNOR U790 ( .A(b[458]), .B(n276), .Z(n277) );
  XNOR U791 ( .A(b[458]), .B(n278), .Z(c[458]) );
  XOR U792 ( .A(n279), .B(n280), .Z(n276) );
  ANDN U793 ( .B(n281), .A(n282), .Z(n279) );
  XNOR U794 ( .A(b[457]), .B(n280), .Z(n281) );
  XNOR U795 ( .A(b[457]), .B(n282), .Z(c[457]) );
  XOR U796 ( .A(n283), .B(n284), .Z(n280) );
  ANDN U797 ( .B(n285), .A(n286), .Z(n283) );
  XNOR U798 ( .A(b[456]), .B(n284), .Z(n285) );
  XNOR U799 ( .A(b[456]), .B(n286), .Z(c[456]) );
  XOR U800 ( .A(n287), .B(n288), .Z(n284) );
  ANDN U801 ( .B(n289), .A(n290), .Z(n287) );
  XNOR U802 ( .A(b[455]), .B(n288), .Z(n289) );
  XNOR U803 ( .A(b[455]), .B(n290), .Z(c[455]) );
  XOR U804 ( .A(n291), .B(n292), .Z(n288) );
  ANDN U805 ( .B(n293), .A(n294), .Z(n291) );
  XNOR U806 ( .A(b[454]), .B(n292), .Z(n293) );
  XNOR U807 ( .A(b[454]), .B(n294), .Z(c[454]) );
  XOR U808 ( .A(n295), .B(n296), .Z(n292) );
  ANDN U809 ( .B(n297), .A(n298), .Z(n295) );
  XNOR U810 ( .A(b[453]), .B(n296), .Z(n297) );
  XNOR U811 ( .A(b[453]), .B(n298), .Z(c[453]) );
  XOR U812 ( .A(n299), .B(n300), .Z(n296) );
  ANDN U813 ( .B(n301), .A(n302), .Z(n299) );
  XNOR U814 ( .A(b[452]), .B(n300), .Z(n301) );
  XNOR U815 ( .A(b[452]), .B(n302), .Z(c[452]) );
  XOR U816 ( .A(n303), .B(n304), .Z(n300) );
  ANDN U817 ( .B(n305), .A(n306), .Z(n303) );
  XNOR U818 ( .A(b[451]), .B(n304), .Z(n305) );
  XNOR U819 ( .A(b[451]), .B(n306), .Z(c[451]) );
  XOR U820 ( .A(n307), .B(n308), .Z(n304) );
  ANDN U821 ( .B(n309), .A(n310), .Z(n307) );
  XNOR U822 ( .A(b[450]), .B(n308), .Z(n309) );
  XNOR U823 ( .A(b[450]), .B(n310), .Z(c[450]) );
  XOR U824 ( .A(n311), .B(n312), .Z(n308) );
  ANDN U825 ( .B(n313), .A(n314), .Z(n311) );
  XNOR U826 ( .A(b[449]), .B(n312), .Z(n313) );
  XNOR U827 ( .A(b[44]), .B(n315), .Z(c[44]) );
  XNOR U828 ( .A(b[449]), .B(n314), .Z(c[449]) );
  XOR U829 ( .A(n316), .B(n317), .Z(n312) );
  ANDN U830 ( .B(n318), .A(n319), .Z(n316) );
  XNOR U831 ( .A(b[448]), .B(n317), .Z(n318) );
  XNOR U832 ( .A(b[448]), .B(n319), .Z(c[448]) );
  XOR U833 ( .A(n320), .B(n321), .Z(n317) );
  ANDN U834 ( .B(n322), .A(n323), .Z(n320) );
  XNOR U835 ( .A(b[447]), .B(n321), .Z(n322) );
  XNOR U836 ( .A(b[447]), .B(n323), .Z(c[447]) );
  XOR U837 ( .A(n324), .B(n325), .Z(n321) );
  ANDN U838 ( .B(n326), .A(n327), .Z(n324) );
  XNOR U839 ( .A(b[446]), .B(n325), .Z(n326) );
  XNOR U840 ( .A(b[446]), .B(n327), .Z(c[446]) );
  XOR U841 ( .A(n328), .B(n329), .Z(n325) );
  ANDN U842 ( .B(n330), .A(n331), .Z(n328) );
  XNOR U843 ( .A(b[445]), .B(n329), .Z(n330) );
  XNOR U844 ( .A(b[445]), .B(n331), .Z(c[445]) );
  XOR U845 ( .A(n332), .B(n333), .Z(n329) );
  ANDN U846 ( .B(n334), .A(n335), .Z(n332) );
  XNOR U847 ( .A(b[444]), .B(n333), .Z(n334) );
  XNOR U848 ( .A(b[444]), .B(n335), .Z(c[444]) );
  XOR U849 ( .A(n336), .B(n337), .Z(n333) );
  ANDN U850 ( .B(n338), .A(n339), .Z(n336) );
  XNOR U851 ( .A(b[443]), .B(n337), .Z(n338) );
  XNOR U852 ( .A(b[443]), .B(n339), .Z(c[443]) );
  XOR U853 ( .A(n340), .B(n341), .Z(n337) );
  ANDN U854 ( .B(n342), .A(n343), .Z(n340) );
  XNOR U855 ( .A(b[442]), .B(n341), .Z(n342) );
  XNOR U856 ( .A(b[442]), .B(n343), .Z(c[442]) );
  XOR U857 ( .A(n344), .B(n345), .Z(n341) );
  ANDN U858 ( .B(n346), .A(n347), .Z(n344) );
  XNOR U859 ( .A(b[441]), .B(n345), .Z(n346) );
  XNOR U860 ( .A(b[441]), .B(n347), .Z(c[441]) );
  XOR U861 ( .A(n348), .B(n349), .Z(n345) );
  ANDN U862 ( .B(n350), .A(n351), .Z(n348) );
  XNOR U863 ( .A(b[440]), .B(n349), .Z(n350) );
  XNOR U864 ( .A(b[440]), .B(n351), .Z(c[440]) );
  XOR U865 ( .A(n352), .B(n353), .Z(n349) );
  ANDN U866 ( .B(n354), .A(n355), .Z(n352) );
  XNOR U867 ( .A(b[439]), .B(n353), .Z(n354) );
  XNOR U868 ( .A(b[43]), .B(n356), .Z(c[43]) );
  XNOR U869 ( .A(b[439]), .B(n355), .Z(c[439]) );
  XOR U870 ( .A(n357), .B(n358), .Z(n353) );
  ANDN U871 ( .B(n359), .A(n360), .Z(n357) );
  XNOR U872 ( .A(b[438]), .B(n358), .Z(n359) );
  XNOR U873 ( .A(b[438]), .B(n360), .Z(c[438]) );
  XOR U874 ( .A(n361), .B(n362), .Z(n358) );
  ANDN U875 ( .B(n363), .A(n364), .Z(n361) );
  XNOR U876 ( .A(b[437]), .B(n362), .Z(n363) );
  XNOR U877 ( .A(b[437]), .B(n364), .Z(c[437]) );
  XOR U878 ( .A(n365), .B(n366), .Z(n362) );
  ANDN U879 ( .B(n367), .A(n368), .Z(n365) );
  XNOR U880 ( .A(b[436]), .B(n366), .Z(n367) );
  XNOR U881 ( .A(b[436]), .B(n368), .Z(c[436]) );
  XOR U882 ( .A(n369), .B(n370), .Z(n366) );
  ANDN U883 ( .B(n371), .A(n372), .Z(n369) );
  XNOR U884 ( .A(b[435]), .B(n370), .Z(n371) );
  XNOR U885 ( .A(b[435]), .B(n372), .Z(c[435]) );
  XOR U886 ( .A(n373), .B(n374), .Z(n370) );
  ANDN U887 ( .B(n375), .A(n376), .Z(n373) );
  XNOR U888 ( .A(b[434]), .B(n374), .Z(n375) );
  XNOR U889 ( .A(b[434]), .B(n376), .Z(c[434]) );
  XOR U890 ( .A(n377), .B(n378), .Z(n374) );
  ANDN U891 ( .B(n379), .A(n380), .Z(n377) );
  XNOR U892 ( .A(b[433]), .B(n378), .Z(n379) );
  XNOR U893 ( .A(b[433]), .B(n380), .Z(c[433]) );
  XOR U894 ( .A(n381), .B(n382), .Z(n378) );
  ANDN U895 ( .B(n383), .A(n384), .Z(n381) );
  XNOR U896 ( .A(b[432]), .B(n382), .Z(n383) );
  XNOR U897 ( .A(b[432]), .B(n384), .Z(c[432]) );
  XOR U898 ( .A(n385), .B(n386), .Z(n382) );
  ANDN U899 ( .B(n387), .A(n388), .Z(n385) );
  XNOR U900 ( .A(b[431]), .B(n386), .Z(n387) );
  XNOR U901 ( .A(b[431]), .B(n388), .Z(c[431]) );
  XOR U902 ( .A(n389), .B(n390), .Z(n386) );
  ANDN U903 ( .B(n391), .A(n392), .Z(n389) );
  XNOR U904 ( .A(b[430]), .B(n390), .Z(n391) );
  XNOR U905 ( .A(b[430]), .B(n392), .Z(c[430]) );
  XOR U906 ( .A(n393), .B(n394), .Z(n390) );
  ANDN U907 ( .B(n395), .A(n396), .Z(n393) );
  XNOR U908 ( .A(b[429]), .B(n394), .Z(n395) );
  XNOR U909 ( .A(b[42]), .B(n397), .Z(c[42]) );
  XNOR U910 ( .A(b[429]), .B(n396), .Z(c[429]) );
  XOR U911 ( .A(n398), .B(n399), .Z(n394) );
  ANDN U912 ( .B(n400), .A(n401), .Z(n398) );
  XNOR U913 ( .A(b[428]), .B(n399), .Z(n400) );
  XNOR U914 ( .A(b[428]), .B(n401), .Z(c[428]) );
  XOR U915 ( .A(n402), .B(n403), .Z(n399) );
  ANDN U916 ( .B(n404), .A(n405), .Z(n402) );
  XNOR U917 ( .A(b[427]), .B(n403), .Z(n404) );
  XNOR U918 ( .A(b[427]), .B(n405), .Z(c[427]) );
  XOR U919 ( .A(n406), .B(n407), .Z(n403) );
  ANDN U920 ( .B(n408), .A(n409), .Z(n406) );
  XNOR U921 ( .A(b[426]), .B(n407), .Z(n408) );
  XNOR U922 ( .A(b[426]), .B(n409), .Z(c[426]) );
  XOR U923 ( .A(n410), .B(n411), .Z(n407) );
  ANDN U924 ( .B(n412), .A(n413), .Z(n410) );
  XNOR U925 ( .A(b[425]), .B(n411), .Z(n412) );
  XNOR U926 ( .A(b[425]), .B(n413), .Z(c[425]) );
  XOR U927 ( .A(n414), .B(n415), .Z(n411) );
  ANDN U928 ( .B(n416), .A(n417), .Z(n414) );
  XNOR U929 ( .A(b[424]), .B(n415), .Z(n416) );
  XNOR U930 ( .A(b[424]), .B(n417), .Z(c[424]) );
  XOR U931 ( .A(n418), .B(n419), .Z(n415) );
  ANDN U932 ( .B(n420), .A(n421), .Z(n418) );
  XNOR U933 ( .A(b[423]), .B(n419), .Z(n420) );
  XNOR U934 ( .A(b[423]), .B(n421), .Z(c[423]) );
  XOR U935 ( .A(n422), .B(n423), .Z(n419) );
  ANDN U936 ( .B(n424), .A(n425), .Z(n422) );
  XNOR U937 ( .A(b[422]), .B(n423), .Z(n424) );
  XNOR U938 ( .A(b[422]), .B(n425), .Z(c[422]) );
  XOR U939 ( .A(n426), .B(n427), .Z(n423) );
  ANDN U940 ( .B(n428), .A(n429), .Z(n426) );
  XNOR U941 ( .A(b[421]), .B(n427), .Z(n428) );
  XNOR U942 ( .A(b[421]), .B(n429), .Z(c[421]) );
  XOR U943 ( .A(n430), .B(n431), .Z(n427) );
  ANDN U944 ( .B(n432), .A(n433), .Z(n430) );
  XNOR U945 ( .A(b[420]), .B(n431), .Z(n432) );
  XNOR U946 ( .A(b[420]), .B(n433), .Z(c[420]) );
  XOR U947 ( .A(n434), .B(n435), .Z(n431) );
  ANDN U948 ( .B(n436), .A(n437), .Z(n434) );
  XNOR U949 ( .A(b[419]), .B(n435), .Z(n436) );
  XNOR U950 ( .A(b[41]), .B(n438), .Z(c[41]) );
  XNOR U951 ( .A(b[419]), .B(n437), .Z(c[419]) );
  XOR U952 ( .A(n439), .B(n440), .Z(n435) );
  ANDN U953 ( .B(n441), .A(n442), .Z(n439) );
  XNOR U954 ( .A(b[418]), .B(n440), .Z(n441) );
  XNOR U955 ( .A(b[418]), .B(n442), .Z(c[418]) );
  XOR U956 ( .A(n443), .B(n444), .Z(n440) );
  ANDN U957 ( .B(n445), .A(n446), .Z(n443) );
  XNOR U958 ( .A(b[417]), .B(n444), .Z(n445) );
  XNOR U959 ( .A(b[417]), .B(n446), .Z(c[417]) );
  XOR U960 ( .A(n447), .B(n448), .Z(n444) );
  ANDN U961 ( .B(n449), .A(n450), .Z(n447) );
  XNOR U962 ( .A(b[416]), .B(n448), .Z(n449) );
  XNOR U963 ( .A(b[416]), .B(n450), .Z(c[416]) );
  XOR U964 ( .A(n451), .B(n452), .Z(n448) );
  ANDN U965 ( .B(n453), .A(n454), .Z(n451) );
  XNOR U966 ( .A(b[415]), .B(n452), .Z(n453) );
  XNOR U967 ( .A(b[415]), .B(n454), .Z(c[415]) );
  XOR U968 ( .A(n455), .B(n456), .Z(n452) );
  ANDN U969 ( .B(n457), .A(n458), .Z(n455) );
  XNOR U970 ( .A(b[414]), .B(n456), .Z(n457) );
  XNOR U971 ( .A(b[414]), .B(n458), .Z(c[414]) );
  XOR U972 ( .A(n459), .B(n460), .Z(n456) );
  ANDN U973 ( .B(n461), .A(n462), .Z(n459) );
  XNOR U974 ( .A(b[413]), .B(n460), .Z(n461) );
  XNOR U975 ( .A(b[413]), .B(n462), .Z(c[413]) );
  XOR U976 ( .A(n463), .B(n464), .Z(n460) );
  ANDN U977 ( .B(n465), .A(n466), .Z(n463) );
  XNOR U978 ( .A(b[412]), .B(n464), .Z(n465) );
  XNOR U979 ( .A(b[412]), .B(n466), .Z(c[412]) );
  XOR U980 ( .A(n467), .B(n468), .Z(n464) );
  ANDN U981 ( .B(n469), .A(n470), .Z(n467) );
  XNOR U982 ( .A(b[411]), .B(n468), .Z(n469) );
  XNOR U983 ( .A(b[411]), .B(n470), .Z(c[411]) );
  XOR U984 ( .A(n471), .B(n472), .Z(n468) );
  ANDN U985 ( .B(n473), .A(n474), .Z(n471) );
  XNOR U986 ( .A(b[410]), .B(n472), .Z(n473) );
  XNOR U987 ( .A(b[410]), .B(n474), .Z(c[410]) );
  XOR U988 ( .A(n475), .B(n476), .Z(n472) );
  ANDN U989 ( .B(n477), .A(n478), .Z(n475) );
  XNOR U990 ( .A(b[409]), .B(n476), .Z(n477) );
  XNOR U991 ( .A(b[40]), .B(n479), .Z(c[40]) );
  XNOR U992 ( .A(b[409]), .B(n478), .Z(c[409]) );
  XOR U993 ( .A(n480), .B(n481), .Z(n476) );
  ANDN U994 ( .B(n482), .A(n483), .Z(n480) );
  XNOR U995 ( .A(b[408]), .B(n481), .Z(n482) );
  XNOR U996 ( .A(b[408]), .B(n483), .Z(c[408]) );
  XOR U997 ( .A(n484), .B(n485), .Z(n481) );
  ANDN U998 ( .B(n486), .A(n487), .Z(n484) );
  XNOR U999 ( .A(b[407]), .B(n485), .Z(n486) );
  XNOR U1000 ( .A(b[407]), .B(n487), .Z(c[407]) );
  XOR U1001 ( .A(n488), .B(n489), .Z(n485) );
  ANDN U1002 ( .B(n490), .A(n491), .Z(n488) );
  XNOR U1003 ( .A(b[406]), .B(n489), .Z(n490) );
  XNOR U1004 ( .A(b[406]), .B(n491), .Z(c[406]) );
  XOR U1005 ( .A(n492), .B(n493), .Z(n489) );
  ANDN U1006 ( .B(n494), .A(n495), .Z(n492) );
  XNOR U1007 ( .A(b[405]), .B(n493), .Z(n494) );
  XNOR U1008 ( .A(b[405]), .B(n495), .Z(c[405]) );
  XOR U1009 ( .A(n496), .B(n497), .Z(n493) );
  ANDN U1010 ( .B(n498), .A(n499), .Z(n496) );
  XNOR U1011 ( .A(b[404]), .B(n497), .Z(n498) );
  XNOR U1012 ( .A(b[404]), .B(n499), .Z(c[404]) );
  XOR U1013 ( .A(n500), .B(n501), .Z(n497) );
  ANDN U1014 ( .B(n502), .A(n503), .Z(n500) );
  XNOR U1015 ( .A(b[403]), .B(n501), .Z(n502) );
  XNOR U1016 ( .A(b[403]), .B(n503), .Z(c[403]) );
  XOR U1017 ( .A(n504), .B(n505), .Z(n501) );
  ANDN U1018 ( .B(n506), .A(n507), .Z(n504) );
  XNOR U1019 ( .A(b[402]), .B(n505), .Z(n506) );
  XNOR U1020 ( .A(b[402]), .B(n507), .Z(c[402]) );
  XOR U1021 ( .A(n508), .B(n509), .Z(n505) );
  ANDN U1022 ( .B(n510), .A(n511), .Z(n508) );
  XNOR U1023 ( .A(b[401]), .B(n509), .Z(n510) );
  XNOR U1024 ( .A(b[401]), .B(n511), .Z(c[401]) );
  XOR U1025 ( .A(n512), .B(n513), .Z(n509) );
  ANDN U1026 ( .B(n514), .A(n515), .Z(n512) );
  XNOR U1027 ( .A(b[400]), .B(n513), .Z(n514) );
  XNOR U1028 ( .A(b[400]), .B(n515), .Z(c[400]) );
  XOR U1029 ( .A(n516), .B(n517), .Z(n513) );
  ANDN U1030 ( .B(n518), .A(n519), .Z(n516) );
  XNOR U1031 ( .A(b[399]), .B(n517), .Z(n518) );
  XNOR U1032 ( .A(b[3]), .B(n520), .Z(c[3]) );
  XNOR U1033 ( .A(b[39]), .B(n521), .Z(c[39]) );
  XNOR U1034 ( .A(b[399]), .B(n519), .Z(c[399]) );
  XOR U1035 ( .A(n522), .B(n523), .Z(n517) );
  ANDN U1036 ( .B(n524), .A(n525), .Z(n522) );
  XNOR U1037 ( .A(b[398]), .B(n523), .Z(n524) );
  XNOR U1038 ( .A(b[398]), .B(n525), .Z(c[398]) );
  XOR U1039 ( .A(n526), .B(n527), .Z(n523) );
  ANDN U1040 ( .B(n528), .A(n529), .Z(n526) );
  XNOR U1041 ( .A(b[397]), .B(n527), .Z(n528) );
  XNOR U1042 ( .A(b[397]), .B(n529), .Z(c[397]) );
  XOR U1043 ( .A(n530), .B(n531), .Z(n527) );
  ANDN U1044 ( .B(n532), .A(n533), .Z(n530) );
  XNOR U1045 ( .A(b[396]), .B(n531), .Z(n532) );
  XNOR U1046 ( .A(b[396]), .B(n533), .Z(c[396]) );
  XOR U1047 ( .A(n534), .B(n535), .Z(n531) );
  ANDN U1048 ( .B(n536), .A(n537), .Z(n534) );
  XNOR U1049 ( .A(b[395]), .B(n535), .Z(n536) );
  XNOR U1050 ( .A(b[395]), .B(n537), .Z(c[395]) );
  XOR U1051 ( .A(n538), .B(n539), .Z(n535) );
  ANDN U1052 ( .B(n540), .A(n541), .Z(n538) );
  XNOR U1053 ( .A(b[394]), .B(n539), .Z(n540) );
  XNOR U1054 ( .A(b[394]), .B(n541), .Z(c[394]) );
  XOR U1055 ( .A(n542), .B(n543), .Z(n539) );
  ANDN U1056 ( .B(n544), .A(n545), .Z(n542) );
  XNOR U1057 ( .A(b[393]), .B(n543), .Z(n544) );
  XNOR U1058 ( .A(b[393]), .B(n545), .Z(c[393]) );
  XOR U1059 ( .A(n546), .B(n547), .Z(n543) );
  ANDN U1060 ( .B(n548), .A(n549), .Z(n546) );
  XNOR U1061 ( .A(b[392]), .B(n547), .Z(n548) );
  XNOR U1062 ( .A(b[392]), .B(n549), .Z(c[392]) );
  XOR U1063 ( .A(n550), .B(n551), .Z(n547) );
  ANDN U1064 ( .B(n552), .A(n553), .Z(n550) );
  XNOR U1065 ( .A(b[391]), .B(n551), .Z(n552) );
  XNOR U1066 ( .A(b[391]), .B(n553), .Z(c[391]) );
  XOR U1067 ( .A(n554), .B(n555), .Z(n551) );
  ANDN U1068 ( .B(n556), .A(n557), .Z(n554) );
  XNOR U1069 ( .A(b[390]), .B(n555), .Z(n556) );
  XNOR U1070 ( .A(b[390]), .B(n557), .Z(c[390]) );
  XOR U1071 ( .A(n558), .B(n559), .Z(n555) );
  ANDN U1072 ( .B(n560), .A(n561), .Z(n558) );
  XNOR U1073 ( .A(b[389]), .B(n559), .Z(n560) );
  XNOR U1074 ( .A(b[38]), .B(n562), .Z(c[38]) );
  XNOR U1075 ( .A(b[389]), .B(n561), .Z(c[389]) );
  XOR U1076 ( .A(n563), .B(n564), .Z(n559) );
  ANDN U1077 ( .B(n565), .A(n566), .Z(n563) );
  XNOR U1078 ( .A(b[388]), .B(n564), .Z(n565) );
  XNOR U1079 ( .A(b[388]), .B(n566), .Z(c[388]) );
  XOR U1080 ( .A(n567), .B(n568), .Z(n564) );
  ANDN U1081 ( .B(n569), .A(n570), .Z(n567) );
  XNOR U1082 ( .A(b[387]), .B(n568), .Z(n569) );
  XNOR U1083 ( .A(b[387]), .B(n570), .Z(c[387]) );
  XOR U1084 ( .A(n571), .B(n572), .Z(n568) );
  ANDN U1085 ( .B(n573), .A(n574), .Z(n571) );
  XNOR U1086 ( .A(b[386]), .B(n572), .Z(n573) );
  XNOR U1087 ( .A(b[386]), .B(n574), .Z(c[386]) );
  XOR U1088 ( .A(n575), .B(n576), .Z(n572) );
  ANDN U1089 ( .B(n577), .A(n578), .Z(n575) );
  XNOR U1090 ( .A(b[385]), .B(n576), .Z(n577) );
  XNOR U1091 ( .A(b[385]), .B(n578), .Z(c[385]) );
  XOR U1092 ( .A(n579), .B(n580), .Z(n576) );
  ANDN U1093 ( .B(n581), .A(n582), .Z(n579) );
  XNOR U1094 ( .A(b[384]), .B(n580), .Z(n581) );
  XNOR U1095 ( .A(b[384]), .B(n582), .Z(c[384]) );
  XOR U1096 ( .A(n583), .B(n584), .Z(n580) );
  ANDN U1097 ( .B(n585), .A(n586), .Z(n583) );
  XNOR U1098 ( .A(b[383]), .B(n584), .Z(n585) );
  XNOR U1099 ( .A(b[383]), .B(n586), .Z(c[383]) );
  XOR U1100 ( .A(n587), .B(n588), .Z(n584) );
  ANDN U1101 ( .B(n589), .A(n590), .Z(n587) );
  XNOR U1102 ( .A(b[382]), .B(n588), .Z(n589) );
  XNOR U1103 ( .A(b[382]), .B(n590), .Z(c[382]) );
  XOR U1104 ( .A(n591), .B(n592), .Z(n588) );
  ANDN U1105 ( .B(n593), .A(n594), .Z(n591) );
  XNOR U1106 ( .A(b[381]), .B(n592), .Z(n593) );
  XNOR U1107 ( .A(b[381]), .B(n594), .Z(c[381]) );
  XOR U1108 ( .A(n595), .B(n596), .Z(n592) );
  ANDN U1109 ( .B(n597), .A(n598), .Z(n595) );
  XNOR U1110 ( .A(b[380]), .B(n596), .Z(n597) );
  XNOR U1111 ( .A(b[380]), .B(n598), .Z(c[380]) );
  XOR U1112 ( .A(n599), .B(n600), .Z(n596) );
  ANDN U1113 ( .B(n601), .A(n602), .Z(n599) );
  XNOR U1114 ( .A(b[379]), .B(n600), .Z(n601) );
  XNOR U1115 ( .A(b[37]), .B(n603), .Z(c[37]) );
  XNOR U1116 ( .A(b[379]), .B(n602), .Z(c[379]) );
  XOR U1117 ( .A(n604), .B(n605), .Z(n600) );
  ANDN U1118 ( .B(n606), .A(n607), .Z(n604) );
  XNOR U1119 ( .A(b[378]), .B(n605), .Z(n606) );
  XNOR U1120 ( .A(b[378]), .B(n607), .Z(c[378]) );
  XOR U1121 ( .A(n608), .B(n609), .Z(n605) );
  ANDN U1122 ( .B(n610), .A(n611), .Z(n608) );
  XNOR U1123 ( .A(b[377]), .B(n609), .Z(n610) );
  XNOR U1124 ( .A(b[377]), .B(n611), .Z(c[377]) );
  XOR U1125 ( .A(n612), .B(n613), .Z(n609) );
  ANDN U1126 ( .B(n614), .A(n615), .Z(n612) );
  XNOR U1127 ( .A(b[376]), .B(n613), .Z(n614) );
  XNOR U1128 ( .A(b[376]), .B(n615), .Z(c[376]) );
  XOR U1129 ( .A(n616), .B(n617), .Z(n613) );
  ANDN U1130 ( .B(n618), .A(n619), .Z(n616) );
  XNOR U1131 ( .A(b[375]), .B(n617), .Z(n618) );
  XNOR U1132 ( .A(b[375]), .B(n619), .Z(c[375]) );
  XOR U1133 ( .A(n620), .B(n621), .Z(n617) );
  ANDN U1134 ( .B(n622), .A(n623), .Z(n620) );
  XNOR U1135 ( .A(b[374]), .B(n621), .Z(n622) );
  XNOR U1136 ( .A(b[374]), .B(n623), .Z(c[374]) );
  XOR U1137 ( .A(n624), .B(n625), .Z(n621) );
  ANDN U1138 ( .B(n626), .A(n627), .Z(n624) );
  XNOR U1139 ( .A(b[373]), .B(n625), .Z(n626) );
  XNOR U1140 ( .A(b[373]), .B(n627), .Z(c[373]) );
  XOR U1141 ( .A(n628), .B(n629), .Z(n625) );
  ANDN U1142 ( .B(n630), .A(n631), .Z(n628) );
  XNOR U1143 ( .A(b[372]), .B(n629), .Z(n630) );
  XNOR U1144 ( .A(b[372]), .B(n631), .Z(c[372]) );
  XOR U1145 ( .A(n632), .B(n633), .Z(n629) );
  ANDN U1146 ( .B(n634), .A(n635), .Z(n632) );
  XNOR U1147 ( .A(b[371]), .B(n633), .Z(n634) );
  XNOR U1148 ( .A(b[371]), .B(n635), .Z(c[371]) );
  XOR U1149 ( .A(n636), .B(n637), .Z(n633) );
  ANDN U1150 ( .B(n638), .A(n639), .Z(n636) );
  XNOR U1151 ( .A(b[370]), .B(n637), .Z(n638) );
  XNOR U1152 ( .A(b[370]), .B(n639), .Z(c[370]) );
  XOR U1153 ( .A(n640), .B(n641), .Z(n637) );
  ANDN U1154 ( .B(n642), .A(n643), .Z(n640) );
  XNOR U1155 ( .A(b[369]), .B(n641), .Z(n642) );
  XNOR U1156 ( .A(b[36]), .B(n644), .Z(c[36]) );
  XNOR U1157 ( .A(b[369]), .B(n643), .Z(c[369]) );
  XOR U1158 ( .A(n645), .B(n646), .Z(n641) );
  ANDN U1159 ( .B(n647), .A(n648), .Z(n645) );
  XNOR U1160 ( .A(b[368]), .B(n646), .Z(n647) );
  XNOR U1161 ( .A(b[368]), .B(n648), .Z(c[368]) );
  XOR U1162 ( .A(n649), .B(n650), .Z(n646) );
  ANDN U1163 ( .B(n651), .A(n652), .Z(n649) );
  XNOR U1164 ( .A(b[367]), .B(n650), .Z(n651) );
  XNOR U1165 ( .A(b[367]), .B(n652), .Z(c[367]) );
  XOR U1166 ( .A(n653), .B(n654), .Z(n650) );
  ANDN U1167 ( .B(n655), .A(n656), .Z(n653) );
  XNOR U1168 ( .A(b[366]), .B(n654), .Z(n655) );
  XNOR U1169 ( .A(b[366]), .B(n656), .Z(c[366]) );
  XOR U1170 ( .A(n657), .B(n658), .Z(n654) );
  ANDN U1171 ( .B(n659), .A(n660), .Z(n657) );
  XNOR U1172 ( .A(b[365]), .B(n658), .Z(n659) );
  XNOR U1173 ( .A(b[365]), .B(n660), .Z(c[365]) );
  XOR U1174 ( .A(n661), .B(n662), .Z(n658) );
  ANDN U1175 ( .B(n663), .A(n664), .Z(n661) );
  XNOR U1176 ( .A(b[364]), .B(n662), .Z(n663) );
  XNOR U1177 ( .A(b[364]), .B(n664), .Z(c[364]) );
  XOR U1178 ( .A(n665), .B(n666), .Z(n662) );
  ANDN U1179 ( .B(n667), .A(n668), .Z(n665) );
  XNOR U1180 ( .A(b[363]), .B(n666), .Z(n667) );
  XNOR U1181 ( .A(b[363]), .B(n668), .Z(c[363]) );
  XOR U1182 ( .A(n669), .B(n670), .Z(n666) );
  ANDN U1183 ( .B(n671), .A(n672), .Z(n669) );
  XNOR U1184 ( .A(b[362]), .B(n670), .Z(n671) );
  XNOR U1185 ( .A(b[362]), .B(n672), .Z(c[362]) );
  XOR U1186 ( .A(n673), .B(n674), .Z(n670) );
  ANDN U1187 ( .B(n675), .A(n676), .Z(n673) );
  XNOR U1188 ( .A(b[361]), .B(n674), .Z(n675) );
  XNOR U1189 ( .A(b[361]), .B(n676), .Z(c[361]) );
  XOR U1190 ( .A(n677), .B(n678), .Z(n674) );
  ANDN U1191 ( .B(n679), .A(n680), .Z(n677) );
  XNOR U1192 ( .A(b[360]), .B(n678), .Z(n679) );
  XNOR U1193 ( .A(b[360]), .B(n680), .Z(c[360]) );
  XOR U1194 ( .A(n681), .B(n682), .Z(n678) );
  ANDN U1195 ( .B(n683), .A(n684), .Z(n681) );
  XNOR U1196 ( .A(b[359]), .B(n682), .Z(n683) );
  XNOR U1197 ( .A(b[35]), .B(n685), .Z(c[35]) );
  XNOR U1198 ( .A(b[359]), .B(n684), .Z(c[359]) );
  XOR U1199 ( .A(n686), .B(n687), .Z(n682) );
  ANDN U1200 ( .B(n688), .A(n689), .Z(n686) );
  XNOR U1201 ( .A(b[358]), .B(n687), .Z(n688) );
  XNOR U1202 ( .A(b[358]), .B(n689), .Z(c[358]) );
  XOR U1203 ( .A(n690), .B(n691), .Z(n687) );
  ANDN U1204 ( .B(n692), .A(n693), .Z(n690) );
  XNOR U1205 ( .A(b[357]), .B(n691), .Z(n692) );
  XNOR U1206 ( .A(b[357]), .B(n693), .Z(c[357]) );
  XOR U1207 ( .A(n694), .B(n695), .Z(n691) );
  ANDN U1208 ( .B(n696), .A(n697), .Z(n694) );
  XNOR U1209 ( .A(b[356]), .B(n695), .Z(n696) );
  XNOR U1210 ( .A(b[356]), .B(n697), .Z(c[356]) );
  XOR U1211 ( .A(n698), .B(n699), .Z(n695) );
  ANDN U1212 ( .B(n700), .A(n701), .Z(n698) );
  XNOR U1213 ( .A(b[355]), .B(n699), .Z(n700) );
  XNOR U1214 ( .A(b[355]), .B(n701), .Z(c[355]) );
  XOR U1215 ( .A(n702), .B(n703), .Z(n699) );
  ANDN U1216 ( .B(n704), .A(n705), .Z(n702) );
  XNOR U1217 ( .A(b[354]), .B(n703), .Z(n704) );
  XNOR U1218 ( .A(b[354]), .B(n705), .Z(c[354]) );
  XOR U1219 ( .A(n706), .B(n707), .Z(n703) );
  ANDN U1220 ( .B(n708), .A(n709), .Z(n706) );
  XNOR U1221 ( .A(b[353]), .B(n707), .Z(n708) );
  XNOR U1222 ( .A(b[353]), .B(n709), .Z(c[353]) );
  XOR U1223 ( .A(n710), .B(n711), .Z(n707) );
  ANDN U1224 ( .B(n712), .A(n713), .Z(n710) );
  XNOR U1225 ( .A(b[352]), .B(n711), .Z(n712) );
  XNOR U1226 ( .A(b[352]), .B(n713), .Z(c[352]) );
  XOR U1227 ( .A(n714), .B(n715), .Z(n711) );
  ANDN U1228 ( .B(n716), .A(n717), .Z(n714) );
  XNOR U1229 ( .A(b[351]), .B(n715), .Z(n716) );
  XNOR U1230 ( .A(b[351]), .B(n717), .Z(c[351]) );
  XOR U1231 ( .A(n718), .B(n719), .Z(n715) );
  ANDN U1232 ( .B(n720), .A(n721), .Z(n718) );
  XNOR U1233 ( .A(b[350]), .B(n719), .Z(n720) );
  XNOR U1234 ( .A(b[350]), .B(n721), .Z(c[350]) );
  XOR U1235 ( .A(n722), .B(n723), .Z(n719) );
  ANDN U1236 ( .B(n724), .A(n725), .Z(n722) );
  XNOR U1237 ( .A(b[349]), .B(n723), .Z(n724) );
  XNOR U1238 ( .A(b[34]), .B(n726), .Z(c[34]) );
  XNOR U1239 ( .A(b[349]), .B(n725), .Z(c[349]) );
  XOR U1240 ( .A(n727), .B(n728), .Z(n723) );
  ANDN U1241 ( .B(n729), .A(n730), .Z(n727) );
  XNOR U1242 ( .A(b[348]), .B(n728), .Z(n729) );
  XNOR U1243 ( .A(b[348]), .B(n730), .Z(c[348]) );
  XOR U1244 ( .A(n731), .B(n732), .Z(n728) );
  ANDN U1245 ( .B(n733), .A(n734), .Z(n731) );
  XNOR U1246 ( .A(b[347]), .B(n732), .Z(n733) );
  XNOR U1247 ( .A(b[347]), .B(n734), .Z(c[347]) );
  XOR U1248 ( .A(n735), .B(n736), .Z(n732) );
  ANDN U1249 ( .B(n737), .A(n738), .Z(n735) );
  XNOR U1250 ( .A(b[346]), .B(n736), .Z(n737) );
  XNOR U1251 ( .A(b[346]), .B(n738), .Z(c[346]) );
  XOR U1252 ( .A(n739), .B(n740), .Z(n736) );
  ANDN U1253 ( .B(n741), .A(n742), .Z(n739) );
  XNOR U1254 ( .A(b[345]), .B(n740), .Z(n741) );
  XNOR U1255 ( .A(b[345]), .B(n742), .Z(c[345]) );
  XOR U1256 ( .A(n743), .B(n744), .Z(n740) );
  ANDN U1257 ( .B(n745), .A(n746), .Z(n743) );
  XNOR U1258 ( .A(b[344]), .B(n744), .Z(n745) );
  XNOR U1259 ( .A(b[344]), .B(n746), .Z(c[344]) );
  XOR U1260 ( .A(n747), .B(n748), .Z(n744) );
  ANDN U1261 ( .B(n749), .A(n750), .Z(n747) );
  XNOR U1262 ( .A(b[343]), .B(n748), .Z(n749) );
  XNOR U1263 ( .A(b[343]), .B(n750), .Z(c[343]) );
  XOR U1264 ( .A(n751), .B(n752), .Z(n748) );
  ANDN U1265 ( .B(n753), .A(n754), .Z(n751) );
  XNOR U1266 ( .A(b[342]), .B(n752), .Z(n753) );
  XNOR U1267 ( .A(b[342]), .B(n754), .Z(c[342]) );
  XOR U1268 ( .A(n755), .B(n756), .Z(n752) );
  ANDN U1269 ( .B(n757), .A(n758), .Z(n755) );
  XNOR U1270 ( .A(b[341]), .B(n756), .Z(n757) );
  XNOR U1271 ( .A(b[341]), .B(n758), .Z(c[341]) );
  XOR U1272 ( .A(n759), .B(n760), .Z(n756) );
  ANDN U1273 ( .B(n761), .A(n762), .Z(n759) );
  XNOR U1274 ( .A(b[340]), .B(n760), .Z(n761) );
  XNOR U1275 ( .A(b[340]), .B(n762), .Z(c[340]) );
  XOR U1276 ( .A(n763), .B(n764), .Z(n760) );
  ANDN U1277 ( .B(n765), .A(n766), .Z(n763) );
  XNOR U1278 ( .A(b[339]), .B(n764), .Z(n765) );
  XNOR U1279 ( .A(b[33]), .B(n767), .Z(c[33]) );
  XNOR U1280 ( .A(b[339]), .B(n766), .Z(c[339]) );
  XOR U1281 ( .A(n768), .B(n769), .Z(n764) );
  ANDN U1282 ( .B(n770), .A(n771), .Z(n768) );
  XNOR U1283 ( .A(b[338]), .B(n769), .Z(n770) );
  XNOR U1284 ( .A(b[338]), .B(n771), .Z(c[338]) );
  XOR U1285 ( .A(n772), .B(n773), .Z(n769) );
  ANDN U1286 ( .B(n774), .A(n775), .Z(n772) );
  XNOR U1287 ( .A(b[337]), .B(n773), .Z(n774) );
  XNOR U1288 ( .A(b[337]), .B(n775), .Z(c[337]) );
  XOR U1289 ( .A(n776), .B(n777), .Z(n773) );
  ANDN U1290 ( .B(n778), .A(n779), .Z(n776) );
  XNOR U1291 ( .A(b[336]), .B(n777), .Z(n778) );
  XNOR U1292 ( .A(b[336]), .B(n779), .Z(c[336]) );
  XOR U1293 ( .A(n780), .B(n781), .Z(n777) );
  ANDN U1294 ( .B(n782), .A(n783), .Z(n780) );
  XNOR U1295 ( .A(b[335]), .B(n781), .Z(n782) );
  XNOR U1296 ( .A(b[335]), .B(n783), .Z(c[335]) );
  XOR U1297 ( .A(n784), .B(n785), .Z(n781) );
  ANDN U1298 ( .B(n786), .A(n787), .Z(n784) );
  XNOR U1299 ( .A(b[334]), .B(n785), .Z(n786) );
  XNOR U1300 ( .A(b[334]), .B(n787), .Z(c[334]) );
  XOR U1301 ( .A(n788), .B(n789), .Z(n785) );
  ANDN U1302 ( .B(n790), .A(n791), .Z(n788) );
  XNOR U1303 ( .A(b[333]), .B(n789), .Z(n790) );
  XNOR U1304 ( .A(b[333]), .B(n791), .Z(c[333]) );
  XOR U1305 ( .A(n792), .B(n793), .Z(n789) );
  ANDN U1306 ( .B(n794), .A(n795), .Z(n792) );
  XNOR U1307 ( .A(b[332]), .B(n793), .Z(n794) );
  XNOR U1308 ( .A(b[332]), .B(n795), .Z(c[332]) );
  XOR U1309 ( .A(n796), .B(n797), .Z(n793) );
  ANDN U1310 ( .B(n798), .A(n799), .Z(n796) );
  XNOR U1311 ( .A(b[331]), .B(n797), .Z(n798) );
  XNOR U1312 ( .A(b[331]), .B(n799), .Z(c[331]) );
  XOR U1313 ( .A(n800), .B(n801), .Z(n797) );
  ANDN U1314 ( .B(n802), .A(n803), .Z(n800) );
  XNOR U1315 ( .A(b[330]), .B(n801), .Z(n802) );
  XNOR U1316 ( .A(b[330]), .B(n803), .Z(c[330]) );
  XOR U1317 ( .A(n804), .B(n805), .Z(n801) );
  ANDN U1318 ( .B(n806), .A(n807), .Z(n804) );
  XNOR U1319 ( .A(b[329]), .B(n805), .Z(n806) );
  XNOR U1320 ( .A(b[32]), .B(n808), .Z(c[32]) );
  XNOR U1321 ( .A(b[329]), .B(n807), .Z(c[329]) );
  XOR U1322 ( .A(n809), .B(n810), .Z(n805) );
  ANDN U1323 ( .B(n811), .A(n812), .Z(n809) );
  XNOR U1324 ( .A(b[328]), .B(n810), .Z(n811) );
  XNOR U1325 ( .A(b[328]), .B(n812), .Z(c[328]) );
  XOR U1326 ( .A(n813), .B(n814), .Z(n810) );
  ANDN U1327 ( .B(n815), .A(n816), .Z(n813) );
  XNOR U1328 ( .A(b[327]), .B(n814), .Z(n815) );
  XNOR U1329 ( .A(b[327]), .B(n816), .Z(c[327]) );
  XOR U1330 ( .A(n817), .B(n818), .Z(n814) );
  ANDN U1331 ( .B(n819), .A(n820), .Z(n817) );
  XNOR U1332 ( .A(b[326]), .B(n818), .Z(n819) );
  XNOR U1333 ( .A(b[326]), .B(n820), .Z(c[326]) );
  XOR U1334 ( .A(n821), .B(n822), .Z(n818) );
  ANDN U1335 ( .B(n823), .A(n824), .Z(n821) );
  XNOR U1336 ( .A(b[325]), .B(n822), .Z(n823) );
  XNOR U1337 ( .A(b[325]), .B(n824), .Z(c[325]) );
  XOR U1338 ( .A(n825), .B(n826), .Z(n822) );
  ANDN U1339 ( .B(n827), .A(n828), .Z(n825) );
  XNOR U1340 ( .A(b[324]), .B(n826), .Z(n827) );
  XNOR U1341 ( .A(b[324]), .B(n828), .Z(c[324]) );
  XOR U1342 ( .A(n829), .B(n830), .Z(n826) );
  ANDN U1343 ( .B(n831), .A(n832), .Z(n829) );
  XNOR U1344 ( .A(b[323]), .B(n830), .Z(n831) );
  XNOR U1345 ( .A(b[323]), .B(n832), .Z(c[323]) );
  XOR U1346 ( .A(n833), .B(n834), .Z(n830) );
  ANDN U1347 ( .B(n835), .A(n836), .Z(n833) );
  XNOR U1348 ( .A(b[322]), .B(n834), .Z(n835) );
  XNOR U1349 ( .A(b[322]), .B(n836), .Z(c[322]) );
  XOR U1350 ( .A(n837), .B(n838), .Z(n834) );
  ANDN U1351 ( .B(n839), .A(n840), .Z(n837) );
  XNOR U1352 ( .A(b[321]), .B(n838), .Z(n839) );
  XNOR U1353 ( .A(b[321]), .B(n840), .Z(c[321]) );
  XOR U1354 ( .A(n841), .B(n842), .Z(n838) );
  ANDN U1355 ( .B(n843), .A(n844), .Z(n841) );
  XNOR U1356 ( .A(b[320]), .B(n842), .Z(n843) );
  XNOR U1357 ( .A(b[320]), .B(n844), .Z(c[320]) );
  XOR U1358 ( .A(n845), .B(n846), .Z(n842) );
  ANDN U1359 ( .B(n847), .A(n848), .Z(n845) );
  XNOR U1360 ( .A(b[319]), .B(n846), .Z(n847) );
  XNOR U1361 ( .A(b[31]), .B(n849), .Z(c[31]) );
  XNOR U1362 ( .A(b[319]), .B(n848), .Z(c[319]) );
  XOR U1363 ( .A(n850), .B(n851), .Z(n846) );
  ANDN U1364 ( .B(n852), .A(n853), .Z(n850) );
  XNOR U1365 ( .A(b[318]), .B(n851), .Z(n852) );
  XNOR U1366 ( .A(b[318]), .B(n853), .Z(c[318]) );
  XOR U1367 ( .A(n854), .B(n855), .Z(n851) );
  ANDN U1368 ( .B(n856), .A(n857), .Z(n854) );
  XNOR U1369 ( .A(b[317]), .B(n855), .Z(n856) );
  XNOR U1370 ( .A(b[317]), .B(n857), .Z(c[317]) );
  XOR U1371 ( .A(n858), .B(n859), .Z(n855) );
  ANDN U1372 ( .B(n860), .A(n861), .Z(n858) );
  XNOR U1373 ( .A(b[316]), .B(n859), .Z(n860) );
  XNOR U1374 ( .A(b[316]), .B(n861), .Z(c[316]) );
  XOR U1375 ( .A(n862), .B(n863), .Z(n859) );
  ANDN U1376 ( .B(n864), .A(n865), .Z(n862) );
  XNOR U1377 ( .A(b[315]), .B(n863), .Z(n864) );
  XNOR U1378 ( .A(b[315]), .B(n865), .Z(c[315]) );
  XOR U1379 ( .A(n866), .B(n867), .Z(n863) );
  ANDN U1380 ( .B(n868), .A(n869), .Z(n866) );
  XNOR U1381 ( .A(b[314]), .B(n867), .Z(n868) );
  XNOR U1382 ( .A(b[314]), .B(n869), .Z(c[314]) );
  XOR U1383 ( .A(n870), .B(n871), .Z(n867) );
  ANDN U1384 ( .B(n872), .A(n873), .Z(n870) );
  XNOR U1385 ( .A(b[313]), .B(n871), .Z(n872) );
  XNOR U1386 ( .A(b[313]), .B(n873), .Z(c[313]) );
  XOR U1387 ( .A(n874), .B(n875), .Z(n871) );
  ANDN U1388 ( .B(n876), .A(n877), .Z(n874) );
  XNOR U1389 ( .A(b[312]), .B(n875), .Z(n876) );
  XNOR U1390 ( .A(b[312]), .B(n877), .Z(c[312]) );
  XOR U1391 ( .A(n878), .B(n879), .Z(n875) );
  ANDN U1392 ( .B(n880), .A(n881), .Z(n878) );
  XNOR U1393 ( .A(b[311]), .B(n879), .Z(n880) );
  XNOR U1394 ( .A(b[311]), .B(n881), .Z(c[311]) );
  XOR U1395 ( .A(n882), .B(n883), .Z(n879) );
  ANDN U1396 ( .B(n884), .A(n885), .Z(n882) );
  XNOR U1397 ( .A(b[310]), .B(n883), .Z(n884) );
  XNOR U1398 ( .A(b[310]), .B(n885), .Z(c[310]) );
  XOR U1399 ( .A(n886), .B(n887), .Z(n883) );
  ANDN U1400 ( .B(n888), .A(n889), .Z(n886) );
  XNOR U1401 ( .A(b[309]), .B(n887), .Z(n888) );
  XNOR U1402 ( .A(b[30]), .B(n890), .Z(c[30]) );
  XNOR U1403 ( .A(b[309]), .B(n889), .Z(c[309]) );
  XOR U1404 ( .A(n891), .B(n892), .Z(n887) );
  ANDN U1405 ( .B(n893), .A(n894), .Z(n891) );
  XNOR U1406 ( .A(b[308]), .B(n892), .Z(n893) );
  XNOR U1407 ( .A(b[308]), .B(n894), .Z(c[308]) );
  XOR U1408 ( .A(n895), .B(n896), .Z(n892) );
  ANDN U1409 ( .B(n897), .A(n898), .Z(n895) );
  XNOR U1410 ( .A(b[307]), .B(n896), .Z(n897) );
  XNOR U1411 ( .A(b[307]), .B(n898), .Z(c[307]) );
  XOR U1412 ( .A(n899), .B(n900), .Z(n896) );
  ANDN U1413 ( .B(n901), .A(n902), .Z(n899) );
  XNOR U1414 ( .A(b[306]), .B(n900), .Z(n901) );
  XNOR U1415 ( .A(b[306]), .B(n902), .Z(c[306]) );
  XOR U1416 ( .A(n903), .B(n904), .Z(n900) );
  ANDN U1417 ( .B(n905), .A(n906), .Z(n903) );
  XNOR U1418 ( .A(b[305]), .B(n904), .Z(n905) );
  XNOR U1419 ( .A(b[305]), .B(n906), .Z(c[305]) );
  XOR U1420 ( .A(n907), .B(n908), .Z(n904) );
  ANDN U1421 ( .B(n909), .A(n910), .Z(n907) );
  XNOR U1422 ( .A(b[304]), .B(n908), .Z(n909) );
  XNOR U1423 ( .A(b[304]), .B(n910), .Z(c[304]) );
  XOR U1424 ( .A(n911), .B(n912), .Z(n908) );
  ANDN U1425 ( .B(n913), .A(n914), .Z(n911) );
  XNOR U1426 ( .A(b[303]), .B(n912), .Z(n913) );
  XNOR U1427 ( .A(b[303]), .B(n914), .Z(c[303]) );
  XOR U1428 ( .A(n915), .B(n916), .Z(n912) );
  ANDN U1429 ( .B(n917), .A(n918), .Z(n915) );
  XNOR U1430 ( .A(b[302]), .B(n916), .Z(n917) );
  XNOR U1431 ( .A(b[302]), .B(n918), .Z(c[302]) );
  XOR U1432 ( .A(n919), .B(n920), .Z(n916) );
  ANDN U1433 ( .B(n921), .A(n922), .Z(n919) );
  XNOR U1434 ( .A(b[301]), .B(n920), .Z(n921) );
  XNOR U1435 ( .A(b[301]), .B(n922), .Z(c[301]) );
  XOR U1436 ( .A(n923), .B(n924), .Z(n920) );
  ANDN U1437 ( .B(n925), .A(n926), .Z(n923) );
  XNOR U1438 ( .A(b[300]), .B(n924), .Z(n925) );
  XNOR U1439 ( .A(b[300]), .B(n926), .Z(c[300]) );
  XOR U1440 ( .A(n927), .B(n928), .Z(n924) );
  ANDN U1441 ( .B(n929), .A(n930), .Z(n927) );
  XNOR U1442 ( .A(b[299]), .B(n928), .Z(n929) );
  XNOR U1443 ( .A(b[2]), .B(n931), .Z(c[2]) );
  XNOR U1444 ( .A(b[29]), .B(n932), .Z(c[29]) );
  XNOR U1445 ( .A(b[299]), .B(n930), .Z(c[299]) );
  XOR U1446 ( .A(n933), .B(n934), .Z(n928) );
  ANDN U1447 ( .B(n935), .A(n936), .Z(n933) );
  XNOR U1448 ( .A(b[298]), .B(n934), .Z(n935) );
  XNOR U1449 ( .A(b[298]), .B(n936), .Z(c[298]) );
  XOR U1450 ( .A(n937), .B(n938), .Z(n934) );
  ANDN U1451 ( .B(n939), .A(n940), .Z(n937) );
  XNOR U1452 ( .A(b[297]), .B(n938), .Z(n939) );
  XNOR U1453 ( .A(b[297]), .B(n940), .Z(c[297]) );
  XOR U1454 ( .A(n941), .B(n942), .Z(n938) );
  ANDN U1455 ( .B(n943), .A(n944), .Z(n941) );
  XNOR U1456 ( .A(b[296]), .B(n942), .Z(n943) );
  XNOR U1457 ( .A(b[296]), .B(n944), .Z(c[296]) );
  XOR U1458 ( .A(n945), .B(n946), .Z(n942) );
  ANDN U1459 ( .B(n947), .A(n948), .Z(n945) );
  XNOR U1460 ( .A(b[295]), .B(n946), .Z(n947) );
  XNOR U1461 ( .A(b[295]), .B(n948), .Z(c[295]) );
  XOR U1462 ( .A(n949), .B(n950), .Z(n946) );
  ANDN U1463 ( .B(n951), .A(n952), .Z(n949) );
  XNOR U1464 ( .A(b[294]), .B(n950), .Z(n951) );
  XNOR U1465 ( .A(b[294]), .B(n952), .Z(c[294]) );
  XOR U1466 ( .A(n953), .B(n954), .Z(n950) );
  ANDN U1467 ( .B(n955), .A(n956), .Z(n953) );
  XNOR U1468 ( .A(b[293]), .B(n954), .Z(n955) );
  XNOR U1469 ( .A(b[293]), .B(n956), .Z(c[293]) );
  XOR U1470 ( .A(n957), .B(n958), .Z(n954) );
  ANDN U1471 ( .B(n959), .A(n960), .Z(n957) );
  XNOR U1472 ( .A(b[292]), .B(n958), .Z(n959) );
  XNOR U1473 ( .A(b[292]), .B(n960), .Z(c[292]) );
  XOR U1474 ( .A(n961), .B(n962), .Z(n958) );
  ANDN U1475 ( .B(n963), .A(n964), .Z(n961) );
  XNOR U1476 ( .A(b[291]), .B(n962), .Z(n963) );
  XNOR U1477 ( .A(b[291]), .B(n964), .Z(c[291]) );
  XOR U1478 ( .A(n965), .B(n966), .Z(n962) );
  ANDN U1479 ( .B(n967), .A(n968), .Z(n965) );
  XNOR U1480 ( .A(b[290]), .B(n966), .Z(n967) );
  XNOR U1481 ( .A(b[290]), .B(n968), .Z(c[290]) );
  XOR U1482 ( .A(n969), .B(n970), .Z(n966) );
  ANDN U1483 ( .B(n971), .A(n972), .Z(n969) );
  XNOR U1484 ( .A(b[289]), .B(n970), .Z(n971) );
  XNOR U1485 ( .A(b[28]), .B(n973), .Z(c[28]) );
  XNOR U1486 ( .A(b[289]), .B(n972), .Z(c[289]) );
  XOR U1487 ( .A(n974), .B(n975), .Z(n970) );
  ANDN U1488 ( .B(n976), .A(n977), .Z(n974) );
  XNOR U1489 ( .A(b[288]), .B(n975), .Z(n976) );
  XNOR U1490 ( .A(b[288]), .B(n977), .Z(c[288]) );
  XOR U1491 ( .A(n978), .B(n979), .Z(n975) );
  ANDN U1492 ( .B(n980), .A(n981), .Z(n978) );
  XNOR U1493 ( .A(b[287]), .B(n979), .Z(n980) );
  XNOR U1494 ( .A(b[287]), .B(n981), .Z(c[287]) );
  XOR U1495 ( .A(n982), .B(n983), .Z(n979) );
  ANDN U1496 ( .B(n984), .A(n985), .Z(n982) );
  XNOR U1497 ( .A(b[286]), .B(n983), .Z(n984) );
  XNOR U1498 ( .A(b[286]), .B(n985), .Z(c[286]) );
  XOR U1499 ( .A(n986), .B(n987), .Z(n983) );
  ANDN U1500 ( .B(n988), .A(n989), .Z(n986) );
  XNOR U1501 ( .A(b[285]), .B(n987), .Z(n988) );
  XNOR U1502 ( .A(b[285]), .B(n989), .Z(c[285]) );
  XOR U1503 ( .A(n990), .B(n991), .Z(n987) );
  ANDN U1504 ( .B(n992), .A(n993), .Z(n990) );
  XNOR U1505 ( .A(b[284]), .B(n991), .Z(n992) );
  XNOR U1506 ( .A(b[284]), .B(n993), .Z(c[284]) );
  XOR U1507 ( .A(n994), .B(n995), .Z(n991) );
  ANDN U1508 ( .B(n996), .A(n997), .Z(n994) );
  XNOR U1509 ( .A(b[283]), .B(n995), .Z(n996) );
  XNOR U1510 ( .A(b[283]), .B(n997), .Z(c[283]) );
  XOR U1511 ( .A(n998), .B(n999), .Z(n995) );
  ANDN U1512 ( .B(n1000), .A(n1001), .Z(n998) );
  XNOR U1513 ( .A(b[282]), .B(n999), .Z(n1000) );
  XNOR U1514 ( .A(b[282]), .B(n1001), .Z(c[282]) );
  XOR U1515 ( .A(n1002), .B(n1003), .Z(n999) );
  ANDN U1516 ( .B(n1004), .A(n1005), .Z(n1002) );
  XNOR U1517 ( .A(b[281]), .B(n1003), .Z(n1004) );
  XNOR U1518 ( .A(b[281]), .B(n1005), .Z(c[281]) );
  XOR U1519 ( .A(n1006), .B(n1007), .Z(n1003) );
  ANDN U1520 ( .B(n1008), .A(n1009), .Z(n1006) );
  XNOR U1521 ( .A(b[280]), .B(n1007), .Z(n1008) );
  XNOR U1522 ( .A(b[280]), .B(n1009), .Z(c[280]) );
  XOR U1523 ( .A(n1010), .B(n1011), .Z(n1007) );
  ANDN U1524 ( .B(n1012), .A(n1013), .Z(n1010) );
  XNOR U1525 ( .A(b[279]), .B(n1011), .Z(n1012) );
  XNOR U1526 ( .A(b[27]), .B(n1014), .Z(c[27]) );
  XNOR U1527 ( .A(b[279]), .B(n1013), .Z(c[279]) );
  XOR U1528 ( .A(n1015), .B(n1016), .Z(n1011) );
  ANDN U1529 ( .B(n1017), .A(n1018), .Z(n1015) );
  XNOR U1530 ( .A(b[278]), .B(n1016), .Z(n1017) );
  XNOR U1531 ( .A(b[278]), .B(n1018), .Z(c[278]) );
  XOR U1532 ( .A(n1019), .B(n1020), .Z(n1016) );
  ANDN U1533 ( .B(n1021), .A(n1022), .Z(n1019) );
  XNOR U1534 ( .A(b[277]), .B(n1020), .Z(n1021) );
  XNOR U1535 ( .A(b[277]), .B(n1022), .Z(c[277]) );
  XOR U1536 ( .A(n1023), .B(n1024), .Z(n1020) );
  ANDN U1537 ( .B(n1025), .A(n1026), .Z(n1023) );
  XNOR U1538 ( .A(b[276]), .B(n1024), .Z(n1025) );
  XNOR U1539 ( .A(b[276]), .B(n1026), .Z(c[276]) );
  XOR U1540 ( .A(n1027), .B(n1028), .Z(n1024) );
  ANDN U1541 ( .B(n1029), .A(n1030), .Z(n1027) );
  XNOR U1542 ( .A(b[275]), .B(n1028), .Z(n1029) );
  XNOR U1543 ( .A(b[275]), .B(n1030), .Z(c[275]) );
  XOR U1544 ( .A(n1031), .B(n1032), .Z(n1028) );
  ANDN U1545 ( .B(n1033), .A(n1034), .Z(n1031) );
  XNOR U1546 ( .A(b[274]), .B(n1032), .Z(n1033) );
  XNOR U1547 ( .A(b[274]), .B(n1034), .Z(c[274]) );
  XOR U1548 ( .A(n1035), .B(n1036), .Z(n1032) );
  ANDN U1549 ( .B(n1037), .A(n1038), .Z(n1035) );
  XNOR U1550 ( .A(b[273]), .B(n1036), .Z(n1037) );
  XNOR U1551 ( .A(b[273]), .B(n1038), .Z(c[273]) );
  XOR U1552 ( .A(n1039), .B(n1040), .Z(n1036) );
  ANDN U1553 ( .B(n1041), .A(n1042), .Z(n1039) );
  XNOR U1554 ( .A(b[272]), .B(n1040), .Z(n1041) );
  XNOR U1555 ( .A(b[272]), .B(n1042), .Z(c[272]) );
  XOR U1556 ( .A(n1043), .B(n1044), .Z(n1040) );
  ANDN U1557 ( .B(n1045), .A(n1046), .Z(n1043) );
  XNOR U1558 ( .A(b[271]), .B(n1044), .Z(n1045) );
  XNOR U1559 ( .A(b[271]), .B(n1046), .Z(c[271]) );
  XOR U1560 ( .A(n1047), .B(n1048), .Z(n1044) );
  ANDN U1561 ( .B(n1049), .A(n1050), .Z(n1047) );
  XNOR U1562 ( .A(b[270]), .B(n1048), .Z(n1049) );
  XNOR U1563 ( .A(b[270]), .B(n1050), .Z(c[270]) );
  XOR U1564 ( .A(n1051), .B(n1052), .Z(n1048) );
  ANDN U1565 ( .B(n1053), .A(n1054), .Z(n1051) );
  XNOR U1566 ( .A(b[269]), .B(n1052), .Z(n1053) );
  XNOR U1567 ( .A(b[26]), .B(n1055), .Z(c[26]) );
  XNOR U1568 ( .A(b[269]), .B(n1054), .Z(c[269]) );
  XOR U1569 ( .A(n1056), .B(n1057), .Z(n1052) );
  ANDN U1570 ( .B(n1058), .A(n1059), .Z(n1056) );
  XNOR U1571 ( .A(b[268]), .B(n1057), .Z(n1058) );
  XNOR U1572 ( .A(b[268]), .B(n1059), .Z(c[268]) );
  XOR U1573 ( .A(n1060), .B(n1061), .Z(n1057) );
  ANDN U1574 ( .B(n1062), .A(n1063), .Z(n1060) );
  XNOR U1575 ( .A(b[267]), .B(n1061), .Z(n1062) );
  XNOR U1576 ( .A(b[267]), .B(n1063), .Z(c[267]) );
  XOR U1577 ( .A(n1064), .B(n1065), .Z(n1061) );
  ANDN U1578 ( .B(n1066), .A(n1067), .Z(n1064) );
  XNOR U1579 ( .A(b[266]), .B(n1065), .Z(n1066) );
  XNOR U1580 ( .A(b[266]), .B(n1067), .Z(c[266]) );
  XOR U1581 ( .A(n1068), .B(n1069), .Z(n1065) );
  ANDN U1582 ( .B(n1070), .A(n1071), .Z(n1068) );
  XNOR U1583 ( .A(b[265]), .B(n1069), .Z(n1070) );
  XNOR U1584 ( .A(b[265]), .B(n1071), .Z(c[265]) );
  XOR U1585 ( .A(n1072), .B(n1073), .Z(n1069) );
  ANDN U1586 ( .B(n1074), .A(n1075), .Z(n1072) );
  XNOR U1587 ( .A(b[264]), .B(n1073), .Z(n1074) );
  XNOR U1588 ( .A(b[264]), .B(n1075), .Z(c[264]) );
  XOR U1589 ( .A(n1076), .B(n1077), .Z(n1073) );
  ANDN U1590 ( .B(n1078), .A(n1079), .Z(n1076) );
  XNOR U1591 ( .A(b[263]), .B(n1077), .Z(n1078) );
  XNOR U1592 ( .A(b[263]), .B(n1079), .Z(c[263]) );
  XOR U1593 ( .A(n1080), .B(n1081), .Z(n1077) );
  ANDN U1594 ( .B(n1082), .A(n1083), .Z(n1080) );
  XNOR U1595 ( .A(b[262]), .B(n1081), .Z(n1082) );
  XNOR U1596 ( .A(b[262]), .B(n1083), .Z(c[262]) );
  XOR U1597 ( .A(n1084), .B(n1085), .Z(n1081) );
  ANDN U1598 ( .B(n1086), .A(n1087), .Z(n1084) );
  XNOR U1599 ( .A(b[261]), .B(n1085), .Z(n1086) );
  XNOR U1600 ( .A(b[261]), .B(n1087), .Z(c[261]) );
  XOR U1601 ( .A(n1088), .B(n1089), .Z(n1085) );
  ANDN U1602 ( .B(n1090), .A(n1091), .Z(n1088) );
  XNOR U1603 ( .A(b[260]), .B(n1089), .Z(n1090) );
  XNOR U1604 ( .A(b[260]), .B(n1091), .Z(c[260]) );
  XOR U1605 ( .A(n1092), .B(n1093), .Z(n1089) );
  ANDN U1606 ( .B(n1094), .A(n1095), .Z(n1092) );
  XNOR U1607 ( .A(b[259]), .B(n1093), .Z(n1094) );
  XNOR U1608 ( .A(b[25]), .B(n1096), .Z(c[25]) );
  XNOR U1609 ( .A(b[259]), .B(n1095), .Z(c[259]) );
  XOR U1610 ( .A(n1097), .B(n1098), .Z(n1093) );
  ANDN U1611 ( .B(n1099), .A(n1100), .Z(n1097) );
  XNOR U1612 ( .A(b[258]), .B(n1098), .Z(n1099) );
  XNOR U1613 ( .A(b[258]), .B(n1100), .Z(c[258]) );
  XOR U1614 ( .A(n1101), .B(n1102), .Z(n1098) );
  ANDN U1615 ( .B(n1103), .A(n1104), .Z(n1101) );
  XNOR U1616 ( .A(b[257]), .B(n1102), .Z(n1103) );
  XNOR U1617 ( .A(b[257]), .B(n1104), .Z(c[257]) );
  XOR U1618 ( .A(n1105), .B(n1106), .Z(n1102) );
  ANDN U1619 ( .B(n1107), .A(n1108), .Z(n1105) );
  XNOR U1620 ( .A(b[256]), .B(n1106), .Z(n1107) );
  XNOR U1621 ( .A(b[256]), .B(n1108), .Z(c[256]) );
  XOR U1622 ( .A(n1109), .B(n1110), .Z(n1106) );
  ANDN U1623 ( .B(n1111), .A(n1112), .Z(n1109) );
  XNOR U1624 ( .A(b[255]), .B(n1110), .Z(n1111) );
  XNOR U1625 ( .A(b[255]), .B(n1112), .Z(c[255]) );
  XOR U1626 ( .A(n1113), .B(n1114), .Z(n1110) );
  ANDN U1627 ( .B(n1115), .A(n1116), .Z(n1113) );
  XNOR U1628 ( .A(b[254]), .B(n1114), .Z(n1115) );
  XNOR U1629 ( .A(b[254]), .B(n1116), .Z(c[254]) );
  XOR U1630 ( .A(n1117), .B(n1118), .Z(n1114) );
  ANDN U1631 ( .B(n1119), .A(n1120), .Z(n1117) );
  XNOR U1632 ( .A(b[253]), .B(n1118), .Z(n1119) );
  XNOR U1633 ( .A(b[253]), .B(n1120), .Z(c[253]) );
  XOR U1634 ( .A(n1121), .B(n1122), .Z(n1118) );
  ANDN U1635 ( .B(n1123), .A(n1124), .Z(n1121) );
  XNOR U1636 ( .A(b[252]), .B(n1122), .Z(n1123) );
  XNOR U1637 ( .A(b[252]), .B(n1124), .Z(c[252]) );
  XOR U1638 ( .A(n1125), .B(n1126), .Z(n1122) );
  ANDN U1639 ( .B(n1127), .A(n1128), .Z(n1125) );
  XNOR U1640 ( .A(b[251]), .B(n1126), .Z(n1127) );
  XNOR U1641 ( .A(b[251]), .B(n1128), .Z(c[251]) );
  XOR U1642 ( .A(n1129), .B(n1130), .Z(n1126) );
  ANDN U1643 ( .B(n1131), .A(n1132), .Z(n1129) );
  XNOR U1644 ( .A(b[250]), .B(n1130), .Z(n1131) );
  XNOR U1645 ( .A(b[250]), .B(n1132), .Z(c[250]) );
  XOR U1646 ( .A(n1133), .B(n1134), .Z(n1130) );
  ANDN U1647 ( .B(n1135), .A(n1136), .Z(n1133) );
  XNOR U1648 ( .A(b[249]), .B(n1134), .Z(n1135) );
  XNOR U1649 ( .A(b[24]), .B(n1137), .Z(c[24]) );
  XNOR U1650 ( .A(b[249]), .B(n1136), .Z(c[249]) );
  XOR U1651 ( .A(n1138), .B(n1139), .Z(n1134) );
  ANDN U1652 ( .B(n1140), .A(n1141), .Z(n1138) );
  XNOR U1653 ( .A(b[248]), .B(n1139), .Z(n1140) );
  XNOR U1654 ( .A(b[248]), .B(n1141), .Z(c[248]) );
  XOR U1655 ( .A(n1142), .B(n1143), .Z(n1139) );
  ANDN U1656 ( .B(n1144), .A(n1145), .Z(n1142) );
  XNOR U1657 ( .A(b[247]), .B(n1143), .Z(n1144) );
  XNOR U1658 ( .A(b[247]), .B(n1145), .Z(c[247]) );
  XOR U1659 ( .A(n1146), .B(n1147), .Z(n1143) );
  ANDN U1660 ( .B(n1148), .A(n1149), .Z(n1146) );
  XNOR U1661 ( .A(b[246]), .B(n1147), .Z(n1148) );
  XNOR U1662 ( .A(b[246]), .B(n1149), .Z(c[246]) );
  XOR U1663 ( .A(n1150), .B(n1151), .Z(n1147) );
  ANDN U1664 ( .B(n1152), .A(n1153), .Z(n1150) );
  XNOR U1665 ( .A(b[245]), .B(n1151), .Z(n1152) );
  XNOR U1666 ( .A(b[245]), .B(n1153), .Z(c[245]) );
  XOR U1667 ( .A(n1154), .B(n1155), .Z(n1151) );
  ANDN U1668 ( .B(n1156), .A(n1157), .Z(n1154) );
  XNOR U1669 ( .A(b[244]), .B(n1155), .Z(n1156) );
  XNOR U1670 ( .A(b[244]), .B(n1157), .Z(c[244]) );
  XOR U1671 ( .A(n1158), .B(n1159), .Z(n1155) );
  ANDN U1672 ( .B(n1160), .A(n1161), .Z(n1158) );
  XNOR U1673 ( .A(b[243]), .B(n1159), .Z(n1160) );
  XNOR U1674 ( .A(b[243]), .B(n1161), .Z(c[243]) );
  XOR U1675 ( .A(n1162), .B(n1163), .Z(n1159) );
  ANDN U1676 ( .B(n1164), .A(n1165), .Z(n1162) );
  XNOR U1677 ( .A(b[242]), .B(n1163), .Z(n1164) );
  XNOR U1678 ( .A(b[242]), .B(n1165), .Z(c[242]) );
  XOR U1679 ( .A(n1166), .B(n1167), .Z(n1163) );
  ANDN U1680 ( .B(n1168), .A(n1169), .Z(n1166) );
  XNOR U1681 ( .A(b[241]), .B(n1167), .Z(n1168) );
  XNOR U1682 ( .A(b[241]), .B(n1169), .Z(c[241]) );
  XOR U1683 ( .A(n1170), .B(n1171), .Z(n1167) );
  ANDN U1684 ( .B(n1172), .A(n1173), .Z(n1170) );
  XNOR U1685 ( .A(b[240]), .B(n1171), .Z(n1172) );
  XNOR U1686 ( .A(b[240]), .B(n1173), .Z(c[240]) );
  XOR U1687 ( .A(n1174), .B(n1175), .Z(n1171) );
  ANDN U1688 ( .B(n1176), .A(n1177), .Z(n1174) );
  XNOR U1689 ( .A(b[239]), .B(n1175), .Z(n1176) );
  XNOR U1690 ( .A(b[23]), .B(n1178), .Z(c[23]) );
  XNOR U1691 ( .A(b[239]), .B(n1177), .Z(c[239]) );
  XOR U1692 ( .A(n1179), .B(n1180), .Z(n1175) );
  ANDN U1693 ( .B(n1181), .A(n1182), .Z(n1179) );
  XNOR U1694 ( .A(b[238]), .B(n1180), .Z(n1181) );
  XNOR U1695 ( .A(b[238]), .B(n1182), .Z(c[238]) );
  XOR U1696 ( .A(n1183), .B(n1184), .Z(n1180) );
  ANDN U1697 ( .B(n1185), .A(n1186), .Z(n1183) );
  XNOR U1698 ( .A(b[237]), .B(n1184), .Z(n1185) );
  XNOR U1699 ( .A(b[237]), .B(n1186), .Z(c[237]) );
  XOR U1700 ( .A(n1187), .B(n1188), .Z(n1184) );
  ANDN U1701 ( .B(n1189), .A(n1190), .Z(n1187) );
  XNOR U1702 ( .A(b[236]), .B(n1188), .Z(n1189) );
  XNOR U1703 ( .A(b[236]), .B(n1190), .Z(c[236]) );
  XOR U1704 ( .A(n1191), .B(n1192), .Z(n1188) );
  ANDN U1705 ( .B(n1193), .A(n1194), .Z(n1191) );
  XNOR U1706 ( .A(b[235]), .B(n1192), .Z(n1193) );
  XNOR U1707 ( .A(b[235]), .B(n1194), .Z(c[235]) );
  XOR U1708 ( .A(n1195), .B(n1196), .Z(n1192) );
  ANDN U1709 ( .B(n1197), .A(n1198), .Z(n1195) );
  XNOR U1710 ( .A(b[234]), .B(n1196), .Z(n1197) );
  XNOR U1711 ( .A(b[234]), .B(n1198), .Z(c[234]) );
  XOR U1712 ( .A(n1199), .B(n1200), .Z(n1196) );
  ANDN U1713 ( .B(n1201), .A(n1202), .Z(n1199) );
  XNOR U1714 ( .A(b[233]), .B(n1200), .Z(n1201) );
  XNOR U1715 ( .A(b[233]), .B(n1202), .Z(c[233]) );
  XOR U1716 ( .A(n1203), .B(n1204), .Z(n1200) );
  ANDN U1717 ( .B(n1205), .A(n1206), .Z(n1203) );
  XNOR U1718 ( .A(b[232]), .B(n1204), .Z(n1205) );
  XNOR U1719 ( .A(b[232]), .B(n1206), .Z(c[232]) );
  XOR U1720 ( .A(n1207), .B(n1208), .Z(n1204) );
  ANDN U1721 ( .B(n1209), .A(n1210), .Z(n1207) );
  XNOR U1722 ( .A(b[231]), .B(n1208), .Z(n1209) );
  XNOR U1723 ( .A(b[231]), .B(n1210), .Z(c[231]) );
  XOR U1724 ( .A(n1211), .B(n1212), .Z(n1208) );
  ANDN U1725 ( .B(n1213), .A(n1214), .Z(n1211) );
  XNOR U1726 ( .A(b[230]), .B(n1212), .Z(n1213) );
  XNOR U1727 ( .A(b[230]), .B(n1214), .Z(c[230]) );
  XOR U1728 ( .A(n1215), .B(n1216), .Z(n1212) );
  ANDN U1729 ( .B(n1217), .A(n1218), .Z(n1215) );
  XNOR U1730 ( .A(b[229]), .B(n1216), .Z(n1217) );
  XNOR U1731 ( .A(b[22]), .B(n1219), .Z(c[22]) );
  XNOR U1732 ( .A(b[229]), .B(n1218), .Z(c[229]) );
  XOR U1733 ( .A(n1220), .B(n1221), .Z(n1216) );
  ANDN U1734 ( .B(n1222), .A(n1223), .Z(n1220) );
  XNOR U1735 ( .A(b[228]), .B(n1221), .Z(n1222) );
  XNOR U1736 ( .A(b[228]), .B(n1223), .Z(c[228]) );
  XOR U1737 ( .A(n1224), .B(n1225), .Z(n1221) );
  ANDN U1738 ( .B(n1226), .A(n1227), .Z(n1224) );
  XNOR U1739 ( .A(b[227]), .B(n1225), .Z(n1226) );
  XNOR U1740 ( .A(b[227]), .B(n1227), .Z(c[227]) );
  XOR U1741 ( .A(n1228), .B(n1229), .Z(n1225) );
  ANDN U1742 ( .B(n1230), .A(n1231), .Z(n1228) );
  XNOR U1743 ( .A(b[226]), .B(n1229), .Z(n1230) );
  XNOR U1744 ( .A(b[226]), .B(n1231), .Z(c[226]) );
  XOR U1745 ( .A(n1232), .B(n1233), .Z(n1229) );
  ANDN U1746 ( .B(n1234), .A(n1235), .Z(n1232) );
  XNOR U1747 ( .A(b[225]), .B(n1233), .Z(n1234) );
  XNOR U1748 ( .A(b[225]), .B(n1235), .Z(c[225]) );
  XOR U1749 ( .A(n1236), .B(n1237), .Z(n1233) );
  ANDN U1750 ( .B(n1238), .A(n1239), .Z(n1236) );
  XNOR U1751 ( .A(b[224]), .B(n1237), .Z(n1238) );
  XNOR U1752 ( .A(b[224]), .B(n1239), .Z(c[224]) );
  XOR U1753 ( .A(n1240), .B(n1241), .Z(n1237) );
  ANDN U1754 ( .B(n1242), .A(n1243), .Z(n1240) );
  XNOR U1755 ( .A(b[223]), .B(n1241), .Z(n1242) );
  XNOR U1756 ( .A(b[223]), .B(n1243), .Z(c[223]) );
  XOR U1757 ( .A(n1244), .B(n1245), .Z(n1241) );
  ANDN U1758 ( .B(n1246), .A(n1247), .Z(n1244) );
  XNOR U1759 ( .A(b[222]), .B(n1245), .Z(n1246) );
  XNOR U1760 ( .A(b[222]), .B(n1247), .Z(c[222]) );
  XOR U1761 ( .A(n1248), .B(n1249), .Z(n1245) );
  ANDN U1762 ( .B(n1250), .A(n1251), .Z(n1248) );
  XNOR U1763 ( .A(b[221]), .B(n1249), .Z(n1250) );
  XNOR U1764 ( .A(b[221]), .B(n1251), .Z(c[221]) );
  XOR U1765 ( .A(n1252), .B(n1253), .Z(n1249) );
  ANDN U1766 ( .B(n1254), .A(n1255), .Z(n1252) );
  XNOR U1767 ( .A(b[220]), .B(n1253), .Z(n1254) );
  XNOR U1768 ( .A(b[220]), .B(n1255), .Z(c[220]) );
  XOR U1769 ( .A(n1256), .B(n1257), .Z(n1253) );
  ANDN U1770 ( .B(n1258), .A(n1259), .Z(n1256) );
  XNOR U1771 ( .A(b[219]), .B(n1257), .Z(n1258) );
  XNOR U1772 ( .A(b[21]), .B(n1260), .Z(c[21]) );
  XNOR U1773 ( .A(b[219]), .B(n1259), .Z(c[219]) );
  XOR U1774 ( .A(n1261), .B(n1262), .Z(n1257) );
  ANDN U1775 ( .B(n1263), .A(n1264), .Z(n1261) );
  XNOR U1776 ( .A(b[218]), .B(n1262), .Z(n1263) );
  XNOR U1777 ( .A(b[218]), .B(n1264), .Z(c[218]) );
  XOR U1778 ( .A(n1265), .B(n1266), .Z(n1262) );
  ANDN U1779 ( .B(n1267), .A(n1268), .Z(n1265) );
  XNOR U1780 ( .A(b[217]), .B(n1266), .Z(n1267) );
  XNOR U1781 ( .A(b[217]), .B(n1268), .Z(c[217]) );
  XOR U1782 ( .A(n1269), .B(n1270), .Z(n1266) );
  ANDN U1783 ( .B(n1271), .A(n1272), .Z(n1269) );
  XNOR U1784 ( .A(b[216]), .B(n1270), .Z(n1271) );
  XNOR U1785 ( .A(b[216]), .B(n1272), .Z(c[216]) );
  XOR U1786 ( .A(n1273), .B(n1274), .Z(n1270) );
  ANDN U1787 ( .B(n1275), .A(n1276), .Z(n1273) );
  XNOR U1788 ( .A(b[215]), .B(n1274), .Z(n1275) );
  XNOR U1789 ( .A(b[215]), .B(n1276), .Z(c[215]) );
  XOR U1790 ( .A(n1277), .B(n1278), .Z(n1274) );
  ANDN U1791 ( .B(n1279), .A(n1280), .Z(n1277) );
  XNOR U1792 ( .A(b[214]), .B(n1278), .Z(n1279) );
  XNOR U1793 ( .A(b[214]), .B(n1280), .Z(c[214]) );
  XOR U1794 ( .A(n1281), .B(n1282), .Z(n1278) );
  ANDN U1795 ( .B(n1283), .A(n1284), .Z(n1281) );
  XNOR U1796 ( .A(b[213]), .B(n1282), .Z(n1283) );
  XNOR U1797 ( .A(b[213]), .B(n1284), .Z(c[213]) );
  XOR U1798 ( .A(n1285), .B(n1286), .Z(n1282) );
  ANDN U1799 ( .B(n1287), .A(n1288), .Z(n1285) );
  XNOR U1800 ( .A(b[212]), .B(n1286), .Z(n1287) );
  XNOR U1801 ( .A(b[212]), .B(n1288), .Z(c[212]) );
  XOR U1802 ( .A(n1289), .B(n1290), .Z(n1286) );
  ANDN U1803 ( .B(n1291), .A(n1292), .Z(n1289) );
  XNOR U1804 ( .A(b[211]), .B(n1290), .Z(n1291) );
  XNOR U1805 ( .A(b[211]), .B(n1292), .Z(c[211]) );
  XOR U1806 ( .A(n1293), .B(n1294), .Z(n1290) );
  ANDN U1807 ( .B(n1295), .A(n1296), .Z(n1293) );
  XNOR U1808 ( .A(b[210]), .B(n1294), .Z(n1295) );
  XNOR U1809 ( .A(b[210]), .B(n1296), .Z(c[210]) );
  XOR U1810 ( .A(n1297), .B(n1298), .Z(n1294) );
  ANDN U1811 ( .B(n1299), .A(n1300), .Z(n1297) );
  XNOR U1812 ( .A(b[209]), .B(n1298), .Z(n1299) );
  XNOR U1813 ( .A(b[20]), .B(n1301), .Z(c[20]) );
  XNOR U1814 ( .A(b[209]), .B(n1300), .Z(c[209]) );
  XOR U1815 ( .A(n1302), .B(n1303), .Z(n1298) );
  ANDN U1816 ( .B(n1304), .A(n1305), .Z(n1302) );
  XNOR U1817 ( .A(b[208]), .B(n1303), .Z(n1304) );
  XNOR U1818 ( .A(b[208]), .B(n1305), .Z(c[208]) );
  XOR U1819 ( .A(n1306), .B(n1307), .Z(n1303) );
  ANDN U1820 ( .B(n1308), .A(n1309), .Z(n1306) );
  XNOR U1821 ( .A(b[207]), .B(n1307), .Z(n1308) );
  XNOR U1822 ( .A(b[207]), .B(n1309), .Z(c[207]) );
  XOR U1823 ( .A(n1310), .B(n1311), .Z(n1307) );
  ANDN U1824 ( .B(n1312), .A(n1313), .Z(n1310) );
  XNOR U1825 ( .A(b[206]), .B(n1311), .Z(n1312) );
  XNOR U1826 ( .A(b[206]), .B(n1313), .Z(c[206]) );
  XOR U1827 ( .A(n1314), .B(n1315), .Z(n1311) );
  ANDN U1828 ( .B(n1316), .A(n1317), .Z(n1314) );
  XNOR U1829 ( .A(b[205]), .B(n1315), .Z(n1316) );
  XNOR U1830 ( .A(b[205]), .B(n1317), .Z(c[205]) );
  XOR U1831 ( .A(n1318), .B(n1319), .Z(n1315) );
  ANDN U1832 ( .B(n1320), .A(n1321), .Z(n1318) );
  XNOR U1833 ( .A(b[204]), .B(n1319), .Z(n1320) );
  XNOR U1834 ( .A(b[204]), .B(n1321), .Z(c[204]) );
  XOR U1835 ( .A(n1322), .B(n1323), .Z(n1319) );
  ANDN U1836 ( .B(n1324), .A(n1325), .Z(n1322) );
  XNOR U1837 ( .A(b[203]), .B(n1323), .Z(n1324) );
  XNOR U1838 ( .A(b[203]), .B(n1325), .Z(c[203]) );
  XOR U1839 ( .A(n1326), .B(n1327), .Z(n1323) );
  ANDN U1840 ( .B(n1328), .A(n1329), .Z(n1326) );
  XNOR U1841 ( .A(b[202]), .B(n1327), .Z(n1328) );
  XNOR U1842 ( .A(b[202]), .B(n1329), .Z(c[202]) );
  XOR U1843 ( .A(n1330), .B(n1331), .Z(n1327) );
  ANDN U1844 ( .B(n1332), .A(n1333), .Z(n1330) );
  XNOR U1845 ( .A(b[201]), .B(n1331), .Z(n1332) );
  XNOR U1846 ( .A(b[201]), .B(n1333), .Z(c[201]) );
  XOR U1847 ( .A(n1334), .B(n1335), .Z(n1331) );
  ANDN U1848 ( .B(n1336), .A(n1337), .Z(n1334) );
  XNOR U1849 ( .A(b[200]), .B(n1335), .Z(n1336) );
  XNOR U1850 ( .A(b[200]), .B(n1337), .Z(c[200]) );
  XOR U1851 ( .A(n1338), .B(n1339), .Z(n1335) );
  ANDN U1852 ( .B(n1340), .A(n1341), .Z(n1338) );
  XNOR U1853 ( .A(b[199]), .B(n1339), .Z(n1340) );
  XNOR U1854 ( .A(b[1]), .B(n1342), .Z(c[1]) );
  XNOR U1855 ( .A(b[19]), .B(n1343), .Z(c[19]) );
  XNOR U1856 ( .A(b[199]), .B(n1341), .Z(c[199]) );
  XOR U1857 ( .A(n1344), .B(n1345), .Z(n1339) );
  ANDN U1858 ( .B(n1346), .A(n1347), .Z(n1344) );
  XNOR U1859 ( .A(b[198]), .B(n1345), .Z(n1346) );
  XNOR U1860 ( .A(b[198]), .B(n1347), .Z(c[198]) );
  XOR U1861 ( .A(n1348), .B(n1349), .Z(n1345) );
  ANDN U1862 ( .B(n1350), .A(n1351), .Z(n1348) );
  XNOR U1863 ( .A(b[197]), .B(n1349), .Z(n1350) );
  XNOR U1864 ( .A(b[197]), .B(n1351), .Z(c[197]) );
  XOR U1865 ( .A(n1352), .B(n1353), .Z(n1349) );
  ANDN U1866 ( .B(n1354), .A(n1355), .Z(n1352) );
  XNOR U1867 ( .A(b[196]), .B(n1353), .Z(n1354) );
  XNOR U1868 ( .A(b[196]), .B(n1355), .Z(c[196]) );
  XOR U1869 ( .A(n1356), .B(n1357), .Z(n1353) );
  ANDN U1870 ( .B(n1358), .A(n1359), .Z(n1356) );
  XNOR U1871 ( .A(b[195]), .B(n1357), .Z(n1358) );
  XNOR U1872 ( .A(b[195]), .B(n1359), .Z(c[195]) );
  XOR U1873 ( .A(n1360), .B(n1361), .Z(n1357) );
  ANDN U1874 ( .B(n1362), .A(n1363), .Z(n1360) );
  XNOR U1875 ( .A(b[194]), .B(n1361), .Z(n1362) );
  XNOR U1876 ( .A(b[194]), .B(n1363), .Z(c[194]) );
  XOR U1877 ( .A(n1364), .B(n1365), .Z(n1361) );
  ANDN U1878 ( .B(n1366), .A(n1367), .Z(n1364) );
  XNOR U1879 ( .A(b[193]), .B(n1365), .Z(n1366) );
  XNOR U1880 ( .A(b[193]), .B(n1367), .Z(c[193]) );
  XOR U1881 ( .A(n1368), .B(n1369), .Z(n1365) );
  ANDN U1882 ( .B(n1370), .A(n1371), .Z(n1368) );
  XNOR U1883 ( .A(b[192]), .B(n1369), .Z(n1370) );
  XNOR U1884 ( .A(b[192]), .B(n1371), .Z(c[192]) );
  XOR U1885 ( .A(n1372), .B(n1373), .Z(n1369) );
  ANDN U1886 ( .B(n1374), .A(n1375), .Z(n1372) );
  XNOR U1887 ( .A(b[191]), .B(n1373), .Z(n1374) );
  XNOR U1888 ( .A(b[191]), .B(n1375), .Z(c[191]) );
  XOR U1889 ( .A(n1376), .B(n1377), .Z(n1373) );
  ANDN U1890 ( .B(n1378), .A(n1379), .Z(n1376) );
  XNOR U1891 ( .A(b[190]), .B(n1377), .Z(n1378) );
  XNOR U1892 ( .A(b[190]), .B(n1379), .Z(c[190]) );
  XOR U1893 ( .A(n1380), .B(n1381), .Z(n1377) );
  ANDN U1894 ( .B(n1382), .A(n1383), .Z(n1380) );
  XNOR U1895 ( .A(b[189]), .B(n1381), .Z(n1382) );
  XNOR U1896 ( .A(b[18]), .B(n1384), .Z(c[18]) );
  XNOR U1897 ( .A(b[189]), .B(n1383), .Z(c[189]) );
  XOR U1898 ( .A(n1385), .B(n1386), .Z(n1381) );
  ANDN U1899 ( .B(n1387), .A(n1388), .Z(n1385) );
  XNOR U1900 ( .A(b[188]), .B(n1386), .Z(n1387) );
  XNOR U1901 ( .A(b[188]), .B(n1388), .Z(c[188]) );
  XOR U1902 ( .A(n1389), .B(n1390), .Z(n1386) );
  ANDN U1903 ( .B(n1391), .A(n1392), .Z(n1389) );
  XNOR U1904 ( .A(b[187]), .B(n1390), .Z(n1391) );
  XNOR U1905 ( .A(b[187]), .B(n1392), .Z(c[187]) );
  XOR U1906 ( .A(n1393), .B(n1394), .Z(n1390) );
  ANDN U1907 ( .B(n1395), .A(n1396), .Z(n1393) );
  XNOR U1908 ( .A(b[186]), .B(n1394), .Z(n1395) );
  XNOR U1909 ( .A(b[186]), .B(n1396), .Z(c[186]) );
  XOR U1910 ( .A(n1397), .B(n1398), .Z(n1394) );
  ANDN U1911 ( .B(n1399), .A(n1400), .Z(n1397) );
  XNOR U1912 ( .A(b[185]), .B(n1398), .Z(n1399) );
  XNOR U1913 ( .A(b[185]), .B(n1400), .Z(c[185]) );
  XOR U1914 ( .A(n1401), .B(n1402), .Z(n1398) );
  ANDN U1915 ( .B(n1403), .A(n1404), .Z(n1401) );
  XNOR U1916 ( .A(b[184]), .B(n1402), .Z(n1403) );
  XNOR U1917 ( .A(b[184]), .B(n1404), .Z(c[184]) );
  XOR U1918 ( .A(n1405), .B(n1406), .Z(n1402) );
  ANDN U1919 ( .B(n1407), .A(n1408), .Z(n1405) );
  XNOR U1920 ( .A(b[183]), .B(n1406), .Z(n1407) );
  XNOR U1921 ( .A(b[183]), .B(n1408), .Z(c[183]) );
  XOR U1922 ( .A(n1409), .B(n1410), .Z(n1406) );
  ANDN U1923 ( .B(n1411), .A(n1412), .Z(n1409) );
  XNOR U1924 ( .A(b[182]), .B(n1410), .Z(n1411) );
  XNOR U1925 ( .A(b[182]), .B(n1412), .Z(c[182]) );
  XOR U1926 ( .A(n1413), .B(n1414), .Z(n1410) );
  ANDN U1927 ( .B(n1415), .A(n1416), .Z(n1413) );
  XNOR U1928 ( .A(b[181]), .B(n1414), .Z(n1415) );
  XNOR U1929 ( .A(b[181]), .B(n1416), .Z(c[181]) );
  XOR U1930 ( .A(n1417), .B(n1418), .Z(n1414) );
  ANDN U1931 ( .B(n1419), .A(n1420), .Z(n1417) );
  XNOR U1932 ( .A(b[180]), .B(n1418), .Z(n1419) );
  XNOR U1933 ( .A(b[180]), .B(n1420), .Z(c[180]) );
  XOR U1934 ( .A(n1421), .B(n1422), .Z(n1418) );
  ANDN U1935 ( .B(n1423), .A(n1424), .Z(n1421) );
  XNOR U1936 ( .A(b[179]), .B(n1422), .Z(n1423) );
  XNOR U1937 ( .A(b[17]), .B(n1425), .Z(c[17]) );
  XNOR U1938 ( .A(b[179]), .B(n1424), .Z(c[179]) );
  XOR U1939 ( .A(n1426), .B(n1427), .Z(n1422) );
  ANDN U1940 ( .B(n1428), .A(n1429), .Z(n1426) );
  XNOR U1941 ( .A(b[178]), .B(n1427), .Z(n1428) );
  XNOR U1942 ( .A(b[178]), .B(n1429), .Z(c[178]) );
  XOR U1943 ( .A(n1430), .B(n1431), .Z(n1427) );
  ANDN U1944 ( .B(n1432), .A(n1433), .Z(n1430) );
  XNOR U1945 ( .A(b[177]), .B(n1431), .Z(n1432) );
  XNOR U1946 ( .A(b[177]), .B(n1433), .Z(c[177]) );
  XOR U1947 ( .A(n1434), .B(n1435), .Z(n1431) );
  ANDN U1948 ( .B(n1436), .A(n1437), .Z(n1434) );
  XNOR U1949 ( .A(b[176]), .B(n1435), .Z(n1436) );
  XNOR U1950 ( .A(b[176]), .B(n1437), .Z(c[176]) );
  XOR U1951 ( .A(n1438), .B(n1439), .Z(n1435) );
  ANDN U1952 ( .B(n1440), .A(n1441), .Z(n1438) );
  XNOR U1953 ( .A(b[175]), .B(n1439), .Z(n1440) );
  XNOR U1954 ( .A(b[175]), .B(n1441), .Z(c[175]) );
  XOR U1955 ( .A(n1442), .B(n1443), .Z(n1439) );
  ANDN U1956 ( .B(n1444), .A(n1445), .Z(n1442) );
  XNOR U1957 ( .A(b[174]), .B(n1443), .Z(n1444) );
  XNOR U1958 ( .A(b[174]), .B(n1445), .Z(c[174]) );
  XOR U1959 ( .A(n1446), .B(n1447), .Z(n1443) );
  ANDN U1960 ( .B(n1448), .A(n1449), .Z(n1446) );
  XNOR U1961 ( .A(b[173]), .B(n1447), .Z(n1448) );
  XNOR U1962 ( .A(b[173]), .B(n1449), .Z(c[173]) );
  XOR U1963 ( .A(n1450), .B(n1451), .Z(n1447) );
  ANDN U1964 ( .B(n1452), .A(n1453), .Z(n1450) );
  XNOR U1965 ( .A(b[172]), .B(n1451), .Z(n1452) );
  XNOR U1966 ( .A(b[172]), .B(n1453), .Z(c[172]) );
  XOR U1967 ( .A(n1454), .B(n1455), .Z(n1451) );
  ANDN U1968 ( .B(n1456), .A(n1457), .Z(n1454) );
  XNOR U1969 ( .A(b[171]), .B(n1455), .Z(n1456) );
  XNOR U1970 ( .A(b[171]), .B(n1457), .Z(c[171]) );
  XOR U1971 ( .A(n1458), .B(n1459), .Z(n1455) );
  ANDN U1972 ( .B(n1460), .A(n1461), .Z(n1458) );
  XNOR U1973 ( .A(b[170]), .B(n1459), .Z(n1460) );
  XNOR U1974 ( .A(b[170]), .B(n1461), .Z(c[170]) );
  XOR U1975 ( .A(n1462), .B(n1463), .Z(n1459) );
  ANDN U1976 ( .B(n1464), .A(n1465), .Z(n1462) );
  XNOR U1977 ( .A(b[169]), .B(n1463), .Z(n1464) );
  XNOR U1978 ( .A(b[16]), .B(n1466), .Z(c[16]) );
  XNOR U1979 ( .A(b[169]), .B(n1465), .Z(c[169]) );
  XOR U1980 ( .A(n1467), .B(n1468), .Z(n1463) );
  ANDN U1981 ( .B(n1469), .A(n1470), .Z(n1467) );
  XNOR U1982 ( .A(b[168]), .B(n1468), .Z(n1469) );
  XNOR U1983 ( .A(b[168]), .B(n1470), .Z(c[168]) );
  XOR U1984 ( .A(n1471), .B(n1472), .Z(n1468) );
  ANDN U1985 ( .B(n1473), .A(n1474), .Z(n1471) );
  XNOR U1986 ( .A(b[167]), .B(n1472), .Z(n1473) );
  XNOR U1987 ( .A(b[167]), .B(n1474), .Z(c[167]) );
  XOR U1988 ( .A(n1475), .B(n1476), .Z(n1472) );
  ANDN U1989 ( .B(n1477), .A(n1478), .Z(n1475) );
  XNOR U1990 ( .A(b[166]), .B(n1476), .Z(n1477) );
  XNOR U1991 ( .A(b[166]), .B(n1478), .Z(c[166]) );
  XOR U1992 ( .A(n1479), .B(n1480), .Z(n1476) );
  ANDN U1993 ( .B(n1481), .A(n1482), .Z(n1479) );
  XNOR U1994 ( .A(b[165]), .B(n1480), .Z(n1481) );
  XNOR U1995 ( .A(b[165]), .B(n1482), .Z(c[165]) );
  XOR U1996 ( .A(n1483), .B(n1484), .Z(n1480) );
  ANDN U1997 ( .B(n1485), .A(n1486), .Z(n1483) );
  XNOR U1998 ( .A(b[164]), .B(n1484), .Z(n1485) );
  XNOR U1999 ( .A(b[164]), .B(n1486), .Z(c[164]) );
  XOR U2000 ( .A(n1487), .B(n1488), .Z(n1484) );
  ANDN U2001 ( .B(n1489), .A(n1490), .Z(n1487) );
  XNOR U2002 ( .A(b[163]), .B(n1488), .Z(n1489) );
  XNOR U2003 ( .A(b[163]), .B(n1490), .Z(c[163]) );
  XOR U2004 ( .A(n1491), .B(n1492), .Z(n1488) );
  ANDN U2005 ( .B(n1493), .A(n1494), .Z(n1491) );
  XNOR U2006 ( .A(b[162]), .B(n1492), .Z(n1493) );
  XNOR U2007 ( .A(b[162]), .B(n1494), .Z(c[162]) );
  XOR U2008 ( .A(n1495), .B(n1496), .Z(n1492) );
  ANDN U2009 ( .B(n1497), .A(n1498), .Z(n1495) );
  XNOR U2010 ( .A(b[161]), .B(n1496), .Z(n1497) );
  XNOR U2011 ( .A(b[161]), .B(n1498), .Z(c[161]) );
  XOR U2012 ( .A(n1499), .B(n1500), .Z(n1496) );
  ANDN U2013 ( .B(n1501), .A(n1502), .Z(n1499) );
  XNOR U2014 ( .A(b[160]), .B(n1500), .Z(n1501) );
  XNOR U2015 ( .A(b[160]), .B(n1502), .Z(c[160]) );
  XOR U2016 ( .A(n1503), .B(n1504), .Z(n1500) );
  ANDN U2017 ( .B(n1505), .A(n1506), .Z(n1503) );
  XNOR U2018 ( .A(b[159]), .B(n1504), .Z(n1505) );
  XNOR U2019 ( .A(b[15]), .B(n1507), .Z(c[15]) );
  XNOR U2020 ( .A(b[159]), .B(n1506), .Z(c[159]) );
  XOR U2021 ( .A(n1508), .B(n1509), .Z(n1504) );
  ANDN U2022 ( .B(n1510), .A(n1511), .Z(n1508) );
  XNOR U2023 ( .A(b[158]), .B(n1509), .Z(n1510) );
  XNOR U2024 ( .A(b[158]), .B(n1511), .Z(c[158]) );
  XOR U2025 ( .A(n1512), .B(n1513), .Z(n1509) );
  ANDN U2026 ( .B(n1514), .A(n1515), .Z(n1512) );
  XNOR U2027 ( .A(b[157]), .B(n1513), .Z(n1514) );
  XNOR U2028 ( .A(b[157]), .B(n1515), .Z(c[157]) );
  XOR U2029 ( .A(n1516), .B(n1517), .Z(n1513) );
  ANDN U2030 ( .B(n1518), .A(n1519), .Z(n1516) );
  XNOR U2031 ( .A(b[156]), .B(n1517), .Z(n1518) );
  XNOR U2032 ( .A(b[156]), .B(n1519), .Z(c[156]) );
  XOR U2033 ( .A(n1520), .B(n1521), .Z(n1517) );
  ANDN U2034 ( .B(n1522), .A(n1523), .Z(n1520) );
  XNOR U2035 ( .A(b[155]), .B(n1521), .Z(n1522) );
  XNOR U2036 ( .A(b[155]), .B(n1523), .Z(c[155]) );
  XOR U2037 ( .A(n1524), .B(n1525), .Z(n1521) );
  ANDN U2038 ( .B(n1526), .A(n1527), .Z(n1524) );
  XNOR U2039 ( .A(b[154]), .B(n1525), .Z(n1526) );
  XNOR U2040 ( .A(b[154]), .B(n1527), .Z(c[154]) );
  XOR U2041 ( .A(n1528), .B(n1529), .Z(n1525) );
  ANDN U2042 ( .B(n1530), .A(n1531), .Z(n1528) );
  XNOR U2043 ( .A(b[153]), .B(n1529), .Z(n1530) );
  XNOR U2044 ( .A(b[153]), .B(n1531), .Z(c[153]) );
  XOR U2045 ( .A(n1532), .B(n1533), .Z(n1529) );
  ANDN U2046 ( .B(n1534), .A(n1535), .Z(n1532) );
  XNOR U2047 ( .A(b[152]), .B(n1533), .Z(n1534) );
  XNOR U2048 ( .A(b[152]), .B(n1535), .Z(c[152]) );
  XOR U2049 ( .A(n1536), .B(n1537), .Z(n1533) );
  ANDN U2050 ( .B(n1538), .A(n1539), .Z(n1536) );
  XNOR U2051 ( .A(b[151]), .B(n1537), .Z(n1538) );
  XNOR U2052 ( .A(b[151]), .B(n1539), .Z(c[151]) );
  XOR U2053 ( .A(n1540), .B(n1541), .Z(n1537) );
  ANDN U2054 ( .B(n1542), .A(n1543), .Z(n1540) );
  XNOR U2055 ( .A(b[150]), .B(n1541), .Z(n1542) );
  XNOR U2056 ( .A(b[150]), .B(n1543), .Z(c[150]) );
  XOR U2057 ( .A(n1544), .B(n1545), .Z(n1541) );
  ANDN U2058 ( .B(n1546), .A(n1547), .Z(n1544) );
  XNOR U2059 ( .A(b[149]), .B(n1545), .Z(n1546) );
  XNOR U2060 ( .A(b[14]), .B(n1548), .Z(c[14]) );
  XNOR U2061 ( .A(b[149]), .B(n1547), .Z(c[149]) );
  XOR U2062 ( .A(n1549), .B(n1550), .Z(n1545) );
  ANDN U2063 ( .B(n1551), .A(n1552), .Z(n1549) );
  XNOR U2064 ( .A(b[148]), .B(n1550), .Z(n1551) );
  XNOR U2065 ( .A(b[148]), .B(n1552), .Z(c[148]) );
  XOR U2066 ( .A(n1553), .B(n1554), .Z(n1550) );
  ANDN U2067 ( .B(n1555), .A(n1556), .Z(n1553) );
  XNOR U2068 ( .A(b[147]), .B(n1554), .Z(n1555) );
  XNOR U2069 ( .A(b[147]), .B(n1556), .Z(c[147]) );
  XOR U2070 ( .A(n1557), .B(n1558), .Z(n1554) );
  ANDN U2071 ( .B(n1559), .A(n1560), .Z(n1557) );
  XNOR U2072 ( .A(b[146]), .B(n1558), .Z(n1559) );
  XNOR U2073 ( .A(b[146]), .B(n1560), .Z(c[146]) );
  XOR U2074 ( .A(n1561), .B(n1562), .Z(n1558) );
  ANDN U2075 ( .B(n1563), .A(n1564), .Z(n1561) );
  XNOR U2076 ( .A(b[145]), .B(n1562), .Z(n1563) );
  XNOR U2077 ( .A(b[145]), .B(n1564), .Z(c[145]) );
  XOR U2078 ( .A(n1565), .B(n1566), .Z(n1562) );
  ANDN U2079 ( .B(n1567), .A(n1568), .Z(n1565) );
  XNOR U2080 ( .A(b[144]), .B(n1566), .Z(n1567) );
  XNOR U2081 ( .A(b[144]), .B(n1568), .Z(c[144]) );
  XOR U2082 ( .A(n1569), .B(n1570), .Z(n1566) );
  ANDN U2083 ( .B(n1571), .A(n1572), .Z(n1569) );
  XNOR U2084 ( .A(b[143]), .B(n1570), .Z(n1571) );
  XNOR U2085 ( .A(b[143]), .B(n1572), .Z(c[143]) );
  XOR U2086 ( .A(n1573), .B(n1574), .Z(n1570) );
  ANDN U2087 ( .B(n1575), .A(n1576), .Z(n1573) );
  XNOR U2088 ( .A(b[142]), .B(n1574), .Z(n1575) );
  XNOR U2089 ( .A(b[142]), .B(n1576), .Z(c[142]) );
  XOR U2090 ( .A(n1577), .B(n1578), .Z(n1574) );
  ANDN U2091 ( .B(n1579), .A(n1580), .Z(n1577) );
  XNOR U2092 ( .A(b[141]), .B(n1578), .Z(n1579) );
  XNOR U2093 ( .A(b[141]), .B(n1580), .Z(c[141]) );
  XOR U2094 ( .A(n1581), .B(n1582), .Z(n1578) );
  ANDN U2095 ( .B(n1583), .A(n1584), .Z(n1581) );
  XNOR U2096 ( .A(b[140]), .B(n1582), .Z(n1583) );
  XNOR U2097 ( .A(b[140]), .B(n1584), .Z(c[140]) );
  XOR U2098 ( .A(n1585), .B(n1586), .Z(n1582) );
  ANDN U2099 ( .B(n1587), .A(n1588), .Z(n1585) );
  XNOR U2100 ( .A(b[139]), .B(n1586), .Z(n1587) );
  XNOR U2101 ( .A(b[13]), .B(n1589), .Z(c[13]) );
  XNOR U2102 ( .A(b[139]), .B(n1588), .Z(c[139]) );
  XOR U2103 ( .A(n1590), .B(n1591), .Z(n1586) );
  ANDN U2104 ( .B(n1592), .A(n1593), .Z(n1590) );
  XNOR U2105 ( .A(b[138]), .B(n1591), .Z(n1592) );
  XNOR U2106 ( .A(b[138]), .B(n1593), .Z(c[138]) );
  XOR U2107 ( .A(n1594), .B(n1595), .Z(n1591) );
  ANDN U2108 ( .B(n1596), .A(n1597), .Z(n1594) );
  XNOR U2109 ( .A(b[137]), .B(n1595), .Z(n1596) );
  XNOR U2110 ( .A(b[137]), .B(n1597), .Z(c[137]) );
  XOR U2111 ( .A(n1598), .B(n1599), .Z(n1595) );
  ANDN U2112 ( .B(n1600), .A(n1601), .Z(n1598) );
  XNOR U2113 ( .A(b[136]), .B(n1599), .Z(n1600) );
  XNOR U2114 ( .A(b[136]), .B(n1601), .Z(c[136]) );
  XOR U2115 ( .A(n1602), .B(n1603), .Z(n1599) );
  ANDN U2116 ( .B(n1604), .A(n1605), .Z(n1602) );
  XNOR U2117 ( .A(b[135]), .B(n1603), .Z(n1604) );
  XNOR U2118 ( .A(b[135]), .B(n1605), .Z(c[135]) );
  XOR U2119 ( .A(n1606), .B(n1607), .Z(n1603) );
  ANDN U2120 ( .B(n1608), .A(n1609), .Z(n1606) );
  XNOR U2121 ( .A(b[134]), .B(n1607), .Z(n1608) );
  XNOR U2122 ( .A(b[134]), .B(n1609), .Z(c[134]) );
  XOR U2123 ( .A(n1610), .B(n1611), .Z(n1607) );
  ANDN U2124 ( .B(n1612), .A(n1613), .Z(n1610) );
  XNOR U2125 ( .A(b[133]), .B(n1611), .Z(n1612) );
  XNOR U2126 ( .A(b[133]), .B(n1613), .Z(c[133]) );
  XOR U2127 ( .A(n1614), .B(n1615), .Z(n1611) );
  ANDN U2128 ( .B(n1616), .A(n1617), .Z(n1614) );
  XNOR U2129 ( .A(b[132]), .B(n1615), .Z(n1616) );
  XNOR U2130 ( .A(b[132]), .B(n1617), .Z(c[132]) );
  XOR U2131 ( .A(n1618), .B(n1619), .Z(n1615) );
  ANDN U2132 ( .B(n1620), .A(n1621), .Z(n1618) );
  XNOR U2133 ( .A(b[131]), .B(n1619), .Z(n1620) );
  XNOR U2134 ( .A(b[131]), .B(n1621), .Z(c[131]) );
  XOR U2135 ( .A(n1622), .B(n1623), .Z(n1619) );
  ANDN U2136 ( .B(n1624), .A(n1625), .Z(n1622) );
  XNOR U2137 ( .A(b[130]), .B(n1623), .Z(n1624) );
  XNOR U2138 ( .A(b[130]), .B(n1625), .Z(c[130]) );
  XOR U2139 ( .A(n1626), .B(n1627), .Z(n1623) );
  ANDN U2140 ( .B(n1628), .A(n1629), .Z(n1626) );
  XNOR U2141 ( .A(b[129]), .B(n1627), .Z(n1628) );
  XNOR U2142 ( .A(b[12]), .B(n1630), .Z(c[12]) );
  XNOR U2143 ( .A(b[129]), .B(n1629), .Z(c[129]) );
  XOR U2144 ( .A(n1631), .B(n1632), .Z(n1627) );
  ANDN U2145 ( .B(n1633), .A(n1634), .Z(n1631) );
  XNOR U2146 ( .A(b[128]), .B(n1632), .Z(n1633) );
  XNOR U2147 ( .A(b[128]), .B(n1634), .Z(c[128]) );
  XOR U2148 ( .A(n1635), .B(n1636), .Z(n1632) );
  ANDN U2149 ( .B(n1637), .A(n1638), .Z(n1635) );
  XNOR U2150 ( .A(b[127]), .B(n1636), .Z(n1637) );
  XNOR U2151 ( .A(b[127]), .B(n1638), .Z(c[127]) );
  XOR U2152 ( .A(n1639), .B(n1640), .Z(n1636) );
  ANDN U2153 ( .B(n1641), .A(n1642), .Z(n1639) );
  XNOR U2154 ( .A(b[126]), .B(n1640), .Z(n1641) );
  XNOR U2155 ( .A(b[126]), .B(n1642), .Z(c[126]) );
  XOR U2156 ( .A(n1643), .B(n1644), .Z(n1640) );
  ANDN U2157 ( .B(n1645), .A(n1646), .Z(n1643) );
  XNOR U2158 ( .A(b[125]), .B(n1644), .Z(n1645) );
  XNOR U2159 ( .A(b[125]), .B(n1646), .Z(c[125]) );
  XOR U2160 ( .A(n1647), .B(n1648), .Z(n1644) );
  ANDN U2161 ( .B(n1649), .A(n1650), .Z(n1647) );
  XNOR U2162 ( .A(b[124]), .B(n1648), .Z(n1649) );
  XNOR U2163 ( .A(b[124]), .B(n1650), .Z(c[124]) );
  XOR U2164 ( .A(n1651), .B(n1652), .Z(n1648) );
  ANDN U2165 ( .B(n1653), .A(n1654), .Z(n1651) );
  XNOR U2166 ( .A(b[123]), .B(n1652), .Z(n1653) );
  XNOR U2167 ( .A(b[123]), .B(n1654), .Z(c[123]) );
  XOR U2168 ( .A(n1655), .B(n1656), .Z(n1652) );
  ANDN U2169 ( .B(n1657), .A(n1658), .Z(n1655) );
  XNOR U2170 ( .A(b[122]), .B(n1656), .Z(n1657) );
  XNOR U2171 ( .A(b[122]), .B(n1658), .Z(c[122]) );
  XOR U2172 ( .A(n1659), .B(n1660), .Z(n1656) );
  ANDN U2173 ( .B(n1661), .A(n1662), .Z(n1659) );
  XNOR U2174 ( .A(b[121]), .B(n1660), .Z(n1661) );
  XNOR U2175 ( .A(b[121]), .B(n1662), .Z(c[121]) );
  XOR U2176 ( .A(n1663), .B(n1664), .Z(n1660) );
  ANDN U2177 ( .B(n1665), .A(n1666), .Z(n1663) );
  XNOR U2178 ( .A(b[120]), .B(n1664), .Z(n1665) );
  XNOR U2179 ( .A(b[120]), .B(n1666), .Z(c[120]) );
  XOR U2180 ( .A(n1667), .B(n1668), .Z(n1664) );
  ANDN U2181 ( .B(n1669), .A(n1670), .Z(n1667) );
  XNOR U2182 ( .A(b[119]), .B(n1668), .Z(n1669) );
  XNOR U2183 ( .A(b[11]), .B(n1671), .Z(c[11]) );
  XNOR U2184 ( .A(b[119]), .B(n1670), .Z(c[119]) );
  XOR U2185 ( .A(n1672), .B(n1673), .Z(n1668) );
  ANDN U2186 ( .B(n1674), .A(n1675), .Z(n1672) );
  XNOR U2187 ( .A(b[118]), .B(n1673), .Z(n1674) );
  XNOR U2188 ( .A(b[118]), .B(n1675), .Z(c[118]) );
  XOR U2189 ( .A(n1676), .B(n1677), .Z(n1673) );
  ANDN U2190 ( .B(n1678), .A(n1679), .Z(n1676) );
  XNOR U2191 ( .A(b[117]), .B(n1677), .Z(n1678) );
  XNOR U2192 ( .A(b[117]), .B(n1679), .Z(c[117]) );
  XOR U2193 ( .A(n1680), .B(n1681), .Z(n1677) );
  ANDN U2194 ( .B(n1682), .A(n1683), .Z(n1680) );
  XNOR U2195 ( .A(b[116]), .B(n1681), .Z(n1682) );
  XNOR U2196 ( .A(b[116]), .B(n1683), .Z(c[116]) );
  XOR U2197 ( .A(n1684), .B(n1685), .Z(n1681) );
  ANDN U2198 ( .B(n1686), .A(n1687), .Z(n1684) );
  XNOR U2199 ( .A(b[115]), .B(n1685), .Z(n1686) );
  XNOR U2200 ( .A(b[115]), .B(n1687), .Z(c[115]) );
  XOR U2201 ( .A(n1688), .B(n1689), .Z(n1685) );
  ANDN U2202 ( .B(n1690), .A(n1691), .Z(n1688) );
  XNOR U2203 ( .A(b[114]), .B(n1689), .Z(n1690) );
  XNOR U2204 ( .A(b[114]), .B(n1691), .Z(c[114]) );
  XOR U2205 ( .A(n1692), .B(n1693), .Z(n1689) );
  ANDN U2206 ( .B(n1694), .A(n1695), .Z(n1692) );
  XNOR U2207 ( .A(b[113]), .B(n1693), .Z(n1694) );
  XNOR U2208 ( .A(b[113]), .B(n1695), .Z(c[113]) );
  XOR U2209 ( .A(n1696), .B(n1697), .Z(n1693) );
  ANDN U2210 ( .B(n1698), .A(n1699), .Z(n1696) );
  XNOR U2211 ( .A(b[112]), .B(n1697), .Z(n1698) );
  XNOR U2212 ( .A(b[112]), .B(n1699), .Z(c[112]) );
  XOR U2213 ( .A(n1700), .B(n1701), .Z(n1697) );
  ANDN U2214 ( .B(n1702), .A(n1703), .Z(n1700) );
  XNOR U2215 ( .A(b[111]), .B(n1701), .Z(n1702) );
  XNOR U2216 ( .A(b[111]), .B(n1703), .Z(c[111]) );
  XOR U2217 ( .A(n1704), .B(n1705), .Z(n1701) );
  ANDN U2218 ( .B(n1706), .A(n1707), .Z(n1704) );
  XNOR U2219 ( .A(b[110]), .B(n1705), .Z(n1706) );
  XNOR U2220 ( .A(b[110]), .B(n1707), .Z(c[110]) );
  XOR U2221 ( .A(n1708), .B(n1709), .Z(n1705) );
  ANDN U2222 ( .B(n1710), .A(n1711), .Z(n1708) );
  XNOR U2223 ( .A(b[109]), .B(n1709), .Z(n1710) );
  XNOR U2224 ( .A(b[10]), .B(n1712), .Z(c[10]) );
  XNOR U2225 ( .A(b[109]), .B(n1711), .Z(c[109]) );
  XOR U2226 ( .A(n1713), .B(n1714), .Z(n1709) );
  ANDN U2227 ( .B(n1715), .A(n1716), .Z(n1713) );
  XNOR U2228 ( .A(b[108]), .B(n1714), .Z(n1715) );
  XNOR U2229 ( .A(b[108]), .B(n1716), .Z(c[108]) );
  XOR U2230 ( .A(n1717), .B(n1718), .Z(n1714) );
  ANDN U2231 ( .B(n1719), .A(n1720), .Z(n1717) );
  XNOR U2232 ( .A(b[107]), .B(n1718), .Z(n1719) );
  XNOR U2233 ( .A(b[107]), .B(n1720), .Z(c[107]) );
  XOR U2234 ( .A(n1721), .B(n1722), .Z(n1718) );
  ANDN U2235 ( .B(n1723), .A(n1724), .Z(n1721) );
  XNOR U2236 ( .A(b[106]), .B(n1722), .Z(n1723) );
  XNOR U2237 ( .A(b[106]), .B(n1724), .Z(c[106]) );
  XOR U2238 ( .A(n1725), .B(n1726), .Z(n1722) );
  ANDN U2239 ( .B(n1727), .A(n1728), .Z(n1725) );
  XNOR U2240 ( .A(b[105]), .B(n1726), .Z(n1727) );
  XNOR U2241 ( .A(b[105]), .B(n1728), .Z(c[105]) );
  XOR U2242 ( .A(n1729), .B(n1730), .Z(n1726) );
  ANDN U2243 ( .B(n1731), .A(n1732), .Z(n1729) );
  XNOR U2244 ( .A(b[104]), .B(n1730), .Z(n1731) );
  XNOR U2245 ( .A(b[104]), .B(n1732), .Z(c[104]) );
  XOR U2246 ( .A(n1733), .B(n1734), .Z(n1730) );
  ANDN U2247 ( .B(n1735), .A(n1736), .Z(n1733) );
  XNOR U2248 ( .A(b[103]), .B(n1734), .Z(n1735) );
  XNOR U2249 ( .A(b[103]), .B(n1736), .Z(c[103]) );
  XOR U2250 ( .A(n1737), .B(n1738), .Z(n1734) );
  ANDN U2251 ( .B(n1739), .A(n1740), .Z(n1737) );
  XNOR U2252 ( .A(b[102]), .B(n1738), .Z(n1739) );
  XNOR U2253 ( .A(b[102]), .B(n1740), .Z(c[102]) );
  XOR U2254 ( .A(n1741), .B(n1742), .Z(n1738) );
  ANDN U2255 ( .B(n1743), .A(n1744), .Z(n1741) );
  XNOR U2256 ( .A(b[101]), .B(n1742), .Z(n1743) );
  XNOR U2257 ( .A(b[101]), .B(n1744), .Z(c[101]) );
  XOR U2258 ( .A(n1745), .B(n1746), .Z(n1742) );
  ANDN U2259 ( .B(n1747), .A(n1748), .Z(n1745) );
  XNOR U2260 ( .A(b[100]), .B(n1746), .Z(n1747) );
  XNOR U2261 ( .A(b[100]), .B(n1748), .Z(c[100]) );
  XOR U2262 ( .A(n1749), .B(n1750), .Z(n1746) );
  ANDN U2263 ( .B(n1751), .A(n7), .Z(n1749) );
  XNOR U2264 ( .A(b[99]), .B(n1750), .Z(n1751) );
  XOR U2265 ( .A(n1752), .B(n1753), .Z(n1750) );
  ANDN U2266 ( .B(n1754), .A(n8), .Z(n1752) );
  XNOR U2267 ( .A(b[98]), .B(n1753), .Z(n1754) );
  XOR U2268 ( .A(n1755), .B(n1756), .Z(n1753) );
  ANDN U2269 ( .B(n1757), .A(n9), .Z(n1755) );
  XNOR U2270 ( .A(b[97]), .B(n1756), .Z(n1757) );
  XOR U2271 ( .A(n1758), .B(n1759), .Z(n1756) );
  ANDN U2272 ( .B(n1760), .A(n10), .Z(n1758) );
  XNOR U2273 ( .A(b[96]), .B(n1759), .Z(n1760) );
  XOR U2274 ( .A(n1761), .B(n1762), .Z(n1759) );
  ANDN U2275 ( .B(n1763), .A(n11), .Z(n1761) );
  XNOR U2276 ( .A(b[95]), .B(n1762), .Z(n1763) );
  XOR U2277 ( .A(n1764), .B(n1765), .Z(n1762) );
  ANDN U2278 ( .B(n1766), .A(n12), .Z(n1764) );
  XNOR U2279 ( .A(b[94]), .B(n1765), .Z(n1766) );
  XOR U2280 ( .A(n1767), .B(n1768), .Z(n1765) );
  ANDN U2281 ( .B(n1769), .A(n13), .Z(n1767) );
  XNOR U2282 ( .A(b[93]), .B(n1768), .Z(n1769) );
  XOR U2283 ( .A(n1770), .B(n1771), .Z(n1768) );
  ANDN U2284 ( .B(n1772), .A(n14), .Z(n1770) );
  XNOR U2285 ( .A(b[92]), .B(n1771), .Z(n1772) );
  XOR U2286 ( .A(n1773), .B(n1774), .Z(n1771) );
  ANDN U2287 ( .B(n1775), .A(n15), .Z(n1773) );
  XNOR U2288 ( .A(b[91]), .B(n1774), .Z(n1775) );
  XOR U2289 ( .A(n1776), .B(n1777), .Z(n1774) );
  ANDN U2290 ( .B(n1778), .A(n16), .Z(n1776) );
  XNOR U2291 ( .A(b[90]), .B(n1777), .Z(n1778) );
  XOR U2292 ( .A(n1779), .B(n1780), .Z(n1777) );
  ANDN U2293 ( .B(n1781), .A(n18), .Z(n1779) );
  XNOR U2294 ( .A(b[89]), .B(n1780), .Z(n1781) );
  XOR U2295 ( .A(n1782), .B(n1783), .Z(n1780) );
  ANDN U2296 ( .B(n1784), .A(n19), .Z(n1782) );
  XNOR U2297 ( .A(b[88]), .B(n1783), .Z(n1784) );
  XOR U2298 ( .A(n1785), .B(n1786), .Z(n1783) );
  ANDN U2299 ( .B(n1787), .A(n20), .Z(n1785) );
  XNOR U2300 ( .A(b[87]), .B(n1786), .Z(n1787) );
  XOR U2301 ( .A(n1788), .B(n1789), .Z(n1786) );
  ANDN U2302 ( .B(n1790), .A(n21), .Z(n1788) );
  XNOR U2303 ( .A(b[86]), .B(n1789), .Z(n1790) );
  XOR U2304 ( .A(n1791), .B(n1792), .Z(n1789) );
  ANDN U2305 ( .B(n1793), .A(n22), .Z(n1791) );
  XNOR U2306 ( .A(b[85]), .B(n1792), .Z(n1793) );
  XOR U2307 ( .A(n1794), .B(n1795), .Z(n1792) );
  ANDN U2308 ( .B(n1796), .A(n23), .Z(n1794) );
  XNOR U2309 ( .A(b[84]), .B(n1795), .Z(n1796) );
  XOR U2310 ( .A(n1797), .B(n1798), .Z(n1795) );
  ANDN U2311 ( .B(n1799), .A(n24), .Z(n1797) );
  XNOR U2312 ( .A(b[83]), .B(n1798), .Z(n1799) );
  XOR U2313 ( .A(n1800), .B(n1801), .Z(n1798) );
  ANDN U2314 ( .B(n1802), .A(n25), .Z(n1800) );
  XNOR U2315 ( .A(b[82]), .B(n1801), .Z(n1802) );
  XOR U2316 ( .A(n1803), .B(n1804), .Z(n1801) );
  ANDN U2317 ( .B(n1805), .A(n26), .Z(n1803) );
  XNOR U2318 ( .A(b[81]), .B(n1804), .Z(n1805) );
  XOR U2319 ( .A(n1806), .B(n1807), .Z(n1804) );
  ANDN U2320 ( .B(n1808), .A(n27), .Z(n1806) );
  XNOR U2321 ( .A(b[80]), .B(n1807), .Z(n1808) );
  XOR U2322 ( .A(n1809), .B(n1810), .Z(n1807) );
  ANDN U2323 ( .B(n1811), .A(n29), .Z(n1809) );
  XNOR U2324 ( .A(b[79]), .B(n1810), .Z(n1811) );
  XOR U2325 ( .A(n1812), .B(n1813), .Z(n1810) );
  ANDN U2326 ( .B(n1814), .A(n30), .Z(n1812) );
  XNOR U2327 ( .A(b[78]), .B(n1813), .Z(n1814) );
  XOR U2328 ( .A(n1815), .B(n1816), .Z(n1813) );
  ANDN U2329 ( .B(n1817), .A(n31), .Z(n1815) );
  XNOR U2330 ( .A(b[77]), .B(n1816), .Z(n1817) );
  XOR U2331 ( .A(n1818), .B(n1819), .Z(n1816) );
  ANDN U2332 ( .B(n1820), .A(n32), .Z(n1818) );
  XNOR U2333 ( .A(b[76]), .B(n1819), .Z(n1820) );
  XOR U2334 ( .A(n1821), .B(n1822), .Z(n1819) );
  ANDN U2335 ( .B(n1823), .A(n33), .Z(n1821) );
  XNOR U2336 ( .A(b[75]), .B(n1822), .Z(n1823) );
  XOR U2337 ( .A(n1824), .B(n1825), .Z(n1822) );
  ANDN U2338 ( .B(n1826), .A(n34), .Z(n1824) );
  XNOR U2339 ( .A(b[74]), .B(n1825), .Z(n1826) );
  XOR U2340 ( .A(n1827), .B(n1828), .Z(n1825) );
  ANDN U2341 ( .B(n1829), .A(n35), .Z(n1827) );
  XNOR U2342 ( .A(b[73]), .B(n1828), .Z(n1829) );
  XOR U2343 ( .A(n1830), .B(n1831), .Z(n1828) );
  ANDN U2344 ( .B(n1832), .A(n36), .Z(n1830) );
  XNOR U2345 ( .A(b[72]), .B(n1831), .Z(n1832) );
  XOR U2346 ( .A(n1833), .B(n1834), .Z(n1831) );
  ANDN U2347 ( .B(n1835), .A(n37), .Z(n1833) );
  XNOR U2348 ( .A(b[71]), .B(n1834), .Z(n1835) );
  XOR U2349 ( .A(n1836), .B(n1837), .Z(n1834) );
  ANDN U2350 ( .B(n1838), .A(n38), .Z(n1836) );
  XNOR U2351 ( .A(b[70]), .B(n1837), .Z(n1838) );
  XOR U2352 ( .A(n1839), .B(n1840), .Z(n1837) );
  ANDN U2353 ( .B(n1841), .A(n40), .Z(n1839) );
  XNOR U2354 ( .A(b[69]), .B(n1840), .Z(n1841) );
  XOR U2355 ( .A(n1842), .B(n1843), .Z(n1840) );
  ANDN U2356 ( .B(n1844), .A(n41), .Z(n1842) );
  XNOR U2357 ( .A(b[68]), .B(n1843), .Z(n1844) );
  XOR U2358 ( .A(n1845), .B(n1846), .Z(n1843) );
  ANDN U2359 ( .B(n1847), .A(n42), .Z(n1845) );
  XNOR U2360 ( .A(b[67]), .B(n1846), .Z(n1847) );
  XOR U2361 ( .A(n1848), .B(n1849), .Z(n1846) );
  ANDN U2362 ( .B(n1850), .A(n43), .Z(n1848) );
  XNOR U2363 ( .A(b[66]), .B(n1849), .Z(n1850) );
  XOR U2364 ( .A(n1851), .B(n1852), .Z(n1849) );
  ANDN U2365 ( .B(n1853), .A(n44), .Z(n1851) );
  XNOR U2366 ( .A(b[65]), .B(n1852), .Z(n1853) );
  XOR U2367 ( .A(n1854), .B(n1855), .Z(n1852) );
  ANDN U2368 ( .B(n1856), .A(n45), .Z(n1854) );
  XNOR U2369 ( .A(b[64]), .B(n1855), .Z(n1856) );
  XOR U2370 ( .A(n1857), .B(n1858), .Z(n1855) );
  ANDN U2371 ( .B(n1859), .A(n46), .Z(n1857) );
  XNOR U2372 ( .A(b[63]), .B(n1858), .Z(n1859) );
  XOR U2373 ( .A(n1860), .B(n1861), .Z(n1858) );
  ANDN U2374 ( .B(n1862), .A(n47), .Z(n1860) );
  XNOR U2375 ( .A(b[62]), .B(n1861), .Z(n1862) );
  XOR U2376 ( .A(n1863), .B(n1864), .Z(n1861) );
  ANDN U2377 ( .B(n1865), .A(n48), .Z(n1863) );
  XNOR U2378 ( .A(b[61]), .B(n1864), .Z(n1865) );
  XOR U2379 ( .A(n1866), .B(n1867), .Z(n1864) );
  ANDN U2380 ( .B(n1868), .A(n49), .Z(n1866) );
  XNOR U2381 ( .A(b[60]), .B(n1867), .Z(n1868) );
  XOR U2382 ( .A(n1869), .B(n1870), .Z(n1867) );
  ANDN U2383 ( .B(n1871), .A(n51), .Z(n1869) );
  XNOR U2384 ( .A(b[59]), .B(n1870), .Z(n1871) );
  XOR U2385 ( .A(n1872), .B(n1873), .Z(n1870) );
  ANDN U2386 ( .B(n1874), .A(n52), .Z(n1872) );
  XNOR U2387 ( .A(b[58]), .B(n1873), .Z(n1874) );
  XOR U2388 ( .A(n1875), .B(n1876), .Z(n1873) );
  ANDN U2389 ( .B(n1877), .A(n53), .Z(n1875) );
  XNOR U2390 ( .A(b[57]), .B(n1876), .Z(n1877) );
  XOR U2391 ( .A(n1878), .B(n1879), .Z(n1876) );
  ANDN U2392 ( .B(n1880), .A(n54), .Z(n1878) );
  XNOR U2393 ( .A(b[56]), .B(n1879), .Z(n1880) );
  XOR U2394 ( .A(n1881), .B(n1882), .Z(n1879) );
  ANDN U2395 ( .B(n1883), .A(n55), .Z(n1881) );
  XNOR U2396 ( .A(b[55]), .B(n1882), .Z(n1883) );
  XOR U2397 ( .A(n1884), .B(n1885), .Z(n1882) );
  ANDN U2398 ( .B(n1886), .A(n56), .Z(n1884) );
  XNOR U2399 ( .A(b[54]), .B(n1885), .Z(n1886) );
  XOR U2400 ( .A(n1887), .B(n1888), .Z(n1885) );
  ANDN U2401 ( .B(n1889), .A(n57), .Z(n1887) );
  XNOR U2402 ( .A(b[53]), .B(n1888), .Z(n1889) );
  XOR U2403 ( .A(n1890), .B(n1891), .Z(n1888) );
  ANDN U2404 ( .B(n1892), .A(n58), .Z(n1890) );
  XNOR U2405 ( .A(b[52]), .B(n1891), .Z(n1892) );
  XOR U2406 ( .A(n1893), .B(n1894), .Z(n1891) );
  ANDN U2407 ( .B(n1895), .A(n59), .Z(n1893) );
  XNOR U2408 ( .A(b[51]), .B(n1894), .Z(n1895) );
  XOR U2409 ( .A(n1896), .B(n1897), .Z(n1894) );
  ANDN U2410 ( .B(n1898), .A(n68), .Z(n1896) );
  XNOR U2411 ( .A(b[50]), .B(n1897), .Z(n1898) );
  XOR U2412 ( .A(n1899), .B(n1900), .Z(n1897) );
  ANDN U2413 ( .B(n1901), .A(n110), .Z(n1899) );
  XNOR U2414 ( .A(b[49]), .B(n1900), .Z(n1901) );
  XOR U2415 ( .A(n1902), .B(n1903), .Z(n1900) );
  ANDN U2416 ( .B(n1904), .A(n151), .Z(n1902) );
  XNOR U2417 ( .A(b[48]), .B(n1903), .Z(n1904) );
  XOR U2418 ( .A(n1905), .B(n1906), .Z(n1903) );
  ANDN U2419 ( .B(n1907), .A(n192), .Z(n1905) );
  XNOR U2420 ( .A(b[47]), .B(n1906), .Z(n1907) );
  XOR U2421 ( .A(n1908), .B(n1909), .Z(n1906) );
  ANDN U2422 ( .B(n1910), .A(n233), .Z(n1908) );
  XNOR U2423 ( .A(b[46]), .B(n1909), .Z(n1910) );
  XOR U2424 ( .A(n1911), .B(n1912), .Z(n1909) );
  ANDN U2425 ( .B(n1913), .A(n274), .Z(n1911) );
  XNOR U2426 ( .A(b[45]), .B(n1912), .Z(n1913) );
  XOR U2427 ( .A(n1914), .B(n1915), .Z(n1912) );
  ANDN U2428 ( .B(n1916), .A(n315), .Z(n1914) );
  XNOR U2429 ( .A(b[44]), .B(n1915), .Z(n1916) );
  XOR U2430 ( .A(n1917), .B(n1918), .Z(n1915) );
  ANDN U2431 ( .B(n1919), .A(n356), .Z(n1917) );
  XNOR U2432 ( .A(b[43]), .B(n1918), .Z(n1919) );
  XOR U2433 ( .A(n1920), .B(n1921), .Z(n1918) );
  ANDN U2434 ( .B(n1922), .A(n397), .Z(n1920) );
  XNOR U2435 ( .A(b[42]), .B(n1921), .Z(n1922) );
  XOR U2436 ( .A(n1923), .B(n1924), .Z(n1921) );
  ANDN U2437 ( .B(n1925), .A(n438), .Z(n1923) );
  XNOR U2438 ( .A(b[41]), .B(n1924), .Z(n1925) );
  XOR U2439 ( .A(n1926), .B(n1927), .Z(n1924) );
  ANDN U2440 ( .B(n1928), .A(n479), .Z(n1926) );
  XNOR U2441 ( .A(b[40]), .B(n1927), .Z(n1928) );
  XOR U2442 ( .A(n1929), .B(n1930), .Z(n1927) );
  ANDN U2443 ( .B(n1931), .A(n521), .Z(n1929) );
  XNOR U2444 ( .A(b[39]), .B(n1930), .Z(n1931) );
  XOR U2445 ( .A(n1932), .B(n1933), .Z(n1930) );
  ANDN U2446 ( .B(n1934), .A(n562), .Z(n1932) );
  XNOR U2447 ( .A(b[38]), .B(n1933), .Z(n1934) );
  XOR U2448 ( .A(n1935), .B(n1936), .Z(n1933) );
  ANDN U2449 ( .B(n1937), .A(n603), .Z(n1935) );
  XNOR U2450 ( .A(b[37]), .B(n1936), .Z(n1937) );
  XOR U2451 ( .A(n1938), .B(n1939), .Z(n1936) );
  ANDN U2452 ( .B(n1940), .A(n644), .Z(n1938) );
  XNOR U2453 ( .A(b[36]), .B(n1939), .Z(n1940) );
  XOR U2454 ( .A(n1941), .B(n1942), .Z(n1939) );
  ANDN U2455 ( .B(n1943), .A(n685), .Z(n1941) );
  XNOR U2456 ( .A(b[35]), .B(n1942), .Z(n1943) );
  XOR U2457 ( .A(n1944), .B(n1945), .Z(n1942) );
  ANDN U2458 ( .B(n1946), .A(n726), .Z(n1944) );
  XNOR U2459 ( .A(b[34]), .B(n1945), .Z(n1946) );
  XOR U2460 ( .A(n1947), .B(n1948), .Z(n1945) );
  ANDN U2461 ( .B(n1949), .A(n767), .Z(n1947) );
  XNOR U2462 ( .A(b[33]), .B(n1948), .Z(n1949) );
  XOR U2463 ( .A(n1950), .B(n1951), .Z(n1948) );
  ANDN U2464 ( .B(n1952), .A(n808), .Z(n1950) );
  XNOR U2465 ( .A(b[32]), .B(n1951), .Z(n1952) );
  XOR U2466 ( .A(n1953), .B(n1954), .Z(n1951) );
  ANDN U2467 ( .B(n1955), .A(n849), .Z(n1953) );
  XNOR U2468 ( .A(b[31]), .B(n1954), .Z(n1955) );
  XOR U2469 ( .A(n1956), .B(n1957), .Z(n1954) );
  ANDN U2470 ( .B(n1958), .A(n890), .Z(n1956) );
  XNOR U2471 ( .A(b[30]), .B(n1957), .Z(n1958) );
  XOR U2472 ( .A(n1959), .B(n1960), .Z(n1957) );
  ANDN U2473 ( .B(n1961), .A(n932), .Z(n1959) );
  XNOR U2474 ( .A(b[29]), .B(n1960), .Z(n1961) );
  XOR U2475 ( .A(n1962), .B(n1963), .Z(n1960) );
  ANDN U2476 ( .B(n1964), .A(n973), .Z(n1962) );
  XNOR U2477 ( .A(b[28]), .B(n1963), .Z(n1964) );
  XOR U2478 ( .A(n1965), .B(n1966), .Z(n1963) );
  ANDN U2479 ( .B(n1967), .A(n1014), .Z(n1965) );
  XNOR U2480 ( .A(b[27]), .B(n1966), .Z(n1967) );
  XOR U2481 ( .A(n1968), .B(n1969), .Z(n1966) );
  ANDN U2482 ( .B(n1970), .A(n1055), .Z(n1968) );
  XNOR U2483 ( .A(b[26]), .B(n1969), .Z(n1970) );
  XOR U2484 ( .A(n1971), .B(n1972), .Z(n1969) );
  ANDN U2485 ( .B(n1973), .A(n1096), .Z(n1971) );
  XNOR U2486 ( .A(b[25]), .B(n1972), .Z(n1973) );
  XOR U2487 ( .A(n1974), .B(n1975), .Z(n1972) );
  ANDN U2488 ( .B(n1976), .A(n1137), .Z(n1974) );
  XNOR U2489 ( .A(b[24]), .B(n1975), .Z(n1976) );
  XOR U2490 ( .A(n1977), .B(n1978), .Z(n1975) );
  ANDN U2491 ( .B(n1979), .A(n1178), .Z(n1977) );
  XNOR U2492 ( .A(b[23]), .B(n1978), .Z(n1979) );
  XOR U2493 ( .A(n1980), .B(n1981), .Z(n1978) );
  ANDN U2494 ( .B(n1982), .A(n1219), .Z(n1980) );
  XNOR U2495 ( .A(b[22]), .B(n1981), .Z(n1982) );
  XOR U2496 ( .A(n1983), .B(n1984), .Z(n1981) );
  ANDN U2497 ( .B(n1985), .A(n1260), .Z(n1983) );
  XNOR U2498 ( .A(b[21]), .B(n1984), .Z(n1985) );
  XOR U2499 ( .A(n1986), .B(n1987), .Z(n1984) );
  ANDN U2500 ( .B(n1988), .A(n1301), .Z(n1986) );
  XNOR U2501 ( .A(b[20]), .B(n1987), .Z(n1988) );
  XOR U2502 ( .A(n1989), .B(n1990), .Z(n1987) );
  ANDN U2503 ( .B(n1991), .A(n1343), .Z(n1989) );
  XNOR U2504 ( .A(b[19]), .B(n1990), .Z(n1991) );
  XOR U2505 ( .A(n1992), .B(n1993), .Z(n1990) );
  ANDN U2506 ( .B(n1994), .A(n1384), .Z(n1992) );
  XNOR U2507 ( .A(b[18]), .B(n1993), .Z(n1994) );
  XOR U2508 ( .A(n1995), .B(n1996), .Z(n1993) );
  ANDN U2509 ( .B(n1997), .A(n1425), .Z(n1995) );
  XNOR U2510 ( .A(b[17]), .B(n1996), .Z(n1997) );
  XOR U2511 ( .A(n1998), .B(n1999), .Z(n1996) );
  ANDN U2512 ( .B(n2000), .A(n1466), .Z(n1998) );
  XNOR U2513 ( .A(b[16]), .B(n1999), .Z(n2000) );
  XOR U2514 ( .A(n2001), .B(n2002), .Z(n1999) );
  ANDN U2515 ( .B(n2003), .A(n1507), .Z(n2001) );
  XNOR U2516 ( .A(b[15]), .B(n2002), .Z(n2003) );
  XOR U2517 ( .A(n2004), .B(n2005), .Z(n2002) );
  ANDN U2518 ( .B(n2006), .A(n1548), .Z(n2004) );
  XNOR U2519 ( .A(b[14]), .B(n2005), .Z(n2006) );
  XOR U2520 ( .A(n2007), .B(n2008), .Z(n2005) );
  ANDN U2521 ( .B(n2009), .A(n1589), .Z(n2007) );
  XNOR U2522 ( .A(b[13]), .B(n2008), .Z(n2009) );
  XOR U2523 ( .A(n2010), .B(n2011), .Z(n2008) );
  ANDN U2524 ( .B(n2012), .A(n1630), .Z(n2010) );
  XNOR U2525 ( .A(b[12]), .B(n2011), .Z(n2012) );
  XOR U2526 ( .A(n2013), .B(n2014), .Z(n2011) );
  ANDN U2527 ( .B(n2015), .A(n1671), .Z(n2013) );
  XNOR U2528 ( .A(b[11]), .B(n2014), .Z(n2015) );
  XOR U2529 ( .A(n2016), .B(n2017), .Z(n2014) );
  ANDN U2530 ( .B(n2018), .A(n1712), .Z(n2016) );
  XNOR U2531 ( .A(b[10]), .B(n2017), .Z(n2018) );
  XOR U2532 ( .A(n2019), .B(n2020), .Z(n2017) );
  ANDN U2533 ( .B(n2021), .A(n6), .Z(n2019) );
  XNOR U2534 ( .A(b[9]), .B(n2020), .Z(n2021) );
  XOR U2535 ( .A(n2022), .B(n2023), .Z(n2020) );
  ANDN U2536 ( .B(n2024), .A(n17), .Z(n2022) );
  XNOR U2537 ( .A(b[8]), .B(n2023), .Z(n2024) );
  XOR U2538 ( .A(n2025), .B(n2026), .Z(n2023) );
  ANDN U2539 ( .B(n2027), .A(n28), .Z(n2025) );
  XNOR U2540 ( .A(b[7]), .B(n2026), .Z(n2027) );
  XOR U2541 ( .A(n2028), .B(n2029), .Z(n2026) );
  ANDN U2542 ( .B(n2030), .A(n39), .Z(n2028) );
  XNOR U2543 ( .A(b[6]), .B(n2029), .Z(n2030) );
  XOR U2544 ( .A(n2031), .B(n2032), .Z(n2029) );
  ANDN U2545 ( .B(n2033), .A(n50), .Z(n2031) );
  XNOR U2546 ( .A(b[5]), .B(n2032), .Z(n2033) );
  XOR U2547 ( .A(n2034), .B(n2035), .Z(n2032) );
  ANDN U2548 ( .B(n2036), .A(n109), .Z(n2034) );
  XNOR U2549 ( .A(b[4]), .B(n2035), .Z(n2036) );
  XOR U2550 ( .A(n2037), .B(n2038), .Z(n2035) );
  ANDN U2551 ( .B(n2039), .A(n520), .Z(n2037) );
  XNOR U2552 ( .A(b[3]), .B(n2038), .Z(n2039) );
  XOR U2553 ( .A(n2040), .B(n2041), .Z(n2038) );
  ANDN U2554 ( .B(n2042), .A(n931), .Z(n2040) );
  XNOR U2555 ( .A(b[2]), .B(n2041), .Z(n2042) );
  XOR U2556 ( .A(n2043), .B(n2044), .Z(n2041) );
  ANDN U2557 ( .B(n2045), .A(n1342), .Z(n2043) );
  XNOR U2558 ( .A(b[1]), .B(n2044), .Z(n2045) );
  XOR U2559 ( .A(carry_on), .B(n2046), .Z(n2044) );
  NANDN U2560 ( .A(n2047), .B(n2048), .Z(n2046) );
  XOR U2561 ( .A(carry_on), .B(b[0]), .Z(n2048) );
  XNOR U2562 ( .A(b[0]), .B(n2047), .Z(c[0]) );
  XNOR U2563 ( .A(a[0]), .B(carry_on), .Z(n2047) );
endmodule

