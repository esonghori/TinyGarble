
module hamming_N1600_CC64 ( clk, rst, x, y, o );
  input [24:0] x;
  input [24:0] y;
  output [10:0] o;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154;
  wire   [10:0] oglobal;

  DFF \oglobal_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .Q(oglobal[10]) );
  DFF \oglobal_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .Q(oglobal[9]) );
  DFF \oglobal_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .Q(oglobal[8]) );
  DFF \oglobal_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .Q(oglobal[7]) );
  DFF \oglobal_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .Q(oglobal[6]) );
  DFF \oglobal_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .Q(oglobal[5]) );
  DFF \oglobal_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .Q(oglobal[4]) );
  DFF \oglobal_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .Q(oglobal[3]) );
  DFF \oglobal_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .Q(oglobal[2]) );
  DFF \oglobal_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .Q(oglobal[1]) );
  DFF \oglobal_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .Q(oglobal[0]) );
  XOR U28 ( .A(n86), .B(n87), .Z(n103) );
  XOR U29 ( .A(n98), .B(n99), .Z(n110) );
  XNOR U30 ( .A(n49), .B(n50), .Z(n42) );
  XOR U31 ( .A(n122), .B(n123), .Z(n117) );
  XNOR U32 ( .A(x[10]), .B(y[10]), .Z(n25) );
  XNOR U33 ( .A(x[8]), .B(y[8]), .Z(n23) );
  XNOR U34 ( .A(x[6]), .B(y[6]), .Z(n22) );
  XNOR U35 ( .A(n23), .B(n22), .Z(n24) );
  XNOR U36 ( .A(n25), .B(n24), .Z(n68) );
  XNOR U37 ( .A(x[16]), .B(y[16]), .Z(n19) );
  XNOR U38 ( .A(x[14]), .B(y[14]), .Z(n17) );
  XNOR U39 ( .A(x[12]), .B(y[12]), .Z(n16) );
  XNOR U40 ( .A(n17), .B(n16), .Z(n18) );
  XNOR U41 ( .A(n19), .B(n18), .Z(n66) );
  XNOR U42 ( .A(x[22]), .B(y[22]), .Z(n65) );
  XNOR U43 ( .A(n66), .B(n65), .Z(n67) );
  XNOR U44 ( .A(n68), .B(n67), .Z(n3) );
  XNOR U45 ( .A(x[15]), .B(y[15]), .Z(n50) );
  XNOR U46 ( .A(x[19]), .B(y[19]), .Z(n48) );
  XNOR U47 ( .A(n48), .B(oglobal[0]), .Z(n49) );
  IV U48 ( .A(n42), .Z(n41) );
  XNOR U49 ( .A(x[23]), .B(y[23]), .Z(n9) );
  XNOR U50 ( .A(x[21]), .B(y[21]), .Z(n8) );
  XNOR U51 ( .A(n9), .B(n8), .Z(n56) );
  XNOR U52 ( .A(x[13]), .B(y[13]), .Z(n54) );
  XNOR U53 ( .A(x[17]), .B(y[17]), .Z(n53) );
  XNOR U54 ( .A(n54), .B(n53), .Z(n55) );
  XNOR U55 ( .A(n56), .B(n55), .Z(n44) );
  XNOR U56 ( .A(x[7]), .B(y[7]), .Z(n62) );
  XNOR U57 ( .A(x[9]), .B(y[9]), .Z(n60) );
  XNOR U58 ( .A(x[11]), .B(y[11]), .Z(n59) );
  XNOR U59 ( .A(n60), .B(n59), .Z(n61) );
  XNOR U60 ( .A(n62), .B(n61), .Z(n40) );
  IV U61 ( .A(n40), .Z(n43) );
  XOR U62 ( .A(n44), .B(n43), .Z(n1) );
  XOR U63 ( .A(n41), .B(n1), .Z(n2) );
  XOR U64 ( .A(n3), .B(n2), .Z(n5) );
  XNOR U65 ( .A(x[20]), .B(y[20]), .Z(n13) );
  XNOR U66 ( .A(x[24]), .B(y[24]), .Z(n11) );
  XNOR U67 ( .A(x[18]), .B(y[18]), .Z(n10) );
  XNOR U68 ( .A(n11), .B(n10), .Z(n12) );
  XNOR U69 ( .A(n13), .B(n12), .Z(n73) );
  XNOR U70 ( .A(x[1]), .B(y[1]), .Z(n31) );
  XNOR U71 ( .A(x[5]), .B(y[5]), .Z(n29) );
  XNOR U72 ( .A(x[3]), .B(y[3]), .Z(n28) );
  XNOR U73 ( .A(n29), .B(n28), .Z(n30) );
  XNOR U74 ( .A(n31), .B(n30), .Z(n71) );
  XNOR U75 ( .A(x[4]), .B(y[4]), .Z(n37) );
  XNOR U76 ( .A(x[2]), .B(y[2]), .Z(n35) );
  XNOR U77 ( .A(x[0]), .B(y[0]), .Z(n34) );
  XNOR U78 ( .A(n35), .B(n34), .Z(n36) );
  XNOR U79 ( .A(n37), .B(n36), .Z(n72) );
  XNOR U80 ( .A(n71), .B(n72), .Z(n74) );
  XNOR U81 ( .A(n73), .B(n74), .Z(n4) );
  XOR U82 ( .A(n5), .B(n4), .Z(o[0]) );
  NANDN U83 ( .A(n3), .B(n2), .Z(n7) );
  OR U84 ( .A(n5), .B(n4), .Z(n6) );
  NAND U85 ( .A(n7), .B(n6), .Z(n77) );
  OR U86 ( .A(n9), .B(n8), .Z(n83) );
  XNOR U87 ( .A(oglobal[1]), .B(n83), .Z(n93) );
  OR U88 ( .A(n11), .B(n10), .Z(n15) );
  OR U89 ( .A(n13), .B(n12), .Z(n14) );
  NAND U90 ( .A(n15), .B(n14), .Z(n91) );
  OR U91 ( .A(n17), .B(n16), .Z(n21) );
  OR U92 ( .A(n19), .B(n18), .Z(n20) );
  NAND U93 ( .A(n21), .B(n20), .Z(n90) );
  XOR U94 ( .A(n91), .B(n90), .Z(n92) );
  XOR U95 ( .A(n93), .B(n92), .Z(n105) );
  OR U96 ( .A(n23), .B(n22), .Z(n27) );
  OR U97 ( .A(n25), .B(n24), .Z(n26) );
  NAND U98 ( .A(n27), .B(n26), .Z(n85) );
  OR U99 ( .A(n29), .B(n28), .Z(n33) );
  OR U100 ( .A(n31), .B(n30), .Z(n32) );
  NAND U101 ( .A(n33), .B(n32), .Z(n84) );
  XOR U102 ( .A(n85), .B(n84), .Z(n86) );
  OR U103 ( .A(n35), .B(n34), .Z(n39) );
  OR U104 ( .A(n37), .B(n36), .Z(n38) );
  NAND U105 ( .A(n39), .B(n38), .Z(n87) );
  NAND U106 ( .A(n41), .B(n40), .Z(n47) );
  AND U107 ( .A(n43), .B(n42), .Z(n45) );
  NANDN U108 ( .A(n45), .B(n44), .Z(n46) );
  NAND U109 ( .A(n47), .B(n46), .Z(n102) );
  XOR U110 ( .A(n103), .B(n102), .Z(n104) );
  XOR U111 ( .A(n105), .B(n104), .Z(n78) );
  XNOR U112 ( .A(n77), .B(n78), .Z(n79) );
  NANDN U113 ( .A(n48), .B(oglobal[0]), .Z(n52) );
  NANDN U114 ( .A(n50), .B(n49), .Z(n51) );
  AND U115 ( .A(n52), .B(n51), .Z(n99) );
  OR U116 ( .A(n54), .B(n53), .Z(n58) );
  OR U117 ( .A(n56), .B(n55), .Z(n57) );
  AND U118 ( .A(n58), .B(n57), .Z(n96) );
  OR U119 ( .A(n60), .B(n59), .Z(n64) );
  OR U120 ( .A(n62), .B(n61), .Z(n63) );
  AND U121 ( .A(n64), .B(n63), .Z(n97) );
  XOR U122 ( .A(n96), .B(n97), .Z(n98) );
  OR U123 ( .A(n66), .B(n65), .Z(n70) );
  OR U124 ( .A(n68), .B(n67), .Z(n69) );
  NAND U125 ( .A(n70), .B(n69), .Z(n109) );
  NAND U126 ( .A(n72), .B(n71), .Z(n76) );
  NANDN U127 ( .A(n74), .B(n73), .Z(n75) );
  AND U128 ( .A(n76), .B(n75), .Z(n108) );
  XNOR U129 ( .A(n109), .B(n108), .Z(n111) );
  XNOR U130 ( .A(n110), .B(n111), .Z(n80) );
  XNOR U131 ( .A(n79), .B(n80), .Z(o[1]) );
  NANDN U132 ( .A(n78), .B(n77), .Z(n82) );
  NANDN U133 ( .A(n80), .B(n79), .Z(n81) );
  NAND U134 ( .A(n82), .B(n81), .Z(n115) );
  NANDN U135 ( .A(n83), .B(oglobal[1]), .Z(n126) );
  XOR U136 ( .A(oglobal[2]), .B(n126), .Z(n129) );
  OR U137 ( .A(n85), .B(n84), .Z(n89) );
  NANDN U138 ( .A(n87), .B(n86), .Z(n88) );
  AND U139 ( .A(n89), .B(n88), .Z(n128) );
  OR U140 ( .A(n91), .B(n90), .Z(n95) );
  NANDN U141 ( .A(n93), .B(n92), .Z(n94) );
  AND U142 ( .A(n95), .B(n94), .Z(n127) );
  XNOR U143 ( .A(n128), .B(n127), .Z(n130) );
  XOR U144 ( .A(n129), .B(n130), .Z(n114) );
  XNOR U145 ( .A(n115), .B(n114), .Z(n116) );
  OR U146 ( .A(n97), .B(n96), .Z(n101) );
  NANDN U147 ( .A(n99), .B(n98), .Z(n100) );
  AND U148 ( .A(n101), .B(n100), .Z(n123) );
  NANDN U149 ( .A(n103), .B(n102), .Z(n107) );
  OR U150 ( .A(n105), .B(n104), .Z(n106) );
  NAND U151 ( .A(n107), .B(n106), .Z(n121) );
  OR U152 ( .A(n109), .B(n108), .Z(n113) );
  NANDN U153 ( .A(n111), .B(n110), .Z(n112) );
  NAND U154 ( .A(n113), .B(n112), .Z(n120) );
  XOR U155 ( .A(n121), .B(n120), .Z(n122) );
  XOR U156 ( .A(n116), .B(n117), .Z(o[2]) );
  NAND U157 ( .A(n115), .B(n114), .Z(n119) );
  OR U158 ( .A(n117), .B(n116), .Z(n118) );
  NAND U159 ( .A(n119), .B(n118), .Z(n133) );
  OR U160 ( .A(n121), .B(n120), .Z(n125) );
  NANDN U161 ( .A(n123), .B(n122), .Z(n124) );
  AND U162 ( .A(n125), .B(n124), .Z(n134) );
  XNOR U163 ( .A(n133), .B(n134), .Z(n135) );
  NANDN U164 ( .A(n126), .B(oglobal[2]), .Z(n139) );
  XOR U165 ( .A(oglobal[3]), .B(n139), .Z(n141) );
  OR U166 ( .A(n128), .B(n127), .Z(n132) );
  NANDN U167 ( .A(n130), .B(n129), .Z(n131) );
  NAND U168 ( .A(n132), .B(n131), .Z(n140) );
  XNOR U169 ( .A(n141), .B(n140), .Z(n136) );
  XNOR U170 ( .A(n135), .B(n136), .Z(o[3]) );
  NANDN U171 ( .A(n134), .B(n133), .Z(n138) );
  NANDN U172 ( .A(n136), .B(n135), .Z(n137) );
  NAND U173 ( .A(n138), .B(n137), .Z(n144) );
  XNOR U174 ( .A(n144), .B(oglobal[4]), .Z(n146) );
  NANDN U175 ( .A(n139), .B(oglobal[3]), .Z(n143) );
  OR U176 ( .A(n141), .B(n140), .Z(n142) );
  AND U177 ( .A(n143), .B(n142), .Z(n145) );
  XOR U178 ( .A(n146), .B(n145), .Z(o[4]) );
  NAND U179 ( .A(n144), .B(oglobal[4]), .Z(n148) );
  OR U180 ( .A(n146), .B(n145), .Z(n147) );
  AND U181 ( .A(n148), .B(n147), .Z(n149) );
  XNOR U182 ( .A(oglobal[5]), .B(n149), .Z(o[5]) );
  NANDN U183 ( .A(n149), .B(oglobal[5]), .Z(n150) );
  XNOR U184 ( .A(n150), .B(oglobal[6]), .Z(o[6]) );
  NANDN U185 ( .A(n150), .B(oglobal[6]), .Z(n151) );
  XNOR U186 ( .A(n151), .B(oglobal[7]), .Z(o[7]) );
  NANDN U187 ( .A(n151), .B(oglobal[7]), .Z(n152) );
  XNOR U188 ( .A(n152), .B(oglobal[8]), .Z(o[8]) );
  NANDN U189 ( .A(n152), .B(oglobal[8]), .Z(n153) );
  XNOR U190 ( .A(oglobal[9]), .B(n153), .Z(o[9]) );
  NANDN U191 ( .A(n153), .B(oglobal[9]), .Z(n154) );
  XNOR U192 ( .A(oglobal[10]), .B(n154), .Z(o[10]) );
endmodule

