
module sum_N1024_CC4 ( clk, rst, a, b, c );
  input [255:0] a;
  input [255:0] b;
  output [255:0] c;
  input clk, rst;
  wire   carry_on, carry_on_d, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023;

  DFF carry_on_reg ( .D(carry_on_d), .CLK(clk), .RST(rst), .Q(carry_on) );
  XOR U3 ( .A(a[0]), .B(b[0]), .Z(n1) );
  XOR U4 ( .A(n1), .B(carry_on), .Z(c[0]) );
  XOR U5 ( .A(a[1]), .B(b[1]), .Z(n5) );
  NAND U6 ( .A(a[0]), .B(b[0]), .Z(n3) );
  NAND U7 ( .A(n1), .B(carry_on), .Z(n2) );
  NAND U8 ( .A(n3), .B(n2), .Z(n4) );
  XOR U9 ( .A(n5), .B(n4), .Z(c[1]) );
  XOR U10 ( .A(a[2]), .B(b[2]), .Z(n9) );
  NAND U11 ( .A(a[1]), .B(b[1]), .Z(n7) );
  NAND U12 ( .A(n5), .B(n4), .Z(n6) );
  NAND U13 ( .A(n7), .B(n6), .Z(n8) );
  XOR U14 ( .A(n9), .B(n8), .Z(c[2]) );
  XOR U15 ( .A(a[3]), .B(b[3]), .Z(n13) );
  NAND U16 ( .A(a[2]), .B(b[2]), .Z(n11) );
  NAND U17 ( .A(n9), .B(n8), .Z(n10) );
  NAND U18 ( .A(n11), .B(n10), .Z(n12) );
  XOR U19 ( .A(n13), .B(n12), .Z(c[3]) );
  XOR U20 ( .A(a[4]), .B(b[4]), .Z(n17) );
  NAND U21 ( .A(a[3]), .B(b[3]), .Z(n15) );
  NAND U22 ( .A(n13), .B(n12), .Z(n14) );
  NAND U23 ( .A(n15), .B(n14), .Z(n16) );
  XOR U24 ( .A(n17), .B(n16), .Z(c[4]) );
  XOR U25 ( .A(a[5]), .B(b[5]), .Z(n21) );
  NAND U26 ( .A(a[4]), .B(b[4]), .Z(n19) );
  NAND U27 ( .A(n17), .B(n16), .Z(n18) );
  NAND U28 ( .A(n19), .B(n18), .Z(n20) );
  XOR U29 ( .A(n21), .B(n20), .Z(c[5]) );
  XOR U30 ( .A(a[6]), .B(b[6]), .Z(n25) );
  NAND U31 ( .A(a[5]), .B(b[5]), .Z(n23) );
  NAND U32 ( .A(n21), .B(n20), .Z(n22) );
  NAND U33 ( .A(n23), .B(n22), .Z(n24) );
  XOR U34 ( .A(n25), .B(n24), .Z(c[6]) );
  XOR U35 ( .A(a[7]), .B(b[7]), .Z(n29) );
  NAND U36 ( .A(a[6]), .B(b[6]), .Z(n27) );
  NAND U37 ( .A(n25), .B(n24), .Z(n26) );
  NAND U38 ( .A(n27), .B(n26), .Z(n28) );
  XOR U39 ( .A(n29), .B(n28), .Z(c[7]) );
  XOR U40 ( .A(a[8]), .B(b[8]), .Z(n33) );
  NAND U41 ( .A(a[7]), .B(b[7]), .Z(n31) );
  NAND U42 ( .A(n29), .B(n28), .Z(n30) );
  NAND U43 ( .A(n31), .B(n30), .Z(n32) );
  XOR U44 ( .A(n33), .B(n32), .Z(c[8]) );
  XOR U45 ( .A(a[9]), .B(b[9]), .Z(n37) );
  NAND U46 ( .A(a[8]), .B(b[8]), .Z(n35) );
  NAND U47 ( .A(n33), .B(n32), .Z(n34) );
  NAND U48 ( .A(n35), .B(n34), .Z(n36) );
  XOR U49 ( .A(n37), .B(n36), .Z(c[9]) );
  XOR U50 ( .A(a[10]), .B(b[10]), .Z(n41) );
  NAND U51 ( .A(a[9]), .B(b[9]), .Z(n39) );
  NAND U52 ( .A(n37), .B(n36), .Z(n38) );
  NAND U53 ( .A(n39), .B(n38), .Z(n40) );
  XOR U54 ( .A(n41), .B(n40), .Z(c[10]) );
  XOR U55 ( .A(a[11]), .B(b[11]), .Z(n45) );
  NAND U56 ( .A(a[10]), .B(b[10]), .Z(n43) );
  NAND U57 ( .A(n41), .B(n40), .Z(n42) );
  NAND U58 ( .A(n43), .B(n42), .Z(n44) );
  XOR U59 ( .A(n45), .B(n44), .Z(c[11]) );
  XOR U60 ( .A(a[12]), .B(b[12]), .Z(n49) );
  NAND U61 ( .A(a[11]), .B(b[11]), .Z(n47) );
  NAND U62 ( .A(n45), .B(n44), .Z(n46) );
  NAND U63 ( .A(n47), .B(n46), .Z(n48) );
  XOR U64 ( .A(n49), .B(n48), .Z(c[12]) );
  XOR U65 ( .A(a[13]), .B(b[13]), .Z(n53) );
  NAND U66 ( .A(a[12]), .B(b[12]), .Z(n51) );
  NAND U67 ( .A(n49), .B(n48), .Z(n50) );
  NAND U68 ( .A(n51), .B(n50), .Z(n52) );
  XOR U69 ( .A(n53), .B(n52), .Z(c[13]) );
  XOR U70 ( .A(a[14]), .B(b[14]), .Z(n57) );
  NAND U71 ( .A(a[13]), .B(b[13]), .Z(n55) );
  NAND U72 ( .A(n53), .B(n52), .Z(n54) );
  NAND U73 ( .A(n55), .B(n54), .Z(n56) );
  XOR U74 ( .A(n57), .B(n56), .Z(c[14]) );
  XOR U75 ( .A(a[15]), .B(b[15]), .Z(n61) );
  NAND U76 ( .A(a[14]), .B(b[14]), .Z(n59) );
  NAND U77 ( .A(n57), .B(n56), .Z(n58) );
  NAND U78 ( .A(n59), .B(n58), .Z(n60) );
  XOR U79 ( .A(n61), .B(n60), .Z(c[15]) );
  XOR U80 ( .A(a[16]), .B(b[16]), .Z(n65) );
  NAND U81 ( .A(a[15]), .B(b[15]), .Z(n63) );
  NAND U82 ( .A(n61), .B(n60), .Z(n62) );
  NAND U83 ( .A(n63), .B(n62), .Z(n64) );
  XOR U84 ( .A(n65), .B(n64), .Z(c[16]) );
  XOR U85 ( .A(a[17]), .B(b[17]), .Z(n69) );
  NAND U86 ( .A(a[16]), .B(b[16]), .Z(n67) );
  NAND U87 ( .A(n65), .B(n64), .Z(n66) );
  NAND U88 ( .A(n67), .B(n66), .Z(n68) );
  XOR U89 ( .A(n69), .B(n68), .Z(c[17]) );
  XOR U90 ( .A(a[18]), .B(b[18]), .Z(n73) );
  NAND U91 ( .A(a[17]), .B(b[17]), .Z(n71) );
  NAND U92 ( .A(n69), .B(n68), .Z(n70) );
  NAND U93 ( .A(n71), .B(n70), .Z(n72) );
  XOR U94 ( .A(n73), .B(n72), .Z(c[18]) );
  XOR U95 ( .A(a[19]), .B(b[19]), .Z(n77) );
  NAND U96 ( .A(a[18]), .B(b[18]), .Z(n75) );
  NAND U97 ( .A(n73), .B(n72), .Z(n74) );
  NAND U98 ( .A(n75), .B(n74), .Z(n76) );
  XOR U99 ( .A(n77), .B(n76), .Z(c[19]) );
  XOR U100 ( .A(a[20]), .B(b[20]), .Z(n81) );
  NAND U101 ( .A(a[19]), .B(b[19]), .Z(n79) );
  NAND U102 ( .A(n77), .B(n76), .Z(n78) );
  NAND U103 ( .A(n79), .B(n78), .Z(n80) );
  XOR U104 ( .A(n81), .B(n80), .Z(c[20]) );
  XOR U105 ( .A(a[21]), .B(b[21]), .Z(n85) );
  NAND U106 ( .A(a[20]), .B(b[20]), .Z(n83) );
  NAND U107 ( .A(n81), .B(n80), .Z(n82) );
  NAND U108 ( .A(n83), .B(n82), .Z(n84) );
  XOR U109 ( .A(n85), .B(n84), .Z(c[21]) );
  XOR U110 ( .A(a[22]), .B(b[22]), .Z(n89) );
  NAND U111 ( .A(a[21]), .B(b[21]), .Z(n87) );
  NAND U112 ( .A(n85), .B(n84), .Z(n86) );
  NAND U113 ( .A(n87), .B(n86), .Z(n88) );
  XOR U114 ( .A(n89), .B(n88), .Z(c[22]) );
  XOR U115 ( .A(a[23]), .B(b[23]), .Z(n93) );
  NAND U116 ( .A(a[22]), .B(b[22]), .Z(n91) );
  NAND U117 ( .A(n89), .B(n88), .Z(n90) );
  NAND U118 ( .A(n91), .B(n90), .Z(n92) );
  XOR U119 ( .A(n93), .B(n92), .Z(c[23]) );
  XOR U120 ( .A(a[24]), .B(b[24]), .Z(n97) );
  NAND U121 ( .A(a[23]), .B(b[23]), .Z(n95) );
  NAND U122 ( .A(n93), .B(n92), .Z(n94) );
  NAND U123 ( .A(n95), .B(n94), .Z(n96) );
  XOR U124 ( .A(n97), .B(n96), .Z(c[24]) );
  XOR U125 ( .A(a[25]), .B(b[25]), .Z(n101) );
  NAND U126 ( .A(a[24]), .B(b[24]), .Z(n99) );
  NAND U127 ( .A(n97), .B(n96), .Z(n98) );
  NAND U128 ( .A(n99), .B(n98), .Z(n100) );
  XOR U129 ( .A(n101), .B(n100), .Z(c[25]) );
  XOR U130 ( .A(a[26]), .B(b[26]), .Z(n105) );
  NAND U131 ( .A(a[25]), .B(b[25]), .Z(n103) );
  NAND U132 ( .A(n101), .B(n100), .Z(n102) );
  NAND U133 ( .A(n103), .B(n102), .Z(n104) );
  XOR U134 ( .A(n105), .B(n104), .Z(c[26]) );
  XOR U135 ( .A(a[27]), .B(b[27]), .Z(n109) );
  NAND U136 ( .A(a[26]), .B(b[26]), .Z(n107) );
  NAND U137 ( .A(n105), .B(n104), .Z(n106) );
  NAND U138 ( .A(n107), .B(n106), .Z(n108) );
  XOR U139 ( .A(n109), .B(n108), .Z(c[27]) );
  XOR U140 ( .A(a[28]), .B(b[28]), .Z(n113) );
  NAND U141 ( .A(a[27]), .B(b[27]), .Z(n111) );
  NAND U142 ( .A(n109), .B(n108), .Z(n110) );
  NAND U143 ( .A(n111), .B(n110), .Z(n112) );
  XOR U144 ( .A(n113), .B(n112), .Z(c[28]) );
  XOR U145 ( .A(a[29]), .B(b[29]), .Z(n117) );
  NAND U146 ( .A(a[28]), .B(b[28]), .Z(n115) );
  NAND U147 ( .A(n113), .B(n112), .Z(n114) );
  NAND U148 ( .A(n115), .B(n114), .Z(n116) );
  XOR U149 ( .A(n117), .B(n116), .Z(c[29]) );
  XOR U150 ( .A(a[30]), .B(b[30]), .Z(n121) );
  NAND U151 ( .A(a[29]), .B(b[29]), .Z(n119) );
  NAND U152 ( .A(n117), .B(n116), .Z(n118) );
  NAND U153 ( .A(n119), .B(n118), .Z(n120) );
  XOR U154 ( .A(n121), .B(n120), .Z(c[30]) );
  XOR U155 ( .A(a[31]), .B(b[31]), .Z(n125) );
  NAND U156 ( .A(a[30]), .B(b[30]), .Z(n123) );
  NAND U157 ( .A(n121), .B(n120), .Z(n122) );
  NAND U158 ( .A(n123), .B(n122), .Z(n124) );
  XOR U159 ( .A(n125), .B(n124), .Z(c[31]) );
  XOR U160 ( .A(a[32]), .B(b[32]), .Z(n129) );
  NAND U161 ( .A(a[31]), .B(b[31]), .Z(n127) );
  NAND U162 ( .A(n125), .B(n124), .Z(n126) );
  NAND U163 ( .A(n127), .B(n126), .Z(n128) );
  XOR U164 ( .A(n129), .B(n128), .Z(c[32]) );
  XOR U165 ( .A(a[33]), .B(b[33]), .Z(n133) );
  NAND U166 ( .A(a[32]), .B(b[32]), .Z(n131) );
  NAND U167 ( .A(n129), .B(n128), .Z(n130) );
  NAND U168 ( .A(n131), .B(n130), .Z(n132) );
  XOR U169 ( .A(n133), .B(n132), .Z(c[33]) );
  XOR U170 ( .A(a[34]), .B(b[34]), .Z(n137) );
  NAND U171 ( .A(a[33]), .B(b[33]), .Z(n135) );
  NAND U172 ( .A(n133), .B(n132), .Z(n134) );
  NAND U173 ( .A(n135), .B(n134), .Z(n136) );
  XOR U174 ( .A(n137), .B(n136), .Z(c[34]) );
  XOR U175 ( .A(a[35]), .B(b[35]), .Z(n141) );
  NAND U176 ( .A(a[34]), .B(b[34]), .Z(n139) );
  NAND U177 ( .A(n137), .B(n136), .Z(n138) );
  NAND U178 ( .A(n139), .B(n138), .Z(n140) );
  XOR U179 ( .A(n141), .B(n140), .Z(c[35]) );
  XOR U180 ( .A(a[36]), .B(b[36]), .Z(n145) );
  NAND U181 ( .A(a[35]), .B(b[35]), .Z(n143) );
  NAND U182 ( .A(n141), .B(n140), .Z(n142) );
  NAND U183 ( .A(n143), .B(n142), .Z(n144) );
  XOR U184 ( .A(n145), .B(n144), .Z(c[36]) );
  XOR U185 ( .A(a[37]), .B(b[37]), .Z(n149) );
  NAND U186 ( .A(a[36]), .B(b[36]), .Z(n147) );
  NAND U187 ( .A(n145), .B(n144), .Z(n146) );
  NAND U188 ( .A(n147), .B(n146), .Z(n148) );
  XOR U189 ( .A(n149), .B(n148), .Z(c[37]) );
  XOR U190 ( .A(a[38]), .B(b[38]), .Z(n153) );
  NAND U191 ( .A(a[37]), .B(b[37]), .Z(n151) );
  NAND U192 ( .A(n149), .B(n148), .Z(n150) );
  NAND U193 ( .A(n151), .B(n150), .Z(n152) );
  XOR U194 ( .A(n153), .B(n152), .Z(c[38]) );
  XOR U195 ( .A(a[39]), .B(b[39]), .Z(n157) );
  NAND U196 ( .A(a[38]), .B(b[38]), .Z(n155) );
  NAND U197 ( .A(n153), .B(n152), .Z(n154) );
  NAND U198 ( .A(n155), .B(n154), .Z(n156) );
  XOR U199 ( .A(n157), .B(n156), .Z(c[39]) );
  XOR U200 ( .A(a[40]), .B(b[40]), .Z(n161) );
  NAND U201 ( .A(a[39]), .B(b[39]), .Z(n159) );
  NAND U202 ( .A(n157), .B(n156), .Z(n158) );
  NAND U203 ( .A(n159), .B(n158), .Z(n160) );
  XOR U204 ( .A(n161), .B(n160), .Z(c[40]) );
  XOR U205 ( .A(a[41]), .B(b[41]), .Z(n165) );
  NAND U206 ( .A(a[40]), .B(b[40]), .Z(n163) );
  NAND U207 ( .A(n161), .B(n160), .Z(n162) );
  NAND U208 ( .A(n163), .B(n162), .Z(n164) );
  XOR U209 ( .A(n165), .B(n164), .Z(c[41]) );
  XOR U210 ( .A(a[42]), .B(b[42]), .Z(n169) );
  NAND U211 ( .A(a[41]), .B(b[41]), .Z(n167) );
  NAND U212 ( .A(n165), .B(n164), .Z(n166) );
  NAND U213 ( .A(n167), .B(n166), .Z(n168) );
  XOR U214 ( .A(n169), .B(n168), .Z(c[42]) );
  XOR U215 ( .A(a[43]), .B(b[43]), .Z(n173) );
  NAND U216 ( .A(a[42]), .B(b[42]), .Z(n171) );
  NAND U217 ( .A(n169), .B(n168), .Z(n170) );
  NAND U218 ( .A(n171), .B(n170), .Z(n172) );
  XOR U219 ( .A(n173), .B(n172), .Z(c[43]) );
  XOR U220 ( .A(a[44]), .B(b[44]), .Z(n177) );
  NAND U221 ( .A(a[43]), .B(b[43]), .Z(n175) );
  NAND U222 ( .A(n173), .B(n172), .Z(n174) );
  NAND U223 ( .A(n175), .B(n174), .Z(n176) );
  XOR U224 ( .A(n177), .B(n176), .Z(c[44]) );
  XOR U225 ( .A(a[45]), .B(b[45]), .Z(n181) );
  NAND U226 ( .A(a[44]), .B(b[44]), .Z(n179) );
  NAND U227 ( .A(n177), .B(n176), .Z(n178) );
  NAND U228 ( .A(n179), .B(n178), .Z(n180) );
  XOR U229 ( .A(n181), .B(n180), .Z(c[45]) );
  XOR U230 ( .A(a[46]), .B(b[46]), .Z(n185) );
  NAND U231 ( .A(a[45]), .B(b[45]), .Z(n183) );
  NAND U232 ( .A(n181), .B(n180), .Z(n182) );
  NAND U233 ( .A(n183), .B(n182), .Z(n184) );
  XOR U234 ( .A(n185), .B(n184), .Z(c[46]) );
  XOR U235 ( .A(a[47]), .B(b[47]), .Z(n189) );
  NAND U236 ( .A(a[46]), .B(b[46]), .Z(n187) );
  NAND U237 ( .A(n185), .B(n184), .Z(n186) );
  NAND U238 ( .A(n187), .B(n186), .Z(n188) );
  XOR U239 ( .A(n189), .B(n188), .Z(c[47]) );
  XOR U240 ( .A(a[48]), .B(b[48]), .Z(n193) );
  NAND U241 ( .A(a[47]), .B(b[47]), .Z(n191) );
  NAND U242 ( .A(n189), .B(n188), .Z(n190) );
  NAND U243 ( .A(n191), .B(n190), .Z(n192) );
  XOR U244 ( .A(n193), .B(n192), .Z(c[48]) );
  XOR U245 ( .A(a[49]), .B(b[49]), .Z(n197) );
  NAND U246 ( .A(a[48]), .B(b[48]), .Z(n195) );
  NAND U247 ( .A(n193), .B(n192), .Z(n194) );
  NAND U248 ( .A(n195), .B(n194), .Z(n196) );
  XOR U249 ( .A(n197), .B(n196), .Z(c[49]) );
  XOR U250 ( .A(a[50]), .B(b[50]), .Z(n201) );
  NAND U251 ( .A(a[49]), .B(b[49]), .Z(n199) );
  NAND U252 ( .A(n197), .B(n196), .Z(n198) );
  NAND U253 ( .A(n199), .B(n198), .Z(n200) );
  XOR U254 ( .A(n201), .B(n200), .Z(c[50]) );
  XOR U255 ( .A(a[51]), .B(b[51]), .Z(n205) );
  NAND U256 ( .A(a[50]), .B(b[50]), .Z(n203) );
  NAND U257 ( .A(n201), .B(n200), .Z(n202) );
  NAND U258 ( .A(n203), .B(n202), .Z(n204) );
  XOR U259 ( .A(n205), .B(n204), .Z(c[51]) );
  XOR U260 ( .A(a[52]), .B(b[52]), .Z(n209) );
  NAND U261 ( .A(a[51]), .B(b[51]), .Z(n207) );
  NAND U262 ( .A(n205), .B(n204), .Z(n206) );
  NAND U263 ( .A(n207), .B(n206), .Z(n208) );
  XOR U264 ( .A(n209), .B(n208), .Z(c[52]) );
  XOR U265 ( .A(a[53]), .B(b[53]), .Z(n213) );
  NAND U266 ( .A(a[52]), .B(b[52]), .Z(n211) );
  NAND U267 ( .A(n209), .B(n208), .Z(n210) );
  NAND U268 ( .A(n211), .B(n210), .Z(n212) );
  XOR U269 ( .A(n213), .B(n212), .Z(c[53]) );
  XOR U270 ( .A(a[54]), .B(b[54]), .Z(n217) );
  NAND U271 ( .A(a[53]), .B(b[53]), .Z(n215) );
  NAND U272 ( .A(n213), .B(n212), .Z(n214) );
  NAND U273 ( .A(n215), .B(n214), .Z(n216) );
  XOR U274 ( .A(n217), .B(n216), .Z(c[54]) );
  XOR U275 ( .A(a[55]), .B(b[55]), .Z(n221) );
  NAND U276 ( .A(a[54]), .B(b[54]), .Z(n219) );
  NAND U277 ( .A(n217), .B(n216), .Z(n218) );
  NAND U278 ( .A(n219), .B(n218), .Z(n220) );
  XOR U279 ( .A(n221), .B(n220), .Z(c[55]) );
  XOR U280 ( .A(a[56]), .B(b[56]), .Z(n225) );
  NAND U281 ( .A(a[55]), .B(b[55]), .Z(n223) );
  NAND U282 ( .A(n221), .B(n220), .Z(n222) );
  NAND U283 ( .A(n223), .B(n222), .Z(n224) );
  XOR U284 ( .A(n225), .B(n224), .Z(c[56]) );
  XOR U285 ( .A(a[57]), .B(b[57]), .Z(n229) );
  NAND U286 ( .A(a[56]), .B(b[56]), .Z(n227) );
  NAND U287 ( .A(n225), .B(n224), .Z(n226) );
  NAND U288 ( .A(n227), .B(n226), .Z(n228) );
  XOR U289 ( .A(n229), .B(n228), .Z(c[57]) );
  XOR U290 ( .A(a[58]), .B(b[58]), .Z(n233) );
  NAND U291 ( .A(a[57]), .B(b[57]), .Z(n231) );
  NAND U292 ( .A(n229), .B(n228), .Z(n230) );
  NAND U293 ( .A(n231), .B(n230), .Z(n232) );
  XOR U294 ( .A(n233), .B(n232), .Z(c[58]) );
  XOR U295 ( .A(a[59]), .B(b[59]), .Z(n237) );
  NAND U296 ( .A(a[58]), .B(b[58]), .Z(n235) );
  NAND U297 ( .A(n233), .B(n232), .Z(n234) );
  NAND U298 ( .A(n235), .B(n234), .Z(n236) );
  XOR U299 ( .A(n237), .B(n236), .Z(c[59]) );
  XOR U300 ( .A(a[60]), .B(b[60]), .Z(n241) );
  NAND U301 ( .A(a[59]), .B(b[59]), .Z(n239) );
  NAND U302 ( .A(n237), .B(n236), .Z(n238) );
  NAND U303 ( .A(n239), .B(n238), .Z(n240) );
  XOR U304 ( .A(n241), .B(n240), .Z(c[60]) );
  XOR U305 ( .A(a[61]), .B(b[61]), .Z(n245) );
  NAND U306 ( .A(a[60]), .B(b[60]), .Z(n243) );
  NAND U307 ( .A(n241), .B(n240), .Z(n242) );
  NAND U308 ( .A(n243), .B(n242), .Z(n244) );
  XOR U309 ( .A(n245), .B(n244), .Z(c[61]) );
  XOR U310 ( .A(a[62]), .B(b[62]), .Z(n249) );
  NAND U311 ( .A(a[61]), .B(b[61]), .Z(n247) );
  NAND U312 ( .A(n245), .B(n244), .Z(n246) );
  NAND U313 ( .A(n247), .B(n246), .Z(n248) );
  XOR U314 ( .A(n249), .B(n248), .Z(c[62]) );
  XOR U315 ( .A(a[63]), .B(b[63]), .Z(n253) );
  NAND U316 ( .A(a[62]), .B(b[62]), .Z(n251) );
  NAND U317 ( .A(n249), .B(n248), .Z(n250) );
  NAND U318 ( .A(n251), .B(n250), .Z(n252) );
  XOR U319 ( .A(n253), .B(n252), .Z(c[63]) );
  XOR U320 ( .A(a[64]), .B(b[64]), .Z(n257) );
  NAND U321 ( .A(a[63]), .B(b[63]), .Z(n255) );
  NAND U322 ( .A(n253), .B(n252), .Z(n254) );
  NAND U323 ( .A(n255), .B(n254), .Z(n256) );
  XOR U324 ( .A(n257), .B(n256), .Z(c[64]) );
  XOR U325 ( .A(a[65]), .B(b[65]), .Z(n261) );
  NAND U326 ( .A(a[64]), .B(b[64]), .Z(n259) );
  NAND U327 ( .A(n257), .B(n256), .Z(n258) );
  NAND U328 ( .A(n259), .B(n258), .Z(n260) );
  XOR U329 ( .A(n261), .B(n260), .Z(c[65]) );
  XOR U330 ( .A(a[66]), .B(b[66]), .Z(n265) );
  NAND U331 ( .A(a[65]), .B(b[65]), .Z(n263) );
  NAND U332 ( .A(n261), .B(n260), .Z(n262) );
  NAND U333 ( .A(n263), .B(n262), .Z(n264) );
  XOR U334 ( .A(n265), .B(n264), .Z(c[66]) );
  XOR U335 ( .A(a[67]), .B(b[67]), .Z(n269) );
  NAND U336 ( .A(a[66]), .B(b[66]), .Z(n267) );
  NAND U337 ( .A(n265), .B(n264), .Z(n266) );
  NAND U338 ( .A(n267), .B(n266), .Z(n268) );
  XOR U339 ( .A(n269), .B(n268), .Z(c[67]) );
  XOR U340 ( .A(a[68]), .B(b[68]), .Z(n273) );
  NAND U341 ( .A(a[67]), .B(b[67]), .Z(n271) );
  NAND U342 ( .A(n269), .B(n268), .Z(n270) );
  NAND U343 ( .A(n271), .B(n270), .Z(n272) );
  XOR U344 ( .A(n273), .B(n272), .Z(c[68]) );
  XOR U345 ( .A(a[69]), .B(b[69]), .Z(n277) );
  NAND U346 ( .A(a[68]), .B(b[68]), .Z(n275) );
  NAND U347 ( .A(n273), .B(n272), .Z(n274) );
  NAND U348 ( .A(n275), .B(n274), .Z(n276) );
  XOR U349 ( .A(n277), .B(n276), .Z(c[69]) );
  XOR U350 ( .A(a[70]), .B(b[70]), .Z(n281) );
  NAND U351 ( .A(a[69]), .B(b[69]), .Z(n279) );
  NAND U352 ( .A(n277), .B(n276), .Z(n278) );
  NAND U353 ( .A(n279), .B(n278), .Z(n280) );
  XOR U354 ( .A(n281), .B(n280), .Z(c[70]) );
  XOR U355 ( .A(a[71]), .B(b[71]), .Z(n285) );
  NAND U356 ( .A(a[70]), .B(b[70]), .Z(n283) );
  NAND U357 ( .A(n281), .B(n280), .Z(n282) );
  NAND U358 ( .A(n283), .B(n282), .Z(n284) );
  XOR U359 ( .A(n285), .B(n284), .Z(c[71]) );
  XOR U360 ( .A(a[72]), .B(b[72]), .Z(n289) );
  NAND U361 ( .A(a[71]), .B(b[71]), .Z(n287) );
  NAND U362 ( .A(n285), .B(n284), .Z(n286) );
  NAND U363 ( .A(n287), .B(n286), .Z(n288) );
  XOR U364 ( .A(n289), .B(n288), .Z(c[72]) );
  XOR U365 ( .A(a[73]), .B(b[73]), .Z(n293) );
  NAND U366 ( .A(a[72]), .B(b[72]), .Z(n291) );
  NAND U367 ( .A(n289), .B(n288), .Z(n290) );
  NAND U368 ( .A(n291), .B(n290), .Z(n292) );
  XOR U369 ( .A(n293), .B(n292), .Z(c[73]) );
  XOR U370 ( .A(a[74]), .B(b[74]), .Z(n297) );
  NAND U371 ( .A(a[73]), .B(b[73]), .Z(n295) );
  NAND U372 ( .A(n293), .B(n292), .Z(n294) );
  NAND U373 ( .A(n295), .B(n294), .Z(n296) );
  XOR U374 ( .A(n297), .B(n296), .Z(c[74]) );
  XOR U375 ( .A(a[75]), .B(b[75]), .Z(n301) );
  NAND U376 ( .A(a[74]), .B(b[74]), .Z(n299) );
  NAND U377 ( .A(n297), .B(n296), .Z(n298) );
  NAND U378 ( .A(n299), .B(n298), .Z(n300) );
  XOR U379 ( .A(n301), .B(n300), .Z(c[75]) );
  XOR U380 ( .A(a[76]), .B(b[76]), .Z(n305) );
  NAND U381 ( .A(a[75]), .B(b[75]), .Z(n303) );
  NAND U382 ( .A(n301), .B(n300), .Z(n302) );
  NAND U383 ( .A(n303), .B(n302), .Z(n304) );
  XOR U384 ( .A(n305), .B(n304), .Z(c[76]) );
  XOR U385 ( .A(a[77]), .B(b[77]), .Z(n309) );
  NAND U386 ( .A(a[76]), .B(b[76]), .Z(n307) );
  NAND U387 ( .A(n305), .B(n304), .Z(n306) );
  NAND U388 ( .A(n307), .B(n306), .Z(n308) );
  XOR U389 ( .A(n309), .B(n308), .Z(c[77]) );
  XOR U390 ( .A(a[78]), .B(b[78]), .Z(n313) );
  NAND U391 ( .A(a[77]), .B(b[77]), .Z(n311) );
  NAND U392 ( .A(n309), .B(n308), .Z(n310) );
  NAND U393 ( .A(n311), .B(n310), .Z(n312) );
  XOR U394 ( .A(n313), .B(n312), .Z(c[78]) );
  XOR U395 ( .A(a[79]), .B(b[79]), .Z(n317) );
  NAND U396 ( .A(a[78]), .B(b[78]), .Z(n315) );
  NAND U397 ( .A(n313), .B(n312), .Z(n314) );
  NAND U398 ( .A(n315), .B(n314), .Z(n316) );
  XOR U399 ( .A(n317), .B(n316), .Z(c[79]) );
  XOR U400 ( .A(a[80]), .B(b[80]), .Z(n321) );
  NAND U401 ( .A(a[79]), .B(b[79]), .Z(n319) );
  NAND U402 ( .A(n317), .B(n316), .Z(n318) );
  NAND U403 ( .A(n319), .B(n318), .Z(n320) );
  XOR U404 ( .A(n321), .B(n320), .Z(c[80]) );
  XOR U405 ( .A(a[81]), .B(b[81]), .Z(n325) );
  NAND U406 ( .A(a[80]), .B(b[80]), .Z(n323) );
  NAND U407 ( .A(n321), .B(n320), .Z(n322) );
  NAND U408 ( .A(n323), .B(n322), .Z(n324) );
  XOR U409 ( .A(n325), .B(n324), .Z(c[81]) );
  XOR U410 ( .A(a[82]), .B(b[82]), .Z(n329) );
  NAND U411 ( .A(a[81]), .B(b[81]), .Z(n327) );
  NAND U412 ( .A(n325), .B(n324), .Z(n326) );
  NAND U413 ( .A(n327), .B(n326), .Z(n328) );
  XOR U414 ( .A(n329), .B(n328), .Z(c[82]) );
  XOR U415 ( .A(a[83]), .B(b[83]), .Z(n333) );
  NAND U416 ( .A(a[82]), .B(b[82]), .Z(n331) );
  NAND U417 ( .A(n329), .B(n328), .Z(n330) );
  NAND U418 ( .A(n331), .B(n330), .Z(n332) );
  XOR U419 ( .A(n333), .B(n332), .Z(c[83]) );
  XOR U420 ( .A(a[84]), .B(b[84]), .Z(n337) );
  NAND U421 ( .A(a[83]), .B(b[83]), .Z(n335) );
  NAND U422 ( .A(n333), .B(n332), .Z(n334) );
  NAND U423 ( .A(n335), .B(n334), .Z(n336) );
  XOR U424 ( .A(n337), .B(n336), .Z(c[84]) );
  XOR U425 ( .A(a[85]), .B(b[85]), .Z(n341) );
  NAND U426 ( .A(a[84]), .B(b[84]), .Z(n339) );
  NAND U427 ( .A(n337), .B(n336), .Z(n338) );
  NAND U428 ( .A(n339), .B(n338), .Z(n340) );
  XOR U429 ( .A(n341), .B(n340), .Z(c[85]) );
  XOR U430 ( .A(a[86]), .B(b[86]), .Z(n345) );
  NAND U431 ( .A(a[85]), .B(b[85]), .Z(n343) );
  NAND U432 ( .A(n341), .B(n340), .Z(n342) );
  NAND U433 ( .A(n343), .B(n342), .Z(n344) );
  XOR U434 ( .A(n345), .B(n344), .Z(c[86]) );
  XOR U435 ( .A(a[87]), .B(b[87]), .Z(n349) );
  NAND U436 ( .A(a[86]), .B(b[86]), .Z(n347) );
  NAND U437 ( .A(n345), .B(n344), .Z(n346) );
  NAND U438 ( .A(n347), .B(n346), .Z(n348) );
  XOR U439 ( .A(n349), .B(n348), .Z(c[87]) );
  XOR U440 ( .A(a[88]), .B(b[88]), .Z(n353) );
  NAND U441 ( .A(a[87]), .B(b[87]), .Z(n351) );
  NAND U442 ( .A(n349), .B(n348), .Z(n350) );
  NAND U443 ( .A(n351), .B(n350), .Z(n352) );
  XOR U444 ( .A(n353), .B(n352), .Z(c[88]) );
  XOR U445 ( .A(a[89]), .B(b[89]), .Z(n357) );
  NAND U446 ( .A(a[88]), .B(b[88]), .Z(n355) );
  NAND U447 ( .A(n353), .B(n352), .Z(n354) );
  NAND U448 ( .A(n355), .B(n354), .Z(n356) );
  XOR U449 ( .A(n357), .B(n356), .Z(c[89]) );
  XOR U450 ( .A(a[90]), .B(b[90]), .Z(n361) );
  NAND U451 ( .A(a[89]), .B(b[89]), .Z(n359) );
  NAND U452 ( .A(n357), .B(n356), .Z(n358) );
  NAND U453 ( .A(n359), .B(n358), .Z(n360) );
  XOR U454 ( .A(n361), .B(n360), .Z(c[90]) );
  XOR U455 ( .A(a[91]), .B(b[91]), .Z(n365) );
  NAND U456 ( .A(a[90]), .B(b[90]), .Z(n363) );
  NAND U457 ( .A(n361), .B(n360), .Z(n362) );
  NAND U458 ( .A(n363), .B(n362), .Z(n364) );
  XOR U459 ( .A(n365), .B(n364), .Z(c[91]) );
  XOR U460 ( .A(a[92]), .B(b[92]), .Z(n369) );
  NAND U461 ( .A(a[91]), .B(b[91]), .Z(n367) );
  NAND U462 ( .A(n365), .B(n364), .Z(n366) );
  NAND U463 ( .A(n367), .B(n366), .Z(n368) );
  XOR U464 ( .A(n369), .B(n368), .Z(c[92]) );
  XOR U465 ( .A(a[93]), .B(b[93]), .Z(n373) );
  NAND U466 ( .A(a[92]), .B(b[92]), .Z(n371) );
  NAND U467 ( .A(n369), .B(n368), .Z(n370) );
  NAND U468 ( .A(n371), .B(n370), .Z(n372) );
  XOR U469 ( .A(n373), .B(n372), .Z(c[93]) );
  XOR U470 ( .A(a[94]), .B(b[94]), .Z(n377) );
  NAND U471 ( .A(a[93]), .B(b[93]), .Z(n375) );
  NAND U472 ( .A(n373), .B(n372), .Z(n374) );
  NAND U473 ( .A(n375), .B(n374), .Z(n376) );
  XOR U474 ( .A(n377), .B(n376), .Z(c[94]) );
  XOR U475 ( .A(a[95]), .B(b[95]), .Z(n381) );
  NAND U476 ( .A(a[94]), .B(b[94]), .Z(n379) );
  NAND U477 ( .A(n377), .B(n376), .Z(n378) );
  NAND U478 ( .A(n379), .B(n378), .Z(n380) );
  XOR U479 ( .A(n381), .B(n380), .Z(c[95]) );
  XOR U480 ( .A(a[96]), .B(b[96]), .Z(n385) );
  NAND U481 ( .A(a[95]), .B(b[95]), .Z(n383) );
  NAND U482 ( .A(n381), .B(n380), .Z(n382) );
  NAND U483 ( .A(n383), .B(n382), .Z(n384) );
  XOR U484 ( .A(n385), .B(n384), .Z(c[96]) );
  XOR U485 ( .A(a[97]), .B(b[97]), .Z(n389) );
  NAND U486 ( .A(a[96]), .B(b[96]), .Z(n387) );
  NAND U487 ( .A(n385), .B(n384), .Z(n386) );
  NAND U488 ( .A(n387), .B(n386), .Z(n388) );
  XOR U489 ( .A(n389), .B(n388), .Z(c[97]) );
  XOR U490 ( .A(a[98]), .B(b[98]), .Z(n393) );
  NAND U491 ( .A(a[97]), .B(b[97]), .Z(n391) );
  NAND U492 ( .A(n389), .B(n388), .Z(n390) );
  NAND U493 ( .A(n391), .B(n390), .Z(n392) );
  XOR U494 ( .A(n393), .B(n392), .Z(c[98]) );
  XOR U495 ( .A(a[99]), .B(b[99]), .Z(n397) );
  NAND U496 ( .A(a[98]), .B(b[98]), .Z(n395) );
  NAND U497 ( .A(n393), .B(n392), .Z(n394) );
  NAND U498 ( .A(n395), .B(n394), .Z(n396) );
  XOR U499 ( .A(n397), .B(n396), .Z(c[99]) );
  XOR U500 ( .A(a[100]), .B(b[100]), .Z(n401) );
  NAND U501 ( .A(a[99]), .B(b[99]), .Z(n399) );
  NAND U502 ( .A(n397), .B(n396), .Z(n398) );
  NAND U503 ( .A(n399), .B(n398), .Z(n400) );
  XOR U504 ( .A(n401), .B(n400), .Z(c[100]) );
  XOR U505 ( .A(a[101]), .B(b[101]), .Z(n405) );
  NAND U506 ( .A(a[100]), .B(b[100]), .Z(n403) );
  NAND U507 ( .A(n401), .B(n400), .Z(n402) );
  NAND U508 ( .A(n403), .B(n402), .Z(n404) );
  XOR U509 ( .A(n405), .B(n404), .Z(c[101]) );
  XOR U510 ( .A(a[102]), .B(b[102]), .Z(n409) );
  NAND U511 ( .A(a[101]), .B(b[101]), .Z(n407) );
  NAND U512 ( .A(n405), .B(n404), .Z(n406) );
  NAND U513 ( .A(n407), .B(n406), .Z(n408) );
  XOR U514 ( .A(n409), .B(n408), .Z(c[102]) );
  XOR U515 ( .A(a[103]), .B(b[103]), .Z(n413) );
  NAND U516 ( .A(a[102]), .B(b[102]), .Z(n411) );
  NAND U517 ( .A(n409), .B(n408), .Z(n410) );
  NAND U518 ( .A(n411), .B(n410), .Z(n412) );
  XOR U519 ( .A(n413), .B(n412), .Z(c[103]) );
  XOR U520 ( .A(a[104]), .B(b[104]), .Z(n417) );
  NAND U521 ( .A(a[103]), .B(b[103]), .Z(n415) );
  NAND U522 ( .A(n413), .B(n412), .Z(n414) );
  NAND U523 ( .A(n415), .B(n414), .Z(n416) );
  XOR U524 ( .A(n417), .B(n416), .Z(c[104]) );
  XOR U525 ( .A(a[105]), .B(b[105]), .Z(n421) );
  NAND U526 ( .A(a[104]), .B(b[104]), .Z(n419) );
  NAND U527 ( .A(n417), .B(n416), .Z(n418) );
  NAND U528 ( .A(n419), .B(n418), .Z(n420) );
  XOR U529 ( .A(n421), .B(n420), .Z(c[105]) );
  XOR U530 ( .A(a[106]), .B(b[106]), .Z(n425) );
  NAND U531 ( .A(a[105]), .B(b[105]), .Z(n423) );
  NAND U532 ( .A(n421), .B(n420), .Z(n422) );
  NAND U533 ( .A(n423), .B(n422), .Z(n424) );
  XOR U534 ( .A(n425), .B(n424), .Z(c[106]) );
  XOR U535 ( .A(a[107]), .B(b[107]), .Z(n429) );
  NAND U536 ( .A(a[106]), .B(b[106]), .Z(n427) );
  NAND U537 ( .A(n425), .B(n424), .Z(n426) );
  NAND U538 ( .A(n427), .B(n426), .Z(n428) );
  XOR U539 ( .A(n429), .B(n428), .Z(c[107]) );
  XOR U540 ( .A(a[108]), .B(b[108]), .Z(n433) );
  NAND U541 ( .A(a[107]), .B(b[107]), .Z(n431) );
  NAND U542 ( .A(n429), .B(n428), .Z(n430) );
  NAND U543 ( .A(n431), .B(n430), .Z(n432) );
  XOR U544 ( .A(n433), .B(n432), .Z(c[108]) );
  XOR U545 ( .A(a[109]), .B(b[109]), .Z(n437) );
  NAND U546 ( .A(a[108]), .B(b[108]), .Z(n435) );
  NAND U547 ( .A(n433), .B(n432), .Z(n434) );
  NAND U548 ( .A(n435), .B(n434), .Z(n436) );
  XOR U549 ( .A(n437), .B(n436), .Z(c[109]) );
  XOR U550 ( .A(a[110]), .B(b[110]), .Z(n441) );
  NAND U551 ( .A(a[109]), .B(b[109]), .Z(n439) );
  NAND U552 ( .A(n437), .B(n436), .Z(n438) );
  NAND U553 ( .A(n439), .B(n438), .Z(n440) );
  XOR U554 ( .A(n441), .B(n440), .Z(c[110]) );
  XOR U555 ( .A(a[111]), .B(b[111]), .Z(n445) );
  NAND U556 ( .A(a[110]), .B(b[110]), .Z(n443) );
  NAND U557 ( .A(n441), .B(n440), .Z(n442) );
  NAND U558 ( .A(n443), .B(n442), .Z(n444) );
  XOR U559 ( .A(n445), .B(n444), .Z(c[111]) );
  XOR U560 ( .A(a[112]), .B(b[112]), .Z(n449) );
  NAND U561 ( .A(a[111]), .B(b[111]), .Z(n447) );
  NAND U562 ( .A(n445), .B(n444), .Z(n446) );
  NAND U563 ( .A(n447), .B(n446), .Z(n448) );
  XOR U564 ( .A(n449), .B(n448), .Z(c[112]) );
  XOR U565 ( .A(a[113]), .B(b[113]), .Z(n453) );
  NAND U566 ( .A(a[112]), .B(b[112]), .Z(n451) );
  NAND U567 ( .A(n449), .B(n448), .Z(n450) );
  NAND U568 ( .A(n451), .B(n450), .Z(n452) );
  XOR U569 ( .A(n453), .B(n452), .Z(c[113]) );
  XOR U570 ( .A(a[114]), .B(b[114]), .Z(n457) );
  NAND U571 ( .A(a[113]), .B(b[113]), .Z(n455) );
  NAND U572 ( .A(n453), .B(n452), .Z(n454) );
  NAND U573 ( .A(n455), .B(n454), .Z(n456) );
  XOR U574 ( .A(n457), .B(n456), .Z(c[114]) );
  XOR U575 ( .A(a[115]), .B(b[115]), .Z(n461) );
  NAND U576 ( .A(a[114]), .B(b[114]), .Z(n459) );
  NAND U577 ( .A(n457), .B(n456), .Z(n458) );
  NAND U578 ( .A(n459), .B(n458), .Z(n460) );
  XOR U579 ( .A(n461), .B(n460), .Z(c[115]) );
  XOR U580 ( .A(a[116]), .B(b[116]), .Z(n465) );
  NAND U581 ( .A(a[115]), .B(b[115]), .Z(n463) );
  NAND U582 ( .A(n461), .B(n460), .Z(n462) );
  NAND U583 ( .A(n463), .B(n462), .Z(n464) );
  XOR U584 ( .A(n465), .B(n464), .Z(c[116]) );
  XOR U585 ( .A(a[117]), .B(b[117]), .Z(n469) );
  NAND U586 ( .A(a[116]), .B(b[116]), .Z(n467) );
  NAND U587 ( .A(n465), .B(n464), .Z(n466) );
  NAND U588 ( .A(n467), .B(n466), .Z(n468) );
  XOR U589 ( .A(n469), .B(n468), .Z(c[117]) );
  XOR U590 ( .A(a[118]), .B(b[118]), .Z(n473) );
  NAND U591 ( .A(a[117]), .B(b[117]), .Z(n471) );
  NAND U592 ( .A(n469), .B(n468), .Z(n470) );
  NAND U593 ( .A(n471), .B(n470), .Z(n472) );
  XOR U594 ( .A(n473), .B(n472), .Z(c[118]) );
  XOR U595 ( .A(a[119]), .B(b[119]), .Z(n477) );
  NAND U596 ( .A(a[118]), .B(b[118]), .Z(n475) );
  NAND U597 ( .A(n473), .B(n472), .Z(n474) );
  NAND U598 ( .A(n475), .B(n474), .Z(n476) );
  XOR U599 ( .A(n477), .B(n476), .Z(c[119]) );
  XOR U600 ( .A(a[120]), .B(b[120]), .Z(n481) );
  NAND U601 ( .A(a[119]), .B(b[119]), .Z(n479) );
  NAND U602 ( .A(n477), .B(n476), .Z(n478) );
  NAND U603 ( .A(n479), .B(n478), .Z(n480) );
  XOR U604 ( .A(n481), .B(n480), .Z(c[120]) );
  XOR U605 ( .A(a[121]), .B(b[121]), .Z(n485) );
  NAND U606 ( .A(a[120]), .B(b[120]), .Z(n483) );
  NAND U607 ( .A(n481), .B(n480), .Z(n482) );
  NAND U608 ( .A(n483), .B(n482), .Z(n484) );
  XOR U609 ( .A(n485), .B(n484), .Z(c[121]) );
  XOR U610 ( .A(a[122]), .B(b[122]), .Z(n489) );
  NAND U611 ( .A(a[121]), .B(b[121]), .Z(n487) );
  NAND U612 ( .A(n485), .B(n484), .Z(n486) );
  NAND U613 ( .A(n487), .B(n486), .Z(n488) );
  XOR U614 ( .A(n489), .B(n488), .Z(c[122]) );
  XOR U615 ( .A(a[123]), .B(b[123]), .Z(n493) );
  NAND U616 ( .A(a[122]), .B(b[122]), .Z(n491) );
  NAND U617 ( .A(n489), .B(n488), .Z(n490) );
  NAND U618 ( .A(n491), .B(n490), .Z(n492) );
  XOR U619 ( .A(n493), .B(n492), .Z(c[123]) );
  XOR U620 ( .A(a[124]), .B(b[124]), .Z(n497) );
  NAND U621 ( .A(a[123]), .B(b[123]), .Z(n495) );
  NAND U622 ( .A(n493), .B(n492), .Z(n494) );
  NAND U623 ( .A(n495), .B(n494), .Z(n496) );
  XOR U624 ( .A(n497), .B(n496), .Z(c[124]) );
  XOR U625 ( .A(a[125]), .B(b[125]), .Z(n501) );
  NAND U626 ( .A(a[124]), .B(b[124]), .Z(n499) );
  NAND U627 ( .A(n497), .B(n496), .Z(n498) );
  NAND U628 ( .A(n499), .B(n498), .Z(n500) );
  XOR U629 ( .A(n501), .B(n500), .Z(c[125]) );
  XOR U630 ( .A(a[126]), .B(b[126]), .Z(n505) );
  NAND U631 ( .A(a[125]), .B(b[125]), .Z(n503) );
  NAND U632 ( .A(n501), .B(n500), .Z(n502) );
  NAND U633 ( .A(n503), .B(n502), .Z(n504) );
  XOR U634 ( .A(n505), .B(n504), .Z(c[126]) );
  XOR U635 ( .A(a[127]), .B(b[127]), .Z(n509) );
  NAND U636 ( .A(a[126]), .B(b[126]), .Z(n507) );
  NAND U637 ( .A(n505), .B(n504), .Z(n506) );
  NAND U638 ( .A(n507), .B(n506), .Z(n508) );
  XOR U639 ( .A(n509), .B(n508), .Z(c[127]) );
  XOR U640 ( .A(a[128]), .B(b[128]), .Z(n513) );
  NAND U641 ( .A(a[127]), .B(b[127]), .Z(n511) );
  NAND U642 ( .A(n509), .B(n508), .Z(n510) );
  NAND U643 ( .A(n511), .B(n510), .Z(n512) );
  XOR U644 ( .A(n513), .B(n512), .Z(c[128]) );
  XOR U645 ( .A(a[129]), .B(b[129]), .Z(n517) );
  NAND U646 ( .A(a[128]), .B(b[128]), .Z(n515) );
  NAND U647 ( .A(n513), .B(n512), .Z(n514) );
  NAND U648 ( .A(n515), .B(n514), .Z(n516) );
  XOR U649 ( .A(n517), .B(n516), .Z(c[129]) );
  XOR U650 ( .A(a[130]), .B(b[130]), .Z(n521) );
  NAND U651 ( .A(a[129]), .B(b[129]), .Z(n519) );
  NAND U652 ( .A(n517), .B(n516), .Z(n518) );
  NAND U653 ( .A(n519), .B(n518), .Z(n520) );
  XOR U654 ( .A(n521), .B(n520), .Z(c[130]) );
  XOR U655 ( .A(a[131]), .B(b[131]), .Z(n525) );
  NAND U656 ( .A(a[130]), .B(b[130]), .Z(n523) );
  NAND U657 ( .A(n521), .B(n520), .Z(n522) );
  NAND U658 ( .A(n523), .B(n522), .Z(n524) );
  XOR U659 ( .A(n525), .B(n524), .Z(c[131]) );
  XOR U660 ( .A(a[132]), .B(b[132]), .Z(n529) );
  NAND U661 ( .A(a[131]), .B(b[131]), .Z(n527) );
  NAND U662 ( .A(n525), .B(n524), .Z(n526) );
  NAND U663 ( .A(n527), .B(n526), .Z(n528) );
  XOR U664 ( .A(n529), .B(n528), .Z(c[132]) );
  XOR U665 ( .A(a[133]), .B(b[133]), .Z(n533) );
  NAND U666 ( .A(a[132]), .B(b[132]), .Z(n531) );
  NAND U667 ( .A(n529), .B(n528), .Z(n530) );
  NAND U668 ( .A(n531), .B(n530), .Z(n532) );
  XOR U669 ( .A(n533), .B(n532), .Z(c[133]) );
  XOR U670 ( .A(a[134]), .B(b[134]), .Z(n537) );
  NAND U671 ( .A(a[133]), .B(b[133]), .Z(n535) );
  NAND U672 ( .A(n533), .B(n532), .Z(n534) );
  NAND U673 ( .A(n535), .B(n534), .Z(n536) );
  XOR U674 ( .A(n537), .B(n536), .Z(c[134]) );
  XOR U675 ( .A(a[135]), .B(b[135]), .Z(n541) );
  NAND U676 ( .A(a[134]), .B(b[134]), .Z(n539) );
  NAND U677 ( .A(n537), .B(n536), .Z(n538) );
  NAND U678 ( .A(n539), .B(n538), .Z(n540) );
  XOR U679 ( .A(n541), .B(n540), .Z(c[135]) );
  XOR U680 ( .A(a[136]), .B(b[136]), .Z(n545) );
  NAND U681 ( .A(a[135]), .B(b[135]), .Z(n543) );
  NAND U682 ( .A(n541), .B(n540), .Z(n542) );
  NAND U683 ( .A(n543), .B(n542), .Z(n544) );
  XOR U684 ( .A(n545), .B(n544), .Z(c[136]) );
  XOR U685 ( .A(a[137]), .B(b[137]), .Z(n549) );
  NAND U686 ( .A(a[136]), .B(b[136]), .Z(n547) );
  NAND U687 ( .A(n545), .B(n544), .Z(n546) );
  NAND U688 ( .A(n547), .B(n546), .Z(n548) );
  XOR U689 ( .A(n549), .B(n548), .Z(c[137]) );
  XOR U690 ( .A(a[138]), .B(b[138]), .Z(n553) );
  NAND U691 ( .A(a[137]), .B(b[137]), .Z(n551) );
  NAND U692 ( .A(n549), .B(n548), .Z(n550) );
  NAND U693 ( .A(n551), .B(n550), .Z(n552) );
  XOR U694 ( .A(n553), .B(n552), .Z(c[138]) );
  XOR U695 ( .A(a[139]), .B(b[139]), .Z(n557) );
  NAND U696 ( .A(a[138]), .B(b[138]), .Z(n555) );
  NAND U697 ( .A(n553), .B(n552), .Z(n554) );
  NAND U698 ( .A(n555), .B(n554), .Z(n556) );
  XOR U699 ( .A(n557), .B(n556), .Z(c[139]) );
  XOR U700 ( .A(a[140]), .B(b[140]), .Z(n561) );
  NAND U701 ( .A(a[139]), .B(b[139]), .Z(n559) );
  NAND U702 ( .A(n557), .B(n556), .Z(n558) );
  NAND U703 ( .A(n559), .B(n558), .Z(n560) );
  XOR U704 ( .A(n561), .B(n560), .Z(c[140]) );
  XOR U705 ( .A(a[141]), .B(b[141]), .Z(n565) );
  NAND U706 ( .A(a[140]), .B(b[140]), .Z(n563) );
  NAND U707 ( .A(n561), .B(n560), .Z(n562) );
  NAND U708 ( .A(n563), .B(n562), .Z(n564) );
  XOR U709 ( .A(n565), .B(n564), .Z(c[141]) );
  XOR U710 ( .A(a[142]), .B(b[142]), .Z(n569) );
  NAND U711 ( .A(a[141]), .B(b[141]), .Z(n567) );
  NAND U712 ( .A(n565), .B(n564), .Z(n566) );
  NAND U713 ( .A(n567), .B(n566), .Z(n568) );
  XOR U714 ( .A(n569), .B(n568), .Z(c[142]) );
  XOR U715 ( .A(a[143]), .B(b[143]), .Z(n573) );
  NAND U716 ( .A(a[142]), .B(b[142]), .Z(n571) );
  NAND U717 ( .A(n569), .B(n568), .Z(n570) );
  NAND U718 ( .A(n571), .B(n570), .Z(n572) );
  XOR U719 ( .A(n573), .B(n572), .Z(c[143]) );
  XOR U720 ( .A(a[144]), .B(b[144]), .Z(n577) );
  NAND U721 ( .A(a[143]), .B(b[143]), .Z(n575) );
  NAND U722 ( .A(n573), .B(n572), .Z(n574) );
  NAND U723 ( .A(n575), .B(n574), .Z(n576) );
  XOR U724 ( .A(n577), .B(n576), .Z(c[144]) );
  XOR U725 ( .A(a[145]), .B(b[145]), .Z(n581) );
  NAND U726 ( .A(a[144]), .B(b[144]), .Z(n579) );
  NAND U727 ( .A(n577), .B(n576), .Z(n578) );
  NAND U728 ( .A(n579), .B(n578), .Z(n580) );
  XOR U729 ( .A(n581), .B(n580), .Z(c[145]) );
  XOR U730 ( .A(a[146]), .B(b[146]), .Z(n585) );
  NAND U731 ( .A(a[145]), .B(b[145]), .Z(n583) );
  NAND U732 ( .A(n581), .B(n580), .Z(n582) );
  NAND U733 ( .A(n583), .B(n582), .Z(n584) );
  XOR U734 ( .A(n585), .B(n584), .Z(c[146]) );
  XOR U735 ( .A(a[147]), .B(b[147]), .Z(n589) );
  NAND U736 ( .A(a[146]), .B(b[146]), .Z(n587) );
  NAND U737 ( .A(n585), .B(n584), .Z(n586) );
  NAND U738 ( .A(n587), .B(n586), .Z(n588) );
  XOR U739 ( .A(n589), .B(n588), .Z(c[147]) );
  XOR U740 ( .A(a[148]), .B(b[148]), .Z(n593) );
  NAND U741 ( .A(a[147]), .B(b[147]), .Z(n591) );
  NAND U742 ( .A(n589), .B(n588), .Z(n590) );
  NAND U743 ( .A(n591), .B(n590), .Z(n592) );
  XOR U744 ( .A(n593), .B(n592), .Z(c[148]) );
  XOR U745 ( .A(a[149]), .B(b[149]), .Z(n597) );
  NAND U746 ( .A(a[148]), .B(b[148]), .Z(n595) );
  NAND U747 ( .A(n593), .B(n592), .Z(n594) );
  NAND U748 ( .A(n595), .B(n594), .Z(n596) );
  XOR U749 ( .A(n597), .B(n596), .Z(c[149]) );
  XOR U750 ( .A(a[150]), .B(b[150]), .Z(n601) );
  NAND U751 ( .A(a[149]), .B(b[149]), .Z(n599) );
  NAND U752 ( .A(n597), .B(n596), .Z(n598) );
  NAND U753 ( .A(n599), .B(n598), .Z(n600) );
  XOR U754 ( .A(n601), .B(n600), .Z(c[150]) );
  XOR U755 ( .A(a[151]), .B(b[151]), .Z(n605) );
  NAND U756 ( .A(a[150]), .B(b[150]), .Z(n603) );
  NAND U757 ( .A(n601), .B(n600), .Z(n602) );
  NAND U758 ( .A(n603), .B(n602), .Z(n604) );
  XOR U759 ( .A(n605), .B(n604), .Z(c[151]) );
  XOR U760 ( .A(a[152]), .B(b[152]), .Z(n609) );
  NAND U761 ( .A(a[151]), .B(b[151]), .Z(n607) );
  NAND U762 ( .A(n605), .B(n604), .Z(n606) );
  NAND U763 ( .A(n607), .B(n606), .Z(n608) );
  XOR U764 ( .A(n609), .B(n608), .Z(c[152]) );
  XOR U765 ( .A(a[153]), .B(b[153]), .Z(n613) );
  NAND U766 ( .A(a[152]), .B(b[152]), .Z(n611) );
  NAND U767 ( .A(n609), .B(n608), .Z(n610) );
  NAND U768 ( .A(n611), .B(n610), .Z(n612) );
  XOR U769 ( .A(n613), .B(n612), .Z(c[153]) );
  XOR U770 ( .A(a[154]), .B(b[154]), .Z(n617) );
  NAND U771 ( .A(a[153]), .B(b[153]), .Z(n615) );
  NAND U772 ( .A(n613), .B(n612), .Z(n614) );
  NAND U773 ( .A(n615), .B(n614), .Z(n616) );
  XOR U774 ( .A(n617), .B(n616), .Z(c[154]) );
  XOR U775 ( .A(a[155]), .B(b[155]), .Z(n621) );
  NAND U776 ( .A(a[154]), .B(b[154]), .Z(n619) );
  NAND U777 ( .A(n617), .B(n616), .Z(n618) );
  NAND U778 ( .A(n619), .B(n618), .Z(n620) );
  XOR U779 ( .A(n621), .B(n620), .Z(c[155]) );
  XOR U780 ( .A(a[156]), .B(b[156]), .Z(n625) );
  NAND U781 ( .A(a[155]), .B(b[155]), .Z(n623) );
  NAND U782 ( .A(n621), .B(n620), .Z(n622) );
  NAND U783 ( .A(n623), .B(n622), .Z(n624) );
  XOR U784 ( .A(n625), .B(n624), .Z(c[156]) );
  XOR U785 ( .A(a[157]), .B(b[157]), .Z(n629) );
  NAND U786 ( .A(a[156]), .B(b[156]), .Z(n627) );
  NAND U787 ( .A(n625), .B(n624), .Z(n626) );
  NAND U788 ( .A(n627), .B(n626), .Z(n628) );
  XOR U789 ( .A(n629), .B(n628), .Z(c[157]) );
  XOR U790 ( .A(a[158]), .B(b[158]), .Z(n633) );
  NAND U791 ( .A(a[157]), .B(b[157]), .Z(n631) );
  NAND U792 ( .A(n629), .B(n628), .Z(n630) );
  NAND U793 ( .A(n631), .B(n630), .Z(n632) );
  XOR U794 ( .A(n633), .B(n632), .Z(c[158]) );
  XOR U795 ( .A(a[159]), .B(b[159]), .Z(n637) );
  NAND U796 ( .A(a[158]), .B(b[158]), .Z(n635) );
  NAND U797 ( .A(n633), .B(n632), .Z(n634) );
  NAND U798 ( .A(n635), .B(n634), .Z(n636) );
  XOR U799 ( .A(n637), .B(n636), .Z(c[159]) );
  XOR U800 ( .A(a[160]), .B(b[160]), .Z(n641) );
  NAND U801 ( .A(a[159]), .B(b[159]), .Z(n639) );
  NAND U802 ( .A(n637), .B(n636), .Z(n638) );
  NAND U803 ( .A(n639), .B(n638), .Z(n640) );
  XOR U804 ( .A(n641), .B(n640), .Z(c[160]) );
  XOR U805 ( .A(a[161]), .B(b[161]), .Z(n645) );
  NAND U806 ( .A(a[160]), .B(b[160]), .Z(n643) );
  NAND U807 ( .A(n641), .B(n640), .Z(n642) );
  NAND U808 ( .A(n643), .B(n642), .Z(n644) );
  XOR U809 ( .A(n645), .B(n644), .Z(c[161]) );
  XOR U810 ( .A(a[162]), .B(b[162]), .Z(n649) );
  NAND U811 ( .A(a[161]), .B(b[161]), .Z(n647) );
  NAND U812 ( .A(n645), .B(n644), .Z(n646) );
  NAND U813 ( .A(n647), .B(n646), .Z(n648) );
  XOR U814 ( .A(n649), .B(n648), .Z(c[162]) );
  XOR U815 ( .A(a[163]), .B(b[163]), .Z(n653) );
  NAND U816 ( .A(a[162]), .B(b[162]), .Z(n651) );
  NAND U817 ( .A(n649), .B(n648), .Z(n650) );
  NAND U818 ( .A(n651), .B(n650), .Z(n652) );
  XOR U819 ( .A(n653), .B(n652), .Z(c[163]) );
  XOR U820 ( .A(a[164]), .B(b[164]), .Z(n657) );
  NAND U821 ( .A(a[163]), .B(b[163]), .Z(n655) );
  NAND U822 ( .A(n653), .B(n652), .Z(n654) );
  NAND U823 ( .A(n655), .B(n654), .Z(n656) );
  XOR U824 ( .A(n657), .B(n656), .Z(c[164]) );
  XOR U825 ( .A(a[165]), .B(b[165]), .Z(n661) );
  NAND U826 ( .A(a[164]), .B(b[164]), .Z(n659) );
  NAND U827 ( .A(n657), .B(n656), .Z(n658) );
  NAND U828 ( .A(n659), .B(n658), .Z(n660) );
  XOR U829 ( .A(n661), .B(n660), .Z(c[165]) );
  XOR U830 ( .A(a[166]), .B(b[166]), .Z(n665) );
  NAND U831 ( .A(a[165]), .B(b[165]), .Z(n663) );
  NAND U832 ( .A(n661), .B(n660), .Z(n662) );
  NAND U833 ( .A(n663), .B(n662), .Z(n664) );
  XOR U834 ( .A(n665), .B(n664), .Z(c[166]) );
  XOR U835 ( .A(a[167]), .B(b[167]), .Z(n669) );
  NAND U836 ( .A(a[166]), .B(b[166]), .Z(n667) );
  NAND U837 ( .A(n665), .B(n664), .Z(n666) );
  NAND U838 ( .A(n667), .B(n666), .Z(n668) );
  XOR U839 ( .A(n669), .B(n668), .Z(c[167]) );
  XOR U840 ( .A(a[168]), .B(b[168]), .Z(n673) );
  NAND U841 ( .A(a[167]), .B(b[167]), .Z(n671) );
  NAND U842 ( .A(n669), .B(n668), .Z(n670) );
  NAND U843 ( .A(n671), .B(n670), .Z(n672) );
  XOR U844 ( .A(n673), .B(n672), .Z(c[168]) );
  XOR U845 ( .A(a[169]), .B(b[169]), .Z(n677) );
  NAND U846 ( .A(a[168]), .B(b[168]), .Z(n675) );
  NAND U847 ( .A(n673), .B(n672), .Z(n674) );
  NAND U848 ( .A(n675), .B(n674), .Z(n676) );
  XOR U849 ( .A(n677), .B(n676), .Z(c[169]) );
  XOR U850 ( .A(a[170]), .B(b[170]), .Z(n681) );
  NAND U851 ( .A(a[169]), .B(b[169]), .Z(n679) );
  NAND U852 ( .A(n677), .B(n676), .Z(n678) );
  NAND U853 ( .A(n679), .B(n678), .Z(n680) );
  XOR U854 ( .A(n681), .B(n680), .Z(c[170]) );
  XOR U855 ( .A(a[171]), .B(b[171]), .Z(n685) );
  NAND U856 ( .A(a[170]), .B(b[170]), .Z(n683) );
  NAND U857 ( .A(n681), .B(n680), .Z(n682) );
  NAND U858 ( .A(n683), .B(n682), .Z(n684) );
  XOR U859 ( .A(n685), .B(n684), .Z(c[171]) );
  XOR U860 ( .A(a[172]), .B(b[172]), .Z(n689) );
  NAND U861 ( .A(a[171]), .B(b[171]), .Z(n687) );
  NAND U862 ( .A(n685), .B(n684), .Z(n686) );
  NAND U863 ( .A(n687), .B(n686), .Z(n688) );
  XOR U864 ( .A(n689), .B(n688), .Z(c[172]) );
  XOR U865 ( .A(a[173]), .B(b[173]), .Z(n693) );
  NAND U866 ( .A(a[172]), .B(b[172]), .Z(n691) );
  NAND U867 ( .A(n689), .B(n688), .Z(n690) );
  NAND U868 ( .A(n691), .B(n690), .Z(n692) );
  XOR U869 ( .A(n693), .B(n692), .Z(c[173]) );
  XOR U870 ( .A(a[174]), .B(b[174]), .Z(n697) );
  NAND U871 ( .A(a[173]), .B(b[173]), .Z(n695) );
  NAND U872 ( .A(n693), .B(n692), .Z(n694) );
  NAND U873 ( .A(n695), .B(n694), .Z(n696) );
  XOR U874 ( .A(n697), .B(n696), .Z(c[174]) );
  XOR U875 ( .A(a[175]), .B(b[175]), .Z(n701) );
  NAND U876 ( .A(a[174]), .B(b[174]), .Z(n699) );
  NAND U877 ( .A(n697), .B(n696), .Z(n698) );
  NAND U878 ( .A(n699), .B(n698), .Z(n700) );
  XOR U879 ( .A(n701), .B(n700), .Z(c[175]) );
  XOR U880 ( .A(a[176]), .B(b[176]), .Z(n705) );
  NAND U881 ( .A(a[175]), .B(b[175]), .Z(n703) );
  NAND U882 ( .A(n701), .B(n700), .Z(n702) );
  NAND U883 ( .A(n703), .B(n702), .Z(n704) );
  XOR U884 ( .A(n705), .B(n704), .Z(c[176]) );
  XOR U885 ( .A(a[177]), .B(b[177]), .Z(n709) );
  NAND U886 ( .A(a[176]), .B(b[176]), .Z(n707) );
  NAND U887 ( .A(n705), .B(n704), .Z(n706) );
  NAND U888 ( .A(n707), .B(n706), .Z(n708) );
  XOR U889 ( .A(n709), .B(n708), .Z(c[177]) );
  XOR U890 ( .A(a[178]), .B(b[178]), .Z(n713) );
  NAND U891 ( .A(a[177]), .B(b[177]), .Z(n711) );
  NAND U892 ( .A(n709), .B(n708), .Z(n710) );
  NAND U893 ( .A(n711), .B(n710), .Z(n712) );
  XOR U894 ( .A(n713), .B(n712), .Z(c[178]) );
  XOR U895 ( .A(a[179]), .B(b[179]), .Z(n717) );
  NAND U896 ( .A(a[178]), .B(b[178]), .Z(n715) );
  NAND U897 ( .A(n713), .B(n712), .Z(n714) );
  NAND U898 ( .A(n715), .B(n714), .Z(n716) );
  XOR U899 ( .A(n717), .B(n716), .Z(c[179]) );
  XOR U900 ( .A(a[180]), .B(b[180]), .Z(n721) );
  NAND U901 ( .A(a[179]), .B(b[179]), .Z(n719) );
  NAND U902 ( .A(n717), .B(n716), .Z(n718) );
  NAND U903 ( .A(n719), .B(n718), .Z(n720) );
  XOR U904 ( .A(n721), .B(n720), .Z(c[180]) );
  XOR U905 ( .A(a[181]), .B(b[181]), .Z(n725) );
  NAND U906 ( .A(a[180]), .B(b[180]), .Z(n723) );
  NAND U907 ( .A(n721), .B(n720), .Z(n722) );
  NAND U908 ( .A(n723), .B(n722), .Z(n724) );
  XOR U909 ( .A(n725), .B(n724), .Z(c[181]) );
  XOR U910 ( .A(a[182]), .B(b[182]), .Z(n729) );
  NAND U911 ( .A(a[181]), .B(b[181]), .Z(n727) );
  NAND U912 ( .A(n725), .B(n724), .Z(n726) );
  NAND U913 ( .A(n727), .B(n726), .Z(n728) );
  XOR U914 ( .A(n729), .B(n728), .Z(c[182]) );
  XOR U915 ( .A(a[183]), .B(b[183]), .Z(n733) );
  NAND U916 ( .A(a[182]), .B(b[182]), .Z(n731) );
  NAND U917 ( .A(n729), .B(n728), .Z(n730) );
  NAND U918 ( .A(n731), .B(n730), .Z(n732) );
  XOR U919 ( .A(n733), .B(n732), .Z(c[183]) );
  XOR U920 ( .A(a[184]), .B(b[184]), .Z(n737) );
  NAND U921 ( .A(a[183]), .B(b[183]), .Z(n735) );
  NAND U922 ( .A(n733), .B(n732), .Z(n734) );
  NAND U923 ( .A(n735), .B(n734), .Z(n736) );
  XOR U924 ( .A(n737), .B(n736), .Z(c[184]) );
  XOR U925 ( .A(a[185]), .B(b[185]), .Z(n741) );
  NAND U926 ( .A(a[184]), .B(b[184]), .Z(n739) );
  NAND U927 ( .A(n737), .B(n736), .Z(n738) );
  NAND U928 ( .A(n739), .B(n738), .Z(n740) );
  XOR U929 ( .A(n741), .B(n740), .Z(c[185]) );
  XOR U930 ( .A(a[186]), .B(b[186]), .Z(n745) );
  NAND U931 ( .A(a[185]), .B(b[185]), .Z(n743) );
  NAND U932 ( .A(n741), .B(n740), .Z(n742) );
  NAND U933 ( .A(n743), .B(n742), .Z(n744) );
  XOR U934 ( .A(n745), .B(n744), .Z(c[186]) );
  XOR U935 ( .A(a[187]), .B(b[187]), .Z(n749) );
  NAND U936 ( .A(a[186]), .B(b[186]), .Z(n747) );
  NAND U937 ( .A(n745), .B(n744), .Z(n746) );
  NAND U938 ( .A(n747), .B(n746), .Z(n748) );
  XOR U939 ( .A(n749), .B(n748), .Z(c[187]) );
  XOR U940 ( .A(a[188]), .B(b[188]), .Z(n753) );
  NAND U941 ( .A(a[187]), .B(b[187]), .Z(n751) );
  NAND U942 ( .A(n749), .B(n748), .Z(n750) );
  NAND U943 ( .A(n751), .B(n750), .Z(n752) );
  XOR U944 ( .A(n753), .B(n752), .Z(c[188]) );
  XOR U945 ( .A(a[189]), .B(b[189]), .Z(n757) );
  NAND U946 ( .A(a[188]), .B(b[188]), .Z(n755) );
  NAND U947 ( .A(n753), .B(n752), .Z(n754) );
  NAND U948 ( .A(n755), .B(n754), .Z(n756) );
  XOR U949 ( .A(n757), .B(n756), .Z(c[189]) );
  XOR U950 ( .A(a[190]), .B(b[190]), .Z(n761) );
  NAND U951 ( .A(a[189]), .B(b[189]), .Z(n759) );
  NAND U952 ( .A(n757), .B(n756), .Z(n758) );
  NAND U953 ( .A(n759), .B(n758), .Z(n760) );
  XOR U954 ( .A(n761), .B(n760), .Z(c[190]) );
  XOR U955 ( .A(a[191]), .B(b[191]), .Z(n765) );
  NAND U956 ( .A(a[190]), .B(b[190]), .Z(n763) );
  NAND U957 ( .A(n761), .B(n760), .Z(n762) );
  NAND U958 ( .A(n763), .B(n762), .Z(n764) );
  XOR U959 ( .A(n765), .B(n764), .Z(c[191]) );
  XOR U960 ( .A(a[192]), .B(b[192]), .Z(n769) );
  NAND U961 ( .A(a[191]), .B(b[191]), .Z(n767) );
  NAND U962 ( .A(n765), .B(n764), .Z(n766) );
  NAND U963 ( .A(n767), .B(n766), .Z(n768) );
  XOR U964 ( .A(n769), .B(n768), .Z(c[192]) );
  XOR U965 ( .A(a[193]), .B(b[193]), .Z(n773) );
  NAND U966 ( .A(a[192]), .B(b[192]), .Z(n771) );
  NAND U967 ( .A(n769), .B(n768), .Z(n770) );
  NAND U968 ( .A(n771), .B(n770), .Z(n772) );
  XOR U969 ( .A(n773), .B(n772), .Z(c[193]) );
  XOR U970 ( .A(a[194]), .B(b[194]), .Z(n777) );
  NAND U971 ( .A(a[193]), .B(b[193]), .Z(n775) );
  NAND U972 ( .A(n773), .B(n772), .Z(n774) );
  NAND U973 ( .A(n775), .B(n774), .Z(n776) );
  XOR U974 ( .A(n777), .B(n776), .Z(c[194]) );
  XOR U975 ( .A(a[195]), .B(b[195]), .Z(n781) );
  NAND U976 ( .A(a[194]), .B(b[194]), .Z(n779) );
  NAND U977 ( .A(n777), .B(n776), .Z(n778) );
  NAND U978 ( .A(n779), .B(n778), .Z(n780) );
  XOR U979 ( .A(n781), .B(n780), .Z(c[195]) );
  XOR U980 ( .A(a[196]), .B(b[196]), .Z(n785) );
  NAND U981 ( .A(a[195]), .B(b[195]), .Z(n783) );
  NAND U982 ( .A(n781), .B(n780), .Z(n782) );
  NAND U983 ( .A(n783), .B(n782), .Z(n784) );
  XOR U984 ( .A(n785), .B(n784), .Z(c[196]) );
  XOR U985 ( .A(a[197]), .B(b[197]), .Z(n789) );
  NAND U986 ( .A(a[196]), .B(b[196]), .Z(n787) );
  NAND U987 ( .A(n785), .B(n784), .Z(n786) );
  NAND U988 ( .A(n787), .B(n786), .Z(n788) );
  XOR U989 ( .A(n789), .B(n788), .Z(c[197]) );
  XOR U990 ( .A(a[198]), .B(b[198]), .Z(n793) );
  NAND U991 ( .A(a[197]), .B(b[197]), .Z(n791) );
  NAND U992 ( .A(n789), .B(n788), .Z(n790) );
  NAND U993 ( .A(n791), .B(n790), .Z(n792) );
  XOR U994 ( .A(n793), .B(n792), .Z(c[198]) );
  XOR U995 ( .A(a[199]), .B(b[199]), .Z(n797) );
  NAND U996 ( .A(a[198]), .B(b[198]), .Z(n795) );
  NAND U997 ( .A(n793), .B(n792), .Z(n794) );
  NAND U998 ( .A(n795), .B(n794), .Z(n796) );
  XOR U999 ( .A(n797), .B(n796), .Z(c[199]) );
  XOR U1000 ( .A(a[200]), .B(b[200]), .Z(n801) );
  NAND U1001 ( .A(a[199]), .B(b[199]), .Z(n799) );
  NAND U1002 ( .A(n797), .B(n796), .Z(n798) );
  NAND U1003 ( .A(n799), .B(n798), .Z(n800) );
  XOR U1004 ( .A(n801), .B(n800), .Z(c[200]) );
  XOR U1005 ( .A(a[201]), .B(b[201]), .Z(n805) );
  NAND U1006 ( .A(a[200]), .B(b[200]), .Z(n803) );
  NAND U1007 ( .A(n801), .B(n800), .Z(n802) );
  NAND U1008 ( .A(n803), .B(n802), .Z(n804) );
  XOR U1009 ( .A(n805), .B(n804), .Z(c[201]) );
  XOR U1010 ( .A(a[202]), .B(b[202]), .Z(n809) );
  NAND U1011 ( .A(a[201]), .B(b[201]), .Z(n807) );
  NAND U1012 ( .A(n805), .B(n804), .Z(n806) );
  NAND U1013 ( .A(n807), .B(n806), .Z(n808) );
  XOR U1014 ( .A(n809), .B(n808), .Z(c[202]) );
  XOR U1015 ( .A(a[203]), .B(b[203]), .Z(n813) );
  NAND U1016 ( .A(a[202]), .B(b[202]), .Z(n811) );
  NAND U1017 ( .A(n809), .B(n808), .Z(n810) );
  NAND U1018 ( .A(n811), .B(n810), .Z(n812) );
  XOR U1019 ( .A(n813), .B(n812), .Z(c[203]) );
  XOR U1020 ( .A(a[204]), .B(b[204]), .Z(n817) );
  NAND U1021 ( .A(a[203]), .B(b[203]), .Z(n815) );
  NAND U1022 ( .A(n813), .B(n812), .Z(n814) );
  NAND U1023 ( .A(n815), .B(n814), .Z(n816) );
  XOR U1024 ( .A(n817), .B(n816), .Z(c[204]) );
  XOR U1025 ( .A(a[205]), .B(b[205]), .Z(n821) );
  NAND U1026 ( .A(a[204]), .B(b[204]), .Z(n819) );
  NAND U1027 ( .A(n817), .B(n816), .Z(n818) );
  NAND U1028 ( .A(n819), .B(n818), .Z(n820) );
  XOR U1029 ( .A(n821), .B(n820), .Z(c[205]) );
  XOR U1030 ( .A(a[206]), .B(b[206]), .Z(n825) );
  NAND U1031 ( .A(a[205]), .B(b[205]), .Z(n823) );
  NAND U1032 ( .A(n821), .B(n820), .Z(n822) );
  NAND U1033 ( .A(n823), .B(n822), .Z(n824) );
  XOR U1034 ( .A(n825), .B(n824), .Z(c[206]) );
  XOR U1035 ( .A(a[207]), .B(b[207]), .Z(n829) );
  NAND U1036 ( .A(a[206]), .B(b[206]), .Z(n827) );
  NAND U1037 ( .A(n825), .B(n824), .Z(n826) );
  NAND U1038 ( .A(n827), .B(n826), .Z(n828) );
  XOR U1039 ( .A(n829), .B(n828), .Z(c[207]) );
  XOR U1040 ( .A(a[208]), .B(b[208]), .Z(n833) );
  NAND U1041 ( .A(a[207]), .B(b[207]), .Z(n831) );
  NAND U1042 ( .A(n829), .B(n828), .Z(n830) );
  NAND U1043 ( .A(n831), .B(n830), .Z(n832) );
  XOR U1044 ( .A(n833), .B(n832), .Z(c[208]) );
  XOR U1045 ( .A(a[209]), .B(b[209]), .Z(n837) );
  NAND U1046 ( .A(a[208]), .B(b[208]), .Z(n835) );
  NAND U1047 ( .A(n833), .B(n832), .Z(n834) );
  NAND U1048 ( .A(n835), .B(n834), .Z(n836) );
  XOR U1049 ( .A(n837), .B(n836), .Z(c[209]) );
  XOR U1050 ( .A(a[210]), .B(b[210]), .Z(n841) );
  NAND U1051 ( .A(a[209]), .B(b[209]), .Z(n839) );
  NAND U1052 ( .A(n837), .B(n836), .Z(n838) );
  NAND U1053 ( .A(n839), .B(n838), .Z(n840) );
  XOR U1054 ( .A(n841), .B(n840), .Z(c[210]) );
  XOR U1055 ( .A(a[211]), .B(b[211]), .Z(n845) );
  NAND U1056 ( .A(a[210]), .B(b[210]), .Z(n843) );
  NAND U1057 ( .A(n841), .B(n840), .Z(n842) );
  NAND U1058 ( .A(n843), .B(n842), .Z(n844) );
  XOR U1059 ( .A(n845), .B(n844), .Z(c[211]) );
  XOR U1060 ( .A(a[212]), .B(b[212]), .Z(n849) );
  NAND U1061 ( .A(a[211]), .B(b[211]), .Z(n847) );
  NAND U1062 ( .A(n845), .B(n844), .Z(n846) );
  NAND U1063 ( .A(n847), .B(n846), .Z(n848) );
  XOR U1064 ( .A(n849), .B(n848), .Z(c[212]) );
  XOR U1065 ( .A(a[213]), .B(b[213]), .Z(n853) );
  NAND U1066 ( .A(a[212]), .B(b[212]), .Z(n851) );
  NAND U1067 ( .A(n849), .B(n848), .Z(n850) );
  NAND U1068 ( .A(n851), .B(n850), .Z(n852) );
  XOR U1069 ( .A(n853), .B(n852), .Z(c[213]) );
  XOR U1070 ( .A(a[214]), .B(b[214]), .Z(n857) );
  NAND U1071 ( .A(a[213]), .B(b[213]), .Z(n855) );
  NAND U1072 ( .A(n853), .B(n852), .Z(n854) );
  NAND U1073 ( .A(n855), .B(n854), .Z(n856) );
  XOR U1074 ( .A(n857), .B(n856), .Z(c[214]) );
  XOR U1075 ( .A(a[215]), .B(b[215]), .Z(n861) );
  NAND U1076 ( .A(a[214]), .B(b[214]), .Z(n859) );
  NAND U1077 ( .A(n857), .B(n856), .Z(n858) );
  NAND U1078 ( .A(n859), .B(n858), .Z(n860) );
  XOR U1079 ( .A(n861), .B(n860), .Z(c[215]) );
  XOR U1080 ( .A(a[216]), .B(b[216]), .Z(n865) );
  NAND U1081 ( .A(a[215]), .B(b[215]), .Z(n863) );
  NAND U1082 ( .A(n861), .B(n860), .Z(n862) );
  NAND U1083 ( .A(n863), .B(n862), .Z(n864) );
  XOR U1084 ( .A(n865), .B(n864), .Z(c[216]) );
  XOR U1085 ( .A(a[217]), .B(b[217]), .Z(n869) );
  NAND U1086 ( .A(a[216]), .B(b[216]), .Z(n867) );
  NAND U1087 ( .A(n865), .B(n864), .Z(n866) );
  NAND U1088 ( .A(n867), .B(n866), .Z(n868) );
  XOR U1089 ( .A(n869), .B(n868), .Z(c[217]) );
  XOR U1090 ( .A(a[218]), .B(b[218]), .Z(n873) );
  NAND U1091 ( .A(a[217]), .B(b[217]), .Z(n871) );
  NAND U1092 ( .A(n869), .B(n868), .Z(n870) );
  NAND U1093 ( .A(n871), .B(n870), .Z(n872) );
  XOR U1094 ( .A(n873), .B(n872), .Z(c[218]) );
  XOR U1095 ( .A(a[219]), .B(b[219]), .Z(n877) );
  NAND U1096 ( .A(a[218]), .B(b[218]), .Z(n875) );
  NAND U1097 ( .A(n873), .B(n872), .Z(n874) );
  NAND U1098 ( .A(n875), .B(n874), .Z(n876) );
  XOR U1099 ( .A(n877), .B(n876), .Z(c[219]) );
  XOR U1100 ( .A(a[220]), .B(b[220]), .Z(n881) );
  NAND U1101 ( .A(a[219]), .B(b[219]), .Z(n879) );
  NAND U1102 ( .A(n877), .B(n876), .Z(n878) );
  NAND U1103 ( .A(n879), .B(n878), .Z(n880) );
  XOR U1104 ( .A(n881), .B(n880), .Z(c[220]) );
  XOR U1105 ( .A(a[221]), .B(b[221]), .Z(n885) );
  NAND U1106 ( .A(a[220]), .B(b[220]), .Z(n883) );
  NAND U1107 ( .A(n881), .B(n880), .Z(n882) );
  NAND U1108 ( .A(n883), .B(n882), .Z(n884) );
  XOR U1109 ( .A(n885), .B(n884), .Z(c[221]) );
  XOR U1110 ( .A(a[222]), .B(b[222]), .Z(n889) );
  NAND U1111 ( .A(a[221]), .B(b[221]), .Z(n887) );
  NAND U1112 ( .A(n885), .B(n884), .Z(n886) );
  NAND U1113 ( .A(n887), .B(n886), .Z(n888) );
  XOR U1114 ( .A(n889), .B(n888), .Z(c[222]) );
  XOR U1115 ( .A(a[223]), .B(b[223]), .Z(n893) );
  NAND U1116 ( .A(a[222]), .B(b[222]), .Z(n891) );
  NAND U1117 ( .A(n889), .B(n888), .Z(n890) );
  NAND U1118 ( .A(n891), .B(n890), .Z(n892) );
  XOR U1119 ( .A(n893), .B(n892), .Z(c[223]) );
  XOR U1120 ( .A(a[224]), .B(b[224]), .Z(n897) );
  NAND U1121 ( .A(a[223]), .B(b[223]), .Z(n895) );
  NAND U1122 ( .A(n893), .B(n892), .Z(n894) );
  NAND U1123 ( .A(n895), .B(n894), .Z(n896) );
  XOR U1124 ( .A(n897), .B(n896), .Z(c[224]) );
  XOR U1125 ( .A(a[225]), .B(b[225]), .Z(n901) );
  NAND U1126 ( .A(a[224]), .B(b[224]), .Z(n899) );
  NAND U1127 ( .A(n897), .B(n896), .Z(n898) );
  NAND U1128 ( .A(n899), .B(n898), .Z(n900) );
  XOR U1129 ( .A(n901), .B(n900), .Z(c[225]) );
  XOR U1130 ( .A(a[226]), .B(b[226]), .Z(n905) );
  NAND U1131 ( .A(a[225]), .B(b[225]), .Z(n903) );
  NAND U1132 ( .A(n901), .B(n900), .Z(n902) );
  NAND U1133 ( .A(n903), .B(n902), .Z(n904) );
  XOR U1134 ( .A(n905), .B(n904), .Z(c[226]) );
  XOR U1135 ( .A(a[227]), .B(b[227]), .Z(n909) );
  NAND U1136 ( .A(a[226]), .B(b[226]), .Z(n907) );
  NAND U1137 ( .A(n905), .B(n904), .Z(n906) );
  NAND U1138 ( .A(n907), .B(n906), .Z(n908) );
  XOR U1139 ( .A(n909), .B(n908), .Z(c[227]) );
  XOR U1140 ( .A(a[228]), .B(b[228]), .Z(n913) );
  NAND U1141 ( .A(a[227]), .B(b[227]), .Z(n911) );
  NAND U1142 ( .A(n909), .B(n908), .Z(n910) );
  NAND U1143 ( .A(n911), .B(n910), .Z(n912) );
  XOR U1144 ( .A(n913), .B(n912), .Z(c[228]) );
  XOR U1145 ( .A(a[229]), .B(b[229]), .Z(n917) );
  NAND U1146 ( .A(a[228]), .B(b[228]), .Z(n915) );
  NAND U1147 ( .A(n913), .B(n912), .Z(n914) );
  NAND U1148 ( .A(n915), .B(n914), .Z(n916) );
  XOR U1149 ( .A(n917), .B(n916), .Z(c[229]) );
  XOR U1150 ( .A(a[230]), .B(b[230]), .Z(n921) );
  NAND U1151 ( .A(a[229]), .B(b[229]), .Z(n919) );
  NAND U1152 ( .A(n917), .B(n916), .Z(n918) );
  NAND U1153 ( .A(n919), .B(n918), .Z(n920) );
  XOR U1154 ( .A(n921), .B(n920), .Z(c[230]) );
  XOR U1155 ( .A(a[231]), .B(b[231]), .Z(n925) );
  NAND U1156 ( .A(a[230]), .B(b[230]), .Z(n923) );
  NAND U1157 ( .A(n921), .B(n920), .Z(n922) );
  NAND U1158 ( .A(n923), .B(n922), .Z(n924) );
  XOR U1159 ( .A(n925), .B(n924), .Z(c[231]) );
  XOR U1160 ( .A(a[232]), .B(b[232]), .Z(n929) );
  NAND U1161 ( .A(a[231]), .B(b[231]), .Z(n927) );
  NAND U1162 ( .A(n925), .B(n924), .Z(n926) );
  NAND U1163 ( .A(n927), .B(n926), .Z(n928) );
  XOR U1164 ( .A(n929), .B(n928), .Z(c[232]) );
  XOR U1165 ( .A(a[233]), .B(b[233]), .Z(n933) );
  NAND U1166 ( .A(a[232]), .B(b[232]), .Z(n931) );
  NAND U1167 ( .A(n929), .B(n928), .Z(n930) );
  NAND U1168 ( .A(n931), .B(n930), .Z(n932) );
  XOR U1169 ( .A(n933), .B(n932), .Z(c[233]) );
  XOR U1170 ( .A(a[234]), .B(b[234]), .Z(n937) );
  NAND U1171 ( .A(a[233]), .B(b[233]), .Z(n935) );
  NAND U1172 ( .A(n933), .B(n932), .Z(n934) );
  NAND U1173 ( .A(n935), .B(n934), .Z(n936) );
  XOR U1174 ( .A(n937), .B(n936), .Z(c[234]) );
  XOR U1175 ( .A(a[235]), .B(b[235]), .Z(n941) );
  NAND U1176 ( .A(a[234]), .B(b[234]), .Z(n939) );
  NAND U1177 ( .A(n937), .B(n936), .Z(n938) );
  NAND U1178 ( .A(n939), .B(n938), .Z(n940) );
  XOR U1179 ( .A(n941), .B(n940), .Z(c[235]) );
  XOR U1180 ( .A(a[236]), .B(b[236]), .Z(n945) );
  NAND U1181 ( .A(a[235]), .B(b[235]), .Z(n943) );
  NAND U1182 ( .A(n941), .B(n940), .Z(n942) );
  NAND U1183 ( .A(n943), .B(n942), .Z(n944) );
  XOR U1184 ( .A(n945), .B(n944), .Z(c[236]) );
  XOR U1185 ( .A(a[237]), .B(b[237]), .Z(n949) );
  NAND U1186 ( .A(a[236]), .B(b[236]), .Z(n947) );
  NAND U1187 ( .A(n945), .B(n944), .Z(n946) );
  NAND U1188 ( .A(n947), .B(n946), .Z(n948) );
  XOR U1189 ( .A(n949), .B(n948), .Z(c[237]) );
  XOR U1190 ( .A(a[238]), .B(b[238]), .Z(n953) );
  NAND U1191 ( .A(a[237]), .B(b[237]), .Z(n951) );
  NAND U1192 ( .A(n949), .B(n948), .Z(n950) );
  NAND U1193 ( .A(n951), .B(n950), .Z(n952) );
  XOR U1194 ( .A(n953), .B(n952), .Z(c[238]) );
  XOR U1195 ( .A(a[239]), .B(b[239]), .Z(n957) );
  NAND U1196 ( .A(a[238]), .B(b[238]), .Z(n955) );
  NAND U1197 ( .A(n953), .B(n952), .Z(n954) );
  NAND U1198 ( .A(n955), .B(n954), .Z(n956) );
  XOR U1199 ( .A(n957), .B(n956), .Z(c[239]) );
  XOR U1200 ( .A(a[240]), .B(b[240]), .Z(n961) );
  NAND U1201 ( .A(a[239]), .B(b[239]), .Z(n959) );
  NAND U1202 ( .A(n957), .B(n956), .Z(n958) );
  NAND U1203 ( .A(n959), .B(n958), .Z(n960) );
  XOR U1204 ( .A(n961), .B(n960), .Z(c[240]) );
  XOR U1205 ( .A(a[241]), .B(b[241]), .Z(n965) );
  NAND U1206 ( .A(a[240]), .B(b[240]), .Z(n963) );
  NAND U1207 ( .A(n961), .B(n960), .Z(n962) );
  NAND U1208 ( .A(n963), .B(n962), .Z(n964) );
  XOR U1209 ( .A(n965), .B(n964), .Z(c[241]) );
  XOR U1210 ( .A(a[242]), .B(b[242]), .Z(n969) );
  NAND U1211 ( .A(a[241]), .B(b[241]), .Z(n967) );
  NAND U1212 ( .A(n965), .B(n964), .Z(n966) );
  NAND U1213 ( .A(n967), .B(n966), .Z(n968) );
  XOR U1214 ( .A(n969), .B(n968), .Z(c[242]) );
  XOR U1215 ( .A(a[243]), .B(b[243]), .Z(n973) );
  NAND U1216 ( .A(a[242]), .B(b[242]), .Z(n971) );
  NAND U1217 ( .A(n969), .B(n968), .Z(n970) );
  NAND U1218 ( .A(n971), .B(n970), .Z(n972) );
  XOR U1219 ( .A(n973), .B(n972), .Z(c[243]) );
  XOR U1220 ( .A(a[244]), .B(b[244]), .Z(n977) );
  NAND U1221 ( .A(a[243]), .B(b[243]), .Z(n975) );
  NAND U1222 ( .A(n973), .B(n972), .Z(n974) );
  NAND U1223 ( .A(n975), .B(n974), .Z(n976) );
  XOR U1224 ( .A(n977), .B(n976), .Z(c[244]) );
  XOR U1225 ( .A(a[245]), .B(b[245]), .Z(n981) );
  NAND U1226 ( .A(a[244]), .B(b[244]), .Z(n979) );
  NAND U1227 ( .A(n977), .B(n976), .Z(n978) );
  NAND U1228 ( .A(n979), .B(n978), .Z(n980) );
  XOR U1229 ( .A(n981), .B(n980), .Z(c[245]) );
  XOR U1230 ( .A(a[246]), .B(b[246]), .Z(n985) );
  NAND U1231 ( .A(a[245]), .B(b[245]), .Z(n983) );
  NAND U1232 ( .A(n981), .B(n980), .Z(n982) );
  NAND U1233 ( .A(n983), .B(n982), .Z(n984) );
  XOR U1234 ( .A(n985), .B(n984), .Z(c[246]) );
  XOR U1235 ( .A(a[247]), .B(b[247]), .Z(n989) );
  NAND U1236 ( .A(a[246]), .B(b[246]), .Z(n987) );
  NAND U1237 ( .A(n985), .B(n984), .Z(n986) );
  NAND U1238 ( .A(n987), .B(n986), .Z(n988) );
  XOR U1239 ( .A(n989), .B(n988), .Z(c[247]) );
  XOR U1240 ( .A(a[248]), .B(b[248]), .Z(n993) );
  NAND U1241 ( .A(a[247]), .B(b[247]), .Z(n991) );
  NAND U1242 ( .A(n989), .B(n988), .Z(n990) );
  NAND U1243 ( .A(n991), .B(n990), .Z(n992) );
  XOR U1244 ( .A(n993), .B(n992), .Z(c[248]) );
  XOR U1245 ( .A(a[249]), .B(b[249]), .Z(n997) );
  NAND U1246 ( .A(a[248]), .B(b[248]), .Z(n995) );
  NAND U1247 ( .A(n993), .B(n992), .Z(n994) );
  NAND U1248 ( .A(n995), .B(n994), .Z(n996) );
  XOR U1249 ( .A(n997), .B(n996), .Z(c[249]) );
  XOR U1250 ( .A(a[250]), .B(b[250]), .Z(n1001) );
  NAND U1251 ( .A(a[249]), .B(b[249]), .Z(n999) );
  NAND U1252 ( .A(n997), .B(n996), .Z(n998) );
  NAND U1253 ( .A(n999), .B(n998), .Z(n1000) );
  XOR U1254 ( .A(n1001), .B(n1000), .Z(c[250]) );
  XOR U1255 ( .A(a[251]), .B(b[251]), .Z(n1005) );
  NAND U1256 ( .A(a[250]), .B(b[250]), .Z(n1003) );
  NAND U1257 ( .A(n1001), .B(n1000), .Z(n1002) );
  NAND U1258 ( .A(n1003), .B(n1002), .Z(n1004) );
  XOR U1259 ( .A(n1005), .B(n1004), .Z(c[251]) );
  XOR U1260 ( .A(a[252]), .B(b[252]), .Z(n1009) );
  NAND U1261 ( .A(a[251]), .B(b[251]), .Z(n1007) );
  NAND U1262 ( .A(n1005), .B(n1004), .Z(n1006) );
  NAND U1263 ( .A(n1007), .B(n1006), .Z(n1008) );
  XOR U1264 ( .A(n1009), .B(n1008), .Z(c[252]) );
  XOR U1265 ( .A(a[253]), .B(b[253]), .Z(n1013) );
  NAND U1266 ( .A(a[252]), .B(b[252]), .Z(n1011) );
  NAND U1267 ( .A(n1009), .B(n1008), .Z(n1010) );
  NAND U1268 ( .A(n1011), .B(n1010), .Z(n1012) );
  XOR U1269 ( .A(n1013), .B(n1012), .Z(c[253]) );
  XOR U1270 ( .A(a[254]), .B(b[254]), .Z(n1017) );
  NAND U1271 ( .A(a[253]), .B(b[253]), .Z(n1015) );
  NAND U1272 ( .A(n1013), .B(n1012), .Z(n1014) );
  NAND U1273 ( .A(n1015), .B(n1014), .Z(n1016) );
  XOR U1274 ( .A(n1017), .B(n1016), .Z(c[254]) );
  NAND U1275 ( .A(a[254]), .B(b[254]), .Z(n1019) );
  NAND U1276 ( .A(n1017), .B(n1016), .Z(n1018) );
  AND U1277 ( .A(n1019), .B(n1018), .Z(n1021) );
  XOR U1278 ( .A(a[255]), .B(b[255]), .Z(n1020) );
  XNOR U1279 ( .A(n1021), .B(n1020), .Z(c[255]) );
  NAND U1280 ( .A(a[255]), .B(b[255]), .Z(n1023) );
  NANDN U1281 ( .A(n1021), .B(n1020), .Z(n1022) );
  NAND U1282 ( .A(n1023), .B(n1022), .Z(carry_on_d) );
endmodule

