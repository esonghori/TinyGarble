
module hamming_N160_CC16 ( clk, rst, x, y, o );
  input [9:0] x;
  input [9:0] y;
  output [7:0] o;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  wire   [7:0] oglobal;

  DFF \oglobal_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .Q(oglobal[7]) );
  DFF \oglobal_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .Q(oglobal[6]) );
  DFF \oglobal_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .Q(oglobal[5]) );
  DFF \oglobal_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .Q(oglobal[4]) );
  DFF \oglobal_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .Q(oglobal[3]) );
  DFF \oglobal_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .Q(oglobal[2]) );
  DFF \oglobal_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .Q(oglobal[1]) );
  DFF \oglobal_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .Q(oglobal[0]) );
  NAND U13 ( .A(n33), .B(n32), .Z(n1) );
  NANDN U14 ( .A(n34), .B(n35), .Z(n2) );
  NAND U15 ( .A(n1), .B(n2), .Z(n47) );
  XOR U16 ( .A(n44), .B(n45), .Z(n3) );
  NANDN U17 ( .A(n46), .B(n3), .Z(n4) );
  NAND U18 ( .A(n44), .B(n45), .Z(n5) );
  AND U19 ( .A(n4), .B(n5), .Z(n51) );
  NAND U20 ( .A(n13), .B(n11), .Z(n6) );
  XOR U21 ( .A(n13), .B(n11), .Z(n7) );
  NANDN U22 ( .A(n12), .B(n7), .Z(n8) );
  NAND U23 ( .A(n6), .B(n8), .Z(n39) );
  NANDN U24 ( .A(n56), .B(n57), .Z(n61) );
  NANDN U25 ( .A(n64), .B(oglobal[6]), .Z(n9) );
  XNOR U26 ( .A(oglobal[7]), .B(n9), .Z(o[7]) );
  XOR U27 ( .A(x[5]), .B(y[5]), .Z(n17) );
  XOR U28 ( .A(x[1]), .B(y[1]), .Z(n14) );
  XNOR U29 ( .A(x[3]), .B(y[3]), .Z(n15) );
  XNOR U30 ( .A(n14), .B(n15), .Z(n16) );
  XNOR U31 ( .A(n17), .B(n16), .Z(n13) );
  XOR U32 ( .A(x[9]), .B(y[9]), .Z(n20) );
  XNOR U33 ( .A(x[7]), .B(y[7]), .Z(n21) );
  XNOR U34 ( .A(n20), .B(n21), .Z(n23) );
  XOR U35 ( .A(x[4]), .B(y[4]), .Z(n35) );
  XOR U36 ( .A(x[8]), .B(y[8]), .Z(n33) );
  XOR U37 ( .A(x[6]), .B(y[6]), .Z(n32) );
  XNOR U38 ( .A(n33), .B(n32), .Z(n34) );
  XNOR U39 ( .A(n35), .B(n34), .Z(n22) );
  XNOR U40 ( .A(n23), .B(n22), .Z(n11) );
  XOR U41 ( .A(x[0]), .B(y[0]), .Z(n28) );
  XNOR U42 ( .A(x[2]), .B(y[2]), .Z(n26) );
  XNOR U43 ( .A(oglobal[0]), .B(n26), .Z(n27) );
  XOR U44 ( .A(n28), .B(n27), .Z(n12) );
  XNOR U45 ( .A(n11), .B(n12), .Z(n10) );
  XNOR U46 ( .A(n13), .B(n10), .Z(o[0]) );
  NANDN U47 ( .A(n15), .B(n14), .Z(n19) );
  NAND U48 ( .A(n17), .B(n16), .Z(n18) );
  NAND U49 ( .A(n19), .B(n18), .Z(n44) );
  NANDN U50 ( .A(n21), .B(n20), .Z(n25) );
  NAND U51 ( .A(n23), .B(n22), .Z(n24) );
  AND U52 ( .A(n25), .B(n24), .Z(n46) );
  NANDN U53 ( .A(n26), .B(oglobal[0]), .Z(n30) );
  NAND U54 ( .A(n28), .B(n27), .Z(n29) );
  NAND U55 ( .A(n30), .B(n29), .Z(n45) );
  XOR U56 ( .A(n46), .B(n45), .Z(n31) );
  XOR U57 ( .A(n44), .B(n31), .Z(n41) );
  XNOR U58 ( .A(oglobal[1]), .B(n47), .Z(n38) );
  IV U59 ( .A(n38), .Z(n37) );
  XNOR U60 ( .A(n41), .B(n37), .Z(n36) );
  XNOR U61 ( .A(n39), .B(n36), .Z(o[1]) );
  NANDN U62 ( .A(n39), .B(n37), .Z(n43) );
  AND U63 ( .A(n39), .B(n38), .Z(n40) );
  OR U64 ( .A(n41), .B(n40), .Z(n42) );
  AND U65 ( .A(n43), .B(n42), .Z(n49) );
  AND U66 ( .A(oglobal[1]), .B(n47), .Z(n54) );
  XOR U67 ( .A(n54), .B(oglobal[2]), .Z(n50) );
  XNOR U68 ( .A(n51), .B(n50), .Z(n48) );
  XNOR U69 ( .A(n49), .B(n48), .Z(o[2]) );
  NANDN U70 ( .A(n49), .B(n50), .Z(n53) );
  NANDN U71 ( .A(n50), .B(n49), .Z(n52) );
  ANDN U72 ( .B(n52), .A(n51), .Z(n57) );
  ANDN U73 ( .B(n53), .A(n57), .Z(n55) );
  NAND U74 ( .A(n54), .B(oglobal[2]), .Z(n56) );
  AND U75 ( .A(n55), .B(n56), .Z(n59) );
  NANDN U76 ( .A(n59), .B(n61), .Z(n58) );
  XNOR U77 ( .A(oglobal[3]), .B(n58), .Z(o[3]) );
  NANDN U78 ( .A(n59), .B(oglobal[3]), .Z(n60) );
  AND U79 ( .A(n61), .B(n60), .Z(n62) );
  XNOR U80 ( .A(n62), .B(oglobal[4]), .Z(o[4]) );
  ANDN U81 ( .B(oglobal[4]), .A(n62), .Z(n63) );
  XOR U82 ( .A(n63), .B(oglobal[5]), .Z(o[5]) );
  NAND U83 ( .A(n63), .B(oglobal[5]), .Z(n64) );
  XNOR U84 ( .A(oglobal[6]), .B(n64), .Z(o[6]) );
endmodule

